magic
tech sky130A
magscale 1 2
timestamp 1731260555
<< checkpaint >>
rect -3418 -3436 35750 26236
<< viali >>
rect 6193 21641 6227 21675
rect 6745 21641 6779 21675
rect 7297 21641 7331 21675
rect 7849 21641 7883 21675
rect 8401 21641 8435 21675
rect 9505 21641 9539 21675
rect 9781 21641 9815 21675
rect 10057 21641 10091 21675
rect 10609 21641 10643 21675
rect 11161 21641 11195 21675
rect 11621 21641 11655 21675
rect 11897 21641 11931 21675
rect 12265 21641 12299 21675
rect 12817 21641 12851 21675
rect 13369 21641 13403 21675
rect 13921 21641 13955 21675
rect 16313 21641 16347 21675
rect 20913 21641 20947 21675
rect 23121 21641 23155 21675
rect 25697 21641 25731 21675
rect 28825 21641 28859 21675
rect 20729 21573 20763 21607
rect 28181 21573 28215 21607
rect 14013 21505 14047 21539
rect 18429 21505 18463 21539
rect 18705 21505 18739 21539
rect 21281 21505 21315 21539
rect 25881 21505 25915 21539
rect 26433 21505 26467 21539
rect 29009 21505 29043 21539
rect 9413 21437 9447 21471
rect 16405 21437 16439 21471
rect 23121 21437 23155 21471
rect 23213 21437 23247 21471
rect 23949 21437 23983 21471
rect 31033 21437 31067 21471
rect 31309 21437 31343 21471
rect 11345 21369 11379 21403
rect 11437 21369 11471 21403
rect 14289 21369 14323 21403
rect 16681 21369 16715 21403
rect 18981 21369 19015 21403
rect 21097 21369 21131 21403
rect 21557 21369 21591 21403
rect 24225 21369 24259 21403
rect 26157 21369 26191 21403
rect 26709 21369 26743 21403
rect 28273 21369 28307 21403
rect 29285 21369 29319 21403
rect 8769 21301 8803 21335
rect 11637 21301 11671 21335
rect 11805 21301 11839 21335
rect 15761 21301 15795 21335
rect 20453 21301 20487 21335
rect 20897 21301 20931 21335
rect 23029 21301 23063 21335
rect 23489 21301 23523 21335
rect 28457 21301 28491 21335
rect 28549 21301 28583 21335
rect 28641 21301 28675 21335
rect 30757 21301 30791 21335
rect 30849 21301 30883 21335
rect 31217 21301 31251 21335
rect 10609 21097 10643 21131
rect 11069 21097 11103 21131
rect 11437 21097 11471 21131
rect 14289 21097 14323 21131
rect 16773 21097 16807 21131
rect 27169 21097 27203 21131
rect 28641 21097 28675 21131
rect 29377 21097 29411 21131
rect 31033 21097 31067 21131
rect 7757 21029 7791 21063
rect 8217 21029 8251 21063
rect 11805 21029 11839 21063
rect 18705 21029 18739 21063
rect 19073 21029 19107 21063
rect 27445 21029 27479 21063
rect 28917 21029 28951 21063
rect 29127 21029 29161 21063
rect 29863 21029 29897 21063
rect 30941 21029 30975 21063
rect 10793 20995 10827 21029
rect 7665 20961 7699 20995
rect 7849 20961 7883 20995
rect 10517 20961 10551 20995
rect 10609 20961 10643 20995
rect 10977 20961 11011 20995
rect 11253 20961 11287 20995
rect 13645 20961 13679 20995
rect 13829 20961 13863 20995
rect 14105 20961 14139 20995
rect 14841 20961 14875 20995
rect 15393 20961 15427 20995
rect 15761 20961 15795 20995
rect 16129 20961 16163 20995
rect 18613 20961 18647 20995
rect 19993 20961 20027 20995
rect 20637 20961 20671 20995
rect 20821 20961 20855 20995
rect 21281 20961 21315 20995
rect 21557 20961 21591 20995
rect 23489 20961 23523 20995
rect 23673 20961 23707 20995
rect 23949 20961 23983 20995
rect 24041 20961 24075 20995
rect 26249 20961 26283 20995
rect 26985 20961 27019 20995
rect 27353 20961 27387 20995
rect 27537 20961 27571 20995
rect 27655 20961 27689 20995
rect 28825 20961 28859 20995
rect 29009 20961 29043 20995
rect 29285 20961 29319 20995
rect 29561 20961 29595 20995
rect 29653 20961 29687 20995
rect 29745 20961 29779 20995
rect 7941 20893 7975 20927
rect 9689 20893 9723 20927
rect 11529 20893 11563 20927
rect 14565 20893 14599 20927
rect 15577 20893 15611 20927
rect 19349 20893 19383 20927
rect 20913 20893 20947 20927
rect 21097 20893 21131 20927
rect 21833 20893 21867 20927
rect 23305 20893 23339 20927
rect 24225 20893 24259 20927
rect 27813 20893 27847 20927
rect 27905 20893 27939 20927
rect 28457 20893 28491 20927
rect 30021 20893 30055 20927
rect 30757 20893 30791 20927
rect 17325 20825 17359 20859
rect 30113 20825 30147 20859
rect 13277 20757 13311 20791
rect 15117 20757 15151 20791
rect 15945 20757 15979 20791
rect 20085 20757 20119 20791
rect 21005 20757 21039 20791
rect 24961 20757 24995 20791
rect 26433 20757 26467 20791
rect 14197 20553 14231 20587
rect 14473 20553 14507 20587
rect 18705 20553 18739 20587
rect 18981 20553 19015 20587
rect 19441 20553 19475 20587
rect 23949 20553 23983 20587
rect 25973 20553 26007 20587
rect 28733 20553 28767 20587
rect 30757 20553 30791 20587
rect 7941 20485 7975 20519
rect 9229 20485 9263 20519
rect 20269 20485 20303 20519
rect 28549 20485 28583 20519
rect 30941 20485 30975 20519
rect 13921 20417 13955 20451
rect 16405 20417 16439 20451
rect 16497 20417 16531 20451
rect 16773 20417 16807 20451
rect 19349 20417 19383 20451
rect 22017 20417 22051 20451
rect 22937 20417 22971 20451
rect 24133 20417 24167 20451
rect 24409 20417 24443 20451
rect 25881 20417 25915 20451
rect 27077 20417 27111 20451
rect 27997 20417 28031 20451
rect 29009 20417 29043 20451
rect 7941 20349 7975 20383
rect 8217 20349 8251 20383
rect 8953 20349 8987 20383
rect 9045 20349 9079 20383
rect 9965 20349 9999 20383
rect 10333 20349 10367 20383
rect 10609 20349 10643 20383
rect 10977 20349 11011 20383
rect 13737 20349 13771 20383
rect 13829 20349 13863 20383
rect 14013 20349 14047 20383
rect 19165 20349 19199 20383
rect 19625 20349 19659 20383
rect 19993 20349 20027 20383
rect 22661 20349 22695 20383
rect 24041 20349 24075 20383
rect 26249 20349 26283 20383
rect 26341 20349 26375 20383
rect 26433 20349 26467 20383
rect 26617 20349 26651 20383
rect 26893 20349 26927 20383
rect 27353 20349 27387 20383
rect 27537 20349 27571 20383
rect 27655 20349 27689 20383
rect 27813 20349 27847 20383
rect 28641 20349 28675 20383
rect 28825 20349 28859 20383
rect 30849 20349 30883 20383
rect 31125 20349 31159 20383
rect 8125 20281 8159 20315
rect 9229 20281 9263 20315
rect 10149 20281 10183 20315
rect 11069 20281 11103 20315
rect 11621 20281 11655 20315
rect 13369 20281 13403 20315
rect 16129 20281 16163 20315
rect 18521 20281 18555 20315
rect 19717 20281 19751 20315
rect 19809 20281 19843 20315
rect 21741 20281 21775 20315
rect 23489 20281 23523 20315
rect 27446 20281 27480 20315
rect 29285 20281 29319 20315
rect 31309 20281 31343 20315
rect 9321 20213 9355 20247
rect 10517 20213 10551 20247
rect 10885 20213 10919 20247
rect 14657 20213 14691 20247
rect 22109 20213 22143 20247
rect 26709 20213 26743 20247
rect 27169 20213 27203 20247
rect 11513 20009 11547 20043
rect 12173 20009 12207 20043
rect 12449 20009 12483 20043
rect 13001 20009 13035 20043
rect 17049 20009 17083 20043
rect 17417 20009 17451 20043
rect 18629 20009 18663 20043
rect 19257 20009 19291 20043
rect 21439 20009 21473 20043
rect 21741 20009 21775 20043
rect 28365 20009 28399 20043
rect 29653 20009 29687 20043
rect 9321 19941 9355 19975
rect 11713 19941 11747 19975
rect 15577 19941 15611 19975
rect 15793 19941 15827 19975
rect 18429 19941 18463 19975
rect 18889 19941 18923 19975
rect 19089 19941 19123 19975
rect 19625 19941 19659 19975
rect 21649 19941 21683 19975
rect 29075 19941 29109 19975
rect 29193 19941 29227 19975
rect 30021 19941 30055 19975
rect 30159 19941 30193 19975
rect 7205 19873 7239 19907
rect 9045 19873 9079 19907
rect 11989 19873 12023 19907
rect 12081 19873 12115 19907
rect 12449 19873 12483 19907
rect 12621 19879 12655 19913
rect 12817 19873 12851 19907
rect 13461 19873 13495 19907
rect 13829 19873 13863 19907
rect 14289 19873 14323 19907
rect 15025 19873 15059 19907
rect 16497 19873 16531 19907
rect 17233 19873 17267 19907
rect 17509 19873 17543 19907
rect 17877 19873 17911 19907
rect 18061 19873 18095 19907
rect 18153 19873 18187 19907
rect 19349 19873 19383 19907
rect 23489 19873 23523 19907
rect 23581 19873 23615 19907
rect 26433 19873 26467 19907
rect 28549 19873 28583 19907
rect 28825 19873 28859 19907
rect 29284 19873 29318 19907
rect 29377 19873 29411 19907
rect 29837 19873 29871 19907
rect 29929 19873 29963 19907
rect 30941 19873 30975 19907
rect 31125 19873 31159 19907
rect 31309 19873 31343 19907
rect 7481 19805 7515 19839
rect 10793 19805 10827 19839
rect 13737 19805 13771 19839
rect 13921 19805 13955 19839
rect 14381 19805 14415 19839
rect 16129 19805 16163 19839
rect 16313 19805 16347 19839
rect 16405 19805 16439 19839
rect 16589 19805 16623 19839
rect 17601 19805 17635 19839
rect 23213 19805 23247 19839
rect 23857 19805 23891 19839
rect 25421 19805 25455 19839
rect 25973 19805 26007 19839
rect 26709 19805 26743 19839
rect 28641 19805 28675 19839
rect 28917 19805 28951 19839
rect 30297 19805 30331 19839
rect 30389 19805 30423 19839
rect 11345 19737 11379 19771
rect 12311 19737 12345 19771
rect 13277 19737 13311 19771
rect 14197 19737 14231 19771
rect 15945 19737 15979 19771
rect 17785 19737 17819 19771
rect 18337 19737 18371 19771
rect 21281 19737 21315 19771
rect 25329 19737 25363 19771
rect 8953 19669 8987 19703
rect 11529 19669 11563 19703
rect 12817 19669 12851 19703
rect 13645 19669 13679 19703
rect 13921 19669 13955 19703
rect 15761 19669 15795 19703
rect 17693 19669 17727 19703
rect 18613 19669 18647 19703
rect 18797 19669 18831 19703
rect 19073 19669 19107 19703
rect 21097 19669 21131 19703
rect 21465 19669 21499 19703
rect 28181 19669 28215 19703
rect 28825 19669 28859 19703
rect 29561 19669 29595 19703
rect 31125 19669 31159 19703
rect 8401 19465 8435 19499
rect 8769 19465 8803 19499
rect 11989 19465 12023 19499
rect 13093 19465 13127 19499
rect 14197 19465 14231 19499
rect 16681 19465 16715 19499
rect 17141 19465 17175 19499
rect 17509 19465 17543 19499
rect 19165 19465 19199 19499
rect 21189 19465 21223 19499
rect 23857 19465 23891 19499
rect 25421 19465 25455 19499
rect 26801 19465 26835 19499
rect 21465 19397 21499 19431
rect 8861 19329 8895 19363
rect 26249 19329 26283 19363
rect 6469 19261 6503 19295
rect 8585 19261 8619 19295
rect 12173 19261 12207 19295
rect 12449 19261 12483 19295
rect 13093 19261 13127 19295
rect 13369 19261 13403 19295
rect 13553 19261 13587 19295
rect 13646 19261 13680 19295
rect 13829 19261 13863 19295
rect 14059 19261 14093 19295
rect 16313 19261 16347 19295
rect 16497 19261 16531 19295
rect 17325 19261 17359 19295
rect 17601 19261 17635 19295
rect 17693 19261 17727 19295
rect 20545 19261 20579 19295
rect 20729 19261 20763 19295
rect 20821 19261 20855 19295
rect 20913 19261 20947 19295
rect 21281 19261 21315 19295
rect 23673 19261 23707 19295
rect 24041 19261 24075 19295
rect 24317 19261 24351 19295
rect 24418 19261 24452 19295
rect 24869 19261 24903 19295
rect 25053 19261 25087 19295
rect 25145 19261 25179 19295
rect 25329 19261 25363 19295
rect 25605 19261 25639 19295
rect 25697 19261 25731 19295
rect 25789 19261 25823 19295
rect 25881 19261 25915 19295
rect 26341 19261 26375 19295
rect 26985 19261 27019 19295
rect 29009 19261 29043 19295
rect 13277 19193 13311 19227
rect 13921 19193 13955 19227
rect 18061 19193 18095 19227
rect 20453 19193 20487 19227
rect 21649 19193 21683 19227
rect 23397 19193 23431 19227
rect 26433 19193 26467 19227
rect 27261 19193 27295 19227
rect 29285 19193 29319 19227
rect 30849 19193 30883 19227
rect 31033 19193 31067 19227
rect 31217 19193 31251 19227
rect 6377 19125 6411 19159
rect 12357 19125 12391 19159
rect 24685 19125 24719 19159
rect 25329 19125 25363 19159
rect 28733 19125 28767 19159
rect 30757 19125 30791 19159
rect 8769 18921 8803 18955
rect 12173 18921 12207 18955
rect 13191 18921 13225 18955
rect 15669 18921 15703 18955
rect 16129 18921 16163 18955
rect 16681 18921 16715 18955
rect 19533 18921 19567 18955
rect 20177 18921 20211 18955
rect 21557 18921 21591 18955
rect 22293 18921 22327 18955
rect 25789 18921 25823 18955
rect 29377 18921 29411 18955
rect 29837 18921 29871 18955
rect 5181 18853 5215 18887
rect 6469 18853 6503 18887
rect 7665 18853 7699 18887
rect 10149 18853 10183 18887
rect 12817 18853 12851 18887
rect 13277 18853 13311 18887
rect 15577 18853 15611 18887
rect 16297 18853 16331 18887
rect 16497 18853 16531 18887
rect 17141 18853 17175 18887
rect 18981 18853 19015 18887
rect 19809 18853 19843 18887
rect 19993 18853 20027 18887
rect 26433 18853 26467 18887
rect 28825 18853 28859 18887
rect 29561 18853 29595 18887
rect 30481 18853 30515 18887
rect 3341 18785 3375 18819
rect 3525 18785 3559 18819
rect 3617 18785 3651 18819
rect 3801 18785 3835 18819
rect 3893 18785 3927 18819
rect 4445 18785 4479 18819
rect 5089 18785 5123 18819
rect 5273 18785 5307 18819
rect 5917 18785 5951 18819
rect 6193 18785 6227 18819
rect 6929 18785 6963 18819
rect 7481 18785 7515 18819
rect 8309 18785 8343 18819
rect 8401 18785 8435 18819
rect 8585 18785 8619 18819
rect 9045 18785 9079 18819
rect 9229 18785 9263 18819
rect 9321 18785 9355 18819
rect 9873 18785 9907 18819
rect 9965 18785 9999 18819
rect 10241 18785 10275 18819
rect 10333 18785 10367 18819
rect 11345 18785 11379 18819
rect 11529 18785 11563 18819
rect 13093 18785 13127 18819
rect 13369 18785 13403 18819
rect 16589 18785 16623 18819
rect 16773 18785 16807 18819
rect 20269 18785 20303 18819
rect 20729 18785 20763 18819
rect 22109 18785 22143 18819
rect 22753 18785 22787 18819
rect 24869 18785 24903 18819
rect 24961 18785 24995 18819
rect 25145 18785 25179 18819
rect 25329 18785 25363 18819
rect 25697 18785 25731 18819
rect 28549 18785 28583 18819
rect 29193 18785 29227 18819
rect 29745 18785 29779 18819
rect 30297 18785 30331 18819
rect 30665 18785 30699 18819
rect 30849 18785 30883 18819
rect 30941 18785 30975 18819
rect 31309 18785 31343 18819
rect 3985 18717 4019 18751
rect 6745 18717 6779 18751
rect 7205 18717 7239 18751
rect 12357 18717 12391 18751
rect 12449 18717 12483 18751
rect 15761 18717 15795 18751
rect 16865 18717 16899 18751
rect 19441 18717 19475 18751
rect 20545 18717 20579 18751
rect 22477 18717 22511 18751
rect 22569 18717 22603 18751
rect 22661 18717 22695 18751
rect 24593 18717 24627 18751
rect 25513 18717 25547 18751
rect 28273 18717 28307 18751
rect 30021 18717 30055 18751
rect 30113 18717 30147 18751
rect 30205 18717 30239 18751
rect 31033 18717 31067 18751
rect 3249 18649 3283 18683
rect 5917 18649 5951 18683
rect 8493 18649 8527 18683
rect 8861 18649 8895 18683
rect 18981 18649 19015 18683
rect 19717 18649 19751 18683
rect 20361 18649 20395 18683
rect 20453 18649 20487 18683
rect 28733 18649 28767 18683
rect 31125 18649 31159 18683
rect 3709 18581 3743 18615
rect 4353 18581 4387 18615
rect 6653 18581 6687 18615
rect 7113 18581 7147 18615
rect 7297 18581 7331 18615
rect 10517 18581 10551 18615
rect 11713 18581 11747 18615
rect 15209 18581 15243 18615
rect 16313 18581 16347 18615
rect 18613 18581 18647 18615
rect 21005 18581 21039 18615
rect 23121 18581 23155 18615
rect 26157 18581 26191 18615
rect 27721 18581 27755 18615
rect 28365 18581 28399 18615
rect 31217 18581 31251 18615
rect 2697 18377 2731 18411
rect 8769 18377 8803 18411
rect 11253 18377 11287 18411
rect 17049 18377 17083 18411
rect 19441 18377 19475 18411
rect 23305 18377 23339 18411
rect 27997 18377 28031 18411
rect 30849 18377 30883 18411
rect 31033 18377 31067 18411
rect 11437 18309 11471 18343
rect 18889 18309 18923 18343
rect 19533 18309 19567 18343
rect 23121 18309 23155 18343
rect 24317 18309 24351 18343
rect 30757 18309 30791 18343
rect 6745 18241 6779 18275
rect 14289 18241 14323 18275
rect 14657 18241 14691 18275
rect 14933 18241 14967 18275
rect 23029 18241 23063 18275
rect 24225 18241 24259 18275
rect 24685 18241 24719 18275
rect 27077 18241 27111 18275
rect 29009 18241 29043 18275
rect 2053 18173 2087 18207
rect 2605 18173 2639 18207
rect 3525 18173 3559 18207
rect 5641 18173 5675 18207
rect 6009 18173 6043 18207
rect 6193 18173 6227 18207
rect 6377 18173 6411 18207
rect 6653 18173 6687 18207
rect 8677 18173 8711 18207
rect 9781 18173 9815 18207
rect 10149 18173 10183 18207
rect 10241 18173 10275 18207
rect 11529 18173 11563 18207
rect 11897 18173 11931 18207
rect 13277 18173 13311 18207
rect 13737 18173 13771 18207
rect 13921 18173 13955 18207
rect 14013 18173 14047 18207
rect 14197 18173 14231 18207
rect 17233 18173 17267 18207
rect 17509 18173 17543 18207
rect 19073 18173 19107 18207
rect 19257 18173 19291 18207
rect 19717 18173 19751 18207
rect 20361 18173 20395 18207
rect 20545 18173 20579 18207
rect 20729 18173 20763 18207
rect 20913 18173 20947 18207
rect 21189 18173 21223 18207
rect 22569 18173 22603 18207
rect 22845 18173 22879 18207
rect 23949 18173 23983 18207
rect 24041 18173 24075 18207
rect 24501 18173 24535 18207
rect 27629 18173 27663 18207
rect 27721 18173 27755 18207
rect 27859 18173 27893 18207
rect 28181 18173 28215 18207
rect 28457 18173 28491 18207
rect 28641 18173 28675 18207
rect 1777 18105 1811 18139
rect 2421 18105 2455 18139
rect 6929 18105 6963 18139
rect 7297 18105 7331 18139
rect 7389 18105 7423 18139
rect 7573 18105 7607 18139
rect 10609 18105 10643 18139
rect 11069 18105 11103 18139
rect 11621 18105 11655 18139
rect 13093 18105 13127 18139
rect 16681 18105 16715 18139
rect 17417 18105 17451 18139
rect 20085 18105 20119 18139
rect 20453 18105 20487 18139
rect 21833 18105 21867 18139
rect 22385 18105 22419 18139
rect 23489 18105 23523 18139
rect 24869 18105 24903 18139
rect 26801 18105 26835 18139
rect 27353 18105 27387 18139
rect 28089 18105 28123 18139
rect 29285 18105 29319 18139
rect 31217 18105 31251 18139
rect 3341 18037 3375 18071
rect 9965 18037 9999 18071
rect 11269 18037 11303 18071
rect 11713 18037 11747 18071
rect 11897 18037 11931 18071
rect 13645 18037 13679 18071
rect 14289 18037 14323 18071
rect 19165 18037 19199 18071
rect 19809 18037 19843 18071
rect 19901 18037 19935 18071
rect 20177 18037 20211 18071
rect 21005 18037 21039 18071
rect 21373 18037 21407 18071
rect 21557 18037 21591 18071
rect 22109 18037 22143 18071
rect 22661 18037 22695 18071
rect 23289 18037 23323 18071
rect 25329 18037 25363 18071
rect 28365 18037 28399 18071
rect 31017 18037 31051 18071
rect 4353 17833 4387 17867
rect 5917 17833 5951 17867
rect 7389 17833 7423 17867
rect 7849 17833 7883 17867
rect 8953 17833 8987 17867
rect 9965 17833 9999 17867
rect 17417 17833 17451 17867
rect 21281 17833 21315 17867
rect 26249 17833 26283 17867
rect 2237 17765 2271 17799
rect 8585 17765 8619 17799
rect 17049 17765 17083 17799
rect 17249 17765 17283 17799
rect 18797 17765 18831 17799
rect 23397 17765 23431 17799
rect 25237 17765 25271 17799
rect 25467 17765 25501 17799
rect 25881 17765 25915 17799
rect 29745 17765 29779 17799
rect 18567 17731 18601 17765
rect 1501 17697 1535 17731
rect 2421 17697 2455 17731
rect 2605 17697 2639 17731
rect 2697 17697 2731 17731
rect 2806 17697 2840 17731
rect 3617 17697 3651 17731
rect 3893 17697 3927 17731
rect 4813 17697 4847 17731
rect 5825 17697 5859 17731
rect 6101 17697 6135 17731
rect 6745 17697 6779 17731
rect 7113 17697 7147 17731
rect 7205 17697 7239 17731
rect 8309 17697 8343 17731
rect 8429 17697 8463 17731
rect 8677 17697 8711 17731
rect 8815 17697 8849 17731
rect 9045 17697 9079 17731
rect 9229 17697 9263 17731
rect 9597 17697 9631 17731
rect 9781 17697 9815 17731
rect 10333 17697 10367 17731
rect 10517 17697 10551 17731
rect 10701 17697 10735 17731
rect 11621 17697 11655 17731
rect 11897 17697 11931 17731
rect 12725 17697 12759 17731
rect 12817 17697 12851 17731
rect 13001 17697 13035 17731
rect 13277 17697 13311 17731
rect 13737 17697 13771 17731
rect 14197 17697 14231 17731
rect 14289 17697 14323 17731
rect 14473 17697 14507 17731
rect 15669 17697 15703 17731
rect 17693 17697 17727 17731
rect 17785 17697 17819 17731
rect 18061 17697 18095 17731
rect 18337 17697 18371 17731
rect 20177 17697 20211 17731
rect 20269 17697 20303 17731
rect 20453 17697 20487 17731
rect 20611 17697 20645 17731
rect 20729 17697 20763 17731
rect 20821 17697 20855 17731
rect 20913 17697 20947 17731
rect 23029 17697 23063 17731
rect 23121 17697 23155 17731
rect 25145 17697 25179 17731
rect 25329 17697 25363 17731
rect 25717 17697 25751 17731
rect 25973 17697 26007 17731
rect 26065 17697 26099 17731
rect 28181 17697 28215 17731
rect 30021 17697 30055 17731
rect 30481 17697 30515 17731
rect 30757 17697 30791 17731
rect 1317 17629 1351 17663
rect 3341 17629 3375 17663
rect 4169 17629 4203 17663
rect 4261 17629 4295 17663
rect 4905 17629 4939 17663
rect 4997 17629 5031 17663
rect 6929 17629 6963 17663
rect 7021 17629 7055 17663
rect 7665 17629 7699 17663
rect 8033 17629 8067 17663
rect 9137 17629 9171 17663
rect 9505 17629 9539 17663
rect 9689 17629 9723 17663
rect 11713 17629 11747 17663
rect 12909 17629 12943 17663
rect 15301 17629 15335 17663
rect 15485 17629 15519 17663
rect 15577 17629 15611 17663
rect 15761 17629 15795 17663
rect 19993 17629 20027 17663
rect 21097 17629 21131 17663
rect 22753 17629 22787 17663
rect 25605 17629 25639 17663
rect 27905 17629 27939 17663
rect 3065 17561 3099 17595
rect 3985 17561 4019 17595
rect 4445 17561 4479 17595
rect 9321 17561 9355 17595
rect 17601 17561 17635 17595
rect 1685 17493 1719 17527
rect 2145 17493 2179 17527
rect 6285 17493 6319 17527
rect 8033 17493 8067 17527
rect 10241 17493 10275 17527
rect 10425 17493 10459 17527
rect 11897 17493 11931 17527
rect 12081 17493 12115 17527
rect 12541 17493 12575 17527
rect 13645 17493 13679 17527
rect 14013 17493 14047 17527
rect 14381 17493 14415 17527
rect 17233 17493 17267 17527
rect 18245 17493 18279 17527
rect 18429 17493 18463 17527
rect 18613 17493 18647 17527
rect 24869 17493 24903 17527
rect 24961 17493 24995 17527
rect 26433 17493 26467 17527
rect 28273 17493 28307 17527
rect 30205 17493 30239 17527
rect 30849 17493 30883 17527
rect 6929 17289 6963 17323
rect 8493 17289 8527 17323
rect 8769 17289 8803 17323
rect 11529 17289 11563 17323
rect 14749 17289 14783 17323
rect 15853 17289 15887 17323
rect 21465 17289 21499 17323
rect 22385 17289 22419 17323
rect 23489 17289 23523 17323
rect 26065 17289 26099 17323
rect 28273 17289 28307 17323
rect 31125 17289 31159 17323
rect 1501 17221 1535 17255
rect 4169 17221 4203 17255
rect 4261 17221 4295 17255
rect 13921 17221 13955 17255
rect 14197 17221 14231 17255
rect 18153 17221 18187 17255
rect 22753 17221 22787 17255
rect 4077 17153 4111 17187
rect 9781 17153 9815 17187
rect 12081 17153 12115 17187
rect 12173 17153 12207 17187
rect 16221 17153 16255 17187
rect 16313 17153 16347 17187
rect 22845 17153 22879 17187
rect 24317 17153 24351 17187
rect 24593 17153 24627 17187
rect 29377 17153 29411 17187
rect 1225 17085 1259 17119
rect 1501 17085 1535 17119
rect 1961 17085 1995 17119
rect 2054 17085 2088 17119
rect 2237 17085 2271 17119
rect 2426 17085 2460 17119
rect 3617 17085 3651 17119
rect 4353 17085 4387 17119
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 5365 17085 5399 17119
rect 5457 17085 5491 17119
rect 7113 17085 7147 17119
rect 7297 17085 7331 17119
rect 7389 17085 7423 17119
rect 8401 17085 8435 17119
rect 8585 17085 8619 17119
rect 10057 17085 10091 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 10517 17085 10551 17119
rect 11713 17085 11747 17119
rect 11805 17085 11839 17119
rect 14105 17085 14139 17119
rect 14289 17085 14323 17119
rect 14381 17085 14415 17119
rect 14565 17085 14599 17119
rect 14657 17085 14691 17119
rect 15025 17085 15059 17119
rect 16037 17085 16071 17119
rect 16129 17085 16163 17119
rect 17233 17085 17267 17119
rect 17417 17085 17451 17119
rect 19027 17085 19061 17119
rect 19165 17085 19199 17119
rect 19257 17085 19291 17119
rect 19440 17085 19474 17119
rect 19533 17085 19567 17119
rect 19901 17085 19935 17119
rect 19993 17085 20027 17119
rect 20177 17085 20211 17119
rect 20269 17085 20303 17119
rect 21373 17085 21407 17119
rect 21557 17085 21591 17119
rect 21925 17085 21959 17119
rect 22109 17085 22143 17119
rect 22569 17085 22603 17119
rect 22937 17085 22971 17119
rect 23029 17085 23063 17119
rect 23121 17085 23155 17119
rect 23857 17085 23891 17119
rect 24041 17085 24075 17119
rect 26433 17085 26467 17119
rect 26893 17085 26927 17119
rect 27077 17085 27111 17119
rect 27721 17085 27755 17119
rect 27905 17085 27939 17119
rect 28089 17085 28123 17119
rect 28365 17085 28399 17119
rect 29285 17085 29319 17119
rect 1317 17017 1351 17051
rect 2329 17017 2363 17051
rect 5181 17017 5215 17051
rect 10149 17017 10183 17051
rect 12817 17017 12851 17051
rect 13001 17017 13035 17051
rect 18521 17017 18555 17051
rect 23581 17017 23615 17051
rect 26157 17017 26191 17051
rect 27537 17017 27571 17051
rect 27997 17017 28031 17051
rect 28641 17017 28675 17051
rect 29653 17017 29687 17051
rect 2605 16949 2639 16983
rect 3341 16949 3375 16983
rect 4813 16949 4847 16983
rect 11989 16949 12023 16983
rect 13093 16949 13127 16983
rect 15209 16949 15243 16983
rect 17325 16949 17359 16983
rect 18061 16949 18095 16983
rect 18889 16949 18923 16983
rect 19717 16949 19751 16983
rect 21741 16949 21775 16983
rect 22201 16949 22235 16983
rect 24225 16949 24259 16983
rect 27445 16949 27479 16983
rect 29101 16949 29135 16983
rect 5457 16745 5491 16779
rect 5917 16745 5951 16779
rect 6561 16745 6595 16779
rect 11713 16745 11747 16779
rect 12357 16745 12391 16779
rect 12725 16745 12759 16779
rect 13369 16745 13403 16779
rect 15761 16745 15795 16779
rect 16681 16745 16715 16779
rect 17417 16745 17451 16779
rect 20729 16745 20763 16779
rect 25053 16745 25087 16779
rect 25881 16745 25915 16779
rect 27813 16745 27847 16779
rect 28825 16745 28859 16779
rect 8217 16677 8251 16711
rect 11529 16677 11563 16711
rect 21281 16677 21315 16711
rect 22753 16677 22787 16711
rect 23489 16677 23523 16711
rect 26709 16677 26743 16711
rect 27261 16677 27295 16711
rect 27629 16677 27663 16711
rect 27997 16677 28031 16711
rect 2789 16609 2823 16643
rect 2881 16609 2915 16643
rect 3157 16609 3191 16643
rect 4997 16609 5031 16643
rect 5273 16609 5307 16643
rect 6101 16609 6135 16643
rect 6285 16609 6319 16643
rect 6377 16609 6411 16643
rect 6745 16609 6779 16643
rect 6837 16609 6871 16643
rect 7021 16609 7055 16643
rect 7849 16609 7883 16643
rect 8033 16609 8067 16643
rect 8125 16609 8159 16643
rect 8401 16609 8435 16643
rect 9321 16609 9355 16643
rect 9413 16609 9447 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 11989 16609 12023 16643
rect 12541 16609 12575 16643
rect 12817 16609 12851 16643
rect 13553 16609 13587 16643
rect 13829 16609 13863 16643
rect 15945 16609 15979 16643
rect 16313 16609 16347 16643
rect 16405 16609 16439 16643
rect 16589 16609 16623 16643
rect 16681 16609 16715 16643
rect 16865 16609 16899 16643
rect 16957 16609 16991 16643
rect 17141 16609 17175 16643
rect 17509 16609 17543 16643
rect 17601 16609 17635 16643
rect 18705 16609 18739 16643
rect 18889 16609 18923 16643
rect 20545 16609 20579 16643
rect 20913 16609 20947 16643
rect 21557 16609 21591 16643
rect 22017 16609 22051 16643
rect 22109 16609 22143 16643
rect 22293 16609 22327 16643
rect 22385 16609 22419 16643
rect 22477 16609 22511 16643
rect 22845 16609 22879 16643
rect 23213 16609 23247 16643
rect 23673 16609 23707 16643
rect 23857 16609 23891 16643
rect 24225 16609 24259 16643
rect 24501 16609 24535 16643
rect 24685 16609 24719 16643
rect 24777 16609 24811 16643
rect 24961 16609 24995 16643
rect 25421 16609 25455 16643
rect 25697 16609 25731 16643
rect 26065 16609 26099 16643
rect 26249 16609 26283 16643
rect 26525 16609 26559 16643
rect 26801 16609 26835 16643
rect 26985 16609 27019 16643
rect 27721 16609 27755 16643
rect 28273 16609 28307 16643
rect 28549 16609 28583 16643
rect 28739 16609 28773 16643
rect 28917 16609 28951 16643
rect 29019 16609 29053 16643
rect 29745 16609 29779 16643
rect 29929 16609 29963 16643
rect 30389 16609 30423 16643
rect 30849 16609 30883 16643
rect 31125 16609 31159 16643
rect 3065 16541 3099 16575
rect 5089 16541 5123 16575
rect 5181 16541 5215 16575
rect 6929 16541 6963 16575
rect 11897 16541 11931 16575
rect 12081 16541 12115 16575
rect 12173 16541 12207 16575
rect 13645 16541 13679 16575
rect 13737 16541 13771 16575
rect 17233 16541 17267 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 24317 16541 24351 16575
rect 29285 16541 29319 16575
rect 16129 16473 16163 16507
rect 18705 16473 18739 16507
rect 24041 16473 24075 16507
rect 2973 16405 3007 16439
rect 16313 16405 16347 16439
rect 21097 16405 21131 16439
rect 26157 16405 26191 16439
rect 26893 16405 26927 16439
rect 28181 16405 28215 16439
rect 29653 16405 29687 16439
rect 31217 16405 31251 16439
rect 2605 16201 2639 16235
rect 3617 16201 3651 16235
rect 5089 16201 5123 16235
rect 6561 16201 6595 16235
rect 10149 16201 10183 16235
rect 11529 16201 11563 16235
rect 14289 16201 14323 16235
rect 14473 16201 14507 16235
rect 19441 16201 19475 16235
rect 19993 16201 20027 16235
rect 22109 16201 22143 16235
rect 22937 16201 22971 16235
rect 23121 16201 23155 16235
rect 26249 16201 26283 16235
rect 28273 16201 28307 16235
rect 29377 16201 29411 16235
rect 30757 16201 30791 16235
rect 9045 16133 9079 16167
rect 12081 16133 12115 16167
rect 22661 16133 22695 16167
rect 23949 16133 23983 16167
rect 25789 16133 25823 16167
rect 27813 16133 27847 16167
rect 29469 16133 29503 16167
rect 1225 16065 1259 16099
rect 1777 16065 1811 16099
rect 5273 16065 5307 16099
rect 7941 16065 7975 16099
rect 12725 16065 12759 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 19073 16065 19107 16099
rect 19901 16065 19935 16099
rect 21097 16065 21131 16099
rect 21281 16065 21315 16099
rect 21833 16065 21867 16099
rect 24317 16065 24351 16099
rect 24685 16065 24719 16099
rect 25145 16065 25179 16099
rect 29561 16065 29595 16099
rect 1409 15997 1443 16031
rect 1869 15997 1903 16031
rect 1961 15997 1995 16031
rect 2145 15997 2179 16031
rect 2237 15997 2271 16031
rect 2513 15997 2547 16031
rect 2697 15997 2731 16031
rect 3801 15997 3835 16031
rect 4261 15997 4295 16031
rect 4997 15997 5031 16031
rect 6469 15997 6503 16031
rect 6653 15997 6687 16031
rect 7757 15997 7791 16031
rect 7849 15997 7883 16031
rect 8033 15997 8067 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 8861 15997 8895 16031
rect 10333 15997 10367 16031
rect 10609 15997 10643 16031
rect 11713 15997 11747 16031
rect 11897 15997 11931 16031
rect 11989 15997 12023 16031
rect 12262 15997 12296 16031
rect 12633 15997 12667 16031
rect 13829 15997 13863 16031
rect 13921 15997 13955 16031
rect 14289 15997 14323 16031
rect 15301 15997 15335 16031
rect 15393 15997 15427 16031
rect 18889 15997 18923 16031
rect 19993 15997 20027 16031
rect 21373 15997 21407 16031
rect 21465 15997 21499 16031
rect 21557 15997 21591 16031
rect 21741 15997 21775 16031
rect 21925 15997 21959 16031
rect 22293 15997 22327 16031
rect 23397 15997 23431 16031
rect 24133 15997 24167 16031
rect 24501 15997 24535 16031
rect 24593 15997 24627 16031
rect 24777 15997 24811 16031
rect 25329 15997 25363 16031
rect 25789 15997 25823 16031
rect 26157 15997 26191 16031
rect 26341 15997 26375 16031
rect 26801 15997 26835 16031
rect 27261 15997 27295 16031
rect 27997 15997 28031 16031
rect 28089 15997 28123 16031
rect 28671 15997 28705 16031
rect 28825 15997 28859 16031
rect 29009 15997 29043 16031
rect 30389 15997 30423 16031
rect 30941 15997 30975 16031
rect 31125 15997 31159 16031
rect 5273 15929 5307 15963
rect 8677 15929 8711 15963
rect 8769 15929 8803 15963
rect 9505 15929 9539 15963
rect 13001 15929 13035 15963
rect 18705 15929 18739 15963
rect 19257 15929 19291 15963
rect 19457 15929 19491 15963
rect 19717 15929 19751 15963
rect 22385 15929 22419 15963
rect 23089 15929 23123 15963
rect 23305 15929 23339 15963
rect 28457 15929 28491 15963
rect 30205 15929 30239 15963
rect 1409 15861 1443 15895
rect 2421 15861 2455 15895
rect 8217 15861 8251 15895
rect 9597 15861 9631 15895
rect 10517 15861 10551 15895
rect 12265 15861 12299 15895
rect 12909 15861 12943 15895
rect 15117 15861 15151 15895
rect 15485 15861 15519 15895
rect 19625 15861 19659 15895
rect 22845 15861 22879 15895
rect 23581 15861 23615 15895
rect 26893 15861 26927 15895
rect 27445 15861 27479 15895
rect 29837 15861 29871 15895
rect 1593 15657 1627 15691
rect 3433 15657 3467 15691
rect 10701 15657 10735 15691
rect 12081 15657 12115 15691
rect 14013 15657 14047 15691
rect 15669 15657 15703 15691
rect 16313 15657 16347 15691
rect 22937 15657 22971 15691
rect 24685 15657 24719 15691
rect 27537 15657 27571 15691
rect 28457 15657 28491 15691
rect 29469 15657 29503 15691
rect 30941 15657 30975 15691
rect 5549 15589 5583 15623
rect 5917 15589 5951 15623
rect 8033 15589 8067 15623
rect 8401 15589 8435 15623
rect 14473 15589 14507 15623
rect 15025 15589 15059 15623
rect 21373 15589 21407 15623
rect 22477 15589 22511 15623
rect 23765 15589 23799 15623
rect 25860 15589 25894 15623
rect 26065 15589 26099 15623
rect 27077 15589 27111 15623
rect 28549 15589 28583 15623
rect 1501 15521 1535 15555
rect 1685 15521 1719 15555
rect 3157 15521 3191 15555
rect 3341 15521 3375 15555
rect 3801 15521 3835 15555
rect 5365 15521 5399 15555
rect 5641 15521 5675 15555
rect 6101 15521 6135 15555
rect 6285 15521 6319 15555
rect 6377 15521 6411 15555
rect 7481 15521 7515 15555
rect 7665 15521 7699 15555
rect 9321 15521 9355 15555
rect 10057 15521 10091 15555
rect 10241 15521 10275 15555
rect 10517 15521 10551 15555
rect 12081 15521 12115 15555
rect 12265 15521 12299 15555
rect 13277 15521 13311 15555
rect 13762 15521 13796 15555
rect 14841 15521 14875 15555
rect 15117 15521 15151 15555
rect 15209 15521 15243 15555
rect 15669 15521 15703 15555
rect 15853 15521 15887 15555
rect 16497 15521 16531 15555
rect 16589 15521 16623 15555
rect 16957 15521 16991 15555
rect 17969 15521 18003 15555
rect 18061 15521 18095 15555
rect 20913 15521 20947 15555
rect 21281 15521 21315 15555
rect 21465 15521 21499 15555
rect 23581 15521 23615 15555
rect 23673 15521 23707 15555
rect 23949 15521 23983 15555
rect 24041 15521 24075 15555
rect 24225 15521 24259 15555
rect 24317 15521 24351 15555
rect 24409 15521 24443 15555
rect 26985 15521 27019 15555
rect 27169 15521 27203 15555
rect 27353 15521 27387 15555
rect 27445 15521 27479 15555
rect 27721 15521 27755 15555
rect 27813 15521 27847 15555
rect 27997 15521 28031 15555
rect 28089 15521 28123 15555
rect 29009 15521 29043 15555
rect 29285 15521 29319 15555
rect 29561 15521 29595 15555
rect 29837 15521 29871 15555
rect 30757 15521 30791 15555
rect 31125 15521 31159 15555
rect 31309 15521 31343 15555
rect 3617 15453 3651 15487
rect 3709 15453 3743 15487
rect 3893 15453 3927 15487
rect 5181 15453 5215 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 9045 15453 9079 15487
rect 9137 15453 9171 15487
rect 9229 15453 9263 15487
rect 9505 15453 9539 15487
rect 10425 15453 10459 15487
rect 13553 15453 13587 15487
rect 16681 15453 16715 15487
rect 16773 15453 16807 15487
rect 17785 15453 17819 15487
rect 21097 15453 21131 15487
rect 23489 15453 23523 15487
rect 24777 15453 24811 15487
rect 25053 15453 25087 15487
rect 29984 15453 30018 15487
rect 30205 15453 30239 15487
rect 31217 15453 31251 15487
rect 7941 15385 7975 15419
rect 10333 15385 10367 15419
rect 20729 15385 20763 15419
rect 22845 15385 22879 15419
rect 25697 15385 25731 15419
rect 3157 15317 3191 15351
rect 13461 15317 13495 15351
rect 13645 15317 13679 15351
rect 14197 15317 14231 15351
rect 15393 15317 15427 15351
rect 17877 15317 17911 15351
rect 23949 15317 23983 15351
rect 25881 15317 25915 15351
rect 26801 15317 26835 15351
rect 28825 15317 28859 15351
rect 29101 15317 29135 15351
rect 30113 15317 30147 15351
rect 30297 15317 30331 15351
rect 5273 15113 5307 15147
rect 7297 15113 7331 15147
rect 7481 15113 7515 15147
rect 9597 15113 9631 15147
rect 11897 15113 11931 15147
rect 14657 15113 14691 15147
rect 14841 15113 14875 15147
rect 21925 15113 21959 15147
rect 29009 15113 29043 15147
rect 29469 15113 29503 15147
rect 29929 15113 29963 15147
rect 31033 15113 31067 15147
rect 3985 15045 4019 15079
rect 5641 15045 5675 15079
rect 6837 15045 6871 15079
rect 8033 15045 8067 15079
rect 9229 15045 9263 15079
rect 11529 15045 11563 15079
rect 24685 15045 24719 15079
rect 27997 15045 28031 15079
rect 5089 14977 5123 15011
rect 5825 14977 5859 15011
rect 7205 14977 7239 15011
rect 8861 14977 8895 15011
rect 9137 14977 9171 15011
rect 9505 14977 9539 15011
rect 14289 14977 14323 15011
rect 17693 14977 17727 15011
rect 17969 14977 18003 15011
rect 19717 14977 19751 15011
rect 20085 14977 20119 15011
rect 20729 14977 20763 15011
rect 20821 14977 20855 15011
rect 1501 14909 1535 14943
rect 1685 14909 1719 14943
rect 3341 14909 3375 14943
rect 3525 14909 3559 14943
rect 3617 14909 3651 14943
rect 3709 14909 3743 14943
rect 4077 14909 4111 14943
rect 4261 14909 4295 14943
rect 4905 14909 4939 14943
rect 5273 14909 5307 14943
rect 5549 14909 5583 14943
rect 5917 14909 5951 14943
rect 6101 14909 6135 14943
rect 7021 14909 7055 14943
rect 7389 14909 7423 14943
rect 7573 14909 7607 14943
rect 8217 14909 8251 14943
rect 8493 14909 8527 14943
rect 8677 14909 8711 14943
rect 8769 14909 8803 14943
rect 8953 14909 8987 14943
rect 9781 14909 9815 14943
rect 11253 14909 11287 14943
rect 11437 14909 11471 14943
rect 11621 14909 11655 14943
rect 11713 14909 11747 14943
rect 13553 14909 13587 14943
rect 13737 14909 13771 14943
rect 13829 14909 13863 14943
rect 13921 14909 13955 14943
rect 14105 14909 14139 14943
rect 17141 14909 17175 14943
rect 17233 14909 17267 14943
rect 17325 14909 17359 14943
rect 17509 14909 17543 14943
rect 17785 14909 17819 14943
rect 17877 14909 17911 14943
rect 19809 14909 19843 14943
rect 20637 14909 20671 14943
rect 20913 14909 20947 14943
rect 21373 14909 21407 14943
rect 21649 14909 21683 14943
rect 22109 14909 22143 14943
rect 22477 14909 22511 14943
rect 22569 14909 22603 14943
rect 23121 14909 23155 14943
rect 23397 14909 23431 14943
rect 24317 14909 24351 14943
rect 24501 14909 24535 14943
rect 24593 14909 24627 14943
rect 24777 14909 24811 14943
rect 26525 14909 26559 14943
rect 27905 14909 27939 14943
rect 28089 14909 28123 14943
rect 29285 14909 29319 14943
rect 29469 14909 29503 14943
rect 29745 14909 29779 14943
rect 30205 14909 30239 14943
rect 30573 14909 30607 14943
rect 30849 14909 30883 14943
rect 4169 14841 4203 14875
rect 6009 14841 6043 14875
rect 7297 14841 7331 14875
rect 14825 14841 14859 14875
rect 15025 14841 15059 14875
rect 20177 14841 20211 14875
rect 21281 14841 21315 14875
rect 22201 14841 22235 14875
rect 22293 14841 22327 14875
rect 23029 14841 23063 14875
rect 25513 14841 25547 14875
rect 25697 14841 25731 14875
rect 26065 14841 26099 14875
rect 29009 14841 29043 14875
rect 29561 14841 29595 14875
rect 30021 14841 30055 14875
rect 1593 14773 1627 14807
rect 4997 14773 5031 14807
rect 5825 14773 5859 14807
rect 16865 14773 16899 14807
rect 18153 14773 18187 14807
rect 19533 14773 19567 14807
rect 20453 14773 20487 14807
rect 24961 14773 24995 14807
rect 25789 14773 25823 14807
rect 25881 14773 25915 14807
rect 26249 14773 26283 14807
rect 29193 14773 29227 14807
rect 30389 14773 30423 14807
rect 30757 14773 30791 14807
rect 6377 14569 6411 14603
rect 7290 14569 7324 14603
rect 9321 14569 9355 14603
rect 14013 14569 14047 14603
rect 14841 14569 14875 14603
rect 16129 14569 16163 14603
rect 18061 14569 18095 14603
rect 22477 14569 22511 14603
rect 22937 14569 22971 14603
rect 29377 14569 29411 14603
rect 30665 14569 30699 14603
rect 3157 14501 3191 14535
rect 9137 14501 9171 14535
rect 12817 14501 12851 14535
rect 15209 14501 15243 14535
rect 25329 14501 25363 14535
rect 27077 14501 27111 14535
rect 28089 14501 28123 14535
rect 1685 14433 1719 14467
rect 1869 14433 1903 14467
rect 1961 14433 1995 14467
rect 2237 14433 2271 14467
rect 3433 14433 3467 14467
rect 5181 14433 5215 14467
rect 5457 14433 5491 14467
rect 6929 14433 6963 14467
rect 7113 14433 7147 14467
rect 7205 14433 7239 14467
rect 7389 14433 7423 14467
rect 7573 14433 7607 14467
rect 7757 14433 7791 14467
rect 8677 14433 8711 14467
rect 8861 14433 8895 14467
rect 9413 14433 9447 14467
rect 10609 14433 10643 14467
rect 10793 14433 10827 14467
rect 10977 14433 11011 14467
rect 11437 14433 11471 14467
rect 11713 14433 11747 14467
rect 11897 14433 11931 14467
rect 12725 14433 12759 14467
rect 13093 14433 13127 14467
rect 13369 14433 13403 14467
rect 13553 14433 13587 14467
rect 13645 14433 13679 14467
rect 13737 14433 13771 14467
rect 14749 14433 14783 14467
rect 15025 14433 15059 14467
rect 15301 14433 15335 14467
rect 15485 14433 15519 14467
rect 15577 14433 15611 14467
rect 15669 14433 15703 14467
rect 16313 14433 16347 14467
rect 16589 14433 16623 14467
rect 16773 14433 16807 14467
rect 18245 14433 18279 14467
rect 18429 14433 18463 14467
rect 18521 14433 18555 14467
rect 19533 14433 19567 14467
rect 19901 14433 19935 14467
rect 19993 14433 20027 14467
rect 22845 14433 22879 14467
rect 23121 14433 23155 14467
rect 23489 14433 23523 14467
rect 23857 14433 23891 14467
rect 24041 14433 24075 14467
rect 24133 14433 24167 14467
rect 24317 14433 24351 14467
rect 24409 14433 24443 14467
rect 24501 14433 24535 14467
rect 25697 14433 25731 14467
rect 25881 14433 25915 14467
rect 26985 14433 27019 14467
rect 27169 14433 27203 14467
rect 27353 14433 27387 14467
rect 27629 14433 27663 14467
rect 27905 14433 27939 14467
rect 28365 14433 28399 14467
rect 28733 14433 28767 14467
rect 28917 14433 28951 14467
rect 29377 14433 29411 14467
rect 29561 14433 29595 14467
rect 29837 14433 29871 14467
rect 30021 14433 30055 14467
rect 30205 14433 30239 14467
rect 30481 14433 30515 14467
rect 30757 14433 30791 14467
rect 30849 14433 30883 14467
rect 2053 14365 2087 14399
rect 3341 14365 3375 14399
rect 5273 14365 5307 14399
rect 5365 14365 5399 14399
rect 5641 14365 5675 14399
rect 5917 14365 5951 14399
rect 6009 14365 6043 14399
rect 6101 14365 6135 14399
rect 6193 14365 6227 14399
rect 11161 14365 11195 14399
rect 11253 14365 11287 14399
rect 11345 14365 11379 14399
rect 11805 14365 11839 14399
rect 12909 14365 12943 14399
rect 19349 14365 19383 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 19809 14365 19843 14399
rect 20177 14365 20211 14399
rect 22753 14365 22787 14399
rect 23949 14365 23983 14399
rect 27261 14365 27295 14399
rect 28089 14365 28123 14399
rect 29653 14365 29687 14399
rect 3617 14297 3651 14331
rect 7757 14297 7791 14331
rect 9045 14297 9079 14331
rect 9137 14297 9171 14331
rect 10793 14297 10827 14331
rect 13093 14297 13127 14331
rect 15945 14297 15979 14331
rect 16405 14297 16439 14331
rect 16497 14297 16531 14331
rect 20085 14297 20119 14331
rect 24961 14297 24995 14331
rect 2421 14229 2455 14263
rect 3157 14229 3191 14263
rect 6653 14229 6687 14263
rect 8677 14229 8711 14263
rect 11621 14229 11655 14263
rect 22845 14229 22879 14263
rect 23397 14229 23431 14263
rect 24777 14229 24811 14263
rect 24869 14229 24903 14263
rect 25697 14229 25731 14263
rect 27813 14229 27847 14263
rect 28273 14229 28307 14263
rect 28825 14229 28859 14263
rect 31033 14229 31067 14263
rect 3801 14025 3835 14059
rect 6837 14025 6871 14059
rect 8401 14025 8435 14059
rect 9413 14025 9447 14059
rect 10149 14025 10183 14059
rect 13553 14025 13587 14059
rect 15301 14025 15335 14059
rect 16865 14025 16899 14059
rect 17509 14025 17543 14059
rect 18705 14025 18739 14059
rect 20821 14025 20855 14059
rect 22293 14025 22327 14059
rect 22937 14025 22971 14059
rect 25605 14025 25639 14059
rect 30297 14025 30331 14059
rect 31125 14025 31159 14059
rect 4537 13957 4571 13991
rect 17233 13957 17267 13991
rect 19073 13957 19107 13991
rect 21005 13957 21039 13991
rect 21833 13957 21867 13991
rect 25789 13957 25823 13991
rect 3617 13889 3651 13923
rect 5273 13889 5307 13923
rect 17785 13889 17819 13923
rect 17969 13889 18003 13923
rect 18981 13889 19015 13923
rect 20453 13889 20487 13923
rect 21741 13889 21775 13923
rect 22109 13889 22143 13923
rect 3341 13821 3375 13855
rect 3433 13821 3467 13855
rect 3709 13821 3743 13855
rect 4721 13821 4755 13855
rect 4813 13821 4847 13855
rect 5089 13821 5123 13855
rect 5181 13821 5215 13855
rect 5457 13821 5491 13855
rect 5733 13821 5767 13855
rect 6193 13821 6227 13855
rect 6285 13821 6319 13855
rect 6469 13821 6503 13855
rect 6561 13821 6595 13855
rect 6745 13821 6779 13855
rect 7021 13821 7055 13855
rect 7113 13821 7147 13855
rect 7297 13821 7331 13855
rect 7389 13821 7423 13855
rect 7757 13821 7791 13855
rect 8125 13821 8159 13855
rect 8401 13821 8435 13855
rect 8585 13821 8619 13855
rect 8769 13821 8803 13855
rect 8953 13821 8987 13855
rect 9045 13821 9079 13855
rect 9137 13821 9171 13855
rect 9505 13821 9539 13855
rect 9689 13821 9723 13855
rect 9781 13821 9815 13855
rect 9873 13821 9907 13855
rect 13829 13821 13863 13855
rect 13921 13821 13955 13855
rect 14013 13821 14047 13855
rect 14197 13821 14231 13855
rect 15117 13821 15151 13855
rect 15301 13821 15335 13855
rect 17049 13821 17083 13855
rect 17141 13821 17175 13855
rect 17325 13821 17359 13855
rect 17693 13821 17727 13855
rect 17877 13821 17911 13855
rect 19165 13821 19199 13855
rect 19257 13821 19291 13855
rect 19441 13821 19475 13855
rect 21097 13821 21131 13855
rect 21281 13821 21315 13855
rect 21373 13821 21407 13855
rect 21465 13821 21499 13855
rect 22017 13821 22051 13855
rect 22293 13821 22327 13855
rect 22385 13821 22419 13855
rect 25697 13821 25731 13855
rect 25973 13821 26007 13855
rect 26065 13821 26099 13855
rect 28273 13821 28307 13855
rect 28365 13821 28399 13855
rect 28549 13821 28583 13855
rect 28641 13821 28675 13855
rect 28825 13821 28859 13855
rect 29929 13821 29963 13855
rect 30389 13821 30423 13855
rect 30941 13821 30975 13855
rect 4905 13753 4939 13787
rect 5641 13753 5675 13787
rect 7573 13753 7607 13787
rect 22569 13753 22603 13787
rect 30113 13753 30147 13787
rect 20821 13685 20855 13719
rect 22661 13685 22695 13719
rect 22753 13685 22787 13719
rect 29653 13685 29687 13719
rect 30021 13685 30055 13719
rect 857 13481 891 13515
rect 1869 13481 1903 13515
rect 2053 13481 2087 13515
rect 8861 13481 8895 13515
rect 12173 13481 12207 13515
rect 13001 13481 13035 13515
rect 16129 13481 16163 13515
rect 18889 13481 18923 13515
rect 22753 13481 22787 13515
rect 23121 13481 23155 13515
rect 25513 13481 25547 13515
rect 28733 13481 28767 13515
rect 1225 13413 1259 13447
rect 6561 13413 6595 13447
rect 7389 13413 7423 13447
rect 10517 13413 10551 13447
rect 22293 13413 22327 13447
rect 26065 13413 26099 13447
rect 26249 13413 26283 13447
rect 28993 13413 29027 13447
rect 29193 13413 29227 13447
rect 1041 13345 1075 13379
rect 1317 13345 1351 13379
rect 1928 13345 1962 13379
rect 2513 13345 2547 13379
rect 2697 13345 2731 13379
rect 2789 13345 2823 13379
rect 2881 13345 2915 13379
rect 3065 13345 3099 13379
rect 6469 13345 6503 13379
rect 6745 13345 6779 13379
rect 7573 13345 7607 13379
rect 8309 13345 8343 13379
rect 8401 13345 8435 13379
rect 8585 13345 8619 13379
rect 8677 13345 8711 13379
rect 10149 13345 10183 13379
rect 10297 13345 10331 13379
rect 10425 13345 10459 13379
rect 10614 13345 10648 13379
rect 11156 13345 11190 13379
rect 11253 13345 11287 13379
rect 11345 13345 11379 13379
rect 11473 13345 11507 13379
rect 11621 13345 11655 13379
rect 12633 13345 12667 13379
rect 13277 13345 13311 13379
rect 15025 13345 15059 13379
rect 15117 13345 15151 13379
rect 15209 13345 15243 13379
rect 15393 13345 15427 13379
rect 15853 13345 15887 13379
rect 16313 13345 16347 13379
rect 16497 13345 16531 13379
rect 17049 13345 17083 13379
rect 17233 13345 17267 13379
rect 17509 13345 17543 13379
rect 18797 13345 18831 13379
rect 19073 13345 19107 13379
rect 19165 13345 19199 13379
rect 19257 13345 19291 13379
rect 19441 13345 19475 13379
rect 20821 13345 20855 13379
rect 20913 13345 20947 13379
rect 21465 13345 21499 13379
rect 21649 13345 21683 13379
rect 21741 13345 21775 13379
rect 22017 13345 22051 13379
rect 22937 13345 22971 13379
rect 23213 13345 23247 13379
rect 24041 13345 24075 13379
rect 24409 13345 24443 13379
rect 24869 13345 24903 13379
rect 25329 13345 25363 13379
rect 25421 13345 25455 13379
rect 25605 13345 25639 13379
rect 25973 13345 26007 13379
rect 26433 13345 26467 13379
rect 26617 13345 26651 13379
rect 26709 13345 26743 13379
rect 26985 13345 27019 13379
rect 28089 13345 28123 13379
rect 28365 13345 28399 13379
rect 28457 13345 28491 13379
rect 28549 13345 28583 13379
rect 29837 13345 29871 13379
rect 30021 13345 30055 13379
rect 1409 13277 1443 13311
rect 12357 13277 12391 13311
rect 12449 13277 12483 13311
rect 12541 13277 12575 13311
rect 13185 13277 13219 13311
rect 13553 13277 13587 13311
rect 13645 13277 13679 13311
rect 14749 13277 14783 13311
rect 18981 13277 19015 13311
rect 21097 13277 21131 13311
rect 22201 13277 22235 13311
rect 25053 13277 25087 13311
rect 25145 13277 25179 13311
rect 26801 13277 26835 13311
rect 28273 13277 28307 13311
rect 7757 13209 7791 13243
rect 10793 13209 10827 13243
rect 10977 13209 11011 13243
rect 15577 13209 15611 13243
rect 17325 13209 17359 13243
rect 17417 13209 17451 13243
rect 21833 13209 21867 13243
rect 24685 13209 24719 13243
rect 24961 13209 24995 13243
rect 1501 13141 1535 13175
rect 2329 13141 2363 13175
rect 2881 13141 2915 13175
rect 3249 13141 3283 13175
rect 6929 13141 6963 13175
rect 16313 13141 16347 13175
rect 19257 13141 19291 13175
rect 21281 13141 21315 13175
rect 22201 13141 22235 13175
rect 24225 13141 24259 13175
rect 24593 13141 24627 13175
rect 26157 13141 26191 13175
rect 27169 13141 27203 13175
rect 28825 13141 28859 13175
rect 29009 13141 29043 13175
rect 29929 13141 29963 13175
rect 4445 12937 4479 12971
rect 5641 12937 5675 12971
rect 6745 12937 6779 12971
rect 8033 12937 8067 12971
rect 13185 12937 13219 12971
rect 13737 12937 13771 12971
rect 13829 12937 13863 12971
rect 16681 12937 16715 12971
rect 17325 12937 17359 12971
rect 17509 12937 17543 12971
rect 21097 12937 21131 12971
rect 22661 12937 22695 12971
rect 22753 12937 22787 12971
rect 29009 12937 29043 12971
rect 29377 12937 29411 12971
rect 4629 12869 4663 12903
rect 7389 12869 7423 12903
rect 8677 12869 8711 12903
rect 8769 12869 8803 12903
rect 10149 12869 10183 12903
rect 12541 12869 12575 12903
rect 12725 12869 12759 12903
rect 14841 12869 14875 12903
rect 17969 12869 18003 12903
rect 18981 12869 19015 12903
rect 22937 12869 22971 12903
rect 29837 12869 29871 12903
rect 29929 12869 29963 12903
rect 4353 12801 4387 12835
rect 6285 12801 6319 12835
rect 6377 12801 6411 12835
rect 6469 12801 6503 12835
rect 6929 12801 6963 12835
rect 7113 12801 7147 12835
rect 8401 12801 8435 12835
rect 10333 12801 10367 12835
rect 13645 12801 13679 12835
rect 15209 12801 15243 12835
rect 18337 12801 18371 12835
rect 19349 12801 19383 12835
rect 20821 12801 20855 12835
rect 22753 12801 22787 12835
rect 24869 12801 24903 12835
rect 26341 12801 26375 12835
rect 30297 12801 30331 12835
rect 30389 12801 30423 12835
rect 4261 12733 4295 12767
rect 4721 12733 4755 12767
rect 4997 12733 5031 12767
rect 5549 12733 5583 12767
rect 5641 12733 5675 12767
rect 6101 12733 6135 12767
rect 6561 12733 6595 12767
rect 7020 12733 7054 12767
rect 7205 12733 7239 12767
rect 7941 12733 7975 12767
rect 8125 12733 8159 12767
rect 8585 12733 8619 12767
rect 8861 12733 8895 12767
rect 10149 12733 10183 12767
rect 11443 12733 11477 12767
rect 11621 12733 11655 12767
rect 12265 12733 12299 12767
rect 12633 12733 12667 12767
rect 12817 12733 12851 12767
rect 13001 12733 13035 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 13921 12733 13955 12767
rect 15025 12733 15059 12767
rect 15301 12733 15335 12767
rect 15393 12733 15427 12767
rect 15577 12733 15611 12767
rect 16865 12733 16899 12767
rect 16957 12733 16991 12767
rect 17141 12733 17175 12767
rect 17233 12733 17267 12767
rect 17509 12733 17543 12767
rect 17877 12733 17911 12767
rect 18153 12733 18187 12767
rect 18429 12733 18463 12767
rect 18889 12733 18923 12767
rect 19165 12733 19199 12767
rect 19625 12733 19659 12767
rect 19717 12733 19751 12767
rect 19809 12733 19843 12767
rect 19993 12733 20027 12767
rect 20453 12733 20487 12767
rect 20913 12733 20947 12767
rect 22569 12733 22603 12767
rect 24041 12733 24075 12767
rect 24133 12733 24167 12767
rect 24501 12733 24535 12767
rect 24777 12733 24811 12767
rect 24961 12733 24995 12767
rect 26433 12733 26467 12767
rect 29196 12733 29230 12767
rect 29285 12733 29319 12767
rect 30573 12733 30607 12767
rect 30849 12733 30883 12767
rect 9781 12665 9815 12699
rect 24225 12665 24259 12699
rect 24343 12665 24377 12699
rect 29653 12665 29687 12699
rect 4813 12597 4847 12631
rect 5181 12597 5215 12631
rect 5273 12597 5307 12631
rect 11529 12597 11563 12631
rect 20545 12597 20579 12631
rect 20729 12597 20763 12631
rect 23857 12597 23891 12631
rect 26801 12597 26835 12631
rect 30757 12597 30791 12631
rect 1777 12393 1811 12427
rect 3249 12393 3283 12427
rect 4997 12393 5031 12427
rect 6837 12393 6871 12427
rect 9137 12393 9171 12427
rect 9873 12393 9907 12427
rect 13001 12393 13035 12427
rect 13737 12393 13771 12427
rect 15025 12393 15059 12427
rect 18245 12393 18279 12427
rect 22109 12393 22143 12427
rect 23673 12393 23707 12427
rect 26433 12393 26467 12427
rect 27445 12393 27479 12427
rect 27537 12393 27571 12427
rect 1593 12325 1627 12359
rect 4813 12325 4847 12359
rect 12449 12325 12483 12359
rect 13487 12325 13521 12359
rect 16865 12325 16899 12359
rect 26709 12325 26743 12359
rect 27721 12325 27755 12359
rect 28365 12325 28399 12359
rect 29101 12325 29135 12359
rect 1869 12257 1903 12291
rect 3433 12257 3467 12291
rect 3525 12257 3559 12291
rect 3709 12257 3743 12291
rect 3893 12257 3927 12291
rect 5089 12257 5123 12291
rect 7021 12257 7055 12291
rect 7205 12257 7239 12291
rect 7297 12257 7331 12291
rect 9321 12257 9355 12291
rect 9597 12257 9631 12291
rect 9781 12257 9815 12291
rect 10057 12257 10091 12291
rect 10517 12257 10551 12291
rect 12173 12257 12207 12291
rect 13185 12257 13219 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 13645 12257 13679 12291
rect 14013 12257 14047 12291
rect 14381 12257 14415 12291
rect 14544 12257 14578 12291
rect 14657 12257 14691 12291
rect 14749 12257 14783 12291
rect 15301 12257 15335 12291
rect 15485 12257 15519 12291
rect 16681 12257 16715 12291
rect 16957 12257 16991 12291
rect 17049 12257 17083 12291
rect 17693 12257 17727 12291
rect 17877 12257 17911 12291
rect 18061 12257 18095 12291
rect 18337 12257 18371 12291
rect 18981 12257 19015 12291
rect 19073 12257 19107 12291
rect 22661 12257 22695 12291
rect 22937 12257 22971 12291
rect 23121 12257 23155 12291
rect 23213 12257 23247 12291
rect 23305 12257 23339 12291
rect 23397 12257 23431 12291
rect 24409 12257 24443 12291
rect 24869 12257 24903 12291
rect 25145 12257 25179 12291
rect 25513 12257 25547 12291
rect 25697 12257 25731 12291
rect 26065 12257 26099 12291
rect 26249 12257 26283 12291
rect 26617 12257 26651 12291
rect 26801 12257 26835 12291
rect 26985 12257 27019 12291
rect 27077 12257 27111 12291
rect 27353 12257 27387 12291
rect 27997 12257 28031 12291
rect 28181 12257 28215 12291
rect 28457 12257 28491 12291
rect 28917 12257 28951 12291
rect 29193 12257 29227 12291
rect 30481 12257 30515 12291
rect 7113 12189 7147 12223
rect 9505 12189 9539 12223
rect 10241 12189 10275 12223
rect 10333 12189 10367 12223
rect 12265 12189 12299 12223
rect 12449 12189 12483 12223
rect 13921 12189 13955 12223
rect 14105 12189 14139 12223
rect 14197 12189 14231 12223
rect 15669 12189 15703 12223
rect 18889 12189 18923 12223
rect 19165 12189 19199 12223
rect 22385 12189 22419 12223
rect 25421 12189 25455 12223
rect 25605 12189 25639 12223
rect 26157 12189 26191 12223
rect 30205 12189 30239 12223
rect 1593 12121 1627 12155
rect 3617 12121 3651 12155
rect 4813 12121 4847 12155
rect 9413 12121 9447 12155
rect 10149 12121 10183 12155
rect 17233 12121 17267 12155
rect 18705 12121 18739 12155
rect 24133 12121 24167 12155
rect 24501 12121 24535 12155
rect 24961 12121 24995 12155
rect 27169 12121 27203 12155
rect 29929 12121 29963 12155
rect 15117 12053 15151 12087
rect 17417 12053 17451 12087
rect 22569 12053 22603 12087
rect 22753 12053 22787 12087
rect 23305 12053 23339 12087
rect 24593 12053 24627 12087
rect 24685 12053 24719 12087
rect 25329 12053 25363 12087
rect 28733 12053 28767 12087
rect 30113 12053 30147 12087
rect 1317 11849 1351 11883
rect 2237 11849 2271 11883
rect 2605 11849 2639 11883
rect 3341 11849 3375 11883
rect 5917 11849 5951 11883
rect 7573 11849 7607 11883
rect 8861 11849 8895 11883
rect 11989 11849 12023 11883
rect 15117 11849 15151 11883
rect 16773 11849 16807 11883
rect 17141 11849 17175 11883
rect 17785 11849 17819 11883
rect 19910 11849 19944 11883
rect 20269 11849 20303 11883
rect 21741 11849 21775 11883
rect 22017 11849 22051 11883
rect 22477 11849 22511 11883
rect 26249 11849 26283 11883
rect 27353 11849 27387 11883
rect 28089 11849 28123 11883
rect 28549 11849 28583 11883
rect 7849 11781 7883 11815
rect 10333 11781 10367 11815
rect 19717 11781 19751 11815
rect 30573 11781 30607 11815
rect 2973 11713 3007 11747
rect 3065 11713 3099 11747
rect 4096 11713 4130 11747
rect 4997 11713 5031 11747
rect 6377 11713 6411 11747
rect 6469 11713 6503 11747
rect 10793 11713 10827 11747
rect 15209 11713 15243 11747
rect 17693 11713 17727 11747
rect 18705 11713 18739 11747
rect 18797 11713 18831 11747
rect 20637 11713 20671 11747
rect 21557 11713 21591 11747
rect 26617 11713 26651 11747
rect 26893 11713 26927 11747
rect 30757 11713 30791 11747
rect 1593 11645 1627 11679
rect 1685 11645 1719 11679
rect 1777 11645 1811 11679
rect 1961 11645 1995 11679
rect 2053 11645 2087 11679
rect 2145 11645 2179 11679
rect 2849 11645 2883 11679
rect 3525 11645 3559 11679
rect 3893 11645 3927 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 5089 11645 5123 11679
rect 5825 11645 5859 11679
rect 6101 11645 6135 11679
rect 6653 11645 6687 11679
rect 7757 11645 7791 11679
rect 7941 11645 7975 11679
rect 8033 11645 8067 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 10241 11645 10275 11679
rect 10517 11645 10551 11679
rect 10609 11645 10643 11679
rect 11069 11645 11103 11679
rect 11161 11645 11195 11679
rect 11253 11645 11287 11679
rect 11437 11645 11471 11679
rect 11529 11645 11563 11679
rect 11621 11645 11655 11679
rect 11805 11645 11839 11679
rect 14473 11645 14507 11679
rect 14749 11645 14783 11679
rect 14841 11645 14875 11679
rect 14933 11645 14967 11679
rect 15393 11645 15427 11679
rect 16773 11645 16807 11679
rect 16865 11645 16899 11679
rect 17785 11645 17819 11679
rect 18981 11645 19015 11679
rect 20177 11645 20211 11679
rect 20453 11645 20487 11679
rect 21465 11645 21499 11679
rect 21741 11645 21775 11679
rect 22293 11645 22327 11679
rect 22385 11645 22419 11679
rect 22569 11645 22603 11679
rect 22753 11645 22787 11679
rect 24225 11645 24259 11679
rect 24593 11645 24627 11679
rect 25329 11645 25363 11679
rect 25605 11645 25639 11679
rect 25697 11645 25731 11679
rect 26408 11645 26442 11679
rect 27077 11645 27111 11679
rect 27169 11645 27203 11679
rect 28365 11645 28399 11679
rect 28641 11645 28675 11679
rect 29469 11645 29503 11679
rect 29561 11645 29595 11679
rect 29745 11645 29779 11679
rect 29929 11645 29963 11679
rect 30205 11645 30239 11679
rect 30941 11645 30975 11679
rect 3801 11577 3835 11611
rect 4169 11577 4203 11611
rect 4629 11577 4663 11611
rect 8861 11577 8895 11611
rect 14611 11577 14645 11611
rect 20085 11577 20119 11611
rect 25421 11577 25455 11611
rect 25973 11577 26007 11611
rect 27353 11577 27387 11611
rect 2421 11509 2455 11543
rect 3709 11509 3743 11543
rect 3985 11509 4019 11543
rect 6285 11509 6319 11543
rect 6837 11509 6871 11543
rect 8401 11509 8435 11543
rect 10701 11509 10735 11543
rect 17233 11509 17267 11543
rect 17417 11509 17451 11543
rect 19165 11509 19199 11543
rect 19875 11509 19909 11543
rect 21281 11509 21315 11543
rect 24041 11509 24075 11543
rect 24409 11509 24443 11543
rect 25506 11509 25540 11543
rect 26525 11509 26559 11543
rect 29285 11509 29319 11543
rect 29653 11509 29687 11543
rect 3617 11305 3651 11339
rect 4629 11305 4663 11339
rect 6745 11305 6779 11339
rect 8033 11305 8067 11339
rect 11621 11305 11655 11339
rect 12265 11305 12299 11339
rect 14289 11305 14323 11339
rect 15209 11305 15243 11339
rect 16865 11305 16899 11339
rect 22937 11305 22971 11339
rect 23489 11305 23523 11339
rect 25697 11305 25731 11339
rect 29469 11305 29503 11339
rect 30297 11305 30331 11339
rect 4077 11237 4111 11271
rect 15025 11237 15059 11271
rect 20361 11237 20395 11271
rect 24777 11237 24811 11271
rect 25191 11237 25225 11271
rect 25421 11237 25455 11271
rect 27629 11237 27663 11271
rect 30849 11237 30883 11271
rect 1409 11169 1443 11203
rect 1501 11169 1535 11203
rect 2145 11169 2179 11203
rect 2513 11169 2547 11203
rect 2881 11169 2915 11203
rect 3065 11169 3099 11203
rect 3157 11169 3191 11203
rect 3341 11169 3375 11203
rect 3433 11169 3467 11203
rect 4629 11169 4663 11203
rect 4997 11169 5031 11203
rect 6929 11169 6963 11203
rect 7205 11169 7239 11203
rect 7941 11169 7975 11203
rect 8125 11169 8159 11203
rect 8953 11169 8987 11203
rect 9137 11169 9171 11203
rect 9413 11169 9447 11203
rect 9597 11169 9631 11203
rect 10977 11169 11011 11203
rect 11161 11169 11195 11203
rect 11345 11169 11379 11203
rect 11437 11169 11471 11203
rect 11529 11169 11563 11203
rect 11805 11169 11839 11203
rect 12633 11169 12667 11203
rect 12909 11169 12943 11203
rect 13093 11169 13127 11203
rect 13185 11169 13219 11203
rect 13369 11169 13403 11203
rect 14105 11169 14139 11203
rect 14289 11169 14323 11203
rect 14749 11169 14783 11203
rect 15301 11169 15335 11203
rect 16359 11169 16393 11203
rect 16497 11169 16531 11203
rect 16589 11169 16623 11203
rect 16681 11169 16715 11203
rect 20269 11169 20303 11203
rect 20453 11169 20487 11203
rect 22845 11169 22879 11203
rect 23029 11169 23063 11203
rect 23673 11169 23707 11203
rect 23765 11169 23799 11203
rect 23949 11169 23983 11203
rect 25053 11169 25087 11203
rect 25329 11169 25363 11203
rect 25513 11169 25547 11203
rect 27169 11169 27203 11203
rect 27261 11169 27295 11203
rect 27353 11169 27387 11203
rect 27445 11169 27479 11203
rect 27905 11169 27939 11203
rect 27997 11169 28031 11203
rect 28089 11169 28123 11203
rect 28273 11169 28307 11203
rect 28457 11169 28491 11203
rect 29101 11169 29135 11203
rect 29745 11169 29779 11203
rect 29837 11169 29871 11203
rect 29929 11169 29963 11203
rect 30113 11169 30147 11203
rect 30573 11169 30607 11203
rect 2237 11101 2271 11135
rect 4445 11101 4479 11135
rect 7113 11101 7147 11135
rect 12449 11101 12483 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 15097 11101 15131 11135
rect 16221 11101 16255 11135
rect 23857 11101 23891 11135
rect 28917 11101 28951 11135
rect 29377 11101 29411 11135
rect 11805 11033 11839 11067
rect 13001 11033 13035 11067
rect 29285 11033 29319 11067
rect 31033 11033 31067 11067
rect 3985 10965 4019 10999
rect 6929 10965 6963 10999
rect 9137 10965 9171 10999
rect 9597 10965 9631 10999
rect 13277 10965 13311 10999
rect 14381 10965 14415 10999
rect 24501 10965 24535 10999
rect 26985 10965 27019 10999
rect 28549 10965 28583 10999
rect 3893 10761 3927 10795
rect 6101 10761 6135 10795
rect 6837 10761 6871 10795
rect 7757 10761 7791 10795
rect 8033 10761 8067 10795
rect 8217 10761 8251 10795
rect 17141 10761 17175 10795
rect 19441 10761 19475 10795
rect 22385 10761 22419 10795
rect 23029 10761 23063 10795
rect 23949 10761 23983 10795
rect 24777 10761 24811 10795
rect 25789 10761 25823 10795
rect 27629 10761 27663 10795
rect 1961 10693 1995 10727
rect 5089 10693 5123 10727
rect 6469 10693 6503 10727
rect 7021 10693 7055 10727
rect 8677 10693 8711 10727
rect 9781 10693 9815 10727
rect 15531 10693 15565 10727
rect 15669 10693 15703 10727
rect 21281 10693 21315 10727
rect 26617 10693 26651 10727
rect 27169 10693 27203 10727
rect 27445 10693 27479 10727
rect 30389 10693 30423 10727
rect 2053 10625 2087 10659
rect 3985 10625 4019 10659
rect 6193 10625 6227 10659
rect 6653 10625 6687 10659
rect 9045 10625 9079 10659
rect 9137 10625 9171 10659
rect 11529 10625 11563 10659
rect 14013 10625 14047 10659
rect 15761 10625 15795 10659
rect 20453 10625 20487 10659
rect 24685 10625 24719 10659
rect 26157 10625 26191 10659
rect 1777 10557 1811 10591
rect 3249 10557 3283 10591
rect 3342 10557 3376 10591
rect 3714 10557 3748 10591
rect 4353 10557 4387 10591
rect 4813 10557 4847 10591
rect 5089 10557 5123 10591
rect 5273 10557 5307 10591
rect 5365 10557 5399 10591
rect 5733 10557 5767 10591
rect 6009 10557 6043 10591
rect 6101 10557 6135 10591
rect 6561 10557 6595 10591
rect 6837 10557 6871 10591
rect 7113 10557 7147 10591
rect 7205 10557 7239 10591
rect 7481 10557 7515 10591
rect 7573 10557 7607 10591
rect 8861 10557 8895 10591
rect 9229 10557 9263 10591
rect 9413 10557 9447 10591
rect 9689 10557 9723 10591
rect 9873 10557 9907 10591
rect 9965 10557 9999 10591
rect 10149 10557 10183 10591
rect 10517 10557 10551 10591
rect 10701 10551 10735 10585
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 11342 10557 11376 10591
rect 11713 10557 11747 10591
rect 11805 10557 11839 10591
rect 13645 10557 13679 10591
rect 13921 10557 13955 10591
rect 14197 10557 14231 10591
rect 14473 10557 14507 10591
rect 14565 10557 14599 10591
rect 14749 10557 14783 10591
rect 15393 10557 15427 10591
rect 15853 10557 15887 10591
rect 17417 10557 17451 10591
rect 17509 10557 17543 10591
rect 17601 10557 17635 10591
rect 17785 10557 17819 10591
rect 18061 10557 18095 10591
rect 18337 10557 18371 10591
rect 18521 10557 18555 10591
rect 18889 10557 18923 10591
rect 19161 10557 19195 10591
rect 19257 10557 19291 10591
rect 19993 10557 20027 10591
rect 21465 10557 21499 10591
rect 21557 10557 21591 10591
rect 21741 10557 21775 10591
rect 21833 10557 21867 10591
rect 22661 10557 22695 10591
rect 23121 10557 23155 10591
rect 24133 10557 24167 10591
rect 24225 10557 24259 10591
rect 24501 10557 24535 10591
rect 24593 10557 24627 10591
rect 24961 10557 24995 10591
rect 25973 10557 26007 10591
rect 26249 10557 26283 10591
rect 26341 10557 26375 10591
rect 26433 10557 26467 10591
rect 26617 10557 26651 10591
rect 26709 10557 26743 10591
rect 27353 10557 27387 10591
rect 28641 10557 28675 10591
rect 29469 10557 29503 10591
rect 30021 10557 30055 10591
rect 30389 10557 30423 10591
rect 30665 10557 30699 10591
rect 31033 10557 31067 10591
rect 3525 10489 3559 10523
rect 3617 10489 3651 10523
rect 4169 10489 4203 10523
rect 7389 10489 7423 10523
rect 7849 10489 7883 10523
rect 8049 10489 8083 10523
rect 9505 10489 9539 10523
rect 18429 10489 18463 10523
rect 19073 10489 19107 10523
rect 20085 10489 20119 10523
rect 20190 10489 20224 10523
rect 20295 10489 20329 10523
rect 24317 10489 24351 10523
rect 25145 10489 25179 10523
rect 27597 10489 27631 10523
rect 27813 10489 27847 10523
rect 29745 10489 29779 10523
rect 1593 10421 1627 10455
rect 5549 10421 5583 10455
rect 5641 10421 5675 10455
rect 11529 10421 11563 10455
rect 11621 10421 11655 10455
rect 14657 10421 14691 10455
rect 17969 10421 18003 10455
rect 18705 10421 18739 10455
rect 19809 10421 19843 10455
rect 22753 10421 22787 10455
rect 22845 10421 22879 10455
rect 26893 10421 26927 10455
rect 28825 10421 28859 10455
rect 29285 10421 29319 10455
rect 3617 10217 3651 10251
rect 3801 10217 3835 10251
rect 6285 10217 6319 10251
rect 8309 10217 8343 10251
rect 9045 10217 9079 10251
rect 10241 10217 10275 10251
rect 10977 10217 11011 10251
rect 21649 10217 21683 10251
rect 23857 10217 23891 10251
rect 24025 10217 24059 10251
rect 24685 10217 24719 10251
rect 26249 10217 26283 10251
rect 3525 10149 3559 10183
rect 9965 10149 9999 10183
rect 14473 10149 14507 10183
rect 14565 10149 14599 10183
rect 16957 10149 16991 10183
rect 17141 10149 17175 10183
rect 22937 10149 22971 10183
rect 24225 10149 24259 10183
rect 29377 10149 29411 10183
rect 3433 10081 3467 10115
rect 3893 10081 3927 10115
rect 4169 10081 4203 10115
rect 6193 10081 6227 10115
rect 6745 10081 6779 10115
rect 7021 10081 7055 10115
rect 7665 10081 7699 10115
rect 8493 10081 8527 10115
rect 8677 10081 8711 10115
rect 9229 10081 9263 10115
rect 9321 10081 9355 10115
rect 9505 10081 9539 10115
rect 9597 10081 9631 10115
rect 9689 10081 9723 10115
rect 9873 10081 9907 10115
rect 10057 10081 10091 10115
rect 11069 10081 11103 10115
rect 11437 10081 11471 10115
rect 12909 10081 12943 10115
rect 13001 10081 13035 10115
rect 13185 10081 13219 10115
rect 13277 10081 13311 10115
rect 14335 10081 14369 10115
rect 14657 10081 14691 10115
rect 16497 10081 16531 10115
rect 17049 10081 17083 10115
rect 17233 10081 17267 10115
rect 18981 10081 19015 10115
rect 19165 10081 19199 10115
rect 20821 10081 20855 10115
rect 20913 10081 20947 10115
rect 21097 10081 21131 10115
rect 21833 10081 21867 10115
rect 22017 10081 22051 10115
rect 22109 10081 22143 10115
rect 23029 10081 23063 10115
rect 23305 10081 23339 10115
rect 24501 10081 24535 10115
rect 24869 10081 24903 10115
rect 25789 10081 25823 10115
rect 26065 10081 26099 10115
rect 27261 10081 27295 10115
rect 27537 10081 27571 10115
rect 28181 10081 28215 10115
rect 28457 10081 28491 10115
rect 28733 10081 28767 10115
rect 29009 10081 29043 10115
rect 29561 10081 29595 10115
rect 29653 10081 29687 10115
rect 29745 10081 29779 10115
rect 29837 10081 29871 10115
rect 30113 10081 30147 10115
rect 30205 10081 30239 10115
rect 30389 10081 30423 10115
rect 30665 10081 30699 10115
rect 30849 10081 30883 10115
rect 30941 10081 30975 10115
rect 31033 10081 31067 10115
rect 4261 10013 4295 10047
rect 6653 10013 6687 10047
rect 8769 10013 8803 10047
rect 11161 10013 11195 10047
rect 12725 10013 12759 10047
rect 14197 10013 14231 10047
rect 14841 10013 14875 10047
rect 16773 10013 16807 10047
rect 16865 10013 16899 10047
rect 19257 10013 19291 10047
rect 19349 10013 19383 10047
rect 19441 10013 19475 10047
rect 21925 10013 21959 10047
rect 24409 10013 24443 10047
rect 24777 10013 24811 10047
rect 25881 10013 25915 10047
rect 25973 10013 26007 10047
rect 26617 10013 26651 10047
rect 26709 10013 26743 10047
rect 26801 10013 26835 10047
rect 26893 10013 26927 10047
rect 27077 10013 27111 10047
rect 27997 10013 28031 10047
rect 28273 10013 28307 10047
rect 28365 10013 28399 10047
rect 3249 9945 3283 9979
rect 16589 9945 16623 9979
rect 19717 9945 19751 9979
rect 26433 9945 26467 9979
rect 27353 9945 27387 9979
rect 27445 9945 27479 9979
rect 7757 9877 7791 9911
rect 11345 9877 11379 9911
rect 24041 9877 24075 9911
rect 25053 9877 25087 9911
rect 29377 9877 29411 9911
rect 31309 9877 31343 9911
rect 1777 9673 1811 9707
rect 3249 9673 3283 9707
rect 5457 9673 5491 9707
rect 5917 9673 5951 9707
rect 8033 9673 8067 9707
rect 11345 9673 11379 9707
rect 12357 9673 12391 9707
rect 13093 9673 13127 9707
rect 20085 9673 20119 9707
rect 22017 9673 22051 9707
rect 22845 9673 22879 9707
rect 26801 9673 26835 9707
rect 27261 9673 27295 9707
rect 28273 9673 28307 9707
rect 1317 9605 1351 9639
rect 4813 9605 4847 9639
rect 7665 9605 7699 9639
rect 8861 9605 8895 9639
rect 8953 9605 8987 9639
rect 12633 9605 12667 9639
rect 14013 9605 14047 9639
rect 15945 9605 15979 9639
rect 17141 9605 17175 9639
rect 21741 9605 21775 9639
rect 22293 9605 22327 9639
rect 25237 9605 25271 9639
rect 26525 9605 26559 9639
rect 27077 9605 27111 9639
rect 29285 9605 29319 9639
rect 5365 9537 5399 9571
rect 5733 9537 5767 9571
rect 6193 9537 6227 9571
rect 8217 9537 8251 9571
rect 9965 9537 9999 9571
rect 10241 9537 10275 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 12725 9537 12759 9571
rect 12817 9537 12851 9571
rect 15301 9537 15335 9571
rect 16221 9537 16255 9571
rect 16497 9537 16531 9571
rect 19349 9537 19383 9571
rect 20269 9537 20303 9571
rect 26709 9537 26743 9571
rect 27537 9537 27571 9571
rect 29561 9537 29595 9571
rect 29929 9537 29963 9571
rect 1501 9469 1535 9503
rect 1593 9469 1627 9503
rect 1869 9469 1903 9503
rect 3433 9469 3467 9503
rect 3525 9469 3559 9503
rect 3709 9469 3743 9503
rect 3801 9469 3835 9503
rect 4721 9469 4755 9503
rect 4905 9469 4939 9503
rect 5181 9469 5215 9503
rect 5641 9469 5675 9503
rect 6009 9469 6043 9503
rect 7021 9469 7055 9503
rect 7205 9469 7239 9503
rect 7481 9469 7515 9503
rect 7941 9469 7975 9503
rect 8769 9469 8803 9503
rect 9045 9469 9079 9503
rect 9229 9469 9263 9503
rect 9781 9469 9815 9503
rect 10149 9469 10183 9503
rect 10609 9469 10643 9503
rect 11529 9469 11563 9503
rect 11805 9469 11839 9503
rect 12541 9469 12575 9503
rect 13001 9469 13035 9503
rect 13093 9469 13127 9503
rect 13277 9469 13311 9503
rect 13921 9469 13955 9503
rect 14105 9469 14139 9503
rect 15485 9469 15519 9503
rect 16359 9469 16393 9503
rect 17417 9469 17451 9503
rect 17601 9469 17635 9503
rect 17693 9469 17727 9503
rect 17877 9469 17911 9503
rect 18061 9469 18095 9503
rect 18705 9469 18739 9503
rect 19165 9469 19199 9503
rect 19441 9469 19475 9503
rect 19625 9469 19659 9503
rect 19717 9469 19751 9503
rect 19829 9469 19863 9503
rect 20453 9469 20487 9503
rect 20545 9469 20579 9503
rect 20729 9469 20763 9503
rect 20821 9469 20855 9503
rect 21741 9469 21775 9503
rect 21925 9469 21959 9503
rect 22201 9469 22235 9503
rect 22385 9469 22419 9503
rect 22477 9469 22511 9503
rect 23029 9469 23063 9503
rect 23305 9469 23339 9503
rect 24133 9469 24167 9503
rect 24409 9469 24443 9503
rect 24501 9469 24535 9503
rect 24777 9469 24811 9503
rect 24961 9469 24995 9503
rect 25237 9469 25271 9503
rect 25513 9469 25547 9503
rect 25605 9469 25639 9503
rect 26249 9469 26283 9503
rect 26617 9469 26651 9503
rect 26893 9469 26927 9503
rect 27169 9469 27203 9503
rect 27353 9469 27387 9503
rect 29469 9469 29503 9503
rect 29653 9469 29687 9503
rect 29745 9469 29779 9503
rect 30205 9469 30239 9503
rect 30297 9469 30331 9503
rect 30389 9469 30423 9503
rect 30573 9469 30607 9503
rect 30849 9469 30883 9503
rect 31033 9469 31067 9503
rect 31125 9469 31159 9503
rect 5457 9401 5491 9435
rect 5549 9401 5583 9435
rect 5917 9401 5951 9435
rect 6745 9401 6779 9435
rect 9505 9401 9539 9435
rect 14289 9401 14323 9435
rect 14841 9401 14875 9435
rect 17969 9401 18003 9435
rect 18863 9401 18897 9435
rect 18981 9401 19015 9435
rect 19073 9401 19107 9435
rect 25881 9401 25915 9435
rect 26525 9401 26559 9435
rect 27813 9401 27847 9435
rect 28365 9401 28399 9435
rect 30665 9401 30699 9435
rect 4997 9333 5031 9367
rect 7297 9333 7331 9367
rect 8217 9333 8251 9367
rect 8585 9333 8619 9367
rect 11713 9333 11747 9367
rect 14381 9333 14415 9367
rect 15117 9333 15151 9367
rect 17233 9333 17267 9367
rect 23213 9333 23247 9367
rect 26341 9333 26375 9367
rect 1041 9129 1075 9163
rect 2605 9129 2639 9163
rect 3525 9129 3559 9163
rect 11345 9129 11379 9163
rect 12173 9129 12207 9163
rect 16129 9129 16163 9163
rect 20453 9129 20487 9163
rect 23029 9129 23063 9163
rect 25881 9129 25915 9163
rect 27629 9129 27663 9163
rect 28457 9129 28491 9163
rect 29837 9129 29871 9163
rect 6561 9061 6595 9095
rect 9597 9061 9631 9095
rect 15485 9061 15519 9095
rect 24777 9061 24811 9095
rect 30665 9061 30699 9095
rect 1225 8993 1259 9027
rect 1409 8993 1443 9027
rect 1501 8993 1535 9027
rect 1961 8993 1995 9027
rect 2697 8993 2731 9027
rect 3065 8993 3099 9027
rect 3433 8993 3467 9027
rect 3617 8993 3651 9027
rect 4537 8993 4571 9027
rect 4721 8993 4755 9027
rect 4997 8993 5031 9027
rect 5181 8993 5215 9027
rect 6285 8993 6319 9027
rect 6929 8993 6963 9027
rect 8677 8993 8711 9027
rect 9137 8993 9171 9027
rect 9229 8993 9263 9027
rect 9413 8993 9447 9027
rect 9505 8993 9539 9027
rect 9689 8993 9723 9027
rect 10977 8993 11011 9027
rect 11161 8993 11195 9027
rect 12081 8993 12115 9027
rect 12265 8993 12299 9027
rect 12725 8993 12759 9027
rect 13829 8993 13863 9027
rect 14013 8993 14047 9027
rect 14289 8993 14323 9027
rect 14473 8993 14507 9027
rect 15025 8993 15059 9027
rect 15669 8993 15703 9027
rect 15761 8993 15795 9027
rect 15945 8993 15979 9027
rect 16497 8993 16531 9027
rect 17325 8993 17359 9027
rect 17785 8993 17819 9027
rect 18429 8993 18463 9027
rect 18613 8993 18647 9027
rect 18981 8993 19015 9027
rect 19717 8993 19751 9027
rect 19993 8993 20027 9027
rect 20177 8993 20211 9027
rect 21281 8993 21315 9027
rect 21557 8993 21591 9027
rect 21649 8993 21683 9027
rect 21833 8993 21867 9027
rect 23305 8993 23339 9027
rect 23397 8993 23431 9027
rect 24041 8993 24075 9027
rect 24225 8993 24259 9027
rect 24501 8993 24535 9027
rect 24869 8993 24903 9027
rect 25421 8993 25455 9027
rect 25697 8993 25731 9027
rect 27169 8993 27203 9027
rect 27445 8993 27479 9027
rect 28089 8993 28123 9027
rect 28273 8993 28307 9027
rect 28917 8993 28951 9027
rect 29101 8993 29135 9027
rect 29377 8993 29411 9027
rect 30113 8993 30147 9027
rect 30205 8993 30239 9027
rect 30297 8993 30331 9027
rect 30481 8993 30515 9027
rect 1869 8925 1903 8959
rect 8769 8925 8803 8959
rect 13001 8925 13035 8959
rect 14657 8925 14691 8959
rect 14841 8925 14875 8959
rect 15577 8925 15611 8959
rect 16405 8925 16439 8959
rect 17509 8925 17543 8959
rect 17601 8925 17635 8959
rect 20453 8925 20487 8959
rect 21373 8925 21407 8959
rect 23213 8925 23247 8959
rect 23489 8925 23523 8959
rect 25513 8925 25547 8959
rect 3249 8857 3283 8891
rect 7113 8857 7147 8891
rect 12909 8857 12943 8891
rect 15301 8857 15335 8891
rect 17417 8857 17451 8891
rect 18521 8857 18555 8891
rect 24409 8857 24443 8891
rect 27261 8857 27295 8891
rect 27353 8857 27387 8891
rect 29377 8857 29411 8891
rect 30849 8857 30883 8891
rect 4629 8789 4663 8823
rect 4997 8789 5031 8823
rect 8677 8789 8711 8823
rect 9045 8789 9079 8823
rect 9413 8789 9447 8823
rect 11161 8789 11195 8823
rect 12541 8789 12575 8823
rect 16497 8789 16531 8823
rect 17141 8789 17175 8823
rect 19165 8789 19199 8823
rect 19809 8789 19843 8823
rect 20269 8789 20303 8823
rect 25053 8789 25087 8823
rect 25697 8789 25731 8823
rect 26893 8789 26927 8823
rect 28641 8789 28675 8823
rect 1777 8585 1811 8619
rect 2053 8585 2087 8619
rect 4261 8585 4295 8619
rect 5457 8585 5491 8619
rect 6469 8585 6503 8619
rect 7481 8585 7515 8619
rect 12081 8585 12115 8619
rect 13185 8585 13219 8619
rect 14381 8585 14415 8619
rect 14565 8585 14599 8619
rect 22017 8585 22051 8619
rect 22385 8585 22419 8619
rect 23121 8585 23155 8619
rect 24409 8585 24443 8619
rect 25605 8585 25639 8619
rect 29929 8585 29963 8619
rect 30665 8585 30699 8619
rect 1593 8517 1627 8551
rect 2237 8517 2271 8551
rect 5549 8517 5583 8551
rect 6837 8517 6871 8551
rect 7205 8517 7239 8551
rect 8401 8517 8435 8551
rect 15025 8517 15059 8551
rect 19073 8517 19107 8551
rect 20177 8517 20211 8551
rect 21557 8517 21591 8551
rect 25237 8517 25271 8551
rect 26065 8517 26099 8551
rect 26433 8517 26467 8551
rect 28457 8517 28491 8551
rect 29285 8517 29319 8551
rect 5365 8449 5399 8483
rect 7113 8449 7147 8483
rect 7573 8449 7607 8483
rect 8677 8449 8711 8483
rect 8769 8449 8803 8483
rect 11161 8449 11195 8483
rect 11345 8449 11379 8483
rect 11529 8449 11563 8483
rect 12541 8449 12575 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 17417 8449 17451 8483
rect 17693 8449 17727 8483
rect 23305 8449 23339 8483
rect 23397 8449 23431 8483
rect 26249 8449 26283 8483
rect 29377 8449 29411 8483
rect 1685 8381 1719 8415
rect 1869 8381 1903 8415
rect 2053 8381 2087 8415
rect 3249 8381 3283 8415
rect 3433 8381 3467 8415
rect 3525 8381 3559 8415
rect 3617 8381 3651 8415
rect 3709 8381 3743 8415
rect 4353 8381 4387 8415
rect 4721 8381 4755 8415
rect 4905 8381 4939 8415
rect 4997 8381 5031 8415
rect 5089 8381 5123 8415
rect 6469 8381 6503 8415
rect 6653 8381 6687 8415
rect 7021 8381 7055 8415
rect 7297 8381 7331 8415
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 8585 8381 8619 8415
rect 8861 8381 8895 8415
rect 9045 8381 9079 8415
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 11437 8381 11471 8415
rect 11621 8381 11655 8415
rect 12265 8381 12299 8415
rect 12357 8381 12391 8415
rect 12449 8381 12483 8415
rect 12725 8381 12759 8415
rect 12817 8381 12851 8415
rect 13001 8381 13035 8415
rect 13737 8381 13771 8415
rect 13921 8381 13955 8415
rect 14013 8381 14047 8415
rect 14105 8381 14139 8415
rect 14473 8381 14507 8415
rect 14749 8381 14783 8415
rect 15301 8381 15335 8415
rect 17509 8381 17543 8415
rect 17877 8381 17911 8415
rect 17969 8381 18003 8415
rect 19901 8381 19935 8415
rect 20545 8381 20579 8415
rect 20821 8381 20855 8415
rect 20913 8381 20947 8415
rect 21189 8381 21223 8415
rect 21465 8381 21499 8415
rect 21833 8381 21867 8415
rect 21925 8381 21959 8415
rect 22109 8381 22143 8415
rect 22293 8381 22327 8415
rect 22661 8381 22695 8415
rect 22753 8381 22787 8415
rect 22845 8381 22879 8415
rect 23029 8381 23063 8415
rect 23489 8381 23523 8415
rect 23581 8381 23615 8415
rect 23949 8381 23983 8415
rect 24225 8381 24259 8415
rect 24409 8381 24443 8415
rect 24593 8381 24627 8415
rect 25237 8381 25271 8415
rect 25421 8381 25455 8415
rect 25513 8381 25547 8415
rect 25789 8381 25823 8415
rect 25881 8381 25915 8415
rect 26157 8381 26191 8415
rect 26525 8381 26559 8415
rect 28181 8381 28215 8415
rect 28365 8381 28399 8415
rect 28549 8381 28583 8415
rect 28641 8381 28675 8415
rect 29193 8381 29227 8415
rect 29469 8381 29503 8415
rect 30113 8381 30147 8415
rect 30297 8381 30331 8415
rect 30849 8381 30883 8415
rect 1317 8313 1351 8347
rect 3893 8313 3927 8347
rect 4537 8313 4571 8347
rect 5917 8313 5951 8347
rect 15117 8313 15151 8347
rect 17693 8313 17727 8347
rect 18705 8313 18739 8347
rect 18889 8313 18923 8347
rect 20177 8313 20211 8347
rect 21373 8313 21407 8347
rect 23857 8313 23891 8347
rect 26249 8313 26283 8347
rect 27077 8313 27111 8347
rect 27253 8313 27287 8347
rect 27445 8313 27479 8347
rect 27721 8313 27755 8347
rect 1409 8245 1443 8279
rect 7941 8245 7975 8279
rect 10425 8245 10459 8279
rect 17049 8245 17083 8279
rect 19993 8245 20027 8279
rect 27813 8245 27847 8279
rect 29009 8245 29043 8279
rect 11437 8041 11471 8075
rect 11529 8041 11563 8075
rect 15577 8041 15611 8075
rect 17141 8041 17175 8075
rect 18521 8041 18555 8075
rect 20637 8041 20671 8075
rect 23029 8041 23063 8075
rect 28089 8041 28123 8075
rect 28733 8041 28767 8075
rect 30757 8041 30791 8075
rect 1593 7973 1627 8007
rect 1961 7973 1995 8007
rect 8861 7973 8895 8007
rect 8953 7973 8987 8007
rect 11897 7973 11931 8007
rect 13553 7973 13587 8007
rect 13737 7973 13771 8007
rect 19349 7973 19383 8007
rect 21833 7973 21867 8007
rect 27261 7973 27295 8007
rect 1225 7905 1259 7939
rect 1409 7905 1443 7939
rect 1501 7905 1535 7939
rect 1777 7905 1811 7939
rect 2421 7905 2455 7939
rect 4629 7905 4663 7939
rect 4905 7905 4939 7939
rect 5273 7905 5307 7939
rect 5457 7905 5491 7939
rect 8585 7905 8619 7939
rect 9229 7905 9263 7939
rect 9413 7905 9447 7939
rect 9689 7905 9723 7939
rect 10977 7905 11011 7939
rect 11253 7905 11287 7939
rect 11713 7905 11747 7939
rect 11805 7905 11839 7939
rect 12081 7905 12115 7939
rect 12173 7905 12207 7939
rect 12357 7905 12391 7939
rect 13185 7905 13219 7939
rect 13645 7905 13679 7939
rect 13829 7905 13863 7939
rect 14105 7905 14139 7939
rect 14197 7905 14231 7939
rect 14381 7905 14415 7939
rect 14473 7905 14507 7939
rect 14749 7905 14783 7939
rect 14933 7905 14967 7939
rect 15025 7905 15059 7939
rect 15117 7905 15151 7939
rect 15297 7915 15331 7949
rect 15393 7939 15427 7973
rect 15669 7905 15703 7939
rect 17049 7905 17083 7939
rect 17325 7905 17359 7939
rect 18705 7905 18739 7939
rect 18797 7905 18831 7939
rect 18889 7905 18923 7939
rect 19007 7905 19041 7939
rect 19165 7905 19199 7939
rect 19257 7905 19291 7939
rect 19441 7905 19475 7939
rect 19533 7905 19567 7939
rect 19717 7905 19751 7939
rect 20361 7905 20395 7939
rect 20545 7905 20579 7939
rect 20637 7905 20671 7939
rect 22017 7905 22051 7939
rect 22109 7905 22143 7939
rect 22661 7905 22695 7939
rect 23213 7905 23247 7939
rect 23489 7905 23523 7939
rect 23673 7905 23707 7939
rect 24501 7905 24535 7939
rect 24593 7905 24627 7939
rect 24777 7905 24811 7939
rect 25145 7905 25179 7939
rect 25329 7905 25363 7939
rect 25421 7905 25455 7939
rect 25697 7905 25731 7939
rect 26065 7905 26099 7939
rect 26709 7905 26743 7939
rect 26985 7905 27019 7939
rect 27169 7905 27203 7939
rect 27537 7905 27571 7939
rect 27905 7905 27939 7939
rect 28273 7905 28307 7939
rect 28549 7905 28583 7939
rect 28947 7905 28981 7939
rect 29101 7905 29135 7939
rect 29377 7905 29411 7939
rect 29561 7905 29595 7939
rect 29929 7905 29963 7939
rect 30481 7905 30515 7939
rect 30849 7905 30883 7939
rect 8493 7837 8527 7871
rect 8861 7837 8895 7871
rect 9321 7837 9355 7871
rect 11161 7837 11195 7871
rect 16589 7837 16623 7871
rect 16681 7837 16715 7871
rect 16773 7837 16807 7871
rect 16865 7837 16899 7871
rect 23305 7837 23339 7871
rect 24961 7837 24995 7871
rect 25237 7837 25271 7871
rect 1409 7769 1443 7803
rect 4905 7769 4939 7803
rect 5457 7769 5491 7803
rect 9505 7769 9539 7803
rect 15393 7769 15427 7803
rect 19625 7769 19659 7803
rect 23397 7769 23431 7803
rect 24685 7769 24719 7803
rect 28365 7769 28399 7803
rect 28457 7769 28491 7803
rect 30297 7769 30331 7803
rect 2237 7701 2271 7735
rect 8677 7701 8711 7735
rect 10977 7701 11011 7735
rect 12633 7701 12667 7735
rect 13921 7701 13955 7735
rect 14565 7701 14599 7735
rect 16405 7701 16439 7735
rect 17325 7701 17359 7735
rect 21833 7701 21867 7735
rect 22293 7701 22327 7735
rect 22477 7701 22511 7735
rect 24317 7701 24351 7735
rect 25973 7701 26007 7735
rect 26249 7701 26283 7735
rect 26525 7701 26559 7735
rect 29469 7701 29503 7735
rect 4905 7497 4939 7531
rect 5089 7497 5123 7531
rect 7021 7497 7055 7531
rect 9137 7497 9171 7531
rect 10241 7497 10275 7531
rect 14473 7497 14507 7531
rect 15209 7497 15243 7531
rect 16129 7497 16163 7531
rect 16773 7497 16807 7531
rect 16957 7497 16991 7531
rect 21465 7497 21499 7531
rect 23857 7497 23891 7531
rect 25973 7497 26007 7531
rect 26157 7497 26191 7531
rect 27445 7497 27479 7531
rect 29285 7497 29319 7531
rect 30389 7497 30423 7531
rect 30757 7497 30791 7531
rect 10333 7429 10367 7463
rect 22293 7429 22327 7463
rect 24685 7429 24719 7463
rect 2789 7361 2823 7395
rect 4537 7361 4571 7395
rect 5549 7361 5583 7395
rect 8953 7361 8987 7395
rect 10057 7361 10091 7395
rect 10241 7361 10275 7395
rect 20729 7361 20763 7395
rect 25421 7361 25455 7395
rect 26065 7361 26099 7395
rect 28089 7361 28123 7395
rect 29929 7361 29963 7395
rect 30021 7361 30055 7395
rect 1501 7293 1535 7327
rect 1777 7293 1811 7327
rect 1961 7293 1995 7327
rect 2053 7293 2087 7327
rect 2237 7293 2271 7327
rect 3893 7293 3927 7327
rect 3985 7293 4019 7327
rect 4169 7293 4203 7327
rect 4353 7293 4387 7327
rect 4445 7293 4479 7327
rect 4629 7293 4663 7327
rect 5273 7293 5307 7327
rect 5365 7293 5399 7327
rect 5457 7293 5491 7327
rect 6561 7293 6595 7327
rect 6837 7293 6871 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 8861 7293 8895 7327
rect 9045 7293 9079 7327
rect 9229 7293 9263 7327
rect 10425 7293 10459 7327
rect 12909 7293 12943 7327
rect 14657 7293 14691 7327
rect 14933 7293 14967 7327
rect 15117 7293 15151 7327
rect 15393 7293 15427 7327
rect 15485 7293 15519 7327
rect 15577 7293 15611 7327
rect 15669 7293 15703 7327
rect 16313 7293 16347 7327
rect 16405 7293 16439 7327
rect 16589 7293 16623 7327
rect 16681 7293 16715 7327
rect 20177 7293 20211 7327
rect 20269 7293 20303 7327
rect 20453 7293 20487 7327
rect 20545 7293 20579 7327
rect 21005 7293 21039 7327
rect 21189 7293 21223 7327
rect 21495 7293 21529 7327
rect 21649 7293 21683 7327
rect 21741 7293 21775 7327
rect 22109 7293 22143 7327
rect 22385 7293 22419 7327
rect 22569 7293 22603 7327
rect 22661 7293 22695 7327
rect 22845 7293 22879 7327
rect 22937 7293 22971 7327
rect 24133 7293 24167 7327
rect 24501 7293 24535 7327
rect 24593 7293 24627 7327
rect 25513 7293 25547 7327
rect 25605 7293 25639 7327
rect 25697 7293 25731 7327
rect 26985 7293 27019 7327
rect 27077 7293 27111 7327
rect 27261 7293 27295 7327
rect 27445 7293 27479 7327
rect 27537 7293 27571 7327
rect 28273 7293 28307 7327
rect 28549 7293 28583 7327
rect 29469 7293 29503 7327
rect 29561 7293 29595 7327
rect 30389 7293 30423 7327
rect 30665 7293 30699 7327
rect 25237 7259 25271 7293
rect 4077 7225 4111 7259
rect 17141 7225 17175 7259
rect 21097 7225 21131 7259
rect 21925 7225 21959 7259
rect 22017 7225 22051 7259
rect 24317 7225 24351 7259
rect 24869 7225 24903 7259
rect 27813 7225 27847 7259
rect 28457 7225 28491 7259
rect 4813 7157 4847 7191
rect 6653 7157 6687 7191
rect 12817 7157 12851 7191
rect 16941 7157 16975 7191
rect 24225 7157 24259 7191
rect 25329 7157 25363 7191
rect 25789 7157 25823 7191
rect 28733 7157 28767 7191
rect 30205 7157 30239 7191
rect 2053 6953 2087 6987
rect 5457 6953 5491 6987
rect 7665 6953 7699 6987
rect 15393 6953 15427 6987
rect 23673 6953 23707 6987
rect 24567 6953 24601 6987
rect 25513 6953 25547 6987
rect 2145 6885 2179 6919
rect 3985 6885 4019 6919
rect 10333 6885 10367 6919
rect 11989 6885 12023 6919
rect 18397 6885 18431 6919
rect 18613 6885 18647 6919
rect 24041 6885 24075 6919
rect 24777 6885 24811 6919
rect 25697 6885 25731 6919
rect 27813 6885 27847 6919
rect 1593 6817 1627 6851
rect 2421 6817 2455 6851
rect 3249 6817 3283 6851
rect 3617 6817 3651 6851
rect 3709 6817 3743 6851
rect 4077 6817 4111 6851
rect 4353 6817 4387 6851
rect 4721 6817 4755 6851
rect 4997 6817 5031 6851
rect 5365 6817 5399 6851
rect 6193 6817 6227 6851
rect 6285 6817 6319 6851
rect 6469 6817 6503 6851
rect 7021 6817 7055 6851
rect 7757 6817 7791 6851
rect 8309 6817 8343 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 8861 6817 8895 6851
rect 8953 6817 8987 6851
rect 9413 6817 9447 6851
rect 9597 6817 9631 6851
rect 10241 6817 10275 6851
rect 10425 6817 10459 6851
rect 10977 6817 11011 6851
rect 11253 6817 11287 6851
rect 11345 6817 11379 6851
rect 11805 6817 11839 6851
rect 12081 6817 12115 6851
rect 12633 6817 12667 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 13001 6817 13035 6851
rect 13277 6817 13311 6851
rect 14565 6817 14599 6851
rect 15025 6817 15059 6851
rect 16313 6817 16347 6851
rect 16497 6817 16531 6851
rect 16773 6817 16807 6851
rect 16865 6817 16899 6851
rect 17049 6817 17083 6851
rect 17141 6817 17175 6851
rect 17325 6817 17359 6851
rect 17509 6817 17543 6851
rect 17693 6817 17727 6851
rect 17877 6817 17911 6851
rect 18061 6817 18095 6851
rect 18153 6817 18187 6851
rect 18797 6817 18831 6851
rect 18981 6817 19015 6851
rect 19809 6817 19843 6851
rect 20269 6817 20303 6851
rect 20545 6817 20579 6851
rect 20729 6817 20763 6851
rect 21373 6817 21407 6851
rect 21557 6817 21591 6851
rect 22201 6817 22235 6851
rect 22293 6817 22327 6851
rect 22385 6817 22419 6851
rect 22569 6817 22603 6851
rect 23305 6817 23339 6851
rect 23489 6817 23523 6851
rect 23581 6817 23615 6851
rect 23857 6817 23891 6851
rect 23949 6817 23983 6851
rect 24225 6817 24259 6851
rect 24317 6817 24351 6851
rect 25145 6817 25179 6851
rect 25421 6817 25455 6851
rect 25881 6817 25915 6851
rect 27537 6817 27571 6851
rect 28549 6817 28583 6851
rect 28641 6817 28675 6851
rect 28825 6817 28859 6851
rect 29469 6817 29503 6851
rect 30113 6817 30147 6851
rect 30573 6817 30607 6851
rect 31125 6817 31159 6851
rect 1777 6749 1811 6783
rect 1869 6749 1903 6783
rect 2237 6749 2271 6783
rect 6929 6749 6963 6783
rect 8401 6749 8435 6783
rect 8769 6749 8803 6783
rect 9229 6749 9263 6783
rect 11529 6749 11563 6783
rect 12449 6749 12483 6783
rect 13553 6749 13587 6783
rect 15117 6749 15151 6783
rect 15301 6749 15335 6783
rect 15393 6749 15427 6783
rect 16681 6749 16715 6783
rect 17601 6749 17635 6783
rect 19993 6749 20027 6783
rect 20085 6749 20119 6783
rect 20177 6749 20211 6783
rect 21925 6749 21959 6783
rect 25053 6749 25087 6783
rect 27629 6749 27663 6783
rect 30021 6749 30055 6783
rect 2605 6681 2639 6715
rect 3893 6681 3927 6715
rect 11621 6681 11655 6715
rect 13461 6681 13495 6715
rect 17049 6681 17083 6715
rect 18981 6681 19015 6715
rect 20453 6681 20487 6715
rect 24409 6681 24443 6715
rect 29193 6681 29227 6715
rect 3709 6613 3743 6647
rect 9137 6613 9171 6647
rect 11069 6613 11103 6647
rect 13093 6613 13127 6647
rect 14657 6613 14691 6647
rect 18245 6613 18279 6647
rect 18429 6613 18463 6647
rect 20637 6613 20671 6647
rect 21373 6613 21407 6647
rect 21741 6613 21775 6647
rect 23305 6613 23339 6647
rect 24593 6613 24627 6647
rect 24961 6613 24995 6647
rect 25329 6613 25363 6647
rect 27353 6613 27387 6647
rect 27629 6613 27663 6647
rect 29009 6613 29043 6647
rect 1777 6409 1811 6443
rect 2881 6409 2915 6443
rect 2973 6409 3007 6443
rect 6653 6409 6687 6443
rect 7113 6409 7147 6443
rect 10609 6409 10643 6443
rect 14381 6409 14415 6443
rect 15485 6409 15519 6443
rect 16129 6409 16163 6443
rect 22109 6409 22143 6443
rect 24041 6409 24075 6443
rect 24409 6409 24443 6443
rect 25145 6409 25179 6443
rect 25513 6409 25547 6443
rect 27353 6409 27387 6443
rect 30389 6409 30423 6443
rect 4261 6341 4295 6375
rect 1409 6273 1443 6307
rect 3065 6273 3099 6307
rect 6745 6273 6779 6307
rect 7205 6273 7239 6307
rect 12817 6273 12851 6307
rect 12909 6273 12943 6307
rect 14473 6273 14507 6307
rect 14841 6273 14875 6307
rect 29009 6273 29043 6307
rect 29561 6273 29595 6307
rect 29653 6273 29687 6307
rect 29837 6273 29871 6307
rect 30021 6273 30055 6307
rect 30113 6273 30147 6307
rect 1593 6205 1627 6239
rect 2789 6205 2823 6239
rect 3249 6205 3283 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 3893 6205 3927 6239
rect 5273 6205 5307 6239
rect 5549 6205 5583 6239
rect 6929 6205 6963 6239
rect 7389 6205 7423 6239
rect 7665 6205 7699 6239
rect 7849 6205 7883 6239
rect 10241 6205 10275 6239
rect 10333 6205 10367 6239
rect 10701 6205 10735 6239
rect 12633 6205 12667 6239
rect 13093 6205 13127 6239
rect 13277 6205 13311 6239
rect 13829 6205 13863 6239
rect 13921 6205 13955 6239
rect 14105 6205 14139 6239
rect 14197 6205 14231 6239
rect 14657 6205 14691 6239
rect 14749 6205 14783 6239
rect 14933 6205 14967 6239
rect 15301 6205 15335 6239
rect 16313 6205 16347 6239
rect 16497 6205 16531 6239
rect 16589 6205 16623 6239
rect 19257 6205 19291 6239
rect 19533 6205 19567 6239
rect 21925 6205 21959 6239
rect 22109 6205 22143 6239
rect 24317 6205 24351 6239
rect 24501 6205 24535 6239
rect 25053 6205 25087 6239
rect 25237 6205 25271 6239
rect 25697 6205 25731 6239
rect 25789 6205 25823 6239
rect 27169 6205 27203 6239
rect 27353 6205 27387 6239
rect 29193 6205 29227 6239
rect 29929 6205 29963 6239
rect 30297 6205 30331 6239
rect 30481 6205 30515 6239
rect 4077 6137 4111 6171
rect 5457 6137 5491 6171
rect 6009 6137 6043 6171
rect 6653 6137 6687 6171
rect 12449 6137 12483 6171
rect 15117 6137 15151 6171
rect 24225 6137 24259 6171
rect 5089 6069 5123 6103
rect 5733 6069 5767 6103
rect 10425 6069 10459 6103
rect 10701 6069 10735 6103
rect 13277 6069 13311 6103
rect 19073 6069 19107 6103
rect 19441 6069 19475 6103
rect 23857 6069 23891 6103
rect 24025 6069 24059 6103
rect 29193 6069 29227 6103
rect 1409 5865 1443 5899
rect 4629 5865 4663 5899
rect 4813 5865 4847 5899
rect 6285 5865 6319 5899
rect 8861 5865 8895 5899
rect 9689 5865 9723 5899
rect 17417 5865 17451 5899
rect 18337 5865 18371 5899
rect 19257 5865 19291 5899
rect 20269 5865 20303 5899
rect 21373 5865 21407 5899
rect 23765 5865 23799 5899
rect 27077 5865 27111 5899
rect 28917 5865 28951 5899
rect 29653 5865 29687 5899
rect 1961 5797 1995 5831
rect 2329 5797 2363 5831
rect 6561 5797 6595 5831
rect 8769 5797 8803 5831
rect 9137 5797 9171 5831
rect 9229 5797 9263 5831
rect 11621 5797 11655 5831
rect 11805 5797 11839 5831
rect 26617 5797 26651 5831
rect 26985 5797 27019 5831
rect 1317 5729 1351 5763
rect 1501 5729 1535 5763
rect 1869 5729 1903 5763
rect 3065 5729 3099 5763
rect 3341 5729 3375 5763
rect 3985 5729 4019 5763
rect 4810 5729 4844 5763
rect 5181 5729 5215 5763
rect 5273 5729 5307 5763
rect 6285 5729 6319 5763
rect 6377 5729 6411 5763
rect 7573 5729 7607 5763
rect 8493 5729 8527 5763
rect 8585 5729 8619 5763
rect 9040 5729 9074 5763
rect 9412 5729 9446 5763
rect 9505 5729 9539 5763
rect 9597 5729 9631 5763
rect 9965 5729 9999 5763
rect 11161 5729 11195 5763
rect 11253 5729 11287 5763
rect 11437 5729 11471 5763
rect 11529 5729 11563 5763
rect 16497 5729 16531 5763
rect 16681 5729 16715 5763
rect 16773 5729 16807 5763
rect 17601 5729 17635 5763
rect 17693 5729 17727 5763
rect 17969 5729 18003 5763
rect 18245 5729 18279 5763
rect 18429 5729 18463 5763
rect 18521 5729 18555 5763
rect 18705 5729 18739 5763
rect 19533 5729 19567 5763
rect 19809 5729 19843 5763
rect 19901 5729 19935 5763
rect 20085 5729 20119 5763
rect 20361 5729 20395 5763
rect 21557 5729 21591 5763
rect 21833 5729 21867 5763
rect 22017 5729 22051 5763
rect 22201 5729 22235 5763
rect 22385 5729 22419 5763
rect 22569 5729 22603 5763
rect 24133 5729 24167 5763
rect 25513 5729 25547 5763
rect 25789 5729 25823 5763
rect 25973 5729 26007 5763
rect 26893 5729 26927 5763
rect 27261 5729 27295 5763
rect 28457 5729 28491 5763
rect 28733 5729 28767 5763
rect 29414 5729 29448 5763
rect 29561 5729 29595 5763
rect 29653 5729 29687 5763
rect 29837 5729 29871 5763
rect 2053 5661 2087 5695
rect 4077 5661 4111 5695
rect 7849 5661 7883 5695
rect 10149 5661 10183 5695
rect 10977 5661 11011 5695
rect 11989 5661 12023 5695
rect 17877 5661 17911 5695
rect 18613 5661 18647 5695
rect 21649 5661 21683 5695
rect 22109 5661 22143 5695
rect 24041 5661 24075 5695
rect 25421 5661 25455 5695
rect 27353 5661 27387 5695
rect 28089 5661 28123 5695
rect 29193 5661 29227 5695
rect 2513 5593 2547 5627
rect 4353 5593 4387 5627
rect 8769 5593 8803 5627
rect 21741 5593 21775 5627
rect 28641 5593 28675 5627
rect 29285 5593 29319 5627
rect 16313 5525 16347 5559
rect 19441 5525 19475 5559
rect 22477 5525 22511 5559
rect 23949 5525 23983 5559
rect 25973 5525 26007 5559
rect 5917 5321 5951 5355
rect 12541 5321 12575 5355
rect 13553 5321 13587 5355
rect 17325 5321 17359 5355
rect 19073 5321 19107 5355
rect 21465 5321 21499 5355
rect 23949 5321 23983 5355
rect 25605 5321 25639 5355
rect 26617 5321 26651 5355
rect 29009 5321 29043 5355
rect 2513 5253 2547 5287
rect 7849 5253 7883 5287
rect 14933 5253 14967 5287
rect 15945 5253 15979 5287
rect 24133 5253 24167 5287
rect 26433 5253 26467 5287
rect 3617 5185 3651 5219
rect 11805 5185 11839 5219
rect 11897 5185 11931 5219
rect 11989 5185 12023 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 14105 5185 14139 5219
rect 23213 5185 23247 5219
rect 23581 5185 23615 5219
rect 26157 5185 26191 5219
rect 27997 5185 28031 5219
rect 1869 5117 1903 5151
rect 2789 5117 2823 5151
rect 3341 5117 3375 5151
rect 3525 5117 3559 5151
rect 6101 5117 6135 5151
rect 6285 5117 6319 5151
rect 6377 5117 6411 5151
rect 6469 5117 6503 5151
rect 6653 5117 6687 5151
rect 7389 5117 7423 5151
rect 7573 5117 7607 5151
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 12081 5117 12115 5151
rect 12725 5117 12759 5151
rect 13678 5117 13712 5151
rect 14197 5117 14231 5151
rect 14749 5117 14783 5151
rect 14841 5117 14875 5151
rect 15209 5117 15243 5151
rect 15301 5117 15335 5151
rect 15393 5117 15427 5151
rect 15761 5117 15795 5151
rect 16037 5117 16071 5151
rect 16221 5117 16255 5151
rect 17049 5117 17083 5151
rect 17141 5117 17175 5151
rect 18705 5117 18739 5151
rect 18797 5117 18831 5151
rect 18981 5117 19015 5151
rect 19073 5117 19107 5151
rect 20637 5117 20671 5151
rect 20729 5117 20763 5151
rect 20913 5117 20947 5151
rect 21097 5117 21131 5151
rect 21189 5117 21223 5151
rect 21465 5117 21499 5151
rect 23397 5117 23431 5151
rect 23673 5117 23707 5151
rect 24409 5117 24443 5151
rect 24777 5117 24811 5151
rect 25053 5117 25087 5151
rect 25421 5117 25455 5151
rect 25605 5117 25639 5151
rect 26709 5117 26743 5151
rect 27353 5117 27387 5151
rect 27721 5117 27755 5151
rect 28549 5117 28583 5151
rect 29285 5117 29319 5151
rect 29377 5117 29411 5151
rect 29745 5117 29779 5151
rect 30205 5117 30239 5151
rect 30849 5117 30883 5151
rect 14473 5049 14507 5083
rect 15577 5049 15611 5083
rect 15669 5049 15703 5083
rect 17325 5049 17359 5083
rect 7389 4981 7423 5015
rect 11621 4981 11655 5015
rect 13737 4981 13771 5015
rect 15117 4981 15151 5015
rect 16129 4981 16163 5015
rect 21281 4981 21315 5015
rect 24593 4981 24627 5015
rect 24961 4981 24995 5015
rect 25237 4981 25271 5015
rect 28549 4981 28583 5015
rect 2421 4777 2455 4811
rect 3249 4777 3283 4811
rect 3985 4777 4019 4811
rect 4997 4777 5031 4811
rect 5825 4777 5859 4811
rect 17233 4777 17267 4811
rect 18705 4777 18739 4811
rect 19441 4777 19475 4811
rect 22385 4777 22419 4811
rect 25053 4777 25087 4811
rect 29377 4777 29411 4811
rect 2053 4709 2087 4743
rect 3617 4709 3651 4743
rect 18521 4709 18555 4743
rect 20361 4709 20395 4743
rect 1869 4641 1903 4675
rect 2421 4641 2455 4675
rect 2605 4641 2639 4675
rect 3433 4641 3467 4675
rect 3525 4641 3559 4675
rect 3801 4641 3835 4675
rect 4353 4641 4387 4675
rect 4905 4641 4939 4675
rect 5089 4641 5123 4675
rect 6009 4641 6043 4675
rect 6377 4641 6411 4675
rect 6561 4641 6595 4675
rect 7389 4641 7423 4675
rect 7757 4641 7791 4675
rect 8217 4641 8251 4675
rect 9505 4641 9539 4675
rect 9597 4641 9631 4675
rect 9781 4641 9815 4675
rect 10333 4641 10367 4675
rect 11713 4641 11747 4675
rect 15577 4641 15611 4675
rect 15761 4641 15795 4675
rect 16497 4641 16531 4675
rect 16681 4641 16715 4675
rect 18061 4641 18095 4675
rect 18245 4641 18279 4675
rect 18337 4641 18371 4675
rect 18797 4641 18831 4675
rect 18981 4641 19015 4675
rect 19073 4641 19107 4675
rect 19165 4641 19199 4675
rect 20575 4641 20609 4675
rect 20729 4641 20763 4675
rect 22661 4641 22695 4675
rect 22753 4641 22787 4675
rect 22845 4641 22879 4675
rect 23029 4641 23063 4675
rect 25053 4641 25087 4675
rect 25237 4641 25271 4675
rect 26801 4641 26835 4675
rect 27445 4641 27479 4675
rect 29469 4641 29503 4675
rect 2145 4573 2179 4607
rect 4261 4573 4295 4607
rect 6193 4573 6227 4607
rect 6285 4573 6319 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 10057 4573 10091 4607
rect 10241 4573 10275 4607
rect 10425 4573 10459 4607
rect 10517 4573 10551 4607
rect 11805 4573 11839 4607
rect 11897 4573 11931 4607
rect 11989 4573 12023 4607
rect 16773 4573 16807 4607
rect 16865 4573 16899 4607
rect 18153 4573 18187 4607
rect 26709 4573 26743 4607
rect 8033 4437 8067 4471
rect 9965 4437 9999 4471
rect 11529 4437 11563 4471
rect 16957 4437 16991 4471
rect 7941 4233 7975 4267
rect 8493 4233 8527 4267
rect 9965 4233 9999 4267
rect 10241 4233 10275 4267
rect 12633 4233 12667 4267
rect 15945 4233 15979 4267
rect 20453 4233 20487 4267
rect 22661 4233 22695 4267
rect 24777 4233 24811 4267
rect 8953 4165 8987 4199
rect 17509 4165 17543 4199
rect 21189 4165 21223 4199
rect 25237 4165 25271 4199
rect 5365 4097 5399 4131
rect 6929 4097 6963 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 9873 4097 9907 4131
rect 11253 4097 11287 4131
rect 11345 4097 11379 4131
rect 13093 4097 13127 4131
rect 13553 4097 13587 4131
rect 19809 4097 19843 4131
rect 20637 4097 20671 4131
rect 22753 4097 22787 4131
rect 24133 4097 24167 4131
rect 25973 4097 26007 4131
rect 3801 4029 3835 4063
rect 4169 4029 4203 4063
rect 5181 4029 5215 4063
rect 6561 4029 6595 4063
rect 7113 4029 7147 4063
rect 7573 4029 7607 4063
rect 8033 4029 8067 4063
rect 8401 4029 8435 4063
rect 9045 4029 9079 4063
rect 9781 4029 9815 4063
rect 10425 4029 10459 4063
rect 10517 4029 10551 4063
rect 10609 4029 10643 4063
rect 10701 4029 10735 4063
rect 11161 4029 11195 4063
rect 11437 4029 11471 4063
rect 12817 4029 12851 4063
rect 13001 4029 13035 4063
rect 13645 4029 13679 4063
rect 13829 4029 13863 4063
rect 14565 4029 14599 4063
rect 14749 4029 14783 4063
rect 14933 4029 14967 4063
rect 15301 4029 15335 4063
rect 15485 4029 15519 4063
rect 15761 4029 15795 4063
rect 15945 4029 15979 4063
rect 17784 4029 17818 4063
rect 17877 4029 17911 4063
rect 19717 4029 19751 4063
rect 19901 4029 19935 4063
rect 19993 4029 20027 4063
rect 20177 4029 20211 4063
rect 21648 4029 21682 4063
rect 21741 4029 21775 4063
rect 21833 4029 21867 4063
rect 22017 4029 22051 4063
rect 22385 4029 22419 4063
rect 22937 4029 22971 4063
rect 23029 4029 23063 4063
rect 23213 4029 23247 4063
rect 23305 4029 23339 4063
rect 24409 4029 24443 4063
rect 24869 4029 24903 4063
rect 25329 4029 25363 4063
rect 25881 4029 25915 4063
rect 4997 3961 5031 3995
rect 8677 3961 8711 3995
rect 8769 3961 8803 3995
rect 15669 3961 15703 3995
rect 19165 3961 19199 3995
rect 19349 3961 19383 3995
rect 19533 3961 19567 3995
rect 20361 3961 20395 3995
rect 21189 3961 21223 3995
rect 21373 3961 21407 3995
rect 22661 3961 22695 3995
rect 24501 3961 24535 3995
rect 4077 3893 4111 3927
rect 10149 3893 10183 3927
rect 11621 3893 11655 3927
rect 20729 3893 20763 3927
rect 22477 3893 22511 3927
rect 24593 3893 24627 3927
rect 3525 3689 3559 3723
rect 14657 3689 14691 3723
rect 3157 3621 3191 3655
rect 8493 3621 8527 3655
rect 10793 3621 10827 3655
rect 3249 3553 3283 3587
rect 3433 3553 3467 3587
rect 3525 3553 3559 3587
rect 6653 3553 6687 3587
rect 7021 3553 7055 3587
rect 10517 3553 10551 3587
rect 10609 3553 10643 3587
rect 12909 3553 12943 3587
rect 13001 3553 13035 3587
rect 13737 3553 13771 3587
rect 13921 3553 13955 3587
rect 14289 3553 14323 3587
rect 14382 3553 14416 3587
rect 14105 3417 14139 3451
rect 3341 3349 3375 3383
rect 10517 3349 10551 3383
<< metal1 >>
rect 11974 21972 11980 22024
rect 12032 22012 12038 22024
rect 26878 22012 26884 22024
rect 12032 21984 26884 22012
rect 12032 21972 12038 21984
rect 26878 21972 26884 21984
rect 26936 21972 26942 22024
rect 13814 21904 13820 21956
rect 13872 21944 13878 21956
rect 26234 21944 26240 21956
rect 13872 21916 26240 21944
rect 13872 21904 13878 21916
rect 26234 21904 26240 21916
rect 26292 21904 26298 21956
rect 27982 21904 27988 21956
rect 28040 21944 28046 21956
rect 30926 21944 30932 21956
rect 28040 21916 30932 21944
rect 28040 21904 28046 21916
rect 30926 21904 30932 21916
rect 30984 21904 30990 21956
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 18782 21876 18788 21888
rect 9180 21848 18788 21876
rect 9180 21836 9186 21848
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 24762 21836 24768 21888
rect 24820 21876 24826 21888
rect 27522 21876 27528 21888
rect 24820 21848 27528 21876
rect 24820 21836 24826 21848
rect 27522 21836 27528 21848
rect 27580 21876 27586 21888
rect 30282 21876 30288 21888
rect 27580 21848 30288 21876
rect 27580 21836 27586 21848
rect 30282 21836 30288 21848
rect 30340 21836 30346 21888
rect 552 21786 31648 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 11436 21786
rect 11488 21734 11500 21786
rect 11552 21734 11564 21786
rect 11616 21734 11628 21786
rect 11680 21734 11692 21786
rect 11744 21734 19210 21786
rect 19262 21734 19274 21786
rect 19326 21734 19338 21786
rect 19390 21734 19402 21786
rect 19454 21734 19466 21786
rect 19518 21734 26984 21786
rect 27036 21734 27048 21786
rect 27100 21734 27112 21786
rect 27164 21734 27176 21786
rect 27228 21734 27240 21786
rect 27292 21734 31648 21786
rect 552 21712 31648 21734
rect 6178 21632 6184 21684
rect 6236 21632 6242 21684
rect 6730 21632 6736 21684
rect 6788 21632 6794 21684
rect 7282 21632 7288 21684
rect 7340 21632 7346 21684
rect 7834 21632 7840 21684
rect 7892 21632 7898 21684
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 9490 21632 9496 21684
rect 9548 21632 9554 21684
rect 9582 21632 9588 21684
rect 9640 21672 9646 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 9640 21644 9781 21672
rect 9640 21632 9646 21644
rect 9769 21641 9781 21644
rect 9815 21641 9827 21675
rect 9769 21635 9827 21641
rect 10042 21632 10048 21684
rect 10100 21632 10106 21684
rect 10594 21632 10600 21684
rect 10652 21632 10658 21684
rect 11146 21632 11152 21684
rect 11204 21632 11210 21684
rect 11422 21632 11428 21684
rect 11480 21672 11486 21684
rect 11609 21675 11667 21681
rect 11609 21672 11621 21675
rect 11480 21644 11621 21672
rect 11480 21632 11486 21644
rect 11609 21641 11621 21644
rect 11655 21641 11667 21675
rect 11609 21635 11667 21641
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12250 21632 12256 21684
rect 12308 21632 12314 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 13354 21632 13360 21684
rect 13412 21632 13418 21684
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 16301 21675 16359 21681
rect 16301 21641 16313 21675
rect 16347 21672 16359 21675
rect 16666 21672 16672 21684
rect 16347 21644 16672 21672
rect 16347 21641 16359 21644
rect 16301 21635 16359 21641
rect 16666 21632 16672 21644
rect 16724 21632 16730 21684
rect 20901 21675 20959 21681
rect 20901 21641 20913 21675
rect 20947 21672 20959 21675
rect 22278 21672 22284 21684
rect 20947 21644 22284 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 23106 21632 23112 21684
rect 23164 21632 23170 21684
rect 25685 21675 25743 21681
rect 25685 21641 25697 21675
rect 25731 21672 25743 21675
rect 26418 21672 26424 21684
rect 25731 21644 26424 21672
rect 25731 21641 25743 21644
rect 25685 21635 25743 21641
rect 26418 21632 26424 21644
rect 26476 21632 26482 21684
rect 28813 21675 28871 21681
rect 28813 21672 28825 21675
rect 26528 21644 28825 21672
rect 10778 21564 10784 21616
rect 10836 21604 10842 21616
rect 13814 21604 13820 21616
rect 10836 21576 13820 21604
rect 10836 21564 10842 21576
rect 13814 21564 13820 21576
rect 13872 21564 13878 21616
rect 20717 21607 20775 21613
rect 20717 21573 20729 21607
rect 20763 21604 20775 21607
rect 21174 21604 21180 21616
rect 20763 21576 21180 21604
rect 20763 21573 20775 21576
rect 20717 21567 20775 21573
rect 21174 21564 21180 21576
rect 21232 21564 21238 21616
rect 25222 21564 25228 21616
rect 25280 21604 25286 21616
rect 26528 21604 26556 21644
rect 28813 21641 28825 21644
rect 28859 21672 28871 21675
rect 28859 21644 31340 21672
rect 28859 21641 28871 21644
rect 28813 21635 28871 21641
rect 25280 21576 26556 21604
rect 28169 21607 28227 21613
rect 25280 21564 25286 21576
rect 28169 21573 28181 21607
rect 28215 21604 28227 21607
rect 28350 21604 28356 21616
rect 28215 21576 28356 21604
rect 28215 21573 28227 21576
rect 28169 21567 28227 21573
rect 28350 21564 28356 21576
rect 28408 21564 28414 21616
rect 28920 21576 29040 21604
rect 11330 21496 11336 21548
rect 11388 21536 11394 21548
rect 14001 21539 14059 21545
rect 14001 21536 14013 21539
rect 11388 21508 14013 21536
rect 11388 21496 11394 21508
rect 14001 21505 14013 21508
rect 14047 21536 14059 21539
rect 14642 21536 14648 21548
rect 14047 21508 14648 21536
rect 14047 21505 14059 21508
rect 14001 21499 14059 21505
rect 14642 21496 14648 21508
rect 14700 21496 14706 21548
rect 14734 21496 14740 21548
rect 14792 21536 14798 21548
rect 17218 21536 17224 21548
rect 14792 21508 17224 21536
rect 14792 21496 14798 21508
rect 17218 21496 17224 21508
rect 17276 21536 17282 21548
rect 17276 21508 17816 21536
rect 17276 21496 17282 21508
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 9950 21468 9956 21480
rect 9447 21440 9956 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 9950 21428 9956 21440
rect 10008 21428 10014 21480
rect 16390 21428 16396 21480
rect 16448 21428 16454 21480
rect 17788 21454 17816 21508
rect 18414 21496 18420 21548
rect 18472 21496 18478 21548
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 19426 21536 19432 21548
rect 18739 21508 19432 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 21315 21508 23980 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 22922 21468 22928 21480
rect 20364 21440 21220 21468
rect 22678 21440 22928 21468
rect 11333 21403 11391 21409
rect 11333 21369 11345 21403
rect 11379 21400 11391 21403
rect 11425 21403 11483 21409
rect 11425 21400 11437 21403
rect 11379 21372 11437 21400
rect 11379 21369 11391 21372
rect 11333 21363 11391 21369
rect 11425 21369 11437 21372
rect 11471 21400 11483 21403
rect 11471 21372 12434 21400
rect 11471 21369 11483 21372
rect 11425 21363 11483 21369
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 8757 21335 8815 21341
rect 8757 21332 8769 21335
rect 7892 21304 8769 21332
rect 7892 21292 7898 21304
rect 8757 21301 8769 21304
rect 8803 21332 8815 21335
rect 9030 21332 9036 21344
rect 8803 21304 9036 21332
rect 8803 21301 8815 21304
rect 8757 21295 8815 21301
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 10594 21292 10600 21344
rect 10652 21332 10658 21344
rect 11625 21335 11683 21341
rect 11625 21332 11637 21335
rect 10652 21304 11637 21332
rect 10652 21292 10658 21304
rect 11625 21301 11637 21304
rect 11671 21301 11683 21335
rect 11625 21295 11683 21301
rect 11790 21292 11796 21344
rect 11848 21292 11854 21344
rect 12406 21332 12434 21372
rect 14274 21360 14280 21412
rect 14332 21360 14338 21412
rect 14734 21360 14740 21412
rect 14792 21360 14798 21412
rect 16669 21403 16727 21409
rect 15580 21372 16620 21400
rect 15580 21332 15608 21372
rect 12406 21304 15608 21332
rect 15749 21335 15807 21341
rect 15749 21301 15761 21335
rect 15795 21332 15807 21335
rect 16114 21332 16120 21344
rect 15795 21304 16120 21332
rect 15795 21301 15807 21304
rect 15749 21295 15807 21301
rect 16114 21292 16120 21304
rect 16172 21292 16178 21344
rect 16592 21332 16620 21372
rect 16669 21369 16681 21403
rect 16715 21400 16727 21403
rect 16758 21400 16764 21412
rect 16715 21372 16764 21400
rect 16715 21369 16727 21372
rect 16669 21363 16727 21369
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 18966 21360 18972 21412
rect 19024 21360 19030 21412
rect 20254 21400 20260 21412
rect 20194 21372 20260 21400
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 17310 21332 17316 21344
rect 16592 21304 17316 21332
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 18322 21292 18328 21344
rect 18380 21332 18386 21344
rect 20364 21332 20392 21440
rect 20622 21400 20628 21412
rect 20456 21372 20628 21400
rect 20456 21341 20484 21372
rect 20622 21360 20628 21372
rect 20680 21400 20686 21412
rect 20680 21372 21036 21400
rect 20680 21360 20686 21372
rect 20898 21341 20904 21344
rect 18380 21304 20392 21332
rect 20441 21335 20499 21341
rect 18380 21292 18386 21304
rect 20441 21301 20453 21335
rect 20487 21301 20499 21335
rect 20441 21295 20499 21301
rect 20885 21335 20904 21341
rect 20885 21301 20897 21335
rect 20885 21295 20904 21301
rect 20898 21292 20904 21295
rect 20956 21292 20962 21344
rect 21008 21332 21036 21372
rect 21082 21360 21088 21412
rect 21140 21360 21146 21412
rect 21192 21400 21220 21440
rect 22922 21428 22928 21440
rect 22980 21428 22986 21480
rect 23014 21428 23020 21480
rect 23072 21468 23078 21480
rect 23952 21477 23980 21508
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 25869 21539 25927 21545
rect 25869 21536 25881 21539
rect 24912 21508 25881 21536
rect 24912 21496 24918 21508
rect 25869 21505 25881 21508
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 26326 21496 26332 21548
rect 26384 21536 26390 21548
rect 26421 21539 26479 21545
rect 26421 21536 26433 21539
rect 26384 21508 26433 21536
rect 26384 21496 26390 21508
rect 26421 21505 26433 21508
rect 26467 21536 26479 21539
rect 28920 21536 28948 21576
rect 29012 21545 29040 21576
rect 26467 21508 28948 21536
rect 26467 21505 26479 21508
rect 26421 21499 26479 21505
rect 23109 21471 23167 21477
rect 23109 21468 23121 21471
rect 23072 21440 23121 21468
rect 23072 21428 23078 21440
rect 23109 21437 23121 21440
rect 23155 21437 23167 21471
rect 23109 21431 23167 21437
rect 23201 21471 23259 21477
rect 23201 21437 23213 21471
rect 23247 21437 23259 21471
rect 23201 21431 23259 21437
rect 23937 21471 23995 21477
rect 23937 21437 23949 21471
rect 23983 21437 23995 21471
rect 26050 21468 26056 21480
rect 25346 21440 26056 21468
rect 23937 21431 23995 21437
rect 21545 21403 21603 21409
rect 21545 21400 21557 21403
rect 21192 21372 21557 21400
rect 21545 21369 21557 21372
rect 21591 21369 21603 21403
rect 23216 21400 23244 21431
rect 21545 21363 21603 21369
rect 22848 21372 23244 21400
rect 23952 21400 23980 21431
rect 26050 21428 26056 21440
rect 26108 21428 26114 21480
rect 24118 21400 24124 21412
rect 23952 21372 24124 21400
rect 22848 21332 22876 21372
rect 24118 21360 24124 21372
rect 24176 21360 24182 21412
rect 24210 21360 24216 21412
rect 24268 21360 24274 21412
rect 25516 21372 26004 21400
rect 21008 21304 22876 21332
rect 23017 21335 23075 21341
rect 23017 21301 23029 21335
rect 23063 21332 23075 21335
rect 23106 21332 23112 21344
rect 23063 21304 23112 21332
rect 23063 21301 23075 21304
rect 23017 21295 23075 21301
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 24026 21332 24032 21344
rect 23523 21304 24032 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24302 21292 24308 21344
rect 24360 21332 24366 21344
rect 25516 21332 25544 21372
rect 24360 21304 25544 21332
rect 25976 21332 26004 21372
rect 26142 21360 26148 21412
rect 26200 21360 26206 21412
rect 26697 21403 26755 21409
rect 26697 21369 26709 21403
rect 26743 21369 26755 21403
rect 27982 21400 27988 21412
rect 27922 21372 27988 21400
rect 26697 21363 26755 21369
rect 26602 21332 26608 21344
rect 25976 21304 26608 21332
rect 24360 21292 24366 21304
rect 26602 21292 26608 21304
rect 26660 21292 26666 21344
rect 26719 21332 26747 21363
rect 27982 21360 27988 21372
rect 28040 21360 28046 21412
rect 28258 21360 28264 21412
rect 28316 21360 28322 21412
rect 28074 21332 28080 21344
rect 26719 21304 28080 21332
rect 28074 21292 28080 21304
rect 28132 21292 28138 21344
rect 28166 21292 28172 21344
rect 28224 21332 28230 21344
rect 28445 21335 28503 21341
rect 28445 21332 28457 21335
rect 28224 21304 28457 21332
rect 28224 21292 28230 21304
rect 28445 21301 28457 21304
rect 28491 21301 28503 21335
rect 28445 21295 28503 21301
rect 28534 21292 28540 21344
rect 28592 21292 28598 21344
rect 28626 21292 28632 21344
rect 28684 21292 28690 21344
rect 28920 21332 28948 21508
rect 28997 21539 29055 21545
rect 28997 21505 29009 21539
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 31021 21471 31079 21477
rect 31021 21437 31033 21471
rect 31067 21468 31079 21471
rect 31202 21468 31208 21480
rect 31067 21440 31208 21468
rect 31067 21437 31079 21440
rect 31021 21431 31079 21437
rect 31202 21428 31208 21440
rect 31260 21428 31266 21480
rect 31312 21477 31340 21644
rect 31297 21471 31355 21477
rect 31297 21437 31309 21471
rect 31343 21468 31355 21471
rect 31386 21468 31392 21480
rect 31343 21440 31392 21468
rect 31343 21437 31355 21440
rect 31297 21431 31355 21437
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 29273 21403 29331 21409
rect 29273 21369 29285 21403
rect 29319 21400 29331 21403
rect 29362 21400 29368 21412
rect 29319 21372 29368 21400
rect 29319 21369 29331 21372
rect 29273 21363 29331 21369
rect 29362 21360 29368 21372
rect 29420 21360 29426 21412
rect 30558 21400 30564 21412
rect 30498 21372 30564 21400
rect 30558 21360 30564 21372
rect 30616 21360 30622 21412
rect 30760 21372 31248 21400
rect 28994 21332 29000 21344
rect 28920 21304 29000 21332
rect 28994 21292 29000 21304
rect 29052 21292 29058 21344
rect 30190 21292 30196 21344
rect 30248 21332 30254 21344
rect 30760 21341 30788 21372
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30248 21304 30757 21332
rect 30248 21292 30254 21304
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 30745 21295 30803 21301
rect 30834 21292 30840 21344
rect 30892 21292 30898 21344
rect 31220 21341 31248 21372
rect 31205 21335 31263 21341
rect 31205 21301 31217 21335
rect 31251 21301 31263 21335
rect 31205 21295 31263 21301
rect 552 21242 31648 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 12096 21242
rect 12148 21190 12160 21242
rect 12212 21190 12224 21242
rect 12276 21190 12288 21242
rect 12340 21190 12352 21242
rect 12404 21190 19870 21242
rect 19922 21190 19934 21242
rect 19986 21190 19998 21242
rect 20050 21190 20062 21242
rect 20114 21190 20126 21242
rect 20178 21190 27644 21242
rect 27696 21190 27708 21242
rect 27760 21190 27772 21242
rect 27824 21190 27836 21242
rect 27888 21190 27900 21242
rect 27952 21190 31648 21242
rect 552 21168 31648 21190
rect 10594 21088 10600 21140
rect 10652 21088 10658 21140
rect 11057 21131 11115 21137
rect 10704 21100 11008 21128
rect 7745 21063 7803 21069
rect 7745 21029 7757 21063
rect 7791 21060 7803 21063
rect 8205 21063 8263 21069
rect 8205 21060 8217 21063
rect 7791 21032 8217 21060
rect 7791 21029 7803 21032
rect 7745 21023 7803 21029
rect 8205 21029 8217 21032
rect 8251 21029 8263 21063
rect 9582 21060 9588 21072
rect 9430 21032 9588 21060
rect 8205 21023 8263 21029
rect 9582 21020 9588 21032
rect 9640 21060 9646 21072
rect 10704 21060 10732 21100
rect 9640 21032 10732 21060
rect 10980 21060 11008 21100
rect 11057 21097 11069 21131
rect 11103 21128 11115 21131
rect 11238 21128 11244 21140
rect 11103 21100 11244 21128
rect 11103 21097 11115 21100
rect 11057 21091 11115 21097
rect 11238 21088 11244 21100
rect 11296 21088 11302 21140
rect 11422 21088 11428 21140
rect 11480 21088 11486 21140
rect 11716 21100 14228 21128
rect 11716 21060 11744 21100
rect 9640 21020 9646 21032
rect 10781 21029 10839 21035
rect 10980 21032 11744 21060
rect 7650 20952 7656 21004
rect 7708 20952 7714 21004
rect 7834 20952 7840 21004
rect 7892 20952 7898 21004
rect 10505 20995 10563 21001
rect 10505 20961 10517 20995
rect 10551 20961 10563 20995
rect 10505 20955 10563 20961
rect 7190 20884 7196 20936
rect 7248 20924 7254 20936
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7248 20896 7941 20924
rect 7248 20884 7254 20896
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 9950 20924 9956 20936
rect 9723 20896 9956 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 9950 20884 9956 20896
rect 10008 20924 10014 20936
rect 10520 20924 10548 20955
rect 10594 20952 10600 21004
rect 10652 20952 10658 21004
rect 10781 20995 10793 21029
rect 10827 21026 10839 21029
rect 10827 20998 10916 21026
rect 11790 21020 11796 21072
rect 11848 21020 11854 21072
rect 12176 21060 12204 21100
rect 14200 21060 14228 21100
rect 14274 21088 14280 21140
rect 14332 21088 14338 21140
rect 16758 21088 16764 21140
rect 16816 21088 16822 21140
rect 17310 21088 17316 21140
rect 17368 21128 17374 21140
rect 21910 21128 21916 21140
rect 17368 21100 21916 21128
rect 17368 21088 17374 21100
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 23106 21128 23112 21140
rect 22066 21100 23112 21128
rect 14734 21060 14740 21072
rect 12176 21032 12282 21060
rect 14200 21032 14740 21060
rect 14734 21020 14740 21032
rect 14792 21020 14798 21072
rect 16482 21060 16488 21072
rect 14844 21032 16488 21060
rect 10827 20995 10839 20998
rect 10781 20989 10839 20995
rect 10008 20896 10548 20924
rect 10888 20924 10916 20998
rect 10962 20952 10968 21004
rect 11020 20952 11026 21004
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11256 20924 11284 20955
rect 13078 20952 13084 21004
rect 13136 20992 13142 21004
rect 13633 20995 13691 21001
rect 13633 20992 13645 20995
rect 13136 20964 13645 20992
rect 13136 20952 13142 20964
rect 13633 20961 13645 20964
rect 13679 20961 13691 20995
rect 13633 20955 13691 20961
rect 13817 20995 13875 21001
rect 13817 20961 13829 20995
rect 13863 20961 13875 20995
rect 13817 20955 13875 20961
rect 10888 20896 11284 20924
rect 10008 20884 10014 20896
rect 10520 20856 10548 20896
rect 11146 20856 11152 20868
rect 10520 20828 11152 20856
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 10594 20748 10600 20800
rect 10652 20788 10658 20800
rect 10962 20788 10968 20800
rect 10652 20760 10968 20788
rect 10652 20748 10658 20760
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 11256 20788 11284 20896
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 11517 20927 11575 20933
rect 11517 20924 11529 20927
rect 11388 20896 11529 20924
rect 11388 20884 11394 20896
rect 11517 20893 11529 20896
rect 11563 20893 11575 20927
rect 11517 20887 11575 20893
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 13832 20924 13860 20955
rect 14090 20952 14096 21004
rect 14148 20952 14154 21004
rect 14844 21001 14872 21032
rect 16482 21020 16488 21032
rect 16540 21020 16546 21072
rect 17218 21020 17224 21072
rect 17276 21060 17282 21072
rect 18138 21060 18144 21072
rect 17276 21032 18144 21060
rect 17276 21020 17282 21032
rect 18138 21020 18144 21032
rect 18196 21060 18202 21072
rect 18693 21063 18751 21069
rect 18693 21060 18705 21063
rect 18196 21032 18705 21060
rect 18196 21020 18202 21032
rect 18693 21029 18705 21032
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 19058 21020 19064 21072
rect 19116 21020 19122 21072
rect 22066 21060 22094 21100
rect 23106 21088 23112 21100
rect 23164 21088 23170 21140
rect 24210 21088 24216 21140
rect 24268 21128 24274 21140
rect 27157 21131 27215 21137
rect 27157 21128 27169 21131
rect 24268 21100 27169 21128
rect 24268 21088 24274 21100
rect 27157 21097 27169 21100
rect 27203 21097 27215 21131
rect 27157 21091 27215 21097
rect 28074 21088 28080 21140
rect 28132 21128 28138 21140
rect 28629 21131 28687 21137
rect 28629 21128 28641 21131
rect 28132 21100 28641 21128
rect 28132 21088 28138 21100
rect 28629 21097 28641 21100
rect 28675 21097 28687 21131
rect 28629 21091 28687 21097
rect 28810 21088 28816 21140
rect 28868 21128 28874 21140
rect 29270 21128 29276 21140
rect 28868 21100 29276 21128
rect 28868 21088 28874 21100
rect 29270 21088 29276 21100
rect 29328 21088 29334 21140
rect 29362 21088 29368 21140
rect 29420 21088 29426 21140
rect 30558 21088 30564 21140
rect 30616 21128 30622 21140
rect 31021 21131 31079 21137
rect 31021 21128 31033 21131
rect 30616 21100 31033 21128
rect 30616 21088 30622 21100
rect 31021 21097 31033 21100
rect 31067 21097 31079 21131
rect 31021 21091 31079 21097
rect 27433 21063 27491 21069
rect 19996 21032 22094 21060
rect 23676 21032 27016 21060
rect 14829 20995 14887 21001
rect 14829 20961 14841 20995
rect 14875 20961 14887 20995
rect 14829 20955 14887 20961
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 15749 20995 15807 21001
rect 15749 20961 15761 20995
rect 15795 20992 15807 20995
rect 16022 20992 16028 21004
rect 15795 20964 16028 20992
rect 15795 20961 15807 20964
rect 15749 20955 15807 20961
rect 16022 20952 16028 20964
rect 16080 20952 16086 21004
rect 16114 20952 16120 21004
rect 16172 20952 16178 21004
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 19996 21001 20024 21032
rect 19981 20995 20039 21001
rect 19981 20961 19993 20995
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 20622 20952 20628 21004
rect 20680 20952 20686 21004
rect 20809 20995 20867 21001
rect 20809 20961 20821 20995
rect 20855 20992 20867 20995
rect 20990 20992 20996 21004
rect 20855 20964 20996 20992
rect 20855 20961 20867 20964
rect 20809 20955 20867 20961
rect 20990 20952 20996 20964
rect 21048 20952 21054 21004
rect 21266 20952 21272 21004
rect 21324 20952 21330 21004
rect 21542 20952 21548 21004
rect 21600 20952 21606 21004
rect 22922 20952 22928 21004
rect 22980 20952 22986 21004
rect 23474 20952 23480 21004
rect 23532 20952 23538 21004
rect 23676 21001 23704 21032
rect 23661 20995 23719 21001
rect 23661 20961 23673 20995
rect 23707 20961 23719 20995
rect 23661 20955 23719 20961
rect 23937 20995 23995 21001
rect 23937 20961 23949 20995
rect 23983 20961 23995 20995
rect 23937 20955 23995 20961
rect 12492 20896 13860 20924
rect 14553 20927 14611 20933
rect 12492 20884 12498 20896
rect 14553 20893 14565 20927
rect 14599 20924 14611 20927
rect 15470 20924 15476 20936
rect 14599 20896 15476 20924
rect 14599 20893 14611 20896
rect 14553 20887 14611 20893
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 17034 20924 17040 20936
rect 15611 20896 17040 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 17034 20884 17040 20896
rect 17092 20884 17098 20936
rect 18046 20884 18052 20936
rect 18104 20924 18110 20936
rect 19337 20927 19395 20933
rect 19337 20924 19349 20927
rect 18104 20896 19349 20924
rect 18104 20884 18110 20896
rect 19337 20893 19349 20896
rect 19383 20893 19395 20927
rect 19337 20887 19395 20893
rect 19610 20884 19616 20936
rect 19668 20924 19674 20936
rect 20901 20927 20959 20933
rect 20901 20924 20913 20927
rect 19668 20896 20913 20924
rect 19668 20884 19674 20896
rect 20901 20893 20913 20896
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20924 21143 20927
rect 21450 20924 21456 20936
rect 21131 20896 21456 20924
rect 21131 20893 21143 20896
rect 21085 20887 21143 20893
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 15378 20816 15384 20868
rect 15436 20856 15442 20868
rect 16482 20856 16488 20868
rect 15436 20828 16488 20856
rect 15436 20816 15442 20828
rect 16482 20816 16488 20828
rect 16540 20856 16546 20868
rect 17313 20859 17371 20865
rect 17313 20856 17325 20859
rect 16540 20828 17325 20856
rect 16540 20816 16546 20828
rect 17313 20825 17325 20828
rect 17359 20856 17371 20859
rect 19426 20856 19432 20868
rect 17359 20828 19432 20856
rect 17359 20825 17371 20828
rect 17313 20819 17371 20825
rect 19426 20816 19432 20828
rect 19484 20856 19490 20868
rect 19794 20856 19800 20868
rect 19484 20828 19800 20856
rect 19484 20816 19490 20828
rect 19794 20816 19800 20828
rect 19852 20856 19858 20868
rect 21560 20856 21588 20952
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20924 21879 20927
rect 23293 20927 23351 20933
rect 21867 20896 23244 20924
rect 21867 20893 21879 20896
rect 21821 20887 21879 20893
rect 19852 20828 21588 20856
rect 23216 20856 23244 20896
rect 23293 20893 23305 20927
rect 23339 20924 23351 20927
rect 23676 20924 23704 20955
rect 23339 20896 23704 20924
rect 23339 20893 23351 20896
rect 23293 20887 23351 20893
rect 23658 20856 23664 20868
rect 23216 20828 23664 20856
rect 19852 20816 19858 20828
rect 23658 20816 23664 20828
rect 23716 20816 23722 20868
rect 23952 20856 23980 20955
rect 24026 20952 24032 21004
rect 24084 20952 24090 21004
rect 26237 20995 26295 21001
rect 26237 20961 26249 20995
rect 26283 20992 26295 20995
rect 26418 20992 26424 21004
rect 26283 20964 26424 20992
rect 26283 20961 26295 20964
rect 26237 20955 26295 20961
rect 26418 20952 26424 20964
rect 26476 20952 26482 21004
rect 26988 21001 27016 21032
rect 27433 21029 27445 21063
rect 27479 21060 27491 21063
rect 28718 21060 28724 21072
rect 27479 21032 28724 21060
rect 27479 21029 27491 21032
rect 27433 21023 27491 21029
rect 28718 21020 28724 21032
rect 28776 21020 28782 21072
rect 28902 21020 28908 21072
rect 28960 21020 28966 21072
rect 29115 21063 29173 21069
rect 29115 21029 29127 21063
rect 29161 21060 29173 21063
rect 29822 21060 29828 21072
rect 29880 21069 29886 21072
rect 29880 21063 29909 21069
rect 29161 21032 29828 21060
rect 29161 21029 29173 21032
rect 29115 21023 29173 21029
rect 29822 21020 29828 21032
rect 29897 21060 29909 21063
rect 29897 21032 29973 21060
rect 29897 21029 29909 21032
rect 29880 21023 29909 21029
rect 29880 21020 29886 21023
rect 30926 21020 30932 21072
rect 30984 21020 30990 21072
rect 26973 20995 27031 21001
rect 26973 20961 26985 20995
rect 27019 20961 27031 20995
rect 26973 20955 27031 20961
rect 27338 20952 27344 21004
rect 27396 20952 27402 21004
rect 27522 20952 27528 21004
rect 27580 20952 27586 21004
rect 27614 20952 27620 21004
rect 27672 21001 27678 21004
rect 27672 20995 27701 21001
rect 27689 20961 27701 20995
rect 27672 20955 27701 20961
rect 27672 20952 27678 20955
rect 28810 20952 28816 21004
rect 28868 20952 28874 21004
rect 28997 20995 29055 21001
rect 28997 20961 29009 20995
rect 29043 20961 29055 20995
rect 28997 20955 29055 20961
rect 29273 20995 29331 21001
rect 29273 20961 29285 20995
rect 29319 20992 29331 20995
rect 29319 20964 29500 20992
rect 29319 20961 29331 20964
rect 29273 20955 29331 20961
rect 24210 20884 24216 20936
rect 24268 20924 24274 20936
rect 24762 20924 24768 20936
rect 24268 20896 24768 20924
rect 24268 20884 24274 20896
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 27801 20927 27859 20933
rect 27801 20924 27813 20927
rect 25832 20896 27813 20924
rect 25832 20884 25838 20896
rect 27801 20893 27813 20896
rect 27847 20924 27859 20927
rect 27893 20927 27951 20933
rect 27893 20924 27905 20927
rect 27847 20896 27905 20924
rect 27847 20893 27859 20896
rect 27801 20887 27859 20893
rect 27893 20893 27905 20896
rect 27939 20893 27951 20927
rect 27893 20887 27951 20893
rect 28442 20884 28448 20936
rect 28500 20884 28506 20936
rect 29012 20924 29040 20955
rect 29472 20924 29500 20964
rect 29546 20952 29552 21004
rect 29604 20952 29610 21004
rect 29638 20952 29644 21004
rect 29696 20952 29702 21004
rect 29730 20952 29736 21004
rect 29788 20952 29794 21004
rect 30009 20927 30067 20933
rect 29012 20896 29315 20924
rect 29472 20896 29684 20924
rect 25958 20856 25964 20868
rect 23952 20828 25964 20856
rect 25958 20816 25964 20828
rect 26016 20816 26022 20868
rect 29287 20856 29315 20896
rect 29454 20856 29460 20868
rect 29287 20828 29460 20856
rect 29454 20816 29460 20828
rect 29512 20816 29518 20868
rect 29656 20856 29684 20896
rect 30009 20893 30021 20927
rect 30055 20924 30067 20927
rect 30190 20924 30196 20936
rect 30055 20896 30196 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 30190 20884 30196 20896
rect 30248 20884 30254 20936
rect 30745 20927 30803 20933
rect 30745 20893 30757 20927
rect 30791 20924 30803 20927
rect 31202 20924 31208 20936
rect 30791 20896 31208 20924
rect 30791 20893 30803 20896
rect 30745 20887 30803 20893
rect 31202 20884 31208 20896
rect 31260 20884 31266 20936
rect 30101 20859 30159 20865
rect 30101 20856 30113 20859
rect 29656 20828 30113 20856
rect 30101 20825 30113 20828
rect 30147 20825 30159 20859
rect 30101 20819 30159 20825
rect 12894 20788 12900 20800
rect 11256 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20788 12958 20800
rect 13265 20791 13323 20797
rect 13265 20788 13277 20791
rect 12952 20760 13277 20788
rect 12952 20748 12958 20760
rect 13265 20757 13277 20760
rect 13311 20757 13323 20791
rect 13265 20751 13323 20757
rect 15105 20791 15163 20797
rect 15105 20757 15117 20791
rect 15151 20788 15163 20791
rect 15194 20788 15200 20800
rect 15151 20760 15200 20788
rect 15151 20757 15163 20760
rect 15105 20751 15163 20757
rect 15194 20748 15200 20760
rect 15252 20748 15258 20800
rect 15933 20791 15991 20797
rect 15933 20757 15945 20791
rect 15979 20788 15991 20791
rect 16758 20788 16764 20800
rect 15979 20760 16764 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 19702 20748 19708 20800
rect 19760 20788 19766 20800
rect 20073 20791 20131 20797
rect 20073 20788 20085 20791
rect 19760 20760 20085 20788
rect 19760 20748 19766 20760
rect 20073 20757 20085 20760
rect 20119 20757 20131 20791
rect 20073 20751 20131 20757
rect 20162 20748 20168 20800
rect 20220 20788 20226 20800
rect 20714 20788 20720 20800
rect 20220 20760 20720 20788
rect 20220 20748 20226 20760
rect 20714 20748 20720 20760
rect 20772 20788 20778 20800
rect 20993 20791 21051 20797
rect 20993 20788 21005 20791
rect 20772 20760 21005 20788
rect 20772 20748 20778 20760
rect 20993 20757 21005 20760
rect 21039 20757 21051 20791
rect 20993 20751 21051 20757
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24176 20760 24961 20788
rect 24176 20748 24182 20760
rect 24949 20757 24961 20760
rect 24995 20788 25007 20791
rect 26326 20788 26332 20800
rect 24995 20760 26332 20788
rect 24995 20757 25007 20760
rect 24949 20751 25007 20757
rect 26326 20748 26332 20760
rect 26384 20748 26390 20800
rect 26421 20791 26479 20797
rect 26421 20757 26433 20791
rect 26467 20788 26479 20791
rect 26602 20788 26608 20800
rect 26467 20760 26608 20788
rect 26467 20757 26479 20760
rect 26421 20751 26479 20757
rect 26602 20748 26608 20760
rect 26660 20748 26666 20800
rect 27338 20748 27344 20800
rect 27396 20788 27402 20800
rect 29086 20788 29092 20800
rect 27396 20760 29092 20788
rect 27396 20748 27402 20760
rect 29086 20748 29092 20760
rect 29144 20748 29150 20800
rect 552 20698 31648 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 11436 20698
rect 11488 20646 11500 20698
rect 11552 20646 11564 20698
rect 11616 20646 11628 20698
rect 11680 20646 11692 20698
rect 11744 20646 19210 20698
rect 19262 20646 19274 20698
rect 19326 20646 19338 20698
rect 19390 20646 19402 20698
rect 19454 20646 19466 20698
rect 19518 20646 26984 20698
rect 27036 20646 27048 20698
rect 27100 20646 27112 20698
rect 27164 20646 27176 20698
rect 27228 20646 27240 20698
rect 27292 20646 31648 20698
rect 552 20624 31648 20646
rect 13722 20544 13728 20596
rect 13780 20584 13786 20596
rect 13780 20556 13952 20584
rect 13780 20544 13786 20556
rect 7929 20519 7987 20525
rect 7929 20485 7941 20519
rect 7975 20516 7987 20519
rect 8478 20516 8484 20528
rect 7975 20488 8484 20516
rect 7975 20485 7987 20488
rect 7929 20479 7987 20485
rect 8478 20476 8484 20488
rect 8536 20476 8542 20528
rect 9214 20476 9220 20528
rect 9272 20476 9278 20528
rect 13924 20516 13952 20556
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14185 20587 14243 20593
rect 14185 20584 14197 20587
rect 14148 20556 14197 20584
rect 14148 20544 14154 20556
rect 14185 20553 14197 20556
rect 14231 20553 14243 20587
rect 14185 20547 14243 20553
rect 14458 20544 14464 20596
rect 14516 20544 14522 20596
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 16448 20556 17816 20584
rect 16448 20544 16454 20556
rect 13924 20488 14320 20516
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 7708 20420 12434 20448
rect 7708 20408 7714 20420
rect 7944 20389 7972 20420
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20349 7987 20383
rect 7929 20343 7987 20349
rect 8205 20383 8263 20389
rect 8205 20349 8217 20383
rect 8251 20380 8263 20383
rect 8846 20380 8852 20392
rect 8251 20352 8852 20380
rect 8251 20349 8263 20352
rect 8205 20343 8263 20349
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 8938 20340 8944 20392
rect 8996 20340 9002 20392
rect 9030 20340 9036 20392
rect 9088 20340 9094 20392
rect 9950 20380 9956 20392
rect 9140 20352 9956 20380
rect 8113 20315 8171 20321
rect 8113 20281 8125 20315
rect 8159 20312 8171 20315
rect 9140 20312 9168 20352
rect 9950 20340 9956 20352
rect 10008 20340 10014 20392
rect 10336 20389 10364 20420
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 10502 20340 10508 20392
rect 10560 20380 10566 20392
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 10560 20352 10609 20380
rect 10560 20340 10566 20352
rect 10597 20349 10609 20352
rect 10643 20349 10655 20383
rect 10597 20343 10655 20349
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 12406 20380 12434 20420
rect 13446 20408 13452 20460
rect 13504 20448 13510 20460
rect 13909 20451 13967 20457
rect 13504 20420 13860 20448
rect 13504 20408 13510 20420
rect 13722 20380 13728 20392
rect 12406 20352 13728 20380
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 13832 20389 13860 20420
rect 13909 20417 13921 20451
rect 13955 20448 13967 20451
rect 14090 20448 14096 20460
rect 13955 20420 14096 20448
rect 13955 20417 13967 20420
rect 13909 20411 13967 20417
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 14292 20448 14320 20488
rect 15378 20448 15384 20460
rect 14292 20420 15384 20448
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 16393 20451 16451 20457
rect 16393 20417 16405 20451
rect 16439 20448 16451 20451
rect 16482 20448 16488 20460
rect 16439 20420 16488 20448
rect 16439 20417 16451 20420
rect 16393 20411 16451 20417
rect 16482 20408 16488 20420
rect 16540 20408 16546 20460
rect 16758 20408 16764 20460
rect 16816 20408 16822 20460
rect 17788 20448 17816 20556
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18693 20587 18751 20593
rect 18693 20584 18705 20587
rect 18012 20556 18705 20584
rect 18012 20544 18018 20556
rect 18693 20553 18705 20556
rect 18739 20553 18751 20587
rect 18693 20547 18751 20553
rect 18966 20544 18972 20596
rect 19024 20544 19030 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 20070 20584 20076 20596
rect 19475 20556 20076 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 20070 20544 20076 20556
rect 20128 20544 20134 20596
rect 20346 20544 20352 20596
rect 20404 20584 20410 20596
rect 21266 20584 21272 20596
rect 20404 20556 21272 20584
rect 20404 20544 20410 20556
rect 21266 20544 21272 20556
rect 21324 20584 21330 20596
rect 22922 20584 22928 20596
rect 21324 20556 22928 20584
rect 21324 20544 21330 20556
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 23934 20544 23940 20596
rect 23992 20544 23998 20596
rect 25958 20544 25964 20596
rect 26016 20544 26022 20596
rect 26510 20544 26516 20596
rect 26568 20584 26574 20596
rect 28442 20584 28448 20596
rect 26568 20556 28448 20584
rect 26568 20544 26574 20556
rect 18874 20476 18880 20528
rect 18932 20516 18938 20528
rect 20257 20519 20315 20525
rect 20257 20516 20269 20519
rect 18932 20488 20269 20516
rect 18932 20476 18938 20488
rect 20257 20485 20269 20488
rect 20303 20485 20315 20519
rect 20257 20479 20315 20485
rect 26620 20488 28028 20516
rect 19337 20451 19395 20457
rect 17788 20420 19288 20448
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 13998 20340 14004 20392
rect 14056 20340 14062 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 14792 20352 15042 20380
rect 14792 20340 14798 20352
rect 19150 20340 19156 20392
rect 19208 20340 19214 20392
rect 19260 20380 19288 20420
rect 19337 20417 19349 20451
rect 19383 20448 19395 20451
rect 19702 20448 19708 20460
rect 19383 20420 19708 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 21358 20448 21364 20460
rect 19904 20420 21364 20448
rect 19260 20352 19472 20380
rect 8159 20284 9168 20312
rect 9217 20315 9275 20321
rect 8159 20281 8171 20284
rect 8113 20275 8171 20281
rect 9217 20281 9229 20315
rect 9263 20312 9275 20315
rect 10137 20315 10195 20321
rect 10137 20312 10149 20315
rect 9263 20284 10149 20312
rect 9263 20281 9275 20284
rect 9217 20275 9275 20281
rect 10137 20281 10149 20284
rect 10183 20281 10195 20315
rect 10137 20275 10195 20281
rect 11054 20272 11060 20324
rect 11112 20312 11118 20324
rect 11330 20312 11336 20324
rect 11112 20284 11336 20312
rect 11112 20272 11118 20284
rect 11330 20272 11336 20284
rect 11388 20312 11394 20324
rect 11609 20315 11667 20321
rect 11609 20312 11621 20315
rect 11388 20284 11621 20312
rect 11388 20272 11394 20284
rect 11609 20281 11621 20284
rect 11655 20281 11667 20315
rect 11609 20275 11667 20281
rect 13357 20315 13415 20321
rect 13357 20281 13369 20315
rect 13403 20312 13415 20315
rect 13403 20284 14872 20312
rect 13403 20281 13415 20284
rect 13357 20275 13415 20281
rect 9306 20204 9312 20256
rect 9364 20204 9370 20256
rect 10505 20247 10563 20253
rect 10505 20213 10517 20247
rect 10551 20244 10563 20247
rect 10873 20247 10931 20253
rect 10873 20244 10885 20247
rect 10551 20216 10885 20244
rect 10551 20213 10563 20216
rect 10505 20207 10563 20213
rect 10873 20213 10885 20216
rect 10919 20213 10931 20247
rect 10873 20207 10931 20213
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 12802 20244 12808 20256
rect 11940 20216 12808 20244
rect 11940 20204 11946 20216
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 14645 20247 14703 20253
rect 14645 20213 14657 20247
rect 14691 20244 14703 20247
rect 14734 20244 14740 20256
rect 14691 20216 14740 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 14844 20244 14872 20284
rect 16114 20272 16120 20324
rect 16172 20272 16178 20324
rect 17218 20272 17224 20324
rect 17276 20272 17282 20324
rect 18230 20272 18236 20324
rect 18288 20312 18294 20324
rect 18509 20315 18567 20321
rect 18509 20312 18521 20315
rect 18288 20284 18521 20312
rect 18288 20272 18294 20284
rect 18509 20281 18521 20284
rect 18555 20312 18567 20315
rect 18690 20312 18696 20324
rect 18555 20284 18696 20312
rect 18555 20281 18567 20284
rect 18509 20275 18567 20281
rect 18690 20272 18696 20284
rect 18748 20272 18754 20324
rect 18598 20244 18604 20256
rect 14844 20216 18604 20244
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 19444 20244 19472 20352
rect 19518 20340 19524 20392
rect 19576 20380 19582 20392
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 19576 20352 19625 20380
rect 19576 20340 19582 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19904 20380 19932 20420
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21692 20420 22017 20448
rect 21692 20408 21698 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22925 20451 22983 20457
rect 22925 20417 22937 20451
rect 22971 20448 22983 20451
rect 23474 20448 23480 20460
rect 22971 20420 23480 20448
rect 22971 20417 22983 20420
rect 22925 20411 22983 20417
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 24118 20408 24124 20460
rect 24176 20408 24182 20460
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20448 24455 20451
rect 25406 20448 25412 20460
rect 24443 20420 25412 20448
rect 24443 20417 24455 20420
rect 24397 20411 24455 20417
rect 25406 20408 25412 20420
rect 25464 20408 25470 20460
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20448 25927 20451
rect 26620 20448 26648 20488
rect 25915 20420 26648 20448
rect 25915 20417 25927 20420
rect 25869 20411 25927 20417
rect 19613 20343 19671 20349
rect 19720 20352 19932 20380
rect 19720 20321 19748 20352
rect 19978 20340 19984 20392
rect 20036 20340 20042 20392
rect 22649 20383 22707 20389
rect 22649 20380 22661 20383
rect 22066 20352 22661 20380
rect 19705 20315 19763 20321
rect 19705 20281 19717 20315
rect 19751 20281 19763 20315
rect 19705 20275 19763 20281
rect 19797 20315 19855 20321
rect 19797 20281 19809 20315
rect 19843 20312 19855 20315
rect 20070 20312 20076 20324
rect 19843 20284 20076 20312
rect 19843 20281 19855 20284
rect 19797 20275 19855 20281
rect 19720 20244 19748 20275
rect 20070 20272 20076 20284
rect 20128 20272 20134 20324
rect 21266 20272 21272 20324
rect 21324 20272 21330 20324
rect 21726 20272 21732 20324
rect 21784 20272 21790 20324
rect 21818 20272 21824 20324
rect 21876 20312 21882 20324
rect 22066 20312 22094 20352
rect 22649 20349 22661 20352
rect 22695 20349 22707 20383
rect 22649 20343 22707 20349
rect 24026 20340 24032 20392
rect 24084 20340 24090 20392
rect 26234 20340 26240 20392
rect 26292 20340 26298 20392
rect 26329 20383 26387 20389
rect 26329 20349 26341 20383
rect 26375 20349 26387 20383
rect 26329 20343 26387 20349
rect 26421 20383 26479 20389
rect 26421 20349 26433 20383
rect 26467 20380 26479 20383
rect 26510 20380 26516 20392
rect 26467 20352 26516 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 21876 20284 22094 20312
rect 23477 20315 23535 20321
rect 21876 20272 21882 20284
rect 23477 20281 23489 20315
rect 23523 20312 23535 20315
rect 24670 20312 24676 20324
rect 23523 20284 24676 20312
rect 23523 20281 23535 20284
rect 23477 20275 23535 20281
rect 24670 20272 24676 20284
rect 24728 20272 24734 20324
rect 26050 20312 26056 20324
rect 25622 20284 26056 20312
rect 26050 20272 26056 20284
rect 26108 20272 26114 20324
rect 26344 20312 26372 20343
rect 26510 20340 26516 20352
rect 26568 20340 26574 20392
rect 26620 20389 26648 20420
rect 27065 20451 27123 20457
rect 27065 20417 27077 20451
rect 27111 20448 27123 20451
rect 27154 20448 27160 20460
rect 27111 20420 27160 20448
rect 27111 20417 27123 20420
rect 27065 20411 27123 20417
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 28000 20457 28028 20488
rect 27985 20451 28043 20457
rect 27264 20420 27568 20448
rect 26605 20383 26663 20389
rect 26605 20349 26617 20383
rect 26651 20349 26663 20383
rect 26605 20343 26663 20349
rect 26878 20340 26884 20392
rect 26936 20340 26942 20392
rect 26970 20312 26976 20324
rect 26344 20284 26976 20312
rect 26970 20272 26976 20284
rect 27028 20272 27034 20324
rect 27264 20312 27292 20420
rect 27338 20340 27344 20392
rect 27396 20340 27402 20392
rect 27540 20389 27568 20420
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 28368 20448 28396 20556
rect 28442 20544 28448 20556
rect 28500 20544 28506 20596
rect 28718 20544 28724 20596
rect 28776 20544 28782 20596
rect 28810 20544 28816 20596
rect 28868 20584 28874 20596
rect 30282 20584 30288 20596
rect 28868 20556 30288 20584
rect 28868 20544 28874 20556
rect 30282 20544 30288 20556
rect 30340 20584 30346 20596
rect 30745 20587 30803 20593
rect 30745 20584 30757 20587
rect 30340 20556 30757 20584
rect 30340 20544 30346 20556
rect 30745 20553 30757 20556
rect 30791 20553 30803 20587
rect 30745 20547 30803 20553
rect 28537 20519 28595 20525
rect 28537 20485 28549 20519
rect 28583 20516 28595 20519
rect 28583 20488 29132 20516
rect 28583 20485 28595 20488
rect 28537 20479 28595 20485
rect 28902 20448 28908 20460
rect 28368 20420 28908 20448
rect 27985 20411 28043 20417
rect 27525 20383 27583 20389
rect 27525 20349 27537 20383
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 27614 20340 27620 20392
rect 27672 20389 27678 20392
rect 27672 20383 27701 20389
rect 27689 20349 27701 20383
rect 27672 20343 27701 20349
rect 27801 20383 27859 20389
rect 27801 20349 27813 20383
rect 27847 20380 27859 20383
rect 28258 20380 28264 20392
rect 27847 20352 28264 20380
rect 27847 20349 27859 20352
rect 27801 20343 27859 20349
rect 27672 20340 27678 20343
rect 28258 20340 28264 20352
rect 28316 20380 28322 20392
rect 28442 20380 28448 20392
rect 28316 20352 28448 20380
rect 28316 20340 28322 20352
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 28644 20389 28672 20420
rect 28902 20408 28908 20420
rect 28960 20408 28966 20460
rect 28994 20408 29000 20460
rect 29052 20408 29058 20460
rect 29104 20448 29132 20488
rect 30374 20476 30380 20528
rect 30432 20516 30438 20528
rect 30929 20519 30987 20525
rect 30929 20516 30941 20519
rect 30432 20488 30941 20516
rect 30432 20476 30438 20488
rect 30929 20485 30941 20488
rect 30975 20485 30987 20519
rect 30929 20479 30987 20485
rect 29104 20420 31156 20448
rect 28629 20383 28687 20389
rect 28629 20349 28641 20383
rect 28675 20349 28687 20383
rect 28629 20343 28687 20349
rect 28718 20340 28724 20392
rect 28776 20380 28782 20392
rect 28813 20383 28871 20389
rect 28813 20380 28825 20383
rect 28776 20352 28825 20380
rect 28776 20340 28782 20352
rect 28813 20349 28825 20352
rect 28859 20349 28871 20383
rect 30558 20380 30564 20392
rect 30406 20352 30564 20380
rect 28813 20343 28871 20349
rect 30558 20340 30564 20352
rect 30616 20340 30622 20392
rect 30834 20340 30840 20392
rect 30892 20340 30898 20392
rect 31128 20389 31156 20420
rect 31113 20383 31171 20389
rect 31113 20349 31125 20383
rect 31159 20349 31171 20383
rect 31113 20343 31171 20349
rect 27080 20284 27292 20312
rect 27434 20315 27492 20321
rect 19444 20216 19748 20244
rect 19978 20204 19984 20256
rect 20036 20244 20042 20256
rect 22097 20247 22155 20253
rect 22097 20244 22109 20247
rect 20036 20216 22109 20244
rect 20036 20204 20042 20216
rect 22097 20213 22109 20216
rect 22143 20213 22155 20247
rect 22097 20207 22155 20213
rect 22738 20204 22744 20256
rect 22796 20244 22802 20256
rect 26697 20247 26755 20253
rect 26697 20244 26709 20247
rect 22796 20216 26709 20244
rect 22796 20204 22802 20216
rect 26697 20213 26709 20216
rect 26743 20213 26755 20247
rect 26697 20207 26755 20213
rect 26786 20204 26792 20256
rect 26844 20244 26850 20256
rect 27080 20244 27108 20284
rect 27434 20281 27446 20315
rect 27480 20281 27492 20315
rect 27434 20275 27492 20281
rect 26844 20216 27108 20244
rect 27157 20247 27215 20253
rect 26844 20204 26850 20216
rect 27157 20213 27169 20247
rect 27203 20244 27215 20247
rect 27338 20244 27344 20256
rect 27203 20216 27344 20244
rect 27203 20213 27215 20216
rect 27157 20207 27215 20213
rect 27338 20204 27344 20216
rect 27396 20204 27402 20256
rect 27448 20244 27476 20275
rect 29270 20272 29276 20324
rect 29328 20272 29334 20324
rect 31297 20315 31355 20321
rect 31297 20312 31309 20315
rect 30576 20284 31309 20312
rect 27522 20244 27528 20256
rect 27448 20216 27528 20244
rect 27522 20204 27528 20216
rect 27580 20204 27586 20256
rect 28994 20204 29000 20256
rect 29052 20244 29058 20256
rect 30576 20244 30604 20284
rect 31297 20281 31309 20284
rect 31343 20281 31355 20315
rect 31297 20275 31355 20281
rect 29052 20216 30604 20244
rect 29052 20204 29058 20216
rect 552 20154 31648 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 12096 20154
rect 12148 20102 12160 20154
rect 12212 20102 12224 20154
rect 12276 20102 12288 20154
rect 12340 20102 12352 20154
rect 12404 20102 19870 20154
rect 19922 20102 19934 20154
rect 19986 20102 19998 20154
rect 20050 20102 20062 20154
rect 20114 20102 20126 20154
rect 20178 20102 27644 20154
rect 27696 20102 27708 20154
rect 27760 20102 27772 20154
rect 27824 20102 27836 20154
rect 27888 20102 27900 20154
rect 27952 20102 31648 20154
rect 552 20080 31648 20102
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 11054 20040 11060 20052
rect 7248 20012 11060 20040
rect 7248 20000 7254 20012
rect 7190 19864 7196 19916
rect 7248 19864 7254 19916
rect 9048 19913 9076 20012
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 11501 20043 11559 20049
rect 11501 20009 11513 20043
rect 11547 20040 11559 20043
rect 12161 20043 12219 20049
rect 11547 20012 11836 20040
rect 11547 20009 11559 20012
rect 11501 20003 11559 20009
rect 9214 19932 9220 19984
rect 9272 19972 9278 19984
rect 9309 19975 9367 19981
rect 9309 19972 9321 19975
rect 9272 19944 9321 19972
rect 9272 19932 9278 19944
rect 9309 19941 9321 19944
rect 9355 19941 9367 19975
rect 9309 19935 9367 19941
rect 9582 19932 9588 19984
rect 9640 19972 9646 19984
rect 10962 19972 10968 19984
rect 9640 19944 9798 19972
rect 10796 19944 10968 19972
rect 9640 19932 9646 19944
rect 9033 19907 9091 19913
rect 7466 19796 7472 19848
rect 7524 19796 7530 19848
rect 8588 19768 8616 19890
rect 9033 19873 9045 19907
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 8938 19796 8944 19848
rect 8996 19836 9002 19848
rect 10796 19845 10824 19944
rect 10962 19932 10968 19944
rect 11020 19972 11026 19984
rect 11516 19972 11544 20003
rect 11020 19944 11544 19972
rect 11701 19975 11759 19981
rect 11020 19932 11026 19944
rect 11701 19941 11713 19975
rect 11747 19941 11759 19975
rect 11808 19972 11836 20012
rect 12161 20009 12173 20043
rect 12207 20040 12219 20043
rect 12342 20040 12348 20052
rect 12207 20012 12348 20040
rect 12207 20009 12219 20012
rect 12161 20003 12219 20009
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 12434 20000 12440 20052
rect 12492 20000 12498 20052
rect 12526 20000 12532 20052
rect 12584 20040 12590 20052
rect 12989 20043 13047 20049
rect 12584 20012 12940 20040
rect 12584 20000 12590 20012
rect 12250 19972 12256 19984
rect 11808 19944 12256 19972
rect 11701 19935 11759 19941
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11716 19904 11744 19935
rect 12250 19932 12256 19944
rect 12308 19932 12314 19984
rect 12912 19972 12940 20012
rect 12989 20009 13001 20043
rect 13035 20040 13047 20043
rect 13998 20040 14004 20052
rect 13035 20012 14004 20040
rect 13035 20009 13047 20012
rect 12989 20003 13047 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 15580 20012 16436 20040
rect 15580 19984 15608 20012
rect 12912 19944 13952 19972
rect 12609 19916 12667 19919
rect 11112 19876 11744 19904
rect 11112 19864 11118 19876
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 12066 19864 12072 19916
rect 12124 19864 12130 19916
rect 12609 19913 12624 19916
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19873 12495 19907
rect 12609 19879 12621 19913
rect 12609 19873 12624 19879
rect 12437 19867 12495 19873
rect 10781 19839 10839 19845
rect 8996 19808 10732 19836
rect 8996 19796 9002 19808
rect 10704 19768 10732 19808
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11296 19808 11468 19836
rect 11296 19796 11302 19808
rect 11330 19768 11336 19780
rect 8588 19740 9076 19768
rect 10704 19740 11336 19768
rect 8938 19660 8944 19712
rect 8996 19660 9002 19712
rect 9048 19700 9076 19740
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 11440 19768 11468 19808
rect 12299 19771 12357 19777
rect 12299 19768 12311 19771
rect 11440 19740 12311 19768
rect 12299 19737 12311 19740
rect 12345 19737 12357 19771
rect 12452 19768 12480 19867
rect 12618 19864 12624 19873
rect 12676 19864 12682 19916
rect 12802 19864 12808 19916
rect 12860 19864 12866 19916
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13538 19904 13544 19916
rect 13495 19876 13544 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 13817 19907 13875 19913
rect 13817 19873 13829 19907
rect 13863 19873 13875 19907
rect 13817 19867 13875 19873
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 13228 19808 13737 19836
rect 13228 19796 13234 19808
rect 13725 19805 13737 19808
rect 13771 19836 13783 19839
rect 13832 19836 13860 19867
rect 13924 19845 13952 19944
rect 15562 19932 15568 19984
rect 15620 19932 15626 19984
rect 15781 19975 15839 19981
rect 15781 19941 15793 19975
rect 15827 19972 15839 19975
rect 16298 19972 16304 19984
rect 15827 19944 16304 19972
rect 15827 19941 15839 19944
rect 15781 19935 15839 19941
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 16408 19972 16436 20012
rect 17034 20000 17040 20052
rect 17092 20000 17098 20052
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17405 20043 17463 20049
rect 17405 20040 17417 20043
rect 17184 20012 17417 20040
rect 17184 20000 17190 20012
rect 17405 20009 17417 20012
rect 17451 20040 17463 20043
rect 18617 20043 18675 20049
rect 18617 20040 18629 20043
rect 17451 20012 18629 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 18617 20009 18629 20012
rect 18663 20009 18675 20043
rect 18617 20003 18675 20009
rect 19245 20043 19303 20049
rect 19245 20009 19257 20043
rect 19291 20040 19303 20043
rect 19426 20040 19432 20052
rect 19291 20012 19432 20040
rect 19291 20009 19303 20012
rect 19245 20003 19303 20009
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 20254 20040 20260 20052
rect 19628 20012 20260 20040
rect 18230 19972 18236 19984
rect 16408 19944 18236 19972
rect 14277 19907 14335 19913
rect 14277 19873 14289 19907
rect 14323 19904 14335 19907
rect 14734 19904 14740 19916
rect 14323 19876 14740 19904
rect 14323 19873 14335 19876
rect 14277 19867 14335 19873
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 15010 19864 15016 19916
rect 15068 19864 15074 19916
rect 17236 19913 17264 19944
rect 18230 19932 18236 19944
rect 18288 19932 18294 19984
rect 18414 19932 18420 19984
rect 18472 19932 18478 19984
rect 18874 19932 18880 19984
rect 18932 19932 18938 19984
rect 18966 19932 18972 19984
rect 19024 19972 19030 19984
rect 19077 19975 19135 19981
rect 19077 19972 19089 19975
rect 19024 19944 19089 19972
rect 19024 19932 19030 19944
rect 19077 19941 19089 19944
rect 19123 19941 19135 19975
rect 19518 19972 19524 19984
rect 19077 19935 19135 19941
rect 19352 19944 19524 19972
rect 16485 19907 16543 19913
rect 16485 19904 16497 19907
rect 15120 19876 16497 19904
rect 13771 19808 13860 19836
rect 13909 19839 13967 19845
rect 13771 19805 13783 19808
rect 13725 19799 13783 19805
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 13955 19808 14381 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 14369 19805 14381 19808
rect 14415 19836 14427 19839
rect 15120 19836 15148 19876
rect 16485 19873 16497 19876
rect 16531 19873 16543 19907
rect 16485 19867 16543 19873
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 17552 19876 17816 19904
rect 17552 19864 17558 19876
rect 14415 19808 15148 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 16114 19796 16120 19848
rect 16172 19796 16178 19848
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 13265 19771 13323 19777
rect 13265 19768 13277 19771
rect 12452 19740 13277 19768
rect 12299 19731 12357 19737
rect 13265 19737 13277 19740
rect 13311 19737 13323 19771
rect 13265 19731 13323 19737
rect 13446 19728 13452 19780
rect 13504 19768 13510 19780
rect 14185 19771 14243 19777
rect 14185 19768 14197 19771
rect 13504 19740 14197 19768
rect 13504 19728 13510 19740
rect 14185 19737 14197 19740
rect 14231 19737 14243 19771
rect 14185 19731 14243 19737
rect 15933 19771 15991 19777
rect 15933 19737 15945 19771
rect 15979 19768 15991 19771
rect 16316 19768 16344 19799
rect 16390 19796 16396 19848
rect 16448 19796 16454 19848
rect 16574 19796 16580 19848
rect 16632 19796 16638 19848
rect 16666 19796 16672 19848
rect 16724 19836 16730 19848
rect 17589 19839 17647 19845
rect 17589 19836 17601 19839
rect 16724 19808 17601 19836
rect 16724 19796 16730 19808
rect 17589 19805 17601 19808
rect 17635 19805 17647 19839
rect 17788 19836 17816 19876
rect 17862 19864 17868 19916
rect 17920 19864 17926 19916
rect 18046 19864 18052 19916
rect 18104 19864 18110 19916
rect 19352 19913 19380 19944
rect 19518 19932 19524 19944
rect 19576 19932 19582 19984
rect 19628 19981 19656 20012
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 21427 20043 21485 20049
rect 21427 20040 21439 20043
rect 21232 20012 21439 20040
rect 21232 20000 21238 20012
rect 21427 20009 21439 20012
rect 21473 20009 21485 20043
rect 21427 20003 21485 20009
rect 21729 20043 21787 20049
rect 21729 20009 21741 20043
rect 21775 20040 21787 20043
rect 23474 20040 23480 20052
rect 21775 20012 23480 20040
rect 21775 20009 21787 20012
rect 21729 20003 21787 20009
rect 23474 20000 23480 20012
rect 23532 20000 23538 20052
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 26878 20040 26884 20052
rect 23992 20012 26884 20040
rect 23992 20000 23998 20012
rect 26878 20000 26884 20012
rect 26936 20000 26942 20052
rect 26970 20000 26976 20052
rect 27028 20040 27034 20052
rect 28353 20043 28411 20049
rect 28353 20040 28365 20043
rect 27028 20012 28365 20040
rect 27028 20000 27034 20012
rect 28353 20009 28365 20012
rect 28399 20009 28411 20043
rect 28353 20003 28411 20009
rect 28534 20000 28540 20052
rect 28592 20040 28598 20052
rect 28810 20040 28816 20052
rect 28592 20012 28816 20040
rect 28592 20000 28598 20012
rect 28810 20000 28816 20012
rect 28868 20000 28874 20052
rect 28902 20000 28908 20052
rect 28960 20040 28966 20052
rect 28960 20012 29106 20040
rect 28960 20000 28966 20012
rect 19613 19975 19671 19981
rect 19613 19941 19625 19975
rect 19659 19941 19671 19975
rect 21266 19972 21272 19984
rect 20838 19944 21272 19972
rect 19613 19935 19671 19941
rect 21266 19932 21272 19944
rect 21324 19932 21330 19984
rect 21634 19932 21640 19984
rect 21692 19932 21698 19984
rect 22922 19972 22928 19984
rect 22770 19944 22928 19972
rect 22922 19932 22928 19944
rect 22980 19972 22986 19984
rect 23290 19972 23296 19984
rect 22980 19944 23296 19972
rect 22980 19932 22986 19944
rect 23290 19932 23296 19944
rect 23348 19932 23354 19984
rect 23750 19972 23756 19984
rect 23584 19944 23756 19972
rect 23584 19913 23612 19944
rect 23750 19932 23756 19944
rect 23808 19972 23814 19984
rect 24118 19972 24124 19984
rect 23808 19944 24124 19972
rect 23808 19932 23814 19944
rect 24118 19932 24124 19944
rect 24176 19932 24182 19984
rect 24854 19932 24860 19984
rect 24912 19932 24918 19984
rect 29078 19981 29106 20012
rect 29270 20000 29276 20052
rect 29328 20040 29334 20052
rect 29641 20043 29699 20049
rect 29641 20040 29653 20043
rect 29328 20012 29653 20040
rect 29328 20000 29334 20012
rect 29641 20009 29653 20012
rect 29687 20009 29699 20043
rect 29641 20003 29699 20009
rect 29822 20000 29828 20052
rect 29880 20040 29886 20052
rect 31754 20040 31760 20052
rect 29880 20012 31760 20040
rect 29880 20000 29886 20012
rect 29063 19975 29121 19981
rect 29063 19941 29075 19975
rect 29109 19941 29121 19975
rect 29063 19935 29121 19941
rect 29181 19975 29239 19981
rect 29181 19941 29193 19975
rect 29227 19972 29239 19975
rect 29454 19972 29460 19984
rect 29227 19944 29460 19972
rect 29227 19941 29239 19944
rect 29181 19935 29239 19941
rect 29454 19932 29460 19944
rect 29512 19972 29518 19984
rect 30162 19981 30190 20012
rect 31754 20000 31760 20012
rect 31812 20000 31818 20052
rect 30009 19975 30067 19981
rect 30009 19972 30021 19975
rect 29512 19944 30021 19972
rect 29512 19932 29518 19944
rect 30009 19941 30021 19944
rect 30055 19941 30067 19975
rect 30009 19935 30067 19941
rect 30147 19975 30205 19981
rect 30147 19941 30159 19975
rect 30193 19941 30205 19975
rect 30147 19935 30205 19941
rect 30282 19932 30288 19984
rect 30340 19972 30346 19984
rect 30340 19944 30972 19972
rect 30340 19932 30346 19944
rect 18141 19907 18199 19913
rect 18141 19873 18153 19907
rect 18187 19904 18199 19907
rect 19337 19907 19395 19913
rect 18187 19876 19288 19904
rect 18187 19873 18199 19876
rect 18141 19867 18199 19873
rect 19260 19836 19288 19876
rect 19337 19873 19349 19907
rect 19383 19873 19395 19907
rect 19337 19867 19395 19873
rect 23477 19907 23535 19913
rect 23477 19873 23489 19907
rect 23523 19904 23535 19907
rect 23569 19907 23627 19913
rect 23569 19904 23581 19907
rect 23523 19876 23581 19904
rect 23523 19873 23535 19876
rect 23477 19867 23535 19873
rect 23569 19873 23581 19876
rect 23615 19873 23627 19907
rect 23569 19867 23627 19873
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 26421 19907 26479 19913
rect 26421 19904 26433 19907
rect 26384 19876 26433 19904
rect 26384 19864 26390 19876
rect 26421 19873 26433 19876
rect 26467 19873 26479 19907
rect 27982 19904 27988 19916
rect 27830 19876 27988 19904
rect 26421 19867 26479 19873
rect 27982 19864 27988 19876
rect 28040 19864 28046 19916
rect 28534 19864 28540 19916
rect 28592 19864 28598 19916
rect 28813 19907 28871 19913
rect 28813 19873 28825 19907
rect 28859 19904 28871 19907
rect 29272 19907 29330 19913
rect 28859 19876 29106 19904
rect 28859 19873 28871 19876
rect 28813 19867 28871 19873
rect 23201 19839 23259 19845
rect 17788 19808 19196 19836
rect 19260 19808 19334 19836
rect 17589 19799 17647 19805
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 15979 19740 17785 19768
rect 15979 19737 15991 19740
rect 15933 19731 15991 19737
rect 17773 19737 17785 19740
rect 17819 19737 17831 19771
rect 17773 19731 17831 19737
rect 18322 19728 18328 19780
rect 18380 19728 18386 19780
rect 9490 19700 9496 19712
rect 9048 19672 9496 19700
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12805 19703 12863 19709
rect 12805 19700 12817 19703
rect 11563 19672 12817 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12805 19669 12817 19672
rect 12851 19700 12863 19703
rect 12894 19700 12900 19712
rect 12851 19672 12900 19700
rect 12851 19669 12863 19672
rect 12805 19663 12863 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13354 19660 13360 19712
rect 13412 19700 13418 19712
rect 13633 19703 13691 19709
rect 13633 19700 13645 19703
rect 13412 19672 13645 19700
rect 13412 19660 13418 19672
rect 13633 19669 13645 19672
rect 13679 19669 13691 19703
rect 13633 19663 13691 19669
rect 13906 19660 13912 19712
rect 13964 19660 13970 19712
rect 15746 19660 15752 19712
rect 15804 19660 15810 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16390 19700 16396 19712
rect 16080 19672 16396 19700
rect 16080 19660 16086 19672
rect 16390 19660 16396 19672
rect 16448 19700 16454 19712
rect 17681 19703 17739 19709
rect 17681 19700 17693 19703
rect 16448 19672 17693 19700
rect 16448 19660 16454 19672
rect 17681 19669 17693 19672
rect 17727 19669 17739 19703
rect 17681 19663 17739 19669
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 18690 19700 18696 19712
rect 18647 19672 18696 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 18785 19703 18843 19709
rect 18785 19669 18797 19703
rect 18831 19700 18843 19703
rect 19058 19700 19064 19712
rect 18831 19672 19064 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 19058 19660 19064 19672
rect 19116 19660 19122 19712
rect 19168 19700 19196 19808
rect 19306 19780 19334 19808
rect 23201 19805 23213 19839
rect 23247 19836 23259 19839
rect 23247 19808 23612 19836
rect 23247 19805 23259 19808
rect 23201 19799 23259 19805
rect 23584 19780 23612 19808
rect 23842 19796 23848 19848
rect 23900 19796 23906 19848
rect 24394 19796 24400 19848
rect 24452 19836 24458 19848
rect 25409 19839 25467 19845
rect 25409 19836 25421 19839
rect 24452 19808 25421 19836
rect 24452 19796 24458 19808
rect 25409 19805 25421 19808
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19805 26019 19839
rect 25961 19799 26019 19805
rect 19306 19740 19340 19780
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 20806 19728 20812 19780
rect 20864 19768 20870 19780
rect 21269 19771 21327 19777
rect 21269 19768 21281 19771
rect 20864 19740 21281 19768
rect 20864 19728 20870 19740
rect 21269 19737 21281 19740
rect 21315 19737 21327 19771
rect 21818 19768 21824 19780
rect 21269 19731 21327 19737
rect 21376 19740 21824 19768
rect 20824 19700 20852 19728
rect 19168 19672 20852 19700
rect 20990 19660 20996 19712
rect 21048 19700 21054 19712
rect 21085 19703 21143 19709
rect 21085 19700 21097 19703
rect 21048 19672 21097 19700
rect 21048 19660 21054 19672
rect 21085 19669 21097 19672
rect 21131 19700 21143 19703
rect 21376 19700 21404 19740
rect 21818 19728 21824 19740
rect 21876 19728 21882 19780
rect 23566 19728 23572 19780
rect 23624 19728 23630 19780
rect 25038 19728 25044 19780
rect 25096 19768 25102 19780
rect 25317 19771 25375 19777
rect 25317 19768 25329 19771
rect 25096 19740 25329 19768
rect 25096 19728 25102 19740
rect 25317 19737 25329 19740
rect 25363 19768 25375 19771
rect 25976 19768 26004 19799
rect 26694 19796 26700 19848
rect 26752 19796 26758 19848
rect 26786 19796 26792 19848
rect 26844 19836 26850 19848
rect 28166 19836 28172 19848
rect 26844 19808 28172 19836
rect 26844 19796 26850 19808
rect 28166 19796 28172 19808
rect 28224 19796 28230 19848
rect 28350 19796 28356 19848
rect 28408 19836 28414 19848
rect 28629 19839 28687 19845
rect 28629 19836 28641 19839
rect 28408 19808 28641 19836
rect 28408 19796 28414 19808
rect 28629 19805 28641 19808
rect 28675 19805 28687 19839
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28629 19799 28687 19805
rect 28828 19808 28917 19836
rect 28442 19768 28448 19780
rect 25363 19740 26004 19768
rect 27724 19740 28448 19768
rect 25363 19737 25375 19740
rect 25317 19731 25375 19737
rect 21131 19672 21404 19700
rect 21453 19703 21511 19709
rect 21131 19669 21143 19672
rect 21085 19663 21143 19669
rect 21453 19669 21465 19703
rect 21499 19700 21511 19703
rect 21542 19700 21548 19712
rect 21499 19672 21548 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 21542 19660 21548 19672
rect 21600 19700 21606 19712
rect 22094 19700 22100 19712
rect 21600 19672 22100 19700
rect 21600 19660 21606 19672
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 24210 19660 24216 19712
rect 24268 19700 24274 19712
rect 25682 19700 25688 19712
rect 24268 19672 25688 19700
rect 24268 19660 24274 19672
rect 25682 19660 25688 19672
rect 25740 19660 25746 19712
rect 26234 19660 26240 19712
rect 26292 19700 26298 19712
rect 27724 19700 27752 19740
rect 28442 19728 28448 19740
rect 28500 19728 28506 19780
rect 28534 19728 28540 19780
rect 28592 19768 28598 19780
rect 28644 19768 28672 19799
rect 28592 19740 28672 19768
rect 28592 19728 28598 19740
rect 28828 19712 28856 19808
rect 28905 19805 28917 19808
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 29078 19768 29106 19876
rect 29272 19873 29284 19907
rect 29318 19873 29330 19907
rect 29272 19867 29330 19873
rect 29288 19836 29316 19867
rect 29362 19864 29368 19916
rect 29420 19864 29426 19916
rect 29825 19907 29883 19913
rect 29825 19873 29837 19907
rect 29871 19873 29883 19907
rect 29825 19867 29883 19873
rect 29638 19836 29644 19848
rect 29288 19808 29644 19836
rect 29638 19796 29644 19808
rect 29696 19796 29702 19848
rect 29454 19768 29460 19780
rect 29078 19740 29460 19768
rect 29454 19728 29460 19740
rect 29512 19728 29518 19780
rect 29840 19768 29868 19867
rect 29914 19864 29920 19916
rect 29972 19864 29978 19916
rect 30944 19913 30972 19944
rect 30929 19907 30987 19913
rect 30929 19873 30941 19907
rect 30975 19873 30987 19907
rect 30929 19867 30987 19873
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19873 31171 19907
rect 31113 19867 31171 19873
rect 30285 19839 30343 19845
rect 30285 19805 30297 19839
rect 30331 19836 30343 19839
rect 30377 19839 30435 19845
rect 30377 19836 30389 19839
rect 30331 19808 30389 19836
rect 30331 19805 30343 19808
rect 30285 19799 30343 19805
rect 30377 19805 30389 19808
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 30466 19796 30472 19848
rect 30524 19836 30530 19848
rect 31128 19836 31156 19867
rect 31294 19864 31300 19916
rect 31352 19864 31358 19916
rect 30524 19808 31156 19836
rect 30524 19796 30530 19808
rect 30650 19768 30656 19780
rect 29840 19740 30656 19768
rect 30650 19728 30656 19740
rect 30708 19728 30714 19780
rect 26292 19672 27752 19700
rect 26292 19660 26298 19672
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 28169 19703 28227 19709
rect 28169 19700 28181 19703
rect 27856 19672 28181 19700
rect 27856 19660 27862 19672
rect 28169 19669 28181 19672
rect 28215 19700 28227 19703
rect 28258 19700 28264 19712
rect 28215 19672 28264 19700
rect 28215 19669 28227 19672
rect 28169 19663 28227 19669
rect 28258 19660 28264 19672
rect 28316 19660 28322 19712
rect 28626 19660 28632 19712
rect 28684 19700 28690 19712
rect 28810 19700 28816 19712
rect 28684 19672 28816 19700
rect 28684 19660 28690 19672
rect 28810 19660 28816 19672
rect 28868 19660 28874 19712
rect 29270 19660 29276 19712
rect 29328 19700 29334 19712
rect 29549 19703 29607 19709
rect 29549 19700 29561 19703
rect 29328 19672 29561 19700
rect 29328 19660 29334 19672
rect 29549 19669 29561 19672
rect 29595 19669 29607 19703
rect 29549 19663 29607 19669
rect 29730 19660 29736 19712
rect 29788 19700 29794 19712
rect 31113 19703 31171 19709
rect 31113 19700 31125 19703
rect 29788 19672 31125 19700
rect 29788 19660 29794 19672
rect 31113 19669 31125 19672
rect 31159 19669 31171 19703
rect 31113 19663 31171 19669
rect 552 19610 31648 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 11436 19610
rect 11488 19558 11500 19610
rect 11552 19558 11564 19610
rect 11616 19558 11628 19610
rect 11680 19558 11692 19610
rect 11744 19558 19210 19610
rect 19262 19558 19274 19610
rect 19326 19558 19338 19610
rect 19390 19558 19402 19610
rect 19454 19558 19466 19610
rect 19518 19558 26984 19610
rect 27036 19558 27048 19610
rect 27100 19558 27112 19610
rect 27164 19558 27176 19610
rect 27228 19558 27240 19610
rect 27292 19558 31648 19610
rect 552 19536 31648 19558
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 7524 19468 8401 19496
rect 7524 19456 7530 19468
rect 8389 19465 8401 19468
rect 8435 19465 8447 19499
rect 8389 19459 8447 19465
rect 8757 19499 8815 19505
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 8938 19496 8944 19508
rect 8803 19468 8944 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 8938 19456 8944 19468
rect 8996 19496 9002 19508
rect 10594 19496 10600 19508
rect 8996 19468 10600 19496
rect 8996 19456 9002 19468
rect 10594 19456 10600 19468
rect 10652 19496 10658 19508
rect 11054 19496 11060 19508
rect 10652 19468 11060 19496
rect 10652 19456 10658 19468
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11977 19499 12035 19505
rect 11977 19465 11989 19499
rect 12023 19496 12035 19499
rect 12066 19496 12072 19508
rect 12023 19468 12072 19496
rect 12023 19465 12035 19468
rect 11977 19459 12035 19465
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 13078 19456 13084 19508
rect 13136 19456 13142 19508
rect 14090 19496 14096 19508
rect 13464 19468 14096 19496
rect 11072 19428 11100 19456
rect 12802 19428 12808 19440
rect 11072 19400 12808 19428
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19360 8907 19363
rect 9306 19360 9312 19372
rect 8895 19332 9312 19360
rect 8895 19329 8907 19332
rect 8849 19323 8907 19329
rect 9306 19320 9312 19332
rect 9364 19320 9370 19372
rect 11330 19320 11336 19372
rect 11388 19360 11394 19372
rect 11388 19332 12756 19360
rect 11388 19320 11394 19332
rect 5442 19252 5448 19304
rect 5500 19292 5506 19304
rect 6457 19295 6515 19301
rect 6457 19292 6469 19295
rect 5500 19264 6469 19292
rect 5500 19252 5506 19264
rect 6457 19261 6469 19264
rect 6503 19261 6515 19295
rect 6457 19255 6515 19261
rect 8478 19252 8484 19304
rect 8536 19292 8542 19304
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8536 19264 8585 19292
rect 8536 19252 8542 19264
rect 8573 19261 8585 19264
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 12161 19295 12219 19301
rect 12161 19261 12173 19295
rect 12207 19261 12219 19295
rect 12161 19255 12219 19261
rect 3878 19184 3884 19236
rect 3936 19224 3942 19236
rect 9030 19224 9036 19236
rect 3936 19196 9036 19224
rect 3936 19184 3942 19196
rect 9030 19184 9036 19196
rect 9088 19184 9094 19236
rect 10042 19224 10048 19236
rect 9232 19196 10048 19224
rect 9232 19168 9260 19196
rect 10042 19184 10048 19196
rect 10100 19224 10106 19236
rect 12066 19224 12072 19236
rect 10100 19196 12072 19224
rect 10100 19184 10106 19196
rect 12066 19184 12072 19196
rect 12124 19184 12130 19236
rect 12176 19224 12204 19255
rect 12434 19252 12440 19304
rect 12492 19252 12498 19304
rect 12728 19292 12756 19332
rect 13262 19320 13268 19372
rect 13320 19320 13326 19372
rect 13081 19295 13139 19301
rect 13081 19294 13093 19295
rect 13004 19292 13093 19294
rect 12728 19266 13093 19292
rect 12728 19264 13032 19266
rect 13081 19261 13093 19266
rect 13127 19261 13139 19295
rect 13280 19292 13308 19320
rect 13081 19255 13139 19261
rect 13188 19264 13308 19292
rect 13357 19295 13415 19301
rect 12986 19224 12992 19236
rect 12176 19196 12992 19224
rect 12986 19184 12992 19196
rect 13044 19184 13050 19236
rect 3418 19116 3424 19168
rect 3476 19156 3482 19168
rect 6270 19156 6276 19168
rect 3476 19128 6276 19156
rect 3476 19116 3482 19128
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 6362 19116 6368 19168
rect 6420 19116 6426 19168
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 9214 19156 9220 19168
rect 6880 19128 9220 19156
rect 6880 19116 6886 19128
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 12345 19159 12403 19165
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 13188 19156 13216 19264
rect 13357 19261 13369 19295
rect 13403 19292 13415 19295
rect 13464 19292 13492 19468
rect 14090 19456 14096 19468
rect 14148 19496 14154 19508
rect 14185 19499 14243 19505
rect 14185 19496 14197 19499
rect 14148 19468 14197 19496
rect 14148 19456 14154 19468
rect 14185 19465 14197 19468
rect 14231 19465 14243 19499
rect 14185 19459 14243 19465
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 16632 19468 16681 19496
rect 16632 19456 16638 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 17126 19456 17132 19508
rect 17184 19456 17190 19508
rect 17494 19456 17500 19508
rect 17552 19456 17558 19508
rect 18598 19456 18604 19508
rect 18656 19496 18662 19508
rect 19153 19499 19211 19505
rect 19153 19496 19165 19499
rect 18656 19468 19165 19496
rect 18656 19456 18662 19468
rect 19153 19465 19165 19468
rect 19199 19496 19211 19499
rect 20438 19496 20444 19508
rect 19199 19468 20444 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 21726 19496 21732 19508
rect 21223 19468 21732 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 23842 19456 23848 19508
rect 23900 19456 23906 19508
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24084 19468 25360 19496
rect 24084 19456 24090 19468
rect 13630 19388 13636 19440
rect 13688 19428 13694 19440
rect 13688 19400 14780 19428
rect 13688 19388 13694 19400
rect 14752 19372 14780 19400
rect 18322 19388 18328 19440
rect 18380 19428 18386 19440
rect 20346 19428 20352 19440
rect 18380 19400 20352 19428
rect 18380 19388 18386 19400
rect 20346 19388 20352 19400
rect 20404 19388 20410 19440
rect 21453 19431 21511 19437
rect 21453 19397 21465 19431
rect 21499 19428 21511 19431
rect 21634 19428 21640 19440
rect 21499 19400 21640 19428
rect 21499 19397 21511 19400
rect 21453 19391 21511 19397
rect 21634 19388 21640 19400
rect 21692 19388 21698 19440
rect 25332 19428 25360 19468
rect 25406 19456 25412 19508
rect 25464 19456 25470 19508
rect 26694 19456 26700 19508
rect 26752 19496 26758 19508
rect 26789 19499 26847 19505
rect 26789 19496 26801 19499
rect 26752 19468 26801 19496
rect 26752 19456 26758 19468
rect 26789 19465 26801 19468
rect 26835 19465 26847 19499
rect 28718 19496 28724 19508
rect 26789 19459 26847 19465
rect 27080 19468 28724 19496
rect 27080 19428 27108 19468
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 28810 19456 28816 19508
rect 28868 19496 28874 19508
rect 30006 19496 30012 19508
rect 28868 19468 30012 19496
rect 28868 19456 28874 19468
rect 30006 19456 30012 19468
rect 30064 19456 30070 19508
rect 24320 19400 24900 19428
rect 25332 19400 27108 19428
rect 13722 19320 13728 19372
rect 13780 19320 13786 19372
rect 13924 19332 14228 19360
rect 13403 19264 13492 19292
rect 13403 19261 13415 19264
rect 13357 19255 13415 19261
rect 13538 19252 13544 19304
rect 13596 19252 13602 19304
rect 13630 19252 13636 19304
rect 13688 19252 13694 19304
rect 13740 19292 13768 19320
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13740 19264 13829 19292
rect 13817 19261 13829 19264
rect 13863 19292 13875 19295
rect 13924 19292 13952 19332
rect 14090 19301 14096 19304
rect 13863 19264 13952 19292
rect 14047 19295 14096 19301
rect 13863 19261 13875 19264
rect 13817 19255 13875 19261
rect 14047 19261 14059 19295
rect 14093 19261 14096 19295
rect 14047 19255 14096 19261
rect 14090 19252 14096 19255
rect 14148 19252 14154 19304
rect 14200 19292 14228 19332
rect 14734 19320 14740 19372
rect 14792 19360 14798 19372
rect 18414 19360 18420 19372
rect 14792 19332 18420 19360
rect 14792 19320 14798 19332
rect 16316 19301 16344 19332
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 21910 19320 21916 19372
rect 21968 19360 21974 19372
rect 24320 19360 24348 19400
rect 21968 19332 24348 19360
rect 21968 19320 21974 19332
rect 16301 19295 16359 19301
rect 14200 19264 15700 19292
rect 13265 19227 13323 19233
rect 13265 19193 13277 19227
rect 13311 19224 13323 19227
rect 13446 19224 13452 19236
rect 13311 19196 13452 19224
rect 13311 19193 13323 19196
rect 13265 19187 13323 19193
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 13722 19184 13728 19236
rect 13780 19224 13786 19236
rect 13909 19227 13967 19233
rect 13909 19224 13921 19227
rect 13780 19196 13921 19224
rect 13780 19184 13786 19196
rect 13909 19193 13921 19196
rect 13955 19224 13967 19227
rect 15562 19224 15568 19236
rect 13955 19196 15568 19224
rect 13955 19193 13967 19196
rect 13909 19187 13967 19193
rect 15562 19184 15568 19196
rect 15620 19184 15626 19236
rect 15672 19224 15700 19264
rect 16301 19261 16313 19295
rect 16347 19261 16359 19295
rect 16301 19255 16359 19261
rect 16390 19252 16396 19304
rect 16448 19292 16454 19304
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 16448 19264 16497 19292
rect 16448 19252 16454 19264
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 16666 19252 16672 19304
rect 16724 19292 16730 19304
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 16724 19264 17325 19292
rect 16724 19252 16730 19264
rect 17313 19261 17325 19264
rect 17359 19261 17371 19295
rect 17313 19255 17371 19261
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 17681 19295 17739 19301
rect 17681 19292 17693 19295
rect 17644 19264 17693 19292
rect 17644 19252 17650 19264
rect 17681 19261 17693 19264
rect 17727 19261 17739 19295
rect 20346 19292 20352 19304
rect 17681 19255 17739 19261
rect 17787 19264 20352 19292
rect 17787 19224 17815 19264
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20530 19252 20536 19304
rect 20588 19252 20594 19304
rect 20714 19252 20720 19304
rect 20772 19252 20778 19304
rect 20806 19252 20812 19304
rect 20864 19252 20870 19304
rect 20898 19252 20904 19304
rect 20956 19252 20962 19304
rect 21269 19295 21327 19301
rect 21269 19261 21281 19295
rect 21315 19292 21327 19295
rect 21450 19292 21456 19304
rect 21315 19264 21456 19292
rect 21315 19261 21327 19264
rect 21269 19255 21327 19261
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 23750 19292 23756 19304
rect 23707 19264 23756 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 23750 19252 23756 19264
rect 23808 19252 23814 19304
rect 23842 19252 23848 19304
rect 23900 19292 23906 19304
rect 24029 19295 24087 19301
rect 24029 19292 24041 19295
rect 23900 19264 24041 19292
rect 23900 19252 23906 19264
rect 24029 19261 24041 19264
rect 24075 19292 24087 19295
rect 24210 19292 24216 19304
rect 24075 19264 24216 19292
rect 24075 19261 24087 19264
rect 24029 19255 24087 19261
rect 24210 19252 24216 19264
rect 24268 19252 24274 19304
rect 24320 19301 24348 19332
rect 24872 19304 24900 19400
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19261 24363 19295
rect 24305 19255 24363 19261
rect 24394 19252 24400 19304
rect 24452 19301 24458 19304
rect 24452 19255 24464 19301
rect 24452 19252 24458 19255
rect 24854 19252 24860 19304
rect 24912 19252 24918 19304
rect 25038 19252 25044 19304
rect 25096 19252 25102 19304
rect 25133 19295 25191 19301
rect 25133 19261 25145 19295
rect 25179 19292 25191 19295
rect 25222 19292 25228 19304
rect 25179 19264 25228 19292
rect 25179 19261 25191 19264
rect 25133 19255 25191 19261
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 25317 19295 25375 19301
rect 25317 19261 25329 19295
rect 25363 19292 25375 19295
rect 25406 19292 25412 19304
rect 25363 19264 25412 19292
rect 25363 19261 25375 19264
rect 25317 19255 25375 19261
rect 25406 19252 25412 19264
rect 25464 19252 25470 19304
rect 25608 19301 25636 19400
rect 28258 19388 28264 19440
rect 28316 19428 28322 19440
rect 28902 19428 28908 19440
rect 28316 19400 28908 19428
rect 28316 19388 28322 19400
rect 28902 19388 28908 19400
rect 28960 19388 28966 19440
rect 26237 19363 26295 19369
rect 26237 19329 26249 19363
rect 26283 19360 26295 19363
rect 27798 19360 27804 19372
rect 26283 19332 27804 19360
rect 26283 19329 26295 19332
rect 26237 19323 26295 19329
rect 27798 19320 27804 19332
rect 27856 19320 27862 19372
rect 27982 19320 27988 19372
rect 28040 19360 28046 19372
rect 28040 19332 30420 19360
rect 28040 19320 28046 19332
rect 25593 19295 25651 19301
rect 25593 19261 25605 19295
rect 25639 19261 25651 19295
rect 25593 19255 25651 19261
rect 25682 19252 25688 19304
rect 25740 19252 25746 19304
rect 25774 19252 25780 19304
rect 25832 19252 25838 19304
rect 25869 19295 25927 19301
rect 25869 19261 25881 19295
rect 25915 19292 25927 19295
rect 25958 19292 25964 19304
rect 25915 19264 25964 19292
rect 25915 19261 25927 19264
rect 25869 19255 25927 19261
rect 25958 19252 25964 19264
rect 26016 19252 26022 19304
rect 26326 19252 26332 19304
rect 26384 19252 26390 19304
rect 26973 19295 27031 19301
rect 26973 19261 26985 19295
rect 27019 19261 27031 19295
rect 28368 19278 28396 19332
rect 26973 19255 27031 19261
rect 15672 19196 17815 19224
rect 18046 19184 18052 19236
rect 18104 19224 18110 19236
rect 18506 19224 18512 19236
rect 18104 19196 18512 19224
rect 18104 19184 18110 19196
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 18782 19184 18788 19236
rect 18840 19224 18846 19236
rect 19794 19224 19800 19236
rect 18840 19196 19800 19224
rect 18840 19184 18846 19196
rect 19794 19184 19800 19196
rect 19852 19184 19858 19236
rect 20441 19227 20499 19233
rect 20441 19193 20453 19227
rect 20487 19224 20499 19227
rect 21358 19224 21364 19236
rect 20487 19196 21364 19224
rect 20487 19193 20499 19196
rect 20441 19187 20499 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 21634 19184 21640 19236
rect 21692 19184 21698 19236
rect 22830 19184 22836 19236
rect 22888 19184 22894 19236
rect 23106 19184 23112 19236
rect 23164 19224 23170 19236
rect 23385 19227 23443 19233
rect 23385 19224 23397 19227
rect 23164 19196 23397 19224
rect 23164 19184 23170 19196
rect 23385 19193 23397 19196
rect 23431 19193 23443 19227
rect 23385 19187 23443 19193
rect 24118 19184 24124 19236
rect 24176 19224 24182 19236
rect 24762 19224 24768 19236
rect 24176 19196 24768 19224
rect 24176 19184 24182 19196
rect 24762 19184 24768 19196
rect 24820 19184 24826 19236
rect 26234 19184 26240 19236
rect 26292 19224 26298 19236
rect 26421 19227 26479 19233
rect 26421 19224 26433 19227
rect 26292 19196 26433 19224
rect 26292 19184 26298 19196
rect 26421 19193 26433 19196
rect 26467 19224 26479 19227
rect 26786 19224 26792 19236
rect 26467 19196 26792 19224
rect 26467 19193 26479 19196
rect 26421 19187 26479 19193
rect 26786 19184 26792 19196
rect 26844 19184 26850 19236
rect 26988 19224 27016 19255
rect 28994 19252 29000 19304
rect 29052 19252 29058 19304
rect 30392 19292 30420 19332
rect 30558 19292 30564 19304
rect 30392 19278 30564 19292
rect 30406 19264 30564 19278
rect 30558 19252 30564 19264
rect 30616 19252 30622 19304
rect 27249 19227 27307 19233
rect 26988 19196 27108 19224
rect 12391 19128 13216 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 19610 19156 19616 19168
rect 15160 19128 19616 19156
rect 15160 19116 15166 19128
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 21082 19156 21088 19168
rect 20312 19128 21088 19156
rect 20312 19116 20318 19128
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 24673 19159 24731 19165
rect 24673 19156 24685 19159
rect 22152 19128 24685 19156
rect 22152 19116 22158 19128
rect 24673 19125 24685 19128
rect 24719 19156 24731 19159
rect 24946 19156 24952 19168
rect 24719 19128 24952 19156
rect 24719 19125 24731 19128
rect 24673 19119 24731 19125
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 25314 19116 25320 19168
rect 25372 19116 25378 19168
rect 27080 19156 27108 19196
rect 27249 19193 27261 19227
rect 27295 19224 27307 19227
rect 27338 19224 27344 19236
rect 27295 19196 27344 19224
rect 27295 19193 27307 19196
rect 27249 19187 27307 19193
rect 27338 19184 27344 19196
rect 27396 19184 27402 19236
rect 28644 19196 29224 19224
rect 27522 19156 27528 19168
rect 27080 19128 27528 19156
rect 27522 19116 27528 19128
rect 27580 19116 27586 19168
rect 27614 19116 27620 19168
rect 27672 19156 27678 19168
rect 28644 19156 28672 19196
rect 27672 19128 28672 19156
rect 28721 19159 28779 19165
rect 27672 19116 27678 19128
rect 28721 19125 28733 19159
rect 28767 19156 28779 19159
rect 28810 19156 28816 19168
rect 28767 19128 28816 19156
rect 28767 19125 28779 19128
rect 28721 19119 28779 19125
rect 28810 19116 28816 19128
rect 28868 19116 28874 19168
rect 29196 19156 29224 19196
rect 29270 19184 29276 19236
rect 29328 19184 29334 19236
rect 30837 19227 30895 19233
rect 30837 19224 30849 19227
rect 30576 19196 30849 19224
rect 30576 19156 30604 19196
rect 30837 19193 30849 19196
rect 30883 19193 30895 19227
rect 30837 19187 30895 19193
rect 31018 19184 31024 19236
rect 31076 19184 31082 19236
rect 31110 19184 31116 19236
rect 31168 19224 31174 19236
rect 31205 19227 31263 19233
rect 31205 19224 31217 19227
rect 31168 19196 31217 19224
rect 31168 19184 31174 19196
rect 31205 19193 31217 19196
rect 31251 19193 31263 19227
rect 31205 19187 31263 19193
rect 29196 19128 30604 19156
rect 30742 19116 30748 19168
rect 30800 19116 30806 19168
rect 552 19066 31648 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 12096 19066
rect 12148 19014 12160 19066
rect 12212 19014 12224 19066
rect 12276 19014 12288 19066
rect 12340 19014 12352 19066
rect 12404 19014 19870 19066
rect 19922 19014 19934 19066
rect 19986 19014 19998 19066
rect 20050 19014 20062 19066
rect 20114 19014 20126 19066
rect 20178 19014 27644 19066
rect 27696 19014 27708 19066
rect 27760 19014 27772 19066
rect 27824 19014 27836 19066
rect 27888 19014 27900 19066
rect 27952 19014 31648 19066
rect 552 18992 31648 19014
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 8757 18955 8815 18961
rect 5500 18924 7604 18952
rect 5500 18912 5506 18924
rect 3436 18856 3648 18884
rect 3436 18828 3464 18856
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 3418 18816 3424 18828
rect 3375 18788 3424 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 3418 18776 3424 18788
rect 3476 18776 3482 18828
rect 3620 18825 3648 18856
rect 3804 18856 4016 18884
rect 3804 18825 3832 18856
rect 3513 18819 3571 18825
rect 3513 18785 3525 18819
rect 3559 18785 3571 18819
rect 3513 18779 3571 18785
rect 3605 18819 3663 18825
rect 3605 18785 3617 18819
rect 3651 18785 3663 18819
rect 3605 18779 3663 18785
rect 3789 18819 3847 18825
rect 3789 18785 3801 18819
rect 3835 18785 3847 18819
rect 3789 18779 3847 18785
rect 3234 18640 3240 18692
rect 3292 18640 3298 18692
rect 3528 18680 3556 18779
rect 3878 18776 3884 18828
rect 3936 18776 3942 18828
rect 3988 18816 4016 18856
rect 4062 18844 4068 18896
rect 4120 18884 4126 18896
rect 5169 18887 5227 18893
rect 4120 18856 5120 18884
rect 4120 18844 4126 18856
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3988 18788 4445 18816
rect 4433 18785 4445 18788
rect 4479 18816 4491 18819
rect 4890 18816 4896 18828
rect 4479 18788 4896 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 5092 18825 5120 18856
rect 5169 18853 5181 18887
rect 5215 18884 5227 18887
rect 6086 18884 6092 18896
rect 5215 18856 6092 18884
rect 5215 18853 5227 18856
rect 5169 18847 5227 18853
rect 6086 18844 6092 18856
rect 6144 18884 6150 18896
rect 6457 18887 6515 18893
rect 6457 18884 6469 18887
rect 6144 18856 6469 18884
rect 6144 18844 6150 18856
rect 6457 18853 6469 18856
rect 6503 18853 6515 18887
rect 6457 18847 6515 18853
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18785 5135 18819
rect 5077 18779 5135 18785
rect 5258 18776 5264 18828
rect 5316 18776 5322 18828
rect 5350 18776 5356 18828
rect 5408 18816 5414 18828
rect 5905 18819 5963 18825
rect 5905 18816 5917 18819
rect 5408 18788 5917 18816
rect 5408 18776 5414 18788
rect 5905 18785 5917 18788
rect 5951 18816 5963 18819
rect 5951 18788 6132 18816
rect 5951 18785 5963 18788
rect 5905 18779 5963 18785
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18748 4031 18751
rect 5994 18748 6000 18760
rect 4019 18720 6000 18748
rect 4019 18717 4031 18720
rect 3973 18711 4031 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 6104 18748 6132 18788
rect 6178 18776 6184 18828
rect 6236 18776 6242 18828
rect 6917 18819 6975 18825
rect 6288 18788 6868 18816
rect 6288 18748 6316 18788
rect 6104 18720 6316 18748
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6512 18720 6745 18748
rect 6512 18708 6518 18720
rect 6733 18717 6745 18720
rect 6779 18717 6791 18751
rect 6840 18748 6868 18788
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 7006 18816 7012 18828
rect 6963 18788 7012 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7469 18819 7527 18825
rect 7469 18785 7481 18819
rect 7515 18785 7527 18819
rect 7576 18816 7604 18924
rect 8757 18921 8769 18955
rect 8803 18952 8815 18955
rect 12161 18955 12219 18961
rect 8803 18924 11928 18952
rect 8803 18921 8815 18924
rect 8757 18915 8815 18921
rect 7653 18887 7711 18893
rect 7653 18853 7665 18887
rect 7699 18884 7711 18887
rect 10137 18887 10195 18893
rect 10137 18884 10149 18887
rect 7699 18856 10149 18884
rect 7699 18853 7711 18856
rect 7653 18847 7711 18853
rect 10137 18853 10149 18856
rect 10183 18884 10195 18887
rect 11238 18884 11244 18896
rect 10183 18856 11244 18884
rect 10183 18853 10195 18856
rect 10137 18847 10195 18853
rect 11238 18844 11244 18856
rect 11296 18844 11302 18896
rect 11900 18884 11928 18924
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 12434 18952 12440 18964
rect 12207 18924 12440 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 13179 18955 13237 18961
rect 13179 18921 13191 18955
rect 13225 18952 13237 18955
rect 13630 18952 13636 18964
rect 13225 18924 13636 18952
rect 13225 18921 13237 18924
rect 13179 18915 13237 18921
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 15657 18955 15715 18961
rect 15657 18921 15669 18955
rect 15703 18952 15715 18955
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15703 18924 16129 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16666 18952 16672 18964
rect 16117 18915 16175 18921
rect 16224 18924 16672 18952
rect 12805 18887 12863 18893
rect 12805 18884 12817 18887
rect 11900 18856 12817 18884
rect 12805 18853 12817 18856
rect 12851 18884 12863 18887
rect 13265 18887 13323 18893
rect 13265 18884 13277 18887
rect 12851 18856 13277 18884
rect 12851 18853 12863 18856
rect 12805 18847 12863 18853
rect 13265 18853 13277 18856
rect 13311 18853 13323 18887
rect 13446 18884 13452 18896
rect 13265 18847 13323 18853
rect 13372 18856 13452 18884
rect 8297 18819 8355 18825
rect 8297 18816 8309 18819
rect 7576 18788 8309 18816
rect 7469 18779 7527 18785
rect 8297 18785 8309 18788
rect 8343 18785 8355 18819
rect 8297 18779 8355 18785
rect 7098 18748 7104 18760
rect 6840 18720 7104 18748
rect 6733 18711 6791 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 7193 18751 7251 18757
rect 7193 18717 7205 18751
rect 7239 18748 7251 18751
rect 7374 18748 7380 18760
rect 7239 18720 7380 18748
rect 7239 18717 7251 18720
rect 7193 18711 7251 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 3528 18652 4384 18680
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 4356 18621 4384 18652
rect 5902 18640 5908 18692
rect 5960 18680 5966 18692
rect 6822 18680 6828 18692
rect 5960 18652 6828 18680
rect 5960 18640 5966 18652
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 7484 18624 7512 18779
rect 8312 18748 8340 18779
rect 8386 18776 8392 18828
rect 8444 18776 8450 18828
rect 8570 18776 8576 18828
rect 8628 18776 8634 18828
rect 8938 18776 8944 18828
rect 8996 18822 9002 18828
rect 9033 18822 9091 18825
rect 8996 18819 9091 18822
rect 8996 18794 9045 18819
rect 8996 18776 9002 18794
rect 9033 18785 9045 18794
rect 9079 18785 9091 18819
rect 9033 18779 9091 18785
rect 9214 18776 9220 18828
rect 9272 18776 9278 18828
rect 9306 18776 9312 18828
rect 9364 18776 9370 18828
rect 9858 18776 9864 18828
rect 9916 18776 9922 18828
rect 9950 18776 9956 18828
rect 10008 18776 10014 18828
rect 10226 18776 10232 18828
rect 10284 18776 10290 18828
rect 10321 18819 10379 18825
rect 10321 18785 10333 18819
rect 10367 18816 10379 18819
rect 11054 18816 11060 18828
rect 10367 18788 11060 18816
rect 10367 18785 10379 18788
rect 10321 18779 10379 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 11204 18788 11345 18816
rect 11204 18776 11210 18788
rect 11333 18785 11345 18788
rect 11379 18785 11391 18819
rect 11333 18779 11391 18785
rect 11517 18819 11575 18825
rect 11517 18785 11529 18819
rect 11563 18816 11575 18819
rect 12158 18816 12164 18828
rect 11563 18788 12164 18816
rect 11563 18785 11575 18788
rect 11517 18779 11575 18785
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 13078 18776 13084 18828
rect 13136 18776 13142 18828
rect 13372 18825 13400 18856
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 15565 18887 15623 18893
rect 15565 18853 15577 18887
rect 15611 18884 15623 18887
rect 16224 18884 16252 18924
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 18046 18952 18052 18964
rect 17052 18924 18052 18952
rect 16298 18893 16304 18896
rect 15611 18856 16252 18884
rect 16285 18887 16304 18893
rect 15611 18853 15623 18856
rect 15565 18847 15623 18853
rect 16285 18853 16297 18887
rect 16285 18847 16304 18853
rect 16298 18844 16304 18847
rect 16356 18844 16362 18896
rect 16485 18887 16543 18893
rect 16485 18853 16497 18887
rect 16531 18884 16543 18887
rect 17052 18884 17080 18924
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 18472 18924 19533 18952
rect 18472 18912 18478 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 19610 18912 19616 18964
rect 19668 18952 19674 18964
rect 19886 18952 19892 18964
rect 19668 18924 19892 18952
rect 19668 18912 19674 18924
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 20165 18955 20223 18961
rect 20165 18921 20177 18955
rect 20211 18952 20223 18955
rect 20530 18952 20536 18964
rect 20211 18924 20536 18952
rect 20211 18921 20223 18924
rect 20165 18915 20223 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21545 18955 21603 18961
rect 21545 18952 21557 18955
rect 20956 18924 21557 18952
rect 20956 18912 20962 18924
rect 21545 18921 21557 18924
rect 21591 18921 21603 18955
rect 21545 18915 21603 18921
rect 22281 18955 22339 18961
rect 22281 18921 22293 18955
rect 22327 18952 22339 18955
rect 23106 18952 23112 18964
rect 22327 18924 23112 18952
rect 22327 18921 22339 18924
rect 22281 18915 22339 18921
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 23750 18912 23756 18964
rect 23808 18952 23814 18964
rect 25777 18955 25835 18961
rect 23808 18924 24900 18952
rect 23808 18912 23814 18924
rect 16531 18856 17080 18884
rect 16531 18853 16543 18856
rect 16485 18847 16543 18853
rect 17126 18844 17132 18896
rect 17184 18844 17190 18896
rect 18138 18844 18144 18896
rect 18196 18844 18202 18896
rect 18782 18844 18788 18896
rect 18840 18884 18846 18896
rect 18969 18887 19027 18893
rect 18969 18884 18981 18887
rect 18840 18856 18981 18884
rect 18840 18844 18846 18856
rect 18969 18853 18981 18856
rect 19015 18853 19027 18887
rect 18969 18847 19027 18853
rect 19058 18844 19064 18896
rect 19116 18884 19122 18896
rect 19797 18887 19855 18893
rect 19797 18884 19809 18887
rect 19116 18856 19809 18884
rect 19116 18844 19122 18856
rect 19797 18853 19809 18856
rect 19843 18853 19855 18887
rect 19797 18847 19855 18853
rect 19981 18887 20039 18893
rect 19981 18853 19993 18887
rect 20027 18884 20039 18887
rect 23290 18884 23296 18896
rect 20027 18856 22140 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 13357 18819 13415 18825
rect 13357 18785 13369 18819
rect 13403 18785 13415 18819
rect 13357 18779 13415 18785
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14274 18816 14280 18828
rect 14148 18788 14280 18816
rect 14148 18776 14154 18788
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 16574 18776 16580 18828
rect 16632 18776 16638 18828
rect 16758 18776 16764 18828
rect 16816 18776 16822 18828
rect 19996 18816 20024 18847
rect 19352 18788 20024 18816
rect 9876 18748 9904 18776
rect 8312 18720 9904 18748
rect 10980 18720 11750 18748
rect 8481 18683 8539 18689
rect 8481 18649 8493 18683
rect 8527 18680 8539 18683
rect 8849 18683 8907 18689
rect 8849 18680 8861 18683
rect 8527 18652 8861 18680
rect 8527 18649 8539 18652
rect 8481 18643 8539 18649
rect 8849 18649 8861 18652
rect 8895 18649 8907 18683
rect 10980 18680 11008 18720
rect 8849 18643 8907 18649
rect 8956 18652 11008 18680
rect 8956 18624 8984 18652
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 11330 18680 11336 18692
rect 11112 18652 11336 18680
rect 11112 18640 11118 18652
rect 11330 18640 11336 18652
rect 11388 18640 11394 18692
rect 11722 18680 11750 18720
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 11974 18748 11980 18760
rect 11848 18720 11980 18748
rect 11848 18708 11854 18720
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 12066 18708 12072 18760
rect 12124 18748 12130 18760
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 12124 18720 12357 18748
rect 12124 18708 12130 18720
rect 12345 18717 12357 18720
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12437 18751 12495 18757
rect 12437 18717 12449 18751
rect 12483 18748 12495 18751
rect 14458 18748 14464 18760
rect 12483 18720 14464 18748
rect 12483 18717 12495 18720
rect 12437 18711 12495 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 15746 18748 15752 18760
rect 14608 18720 15752 18748
rect 14608 18708 14614 18720
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 16482 18708 16488 18760
rect 16540 18748 16546 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16540 18720 16865 18748
rect 16540 18708 16546 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 19242 18748 19248 18760
rect 18656 18720 19248 18748
rect 18656 18708 18662 18720
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 16390 18680 16396 18692
rect 11722 18652 16396 18680
rect 16390 18640 16396 18652
rect 16448 18640 16454 18692
rect 18432 18652 18828 18680
rect 3697 18615 3755 18621
rect 3697 18612 3709 18615
rect 3568 18584 3709 18612
rect 3568 18572 3574 18584
rect 3697 18581 3709 18584
rect 3743 18581 3755 18615
rect 3697 18575 3755 18581
rect 4341 18615 4399 18621
rect 4341 18581 4353 18615
rect 4387 18612 4399 18615
rect 6638 18612 6644 18624
rect 4387 18584 6644 18612
rect 4387 18581 4399 18584
rect 4341 18575 4399 18581
rect 6638 18572 6644 18584
rect 6696 18572 6702 18624
rect 7101 18615 7159 18621
rect 7101 18581 7113 18615
rect 7147 18612 7159 18615
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 7147 18584 7297 18612
rect 7147 18581 7159 18584
rect 7101 18575 7159 18581
rect 7285 18581 7297 18584
rect 7331 18581 7343 18615
rect 7285 18575 7343 18581
rect 7466 18572 7472 18624
rect 7524 18612 7530 18624
rect 8938 18612 8944 18624
rect 7524 18584 8944 18612
rect 7524 18572 7530 18584
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 10505 18615 10563 18621
rect 10505 18581 10517 18615
rect 10551 18612 10563 18615
rect 11146 18612 11152 18624
rect 10551 18584 11152 18612
rect 10551 18581 10563 18584
rect 10505 18575 10563 18581
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 11701 18615 11759 18621
rect 11701 18581 11713 18615
rect 11747 18612 11759 18615
rect 11790 18612 11796 18624
rect 11747 18584 11796 18612
rect 11747 18581 11759 18584
rect 11701 18575 11759 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 14734 18612 14740 18624
rect 12216 18584 14740 18612
rect 12216 18572 12222 18584
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 15197 18615 15255 18621
rect 15197 18612 15209 18615
rect 14976 18584 15209 18612
rect 14976 18572 14982 18584
rect 15197 18581 15209 18584
rect 15243 18581 15255 18615
rect 15197 18575 15255 18581
rect 16206 18572 16212 18624
rect 16264 18612 16270 18624
rect 16301 18615 16359 18621
rect 16301 18612 16313 18615
rect 16264 18584 16313 18612
rect 16264 18572 16270 18584
rect 16301 18581 16313 18584
rect 16347 18581 16359 18615
rect 16301 18575 16359 18581
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 18432 18612 18460 18652
rect 16632 18584 18460 18612
rect 16632 18572 16638 18584
rect 18506 18572 18512 18624
rect 18564 18612 18570 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18564 18584 18613 18612
rect 18564 18572 18570 18584
rect 18601 18581 18613 18584
rect 18647 18581 18659 18615
rect 18800 18612 18828 18652
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 18969 18683 19027 18689
rect 18969 18680 18981 18683
rect 18932 18652 18981 18680
rect 18932 18640 18938 18652
rect 18969 18649 18981 18652
rect 19015 18680 19027 18683
rect 19352 18680 19380 18788
rect 20254 18776 20260 18828
rect 20312 18776 20318 18828
rect 20346 18776 20352 18828
rect 20404 18816 20410 18828
rect 20717 18819 20775 18825
rect 20404 18788 20668 18816
rect 20404 18776 20410 18788
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19015 18652 19380 18680
rect 19444 18680 19472 18711
rect 19518 18708 19524 18760
rect 19576 18748 19582 18760
rect 20070 18748 20076 18760
rect 19576 18720 20076 18748
rect 19576 18708 19582 18720
rect 20070 18708 20076 18720
rect 20128 18708 20134 18760
rect 20533 18751 20591 18757
rect 20533 18748 20545 18751
rect 20180 18720 20545 18748
rect 19610 18680 19616 18692
rect 19444 18652 19616 18680
rect 19015 18649 19027 18652
rect 18969 18643 19027 18649
rect 19610 18640 19616 18652
rect 19668 18640 19674 18692
rect 19705 18683 19763 18689
rect 19705 18649 19717 18683
rect 19751 18680 19763 18683
rect 19978 18680 19984 18692
rect 19751 18652 19984 18680
rect 19751 18649 19763 18652
rect 19705 18643 19763 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 20180 18612 20208 18720
rect 20533 18717 20545 18720
rect 20579 18717 20591 18751
rect 20640 18748 20668 18788
rect 20717 18785 20729 18819
rect 20763 18816 20775 18819
rect 20806 18816 20812 18828
rect 20763 18788 20812 18816
rect 20763 18785 20775 18788
rect 20717 18779 20775 18785
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 22112 18825 22140 18856
rect 22204 18856 23296 18884
rect 22097 18819 22155 18825
rect 21140 18788 21864 18816
rect 21140 18776 21146 18788
rect 21174 18748 21180 18760
rect 20640 18720 21180 18748
rect 20533 18711 20591 18717
rect 21174 18708 21180 18720
rect 21232 18748 21238 18760
rect 21836 18748 21864 18788
rect 22097 18785 22109 18819
rect 22143 18785 22155 18819
rect 22097 18779 22155 18785
rect 22204 18748 22232 18856
rect 23290 18844 23296 18856
rect 23348 18844 23354 18896
rect 24026 18844 24032 18896
rect 24084 18844 24090 18896
rect 22738 18776 22744 18828
rect 22796 18776 22802 18828
rect 24872 18825 24900 18924
rect 25777 18921 25789 18955
rect 25823 18952 25835 18955
rect 25866 18952 25872 18964
rect 25823 18924 25872 18952
rect 25823 18921 25835 18924
rect 25777 18915 25835 18921
rect 25866 18912 25872 18924
rect 25924 18912 25930 18964
rect 27706 18952 27712 18964
rect 25976 18924 27712 18952
rect 25222 18844 25228 18896
rect 25280 18884 25286 18896
rect 25976 18884 26004 18924
rect 27706 18912 27712 18924
rect 27764 18912 27770 18964
rect 29178 18912 29184 18964
rect 29236 18952 29242 18964
rect 29365 18955 29423 18961
rect 29365 18952 29377 18955
rect 29236 18924 29377 18952
rect 29236 18912 29242 18924
rect 29365 18921 29377 18924
rect 29411 18921 29423 18955
rect 29365 18915 29423 18921
rect 29825 18955 29883 18961
rect 29825 18921 29837 18955
rect 29871 18952 29883 18955
rect 29914 18952 29920 18964
rect 29871 18924 29920 18952
rect 29871 18921 29883 18924
rect 29825 18915 29883 18921
rect 29914 18912 29920 18924
rect 29972 18912 29978 18964
rect 30006 18912 30012 18964
rect 30064 18952 30070 18964
rect 30742 18952 30748 18964
rect 30064 18924 30748 18952
rect 30064 18912 30070 18924
rect 25280 18856 26004 18884
rect 25280 18844 25286 18856
rect 26418 18844 26424 18896
rect 26476 18844 26482 18896
rect 28813 18887 28871 18893
rect 28813 18884 28825 18887
rect 28000 18856 28825 18884
rect 24857 18819 24915 18825
rect 24857 18785 24869 18819
rect 24903 18785 24915 18819
rect 24857 18779 24915 18785
rect 24949 18819 25007 18825
rect 24949 18785 24961 18819
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 21232 18720 21772 18748
rect 21836 18720 22232 18748
rect 22465 18751 22523 18757
rect 21232 18708 21238 18720
rect 20346 18640 20352 18692
rect 20404 18640 20410 18692
rect 20441 18683 20499 18689
rect 20441 18649 20453 18683
rect 20487 18680 20499 18683
rect 21634 18680 21640 18692
rect 20487 18652 21640 18680
rect 20487 18649 20499 18652
rect 20441 18643 20499 18649
rect 21634 18640 21640 18652
rect 21692 18640 21698 18692
rect 21744 18680 21772 18720
rect 22465 18717 22477 18751
rect 22511 18717 22523 18751
rect 22465 18711 22523 18717
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 22480 18680 22508 18711
rect 21744 18652 22508 18680
rect 22572 18680 22600 18711
rect 22646 18708 22652 18760
rect 22704 18708 22710 18760
rect 23382 18708 23388 18760
rect 23440 18748 23446 18760
rect 24026 18748 24032 18760
rect 23440 18720 24032 18748
rect 23440 18708 23446 18720
rect 24026 18708 24032 18720
rect 24084 18708 24090 18760
rect 24486 18708 24492 18760
rect 24544 18748 24550 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24544 18720 24593 18748
rect 24544 18708 24550 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24964 18748 24992 18779
rect 25038 18776 25044 18828
rect 25096 18816 25102 18828
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 25096 18788 25145 18816
rect 25096 18776 25102 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 25317 18819 25375 18825
rect 25317 18785 25329 18819
rect 25363 18816 25375 18819
rect 25685 18819 25743 18825
rect 25685 18816 25697 18819
rect 25363 18788 25697 18816
rect 25363 18785 25375 18788
rect 25317 18779 25375 18785
rect 25685 18785 25697 18788
rect 25731 18816 25743 18819
rect 27890 18816 27896 18828
rect 25731 18788 27896 18816
rect 25731 18785 25743 18788
rect 25685 18779 25743 18785
rect 26436 18760 26464 18788
rect 27890 18776 27896 18788
rect 27948 18776 27954 18828
rect 25406 18748 25412 18760
rect 24581 18711 24639 18717
rect 24872 18720 25412 18748
rect 24872 18692 24900 18720
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 25498 18708 25504 18760
rect 25556 18708 25562 18760
rect 26418 18708 26424 18760
rect 26476 18708 26482 18760
rect 27338 18708 27344 18760
rect 27396 18748 27402 18760
rect 28000 18748 28028 18856
rect 28813 18853 28825 18856
rect 28859 18853 28871 18887
rect 28813 18847 28871 18853
rect 29086 18844 29092 18896
rect 29144 18884 29150 18896
rect 29549 18887 29607 18893
rect 29549 18884 29561 18887
rect 29144 18856 29561 18884
rect 29144 18844 29150 18856
rect 29549 18853 29561 18856
rect 29595 18853 29607 18887
rect 29549 18847 29607 18853
rect 29638 18844 29644 18896
rect 29696 18884 29702 18896
rect 30469 18887 30527 18893
rect 30469 18884 30481 18887
rect 29696 18856 30481 18884
rect 29696 18844 29702 18856
rect 30469 18853 30481 18856
rect 30515 18853 30527 18887
rect 30469 18847 30527 18853
rect 28074 18776 28080 18828
rect 28132 18816 28138 18828
rect 28537 18819 28595 18825
rect 28537 18816 28549 18819
rect 28132 18788 28549 18816
rect 28132 18776 28138 18788
rect 28537 18785 28549 18788
rect 28583 18785 28595 18819
rect 28537 18779 28595 18785
rect 29181 18822 29239 18825
rect 29270 18822 29276 18828
rect 29181 18819 29276 18822
rect 29181 18785 29193 18819
rect 29227 18794 29276 18819
rect 29227 18785 29239 18794
rect 29181 18779 29239 18785
rect 28261 18751 28319 18757
rect 28261 18748 28273 18751
rect 27396 18720 28273 18748
rect 27396 18708 27402 18720
rect 28261 18717 28273 18720
rect 28307 18717 28319 18751
rect 28552 18748 28580 18779
rect 29270 18776 29276 18794
rect 29328 18776 29334 18828
rect 29730 18776 29736 18828
rect 29788 18776 29794 18828
rect 30282 18776 30288 18828
rect 30340 18776 30346 18828
rect 30576 18816 30604 18924
rect 30742 18912 30748 18924
rect 30800 18912 30806 18964
rect 30834 18912 30840 18964
rect 30892 18952 30898 18964
rect 30892 18924 31248 18952
rect 30892 18912 30898 18924
rect 31018 18884 31024 18896
rect 30852 18856 31024 18884
rect 30852 18825 30880 18856
rect 31018 18844 31024 18856
rect 31076 18844 31082 18896
rect 30653 18819 30711 18825
rect 30653 18816 30665 18819
rect 30576 18788 30665 18816
rect 30653 18785 30665 18788
rect 30699 18785 30711 18819
rect 30653 18779 30711 18785
rect 30837 18819 30895 18825
rect 30837 18785 30849 18819
rect 30883 18785 30895 18819
rect 30837 18779 30895 18785
rect 30929 18819 30987 18825
rect 30929 18785 30941 18819
rect 30975 18816 30987 18819
rect 31110 18816 31116 18828
rect 30975 18788 31116 18816
rect 30975 18785 30987 18788
rect 30929 18779 30987 18785
rect 28552 18720 29776 18748
rect 28261 18711 28319 18717
rect 22572 18652 23244 18680
rect 20898 18612 20904 18624
rect 18800 18584 20904 18612
rect 18601 18575 18659 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 20993 18615 21051 18621
rect 20993 18581 21005 18615
rect 21039 18612 21051 18615
rect 21450 18612 21456 18624
rect 21039 18584 21456 18612
rect 21039 18581 21051 18584
rect 20993 18575 21051 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 21542 18572 21548 18624
rect 21600 18612 21606 18624
rect 22572 18612 22600 18652
rect 21600 18584 22600 18612
rect 21600 18572 21606 18584
rect 23106 18572 23112 18624
rect 23164 18572 23170 18624
rect 23216 18612 23244 18652
rect 24854 18640 24860 18692
rect 24912 18640 24918 18692
rect 24946 18640 24952 18692
rect 25004 18680 25010 18692
rect 28721 18683 28779 18689
rect 25004 18652 28672 18680
rect 25004 18640 25010 18652
rect 25130 18612 25136 18624
rect 23216 18584 25136 18612
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 26142 18572 26148 18624
rect 26200 18572 26206 18624
rect 27522 18572 27528 18624
rect 27580 18612 27586 18624
rect 27709 18615 27767 18621
rect 27709 18612 27721 18615
rect 27580 18584 27721 18612
rect 27580 18572 27586 18584
rect 27709 18581 27721 18584
rect 27755 18581 27767 18615
rect 27709 18575 27767 18581
rect 28166 18572 28172 18624
rect 28224 18612 28230 18624
rect 28353 18615 28411 18621
rect 28353 18612 28365 18615
rect 28224 18584 28365 18612
rect 28224 18572 28230 18584
rect 28353 18581 28365 18584
rect 28399 18581 28411 18615
rect 28644 18612 28672 18652
rect 28721 18649 28733 18683
rect 28767 18680 28779 18683
rect 29638 18680 29644 18692
rect 28767 18652 29644 18680
rect 28767 18649 28779 18652
rect 28721 18643 28779 18649
rect 29638 18640 29644 18652
rect 29696 18640 29702 18692
rect 29748 18680 29776 18720
rect 29914 18708 29920 18760
rect 29972 18748 29978 18760
rect 30009 18751 30067 18757
rect 30009 18748 30021 18751
rect 29972 18720 30021 18748
rect 29972 18708 29978 18720
rect 30009 18717 30021 18720
rect 30055 18717 30067 18751
rect 30009 18711 30067 18717
rect 30098 18708 30104 18760
rect 30156 18708 30162 18760
rect 30190 18708 30196 18760
rect 30248 18748 30254 18760
rect 30852 18748 30880 18779
rect 31110 18776 31116 18788
rect 31168 18776 31174 18828
rect 30248 18720 30880 18748
rect 30248 18708 30254 18720
rect 31018 18708 31024 18760
rect 31076 18708 31082 18760
rect 30834 18680 30840 18692
rect 29748 18652 30840 18680
rect 30834 18640 30840 18652
rect 30892 18640 30898 18692
rect 31113 18683 31171 18689
rect 31113 18649 31125 18683
rect 31159 18680 31171 18683
rect 31220 18680 31248 18924
rect 31297 18819 31355 18825
rect 31297 18785 31309 18819
rect 31343 18816 31355 18819
rect 31478 18816 31484 18828
rect 31343 18788 31484 18816
rect 31343 18785 31355 18788
rect 31297 18779 31355 18785
rect 31478 18776 31484 18788
rect 31536 18776 31542 18828
rect 31159 18652 31248 18680
rect 31159 18649 31171 18652
rect 31113 18643 31171 18649
rect 31018 18612 31024 18624
rect 28644 18584 31024 18612
rect 28353 18575 28411 18581
rect 31018 18572 31024 18584
rect 31076 18572 31082 18624
rect 31205 18615 31263 18621
rect 31205 18581 31217 18615
rect 31251 18612 31263 18615
rect 31294 18612 31300 18624
rect 31251 18584 31300 18612
rect 31251 18581 31263 18584
rect 31205 18575 31263 18581
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 552 18522 31648 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 11436 18522
rect 11488 18470 11500 18522
rect 11552 18470 11564 18522
rect 11616 18470 11628 18522
rect 11680 18470 11692 18522
rect 11744 18470 19210 18522
rect 19262 18470 19274 18522
rect 19326 18470 19338 18522
rect 19390 18470 19402 18522
rect 19454 18470 19466 18522
rect 19518 18470 26984 18522
rect 27036 18470 27048 18522
rect 27100 18470 27112 18522
rect 27164 18470 27176 18522
rect 27228 18470 27240 18522
rect 27292 18470 31648 18522
rect 552 18448 31648 18470
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 2685 18411 2743 18417
rect 2685 18408 2697 18411
rect 2556 18380 2697 18408
rect 2556 18368 2562 18380
rect 2685 18377 2697 18380
rect 2731 18377 2743 18411
rect 2685 18371 2743 18377
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 7466 18408 7472 18420
rect 5868 18380 7472 18408
rect 5868 18368 5874 18380
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 8662 18408 8668 18420
rect 8076 18380 8668 18408
rect 8076 18368 8082 18380
rect 8662 18368 8668 18380
rect 8720 18408 8726 18420
rect 8757 18411 8815 18417
rect 8757 18408 8769 18411
rect 8720 18380 8769 18408
rect 8720 18368 8726 18380
rect 8757 18377 8769 18380
rect 8803 18377 8815 18411
rect 8757 18371 8815 18377
rect 11238 18368 11244 18420
rect 11296 18368 11302 18420
rect 15378 18408 15384 18420
rect 11348 18380 15384 18408
rect 6822 18300 6828 18352
rect 6880 18340 6886 18352
rect 11348 18340 11376 18380
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 16758 18368 16764 18420
rect 16816 18408 16822 18420
rect 17037 18411 17095 18417
rect 17037 18408 17049 18411
rect 16816 18380 17049 18408
rect 16816 18368 16822 18380
rect 17037 18377 17049 18380
rect 17083 18377 17095 18411
rect 17037 18371 17095 18377
rect 17218 18368 17224 18420
rect 17276 18408 17282 18420
rect 17862 18408 17868 18420
rect 17276 18380 17868 18408
rect 17276 18368 17282 18380
rect 17862 18368 17868 18380
rect 17920 18408 17926 18420
rect 19429 18411 19487 18417
rect 17920 18380 19334 18408
rect 17920 18368 17926 18380
rect 6880 18312 11376 18340
rect 11425 18343 11483 18349
rect 6880 18300 6886 18312
rect 11425 18309 11437 18343
rect 11471 18340 11483 18343
rect 11471 18312 12434 18340
rect 11471 18309 11483 18312
rect 11425 18303 11483 18309
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 4062 18272 4068 18284
rect 2464 18244 4068 18272
rect 2464 18232 2470 18244
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 5166 18232 5172 18284
rect 5224 18272 5230 18284
rect 6270 18272 6276 18284
rect 5224 18244 6276 18272
rect 5224 18232 5230 18244
rect 6270 18232 6276 18244
rect 6328 18272 6334 18284
rect 6733 18275 6791 18281
rect 6328 18244 6408 18272
rect 6328 18232 6334 18244
rect 1946 18164 1952 18216
rect 2004 18204 2010 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 2004 18176 2053 18204
rect 2004 18164 2010 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 2130 18164 2136 18216
rect 2188 18204 2194 18216
rect 2593 18207 2651 18213
rect 2593 18204 2605 18207
rect 2188 18176 2605 18204
rect 2188 18164 2194 18176
rect 2593 18173 2605 18176
rect 2639 18204 2651 18207
rect 3513 18207 3571 18213
rect 2639 18176 2774 18204
rect 2639 18173 2651 18176
rect 2593 18167 2651 18173
rect 1762 18096 1768 18148
rect 1820 18096 1826 18148
rect 2406 18096 2412 18148
rect 2464 18096 2470 18148
rect 2038 18028 2044 18080
rect 2096 18068 2102 18080
rect 2424 18068 2452 18096
rect 2096 18040 2452 18068
rect 2746 18068 2774 18176
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3970 18204 3976 18216
rect 3559 18176 3976 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 4764 18176 5641 18204
rect 4764 18164 4770 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 5997 18207 6055 18213
rect 5997 18173 6009 18207
rect 6043 18173 6055 18207
rect 5997 18167 6055 18173
rect 3786 18096 3792 18148
rect 3844 18136 3850 18148
rect 5258 18136 5264 18148
rect 3844 18108 5264 18136
rect 3844 18096 3850 18108
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 6012 18136 6040 18167
rect 6178 18164 6184 18216
rect 6236 18164 6242 18216
rect 6380 18213 6408 18244
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 12066 18272 12072 18284
rect 6779 18244 12072 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 12406 18272 12434 18312
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 14366 18340 14372 18352
rect 12676 18312 14372 18340
rect 12676 18300 12682 18312
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 18138 18340 18144 18352
rect 16040 18312 18144 18340
rect 12406 18244 13952 18272
rect 6365 18207 6423 18213
rect 6365 18173 6377 18207
rect 6411 18173 6423 18207
rect 6365 18167 6423 18173
rect 6638 18164 6644 18216
rect 6696 18164 6702 18216
rect 8478 18204 8484 18216
rect 6840 18176 8484 18204
rect 6840 18136 6868 18176
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 8665 18207 8723 18213
rect 8665 18173 8677 18207
rect 8711 18204 8723 18207
rect 8846 18204 8852 18216
rect 8711 18176 8852 18204
rect 8711 18173 8723 18176
rect 8665 18167 8723 18173
rect 8846 18164 8852 18176
rect 8904 18204 8910 18216
rect 9769 18207 9827 18213
rect 8904 18176 9168 18204
rect 8904 18164 8910 18176
rect 6012 18108 6868 18136
rect 6917 18139 6975 18145
rect 6917 18105 6929 18139
rect 6963 18105 6975 18139
rect 6917 18099 6975 18105
rect 3329 18071 3387 18077
rect 3329 18068 3341 18071
rect 2746 18040 3341 18068
rect 2096 18028 2102 18040
rect 3329 18037 3341 18040
rect 3375 18037 3387 18071
rect 3329 18031 3387 18037
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 5350 18068 5356 18080
rect 4304 18040 5356 18068
rect 4304 18028 4310 18040
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6932 18068 6960 18099
rect 7006 18096 7012 18148
rect 7064 18136 7070 18148
rect 7282 18136 7288 18148
rect 7064 18108 7288 18136
rect 7064 18096 7070 18108
rect 7282 18096 7288 18108
rect 7340 18096 7346 18148
rect 7374 18096 7380 18148
rect 7432 18096 7438 18148
rect 7558 18096 7564 18148
rect 7616 18136 7622 18148
rect 8294 18136 8300 18148
rect 7616 18108 8300 18136
rect 7616 18096 7622 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 9140 18136 9168 18176
rect 9769 18173 9781 18207
rect 9815 18204 9827 18207
rect 10134 18204 10140 18216
rect 9815 18176 10140 18204
rect 9815 18173 9827 18176
rect 9769 18167 9827 18173
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18204 10287 18207
rect 10318 18204 10324 18216
rect 10275 18176 10324 18204
rect 10275 18173 10287 18176
rect 10229 18167 10287 18173
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 11517 18207 11575 18213
rect 11517 18173 11529 18207
rect 11563 18204 11575 18207
rect 11790 18204 11796 18216
rect 11563 18176 11796 18204
rect 11563 18173 11575 18176
rect 11517 18167 11575 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 13265 18207 13323 18213
rect 11931 18176 13225 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 10502 18136 10508 18148
rect 9140 18108 10508 18136
rect 10502 18096 10508 18108
rect 10560 18096 10566 18148
rect 10594 18096 10600 18148
rect 10652 18096 10658 18148
rect 11054 18096 11060 18148
rect 11112 18096 11118 18148
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 11609 18139 11667 18145
rect 11609 18136 11621 18139
rect 11204 18108 11621 18136
rect 11204 18096 11210 18108
rect 11609 18105 11621 18108
rect 11655 18105 11667 18139
rect 12618 18136 12624 18148
rect 11609 18099 11667 18105
rect 11716 18108 12624 18136
rect 6328 18040 6960 18068
rect 6328 18028 6334 18040
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 8386 18068 8392 18080
rect 7156 18040 8392 18068
rect 7156 18028 7162 18040
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 9953 18071 10011 18077
rect 9953 18068 9965 18071
rect 9272 18040 9965 18068
rect 9272 18028 9278 18040
rect 9953 18037 9965 18040
rect 9999 18068 10011 18071
rect 10612 18068 10640 18096
rect 9999 18040 10640 18068
rect 9999 18037 10011 18040
rect 9953 18031 10011 18037
rect 11238 18028 11244 18080
rect 11296 18077 11302 18080
rect 11716 18077 11744 18108
rect 12618 18096 12624 18108
rect 12676 18096 12682 18148
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 13081 18139 13139 18145
rect 13081 18136 13093 18139
rect 12860 18108 13093 18136
rect 12860 18096 12866 18108
rect 13081 18105 13093 18108
rect 13127 18105 13139 18139
rect 13197 18136 13225 18176
rect 13265 18173 13277 18207
rect 13311 18204 13323 18207
rect 13630 18204 13636 18216
rect 13311 18176 13636 18204
rect 13311 18173 13323 18176
rect 13265 18167 13323 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 13725 18207 13783 18213
rect 13725 18173 13737 18207
rect 13771 18204 13783 18207
rect 13814 18204 13820 18216
rect 13771 18176 13820 18204
rect 13771 18173 13783 18176
rect 13725 18167 13783 18173
rect 13740 18136 13768 18167
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 13924 18213 13952 18244
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14148 18244 14289 18272
rect 14148 18232 14154 18244
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 14642 18232 14648 18284
rect 14700 18232 14706 18284
rect 14918 18232 14924 18284
rect 14976 18232 14982 18284
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 13998 18164 14004 18216
rect 14056 18164 14062 18216
rect 14185 18207 14243 18213
rect 14185 18173 14197 18207
rect 14231 18204 14243 18207
rect 14366 18204 14372 18216
rect 14231 18176 14372 18204
rect 14231 18173 14243 18176
rect 14185 18167 14243 18173
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 16040 18190 16068 18312
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 18690 18300 18696 18352
rect 18748 18340 18754 18352
rect 18877 18343 18935 18349
rect 18877 18340 18889 18343
rect 18748 18312 18889 18340
rect 18748 18300 18754 18312
rect 18877 18309 18889 18312
rect 18923 18309 18935 18343
rect 19306 18340 19334 18380
rect 19429 18377 19441 18411
rect 19475 18408 19487 18411
rect 19610 18408 19616 18420
rect 19475 18380 19616 18408
rect 19475 18377 19487 18380
rect 19429 18371 19487 18377
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 22370 18408 22376 18420
rect 20916 18380 22376 18408
rect 19521 18343 19579 18349
rect 19521 18340 19533 18343
rect 19306 18312 19533 18340
rect 18877 18303 18935 18309
rect 19521 18309 19533 18312
rect 19567 18340 19579 18343
rect 20254 18340 20260 18352
rect 19567 18312 20260 18340
rect 19567 18309 19579 18312
rect 19521 18303 19579 18309
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 20438 18300 20444 18352
rect 20496 18340 20502 18352
rect 20622 18340 20628 18352
rect 20496 18312 20628 18340
rect 20496 18300 20502 18312
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16356 18244 17540 18272
rect 16356 18232 16362 18244
rect 16390 18164 16396 18216
rect 16448 18204 16454 18216
rect 16448 18176 16804 18204
rect 16448 18164 16454 18176
rect 16669 18139 16727 18145
rect 16669 18136 16681 18139
rect 13197 18108 13768 18136
rect 16224 18108 16681 18136
rect 13081 18099 13139 18105
rect 11296 18071 11315 18077
rect 11303 18037 11315 18071
rect 11296 18031 11315 18037
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18037 11759 18071
rect 11701 18031 11759 18037
rect 11885 18071 11943 18077
rect 11885 18037 11897 18071
rect 11931 18068 11943 18071
rect 12250 18068 12256 18080
rect 11931 18040 12256 18068
rect 11931 18037 11943 18040
rect 11885 18031 11943 18037
rect 11296 18028 11302 18031
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 13633 18071 13691 18077
rect 13633 18068 13645 18071
rect 13504 18040 13645 18068
rect 13504 18028 13510 18040
rect 13633 18037 13645 18040
rect 13679 18037 13691 18071
rect 13633 18031 13691 18037
rect 14274 18028 14280 18080
rect 14332 18028 14338 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 16224 18068 16252 18108
rect 16669 18105 16681 18108
rect 16715 18105 16727 18139
rect 16776 18136 16804 18176
rect 17218 18164 17224 18216
rect 17276 18164 17282 18216
rect 17512 18213 17540 18244
rect 19076 18244 20760 18272
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18204 17555 18207
rect 18966 18204 18972 18216
rect 17543 18176 18972 18204
rect 17543 18173 17555 18176
rect 17497 18167 17555 18173
rect 18966 18164 18972 18176
rect 19024 18164 19030 18216
rect 19076 18213 19104 18244
rect 19061 18207 19119 18213
rect 19061 18173 19073 18207
rect 19107 18173 19119 18207
rect 19061 18167 19119 18173
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 19208 18176 19257 18204
rect 19208 18164 19214 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 19978 18204 19984 18216
rect 19751 18176 19984 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 19978 18164 19984 18176
rect 20036 18204 20042 18216
rect 20349 18207 20407 18213
rect 20349 18204 20361 18207
rect 20036 18176 20361 18204
rect 20036 18164 20042 18176
rect 20349 18173 20361 18176
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 20530 18164 20536 18216
rect 20588 18164 20594 18216
rect 20732 18213 20760 18244
rect 20717 18207 20775 18213
rect 20717 18173 20729 18207
rect 20763 18204 20775 18207
rect 20806 18204 20812 18216
rect 20763 18176 20812 18204
rect 20763 18173 20775 18176
rect 20717 18167 20775 18173
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 20916 18213 20944 18380
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 23198 18368 23204 18420
rect 23256 18408 23262 18420
rect 23293 18411 23351 18417
rect 23293 18408 23305 18411
rect 23256 18380 23305 18408
rect 23256 18368 23262 18380
rect 23293 18377 23305 18380
rect 23339 18377 23351 18411
rect 23293 18371 23351 18377
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 27985 18411 28043 18417
rect 27985 18408 27997 18411
rect 23440 18380 27997 18408
rect 23440 18368 23446 18380
rect 27985 18377 27997 18380
rect 28031 18408 28043 18411
rect 28442 18408 28448 18420
rect 28031 18380 28448 18408
rect 28031 18377 28043 18380
rect 27985 18371 28043 18377
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 29086 18408 29092 18420
rect 28552 18380 29092 18408
rect 21174 18300 21180 18352
rect 21232 18340 21238 18352
rect 21542 18340 21548 18352
rect 21232 18312 21548 18340
rect 21232 18300 21238 18312
rect 21542 18300 21548 18312
rect 21600 18300 21606 18352
rect 22738 18340 22744 18352
rect 22572 18312 22744 18340
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 21818 18272 21824 18284
rect 21140 18244 21824 18272
rect 21140 18232 21146 18244
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22572 18213 22600 18312
rect 22738 18300 22744 18312
rect 22796 18340 22802 18352
rect 23109 18343 23167 18349
rect 23109 18340 23121 18343
rect 22796 18312 23121 18340
rect 22796 18300 22802 18312
rect 23109 18309 23121 18312
rect 23155 18309 23167 18343
rect 23109 18303 23167 18309
rect 23566 18300 23572 18352
rect 23624 18340 23630 18352
rect 24305 18343 24363 18349
rect 24305 18340 24317 18343
rect 23624 18312 24317 18340
rect 23624 18300 23630 18312
rect 24305 18309 24317 18312
rect 24351 18309 24363 18343
rect 24305 18303 24363 18309
rect 24486 18300 24492 18352
rect 24544 18300 24550 18352
rect 28258 18300 28264 18352
rect 28316 18340 28322 18352
rect 28552 18340 28580 18380
rect 29086 18368 29092 18380
rect 29144 18368 29150 18420
rect 29270 18368 29276 18420
rect 29328 18408 29334 18420
rect 29454 18408 29460 18420
rect 29328 18380 29460 18408
rect 29328 18368 29334 18380
rect 29454 18368 29460 18380
rect 29512 18368 29518 18420
rect 29730 18368 29736 18420
rect 29788 18408 29794 18420
rect 30837 18411 30895 18417
rect 30837 18408 30849 18411
rect 29788 18380 30849 18408
rect 29788 18368 29794 18380
rect 30837 18377 30849 18380
rect 30883 18377 30895 18411
rect 30837 18371 30895 18377
rect 30926 18368 30932 18420
rect 30984 18408 30990 18420
rect 31021 18411 31079 18417
rect 31021 18408 31033 18411
rect 30984 18380 31033 18408
rect 30984 18368 30990 18380
rect 31021 18377 31033 18380
rect 31067 18377 31079 18411
rect 31021 18371 31079 18377
rect 28316 18312 28580 18340
rect 28316 18300 28322 18312
rect 28902 18300 28908 18352
rect 28960 18340 28966 18352
rect 28960 18312 29132 18340
rect 28960 18300 28966 18312
rect 23017 18275 23075 18281
rect 23017 18241 23029 18275
rect 23063 18272 23075 18275
rect 24213 18275 24271 18281
rect 23063 18244 24072 18272
rect 23063 18241 23075 18244
rect 23017 18235 23075 18241
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 21177 18207 21235 18213
rect 21177 18173 21189 18207
rect 21223 18204 21235 18207
rect 22557 18207 22615 18213
rect 21223 18176 22508 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 17405 18139 17463 18145
rect 17405 18136 17417 18139
rect 16776 18108 17417 18136
rect 16669 18099 16727 18105
rect 17405 18105 17417 18108
rect 17451 18136 17463 18139
rect 17586 18136 17592 18148
rect 17451 18108 17592 18136
rect 17451 18105 17463 18108
rect 17405 18099 17463 18105
rect 17586 18096 17592 18108
rect 17644 18096 17650 18148
rect 18984 18136 19012 18164
rect 19518 18136 19524 18148
rect 18984 18108 19524 18136
rect 19518 18096 19524 18108
rect 19576 18096 19582 18148
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20119 18108 20208 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 15896 18040 16252 18068
rect 15896 18028 15902 18040
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 17770 18068 17776 18080
rect 16356 18040 17776 18068
rect 16356 18028 16362 18040
rect 17770 18028 17776 18040
rect 17828 18068 17834 18080
rect 19153 18071 19211 18077
rect 19153 18068 19165 18071
rect 17828 18040 19165 18068
rect 17828 18028 17834 18040
rect 19153 18037 19165 18040
rect 19199 18068 19211 18071
rect 19610 18068 19616 18080
rect 19199 18040 19616 18068
rect 19199 18037 19211 18040
rect 19153 18031 19211 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 19794 18028 19800 18080
rect 19852 18028 19858 18080
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18068 19947 18071
rect 19978 18068 19984 18080
rect 19935 18040 19984 18068
rect 19935 18037 19947 18040
rect 19889 18031 19947 18037
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20180 18077 20208 18108
rect 20438 18096 20444 18148
rect 20496 18096 20502 18148
rect 21192 18136 21220 18167
rect 20548 18108 21220 18136
rect 21821 18139 21879 18145
rect 20165 18071 20223 18077
rect 20165 18037 20177 18071
rect 20211 18068 20223 18071
rect 20548 18068 20576 18108
rect 21821 18105 21833 18139
rect 21867 18105 21879 18139
rect 21821 18099 21879 18105
rect 20211 18040 20576 18068
rect 20211 18037 20223 18040
rect 20165 18031 20223 18037
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20990 18068 20996 18080
rect 20772 18040 20996 18068
rect 20772 18028 20778 18040
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21358 18028 21364 18080
rect 21416 18028 21422 18080
rect 21542 18028 21548 18080
rect 21600 18028 21606 18080
rect 21836 18068 21864 18099
rect 21910 18096 21916 18148
rect 21968 18136 21974 18148
rect 22373 18139 22431 18145
rect 22373 18136 22385 18139
rect 21968 18108 22385 18136
rect 21968 18096 21974 18108
rect 22373 18105 22385 18108
rect 22419 18105 22431 18139
rect 22480 18136 22508 18176
rect 22557 18173 22569 18207
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 22833 18207 22891 18213
rect 22833 18173 22845 18207
rect 22879 18204 22891 18207
rect 23290 18204 23296 18216
rect 22879 18176 23296 18204
rect 22879 18173 22891 18176
rect 22833 18167 22891 18173
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 23842 18204 23848 18216
rect 23400 18176 23848 18204
rect 23400 18136 23428 18176
rect 23842 18164 23848 18176
rect 23900 18164 23906 18216
rect 23934 18164 23940 18216
rect 23992 18164 23998 18216
rect 24044 18213 24072 18244
rect 24213 18241 24225 18275
rect 24259 18272 24271 18275
rect 24504 18272 24532 18300
rect 24259 18244 24532 18272
rect 24259 18241 24271 18244
rect 24213 18235 24271 18241
rect 24670 18232 24676 18284
rect 24728 18232 24734 18284
rect 27065 18275 27123 18281
rect 27065 18272 27077 18275
rect 24872 18244 27077 18272
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18173 24087 18207
rect 24029 18167 24087 18173
rect 24394 18164 24400 18216
rect 24452 18204 24458 18216
rect 24489 18207 24547 18213
rect 24489 18204 24501 18207
rect 24452 18176 24501 18204
rect 24452 18164 24458 18176
rect 24489 18173 24501 18176
rect 24535 18204 24547 18207
rect 24578 18204 24584 18216
rect 24535 18176 24584 18204
rect 24535 18173 24547 18176
rect 24489 18167 24547 18173
rect 24578 18164 24584 18176
rect 24636 18164 24642 18216
rect 22480 18108 23428 18136
rect 22373 18099 22431 18105
rect 23474 18096 23480 18148
rect 23532 18096 23538 18148
rect 24118 18096 24124 18148
rect 24176 18136 24182 18148
rect 24872 18145 24900 18244
rect 27065 18241 27077 18244
rect 27111 18272 27123 18275
rect 27522 18272 27528 18284
rect 27111 18244 27528 18272
rect 27111 18241 27123 18244
rect 27065 18235 27123 18241
rect 27522 18232 27528 18244
rect 27580 18232 27586 18284
rect 28718 18272 28724 18284
rect 27632 18244 28724 18272
rect 27632 18213 27660 18244
rect 28718 18232 28724 18244
rect 28776 18232 28782 18284
rect 28994 18232 29000 18284
rect 29052 18232 29058 18284
rect 29104 18272 29132 18312
rect 30742 18300 30748 18352
rect 30800 18300 30806 18352
rect 30006 18272 30012 18284
rect 29104 18244 30012 18272
rect 30006 18232 30012 18244
rect 30064 18272 30070 18284
rect 31110 18272 31116 18284
rect 30064 18244 31116 18272
rect 30064 18232 30070 18244
rect 31110 18232 31116 18244
rect 31168 18232 31174 18284
rect 27617 18207 27675 18213
rect 27617 18173 27629 18207
rect 27663 18173 27675 18207
rect 27617 18167 27675 18173
rect 27706 18164 27712 18216
rect 27764 18164 27770 18216
rect 27890 18213 27896 18216
rect 27847 18207 27896 18213
rect 27847 18173 27859 18207
rect 27893 18173 27896 18207
rect 27847 18167 27896 18173
rect 27890 18164 27896 18167
rect 27948 18164 27954 18216
rect 28169 18207 28227 18213
rect 28169 18173 28181 18207
rect 28215 18204 28227 18207
rect 28258 18204 28264 18216
rect 28215 18176 28264 18204
rect 28215 18173 28227 18176
rect 28169 18167 28227 18173
rect 28258 18164 28264 18176
rect 28316 18164 28322 18216
rect 28442 18164 28448 18216
rect 28500 18164 28506 18216
rect 28626 18164 28632 18216
rect 28684 18164 28690 18216
rect 24857 18139 24915 18145
rect 24857 18136 24869 18139
rect 24176 18108 24869 18136
rect 24176 18096 24182 18108
rect 24857 18105 24869 18108
rect 24903 18105 24915 18139
rect 24857 18099 24915 18105
rect 25130 18096 25136 18148
rect 25188 18136 25194 18148
rect 25188 18108 25452 18136
rect 25188 18096 25194 18108
rect 22094 18068 22100 18080
rect 21836 18040 22100 18068
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 22649 18071 22707 18077
rect 22649 18037 22661 18071
rect 22695 18068 22707 18071
rect 22830 18068 22836 18080
rect 22695 18040 22836 18068
rect 22695 18037 22707 18040
rect 22649 18031 22707 18037
rect 22830 18028 22836 18040
rect 22888 18028 22894 18080
rect 23277 18071 23335 18077
rect 23277 18037 23289 18071
rect 23323 18068 23335 18071
rect 24946 18068 24952 18080
rect 23323 18040 24952 18068
rect 23323 18037 23335 18040
rect 23277 18031 23335 18037
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 25317 18071 25375 18077
rect 25317 18068 25329 18071
rect 25280 18040 25329 18068
rect 25280 18028 25286 18040
rect 25317 18037 25329 18040
rect 25363 18037 25375 18071
rect 25424 18068 25452 18108
rect 26326 18096 26332 18148
rect 26384 18096 26390 18148
rect 26510 18096 26516 18148
rect 26568 18136 26574 18148
rect 26789 18139 26847 18145
rect 26789 18136 26801 18139
rect 26568 18108 26801 18136
rect 26568 18096 26574 18108
rect 26789 18105 26801 18108
rect 26835 18105 26847 18139
rect 26789 18099 26847 18105
rect 26878 18096 26884 18148
rect 26936 18136 26942 18148
rect 27341 18139 27399 18145
rect 27341 18136 27353 18139
rect 26936 18108 27353 18136
rect 26936 18096 26942 18108
rect 27341 18105 27353 18108
rect 27387 18105 27399 18139
rect 27341 18099 27399 18105
rect 28077 18139 28135 18145
rect 28077 18105 28089 18139
rect 28123 18136 28135 18139
rect 29178 18136 29184 18148
rect 28123 18108 29184 18136
rect 28123 18105 28135 18108
rect 28077 18099 28135 18105
rect 29178 18096 29184 18108
rect 29236 18096 29242 18148
rect 29270 18096 29276 18148
rect 29328 18096 29334 18148
rect 29730 18096 29736 18148
rect 29788 18096 29794 18148
rect 31202 18096 31208 18148
rect 31260 18096 31266 18148
rect 25866 18068 25872 18080
rect 25424 18040 25872 18068
rect 25317 18031 25375 18037
rect 25866 18028 25872 18040
rect 25924 18068 25930 18080
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 25924 18040 28365 18068
rect 25924 18028 25930 18040
rect 28353 18037 28365 18040
rect 28399 18037 28411 18071
rect 28353 18031 28411 18037
rect 28534 18028 28540 18080
rect 28592 18068 28598 18080
rect 30190 18068 30196 18080
rect 28592 18040 30196 18068
rect 28592 18028 28598 18040
rect 30190 18028 30196 18040
rect 30248 18028 30254 18080
rect 31005 18071 31063 18077
rect 31005 18037 31017 18071
rect 31051 18068 31063 18071
rect 31386 18068 31392 18080
rect 31051 18040 31392 18068
rect 31051 18037 31063 18040
rect 31005 18031 31063 18037
rect 31386 18028 31392 18040
rect 31444 18028 31450 18080
rect 552 17978 31648 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 12096 17978
rect 12148 17926 12160 17978
rect 12212 17926 12224 17978
rect 12276 17926 12288 17978
rect 12340 17926 12352 17978
rect 12404 17926 19870 17978
rect 19922 17926 19934 17978
rect 19986 17926 19998 17978
rect 20050 17926 20062 17978
rect 20114 17926 20126 17978
rect 20178 17926 27644 17978
rect 27696 17926 27708 17978
rect 27760 17926 27772 17978
rect 27824 17926 27836 17978
rect 27888 17926 27900 17978
rect 27952 17926 31648 17978
rect 552 17904 31648 17926
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 4341 17867 4399 17873
rect 3016 17836 4292 17864
rect 3016 17824 3022 17836
rect 2222 17756 2228 17808
rect 2280 17756 2286 17808
rect 3786 17796 3792 17808
rect 2608 17768 3792 17796
rect 2608 17740 2636 17768
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 4062 17796 4068 17808
rect 3896 17768 4068 17796
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17728 1547 17731
rect 1762 17728 1768 17740
rect 1535 17700 1768 17728
rect 1535 17697 1547 17700
rect 1489 17691 1547 17697
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 1854 17688 1860 17740
rect 1912 17728 1918 17740
rect 2409 17731 2467 17737
rect 2409 17728 2421 17731
rect 1912 17700 2421 17728
rect 1912 17688 1918 17700
rect 2409 17697 2421 17700
rect 2455 17697 2467 17731
rect 2409 17691 2467 17697
rect 2590 17688 2596 17740
rect 2648 17688 2654 17740
rect 3896 17737 3924 17768
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 4264 17796 4292 17836
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 4706 17864 4712 17876
rect 4387 17836 4712 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 5626 17824 5632 17876
rect 5684 17864 5690 17876
rect 5905 17867 5963 17873
rect 5905 17864 5917 17867
rect 5684 17836 5917 17864
rect 5684 17824 5690 17836
rect 5905 17833 5917 17836
rect 5951 17864 5963 17867
rect 6638 17864 6644 17876
rect 5951 17836 6644 17864
rect 5951 17833 5963 17836
rect 5905 17827 5963 17833
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 7466 17864 7472 17876
rect 7423 17836 7472 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 7837 17867 7895 17873
rect 7837 17833 7849 17867
rect 7883 17864 7895 17867
rect 8202 17864 8208 17876
rect 7883 17836 8208 17864
rect 7883 17833 7895 17836
rect 7837 17827 7895 17833
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 8941 17867 8999 17873
rect 8588 17836 8800 17864
rect 8110 17796 8116 17808
rect 4264 17768 8116 17796
rect 8110 17756 8116 17768
rect 8168 17756 8174 17808
rect 8588 17805 8616 17836
rect 8573 17799 8631 17805
rect 8573 17765 8585 17799
rect 8619 17765 8631 17799
rect 8772 17796 8800 17836
rect 8941 17833 8953 17867
rect 8987 17864 8999 17867
rect 9214 17864 9220 17876
rect 8987 17836 9220 17864
rect 8987 17833 8999 17836
rect 8941 17827 8999 17833
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 9953 17867 10011 17873
rect 9953 17864 9965 17867
rect 9324 17836 9965 17864
rect 9122 17796 9128 17808
rect 8772 17768 9128 17796
rect 8573 17759 8631 17765
rect 9122 17756 9128 17768
rect 9180 17756 9186 17808
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17697 2743 17731
rect 2685 17691 2743 17697
rect 2794 17731 2852 17737
rect 2794 17697 2806 17731
rect 2840 17728 2852 17731
rect 3605 17731 3663 17737
rect 2840 17700 2912 17728
rect 2840 17697 2852 17700
rect 2794 17691 2852 17697
rect 1302 17620 1308 17672
rect 1360 17620 1366 17672
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2700 17660 2728 17691
rect 2280 17632 2728 17660
rect 2884 17660 2912 17700
rect 3605 17697 3617 17731
rect 3651 17697 3663 17731
rect 3605 17691 3663 17697
rect 3881 17731 3939 17737
rect 3881 17697 3893 17731
rect 3927 17697 3939 17731
rect 3881 17691 3939 17697
rect 3329 17663 3387 17669
rect 3329 17660 3341 17663
rect 2884 17632 3341 17660
rect 2280 17620 2286 17632
rect 1320 17592 1348 17620
rect 2884 17592 2912 17632
rect 3329 17629 3341 17632
rect 3375 17629 3387 17663
rect 3329 17623 3387 17629
rect 1320 17564 2912 17592
rect 2958 17552 2964 17604
rect 3016 17592 3022 17604
rect 3053 17595 3111 17601
rect 3053 17592 3065 17595
rect 3016 17564 3065 17592
rect 3016 17552 3022 17564
rect 3053 17561 3065 17564
rect 3099 17561 3111 17595
rect 3053 17555 3111 17561
rect 1670 17484 1676 17536
rect 1728 17484 1734 17536
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17524 2191 17527
rect 2222 17524 2228 17536
rect 2179 17496 2228 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 3620 17524 3648 17691
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 4028 17700 4752 17728
rect 4028 17688 4034 17700
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4157 17663 4215 17669
rect 4157 17660 4169 17663
rect 4120 17632 4169 17660
rect 4120 17620 4126 17632
rect 4157 17629 4169 17632
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4246 17620 4252 17672
rect 4304 17620 4310 17672
rect 3973 17595 4031 17601
rect 3973 17561 3985 17595
rect 4019 17592 4031 17595
rect 4433 17595 4491 17601
rect 4433 17592 4445 17595
rect 4019 17564 4445 17592
rect 4019 17561 4031 17564
rect 3973 17555 4031 17561
rect 4433 17561 4445 17564
rect 4479 17561 4491 17595
rect 4724 17592 4752 17700
rect 4798 17688 4804 17740
rect 4856 17688 4862 17740
rect 4908 17700 5764 17728
rect 4908 17669 4936 17700
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 4985 17663 5043 17669
rect 4985 17629 4997 17663
rect 5031 17629 5043 17663
rect 5736 17660 5764 17700
rect 5810 17688 5816 17740
rect 5868 17688 5874 17740
rect 5994 17688 6000 17740
rect 6052 17728 6058 17740
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 6052 17700 6101 17728
rect 6052 17688 6058 17700
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 6733 17731 6791 17737
rect 6733 17697 6745 17731
rect 6779 17728 6791 17731
rect 6822 17728 6828 17740
rect 6779 17700 6828 17728
rect 6779 17697 6791 17700
rect 6733 17691 6791 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7098 17688 7104 17740
rect 7156 17688 7162 17740
rect 7193 17731 7251 17737
rect 7193 17697 7205 17731
rect 7239 17728 7251 17731
rect 7374 17728 7380 17740
rect 7239 17700 7380 17728
rect 7239 17697 7251 17700
rect 7193 17691 7251 17697
rect 6546 17660 6552 17672
rect 5736 17632 6552 17660
rect 4985 17623 5043 17629
rect 5000 17592 5028 17623
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 6914 17620 6920 17672
rect 6972 17620 6978 17672
rect 7006 17620 7012 17672
rect 7064 17620 7070 17672
rect 7208 17592 7236 17691
rect 7374 17688 7380 17700
rect 7432 17728 7438 17740
rect 7834 17728 7840 17740
rect 7432 17700 7840 17728
rect 7432 17688 7438 17700
rect 7834 17688 7840 17700
rect 7892 17688 7898 17740
rect 8297 17731 8355 17737
rect 8297 17697 8309 17731
rect 8343 17697 8355 17731
rect 8297 17691 8355 17697
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 8018 17620 8024 17672
rect 8076 17620 8082 17672
rect 7926 17592 7932 17604
rect 4724 17564 7236 17592
rect 7300 17564 7932 17592
rect 4433 17555 4491 17561
rect 5902 17524 5908 17536
rect 3620 17496 5908 17524
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6270 17524 6276 17536
rect 6052 17496 6276 17524
rect 6052 17484 6058 17496
rect 6270 17484 6276 17496
rect 6328 17484 6334 17536
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 7300 17524 7328 17564
rect 7926 17552 7932 17564
rect 7984 17552 7990 17604
rect 8319 17592 8347 17691
rect 8386 17688 8392 17740
rect 8444 17737 8450 17740
rect 8846 17737 8852 17740
rect 8444 17731 8475 17737
rect 8463 17697 8475 17731
rect 8444 17691 8475 17697
rect 8665 17731 8723 17737
rect 8665 17697 8677 17731
rect 8711 17697 8723 17731
rect 8665 17691 8723 17697
rect 8803 17731 8852 17737
rect 8803 17697 8815 17731
rect 8849 17697 8852 17731
rect 8803 17691 8852 17697
rect 8444 17688 8450 17691
rect 8680 17660 8708 17691
rect 8846 17688 8852 17691
rect 8904 17688 8910 17740
rect 9033 17731 9091 17737
rect 9033 17697 9045 17731
rect 9079 17728 9091 17731
rect 9140 17728 9168 17756
rect 9079 17700 9168 17728
rect 9217 17731 9275 17737
rect 9079 17697 9091 17700
rect 9033 17691 9091 17697
rect 9217 17697 9229 17731
rect 9263 17728 9275 17731
rect 9324 17728 9352 17836
rect 9953 17833 9965 17836
rect 9999 17833 10011 17867
rect 9953 17827 10011 17833
rect 10226 17824 10232 17876
rect 10284 17864 10290 17876
rect 10410 17864 10416 17876
rect 10284 17836 10416 17864
rect 10284 17824 10290 17836
rect 10410 17824 10416 17836
rect 10468 17824 10474 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 17405 17867 17463 17873
rect 10652 17836 16712 17864
rect 10652 17824 10658 17836
rect 9398 17756 9404 17808
rect 9456 17796 9462 17808
rect 9858 17796 9864 17808
rect 9456 17768 9864 17796
rect 9456 17756 9462 17768
rect 9858 17756 9864 17768
rect 9916 17796 9922 17808
rect 16390 17796 16396 17808
rect 9916 17768 10364 17796
rect 9916 17756 9922 17768
rect 9263 17700 9352 17728
rect 9263 17697 9275 17700
rect 9217 17691 9275 17697
rect 9582 17688 9588 17740
rect 9640 17688 9646 17740
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17728 9827 17731
rect 10134 17728 10140 17740
rect 9815 17700 10140 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 10336 17737 10364 17768
rect 10704 17768 16396 17796
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17697 10379 17731
rect 10321 17691 10379 17697
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 10704 17737 10732 17768
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 10468 17700 10517 17728
rect 10468 17688 10474 17700
rect 10505 17697 10517 17700
rect 10551 17697 10563 17731
rect 10505 17691 10563 17697
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11296 17700 11621 17728
rect 11296 17688 11302 17700
rect 11609 17697 11621 17700
rect 11655 17728 11667 17731
rect 11790 17728 11796 17740
rect 11655 17700 11796 17728
rect 11655 17697 11667 17700
rect 11609 17691 11667 17697
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 11900 17737 11928 17768
rect 16390 17756 16396 17768
rect 16448 17756 16454 17808
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17697 11943 17731
rect 11885 17691 11943 17697
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 12802 17688 12808 17740
rect 12860 17688 12866 17740
rect 12989 17731 13047 17737
rect 12989 17697 13001 17731
rect 13035 17728 13047 17731
rect 13078 17728 13084 17740
rect 13035 17700 13084 17728
rect 13035 17697 13047 17700
rect 12989 17691 13047 17697
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 13265 17731 13323 17737
rect 13265 17697 13277 17731
rect 13311 17728 13323 17731
rect 13722 17728 13728 17740
rect 13311 17700 13728 17728
rect 13311 17697 13323 17700
rect 13265 17691 13323 17697
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 14182 17688 14188 17740
rect 14240 17688 14246 17740
rect 14274 17688 14280 17740
rect 14332 17688 14338 17740
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17728 14519 17731
rect 14642 17728 14648 17740
rect 14507 17700 14648 17728
rect 14507 17697 14519 17700
rect 14461 17691 14519 17697
rect 14642 17688 14648 17700
rect 14700 17728 14706 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 14700 17700 15669 17728
rect 14700 17688 14706 17700
rect 15657 17697 15669 17700
rect 15703 17728 15715 17731
rect 16574 17728 16580 17740
rect 15703 17700 16580 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 8938 17660 8944 17672
rect 8680 17632 8944 17660
rect 8938 17620 8944 17632
rect 8996 17620 9002 17672
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 9171 17632 9505 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 9493 17629 9505 17632
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17660 9735 17663
rect 10226 17660 10232 17672
rect 9723 17632 10232 17660
rect 9723 17629 9735 17632
rect 9677 17623 9735 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 11747 17632 12572 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 9214 17592 9220 17604
rect 8319 17564 9220 17592
rect 9214 17552 9220 17564
rect 9272 17552 9278 17604
rect 9306 17552 9312 17604
rect 9364 17552 9370 17604
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 12434 17592 12440 17604
rect 10192 17564 12440 17592
rect 10192 17552 10198 17564
rect 12434 17552 12440 17564
rect 12492 17552 12498 17604
rect 12544 17536 12572 17632
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 12897 17663 12955 17669
rect 12897 17660 12909 17663
rect 12676 17632 12909 17660
rect 12676 17620 12682 17632
rect 12897 17629 12909 17632
rect 12943 17629 12955 17663
rect 12897 17623 12955 17629
rect 12912 17592 12940 17623
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 14056 17632 15301 17660
rect 14056 17620 14062 17632
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 15838 17660 15844 17672
rect 15795 17632 15844 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16684 17660 16712 17836
rect 17405 17833 17417 17867
rect 17451 17864 17463 17867
rect 17678 17864 17684 17876
rect 17451 17836 17684 17864
rect 17451 17833 17463 17836
rect 17405 17827 17463 17833
rect 17678 17824 17684 17836
rect 17736 17824 17742 17876
rect 17788 17836 18828 17864
rect 17034 17756 17040 17808
rect 17092 17756 17098 17808
rect 17218 17756 17224 17808
rect 17276 17805 17282 17808
rect 17276 17799 17295 17805
rect 17283 17765 17295 17799
rect 17276 17759 17295 17765
rect 17276 17756 17282 17759
rect 17678 17688 17684 17740
rect 17736 17688 17742 17740
rect 17788 17737 17816 17836
rect 18800 17805 18828 17836
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 19886 17864 19892 17876
rect 19576 17836 19892 17864
rect 19576 17824 19582 17836
rect 19886 17824 19892 17836
rect 19944 17824 19950 17876
rect 21082 17864 21088 17876
rect 19996 17836 21088 17864
rect 18785 17799 18843 17805
rect 18555 17765 18613 17771
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17697 17831 17731
rect 17773 17691 17831 17697
rect 18046 17688 18052 17740
rect 18104 17688 18110 17740
rect 18322 17688 18328 17740
rect 18380 17688 18386 17740
rect 18555 17731 18567 17765
rect 18601 17740 18613 17765
rect 18785 17765 18797 17799
rect 18831 17765 18843 17799
rect 18785 17759 18843 17765
rect 18601 17731 18604 17740
rect 18555 17725 18604 17731
rect 18584 17688 18604 17725
rect 18656 17688 18662 17740
rect 18800 17728 18828 17759
rect 19610 17756 19616 17808
rect 19668 17796 19674 17808
rect 19996 17796 20024 17836
rect 19668 17768 20024 17796
rect 19668 17756 19674 17768
rect 20070 17728 20076 17740
rect 18800 17700 20076 17728
rect 20070 17688 20076 17700
rect 20128 17688 20134 17740
rect 20272 17737 20300 17836
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21269 17867 21327 17873
rect 21269 17833 21281 17867
rect 21315 17864 21327 17867
rect 21910 17864 21916 17876
rect 21315 17836 21916 17864
rect 21315 17833 21327 17836
rect 21269 17827 21327 17833
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 24026 17864 24032 17876
rect 23308 17836 24032 17864
rect 21450 17796 21456 17808
rect 20456 17768 21456 17796
rect 20456 17740 20484 17768
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 23308 17796 23336 17836
rect 22310 17768 23336 17796
rect 23385 17799 23443 17805
rect 23385 17765 23397 17799
rect 23431 17796 23443 17799
rect 23474 17796 23480 17808
rect 23431 17768 23480 17796
rect 23431 17765 23443 17768
rect 23385 17759 23443 17765
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 23584 17796 23612 17836
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 24210 17824 24216 17876
rect 24268 17864 24274 17876
rect 24394 17864 24400 17876
rect 24268 17836 24400 17864
rect 24268 17824 24274 17836
rect 24394 17824 24400 17836
rect 24452 17824 24458 17876
rect 26237 17867 26295 17873
rect 25470 17836 26096 17864
rect 25470 17805 25498 17836
rect 25225 17799 25283 17805
rect 25225 17796 25237 17799
rect 23584 17768 23874 17796
rect 24688 17768 25237 17796
rect 20165 17731 20223 17737
rect 20165 17697 20177 17731
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 18584 17660 18612 17688
rect 16684 17632 18612 17660
rect 19886 17620 19892 17672
rect 19944 17660 19950 17672
rect 19981 17663 20039 17669
rect 19981 17660 19993 17663
rect 19944 17632 19993 17660
rect 19944 17620 19950 17632
rect 19981 17629 19993 17632
rect 20027 17629 20039 17663
rect 20180 17660 20208 17691
rect 20438 17688 20444 17740
rect 20496 17688 20502 17740
rect 20622 17737 20628 17740
rect 20599 17731 20628 17737
rect 20599 17697 20611 17731
rect 20599 17691 20628 17697
rect 20622 17688 20628 17691
rect 20680 17688 20686 17740
rect 20714 17688 20720 17740
rect 20772 17688 20778 17740
rect 20809 17731 20867 17737
rect 20809 17697 20821 17731
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21174 17728 21180 17740
rect 20947 17700 21180 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 20346 17660 20352 17672
rect 20180 17632 20352 17660
rect 19981 17623 20039 17629
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20824 17660 20852 17691
rect 21174 17688 21180 17700
rect 21232 17688 21238 17740
rect 23017 17731 23075 17737
rect 23017 17697 23029 17731
rect 23063 17728 23075 17731
rect 23109 17731 23167 17737
rect 23109 17728 23121 17731
rect 23063 17700 23121 17728
rect 23063 17697 23075 17700
rect 23017 17691 23075 17697
rect 23109 17697 23121 17700
rect 23155 17697 23167 17731
rect 24688 17728 24716 17768
rect 25225 17765 25237 17768
rect 25271 17765 25283 17799
rect 25225 17759 25283 17765
rect 25455 17799 25513 17805
rect 25455 17765 25467 17799
rect 25501 17765 25513 17799
rect 25455 17759 25513 17765
rect 25866 17756 25872 17808
rect 25924 17756 25930 17808
rect 23109 17691 23167 17697
rect 24596 17700 24716 17728
rect 20732 17632 20852 17660
rect 21085 17663 21143 17669
rect 12912 17564 14044 17592
rect 14016 17536 14044 17564
rect 14182 17552 14188 17604
rect 14240 17592 14246 17604
rect 16206 17592 16212 17604
rect 14240 17564 16212 17592
rect 14240 17552 14246 17564
rect 16206 17552 16212 17564
rect 16264 17592 16270 17604
rect 17589 17595 17647 17601
rect 17589 17592 17601 17595
rect 16264 17564 17601 17592
rect 16264 17552 16270 17564
rect 17589 17561 17601 17564
rect 17635 17561 17647 17595
rect 17589 17555 17647 17561
rect 17678 17552 17684 17604
rect 17736 17592 17742 17604
rect 18046 17592 18052 17604
rect 17736 17564 18052 17592
rect 17736 17552 17742 17564
rect 18046 17552 18052 17564
rect 18104 17552 18110 17604
rect 20254 17592 20260 17604
rect 18156 17564 20260 17592
rect 6512 17496 7328 17524
rect 6512 17484 6518 17496
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7432 17496 8033 17524
rect 7432 17484 7438 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 9398 17524 9404 17536
rect 8168 17496 9404 17524
rect 8168 17484 8174 17496
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10229 17527 10287 17533
rect 10229 17524 10241 17527
rect 9732 17496 10241 17524
rect 9732 17484 9738 17496
rect 10229 17493 10241 17496
rect 10275 17524 10287 17527
rect 10318 17524 10324 17536
rect 10275 17496 10324 17524
rect 10275 17493 10287 17496
rect 10229 17487 10287 17493
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 10413 17527 10471 17533
rect 10413 17493 10425 17527
rect 10459 17524 10471 17527
rect 10594 17524 10600 17536
rect 10459 17496 10600 17524
rect 10459 17493 10471 17496
rect 10413 17487 10471 17493
rect 10594 17484 10600 17496
rect 10652 17484 10658 17536
rect 10686 17484 10692 17536
rect 10744 17524 10750 17536
rect 11885 17527 11943 17533
rect 11885 17524 11897 17527
rect 10744 17496 11897 17524
rect 10744 17484 10750 17496
rect 11885 17493 11897 17496
rect 11931 17524 11943 17527
rect 11974 17524 11980 17536
rect 11931 17496 11980 17524
rect 11931 17493 11943 17496
rect 11885 17487 11943 17493
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12069 17527 12127 17533
rect 12069 17493 12081 17527
rect 12115 17524 12127 17527
rect 12158 17524 12164 17536
rect 12115 17496 12164 17524
rect 12115 17493 12127 17496
rect 12069 17487 12127 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12526 17484 12532 17536
rect 12584 17484 12590 17536
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13633 17527 13691 17533
rect 13633 17524 13645 17527
rect 13136 17496 13645 17524
rect 13136 17484 13142 17496
rect 13633 17493 13645 17496
rect 13679 17524 13691 17527
rect 13722 17524 13728 17536
rect 13679 17496 13728 17524
rect 13679 17493 13691 17496
rect 13633 17487 13691 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 13998 17484 14004 17536
rect 14056 17484 14062 17536
rect 14369 17527 14427 17533
rect 14369 17493 14381 17527
rect 14415 17524 14427 17527
rect 14734 17524 14740 17536
rect 14415 17496 14740 17524
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 16758 17524 16764 17536
rect 15804 17496 16764 17524
rect 15804 17484 15810 17496
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 17221 17527 17279 17533
rect 17221 17493 17233 17527
rect 17267 17524 17279 17527
rect 18156 17524 18184 17564
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 17267 17496 18184 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 18230 17484 18236 17536
rect 18288 17484 18294 17536
rect 18414 17484 18420 17536
rect 18472 17484 18478 17536
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 19702 17524 19708 17536
rect 19024 17496 19708 17524
rect 19024 17484 19030 17496
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19794 17484 19800 17536
rect 19852 17524 19858 17536
rect 20732 17524 20760 17632
rect 21085 17629 21097 17663
rect 21131 17660 21143 17663
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 21131 17632 22753 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 23124 17660 23152 17691
rect 23934 17660 23940 17672
rect 23124 17632 23940 17660
rect 22741 17623 22799 17629
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 24394 17620 24400 17672
rect 24452 17660 24458 17672
rect 24596 17660 24624 17700
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 26068 17737 26096 17836
rect 26237 17833 26249 17867
rect 26283 17864 26295 17867
rect 26510 17864 26516 17876
rect 26283 17836 26516 17864
rect 26283 17833 26295 17836
rect 26237 17827 26295 17833
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 27982 17864 27988 17876
rect 26620 17836 27988 17864
rect 26326 17756 26332 17808
rect 26384 17796 26390 17808
rect 26620 17796 26648 17836
rect 27540 17796 27568 17836
rect 27982 17824 27988 17836
rect 28040 17824 28046 17876
rect 28994 17864 29000 17876
rect 28184 17836 29000 17864
rect 26384 17768 26648 17796
rect 27462 17768 27568 17796
rect 26384 17756 26390 17768
rect 27614 17756 27620 17808
rect 27672 17796 27678 17808
rect 28184 17796 28212 17836
rect 28994 17824 29000 17836
rect 29052 17864 29058 17876
rect 29052 17836 30052 17864
rect 29052 17824 29058 17836
rect 27672 17768 28212 17796
rect 27672 17756 27678 17768
rect 25317 17731 25375 17737
rect 25317 17697 25329 17731
rect 25363 17697 25375 17731
rect 25705 17731 25763 17737
rect 25705 17728 25717 17731
rect 25317 17691 25375 17697
rect 25700 17697 25717 17728
rect 25751 17697 25763 17731
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 25700 17691 25763 17697
rect 25884 17700 25973 17728
rect 24452 17632 24624 17660
rect 24452 17620 24458 17632
rect 25038 17620 25044 17672
rect 25096 17660 25102 17672
rect 25332 17660 25360 17691
rect 25593 17663 25651 17669
rect 25593 17660 25605 17663
rect 25096 17632 25360 17660
rect 25424 17632 25605 17660
rect 25096 17620 25102 17632
rect 25130 17552 25136 17604
rect 25188 17592 25194 17604
rect 25424 17592 25452 17632
rect 25593 17629 25605 17632
rect 25639 17629 25651 17663
rect 25593 17623 25651 17629
rect 25188 17564 25452 17592
rect 25188 17552 25194 17564
rect 19852 17496 20760 17524
rect 19852 17484 19858 17496
rect 21634 17484 21640 17536
rect 21692 17524 21698 17536
rect 23842 17524 23848 17536
rect 21692 17496 23848 17524
rect 21692 17484 21698 17496
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 24118 17484 24124 17536
rect 24176 17524 24182 17536
rect 24857 17527 24915 17533
rect 24857 17524 24869 17527
rect 24176 17496 24869 17524
rect 24176 17484 24182 17496
rect 24857 17493 24869 17496
rect 24903 17493 24915 17527
rect 24857 17487 24915 17493
rect 24946 17484 24952 17536
rect 25004 17484 25010 17536
rect 25424 17524 25452 17564
rect 25498 17552 25504 17604
rect 25556 17592 25562 17604
rect 25700 17592 25728 17691
rect 25884 17672 25912 17700
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 26053 17731 26111 17737
rect 26053 17697 26065 17731
rect 26099 17728 26111 17731
rect 26418 17728 26424 17740
rect 26099 17700 26424 17728
rect 26099 17697 26111 17700
rect 26053 17691 26111 17697
rect 26418 17688 26424 17700
rect 26476 17688 26482 17740
rect 28184 17737 28212 17768
rect 28350 17756 28356 17808
rect 28408 17796 28414 17808
rect 28408 17768 28566 17796
rect 28408 17756 28414 17768
rect 29638 17756 29644 17808
rect 29696 17796 29702 17808
rect 29733 17799 29791 17805
rect 29733 17796 29745 17799
rect 29696 17768 29745 17796
rect 29696 17756 29702 17768
rect 29733 17765 29745 17768
rect 29779 17765 29791 17799
rect 29733 17759 29791 17765
rect 30024 17740 30052 17836
rect 28169 17731 28227 17737
rect 28169 17697 28181 17731
rect 28215 17697 28227 17731
rect 28169 17691 28227 17697
rect 30006 17688 30012 17740
rect 30064 17688 30070 17740
rect 30190 17688 30196 17740
rect 30248 17728 30254 17740
rect 30469 17731 30527 17737
rect 30469 17728 30481 17731
rect 30248 17700 30481 17728
rect 30248 17688 30254 17700
rect 30469 17697 30481 17700
rect 30515 17728 30527 17731
rect 30745 17731 30803 17737
rect 30745 17728 30757 17731
rect 30515 17700 30757 17728
rect 30515 17697 30527 17700
rect 30469 17691 30527 17697
rect 30745 17697 30757 17700
rect 30791 17697 30803 17731
rect 30745 17691 30803 17697
rect 25866 17620 25872 17672
rect 25924 17620 25930 17672
rect 26142 17620 26148 17672
rect 26200 17660 26206 17672
rect 27893 17663 27951 17669
rect 27893 17660 27905 17663
rect 26200 17632 27905 17660
rect 26200 17620 26206 17632
rect 27893 17629 27905 17632
rect 27939 17629 27951 17663
rect 27893 17623 27951 17629
rect 29638 17620 29644 17672
rect 29696 17660 29702 17672
rect 30098 17660 30104 17672
rect 29696 17632 30104 17660
rect 29696 17620 29702 17632
rect 30098 17620 30104 17632
rect 30156 17620 30162 17672
rect 26878 17592 26884 17604
rect 25556 17564 25728 17592
rect 26344 17564 26884 17592
rect 25556 17552 25562 17564
rect 26344 17524 26372 17564
rect 26878 17552 26884 17564
rect 26936 17552 26942 17604
rect 28350 17592 28356 17604
rect 28184 17564 28356 17592
rect 25424 17496 26372 17524
rect 26418 17484 26424 17536
rect 26476 17484 26482 17536
rect 26602 17484 26608 17536
rect 26660 17524 26666 17536
rect 28184 17524 28212 17564
rect 28350 17552 28356 17564
rect 28408 17552 28414 17604
rect 26660 17496 28212 17524
rect 26660 17484 26666 17496
rect 28258 17484 28264 17536
rect 28316 17484 28322 17536
rect 28626 17484 28632 17536
rect 28684 17524 28690 17536
rect 30193 17527 30251 17533
rect 30193 17524 30205 17527
rect 28684 17496 30205 17524
rect 28684 17484 28690 17496
rect 30193 17493 30205 17496
rect 30239 17493 30251 17527
rect 30193 17487 30251 17493
rect 30282 17484 30288 17536
rect 30340 17524 30346 17536
rect 30837 17527 30895 17533
rect 30837 17524 30849 17527
rect 30340 17496 30849 17524
rect 30340 17484 30346 17496
rect 30837 17493 30849 17496
rect 30883 17493 30895 17527
rect 30837 17487 30895 17493
rect 552 17434 31648 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 11436 17434
rect 11488 17382 11500 17434
rect 11552 17382 11564 17434
rect 11616 17382 11628 17434
rect 11680 17382 11692 17434
rect 11744 17382 19210 17434
rect 19262 17382 19274 17434
rect 19326 17382 19338 17434
rect 19390 17382 19402 17434
rect 19454 17382 19466 17434
rect 19518 17382 26984 17434
rect 27036 17382 27048 17434
rect 27100 17382 27112 17434
rect 27164 17382 27176 17434
rect 27228 17382 27240 17434
rect 27292 17382 31648 17434
rect 552 17360 31648 17382
rect 2406 17320 2412 17332
rect 1412 17292 2412 17320
rect 1213 17119 1271 17125
rect 1213 17085 1225 17119
rect 1259 17116 1271 17119
rect 1412 17116 1440 17292
rect 2406 17280 2412 17292
rect 2464 17280 2470 17332
rect 2498 17280 2504 17332
rect 2556 17320 2562 17332
rect 2556 17292 4292 17320
rect 2556 17280 2562 17292
rect 1489 17255 1547 17261
rect 1489 17221 1501 17255
rect 1535 17252 1547 17255
rect 3050 17252 3056 17264
rect 1535 17224 3056 17252
rect 1535 17221 1547 17224
rect 1489 17215 1547 17221
rect 3050 17212 3056 17224
rect 3108 17212 3114 17264
rect 4264 17261 4292 17292
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 6086 17320 6092 17332
rect 5316 17292 6092 17320
rect 5316 17280 5322 17292
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 6822 17320 6828 17332
rect 6696 17292 6828 17320
rect 6696 17280 6702 17292
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 7006 17320 7012 17332
rect 6963 17292 7012 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 8294 17320 8300 17332
rect 7340 17292 8300 17320
rect 7340 17280 7346 17292
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 8481 17323 8539 17329
rect 8481 17320 8493 17323
rect 8444 17292 8493 17320
rect 8444 17280 8450 17292
rect 8481 17289 8493 17292
rect 8527 17289 8539 17323
rect 8481 17283 8539 17289
rect 8754 17280 8760 17332
rect 8812 17280 8818 17332
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 11388 17292 11529 17320
rect 11388 17280 11394 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 11790 17280 11796 17332
rect 11848 17320 11854 17332
rect 14550 17320 14556 17332
rect 11848 17292 14556 17320
rect 11848 17280 11854 17292
rect 14550 17280 14556 17292
rect 14608 17320 14614 17332
rect 14737 17323 14795 17329
rect 14737 17320 14749 17323
rect 14608 17292 14749 17320
rect 14608 17280 14614 17292
rect 14737 17289 14749 17292
rect 14783 17289 14795 17323
rect 14737 17283 14795 17289
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 15620 17292 15853 17320
rect 15620 17280 15626 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 17218 17280 17224 17332
rect 17276 17320 17282 17332
rect 18414 17320 18420 17332
rect 17276 17292 18420 17320
rect 17276 17280 17282 17292
rect 18414 17280 18420 17292
rect 18472 17320 18478 17332
rect 19794 17320 19800 17332
rect 18472 17292 19800 17320
rect 18472 17280 18478 17292
rect 19794 17280 19800 17292
rect 19852 17280 19858 17332
rect 20622 17280 20628 17332
rect 20680 17320 20686 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 20680 17292 21465 17320
rect 20680 17280 20686 17292
rect 21453 17289 21465 17292
rect 21499 17320 21511 17323
rect 22373 17323 22431 17329
rect 21499 17292 22324 17320
rect 21499 17289 21511 17292
rect 21453 17283 21511 17289
rect 4157 17255 4215 17261
rect 4157 17221 4169 17255
rect 4203 17221 4215 17255
rect 4157 17215 4215 17221
rect 4249 17255 4307 17261
rect 4249 17221 4261 17255
rect 4295 17252 4307 17255
rect 5442 17252 5448 17264
rect 4295 17224 5448 17252
rect 4295 17221 4307 17224
rect 4249 17215 4307 17221
rect 2314 17184 2320 17196
rect 2240 17156 2320 17184
rect 1259 17088 1440 17116
rect 1489 17119 1547 17125
rect 1259 17085 1271 17088
rect 1213 17079 1271 17085
rect 1489 17085 1501 17119
rect 1535 17116 1547 17119
rect 1578 17116 1584 17128
rect 1535 17088 1584 17116
rect 1535 17085 1547 17088
rect 1489 17079 1547 17085
rect 1578 17076 1584 17088
rect 1636 17116 1642 17128
rect 1949 17119 2007 17125
rect 1949 17116 1961 17119
rect 1636 17088 1961 17116
rect 1636 17076 1642 17088
rect 1949 17085 1961 17088
rect 1995 17085 2007 17119
rect 1949 17079 2007 17085
rect 2038 17076 2044 17128
rect 2096 17116 2102 17128
rect 2240 17125 2268 17156
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 4062 17144 4068 17196
rect 4120 17144 4126 17196
rect 4172 17184 4200 17215
rect 5442 17212 5448 17224
rect 5500 17212 5506 17264
rect 5902 17212 5908 17264
rect 5960 17252 5966 17264
rect 12710 17252 12716 17264
rect 5960 17224 12716 17252
rect 5960 17212 5966 17224
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 13909 17255 13967 17261
rect 13909 17252 13921 17255
rect 13136 17224 13921 17252
rect 13136 17212 13142 17224
rect 13909 17221 13921 17224
rect 13955 17221 13967 17255
rect 13909 17215 13967 17221
rect 14182 17212 14188 17264
rect 14240 17212 14246 17264
rect 14660 17224 17540 17252
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 4172 17156 5028 17184
rect 2225 17119 2283 17125
rect 2096 17088 2141 17116
rect 2096 17076 2102 17088
rect 2225 17085 2237 17119
rect 2271 17085 2283 17119
rect 2225 17079 2283 17085
rect 2406 17076 2412 17128
rect 2464 17125 2470 17128
rect 2464 17116 2472 17125
rect 2464 17088 2509 17116
rect 2464 17079 2472 17088
rect 2464 17076 2470 17079
rect 3234 17076 3240 17128
rect 3292 17116 3298 17128
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 3292 17088 3617 17116
rect 3292 17076 3298 17088
rect 3605 17085 3617 17088
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4338 17116 4344 17128
rect 4212 17088 4344 17116
rect 4212 17076 4218 17088
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 5000 17125 5028 17156
rect 5368 17156 9781 17184
rect 4985 17119 5043 17125
rect 4985 17085 4997 17119
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5074 17076 5080 17128
rect 5132 17076 5138 17128
rect 5368 17125 5396 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10336 17156 11920 17184
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17116 5503 17119
rect 5626 17116 5632 17128
rect 5491 17088 5632 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 6086 17076 6092 17128
rect 6144 17116 6150 17128
rect 7101 17119 7159 17125
rect 6144 17088 6592 17116
rect 6144 17076 6150 17088
rect 1305 17051 1363 17057
rect 1305 17017 1317 17051
rect 1351 17048 1363 17051
rect 2130 17048 2136 17060
rect 1351 17020 2136 17048
rect 1351 17017 1363 17020
rect 1305 17011 1363 17017
rect 1210 16940 1216 16992
rect 1268 16980 1274 16992
rect 1320 16980 1348 17011
rect 2130 17008 2136 17020
rect 2188 17048 2194 17060
rect 2317 17051 2375 17057
rect 2317 17048 2329 17051
rect 2188 17020 2329 17048
rect 2188 17008 2194 17020
rect 2317 17017 2329 17020
rect 2363 17017 2375 17051
rect 2317 17011 2375 17017
rect 4706 17008 4712 17060
rect 4764 17048 4770 17060
rect 5166 17048 5172 17060
rect 4764 17020 5172 17048
rect 4764 17008 4770 17020
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 6454 17048 6460 17060
rect 5592 17020 6460 17048
rect 5592 17008 5598 17020
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 6564 17048 6592 17088
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 7190 17116 7196 17128
rect 7147 17088 7196 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 7282 17076 7288 17128
rect 7340 17076 7346 17128
rect 7377 17119 7435 17125
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 7466 17116 7472 17128
rect 7423 17088 7472 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 8386 17076 8392 17128
rect 8444 17076 8450 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8754 17116 8760 17128
rect 8619 17088 8760 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 10042 17076 10048 17128
rect 10100 17076 10106 17128
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 8478 17048 8484 17060
rect 6564 17020 8484 17048
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 9582 17008 9588 17060
rect 9640 17048 9646 17060
rect 10137 17051 10195 17057
rect 10137 17048 10149 17051
rect 9640 17020 10149 17048
rect 9640 17008 9646 17020
rect 10137 17017 10149 17020
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 1268 16952 1348 16980
rect 2593 16983 2651 16989
rect 1268 16940 1274 16952
rect 2593 16949 2605 16983
rect 2639 16980 2651 16983
rect 2866 16980 2872 16992
rect 2639 16952 2872 16980
rect 2639 16949 2651 16952
rect 2593 16943 2651 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3142 16940 3148 16992
rect 3200 16980 3206 16992
rect 3329 16983 3387 16989
rect 3329 16980 3341 16983
rect 3200 16952 3341 16980
rect 3200 16940 3206 16952
rect 3329 16949 3341 16952
rect 3375 16949 3387 16983
rect 3329 16943 3387 16949
rect 4798 16940 4804 16992
rect 4856 16940 4862 16992
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 5258 16980 5264 16992
rect 5040 16952 5264 16980
rect 5040 16940 5046 16952
rect 5258 16940 5264 16952
rect 5316 16980 5322 16992
rect 7282 16980 7288 16992
rect 5316 16952 7288 16980
rect 5316 16940 5322 16952
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 7466 16940 7472 16992
rect 7524 16980 7530 16992
rect 10336 16980 10364 17156
rect 10410 17076 10416 17128
rect 10468 17076 10474 17128
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17116 10563 17119
rect 10870 17116 10876 17128
rect 10551 17088 10876 17116
rect 10551 17085 10563 17088
rect 10505 17079 10563 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 11701 17119 11759 17125
rect 11701 17116 11713 17119
rect 11388 17088 11713 17116
rect 11388 17076 11394 17088
rect 11701 17085 11713 17088
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 11892 17116 11920 17156
rect 11974 17144 11980 17196
rect 12032 17184 12038 17196
rect 12069 17187 12127 17193
rect 12069 17184 12081 17187
rect 12032 17156 12081 17184
rect 12032 17144 12038 17156
rect 12069 17153 12081 17156
rect 12115 17153 12127 17187
rect 12069 17147 12127 17153
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 14660 17184 14688 17224
rect 12268 17156 14688 17184
rect 12268 17116 12296 17156
rect 11892 17088 12296 17116
rect 14093 17119 14151 17125
rect 14093 17085 14105 17119
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 12434 17048 12440 17060
rect 11992 17020 12440 17048
rect 7524 16952 10364 16980
rect 7524 16940 7530 16952
rect 11054 16940 11060 16992
rect 11112 16980 11118 16992
rect 11514 16980 11520 16992
rect 11112 16952 11520 16980
rect 11112 16940 11118 16952
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11992 16989 12020 17020
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 12805 17051 12863 17057
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 12989 17051 13047 17057
rect 12989 17048 13001 17051
rect 12851 17020 13001 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 12989 17017 13001 17020
rect 13035 17048 13047 17051
rect 13035 17020 13492 17048
rect 13035 17017 13047 17020
rect 12989 17011 13047 17017
rect 11977 16983 12035 16989
rect 11977 16949 11989 16983
rect 12023 16949 12035 16983
rect 11977 16943 12035 16949
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12768 16952 13093 16980
rect 12768 16940 12774 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13464 16980 13492 17020
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 14108 17048 14136 17079
rect 14274 17076 14280 17128
rect 14332 17076 14338 17128
rect 14366 17076 14372 17128
rect 14424 17076 14430 17128
rect 14550 17076 14556 17128
rect 14608 17076 14614 17128
rect 14660 17125 14688 17156
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 14884 17156 16221 17184
rect 14884 17144 14890 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16298 17144 16304 17196
rect 16356 17144 16362 17196
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 16816 17156 17448 17184
rect 16816 17144 16822 17156
rect 17420 17128 17448 17156
rect 14645 17119 14703 17125
rect 14645 17085 14657 17119
rect 14691 17085 14703 17119
rect 14645 17079 14703 17085
rect 15010 17076 15016 17128
rect 15068 17076 15074 17128
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15804 17088 16037 17116
rect 15804 17076 15810 17088
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 16632 17088 17233 17116
rect 16632 17076 16638 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 17402 17076 17408 17128
rect 17460 17076 17466 17128
rect 17512 17116 17540 17224
rect 18138 17212 18144 17264
rect 18196 17212 18202 17264
rect 20990 17252 20996 17264
rect 19260 17224 20996 17252
rect 18046 17144 18052 17196
rect 18104 17184 18110 17196
rect 18104 17156 19196 17184
rect 18104 17144 18110 17156
rect 18966 17116 18972 17128
rect 17512 17088 18972 17116
rect 18966 17076 18972 17088
rect 19024 17125 19030 17128
rect 19168 17125 19196 17156
rect 19260 17125 19288 17224
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 22186 17252 22192 17264
rect 22112 17224 22192 17252
rect 21634 17184 21640 17196
rect 19536 17156 21640 17184
rect 19024 17119 19073 17125
rect 19024 17085 19027 17119
rect 19061 17085 19073 17119
rect 19024 17079 19073 17085
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 19245 17119 19303 17125
rect 19245 17085 19257 17119
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 19024 17076 19030 17079
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19536 17125 19564 17156
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 19428 17119 19486 17125
rect 19428 17116 19440 17119
rect 19392 17088 19440 17116
rect 19392 17076 19398 17088
rect 19428 17085 19440 17088
rect 19474 17085 19486 17119
rect 19428 17079 19486 17085
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 15102 17048 15108 17060
rect 13596 17020 13860 17048
rect 14108 17020 15108 17048
rect 13596 17008 13602 17020
rect 13722 16980 13728 16992
rect 13464 16952 13728 16980
rect 13081 16943 13139 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 13832 16980 13860 17020
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 15378 17008 15384 17060
rect 15436 17048 15442 17060
rect 16758 17048 16764 17060
rect 15436 17020 16764 17048
rect 15436 17008 15442 17020
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 16850 17008 16856 17060
rect 16908 17048 16914 17060
rect 16908 17020 17356 17048
rect 16908 17008 16914 17020
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 13832 16952 15209 16980
rect 15197 16949 15209 16952
rect 15243 16980 15255 16983
rect 16942 16980 16948 16992
rect 15243 16952 16948 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17328 16989 17356 17020
rect 17494 17008 17500 17060
rect 17552 17048 17558 17060
rect 18509 17051 18567 17057
rect 17552 17020 18276 17048
rect 17552 17008 17558 17020
rect 17313 16983 17371 16989
rect 17313 16949 17325 16983
rect 17359 16949 17371 16983
rect 17313 16943 17371 16949
rect 18046 16940 18052 16992
rect 18104 16940 18110 16992
rect 18248 16980 18276 17020
rect 18509 17017 18521 17051
rect 18555 17048 18567 17051
rect 18598 17048 18604 17060
rect 18555 17020 18604 17048
rect 18555 17017 18567 17020
rect 18509 17011 18567 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 19447 17048 19475 17079
rect 19610 17076 19616 17128
rect 19668 17116 19674 17128
rect 19794 17116 19800 17128
rect 19668 17088 19800 17116
rect 19668 17076 19674 17088
rect 19794 17076 19800 17088
rect 19852 17116 19858 17128
rect 19889 17119 19947 17125
rect 19889 17116 19901 17119
rect 19852 17088 19901 17116
rect 19852 17076 19858 17088
rect 19889 17085 19901 17088
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 19978 17076 19984 17128
rect 20036 17076 20042 17128
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 20128 17088 20177 17116
rect 20128 17076 20134 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 20180 17048 20208 17079
rect 20254 17076 20260 17128
rect 20312 17076 20318 17128
rect 21358 17076 21364 17128
rect 21416 17076 21422 17128
rect 21545 17119 21603 17125
rect 21545 17085 21557 17119
rect 21591 17116 21603 17119
rect 21726 17116 21732 17128
rect 21591 17088 21732 17116
rect 21591 17085 21603 17088
rect 21545 17079 21603 17085
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 21818 17076 21824 17128
rect 21876 17116 21882 17128
rect 22112 17125 22140 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22296 17252 22324 17292
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 23382 17320 23388 17332
rect 22419 17292 23388 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 24026 17320 24032 17332
rect 23523 17292 24032 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 24026 17280 24032 17292
rect 24084 17280 24090 17332
rect 24762 17320 24768 17332
rect 24421 17292 24768 17320
rect 22296 17224 22600 17252
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 21876 17088 21925 17116
rect 21876 17076 21882 17088
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17085 22155 17119
rect 22462 17116 22468 17128
rect 22097 17079 22155 17085
rect 22204 17088 22468 17116
rect 22204 17048 22232 17088
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 22572 17125 22600 17224
rect 22738 17212 22744 17264
rect 22796 17212 22802 17264
rect 23842 17212 23848 17264
rect 23900 17252 23906 17264
rect 24421 17252 24449 17292
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 25958 17280 25964 17332
rect 26016 17320 26022 17332
rect 26053 17323 26111 17329
rect 26053 17320 26065 17323
rect 26016 17292 26065 17320
rect 26016 17280 26022 17292
rect 26053 17289 26065 17292
rect 26099 17320 26111 17323
rect 27154 17320 27160 17332
rect 26099 17292 27160 17320
rect 26099 17289 26111 17292
rect 26053 17283 26111 17289
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 27522 17280 27528 17332
rect 27580 17280 27586 17332
rect 28261 17323 28319 17329
rect 28261 17289 28273 17323
rect 28307 17320 28319 17323
rect 29270 17320 29276 17332
rect 28307 17292 29276 17320
rect 28307 17289 28319 17292
rect 28261 17283 28319 17289
rect 29270 17280 29276 17292
rect 29328 17280 29334 17332
rect 29454 17320 29460 17332
rect 29380 17292 29460 17320
rect 23900 17224 24449 17252
rect 23900 17212 23906 17224
rect 26234 17212 26240 17264
rect 26292 17252 26298 17264
rect 27540 17252 27568 17280
rect 29380 17252 29408 17292
rect 29454 17280 29460 17292
rect 29512 17320 29518 17332
rect 30742 17320 30748 17332
rect 29512 17292 30748 17320
rect 29512 17280 29518 17292
rect 30742 17280 30748 17292
rect 30800 17280 30806 17332
rect 31110 17280 31116 17332
rect 31168 17280 31174 17332
rect 26292 17224 27568 17252
rect 28736 17224 29408 17252
rect 26292 17212 26298 17224
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17184 22891 17187
rect 23474 17184 23480 17196
rect 22879 17156 23480 17184
rect 22879 17153 22891 17156
rect 22833 17147 22891 17153
rect 23474 17144 23480 17156
rect 23532 17144 23538 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24305 17187 24363 17193
rect 24305 17184 24317 17187
rect 23992 17156 24317 17184
rect 23992 17144 23998 17156
rect 24305 17153 24317 17156
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 24581 17187 24639 17193
rect 24581 17153 24593 17187
rect 24627 17184 24639 17187
rect 24946 17184 24952 17196
rect 24627 17156 24952 17184
rect 24627 17153 24639 17156
rect 24581 17147 24639 17153
rect 24946 17144 24952 17156
rect 25004 17144 25010 17196
rect 27338 17184 27344 17196
rect 26436 17156 27344 17184
rect 22557 17119 22615 17125
rect 22557 17085 22569 17119
rect 22603 17085 22615 17119
rect 22557 17079 22615 17085
rect 22738 17076 22744 17128
rect 22796 17116 22802 17128
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22796 17088 22937 17116
rect 22796 17076 22802 17088
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 22925 17079 22983 17085
rect 23014 17076 23020 17128
rect 23072 17076 23078 17128
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17085 23167 17119
rect 23109 17079 23167 17085
rect 18708 17020 19334 17048
rect 19447 17020 19840 17048
rect 20180 17020 22232 17048
rect 18708 16980 18736 17020
rect 18248 16952 18736 16980
rect 18782 16940 18788 16992
rect 18840 16980 18846 16992
rect 18877 16983 18935 16989
rect 18877 16980 18889 16983
rect 18840 16952 18889 16980
rect 18840 16940 18846 16952
rect 18877 16949 18889 16952
rect 18923 16949 18935 16983
rect 19306 16980 19334 17020
rect 19610 16980 19616 16992
rect 19306 16952 19616 16980
rect 18877 16943 18935 16949
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 19702 16940 19708 16992
rect 19760 16940 19766 16992
rect 19812 16980 19840 17020
rect 22278 17008 22284 17060
rect 22336 17048 22342 17060
rect 23124 17048 23152 17079
rect 23842 17076 23848 17128
rect 23900 17076 23906 17128
rect 24026 17076 24032 17128
rect 24084 17076 24090 17128
rect 26050 17116 26056 17128
rect 25714 17088 26056 17116
rect 26050 17076 26056 17088
rect 26108 17076 26114 17128
rect 26436 17125 26464 17156
rect 27338 17144 27344 17156
rect 27396 17184 27402 17196
rect 27522 17184 27528 17196
rect 27396 17156 27528 17184
rect 27396 17144 27402 17156
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 27982 17144 27988 17196
rect 28040 17144 28046 17196
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 28736 17184 28764 17224
rect 28500 17156 28764 17184
rect 29365 17187 29423 17193
rect 28500 17144 28506 17156
rect 29365 17153 29377 17187
rect 29411 17184 29423 17187
rect 30006 17184 30012 17196
rect 29411 17156 30012 17184
rect 29411 17153 29423 17156
rect 29365 17147 29423 17153
rect 30006 17144 30012 17156
rect 30064 17144 30070 17196
rect 26421 17119 26479 17125
rect 26421 17085 26433 17119
rect 26467 17085 26479 17119
rect 26421 17079 26479 17085
rect 26881 17119 26939 17125
rect 26881 17085 26893 17119
rect 26927 17085 26939 17119
rect 26881 17079 26939 17085
rect 23382 17048 23388 17060
rect 22336 17020 23060 17048
rect 23124 17020 23388 17048
rect 22336 17008 22342 17020
rect 21082 16980 21088 16992
rect 19812 16952 21088 16980
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21358 16940 21364 16992
rect 21416 16980 21422 16992
rect 21729 16983 21787 16989
rect 21729 16980 21741 16983
rect 21416 16952 21741 16980
rect 21416 16940 21422 16952
rect 21729 16949 21741 16952
rect 21775 16980 21787 16983
rect 22002 16980 22008 16992
rect 21775 16952 22008 16980
rect 21775 16949 21787 16952
rect 21729 16943 21787 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22189 16983 22247 16989
rect 22189 16949 22201 16983
rect 22235 16980 22247 16983
rect 22922 16980 22928 16992
rect 22235 16952 22928 16980
rect 22235 16949 22247 16952
rect 22189 16943 22247 16949
rect 22922 16940 22928 16952
rect 22980 16940 22986 16992
rect 23032 16980 23060 17020
rect 23382 17008 23388 17020
rect 23440 17008 23446 17060
rect 23566 17008 23572 17060
rect 23624 17008 23630 17060
rect 26145 17051 26203 17057
rect 26145 17048 26157 17051
rect 24136 17020 24992 17048
rect 24136 16980 24164 17020
rect 23032 16952 24164 16980
rect 24213 16983 24271 16989
rect 24213 16949 24225 16983
rect 24259 16980 24271 16983
rect 24670 16980 24676 16992
rect 24259 16952 24676 16980
rect 24259 16949 24271 16952
rect 24213 16943 24271 16949
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 24964 16980 24992 17020
rect 25976 17020 26157 17048
rect 25590 16980 25596 16992
rect 24964 16952 25596 16980
rect 25590 16940 25596 16952
rect 25648 16980 25654 16992
rect 25976 16980 26004 17020
rect 26145 17017 26157 17020
rect 26191 17017 26203 17051
rect 26896 17048 26924 17079
rect 26970 17076 26976 17128
rect 27028 17116 27034 17128
rect 27065 17119 27123 17125
rect 27065 17116 27077 17119
rect 27028 17088 27077 17116
rect 27028 17076 27034 17088
rect 27065 17085 27077 17088
rect 27111 17085 27123 17119
rect 27709 17119 27767 17125
rect 27065 17079 27123 17085
rect 27172 17088 27660 17116
rect 27172 17048 27200 17088
rect 26145 17011 26203 17017
rect 26528 17020 27200 17048
rect 25648 16952 26004 16980
rect 25648 16940 25654 16952
rect 26050 16940 26056 16992
rect 26108 16980 26114 16992
rect 26528 16980 26556 17020
rect 27338 17008 27344 17060
rect 27396 17048 27402 17060
rect 27525 17051 27583 17057
rect 27525 17048 27537 17051
rect 27396 17020 27537 17048
rect 27396 17008 27402 17020
rect 27525 17017 27537 17020
rect 27571 17017 27583 17051
rect 27525 17011 27583 17017
rect 26108 16952 26556 16980
rect 26108 16940 26114 16952
rect 26602 16940 26608 16992
rect 26660 16980 26666 16992
rect 27433 16983 27491 16989
rect 27433 16980 27445 16983
rect 26660 16952 27445 16980
rect 26660 16940 26666 16952
rect 27433 16949 27445 16952
rect 27479 16949 27491 16983
rect 27632 16980 27660 17088
rect 27709 17085 27721 17119
rect 27755 17085 27767 17119
rect 27709 17079 27767 17085
rect 27724 17048 27752 17079
rect 27890 17076 27896 17128
rect 27948 17076 27954 17128
rect 28000 17116 28028 17144
rect 28077 17119 28135 17125
rect 28077 17116 28089 17119
rect 28000 17088 28089 17116
rect 28077 17085 28089 17088
rect 28123 17085 28135 17119
rect 28077 17079 28135 17085
rect 28353 17119 28411 17125
rect 28353 17085 28365 17119
rect 28399 17116 28411 17119
rect 28399 17088 29132 17116
rect 28399 17085 28411 17088
rect 28353 17079 28411 17085
rect 27985 17051 28043 17057
rect 27724 17020 27936 17048
rect 27798 16980 27804 16992
rect 27632 16952 27804 16980
rect 27433 16943 27491 16949
rect 27798 16940 27804 16952
rect 27856 16940 27862 16992
rect 27908 16980 27936 17020
rect 27985 17017 27997 17051
rect 28031 17048 28043 17051
rect 28442 17048 28448 17060
rect 28031 17020 28448 17048
rect 28031 17017 28043 17020
rect 27985 17011 28043 17017
rect 28442 17008 28448 17020
rect 28500 17008 28506 17060
rect 28629 17051 28687 17057
rect 28629 17017 28641 17051
rect 28675 17048 28687 17051
rect 28902 17048 28908 17060
rect 28675 17020 28908 17048
rect 28675 17017 28687 17020
rect 28629 17011 28687 17017
rect 28902 17008 28908 17020
rect 28960 17008 28966 17060
rect 28810 16980 28816 16992
rect 27908 16952 28816 16980
rect 28810 16940 28816 16952
rect 28868 16940 28874 16992
rect 29104 16989 29132 17088
rect 29270 17076 29276 17128
rect 29328 17076 29334 17128
rect 29178 17008 29184 17060
rect 29236 17048 29242 17060
rect 29641 17051 29699 17057
rect 29641 17048 29653 17051
rect 29236 17020 29653 17048
rect 29236 17008 29242 17020
rect 29641 17017 29653 17020
rect 29687 17017 29699 17051
rect 29641 17011 29699 17017
rect 29730 17008 29736 17060
rect 29788 17048 29794 17060
rect 30098 17048 30104 17060
rect 29788 17020 30104 17048
rect 29788 17008 29794 17020
rect 30098 17008 30104 17020
rect 30156 17008 30162 17060
rect 29089 16983 29147 16989
rect 29089 16949 29101 16983
rect 29135 16980 29147 16983
rect 30466 16980 30472 16992
rect 29135 16952 30472 16980
rect 29135 16949 29147 16952
rect 29089 16943 29147 16949
rect 30466 16940 30472 16952
rect 30524 16940 30530 16992
rect 552 16890 31648 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 12096 16890
rect 12148 16838 12160 16890
rect 12212 16838 12224 16890
rect 12276 16838 12288 16890
rect 12340 16838 12352 16890
rect 12404 16838 19870 16890
rect 19922 16838 19934 16890
rect 19986 16838 19998 16890
rect 20050 16838 20062 16890
rect 20114 16838 20126 16890
rect 20178 16838 27644 16890
rect 27696 16838 27708 16890
rect 27760 16838 27772 16890
rect 27824 16838 27836 16890
rect 27888 16838 27900 16890
rect 27952 16838 31648 16890
rect 552 16816 31648 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 4982 16776 4988 16788
rect 1728 16748 4988 16776
rect 1728 16736 1734 16748
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 5132 16748 5457 16776
rect 5132 16736 5138 16748
rect 5445 16745 5457 16748
rect 5491 16745 5503 16779
rect 5445 16739 5503 16745
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 6178 16776 6184 16788
rect 5951 16748 6184 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 6638 16776 6644 16788
rect 6595 16748 6644 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 8662 16776 8668 16788
rect 6748 16748 8668 16776
rect 658 16668 664 16720
rect 716 16708 722 16720
rect 4154 16708 4160 16720
rect 716 16680 4160 16708
rect 716 16668 722 16680
rect 4154 16668 4160 16680
rect 4212 16668 4218 16720
rect 5166 16708 5172 16720
rect 4908 16680 5172 16708
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 2792 16504 2820 16603
rect 2866 16600 2872 16652
rect 2924 16600 2930 16652
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 4908 16640 4936 16680
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 6748 16708 6776 16748
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 11606 16736 11612 16788
rect 11664 16776 11670 16788
rect 11701 16779 11759 16785
rect 11701 16776 11713 16779
rect 11664 16748 11713 16776
rect 11664 16736 11670 16748
rect 11701 16745 11713 16748
rect 11747 16745 11759 16779
rect 11701 16739 11759 16745
rect 11974 16736 11980 16788
rect 12032 16776 12038 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 12032 16748 12357 16776
rect 12032 16736 12038 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 12492 16748 12725 16776
rect 12492 16736 12498 16748
rect 12713 16745 12725 16748
rect 12759 16776 12771 16779
rect 12894 16776 12900 16788
rect 12759 16748 12900 16776
rect 12759 16745 12771 16748
rect 12713 16739 12771 16745
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13354 16736 13360 16788
rect 13412 16736 13418 16788
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16745 15807 16779
rect 15749 16739 15807 16745
rect 7190 16708 7196 16720
rect 5276 16680 6316 16708
rect 3191 16612 4936 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 4982 16600 4988 16652
rect 5040 16600 5046 16652
rect 5276 16649 5304 16680
rect 6288 16652 6316 16680
rect 6472 16680 6776 16708
rect 6840 16680 7196 16708
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 5994 16600 6000 16652
rect 6052 16640 6058 16652
rect 6089 16643 6147 16649
rect 6089 16640 6101 16643
rect 6052 16612 6101 16640
rect 6052 16600 6058 16612
rect 6089 16609 6101 16612
rect 6135 16609 6147 16643
rect 6089 16603 6147 16609
rect 6270 16600 6276 16652
rect 6328 16600 6334 16652
rect 6362 16600 6368 16652
rect 6420 16600 6426 16652
rect 3050 16532 3056 16584
rect 3108 16532 3114 16584
rect 4890 16532 4896 16584
rect 4948 16572 4954 16584
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 4948 16544 5089 16572
rect 4948 16532 4954 16544
rect 5077 16541 5089 16544
rect 5123 16541 5135 16575
rect 5077 16535 5135 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16572 5227 16575
rect 5534 16572 5540 16584
rect 5215 16544 5540 16572
rect 5215 16541 5227 16544
rect 5169 16535 5227 16541
rect 2866 16504 2872 16516
rect 2792 16476 2872 16504
rect 2866 16464 2872 16476
rect 2924 16504 2930 16516
rect 3142 16504 3148 16516
rect 2924 16476 3148 16504
rect 2924 16464 2930 16476
rect 3142 16464 3148 16476
rect 3200 16464 3206 16516
rect 5092 16504 5120 16535
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 6472 16504 6500 16680
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6840 16649 6868 16680
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 8202 16668 8208 16720
rect 8260 16668 8266 16720
rect 10134 16708 10140 16720
rect 9324 16680 10140 16708
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6604 16612 6745 16640
rect 6604 16600 6610 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 6733 16603 6791 16609
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16609 6883 16643
rect 6825 16603 6883 16609
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16640 7067 16643
rect 7837 16643 7895 16649
rect 7837 16640 7849 16643
rect 7055 16612 7849 16640
rect 7055 16609 7067 16612
rect 7009 16603 7067 16609
rect 7837 16609 7849 16612
rect 7883 16609 7895 16643
rect 7837 16603 7895 16609
rect 8018 16600 8024 16652
rect 8076 16600 8082 16652
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 8478 16640 8484 16652
rect 8435 16612 8484 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 9324 16649 9352 16680
rect 10134 16668 10140 16680
rect 10192 16668 10198 16720
rect 11517 16711 11575 16717
rect 11517 16677 11529 16711
rect 11563 16708 11575 16711
rect 14918 16708 14924 16720
rect 11563 16680 11924 16708
rect 11563 16677 11575 16680
rect 11517 16671 11575 16677
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16609 9367 16643
rect 9309 16603 9367 16609
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16609 9459 16643
rect 9401 16603 9459 16609
rect 6914 16532 6920 16584
rect 6972 16532 6978 16584
rect 7558 16532 7564 16584
rect 7616 16572 7622 16584
rect 9416 16572 9444 16603
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 11146 16640 11152 16652
rect 9815 16612 11152 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 11896 16640 11924 16680
rect 12452 16680 14924 16708
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11896 16612 11989 16640
rect 11977 16609 11989 16612
rect 12023 16640 12035 16643
rect 12452 16640 12480 16680
rect 14918 16668 14924 16680
rect 14976 16668 14982 16720
rect 15764 16708 15792 16739
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16172 16748 16681 16776
rect 16172 16736 16178 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 16816 16748 17417 16776
rect 16816 16736 16822 16748
rect 17405 16745 17417 16748
rect 17451 16776 17463 16779
rect 18230 16776 18236 16788
rect 17451 16748 18236 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 18230 16736 18236 16748
rect 18288 16776 18294 16788
rect 18414 16776 18420 16788
rect 18288 16748 18420 16776
rect 18288 16736 18294 16748
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 18598 16776 18604 16788
rect 18524 16748 18604 16776
rect 16022 16708 16028 16720
rect 15764 16680 16028 16708
rect 16022 16668 16028 16680
rect 16080 16708 16086 16720
rect 16080 16680 16344 16708
rect 16080 16668 16086 16680
rect 12023 16612 12480 16640
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 12526 16600 12532 16652
rect 12584 16600 12590 16652
rect 12802 16600 12808 16652
rect 12860 16600 12866 16652
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13136 16612 13553 16640
rect 13136 16600 13142 16612
rect 13541 16609 13553 16612
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13814 16600 13820 16652
rect 13872 16600 13878 16652
rect 15930 16600 15936 16652
rect 15988 16600 15994 16652
rect 16316 16649 16344 16680
rect 16500 16680 17632 16708
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16390 16600 16396 16652
rect 16448 16600 16454 16652
rect 7616 16544 9444 16572
rect 7616 16532 7622 16544
rect 10042 16532 10048 16584
rect 10100 16572 10106 16584
rect 11054 16572 11060 16584
rect 10100 16544 11060 16572
rect 10100 16532 10106 16544
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 11885 16575 11943 16581
rect 11885 16572 11897 16575
rect 11388 16544 11897 16572
rect 11388 16532 11394 16544
rect 11885 16541 11897 16544
rect 11931 16541 11943 16575
rect 11885 16535 11943 16541
rect 12066 16532 12072 16584
rect 12124 16532 12130 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16541 12219 16575
rect 12161 16535 12219 16541
rect 7466 16504 7472 16516
rect 5092 16476 6500 16504
rect 6748 16476 7472 16504
rect 2961 16439 3019 16445
rect 2961 16405 2973 16439
rect 3007 16436 3019 16439
rect 4798 16436 4804 16448
rect 3007 16408 4804 16436
rect 3007 16405 3019 16408
rect 2961 16399 3019 16405
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 6748 16436 6776 16476
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 8294 16464 8300 16516
rect 8352 16504 8358 16516
rect 10318 16504 10324 16516
rect 8352 16476 10324 16504
rect 8352 16464 8358 16476
rect 10318 16464 10324 16476
rect 10376 16504 10382 16516
rect 11698 16504 11704 16516
rect 10376 16476 11704 16504
rect 10376 16464 10382 16476
rect 11698 16464 11704 16476
rect 11756 16504 11762 16516
rect 12176 16504 12204 16535
rect 13630 16532 13636 16584
rect 13688 16532 13694 16584
rect 13722 16532 13728 16584
rect 13780 16532 13786 16584
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 16022 16572 16028 16584
rect 14424 16544 16028 16572
rect 14424 16532 14430 16544
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 16500 16572 16528 16680
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 16132 16544 16528 16572
rect 16592 16572 16620 16603
rect 16666 16600 16672 16652
rect 16724 16600 16730 16652
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16899 16612 16957 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 16945 16609 16957 16612
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 17092 16612 17141 16640
rect 17092 16600 17098 16612
rect 17129 16609 17141 16612
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17494 16600 17500 16652
rect 17552 16600 17558 16652
rect 17604 16649 17632 16680
rect 18322 16668 18328 16720
rect 18380 16708 18386 16720
rect 18524 16708 18552 16748
rect 18598 16736 18604 16748
rect 18656 16776 18662 16788
rect 19702 16776 19708 16788
rect 18656 16748 19708 16776
rect 18656 16736 18662 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 21082 16776 21088 16788
rect 20763 16748 21088 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 20732 16708 20760 16739
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 22066 16748 24808 16776
rect 18380 16680 18552 16708
rect 18708 16680 20760 16708
rect 18380 16668 18386 16680
rect 18708 16649 18736 16680
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 21269 16711 21327 16717
rect 21269 16708 21281 16711
rect 20864 16680 21281 16708
rect 20864 16668 20870 16680
rect 21269 16677 21281 16680
rect 21315 16677 21327 16711
rect 22066 16708 22094 16748
rect 21269 16671 21327 16677
rect 21376 16680 22094 16708
rect 22741 16711 22799 16717
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 18693 16643 18751 16649
rect 18693 16609 18705 16643
rect 18739 16609 18751 16643
rect 18693 16603 18751 16609
rect 18877 16643 18935 16649
rect 18877 16609 18889 16643
rect 18923 16640 18935 16643
rect 19334 16640 19340 16652
rect 18923 16612 19340 16640
rect 18923 16609 18935 16612
rect 18877 16603 18935 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 20530 16640 20536 16652
rect 19852 16612 20536 16640
rect 19852 16600 19858 16612
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 20898 16640 20904 16652
rect 20680 16612 20904 16640
rect 20680 16600 20686 16612
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 17221 16575 17279 16581
rect 16592 16544 17172 16572
rect 11756 16476 12204 16504
rect 11756 16464 11762 16476
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 14642 16504 14648 16516
rect 12400 16476 14648 16504
rect 12400 16464 12406 16476
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 15654 16464 15660 16516
rect 15712 16504 15718 16516
rect 16132 16513 16160 16544
rect 17144 16516 17172 16544
rect 17221 16541 17233 16575
rect 17267 16572 17279 16575
rect 18046 16572 18052 16584
rect 17267 16544 18052 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 18046 16532 18052 16544
rect 18104 16572 18110 16584
rect 21376 16572 21404 16680
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 21910 16640 21916 16652
rect 21600 16612 21916 16640
rect 21600 16600 21606 16612
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 22020 16649 22048 16680
rect 22741 16677 22753 16711
rect 22787 16708 22799 16711
rect 23477 16711 23535 16717
rect 22787 16680 23244 16708
rect 22787 16677 22799 16680
rect 22741 16671 22799 16677
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 22094 16600 22100 16652
rect 22152 16600 22158 16652
rect 22278 16600 22284 16652
rect 22336 16600 22342 16652
rect 22370 16600 22376 16652
rect 22428 16600 22434 16652
rect 22462 16600 22468 16652
rect 22520 16600 22526 16652
rect 22554 16600 22560 16652
rect 22612 16640 22618 16652
rect 22830 16640 22836 16652
rect 22612 16612 22836 16640
rect 22612 16600 22618 16612
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 23216 16649 23244 16680
rect 23477 16677 23489 16711
rect 23523 16708 23535 16711
rect 23750 16708 23756 16720
rect 23523 16680 23756 16708
rect 23523 16677 23535 16680
rect 23477 16671 23535 16677
rect 23750 16668 23756 16680
rect 23808 16668 23814 16720
rect 24302 16708 24308 16720
rect 23860 16680 24308 16708
rect 23860 16649 23888 16680
rect 24302 16668 24308 16680
rect 24360 16668 24366 16720
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16609 23259 16643
rect 23201 16603 23259 16609
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16640 23719 16643
rect 23845 16643 23903 16649
rect 23707 16612 23796 16640
rect 23707 16609 23719 16612
rect 23661 16603 23719 16609
rect 18104 16544 21404 16572
rect 18104 16532 18110 16544
rect 21726 16532 21732 16584
rect 21784 16572 21790 16584
rect 21784 16544 22876 16572
rect 21784 16532 21790 16544
rect 22848 16516 22876 16544
rect 22922 16532 22928 16584
rect 22980 16532 22986 16584
rect 23014 16532 23020 16584
rect 23072 16532 23078 16584
rect 23768 16572 23796 16612
rect 23845 16609 23857 16643
rect 23891 16609 23903 16643
rect 23845 16603 23903 16609
rect 23934 16600 23940 16652
rect 23992 16640 23998 16652
rect 24213 16643 24271 16649
rect 24213 16640 24225 16643
rect 23992 16612 24225 16640
rect 23992 16600 23998 16612
rect 24213 16609 24225 16612
rect 24259 16609 24271 16643
rect 24213 16603 24271 16609
rect 24486 16600 24492 16652
rect 24544 16600 24550 16652
rect 24780 16649 24808 16748
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 25041 16779 25099 16785
rect 25041 16776 25053 16779
rect 24912 16748 25053 16776
rect 24912 16736 24918 16748
rect 25041 16745 25053 16748
rect 25087 16776 25099 16779
rect 25774 16776 25780 16788
rect 25087 16748 25780 16776
rect 25087 16745 25099 16748
rect 25041 16739 25099 16745
rect 25774 16736 25780 16748
rect 25832 16736 25838 16788
rect 25866 16736 25872 16788
rect 25924 16736 25930 16788
rect 26786 16776 26792 16788
rect 26068 16748 26792 16776
rect 26068 16708 26096 16748
rect 26786 16736 26792 16748
rect 26844 16736 26850 16788
rect 26970 16736 26976 16788
rect 27028 16776 27034 16788
rect 27028 16748 27292 16776
rect 27028 16736 27034 16748
rect 27264 16717 27292 16748
rect 27798 16736 27804 16788
rect 27856 16736 27862 16788
rect 28718 16776 28724 16788
rect 27908 16748 28724 16776
rect 26697 16711 26755 16717
rect 24964 16680 26096 16708
rect 26142 16680 26648 16708
rect 24964 16652 24992 16680
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 24765 16643 24823 16649
rect 24765 16609 24777 16643
rect 24811 16609 24823 16643
rect 24765 16603 24823 16609
rect 24305 16575 24363 16581
rect 23768 16544 24256 16572
rect 24228 16516 24256 16544
rect 24305 16541 24317 16575
rect 24351 16572 24363 16575
rect 24394 16572 24400 16584
rect 24351 16544 24400 16572
rect 24351 16541 24363 16544
rect 24305 16535 24363 16541
rect 24394 16532 24400 16544
rect 24452 16532 24458 16584
rect 24688 16572 24716 16603
rect 24946 16600 24952 16652
rect 25004 16600 25010 16652
rect 25314 16600 25320 16652
rect 25372 16640 25378 16652
rect 25409 16643 25467 16649
rect 25409 16640 25421 16643
rect 25372 16612 25421 16640
rect 25372 16600 25378 16612
rect 25409 16609 25421 16612
rect 25455 16609 25467 16643
rect 25685 16643 25743 16649
rect 25685 16640 25697 16643
rect 25409 16603 25467 16609
rect 25516 16612 25697 16640
rect 25130 16572 25136 16584
rect 24688 16544 25136 16572
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 16117 16507 16175 16513
rect 16117 16504 16129 16507
rect 15712 16476 16129 16504
rect 15712 16464 15718 16476
rect 16117 16473 16129 16476
rect 16163 16473 16175 16507
rect 16117 16467 16175 16473
rect 17126 16464 17132 16516
rect 17184 16464 17190 16516
rect 17954 16464 17960 16516
rect 18012 16504 18018 16516
rect 18693 16507 18751 16513
rect 18693 16504 18705 16507
rect 18012 16476 18705 16504
rect 18012 16464 18018 16476
rect 18693 16473 18705 16476
rect 18739 16473 18751 16507
rect 18693 16467 18751 16473
rect 19794 16464 19800 16516
rect 19852 16504 19858 16516
rect 20622 16504 20628 16516
rect 19852 16476 20628 16504
rect 19852 16464 19858 16476
rect 20622 16464 20628 16476
rect 20680 16504 20686 16516
rect 22554 16504 22560 16516
rect 20680 16476 22560 16504
rect 20680 16464 20686 16476
rect 22554 16464 22560 16476
rect 22612 16464 22618 16516
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 23842 16504 23848 16516
rect 22888 16476 23848 16504
rect 22888 16464 22894 16476
rect 23842 16464 23848 16476
rect 23900 16504 23906 16516
rect 24029 16507 24087 16513
rect 24029 16504 24041 16507
rect 23900 16476 24041 16504
rect 23900 16464 23906 16476
rect 24029 16473 24041 16476
rect 24075 16473 24087 16507
rect 24029 16467 24087 16473
rect 24210 16464 24216 16516
rect 24268 16464 24274 16516
rect 24421 16476 24900 16504
rect 5040 16408 6776 16436
rect 5040 16396 5046 16408
rect 6822 16396 6828 16448
rect 6880 16436 6886 16448
rect 10226 16436 10232 16448
rect 6880 16408 10232 16436
rect 6880 16396 6886 16408
rect 10226 16396 10232 16408
rect 10284 16396 10290 16448
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11882 16436 11888 16448
rect 11112 16408 11888 16436
rect 11112 16396 11118 16408
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 14274 16436 14280 16448
rect 12032 16408 14280 16436
rect 12032 16396 12038 16408
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16301 16439 16359 16445
rect 16301 16436 16313 16439
rect 15988 16408 16313 16436
rect 15988 16396 15994 16408
rect 16301 16405 16313 16408
rect 16347 16405 16359 16439
rect 16301 16399 16359 16405
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 20898 16436 20904 16448
rect 16448 16408 20904 16436
rect 16448 16396 16454 16408
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 21085 16439 21143 16445
rect 21085 16405 21097 16439
rect 21131 16436 21143 16439
rect 21358 16436 21364 16448
rect 21131 16408 21364 16436
rect 21131 16405 21143 16408
rect 21085 16399 21143 16405
rect 21358 16396 21364 16408
rect 21416 16396 21422 16448
rect 22462 16396 22468 16448
rect 22520 16436 22526 16448
rect 23106 16436 23112 16448
rect 22520 16408 23112 16436
rect 22520 16396 22526 16408
rect 23106 16396 23112 16408
rect 23164 16436 23170 16448
rect 23382 16436 23388 16448
rect 23164 16408 23388 16436
rect 23164 16396 23170 16408
rect 23382 16396 23388 16408
rect 23440 16396 23446 16448
rect 23474 16396 23480 16448
rect 23532 16436 23538 16448
rect 24421 16436 24449 16476
rect 23532 16408 24449 16436
rect 24872 16436 24900 16476
rect 25516 16436 25544 16612
rect 25685 16609 25697 16612
rect 25731 16609 25743 16643
rect 25685 16603 25743 16609
rect 26053 16643 26111 16649
rect 26053 16609 26065 16643
rect 26099 16609 26111 16643
rect 26053 16603 26111 16609
rect 26068 16572 26096 16603
rect 25884 16544 26096 16572
rect 25590 16464 25596 16516
rect 25648 16504 25654 16516
rect 25884 16504 25912 16544
rect 26142 16504 26170 16680
rect 26237 16643 26295 16649
rect 26237 16609 26249 16643
rect 26283 16640 26295 16643
rect 26418 16640 26424 16652
rect 26283 16612 26424 16640
rect 26283 16609 26295 16612
rect 26237 16603 26295 16609
rect 26418 16600 26424 16612
rect 26476 16600 26482 16652
rect 26510 16600 26516 16652
rect 26568 16600 26574 16652
rect 26326 16532 26332 16584
rect 26384 16532 26390 16584
rect 26620 16572 26648 16680
rect 26697 16677 26709 16711
rect 26743 16708 26755 16711
rect 27249 16711 27307 16717
rect 26743 16680 27200 16708
rect 26743 16677 26755 16680
rect 26697 16671 26755 16677
rect 26786 16600 26792 16652
rect 26844 16600 26850 16652
rect 26973 16643 27031 16649
rect 26973 16609 26985 16643
rect 27019 16609 27031 16643
rect 27172 16640 27200 16680
rect 27249 16677 27261 16711
rect 27295 16677 27307 16711
rect 27249 16671 27307 16677
rect 27617 16711 27675 16717
rect 27617 16677 27629 16711
rect 27663 16708 27675 16711
rect 27908 16708 27936 16748
rect 28718 16736 28724 16748
rect 28776 16736 28782 16788
rect 28810 16736 28816 16788
rect 28868 16736 28874 16788
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 31018 16776 31024 16788
rect 28960 16748 31024 16776
rect 28960 16736 28966 16748
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 27663 16680 27936 16708
rect 27985 16711 28043 16717
rect 27663 16677 27675 16680
rect 27617 16671 27675 16677
rect 27985 16677 27997 16711
rect 28031 16708 28043 16711
rect 28074 16708 28080 16720
rect 28031 16680 28080 16708
rect 28031 16677 28043 16680
rect 27985 16671 28043 16677
rect 27632 16640 27660 16671
rect 28074 16668 28080 16680
rect 28132 16668 28138 16720
rect 29546 16708 29552 16720
rect 28828 16680 29552 16708
rect 28828 16662 28856 16680
rect 29546 16668 29552 16680
rect 29604 16668 29610 16720
rect 27172 16612 27660 16640
rect 27709 16643 27767 16649
rect 26973 16603 27031 16609
rect 27709 16609 27721 16643
rect 27755 16640 27767 16643
rect 28166 16640 28172 16652
rect 27755 16612 28172 16640
rect 27755 16609 27767 16612
rect 27709 16603 27767 16609
rect 26988 16572 27016 16603
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 28261 16643 28319 16649
rect 28261 16609 28273 16643
rect 28307 16640 28319 16643
rect 28350 16640 28356 16652
rect 28307 16612 28356 16640
rect 28307 16609 28319 16612
rect 28261 16603 28319 16609
rect 28350 16600 28356 16612
rect 28408 16600 28414 16652
rect 28736 16649 28856 16662
rect 28537 16643 28595 16649
rect 28537 16609 28549 16643
rect 28583 16609 28595 16643
rect 28537 16603 28595 16609
rect 28727 16643 28856 16649
rect 28727 16609 28739 16643
rect 28773 16634 28856 16643
rect 28905 16646 28963 16649
rect 28905 16643 28978 16646
rect 28773 16609 28785 16634
rect 28727 16603 28785 16609
rect 28905 16609 28917 16643
rect 28951 16609 28978 16643
rect 28905 16603 28978 16609
rect 29007 16643 29065 16649
rect 29007 16609 29019 16643
rect 29053 16609 29065 16643
rect 29007 16603 29065 16609
rect 26620 16544 27016 16572
rect 27154 16532 27160 16584
rect 27212 16572 27218 16584
rect 27798 16572 27804 16584
rect 27212 16544 27804 16572
rect 27212 16532 27218 16544
rect 27798 16532 27804 16544
rect 27856 16532 27862 16584
rect 27982 16532 27988 16584
rect 28040 16572 28046 16584
rect 28552 16572 28580 16603
rect 28950 16572 28978 16603
rect 28040 16544 28580 16572
rect 28644 16544 28978 16572
rect 28040 16532 28046 16544
rect 25648 16476 25912 16504
rect 26068 16476 26170 16504
rect 26344 16504 26372 16532
rect 26970 16504 26976 16516
rect 26344 16476 26976 16504
rect 25648 16464 25654 16476
rect 26068 16436 26096 16476
rect 26970 16464 26976 16476
rect 27028 16504 27034 16516
rect 28074 16504 28080 16516
rect 27028 16476 28080 16504
rect 27028 16464 27034 16476
rect 28074 16464 28080 16476
rect 28132 16464 28138 16516
rect 28644 16504 28672 16544
rect 29012 16516 29040 16603
rect 29730 16600 29736 16652
rect 29788 16600 29794 16652
rect 29917 16643 29975 16649
rect 29917 16609 29929 16643
rect 29963 16640 29975 16643
rect 29963 16612 29997 16640
rect 29963 16609 29975 16612
rect 29917 16603 29975 16609
rect 29273 16575 29331 16581
rect 29273 16541 29285 16575
rect 29319 16572 29331 16575
rect 29454 16572 29460 16584
rect 29319 16544 29460 16572
rect 29319 16541 29331 16544
rect 29273 16535 29331 16541
rect 29454 16532 29460 16544
rect 29512 16572 29518 16584
rect 29932 16572 29960 16603
rect 30282 16600 30288 16652
rect 30340 16640 30346 16652
rect 30377 16643 30435 16649
rect 30377 16640 30389 16643
rect 30340 16612 30389 16640
rect 30340 16600 30346 16612
rect 30377 16609 30389 16612
rect 30423 16609 30435 16643
rect 30377 16603 30435 16609
rect 30466 16600 30472 16652
rect 30524 16640 30530 16652
rect 30837 16643 30895 16649
rect 30837 16640 30849 16643
rect 30524 16612 30849 16640
rect 30524 16600 30530 16612
rect 30837 16609 30849 16612
rect 30883 16609 30895 16643
rect 30837 16603 30895 16609
rect 31110 16600 31116 16652
rect 31168 16600 31174 16652
rect 30006 16572 30012 16584
rect 29512 16544 30012 16572
rect 29512 16532 29518 16544
rect 30006 16532 30012 16544
rect 30064 16532 30070 16584
rect 28184 16476 28672 16504
rect 24872 16408 26096 16436
rect 26145 16439 26203 16445
rect 23532 16396 23538 16408
rect 26145 16405 26157 16439
rect 26191 16436 26203 16439
rect 26326 16436 26332 16448
rect 26191 16408 26332 16436
rect 26191 16405 26203 16408
rect 26145 16399 26203 16405
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 26786 16396 26792 16448
rect 26844 16436 26850 16448
rect 26881 16439 26939 16445
rect 26881 16436 26893 16439
rect 26844 16408 26893 16436
rect 26844 16396 26850 16408
rect 26881 16405 26893 16408
rect 26927 16405 26939 16439
rect 26881 16399 26939 16405
rect 27062 16396 27068 16448
rect 27120 16436 27126 16448
rect 27890 16436 27896 16448
rect 27120 16408 27896 16436
rect 27120 16396 27126 16408
rect 27890 16396 27896 16408
rect 27948 16436 27954 16448
rect 28184 16445 28212 16476
rect 28994 16464 29000 16516
rect 29052 16464 29058 16516
rect 31294 16504 31300 16516
rect 29656 16476 31300 16504
rect 28169 16439 28227 16445
rect 28169 16436 28181 16439
rect 27948 16408 28181 16436
rect 27948 16396 27954 16408
rect 28169 16405 28181 16408
rect 28215 16405 28227 16439
rect 28169 16399 28227 16405
rect 28442 16396 28448 16448
rect 28500 16436 28506 16448
rect 29178 16436 29184 16448
rect 28500 16408 29184 16436
rect 28500 16396 28506 16408
rect 29178 16396 29184 16408
rect 29236 16396 29242 16448
rect 29546 16396 29552 16448
rect 29604 16436 29610 16448
rect 29656 16445 29684 16476
rect 31294 16464 31300 16476
rect 31352 16464 31358 16516
rect 29641 16439 29699 16445
rect 29641 16436 29653 16439
rect 29604 16408 29653 16436
rect 29604 16396 29610 16408
rect 29641 16405 29653 16408
rect 29687 16405 29699 16439
rect 29641 16399 29699 16405
rect 31202 16396 31208 16448
rect 31260 16396 31266 16448
rect 552 16346 31648 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 11436 16346
rect 11488 16294 11500 16346
rect 11552 16294 11564 16346
rect 11616 16294 11628 16346
rect 11680 16294 11692 16346
rect 11744 16294 19210 16346
rect 19262 16294 19274 16346
rect 19326 16294 19338 16346
rect 19390 16294 19402 16346
rect 19454 16294 19466 16346
rect 19518 16294 26984 16346
rect 27036 16294 27048 16346
rect 27100 16294 27112 16346
rect 27164 16294 27176 16346
rect 27228 16294 27240 16346
rect 27292 16294 31648 16346
rect 552 16272 31648 16294
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 2406 16232 2412 16244
rect 2188 16204 2412 16232
rect 2188 16192 2194 16204
rect 2406 16192 2412 16204
rect 2464 16232 2470 16244
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2464 16204 2605 16232
rect 2464 16192 2470 16204
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 2593 16195 2651 16201
rect 3510 16192 3516 16244
rect 3568 16232 3574 16244
rect 3605 16235 3663 16241
rect 3605 16232 3617 16235
rect 3568 16204 3617 16232
rect 3568 16192 3574 16204
rect 3605 16201 3617 16204
rect 3651 16201 3663 16235
rect 3605 16195 3663 16201
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5258 16232 5264 16244
rect 5123 16204 5264 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6420 16204 6561 16232
rect 6420 16192 6426 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 6549 16195 6607 16201
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 10042 16232 10048 16244
rect 7156 16204 10048 16232
rect 7156 16192 7162 16204
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 10134 16192 10140 16244
rect 10192 16192 10198 16244
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 11388 16204 11529 16232
rect 11388 16192 11394 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 11517 16195 11575 16201
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 11882 16232 11888 16244
rect 11664 16204 11888 16232
rect 11664 16192 11670 16204
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 11992 16204 14136 16232
rect 566 16124 572 16176
rect 624 16164 630 16176
rect 1946 16164 1952 16176
rect 624 16136 1952 16164
rect 624 16124 630 16136
rect 1946 16124 1952 16136
rect 2004 16164 2010 16176
rect 2004 16136 2176 16164
rect 2004 16124 2010 16136
rect 1213 16099 1271 16105
rect 1213 16065 1225 16099
rect 1259 16096 1271 16099
rect 1765 16099 1823 16105
rect 1259 16068 1532 16096
rect 1259 16065 1271 16068
rect 1213 16059 1271 16065
rect 1504 16040 1532 16068
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 1811 16068 2085 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 1397 16031 1455 16037
rect 1397 16028 1409 16031
rect 1360 16000 1409 16028
rect 1360 15988 1366 16000
rect 1397 15997 1409 16000
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1412 15960 1440 15991
rect 1486 15988 1492 16040
rect 1544 16028 1550 16040
rect 1854 16028 1860 16040
rect 1544 16000 1860 16028
rect 1544 15988 1550 16000
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 15997 2007 16031
rect 1949 15991 2007 15997
rect 1964 15960 1992 15991
rect 1412 15932 1992 15960
rect 2057 15960 2085 16068
rect 2148 16037 2176 16136
rect 2222 16124 2228 16176
rect 2280 16164 2286 16176
rect 9033 16167 9091 16173
rect 2280 16136 8892 16164
rect 2280 16124 2286 16136
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 15997 2191 16031
rect 2133 15991 2191 15997
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 2314 16028 2320 16040
rect 2271 16000 2320 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2516 16037 2544 16136
rect 3510 16056 3516 16108
rect 3568 16096 3574 16108
rect 5261 16099 5319 16105
rect 3568 16068 5212 16096
rect 3568 16056 3574 16068
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 15997 2559 16031
rect 2501 15991 2559 15997
rect 2590 15988 2596 16040
rect 2648 16028 2654 16040
rect 2685 16031 2743 16037
rect 2685 16028 2697 16031
rect 2648 16000 2697 16028
rect 2648 15988 2654 16000
rect 2685 15997 2697 16000
rect 2731 15997 2743 16031
rect 2685 15991 2743 15997
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 3804 15960 3832 15991
rect 4246 15988 4252 16040
rect 4304 15988 4310 16040
rect 4982 15988 4988 16040
rect 5040 15988 5046 16040
rect 5184 16028 5212 16068
rect 5261 16065 5273 16099
rect 5307 16096 5319 16099
rect 6914 16096 6920 16108
rect 5307 16068 6920 16096
rect 5307 16065 5319 16068
rect 5261 16059 5319 16065
rect 5994 16028 6000 16040
rect 5184 16000 6000 16028
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 6472 16037 6500 16068
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7929 16099 7987 16105
rect 7064 16068 7880 16096
rect 7064 16056 7070 16068
rect 6457 16031 6515 16037
rect 6457 15997 6469 16031
rect 6503 15997 6515 16031
rect 6457 15991 6515 15997
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 7190 16028 7196 16040
rect 6687 16000 7196 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7852 16037 7880 16068
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8110 16096 8116 16108
rect 7975 16068 8116 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8110 16056 8116 16068
rect 8168 16096 8174 16108
rect 8168 16068 8800 16096
rect 8168 16056 8174 16068
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 5261 15963 5319 15969
rect 2057 15932 2636 15960
rect 3804 15932 3924 15960
rect 2608 15904 2636 15932
rect 1397 15895 1455 15901
rect 1397 15861 1409 15895
rect 1443 15892 1455 15895
rect 1486 15892 1492 15904
rect 1443 15864 1492 15892
rect 1443 15861 1455 15864
rect 1397 15855 1455 15861
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2222 15892 2228 15904
rect 1820 15864 2228 15892
rect 1820 15852 1826 15864
rect 2222 15852 2228 15864
rect 2280 15892 2286 15904
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 2280 15864 2421 15892
rect 2280 15852 2286 15864
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 2590 15852 2596 15904
rect 2648 15852 2654 15904
rect 3896 15892 3924 15932
rect 5261 15929 5273 15963
rect 5307 15960 5319 15963
rect 5626 15960 5632 15972
rect 5307 15932 5632 15960
rect 5307 15929 5319 15932
rect 5261 15923 5319 15929
rect 5626 15920 5632 15932
rect 5684 15960 5690 15972
rect 7760 15960 7788 15991
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 8202 16028 8208 16040
rect 8076 16000 8208 16028
rect 8076 15988 8082 16000
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8294 15988 8300 16040
rect 8352 16028 8358 16040
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 8352 16000 8401 16028
rect 8352 15988 8358 16000
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8481 16031 8539 16037
rect 8481 15997 8493 16031
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 5684 15932 7788 15960
rect 5684 15920 5690 15932
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 8496 15960 8524 15991
rect 7984 15932 8524 15960
rect 7984 15920 7990 15932
rect 8570 15920 8576 15972
rect 8628 15960 8634 15972
rect 8772 15969 8800 16068
rect 8864 16037 8892 16136
rect 9033 16133 9045 16167
rect 9079 16164 9091 16167
rect 11992 16164 12020 16204
rect 9079 16136 12020 16164
rect 9079 16133 9091 16136
rect 9033 16127 9091 16133
rect 12066 16124 12072 16176
rect 12124 16124 12130 16176
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 12434 16096 12440 16108
rect 9364 16068 11744 16096
rect 9364 16056 9370 16068
rect 11716 16040 11744 16068
rect 11992 16068 12440 16096
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 16028 8907 16031
rect 8938 16028 8944 16040
rect 8895 16000 8944 16028
rect 8895 15997 8907 16000
rect 8849 15991 8907 15997
rect 8938 15988 8944 16000
rect 8996 15988 9002 16040
rect 9416 16000 9996 16028
rect 8665 15963 8723 15969
rect 8665 15960 8677 15963
rect 8628 15932 8677 15960
rect 8628 15920 8634 15932
rect 8665 15929 8677 15932
rect 8711 15929 8723 15963
rect 8665 15923 8723 15929
rect 8757 15963 8815 15969
rect 8757 15929 8769 15963
rect 8803 15960 8815 15963
rect 9416 15960 9444 16000
rect 8803 15932 9444 15960
rect 8803 15929 8815 15932
rect 8757 15923 8815 15929
rect 9490 15920 9496 15972
rect 9548 15920 9554 15972
rect 9968 15960 9996 16000
rect 10042 15988 10048 16040
rect 10100 16028 10106 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 10100 16000 10333 16028
rect 10100 15988 10106 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 10597 16031 10655 16037
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 11330 16028 11336 16040
rect 10643 16000 11336 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 11882 15988 11888 16040
rect 11940 15988 11946 16040
rect 11992 16037 12020 16068
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 14108 16096 14136 16204
rect 14274 16192 14280 16244
rect 14332 16192 14338 16244
rect 14458 16192 14464 16244
rect 14516 16192 14522 16244
rect 15010 16192 15016 16244
rect 15068 16232 15074 16244
rect 19429 16235 19487 16241
rect 15068 16204 19334 16232
rect 15068 16192 15074 16204
rect 14292 16136 15792 16164
rect 14292 16096 14320 16136
rect 12912 16068 14044 16096
rect 14108 16068 14320 16096
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12250 16031 12308 16037
rect 12250 15997 12262 16031
rect 12296 16028 12308 16031
rect 12526 16028 12532 16040
rect 12296 16000 12532 16028
rect 12296 15997 12308 16000
rect 12250 15991 12308 15997
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12618 15988 12624 16040
rect 12676 15988 12682 16040
rect 9968 15932 10548 15960
rect 5534 15892 5540 15904
rect 3896 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 7466 15892 7472 15904
rect 6052 15864 7472 15892
rect 6052 15852 6058 15864
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 7650 15852 7656 15904
rect 7708 15892 7714 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7708 15864 8217 15892
rect 7708 15852 7714 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 9030 15852 9036 15904
rect 9088 15892 9094 15904
rect 9585 15895 9643 15901
rect 9585 15892 9597 15895
rect 9088 15864 9597 15892
rect 9088 15852 9094 15864
rect 9585 15861 9597 15864
rect 9631 15892 9643 15895
rect 10134 15892 10140 15904
rect 9631 15864 10140 15892
rect 9631 15861 9643 15864
rect 9585 15855 9643 15861
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10520 15901 10548 15932
rect 10870 15920 10876 15972
rect 10928 15960 10934 15972
rect 12066 15960 12072 15972
rect 10928 15932 12072 15960
rect 10928 15920 10934 15932
rect 12066 15920 12072 15932
rect 12124 15920 12130 15972
rect 12912 15960 12940 16068
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 14016 16028 14044 16068
rect 15654 16056 15660 16108
rect 15712 16056 15718 16108
rect 15764 16105 15792 16136
rect 16022 16124 16028 16176
rect 16080 16164 16086 16176
rect 19306 16164 19334 16204
rect 19429 16201 19441 16235
rect 19475 16232 19487 16235
rect 19794 16232 19800 16244
rect 19475 16204 19800 16232
rect 19475 16201 19487 16204
rect 19429 16195 19487 16201
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 19978 16192 19984 16244
rect 20036 16192 20042 16244
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 22094 16232 22100 16244
rect 20312 16204 22100 16232
rect 20312 16192 20318 16204
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22186 16192 22192 16244
rect 22244 16232 22250 16244
rect 22554 16232 22560 16244
rect 22244 16204 22560 16232
rect 22244 16192 22250 16204
rect 22554 16192 22560 16204
rect 22612 16232 22618 16244
rect 22925 16235 22983 16241
rect 22612 16204 22692 16232
rect 22612 16192 22618 16204
rect 22664 16173 22692 16204
rect 22925 16201 22937 16235
rect 22971 16232 22983 16235
rect 23014 16232 23020 16244
rect 22971 16204 23020 16232
rect 22971 16201 22983 16204
rect 22925 16195 22983 16201
rect 23014 16192 23020 16204
rect 23072 16192 23078 16244
rect 23109 16235 23167 16241
rect 23109 16201 23121 16235
rect 23155 16232 23167 16235
rect 23198 16232 23204 16244
rect 23155 16204 23204 16232
rect 23155 16201 23167 16204
rect 23109 16195 23167 16201
rect 23198 16192 23204 16204
rect 23256 16192 23262 16244
rect 23382 16192 23388 16244
rect 23440 16232 23446 16244
rect 25038 16232 25044 16244
rect 23440 16204 25044 16232
rect 23440 16192 23446 16204
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 26234 16192 26240 16244
rect 26292 16192 26298 16244
rect 26510 16192 26516 16244
rect 26568 16232 26574 16244
rect 28261 16235 28319 16241
rect 28261 16232 28273 16235
rect 26568 16204 28273 16232
rect 26568 16192 26574 16204
rect 28261 16201 28273 16204
rect 28307 16201 28319 16235
rect 28261 16195 28319 16201
rect 28718 16192 28724 16244
rect 28776 16232 28782 16244
rect 29365 16235 29423 16241
rect 29365 16232 29377 16235
rect 28776 16204 29377 16232
rect 28776 16192 28782 16204
rect 29365 16201 29377 16204
rect 29411 16201 29423 16235
rect 29365 16195 29423 16201
rect 29822 16192 29828 16244
rect 29880 16232 29886 16244
rect 30745 16235 30803 16241
rect 30745 16232 30757 16235
rect 29880 16204 30757 16232
rect 29880 16192 29886 16204
rect 30745 16201 30757 16204
rect 30791 16201 30803 16235
rect 30745 16195 30803 16201
rect 22649 16167 22707 16173
rect 16080 16136 18736 16164
rect 19306 16136 22600 16164
rect 16080 16124 16086 16136
rect 18708 16108 18736 16136
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 15988 16068 17908 16096
rect 15988 16056 15994 16068
rect 14016 16000 14228 16028
rect 13909 15991 13967 15997
rect 12268 15932 12940 15960
rect 10505 15895 10563 15901
rect 10505 15861 10517 15895
rect 10551 15892 10563 15895
rect 12158 15892 12164 15904
rect 10551 15864 12164 15892
rect 10551 15861 10563 15864
rect 10505 15855 10563 15861
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 12268 15901 12296 15932
rect 12986 15920 12992 15972
rect 13044 15920 13050 15972
rect 13630 15920 13636 15972
rect 13688 15960 13694 15972
rect 13924 15960 13952 15991
rect 13688 15932 13952 15960
rect 14200 15960 14228 16000
rect 14274 15988 14280 16040
rect 14332 15988 14338 16040
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 15381 16031 15439 16037
rect 15381 15997 15393 16031
rect 15427 16028 15439 16031
rect 16482 16028 16488 16040
rect 15427 16000 16488 16028
rect 15427 15997 15439 16000
rect 15381 15991 15439 15997
rect 15305 15960 15333 15991
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 17880 16028 17908 16068
rect 18690 16056 18696 16108
rect 18748 16096 18754 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18748 16068 19073 16096
rect 18748 16056 18754 16068
rect 19061 16065 19073 16068
rect 19107 16096 19119 16099
rect 19242 16096 19248 16108
rect 19107 16068 19248 16096
rect 19107 16065 19119 16068
rect 19061 16059 19119 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19852 16068 19901 16096
rect 19852 16056 19858 16068
rect 19889 16065 19901 16068
rect 19935 16065 19947 16099
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 19889 16059 19947 16065
rect 19996 16068 21097 16096
rect 19996 16037 20024 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 21821 16099 21879 16105
rect 21821 16096 21833 16099
rect 21315 16068 21833 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21821 16065 21833 16068
rect 21867 16065 21879 16099
rect 22462 16096 22468 16108
rect 21821 16059 21879 16065
rect 21928 16068 22468 16096
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 17880 16000 18889 16028
rect 18877 15997 18889 16000
rect 18923 16028 18935 16031
rect 19981 16031 20039 16037
rect 18923 16000 19840 16028
rect 18923 15997 18935 16000
rect 18877 15991 18935 15997
rect 16114 15960 16120 15972
rect 14200 15932 15148 15960
rect 15305 15932 16120 15960
rect 13688 15920 13694 15932
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12492 15864 12909 15892
rect 12492 15852 12498 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 13998 15892 14004 15904
rect 13872 15864 14004 15892
rect 13872 15852 13878 15864
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 15120 15901 15148 15932
rect 16114 15920 16120 15932
rect 16172 15960 16178 15972
rect 17034 15960 17040 15972
rect 16172 15932 17040 15960
rect 16172 15920 16178 15932
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 18598 15920 18604 15972
rect 18656 15960 18662 15972
rect 18693 15963 18751 15969
rect 18693 15960 18705 15963
rect 18656 15932 18705 15960
rect 18656 15920 18662 15932
rect 18693 15929 18705 15932
rect 18739 15929 18751 15963
rect 18693 15923 18751 15929
rect 19242 15920 19248 15972
rect 19300 15920 19306 15972
rect 19426 15920 19432 15972
rect 19484 15969 19490 15972
rect 19484 15963 19503 15969
rect 19491 15929 19503 15963
rect 19484 15923 19503 15929
rect 19705 15963 19763 15969
rect 19705 15929 19717 15963
rect 19751 15929 19763 15963
rect 19812 15960 19840 16000
rect 19981 15997 19993 16031
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 21361 16031 21419 16037
rect 21361 16028 21373 16031
rect 21232 16000 21373 16028
rect 21232 15988 21238 16000
rect 21361 15997 21373 16000
rect 21407 15997 21419 16031
rect 21361 15991 21419 15997
rect 21450 15988 21456 16040
rect 21508 15988 21514 16040
rect 21542 15988 21548 16040
rect 21600 15988 21606 16040
rect 21726 15988 21732 16040
rect 21784 15988 21790 16040
rect 21928 16037 21956 16068
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 21913 16031 21971 16037
rect 21913 15997 21925 16031
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 22278 15988 22284 16040
rect 22336 15988 22342 16040
rect 22002 15960 22008 15972
rect 19812 15932 22008 15960
rect 19705 15923 19763 15929
rect 19484 15920 19490 15923
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15861 15163 15895
rect 15105 15855 15163 15861
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 15436 15864 15485 15892
rect 15436 15852 15442 15864
rect 15473 15861 15485 15864
rect 15519 15861 15531 15895
rect 15473 15855 15531 15861
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 19334 15892 19340 15904
rect 15620 15864 19340 15892
rect 15620 15852 15626 15864
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 19720 15892 19748 15923
rect 22002 15920 22008 15932
rect 22060 15920 22066 15972
rect 22094 15920 22100 15972
rect 22152 15960 22158 15972
rect 22373 15963 22431 15969
rect 22373 15960 22385 15963
rect 22152 15932 22385 15960
rect 22152 15920 22158 15932
rect 22373 15929 22385 15932
rect 22419 15929 22431 15963
rect 22572 15960 22600 16136
rect 22649 16133 22661 16167
rect 22695 16133 22707 16167
rect 22649 16127 22707 16133
rect 23937 16167 23995 16173
rect 23937 16133 23949 16167
rect 23983 16133 23995 16167
rect 23937 16127 23995 16133
rect 24028 16136 25176 16164
rect 23014 16056 23020 16108
rect 23072 16096 23078 16108
rect 23566 16096 23572 16108
rect 23072 16068 23572 16096
rect 23072 16056 23078 16068
rect 23400 16037 23428 16068
rect 23566 16056 23572 16068
rect 23624 16096 23630 16108
rect 23952 16096 23980 16127
rect 23624 16068 23980 16096
rect 23624 16056 23630 16068
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 16028 23443 16031
rect 23431 16000 23465 16028
rect 23431 15997 23443 16000
rect 23385 15991 23443 15997
rect 23658 15988 23664 16040
rect 23716 15988 23722 16040
rect 23750 15988 23756 16040
rect 23808 16028 23814 16040
rect 24028 16028 24056 16136
rect 24302 16056 24308 16108
rect 24360 16056 24366 16108
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 24854 16096 24860 16108
rect 24719 16068 24860 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 25038 16056 25044 16108
rect 25096 16056 25102 16108
rect 25148 16105 25176 16136
rect 25682 16124 25688 16176
rect 25740 16164 25746 16176
rect 25777 16167 25835 16173
rect 25777 16164 25789 16167
rect 25740 16136 25789 16164
rect 25740 16124 25746 16136
rect 25777 16133 25789 16136
rect 25823 16164 25835 16167
rect 25866 16164 25872 16176
rect 25823 16136 25872 16164
rect 25823 16133 25835 16136
rect 25777 16127 25835 16133
rect 25866 16124 25872 16136
rect 25924 16124 25930 16176
rect 26878 16164 26884 16176
rect 25976 16136 26884 16164
rect 25976 16108 26004 16136
rect 26878 16124 26884 16136
rect 26936 16124 26942 16176
rect 27062 16124 27068 16176
rect 27120 16164 27126 16176
rect 27120 16136 27476 16164
rect 27120 16124 27126 16136
rect 25133 16099 25191 16105
rect 25133 16065 25145 16099
rect 25179 16096 25191 16099
rect 25958 16096 25964 16108
rect 25179 16068 25964 16096
rect 25179 16065 25191 16068
rect 25133 16059 25191 16065
rect 25958 16056 25964 16068
rect 26016 16056 26022 16108
rect 26418 16056 26424 16108
rect 26476 16056 26482 16108
rect 26694 16056 26700 16108
rect 26752 16096 26758 16108
rect 27154 16096 27160 16108
rect 26752 16068 27160 16096
rect 26752 16056 26758 16068
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27448 16096 27476 16136
rect 27522 16124 27528 16176
rect 27580 16164 27586 16176
rect 27614 16164 27620 16176
rect 27580 16136 27620 16164
rect 27580 16124 27586 16136
rect 27614 16124 27620 16136
rect 27672 16124 27678 16176
rect 27801 16167 27859 16173
rect 27801 16164 27813 16167
rect 27724 16136 27813 16164
rect 27724 16096 27752 16136
rect 27801 16133 27813 16136
rect 27847 16133 27859 16167
rect 27801 16127 27859 16133
rect 27982 16124 27988 16176
rect 28040 16164 28046 16176
rect 28040 16136 28856 16164
rect 28040 16124 28046 16136
rect 27448 16068 27752 16096
rect 27816 16068 28120 16096
rect 23808 16000 24056 16028
rect 23808 15988 23814 16000
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 24210 15988 24216 16040
rect 24268 16028 24274 16040
rect 24489 16031 24547 16037
rect 24489 16028 24501 16031
rect 24268 16000 24501 16028
rect 24268 15988 24274 16000
rect 24489 15997 24501 16000
rect 24535 15997 24547 16031
rect 24489 15991 24547 15997
rect 24578 15988 24584 16040
rect 24636 15988 24642 16040
rect 24762 15988 24768 16040
rect 24820 15988 24826 16040
rect 25056 16028 25084 16056
rect 25317 16031 25375 16037
rect 25317 16028 25329 16031
rect 25056 16000 25329 16028
rect 25317 15997 25329 16000
rect 25363 15997 25375 16031
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25317 15991 25375 15997
rect 25608 16000 25789 16028
rect 22922 15960 22928 15972
rect 22572 15932 22928 15960
rect 22373 15923 22431 15929
rect 22922 15920 22928 15932
rect 22980 15960 22986 15972
rect 23077 15963 23135 15969
rect 23077 15960 23089 15963
rect 22980 15932 23089 15960
rect 22980 15920 22986 15932
rect 23077 15929 23089 15932
rect 23123 15929 23135 15963
rect 23077 15923 23135 15929
rect 23293 15963 23351 15969
rect 23293 15929 23305 15963
rect 23339 15929 23351 15963
rect 23293 15923 23351 15929
rect 19659 15864 19748 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 20806 15852 20812 15904
rect 20864 15892 20870 15904
rect 21634 15892 21640 15904
rect 20864 15864 21640 15892
rect 20864 15852 20870 15864
rect 21634 15852 21640 15864
rect 21692 15852 21698 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 22833 15895 22891 15901
rect 22833 15892 22845 15895
rect 22612 15864 22845 15892
rect 22612 15852 22618 15864
rect 22833 15861 22845 15864
rect 22879 15892 22891 15895
rect 23198 15892 23204 15904
rect 22879 15864 23204 15892
rect 22879 15861 22891 15864
rect 22833 15855 22891 15861
rect 23198 15852 23204 15864
rect 23256 15852 23262 15904
rect 23308 15892 23336 15923
rect 23474 15892 23480 15904
rect 23308 15864 23480 15892
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 23566 15852 23572 15904
rect 23624 15852 23630 15904
rect 23676 15892 23704 15988
rect 23934 15920 23940 15972
rect 23992 15960 23998 15972
rect 25038 15960 25044 15972
rect 23992 15932 25044 15960
rect 23992 15920 23998 15932
rect 25038 15920 25044 15932
rect 25096 15960 25102 15972
rect 25608 15960 25636 16000
rect 25777 15997 25789 16000
rect 25823 16028 25835 16031
rect 26050 16028 26056 16040
rect 25823 16000 26056 16028
rect 25823 15997 25835 16000
rect 25777 15991 25835 15997
rect 26050 15988 26056 16000
rect 26108 15988 26114 16040
rect 26145 16031 26203 16037
rect 26145 15997 26157 16031
rect 26191 15997 26203 16031
rect 26145 15991 26203 15997
rect 25096 15932 25636 15960
rect 25096 15920 25102 15932
rect 25682 15920 25688 15972
rect 25740 15960 25746 15972
rect 26160 15960 26188 15991
rect 26326 15988 26332 16040
rect 26384 15988 26390 16040
rect 26436 16028 26464 16056
rect 27816 16040 27844 16068
rect 26789 16031 26847 16037
rect 26789 16028 26801 16031
rect 26436 16000 26801 16028
rect 26789 15997 26801 16000
rect 26835 15997 26847 16031
rect 26789 15991 26847 15997
rect 26878 15988 26884 16040
rect 26936 16028 26942 16040
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26936 16000 27261 16028
rect 26936 15988 26942 16000
rect 27249 15997 27261 16000
rect 27295 15997 27307 16031
rect 27249 15991 27307 15997
rect 27798 15988 27804 16040
rect 27856 15988 27862 16040
rect 28092 16037 28120 16068
rect 28258 16056 28264 16108
rect 28316 16056 28322 16108
rect 28828 16096 28856 16136
rect 29178 16124 29184 16176
rect 29236 16164 29242 16176
rect 29457 16167 29515 16173
rect 29457 16164 29469 16167
rect 29236 16136 29469 16164
rect 29236 16124 29242 16136
rect 29457 16133 29469 16136
rect 29503 16133 29515 16167
rect 29457 16127 29515 16133
rect 29546 16096 29552 16108
rect 28828 16068 29552 16096
rect 27985 16031 28043 16037
rect 27985 15997 27997 16031
rect 28031 15997 28043 16031
rect 27985 15991 28043 15997
rect 28077 16031 28135 16037
rect 28077 15997 28089 16031
rect 28123 15997 28135 16031
rect 28077 15991 28135 15997
rect 28000 15960 28028 15991
rect 28276 15960 28304 16056
rect 28626 15988 28632 16040
rect 28684 16037 28690 16040
rect 28828 16037 28856 16068
rect 29546 16056 29552 16068
rect 29604 16056 29610 16108
rect 28684 16031 28717 16037
rect 28705 15997 28717 16031
rect 28684 15991 28717 15997
rect 28813 16031 28871 16037
rect 28813 15997 28825 16031
rect 28859 15997 28871 16031
rect 28813 15991 28871 15997
rect 28684 15988 28690 15991
rect 28902 15988 28908 16040
rect 28960 16028 28966 16040
rect 28997 16031 29055 16037
rect 28997 16028 29009 16031
rect 28960 16000 29009 16028
rect 28960 15988 28966 16000
rect 28997 15997 29009 16000
rect 29043 15997 29055 16031
rect 28997 15991 29055 15997
rect 30374 15988 30380 16040
rect 30432 15988 30438 16040
rect 30926 15988 30932 16040
rect 30984 15988 30990 16040
rect 31110 15988 31116 16040
rect 31168 16028 31174 16040
rect 31386 16028 31392 16040
rect 31168 16000 31392 16028
rect 31168 15988 31174 16000
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 25740 15932 26188 15960
rect 26252 15932 27614 15960
rect 28000 15932 28304 15960
rect 28445 15963 28503 15969
rect 25740 15920 25746 15932
rect 26252 15892 26280 15932
rect 23676 15864 26280 15892
rect 26878 15852 26884 15904
rect 26936 15852 26942 15904
rect 27154 15852 27160 15904
rect 27212 15892 27218 15904
rect 27433 15895 27491 15901
rect 27433 15892 27445 15895
rect 27212 15864 27445 15892
rect 27212 15852 27218 15864
rect 27433 15861 27445 15864
rect 27479 15861 27491 15895
rect 27586 15892 27614 15932
rect 28445 15929 28457 15963
rect 28491 15929 28503 15963
rect 28445 15923 28503 15929
rect 28460 15892 28488 15923
rect 29454 15920 29460 15972
rect 29512 15960 29518 15972
rect 30190 15960 30196 15972
rect 29512 15932 30196 15960
rect 29512 15920 29518 15932
rect 30190 15920 30196 15932
rect 30248 15920 30254 15972
rect 27586 15864 28488 15892
rect 27433 15855 27491 15861
rect 28626 15852 28632 15904
rect 28684 15892 28690 15904
rect 29825 15895 29883 15901
rect 29825 15892 29837 15895
rect 28684 15864 29837 15892
rect 28684 15852 28690 15864
rect 29825 15861 29837 15864
rect 29871 15861 29883 15895
rect 29825 15855 29883 15861
rect 552 15802 31648 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 12096 15802
rect 12148 15750 12160 15802
rect 12212 15750 12224 15802
rect 12276 15750 12288 15802
rect 12340 15750 12352 15802
rect 12404 15750 19870 15802
rect 19922 15750 19934 15802
rect 19986 15750 19998 15802
rect 20050 15750 20062 15802
rect 20114 15750 20126 15802
rect 20178 15750 27644 15802
rect 27696 15750 27708 15802
rect 27760 15750 27772 15802
rect 27824 15750 27836 15802
rect 27888 15750 27900 15802
rect 27952 15750 31648 15802
rect 552 15728 31648 15750
rect 1578 15648 1584 15700
rect 1636 15648 1642 15700
rect 3421 15691 3479 15697
rect 3421 15657 3433 15691
rect 3467 15688 3479 15691
rect 4062 15688 4068 15700
rect 3467 15660 4068 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 5500 15660 6132 15688
rect 5500 15648 5506 15660
rect 4706 15620 4712 15632
rect 3344 15592 4712 15620
rect 1210 15512 1216 15564
rect 1268 15552 1274 15564
rect 1489 15555 1547 15561
rect 1489 15552 1501 15555
rect 1268 15524 1501 15552
rect 1268 15512 1274 15524
rect 1489 15521 1501 15524
rect 1535 15521 1547 15555
rect 1489 15515 1547 15521
rect 1578 15512 1584 15564
rect 1636 15552 1642 15564
rect 1673 15555 1731 15561
rect 1673 15552 1685 15555
rect 1636 15524 1685 15552
rect 1636 15512 1642 15524
rect 1673 15521 1685 15524
rect 1719 15521 1731 15555
rect 1673 15515 1731 15521
rect 3142 15512 3148 15564
rect 3200 15512 3206 15564
rect 3234 15512 3240 15564
rect 3292 15552 3298 15564
rect 3344 15561 3372 15592
rect 4706 15580 4712 15592
rect 4764 15580 4770 15632
rect 5537 15623 5595 15629
rect 5537 15589 5549 15623
rect 5583 15620 5595 15623
rect 5905 15623 5963 15629
rect 5905 15620 5917 15623
rect 5583 15592 5917 15620
rect 5583 15589 5595 15592
rect 5537 15583 5595 15589
rect 5905 15589 5917 15592
rect 5951 15589 5963 15623
rect 5905 15583 5963 15589
rect 3329 15555 3387 15561
rect 3329 15552 3341 15555
rect 3292 15524 3341 15552
rect 3292 15512 3298 15524
rect 3329 15521 3341 15524
rect 3375 15521 3387 15555
rect 3329 15515 3387 15521
rect 3418 15512 3424 15564
rect 3476 15552 3482 15564
rect 3789 15555 3847 15561
rect 3476 15524 3740 15552
rect 3476 15512 3482 15524
rect 2682 15444 2688 15496
rect 2740 15484 2746 15496
rect 3712 15493 3740 15524
rect 3789 15521 3801 15555
rect 3835 15552 3847 15555
rect 4062 15552 4068 15564
rect 3835 15524 4068 15552
rect 3835 15521 3847 15524
rect 3789 15515 3847 15521
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 3605 15487 3663 15493
rect 3605 15484 3617 15487
rect 2740 15456 3617 15484
rect 2740 15444 2746 15456
rect 3605 15453 3617 15456
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3697 15487 3755 15493
rect 3697 15453 3709 15487
rect 3743 15453 3755 15487
rect 3697 15447 3755 15453
rect 3881 15487 3939 15493
rect 3881 15453 3893 15487
rect 3927 15453 3939 15487
rect 3881 15447 3939 15453
rect 3145 15351 3203 15357
rect 3145 15317 3157 15351
rect 3191 15348 3203 15351
rect 3326 15348 3332 15360
rect 3191 15320 3332 15348
rect 3191 15317 3203 15320
rect 3145 15311 3203 15317
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 3712 15348 3740 15447
rect 3896 15416 3924 15447
rect 5074 15444 5080 15496
rect 5132 15484 5138 15496
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 5132 15456 5181 15484
rect 5132 15444 5138 15456
rect 5169 15453 5181 15456
rect 5215 15453 5227 15487
rect 5368 15484 5396 15515
rect 5626 15512 5632 15564
rect 5684 15512 5690 15564
rect 6104 15561 6132 15660
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 9582 15688 9588 15700
rect 7524 15660 9588 15688
rect 7524 15648 7530 15660
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10689 15691 10747 15697
rect 10689 15688 10701 15691
rect 10008 15660 10701 15688
rect 10008 15648 10014 15660
rect 10689 15657 10701 15660
rect 10735 15657 10747 15691
rect 10689 15651 10747 15657
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 11940 15660 12081 15688
rect 11940 15648 11946 15660
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12069 15651 12127 15657
rect 13538 15648 13544 15700
rect 13596 15648 13602 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 14001 15691 14059 15697
rect 14001 15688 14013 15691
rect 13872 15660 14013 15688
rect 13872 15648 13878 15660
rect 14001 15657 14013 15660
rect 14047 15657 14059 15691
rect 14001 15651 14059 15657
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15657 15691 15715 15697
rect 15657 15688 15669 15691
rect 15252 15660 15669 15688
rect 15252 15648 15258 15660
rect 15657 15657 15669 15660
rect 15703 15657 15715 15691
rect 15657 15651 15715 15657
rect 15746 15648 15752 15700
rect 15804 15688 15810 15700
rect 16301 15691 16359 15697
rect 16301 15688 16313 15691
rect 15804 15660 16313 15688
rect 15804 15648 15810 15660
rect 16301 15657 16313 15660
rect 16347 15657 16359 15691
rect 16301 15651 16359 15657
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 20162 15688 20168 15700
rect 16540 15660 20168 15688
rect 16540 15648 16546 15660
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 20806 15688 20812 15700
rect 20312 15660 20812 15688
rect 20312 15648 20318 15660
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 22646 15688 22652 15700
rect 20956 15660 22652 15688
rect 20956 15648 20962 15660
rect 22646 15648 22652 15660
rect 22704 15648 22710 15700
rect 22922 15648 22928 15700
rect 22980 15648 22986 15700
rect 24578 15688 24584 15700
rect 23400 15660 24584 15688
rect 7006 15620 7012 15632
rect 6288 15592 7012 15620
rect 6288 15561 6316 15592
rect 7006 15580 7012 15592
rect 7064 15620 7070 15632
rect 8021 15623 8079 15629
rect 8021 15620 8033 15623
rect 7064 15592 8033 15620
rect 7064 15580 7070 15592
rect 8021 15589 8033 15592
rect 8067 15589 8079 15623
rect 8021 15583 8079 15589
rect 8389 15623 8447 15629
rect 8389 15589 8401 15623
rect 8435 15620 8447 15623
rect 8478 15620 8484 15632
rect 8435 15592 8484 15620
rect 8435 15589 8447 15592
rect 8389 15583 8447 15589
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 9030 15580 9036 15632
rect 9088 15580 9094 15632
rect 10870 15620 10876 15632
rect 9324 15592 10876 15620
rect 6089 15555 6147 15561
rect 6089 15521 6101 15555
rect 6135 15521 6147 15555
rect 6089 15515 6147 15521
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15552 6423 15555
rect 6822 15552 6828 15564
rect 6411 15524 6828 15552
rect 6411 15521 6423 15524
rect 6365 15515 6423 15521
rect 5534 15484 5540 15496
rect 5368 15456 5540 15484
rect 5169 15447 5227 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 5994 15444 6000 15496
rect 6052 15484 6058 15496
rect 6288 15484 6316 15515
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 7466 15512 7472 15564
rect 7524 15512 7530 15564
rect 7650 15512 7656 15564
rect 7708 15512 7714 15564
rect 6052 15456 6316 15484
rect 6052 15444 6058 15456
rect 7558 15444 7564 15496
rect 7616 15444 7622 15496
rect 7742 15444 7748 15496
rect 7800 15444 7806 15496
rect 8938 15484 8944 15496
rect 7852 15456 8944 15484
rect 7852 15416 7880 15456
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9048 15493 9076 15580
rect 9324 15561 9352 15592
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 11974 15620 11980 15632
rect 11664 15592 11980 15620
rect 11664 15580 11670 15592
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 12434 15620 12440 15632
rect 12084 15592 12440 15620
rect 9309 15555 9367 15561
rect 9309 15521 9321 15555
rect 9355 15521 9367 15555
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9309 15515 9367 15521
rect 9508 15524 10057 15552
rect 9033 15487 9091 15493
rect 9033 15453 9045 15487
rect 9079 15453 9091 15487
rect 9033 15447 9091 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 3896 15388 7880 15416
rect 7929 15419 7987 15425
rect 7929 15385 7941 15419
rect 7975 15416 7987 15419
rect 9140 15416 9168 15447
rect 9214 15444 9220 15496
rect 9272 15444 9278 15496
rect 9508 15493 9536 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 10226 15512 10232 15564
rect 10284 15512 10290 15564
rect 10318 15512 10324 15564
rect 10376 15552 10382 15564
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 10376 15524 10517 15552
rect 10376 15512 10382 15524
rect 10505 15521 10517 15524
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 12084 15561 12112 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 13556 15620 13584 15648
rect 14461 15623 14519 15629
rect 13556 15592 13768 15620
rect 12069 15555 12127 15561
rect 12069 15552 12081 15555
rect 11296 15524 12081 15552
rect 11296 15512 11302 15524
rect 12069 15521 12081 15524
rect 12115 15521 12127 15555
rect 12069 15515 12127 15521
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15552 12311 15555
rect 12526 15552 12532 15564
rect 12299 15524 12532 15552
rect 12299 15521 12311 15524
rect 12253 15515 12311 15521
rect 12526 15512 12532 15524
rect 12584 15552 12590 15564
rect 12894 15552 12900 15564
rect 12584 15524 12900 15552
rect 12584 15512 12590 15524
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 13044 15524 13277 15552
rect 13044 15512 13050 15524
rect 13265 15521 13277 15524
rect 13311 15552 13323 15555
rect 13630 15552 13636 15564
rect 13311 15524 13636 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 13740 15561 13768 15592
rect 14461 15589 14473 15623
rect 14507 15620 14519 15623
rect 14550 15620 14556 15632
rect 14507 15592 14556 15620
rect 14507 15589 14519 15592
rect 14461 15583 14519 15589
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 14642 15580 14648 15632
rect 14700 15620 14706 15632
rect 14700 15592 14964 15620
rect 14700 15580 14706 15592
rect 13740 15555 13808 15561
rect 13740 15524 13762 15555
rect 13750 15521 13762 15524
rect 13796 15521 13808 15555
rect 13750 15515 13808 15521
rect 14826 15512 14832 15564
rect 14884 15512 14890 15564
rect 14936 15552 14964 15592
rect 15010 15580 15016 15632
rect 15068 15580 15074 15632
rect 15120 15592 17724 15620
rect 15120 15561 15148 15592
rect 15105 15555 15163 15561
rect 15105 15552 15117 15555
rect 14936 15524 15117 15552
rect 15105 15521 15117 15524
rect 15151 15521 15163 15555
rect 15105 15515 15163 15521
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15552 15255 15555
rect 15562 15552 15568 15564
rect 15243 15524 15568 15552
rect 15243 15521 15255 15524
rect 15197 15515 15255 15521
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 15654 15512 15660 15564
rect 15712 15512 15718 15564
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 15804 15524 15853 15552
rect 15804 15512 15810 15524
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 16623 15524 16896 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10778 15484 10784 15496
rect 10459 15456 10784 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 13078 15484 13084 15496
rect 10928 15456 13084 15484
rect 10928 15444 10934 15456
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 15672 15484 15700 15512
rect 16500 15484 16528 15515
rect 13587 15476 13814 15484
rect 13924 15476 15608 15484
rect 13587 15456 15608 15476
rect 15672 15456 16528 15484
rect 16669 15487 16727 15493
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 13786 15448 13952 15456
rect 7975 15388 9168 15416
rect 7975 15385 7987 15388
rect 7929 15379 7987 15385
rect 10318 15376 10324 15428
rect 10376 15376 10382 15428
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 11054 15416 11060 15428
rect 11020 15388 11060 15416
rect 11020 15376 11026 15388
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 15580 15416 15608 15456
rect 16669 15453 16681 15487
rect 16715 15453 16727 15487
rect 16669 15447 16727 15453
rect 16390 15416 16396 15428
rect 15580 15388 16396 15416
rect 16390 15376 16396 15388
rect 16448 15376 16454 15428
rect 16684 15416 16712 15447
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 16868 15484 16896 15524
rect 16942 15512 16948 15564
rect 17000 15512 17006 15564
rect 17696 15552 17724 15592
rect 17770 15580 17776 15632
rect 17828 15620 17834 15632
rect 18138 15620 18144 15632
rect 17828 15592 18144 15620
rect 17828 15580 17834 15592
rect 18138 15580 18144 15592
rect 18196 15620 18202 15632
rect 20714 15620 20720 15632
rect 18196 15592 20720 15620
rect 18196 15580 18202 15592
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 21361 15623 21419 15629
rect 21361 15620 21373 15623
rect 20916 15592 21373 15620
rect 17696 15524 17908 15552
rect 17310 15484 17316 15496
rect 16868 15456 17316 15484
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17736 15456 17785 15484
rect 17736 15444 17742 15456
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17880 15484 17908 15524
rect 17954 15512 17960 15564
rect 18012 15512 18018 15564
rect 18049 15555 18107 15561
rect 18049 15521 18061 15555
rect 18095 15552 18107 15555
rect 19518 15552 19524 15564
rect 18095 15524 19524 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 20070 15512 20076 15564
rect 20128 15552 20134 15564
rect 20916 15561 20944 15592
rect 21361 15589 21373 15592
rect 21407 15589 21419 15623
rect 21361 15583 21419 15589
rect 22370 15580 22376 15632
rect 22428 15620 22434 15632
rect 22465 15623 22523 15629
rect 22465 15620 22477 15623
rect 22428 15592 22477 15620
rect 22428 15580 22434 15592
rect 22465 15589 22477 15592
rect 22511 15589 22523 15623
rect 23400 15620 23428 15660
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 24673 15691 24731 15697
rect 24673 15657 24685 15691
rect 24719 15688 24731 15691
rect 24762 15688 24768 15700
rect 24719 15660 24768 15688
rect 24719 15657 24731 15660
rect 24673 15651 24731 15657
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 26510 15688 26516 15700
rect 25792 15660 26516 15688
rect 22465 15583 22523 15589
rect 22664 15592 23428 15620
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20128 15524 20913 15552
rect 20128 15512 20134 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 21174 15512 21180 15564
rect 21232 15552 21238 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 21232 15524 21281 15552
rect 21232 15512 21238 15524
rect 21269 15521 21281 15524
rect 21315 15521 21327 15555
rect 21269 15515 21327 15521
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15521 21511 15555
rect 22664 15552 22692 15592
rect 23474 15580 23480 15632
rect 23532 15620 23538 15632
rect 23532 15592 23704 15620
rect 23532 15580 23538 15592
rect 21453 15515 21511 15521
rect 22296 15524 22692 15552
rect 19702 15484 19708 15496
rect 17880 15456 19708 15484
rect 17773 15447 17831 15453
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20220 15456 21097 15484
rect 20220 15444 20226 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 21468 15484 21496 15515
rect 22296 15484 22324 15524
rect 23198 15512 23204 15564
rect 23256 15552 23262 15564
rect 23676 15561 23704 15592
rect 23750 15580 23756 15632
rect 23808 15580 23814 15632
rect 25792 15620 25820 15660
rect 26510 15648 26516 15660
rect 26568 15648 26574 15700
rect 27525 15691 27583 15697
rect 27525 15688 27537 15691
rect 27080 15660 27537 15688
rect 23860 15592 25820 15620
rect 25848 15623 25906 15629
rect 23569 15555 23627 15561
rect 23569 15552 23581 15555
rect 23256 15524 23581 15552
rect 23256 15512 23262 15524
rect 23569 15521 23581 15524
rect 23615 15521 23627 15555
rect 23569 15515 23627 15521
rect 23661 15555 23719 15561
rect 23661 15521 23673 15555
rect 23707 15521 23719 15555
rect 23661 15515 23719 15521
rect 21468 15456 22324 15484
rect 20717 15419 20775 15425
rect 20717 15416 20729 15419
rect 16684 15388 20729 15416
rect 20717 15385 20729 15388
rect 20763 15416 20775 15419
rect 20806 15416 20812 15428
rect 20763 15388 20812 15416
rect 20763 15385 20775 15388
rect 20717 15379 20775 15385
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 21468 15416 21496 15456
rect 23474 15444 23480 15496
rect 23532 15444 23538 15496
rect 23584 15484 23612 15515
rect 23860 15484 23888 15592
rect 25848 15589 25860 15623
rect 25894 15589 25906 15623
rect 25848 15583 25906 15589
rect 26053 15623 26111 15629
rect 26053 15589 26065 15623
rect 26099 15620 26111 15623
rect 26142 15620 26148 15632
rect 26099 15592 26148 15620
rect 26099 15589 26111 15592
rect 26053 15583 26111 15589
rect 23934 15512 23940 15564
rect 23992 15512 23998 15564
rect 24029 15555 24087 15561
rect 24029 15521 24041 15555
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 23584 15456 23888 15484
rect 20917 15388 21496 15416
rect 6546 15348 6552 15360
rect 3712 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 8018 15308 8024 15360
rect 8076 15348 8082 15360
rect 8846 15348 8852 15360
rect 8076 15320 8852 15348
rect 8076 15308 8082 15320
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 9582 15308 9588 15360
rect 9640 15348 9646 15360
rect 11606 15348 11612 15360
rect 9640 15320 11612 15348
rect 9640 15308 9646 15320
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 13354 15308 13360 15360
rect 13412 15348 13418 15360
rect 13449 15351 13507 15357
rect 13449 15348 13461 15351
rect 13412 15320 13461 15348
rect 13412 15308 13418 15320
rect 13449 15317 13461 15320
rect 13495 15317 13507 15351
rect 13449 15311 13507 15317
rect 13630 15308 13636 15360
rect 13688 15308 13694 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14185 15351 14243 15357
rect 14185 15348 14197 15351
rect 13872 15320 14197 15348
rect 13872 15308 13878 15320
rect 14185 15317 14197 15320
rect 14231 15317 14243 15351
rect 14185 15311 14243 15317
rect 15378 15308 15384 15360
rect 15436 15308 15442 15360
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 17770 15348 17776 15360
rect 15804 15320 17776 15348
rect 15804 15308 15810 15320
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 17862 15308 17868 15360
rect 17920 15308 17926 15360
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 20917 15348 20945 15388
rect 22830 15376 22836 15428
rect 22888 15376 22894 15428
rect 24044 15416 24072 15515
rect 24118 15512 24124 15564
rect 24176 15552 24182 15564
rect 24213 15555 24271 15561
rect 24213 15552 24225 15555
rect 24176 15524 24225 15552
rect 24176 15512 24182 15524
rect 24213 15521 24225 15524
rect 24259 15521 24271 15555
rect 24213 15515 24271 15521
rect 24305 15555 24363 15561
rect 24305 15521 24317 15555
rect 24351 15521 24363 15555
rect 24305 15515 24363 15521
rect 24320 15484 24348 15515
rect 24394 15512 24400 15564
rect 24452 15512 24458 15564
rect 24578 15512 24584 15564
rect 24636 15552 24642 15564
rect 25590 15552 25596 15564
rect 24636 15524 25596 15552
rect 24636 15512 24642 15524
rect 25590 15512 25596 15524
rect 25648 15552 25654 15564
rect 25863 15552 25891 15583
rect 26142 15580 26148 15592
rect 26200 15620 26206 15632
rect 26418 15620 26424 15632
rect 26200 15592 26424 15620
rect 26200 15580 26206 15592
rect 26418 15580 26424 15592
rect 26476 15580 26482 15632
rect 27080 15629 27108 15660
rect 27525 15657 27537 15660
rect 27571 15657 27583 15691
rect 27525 15651 27583 15657
rect 27614 15648 27620 15700
rect 27672 15688 27678 15700
rect 27672 15660 27752 15688
rect 27672 15648 27678 15660
rect 27065 15623 27123 15629
rect 27065 15589 27077 15623
rect 27111 15589 27123 15623
rect 27724 15620 27752 15660
rect 27890 15648 27896 15700
rect 27948 15688 27954 15700
rect 28074 15688 28080 15700
rect 27948 15660 28080 15688
rect 27948 15648 27954 15660
rect 28074 15648 28080 15660
rect 28132 15648 28138 15700
rect 28442 15648 28448 15700
rect 28500 15648 28506 15700
rect 29270 15688 29276 15700
rect 28552 15660 29276 15688
rect 28552 15629 28580 15660
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 29457 15691 29515 15697
rect 29457 15657 29469 15691
rect 29503 15688 29515 15691
rect 29546 15688 29552 15700
rect 29503 15660 29552 15688
rect 29503 15657 29515 15660
rect 29457 15651 29515 15657
rect 29546 15648 29552 15660
rect 29604 15688 29610 15700
rect 30098 15688 30104 15700
rect 29604 15660 30104 15688
rect 29604 15648 29610 15660
rect 30098 15648 30104 15660
rect 30156 15648 30162 15700
rect 30190 15648 30196 15700
rect 30248 15688 30254 15700
rect 30929 15691 30987 15697
rect 30929 15688 30941 15691
rect 30248 15660 30941 15688
rect 30248 15648 30254 15660
rect 30929 15657 30941 15660
rect 30975 15657 30987 15691
rect 30929 15651 30987 15657
rect 28537 15623 28595 15629
rect 27065 15583 27123 15589
rect 27356 15592 27660 15620
rect 27724 15592 27844 15620
rect 25648 15524 25891 15552
rect 25648 15512 25654 15524
rect 26326 15512 26332 15564
rect 26384 15552 26390 15564
rect 26973 15555 27031 15561
rect 26973 15552 26985 15555
rect 26384 15524 26985 15552
rect 26384 15512 26390 15524
rect 26973 15521 26985 15524
rect 27019 15521 27031 15555
rect 26973 15515 27031 15521
rect 27154 15512 27160 15564
rect 27212 15512 27218 15564
rect 27356 15561 27384 15592
rect 27632 15564 27660 15592
rect 27341 15555 27399 15561
rect 27341 15521 27353 15555
rect 27387 15521 27399 15555
rect 27341 15515 27399 15521
rect 27433 15555 27491 15561
rect 27433 15521 27445 15555
rect 27479 15521 27491 15555
rect 27433 15515 27491 15521
rect 24320 15456 24608 15484
rect 24580 15428 24608 15456
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24728 15456 24777 15484
rect 24728 15444 24734 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 25041 15487 25099 15493
rect 25041 15484 25053 15487
rect 24912 15456 25053 15484
rect 24912 15444 24918 15456
rect 25041 15453 25053 15456
rect 25087 15453 25099 15487
rect 25041 15447 25099 15453
rect 25314 15444 25320 15496
rect 25372 15484 25378 15496
rect 27448 15484 27476 15515
rect 27614 15512 27620 15564
rect 27672 15512 27678 15564
rect 27816 15561 27844 15592
rect 28000 15592 28488 15620
rect 28000 15561 28028 15592
rect 28460 15564 28488 15592
rect 28537 15589 28549 15623
rect 28583 15589 28595 15623
rect 31202 15620 31208 15632
rect 28537 15583 28595 15589
rect 29012 15592 31208 15620
rect 27709 15555 27767 15561
rect 27709 15521 27721 15555
rect 27755 15521 27767 15555
rect 27709 15515 27767 15521
rect 27801 15555 27859 15561
rect 27801 15521 27813 15555
rect 27847 15521 27859 15555
rect 27801 15515 27859 15521
rect 27985 15555 28043 15561
rect 27985 15521 27997 15555
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28077 15555 28135 15561
rect 28077 15521 28089 15555
rect 28123 15552 28135 15555
rect 28350 15552 28356 15564
rect 28123 15524 28356 15552
rect 28123 15521 28135 15524
rect 28077 15515 28135 15521
rect 25372 15456 27476 15484
rect 27724 15484 27752 15515
rect 28350 15512 28356 15524
rect 28408 15512 28414 15564
rect 28442 15512 28448 15564
rect 28500 15512 28506 15564
rect 29012 15561 29040 15592
rect 31202 15580 31208 15592
rect 31260 15580 31266 15632
rect 28997 15555 29055 15561
rect 28997 15521 29009 15555
rect 29043 15521 29055 15555
rect 28997 15515 29055 15521
rect 29178 15512 29184 15564
rect 29236 15552 29242 15564
rect 29273 15555 29331 15561
rect 29273 15552 29285 15555
rect 29236 15524 29285 15552
rect 29236 15512 29242 15524
rect 29273 15521 29285 15524
rect 29319 15521 29331 15555
rect 29273 15515 29331 15521
rect 29546 15512 29552 15564
rect 29604 15512 29610 15564
rect 29822 15512 29828 15564
rect 29880 15512 29886 15564
rect 30374 15512 30380 15564
rect 30432 15552 30438 15564
rect 30745 15555 30803 15561
rect 30745 15552 30757 15555
rect 30432 15524 30757 15552
rect 30432 15512 30438 15524
rect 30745 15521 30757 15524
rect 30791 15521 30803 15555
rect 30745 15515 30803 15521
rect 30834 15512 30840 15564
rect 30892 15552 30898 15564
rect 31113 15555 31171 15561
rect 31113 15552 31125 15555
rect 30892 15524 31125 15552
rect 30892 15512 30898 15524
rect 31113 15521 31125 15524
rect 31159 15521 31171 15555
rect 31113 15515 31171 15521
rect 31294 15512 31300 15564
rect 31352 15512 31358 15564
rect 28166 15484 28172 15496
rect 27724 15456 28172 15484
rect 25372 15444 25378 15456
rect 24044 15388 24532 15416
rect 19392 15320 20945 15348
rect 19392 15308 19398 15320
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 23842 15348 23848 15360
rect 21048 15320 23848 15348
rect 21048 15308 21054 15320
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 23937 15351 23995 15357
rect 23937 15317 23949 15351
rect 23983 15348 23995 15351
rect 24302 15348 24308 15360
rect 23983 15320 24308 15348
rect 23983 15317 23995 15320
rect 23937 15311 23995 15317
rect 24302 15308 24308 15320
rect 24360 15308 24366 15360
rect 24504 15348 24532 15388
rect 24578 15376 24584 15428
rect 24636 15416 24642 15428
rect 25685 15419 25743 15425
rect 25685 15416 25697 15419
rect 24636 15388 25697 15416
rect 24636 15376 24642 15388
rect 25685 15385 25697 15388
rect 25731 15385 25743 15419
rect 27448 15416 27476 15456
rect 28166 15444 28172 15456
rect 28224 15444 28230 15496
rect 28258 15444 28264 15496
rect 28316 15484 28322 15496
rect 28626 15484 28632 15496
rect 28316 15456 28632 15484
rect 28316 15444 28322 15456
rect 28626 15444 28632 15456
rect 28684 15444 28690 15496
rect 30006 15493 30012 15496
rect 29972 15487 30012 15493
rect 29972 15453 29984 15487
rect 29972 15447 30012 15453
rect 30006 15444 30012 15447
rect 30064 15444 30070 15496
rect 30193 15487 30251 15493
rect 30193 15453 30205 15487
rect 30239 15484 30251 15487
rect 31205 15487 31263 15493
rect 30239 15456 30328 15484
rect 30239 15453 30251 15456
rect 30193 15447 30251 15453
rect 28902 15416 28908 15428
rect 25685 15379 25743 15385
rect 25792 15388 27200 15416
rect 27448 15388 28908 15416
rect 24946 15348 24952 15360
rect 24504 15320 24952 15348
rect 24946 15308 24952 15320
rect 25004 15308 25010 15360
rect 25314 15308 25320 15360
rect 25372 15348 25378 15360
rect 25792 15348 25820 15388
rect 27172 15360 27200 15388
rect 28902 15376 28908 15388
rect 28960 15376 28966 15428
rect 29546 15376 29552 15428
rect 29604 15416 29610 15428
rect 30300 15416 30328 15456
rect 31205 15453 31217 15487
rect 31251 15484 31263 15487
rect 31662 15484 31668 15496
rect 31251 15456 31668 15484
rect 31251 15453 31263 15456
rect 31205 15447 31263 15453
rect 31662 15444 31668 15456
rect 31720 15444 31726 15496
rect 30466 15416 30472 15428
rect 29604 15388 30236 15416
rect 30300 15388 30472 15416
rect 29604 15376 29610 15388
rect 25372 15320 25820 15348
rect 25372 15308 25378 15320
rect 25866 15308 25872 15360
rect 25924 15308 25930 15360
rect 26694 15308 26700 15360
rect 26752 15348 26758 15360
rect 26789 15351 26847 15357
rect 26789 15348 26801 15351
rect 26752 15320 26801 15348
rect 26752 15308 26758 15320
rect 26789 15317 26801 15320
rect 26835 15317 26847 15351
rect 26789 15311 26847 15317
rect 27154 15308 27160 15360
rect 27212 15348 27218 15360
rect 28350 15348 28356 15360
rect 27212 15320 28356 15348
rect 27212 15308 27218 15320
rect 28350 15308 28356 15320
rect 28408 15308 28414 15360
rect 28813 15351 28871 15357
rect 28813 15317 28825 15351
rect 28859 15348 28871 15351
rect 28994 15348 29000 15360
rect 28859 15320 29000 15348
rect 28859 15317 28871 15320
rect 28813 15311 28871 15317
rect 28994 15308 29000 15320
rect 29052 15308 29058 15360
rect 29089 15351 29147 15357
rect 29089 15317 29101 15351
rect 29135 15348 29147 15351
rect 29270 15348 29276 15360
rect 29135 15320 29276 15348
rect 29135 15317 29147 15320
rect 29089 15311 29147 15317
rect 29270 15308 29276 15320
rect 29328 15308 29334 15360
rect 29730 15308 29736 15360
rect 29788 15348 29794 15360
rect 30101 15351 30159 15357
rect 30101 15348 30113 15351
rect 29788 15320 30113 15348
rect 29788 15308 29794 15320
rect 30101 15317 30113 15320
rect 30147 15317 30159 15351
rect 30208 15348 30236 15388
rect 30466 15376 30472 15388
rect 30524 15376 30530 15428
rect 30282 15348 30288 15360
rect 30208 15320 30288 15348
rect 30101 15311 30159 15317
rect 30282 15308 30288 15320
rect 30340 15308 30346 15360
rect 552 15258 31648 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 11436 15258
rect 11488 15206 11500 15258
rect 11552 15206 11564 15258
rect 11616 15206 11628 15258
rect 11680 15206 11692 15258
rect 11744 15206 19210 15258
rect 19262 15206 19274 15258
rect 19326 15206 19338 15258
rect 19390 15206 19402 15258
rect 19454 15206 19466 15258
rect 19518 15206 26984 15258
rect 27036 15206 27048 15258
rect 27100 15206 27112 15258
rect 27164 15206 27176 15258
rect 27228 15206 27240 15258
rect 27292 15206 31648 15258
rect 552 15184 31648 15206
rect 5261 15147 5319 15153
rect 5261 15113 5273 15147
rect 5307 15144 5319 15147
rect 5442 15144 5448 15156
rect 5307 15116 5448 15144
rect 5307 15113 5319 15116
rect 5261 15107 5319 15113
rect 5442 15104 5448 15116
rect 5500 15144 5506 15156
rect 6086 15144 6092 15156
rect 5500 15116 6092 15144
rect 5500 15104 5506 15116
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 6362 15104 6368 15156
rect 6420 15144 6426 15156
rect 7285 15147 7343 15153
rect 7285 15144 7297 15147
rect 6420 15116 7297 15144
rect 6420 15104 6426 15116
rect 7285 15113 7297 15116
rect 7331 15113 7343 15147
rect 7285 15107 7343 15113
rect 7469 15147 7527 15153
rect 7469 15113 7481 15147
rect 7515 15144 7527 15147
rect 7650 15144 7656 15156
rect 7515 15116 7656 15144
rect 7515 15113 7527 15116
rect 7469 15107 7527 15113
rect 3510 15036 3516 15088
rect 3568 15036 3574 15088
rect 3973 15079 4031 15085
rect 3973 15045 3985 15079
rect 4019 15076 4031 15079
rect 5629 15079 5687 15085
rect 5629 15076 5641 15079
rect 4019 15048 5641 15076
rect 4019 15045 4031 15048
rect 3973 15039 4031 15045
rect 5629 15045 5641 15048
rect 5675 15045 5687 15079
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 5629 15039 5687 15045
rect 5736 15048 6837 15076
rect 1210 14968 1216 15020
rect 1268 15008 1274 15020
rect 3528 15008 3556 15036
rect 1268 14980 3740 15008
rect 1268 14968 1274 14980
rect 1486 14900 1492 14952
rect 1544 14900 1550 14952
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 1719 14912 2176 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 1854 14804 1860 14816
rect 1627 14776 1860 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 2148 14804 2176 14912
rect 3326 14900 3332 14952
rect 3384 14900 3390 14952
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 3528 14872 3556 14903
rect 3602 14900 3608 14952
rect 3660 14900 3666 14952
rect 3712 14949 3740 14980
rect 5074 14968 5080 15020
rect 5132 14968 5138 15020
rect 5736 15008 5764 15048
rect 6825 15045 6837 15048
rect 6871 15045 6883 15079
rect 7300 15076 7328 15107
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 7760 15116 9536 15144
rect 7760 15076 7788 15116
rect 7300 15048 7788 15076
rect 6825 15039 6883 15045
rect 8018 15036 8024 15088
rect 8076 15036 8082 15088
rect 8570 15036 8576 15088
rect 8628 15076 8634 15088
rect 8628 15048 8984 15076
rect 8628 15036 8634 15048
rect 5184 14980 5764 15008
rect 3697 14943 3755 14949
rect 3697 14909 3709 14943
rect 3743 14909 3755 14943
rect 3697 14903 3755 14909
rect 4062 14900 4068 14952
rect 4120 14900 4126 14952
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 4157 14875 4215 14881
rect 4157 14872 4169 14875
rect 3528 14844 4169 14872
rect 4157 14841 4169 14844
rect 4203 14841 4215 14875
rect 4264 14872 4292 14903
rect 4890 14900 4896 14952
rect 4948 14900 4954 14952
rect 5184 14872 5212 14980
rect 5810 14968 5816 15020
rect 5868 14968 5874 15020
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7193 15011 7251 15017
rect 6972 14980 7144 15008
rect 6972 14968 6978 14980
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14909 5319 14943
rect 5261 14903 5319 14909
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 4264 14844 5212 14872
rect 4157 14835 4215 14841
rect 3970 14804 3976 14816
rect 2148 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5166 14804 5172 14816
rect 5031 14776 5172 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5276 14804 5304 14903
rect 5552 14872 5580 14903
rect 5718 14900 5724 14952
rect 5776 14940 5782 14952
rect 5905 14943 5963 14949
rect 5905 14940 5917 14943
rect 5776 14912 5917 14940
rect 5776 14900 5782 14912
rect 5905 14909 5917 14912
rect 5951 14909 5963 14943
rect 5905 14903 5963 14909
rect 6086 14900 6092 14952
rect 6144 14900 6150 14952
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7006 14940 7012 14952
rect 6880 14912 7012 14940
rect 6880 14900 6886 14912
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 5997 14875 6055 14881
rect 5997 14872 6009 14875
rect 5552 14844 6009 14872
rect 5997 14841 6009 14844
rect 6043 14841 6055 14875
rect 5997 14835 6055 14841
rect 5534 14804 5540 14816
rect 5276 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 6822 14804 6828 14816
rect 5859 14776 6828 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7116 14804 7144 14980
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7282 15008 7288 15020
rect 7239 14980 7288 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 8846 14968 8852 15020
rect 8904 14968 8910 15020
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 7282 14832 7288 14884
rect 7340 14872 7346 14884
rect 7392 14872 7420 14903
rect 7558 14900 7564 14952
rect 7616 14900 7622 14952
rect 8202 14900 8208 14952
rect 8260 14900 8266 14952
rect 8478 14900 8484 14952
rect 8536 14900 8542 14952
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 8956 14949 8984 15048
rect 9214 15036 9220 15088
rect 9272 15036 9278 15088
rect 9508 15076 9536 15116
rect 9582 15104 9588 15156
rect 9640 15104 9646 15156
rect 11885 15147 11943 15153
rect 9692 15116 11836 15144
rect 9692 15076 9720 15116
rect 9508 15048 9720 15076
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 11054 15076 11060 15088
rect 10284 15048 11060 15076
rect 10284 15036 10290 15048
rect 11054 15036 11060 15048
rect 11112 15076 11118 15088
rect 11238 15076 11244 15088
rect 11112 15048 11244 15076
rect 11112 15036 11118 15048
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11388 15048 11529 15076
rect 11388 15036 11394 15048
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 11808 15076 11836 15116
rect 11885 15113 11897 15147
rect 11931 15144 11943 15147
rect 14182 15144 14188 15156
rect 11931 15116 14188 15144
rect 11931 15113 11943 15116
rect 11885 15107 11943 15113
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 14274 15104 14280 15156
rect 14332 15144 14338 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14332 15116 14657 15144
rect 14332 15104 14338 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 14829 15147 14887 15153
rect 14829 15113 14841 15147
rect 14875 15113 14887 15147
rect 14829 15107 14887 15113
rect 11808 15048 13114 15076
rect 11517 15039 11575 15045
rect 9125 15011 9183 15017
rect 9125 14977 9137 15011
rect 9171 15008 9183 15011
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 9171 14980 9505 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 12986 15008 12992 15020
rect 10008 14980 12992 15008
rect 10008 14968 10014 14980
rect 12986 14968 12992 14980
rect 13044 14968 13050 15020
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8628 14912 8677 14940
rect 8628 14900 8634 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 8987 14912 9076 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 7340 14844 7420 14872
rect 8772 14872 8800 14903
rect 9048 14884 9076 14912
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9640 14912 9781 14940
rect 9640 14900 9646 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 10560 14912 11253 14940
rect 10560 14900 10566 14912
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 8846 14872 8852 14884
rect 8772 14844 8852 14872
rect 7340 14832 7346 14844
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 9030 14832 9036 14884
rect 9088 14832 9094 14884
rect 9950 14832 9956 14884
rect 10008 14872 10014 14884
rect 10870 14872 10876 14884
rect 10008 14844 10876 14872
rect 10008 14832 10014 14844
rect 10870 14832 10876 14844
rect 10928 14832 10934 14884
rect 11256 14872 11284 14903
rect 11422 14900 11428 14952
rect 11480 14900 11486 14952
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 11609 14943 11667 14949
rect 11609 14940 11621 14943
rect 11572 14912 11621 14940
rect 11572 14900 11578 14912
rect 11609 14909 11621 14912
rect 11655 14909 11667 14943
rect 11609 14903 11667 14909
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14940 11759 14943
rect 12066 14940 12072 14952
rect 11747 14912 12072 14940
rect 11747 14909 11759 14912
rect 11701 14903 11759 14909
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 12158 14900 12164 14952
rect 12216 14940 12222 14952
rect 12710 14940 12716 14952
rect 12216 14912 12716 14940
rect 12216 14900 12222 14912
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 12894 14872 12900 14884
rect 11256 14844 12900 14872
rect 12894 14832 12900 14844
rect 12952 14832 12958 14884
rect 13086 14872 13114 15048
rect 13262 15036 13268 15088
rect 13320 15076 13326 15088
rect 13320 15048 14320 15076
rect 13320 15036 13326 15048
rect 13446 14968 13452 15020
rect 13504 14968 13510 15020
rect 14292 15017 14320 15048
rect 14366 15036 14372 15088
rect 14424 15076 14430 15088
rect 14844 15076 14872 15107
rect 15010 15104 15016 15156
rect 15068 15144 15074 15156
rect 21174 15144 21180 15156
rect 15068 15116 21180 15144
rect 15068 15104 15074 15116
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 21634 15104 21640 15156
rect 21692 15144 21698 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21692 15116 21925 15144
rect 21692 15104 21698 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 21913 15107 21971 15113
rect 22738 15104 22744 15156
rect 22796 15144 22802 15156
rect 23750 15144 23756 15156
rect 22796 15116 23756 15144
rect 22796 15104 22802 15116
rect 23750 15104 23756 15116
rect 23808 15104 23814 15156
rect 24026 15104 24032 15156
rect 24084 15144 24090 15156
rect 25314 15144 25320 15156
rect 24084 15116 25320 15144
rect 24084 15104 24090 15116
rect 25314 15104 25320 15116
rect 25372 15104 25378 15156
rect 26050 15104 26056 15156
rect 26108 15144 26114 15156
rect 26108 15116 26464 15144
rect 26108 15104 26114 15116
rect 14424 15048 14872 15076
rect 14424 15036 14430 15048
rect 15194 15036 15200 15088
rect 15252 15076 15258 15088
rect 15252 15048 23244 15076
rect 15252 15036 15258 15048
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 15286 15008 15292 15020
rect 14700 14980 15292 15008
rect 14700 14968 14706 14980
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16206 15008 16212 15020
rect 15804 14980 16212 15008
rect 15804 14968 15810 14980
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16942 14968 16948 15020
rect 17000 15008 17006 15020
rect 17000 14980 17356 15008
rect 17000 14968 17006 14980
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13464 14940 13492 14968
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13320 14912 13553 14940
rect 13320 14900 13326 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13722 14900 13728 14952
rect 13780 14900 13786 14952
rect 13814 14900 13820 14952
rect 13872 14900 13878 14952
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 13924 14872 13952 14903
rect 14090 14900 14096 14952
rect 14148 14940 14154 14952
rect 14148 14912 15333 14940
rect 14148 14900 14154 14912
rect 14642 14872 14648 14884
rect 13086 14844 13676 14872
rect 13924 14844 14648 14872
rect 7650 14804 7656 14816
rect 7116 14776 7656 14804
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 13538 14804 13544 14816
rect 8168 14776 13544 14804
rect 8168 14764 8174 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 13648 14804 13676 14844
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 14813 14875 14871 14881
rect 14813 14841 14825 14875
rect 14859 14872 14871 14875
rect 14918 14872 14924 14884
rect 14859 14844 14924 14872
rect 14859 14841 14871 14844
rect 14813 14835 14871 14841
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 15013 14875 15071 14881
rect 15013 14841 15025 14875
rect 15059 14872 15071 14875
rect 15102 14872 15108 14884
rect 15059 14844 15108 14872
rect 15059 14841 15071 14844
rect 15013 14835 15071 14841
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15305 14872 15333 14912
rect 15654 14900 15660 14952
rect 15712 14940 15718 14952
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 15712 14912 17141 14940
rect 15712 14900 15718 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17218 14900 17224 14952
rect 17276 14900 17282 14952
rect 17328 14949 17356 14980
rect 17402 14968 17408 15020
rect 17460 15008 17466 15020
rect 17681 15011 17739 15017
rect 17681 15008 17693 15011
rect 17460 14980 17693 15008
rect 17460 14968 17466 14980
rect 17681 14977 17693 14980
rect 17727 14977 17739 15011
rect 17681 14971 17739 14977
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19392 14980 19717 15008
rect 19392 14968 19398 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20128 14980 20729 15008
rect 20128 14968 20134 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 15008 20867 15011
rect 21450 15008 21456 15020
rect 20855 14980 21456 15008
rect 20855 14977 20867 14980
rect 20809 14971 20867 14977
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 17497 14943 17555 14949
rect 17497 14909 17509 14943
rect 17543 14909 17555 14943
rect 17497 14903 17555 14909
rect 17512 14872 17540 14903
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 17773 14943 17831 14949
rect 17773 14940 17785 14943
rect 17644 14912 17785 14940
rect 17644 14900 17650 14912
rect 17773 14909 17785 14912
rect 17819 14909 17831 14943
rect 17773 14903 17831 14909
rect 17862 14900 17868 14952
rect 17920 14900 17926 14952
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14940 19855 14943
rect 20254 14940 20260 14952
rect 19843 14912 20260 14940
rect 19843 14909 19855 14912
rect 19797 14903 19855 14909
rect 20254 14900 20260 14912
rect 20312 14900 20318 14952
rect 20625 14943 20683 14949
rect 20625 14909 20637 14943
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 15305 14844 17356 14872
rect 17512 14844 19656 14872
rect 14182 14804 14188 14816
rect 13648 14776 14188 14804
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 14274 14764 14280 14816
rect 14332 14804 14338 14816
rect 16758 14804 16764 14816
rect 14332 14776 16764 14804
rect 14332 14764 14338 14776
rect 16758 14764 16764 14776
rect 16816 14764 16822 14816
rect 16853 14807 16911 14813
rect 16853 14773 16865 14807
rect 16899 14804 16911 14807
rect 17218 14804 17224 14816
rect 16899 14776 17224 14804
rect 16899 14773 16911 14776
rect 16853 14767 16911 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17328 14804 17356 14844
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 17328 14776 18153 14804
rect 18141 14773 18153 14776
rect 18187 14773 18199 14807
rect 18141 14767 18199 14773
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 19521 14807 19579 14813
rect 19521 14804 19533 14807
rect 19392 14776 19533 14804
rect 19392 14764 19398 14776
rect 19521 14773 19533 14776
rect 19567 14773 19579 14807
rect 19628 14804 19656 14844
rect 19886 14832 19892 14884
rect 19944 14872 19950 14884
rect 20162 14872 20168 14884
rect 19944 14844 20168 14872
rect 19944 14832 19950 14844
rect 20162 14832 20168 14844
rect 20220 14832 20226 14884
rect 20441 14807 20499 14813
rect 20441 14804 20453 14807
rect 19628 14776 20453 14804
rect 19521 14767 19579 14773
rect 20441 14773 20453 14776
rect 20487 14773 20499 14807
rect 20640 14804 20668 14903
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 20824 14872 20852 14971
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 21818 14968 21824 15020
rect 21876 15008 21882 15020
rect 21876 14980 22600 15008
rect 21876 14968 21882 14980
rect 20901 14943 20959 14949
rect 20901 14909 20913 14943
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 21361 14943 21419 14949
rect 21361 14909 21373 14943
rect 21407 14940 21419 14943
rect 21468 14940 21496 14968
rect 21407 14912 21496 14940
rect 21407 14909 21419 14912
rect 21361 14903 21419 14909
rect 20772 14844 20852 14872
rect 20916 14872 20944 14903
rect 21634 14900 21640 14952
rect 21692 14900 21698 14952
rect 21726 14900 21732 14952
rect 21784 14940 21790 14952
rect 22097 14943 22155 14949
rect 22097 14940 22109 14943
rect 21784 14912 22109 14940
rect 21784 14900 21790 14912
rect 22097 14909 22109 14912
rect 22143 14909 22155 14943
rect 22097 14903 22155 14909
rect 22370 14900 22376 14952
rect 22428 14940 22434 14952
rect 22572 14949 22600 14980
rect 22646 14968 22652 15020
rect 22704 15008 22710 15020
rect 22704 14980 23152 15008
rect 22704 14968 22710 14980
rect 23124 14952 23152 14980
rect 22465 14943 22523 14949
rect 22465 14940 22477 14943
rect 22428 14912 22477 14940
rect 22428 14900 22434 14912
rect 22465 14909 22477 14912
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14940 22615 14943
rect 22738 14940 22744 14952
rect 22603 14912 22744 14940
rect 22603 14909 22615 14912
rect 22557 14903 22615 14909
rect 22738 14900 22744 14912
rect 22796 14900 22802 14952
rect 23106 14900 23112 14952
rect 23164 14900 23170 14952
rect 21082 14872 21088 14884
rect 20916 14844 21088 14872
rect 20772 14832 20778 14844
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 21269 14875 21327 14881
rect 21269 14841 21281 14875
rect 21315 14872 21327 14875
rect 21450 14872 21456 14884
rect 21315 14844 21456 14872
rect 21315 14841 21327 14844
rect 21269 14835 21327 14841
rect 21450 14832 21456 14844
rect 21508 14832 21514 14884
rect 22186 14832 22192 14884
rect 22244 14832 22250 14884
rect 22281 14875 22339 14881
rect 22281 14841 22293 14875
rect 22327 14841 22339 14875
rect 22281 14835 22339 14841
rect 21634 14804 21640 14816
rect 20640 14776 21640 14804
rect 20441 14767 20499 14773
rect 21634 14764 21640 14776
rect 21692 14764 21698 14816
rect 21818 14764 21824 14816
rect 21876 14804 21882 14816
rect 22296 14804 22324 14835
rect 23014 14832 23020 14884
rect 23072 14832 23078 14884
rect 23216 14872 23244 15048
rect 23566 15036 23572 15088
rect 23624 15076 23630 15088
rect 24673 15079 24731 15085
rect 24673 15076 24685 15079
rect 23624 15048 24685 15076
rect 23624 15036 23630 15048
rect 24673 15045 24685 15048
rect 24719 15045 24731 15079
rect 24673 15039 24731 15045
rect 24946 14968 24952 15020
rect 25004 14968 25010 15020
rect 25130 14968 25136 15020
rect 25188 15008 25194 15020
rect 26326 15008 26332 15020
rect 25188 14980 26332 15008
rect 25188 14968 25194 14980
rect 23382 14900 23388 14952
rect 23440 14900 23446 14952
rect 24302 14900 24308 14952
rect 24360 14900 24366 14952
rect 24486 14900 24492 14952
rect 24544 14900 24550 14952
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24765 14943 24823 14949
rect 24765 14909 24777 14943
rect 24811 14940 24823 14943
rect 24964 14940 24992 14968
rect 24811 14912 24992 14940
rect 24811 14909 24823 14912
rect 24765 14903 24823 14909
rect 24854 14872 24860 14884
rect 23216 14844 24860 14872
rect 24854 14832 24860 14844
rect 24912 14832 24918 14884
rect 24964 14872 24992 14912
rect 25130 14872 25136 14884
rect 24964 14844 25136 14872
rect 25130 14832 25136 14844
rect 25188 14832 25194 14884
rect 25501 14875 25559 14881
rect 25501 14841 25513 14875
rect 25547 14872 25559 14875
rect 25590 14872 25596 14884
rect 25547 14844 25596 14872
rect 25547 14841 25559 14844
rect 25501 14835 25559 14841
rect 25590 14832 25596 14844
rect 25648 14832 25654 14884
rect 25700 14881 25728 14980
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 25685 14875 25743 14881
rect 25685 14841 25697 14875
rect 25731 14841 25743 14875
rect 26053 14875 26111 14881
rect 25685 14835 25743 14841
rect 25792 14844 26004 14872
rect 22462 14804 22468 14816
rect 21876 14776 22468 14804
rect 21876 14764 21882 14776
rect 22462 14764 22468 14776
rect 22520 14804 22526 14816
rect 23934 14804 23940 14816
rect 22520 14776 23940 14804
rect 22520 14764 22526 14776
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 24949 14807 25007 14813
rect 24949 14773 24961 14807
rect 24995 14804 25007 14807
rect 25314 14804 25320 14816
rect 24995 14776 25320 14804
rect 24995 14773 25007 14776
rect 24949 14767 25007 14773
rect 25314 14764 25320 14776
rect 25372 14764 25378 14816
rect 25406 14764 25412 14816
rect 25464 14804 25470 14816
rect 25792 14813 25820 14844
rect 25777 14807 25835 14813
rect 25777 14804 25789 14807
rect 25464 14776 25789 14804
rect 25464 14764 25470 14776
rect 25777 14773 25789 14776
rect 25823 14773 25835 14807
rect 25777 14767 25835 14773
rect 25866 14764 25872 14816
rect 25924 14764 25930 14816
rect 25976 14804 26004 14844
rect 26053 14841 26065 14875
rect 26099 14872 26111 14875
rect 26436 14872 26464 15116
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 28997 15147 29055 15153
rect 28997 15144 29009 15147
rect 27672 15116 29009 15144
rect 27672 15104 27678 15116
rect 28997 15113 29009 15116
rect 29043 15113 29055 15147
rect 28997 15107 29055 15113
rect 29362 15104 29368 15156
rect 29420 15144 29426 15156
rect 29457 15147 29515 15153
rect 29457 15144 29469 15147
rect 29420 15116 29469 15144
rect 29420 15104 29426 15116
rect 29457 15113 29469 15116
rect 29503 15113 29515 15147
rect 29457 15107 29515 15113
rect 29917 15147 29975 15153
rect 29917 15113 29929 15147
rect 29963 15144 29975 15147
rect 30926 15144 30932 15156
rect 29963 15116 30932 15144
rect 29963 15113 29975 15116
rect 29917 15107 29975 15113
rect 27430 15036 27436 15088
rect 27488 15076 27494 15088
rect 27985 15079 28043 15085
rect 27985 15076 27997 15079
rect 27488 15048 27997 15076
rect 27488 15036 27494 15048
rect 27985 15045 27997 15048
rect 28031 15045 28043 15079
rect 27985 15039 28043 15045
rect 28442 15036 28448 15088
rect 28500 15076 28506 15088
rect 29932 15076 29960 15107
rect 30926 15104 30932 15116
rect 30984 15104 30990 15156
rect 31021 15147 31079 15153
rect 31021 15113 31033 15147
rect 31067 15144 31079 15147
rect 31754 15144 31760 15156
rect 31067 15116 31760 15144
rect 31067 15113 31079 15116
rect 31021 15107 31079 15113
rect 31754 15104 31760 15116
rect 31812 15104 31818 15156
rect 28500 15048 29960 15076
rect 28500 15036 28506 15048
rect 30282 15036 30288 15088
rect 30340 15076 30346 15088
rect 30340 15048 30880 15076
rect 30340 15036 30346 15048
rect 28534 15008 28540 15020
rect 27908 14980 28540 15008
rect 26513 14943 26571 14949
rect 26513 14909 26525 14943
rect 26559 14940 26571 14943
rect 27338 14940 27344 14952
rect 26559 14912 27344 14940
rect 26559 14909 26571 14912
rect 26513 14903 26571 14909
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 27908 14949 27936 14980
rect 28534 14968 28540 14980
rect 28592 15008 28598 15020
rect 28592 14980 29500 15008
rect 28592 14968 28598 14980
rect 27893 14943 27951 14949
rect 27893 14909 27905 14943
rect 27939 14909 27951 14943
rect 27893 14903 27951 14909
rect 28077 14943 28135 14949
rect 28077 14909 28089 14943
rect 28123 14909 28135 14943
rect 28077 14903 28135 14909
rect 26099 14844 26464 14872
rect 26099 14841 26111 14844
rect 26053 14835 26111 14841
rect 26142 14804 26148 14816
rect 25976 14776 26148 14804
rect 26142 14764 26148 14776
rect 26200 14764 26206 14816
rect 26234 14764 26240 14816
rect 26292 14764 26298 14816
rect 27338 14764 27344 14816
rect 27396 14804 27402 14816
rect 27706 14804 27712 14816
rect 27396 14776 27712 14804
rect 27396 14764 27402 14776
rect 27706 14764 27712 14776
rect 27764 14764 27770 14816
rect 28092 14804 28120 14903
rect 28166 14900 28172 14952
rect 28224 14940 28230 14952
rect 29270 14940 29276 14952
rect 28224 14912 29276 14940
rect 28224 14900 28230 14912
rect 29270 14900 29276 14912
rect 29328 14900 29334 14952
rect 29472 14949 29500 14980
rect 29546 14968 29552 15020
rect 29604 15008 29610 15020
rect 29604 14980 30236 15008
rect 29604 14968 29610 14980
rect 29457 14943 29515 14949
rect 29457 14909 29469 14943
rect 29503 14909 29515 14943
rect 29457 14903 29515 14909
rect 29733 14943 29791 14949
rect 29733 14909 29745 14943
rect 29779 14940 29791 14943
rect 29914 14940 29920 14952
rect 29779 14912 29920 14940
rect 29779 14909 29791 14912
rect 29733 14903 29791 14909
rect 29914 14900 29920 14912
rect 29972 14900 29978 14952
rect 30208 14949 30236 14980
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14909 30251 14943
rect 30193 14903 30251 14909
rect 30374 14900 30380 14952
rect 30432 14940 30438 14952
rect 30432 14912 30512 14940
rect 30432 14900 30438 14912
rect 28350 14832 28356 14884
rect 28408 14872 28414 14884
rect 28997 14875 29055 14881
rect 28997 14872 29009 14875
rect 28408 14844 29009 14872
rect 28408 14832 28414 14844
rect 28997 14841 29009 14844
rect 29043 14841 29055 14875
rect 29549 14875 29607 14881
rect 29549 14872 29561 14875
rect 28997 14835 29055 14841
rect 29104 14844 29561 14872
rect 29104 14804 29132 14844
rect 29549 14841 29561 14844
rect 29595 14872 29607 14875
rect 29638 14872 29644 14884
rect 29595 14844 29644 14872
rect 29595 14841 29607 14844
rect 29549 14835 29607 14841
rect 29638 14832 29644 14844
rect 29696 14832 29702 14884
rect 30009 14875 30067 14881
rect 30009 14872 30021 14875
rect 29932 14844 30021 14872
rect 29932 14816 29960 14844
rect 30009 14841 30021 14844
rect 30055 14841 30067 14875
rect 30009 14835 30067 14841
rect 28092 14776 29132 14804
rect 29178 14764 29184 14816
rect 29236 14764 29242 14816
rect 29914 14764 29920 14816
rect 29972 14764 29978 14816
rect 30374 14764 30380 14816
rect 30432 14764 30438 14816
rect 30484 14804 30512 14912
rect 30558 14900 30564 14952
rect 30616 14900 30622 14952
rect 30852 14949 30880 15048
rect 30837 14943 30895 14949
rect 30837 14909 30849 14943
rect 30883 14940 30895 14943
rect 31570 14940 31576 14952
rect 30883 14912 31576 14940
rect 30883 14909 30895 14912
rect 30837 14903 30895 14909
rect 31570 14900 31576 14912
rect 31628 14900 31634 14952
rect 30745 14807 30803 14813
rect 30745 14804 30757 14807
rect 30484 14776 30757 14804
rect 30745 14773 30757 14776
rect 30791 14773 30803 14807
rect 30745 14767 30803 14773
rect 552 14714 31648 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 12096 14714
rect 12148 14662 12160 14714
rect 12212 14662 12224 14714
rect 12276 14662 12288 14714
rect 12340 14662 12352 14714
rect 12404 14662 19870 14714
rect 19922 14662 19934 14714
rect 19986 14662 19998 14714
rect 20050 14662 20062 14714
rect 20114 14662 20126 14714
rect 20178 14662 27644 14714
rect 27696 14662 27708 14714
rect 27760 14662 27772 14714
rect 27824 14662 27836 14714
rect 27888 14662 27900 14714
rect 27952 14662 31648 14714
rect 552 14640 31648 14662
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 6365 14603 6423 14609
rect 3292 14572 3464 14600
rect 3292 14560 3298 14572
rect 1688 14504 2774 14532
rect 1688 14473 1716 14504
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14433 1731 14467
rect 1673 14427 1731 14433
rect 1854 14424 1860 14476
rect 1912 14424 1918 14476
rect 1946 14424 1952 14476
rect 2004 14424 2010 14476
rect 2222 14424 2228 14476
rect 2280 14424 2286 14476
rect 2746 14464 2774 14504
rect 3142 14492 3148 14544
rect 3200 14492 3206 14544
rect 2866 14464 2872 14476
rect 2746 14436 2872 14464
rect 2866 14424 2872 14436
rect 2924 14464 2930 14476
rect 3234 14464 3240 14476
rect 2924 14436 3240 14464
rect 2924 14424 2930 14436
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 3436 14473 3464 14572
rect 6365 14569 6377 14603
rect 6411 14569 6423 14603
rect 6365 14563 6423 14569
rect 5350 14532 5356 14544
rect 5184 14504 5356 14532
rect 3421 14467 3479 14473
rect 3421 14433 3433 14467
rect 3467 14464 3479 14467
rect 4154 14464 4160 14476
rect 3467 14436 4160 14464
rect 3467 14433 3479 14436
rect 3421 14427 3479 14433
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 5184 14473 5212 14504
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 5994 14492 6000 14544
rect 6052 14492 6058 14544
rect 6380 14532 6408 14563
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 7006 14600 7012 14612
rect 6604 14572 7012 14600
rect 6604 14560 6610 14572
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7282 14609 7288 14612
rect 7278 14563 7288 14609
rect 7282 14560 7288 14563
rect 7340 14560 7346 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7432 14572 8708 14600
rect 7432 14560 7438 14572
rect 8110 14532 8116 14544
rect 6380 14504 8116 14532
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 8680 14532 8708 14572
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 8812 14572 9168 14600
rect 8812 14560 8818 14572
rect 8938 14532 8944 14544
rect 8680 14504 8944 14532
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 5442 14424 5448 14476
rect 5500 14424 5506 14476
rect 5718 14464 5724 14476
rect 5552 14436 5724 14464
rect 2041 14399 2099 14405
rect 2041 14365 2053 14399
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14396 3387 14399
rect 4062 14396 4068 14408
rect 3375 14368 4068 14396
rect 3375 14365 3387 14368
rect 3329 14359 3387 14365
rect 1026 14288 1032 14340
rect 1084 14328 1090 14340
rect 2056 14328 2084 14359
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 1084 14300 2084 14328
rect 1084 14288 1090 14300
rect 3234 14288 3240 14340
rect 3292 14328 3298 14340
rect 3418 14328 3424 14340
rect 3292 14300 3424 14328
rect 3292 14288 3298 14300
rect 3418 14288 3424 14300
rect 3476 14288 3482 14340
rect 3605 14331 3663 14337
rect 3605 14297 3617 14331
rect 3651 14328 3663 14331
rect 5276 14328 5304 14359
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5552 14396 5580 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 6012 14464 6040 14492
rect 6012 14436 6868 14464
rect 5408 14368 5580 14396
rect 5629 14399 5687 14405
rect 5408 14356 5414 14368
rect 5629 14365 5641 14399
rect 5675 14396 5687 14399
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 5675 14368 5917 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 5905 14365 5917 14368
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 3651 14300 5304 14328
rect 3651 14297 3663 14300
rect 3605 14291 3663 14297
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 6012 14328 6040 14359
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6178 14356 6184 14408
rect 6236 14356 6242 14408
rect 6840 14396 6868 14436
rect 6914 14424 6920 14476
rect 6972 14424 6978 14476
rect 7098 14424 7104 14476
rect 7156 14424 7162 14476
rect 7193 14467 7251 14473
rect 7193 14433 7205 14467
rect 7239 14433 7251 14467
rect 7193 14427 7251 14433
rect 7208 14396 7236 14427
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7340 14436 7389 14464
rect 7340 14424 7346 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 7466 14424 7472 14476
rect 7524 14464 7530 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 7524 14436 7573 14464
rect 7524 14424 7530 14436
rect 7561 14433 7573 14436
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 6840 14368 7236 14396
rect 7760 14396 7788 14427
rect 8570 14424 8576 14476
rect 8628 14464 8634 14476
rect 8665 14467 8723 14473
rect 8665 14464 8677 14467
rect 8628 14436 8677 14464
rect 8628 14424 8634 14436
rect 8665 14433 8677 14436
rect 8711 14464 8723 14467
rect 8754 14464 8760 14476
rect 8711 14436 8760 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 8864 14473 8892 14504
rect 8938 14492 8944 14504
rect 8996 14492 9002 14544
rect 9140 14541 9168 14572
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9272 14572 9321 14600
rect 9272 14560 9278 14572
rect 9309 14569 9321 14572
rect 9355 14600 9367 14603
rect 10226 14600 10232 14612
rect 9355 14572 10232 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10778 14560 10784 14612
rect 10836 14560 10842 14612
rect 13722 14600 13728 14612
rect 11072 14572 13728 14600
rect 9125 14535 9183 14541
rect 9125 14501 9137 14535
rect 9171 14501 9183 14535
rect 9582 14532 9588 14544
rect 9125 14495 9183 14501
rect 9324 14504 9588 14532
rect 8849 14467 8907 14473
rect 8849 14433 8861 14467
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9324 14464 9352 14504
rect 9582 14492 9588 14504
rect 9640 14492 9646 14544
rect 10502 14492 10508 14544
rect 10560 14532 10566 14544
rect 10796 14532 10824 14560
rect 10560 14504 11008 14532
rect 10560 14492 10566 14504
rect 9088 14436 9352 14464
rect 9401 14467 9459 14473
rect 9088 14424 9094 14436
rect 9401 14433 9413 14467
rect 9447 14464 9459 14467
rect 10410 14464 10416 14476
rect 9447 14436 10416 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 8110 14396 8116 14408
rect 7760 14368 8116 14396
rect 6932 14340 6960 14368
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 9416 14396 9444 14427
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 10594 14424 10600 14476
rect 10652 14424 10658 14476
rect 10778 14424 10784 14476
rect 10836 14424 10842 14476
rect 10980 14473 11008 14504
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 8772 14368 9444 14396
rect 6822 14328 6828 14340
rect 5592 14300 6828 14328
rect 5592 14288 5598 14300
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 6914 14288 6920 14340
rect 6972 14288 6978 14340
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 7745 14331 7803 14337
rect 7745 14328 7757 14331
rect 7432 14300 7757 14328
rect 7432 14288 7438 14300
rect 7745 14297 7757 14300
rect 7791 14328 7803 14331
rect 8772 14328 8800 14368
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 11072 14396 11100 14572
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 14001 14603 14059 14609
rect 14001 14600 14013 14603
rect 13964 14572 14013 14600
rect 13964 14560 13970 14572
rect 14001 14569 14013 14572
rect 14047 14569 14059 14603
rect 14001 14563 14059 14569
rect 14826 14560 14832 14612
rect 14884 14560 14890 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 16117 14603 16175 14609
rect 16117 14600 16129 14603
rect 15344 14572 16129 14600
rect 15344 14560 15350 14572
rect 16117 14569 16129 14572
rect 16163 14569 16175 14603
rect 16117 14563 16175 14569
rect 16390 14560 16396 14612
rect 16448 14600 16454 14612
rect 17770 14600 17776 14612
rect 16448 14572 17776 14600
rect 16448 14560 16454 14572
rect 17770 14560 17776 14572
rect 17828 14560 17834 14612
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 18049 14603 18107 14609
rect 18049 14600 18061 14603
rect 17920 14572 18061 14600
rect 17920 14560 17926 14572
rect 18049 14569 18061 14572
rect 18095 14569 18107 14603
rect 18049 14563 18107 14569
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 19426 14600 19432 14612
rect 18288 14572 19432 14600
rect 18288 14560 18294 14572
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 19702 14560 19708 14612
rect 19760 14600 19766 14612
rect 19978 14600 19984 14612
rect 19760 14572 19984 14600
rect 19760 14560 19766 14572
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 22186 14600 22192 14612
rect 20864 14572 22192 14600
rect 20864 14560 20870 14572
rect 22186 14560 22192 14572
rect 22244 14560 22250 14612
rect 22462 14560 22468 14612
rect 22520 14560 22526 14612
rect 22925 14603 22983 14609
rect 22925 14569 22937 14603
rect 22971 14569 22983 14603
rect 25958 14600 25964 14612
rect 22925 14563 22983 14569
rect 23492 14572 25964 14600
rect 12805 14535 12863 14541
rect 11716 14504 12020 14532
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14464 11483 14467
rect 11606 14464 11612 14476
rect 11471 14436 11612 14464
rect 11471 14433 11483 14436
rect 11425 14427 11483 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 11716 14473 11744 14504
rect 11701 14467 11759 14473
rect 11701 14433 11713 14467
rect 11747 14433 11759 14467
rect 11701 14427 11759 14433
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14433 11943 14467
rect 11992 14462 12020 14504
rect 12805 14501 12817 14535
rect 12851 14532 12863 14535
rect 14274 14532 14280 14544
rect 12851 14504 14280 14532
rect 12851 14501 12863 14504
rect 12805 14495 12863 14501
rect 14274 14492 14280 14504
rect 14332 14492 14338 14544
rect 14642 14492 14648 14544
rect 14700 14532 14706 14544
rect 15197 14535 15255 14541
rect 14700 14504 15148 14532
rect 14700 14492 14706 14504
rect 12066 14462 12072 14476
rect 11992 14434 12072 14462
rect 11885 14427 11943 14433
rect 9640 14368 11100 14396
rect 9640 14356 9646 14368
rect 11146 14356 11152 14408
rect 11204 14356 11210 14408
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 7791 14300 8800 14328
rect 7791 14297 7803 14300
rect 7745 14291 7803 14297
rect 9030 14288 9036 14340
rect 9088 14288 9094 14340
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9490 14328 9496 14340
rect 9171 14300 9496 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 10781 14331 10839 14337
rect 10781 14297 10793 14331
rect 10827 14328 10839 14331
rect 11348 14328 11376 14359
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 11793 14399 11851 14405
rect 11572 14388 11652 14396
rect 11793 14388 11805 14399
rect 11572 14368 11805 14388
rect 11572 14356 11578 14368
rect 11624 14365 11805 14368
rect 11839 14365 11851 14399
rect 11900 14396 11928 14427
rect 12066 14424 12072 14434
rect 12124 14424 12130 14476
rect 12618 14464 12624 14476
rect 12176 14436 12624 14464
rect 11900 14388 12020 14396
rect 12176 14388 12204 14436
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 13081 14467 13139 14473
rect 12759 14436 13032 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 11900 14368 12204 14388
rect 11624 14360 11851 14365
rect 11992 14360 12204 14368
rect 11793 14359 11851 14360
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 12308 14368 12560 14396
rect 12308 14356 12314 14368
rect 12434 14328 12440 14340
rect 10827 14300 11376 14328
rect 11532 14300 12440 14328
rect 10827 14297 10839 14300
rect 10781 14291 10839 14297
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 3145 14263 3203 14269
rect 3145 14260 3157 14263
rect 2455 14232 3157 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 3145 14229 3157 14232
rect 3191 14229 3203 14263
rect 3145 14223 3203 14229
rect 3970 14220 3976 14272
rect 4028 14260 4034 14272
rect 5718 14260 5724 14272
rect 4028 14232 5724 14260
rect 4028 14220 4034 14232
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 6454 14220 6460 14272
rect 6512 14260 6518 14272
rect 6641 14263 6699 14269
rect 6641 14260 6653 14263
rect 6512 14232 6653 14260
rect 6512 14220 6518 14232
rect 6641 14229 6653 14232
rect 6687 14229 6699 14263
rect 6641 14223 6699 14229
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 8386 14260 8392 14272
rect 7524 14232 8392 14260
rect 7524 14220 7530 14232
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 11532 14260 11560 14300
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 12532 14328 12560 14368
rect 12894 14356 12900 14408
rect 12952 14356 12958 14408
rect 13004 14396 13032 14436
rect 13081 14433 13093 14467
rect 13127 14464 13139 14467
rect 13262 14464 13268 14476
rect 13127 14436 13268 14464
rect 13127 14433 13139 14436
rect 13081 14427 13139 14433
rect 13262 14424 13268 14436
rect 13320 14464 13326 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 13320 14436 13369 14464
rect 13320 14424 13326 14436
rect 13357 14433 13369 14436
rect 13403 14433 13415 14467
rect 13357 14427 13415 14433
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14433 13691 14467
rect 13633 14427 13691 14433
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14464 13783 14467
rect 14090 14464 14096 14476
rect 13771 14436 14096 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 13648 14396 13676 14427
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14464 14795 14467
rect 14918 14464 14924 14476
rect 14783 14436 14924 14464
rect 14783 14433 14795 14436
rect 14737 14427 14795 14433
rect 14918 14424 14924 14436
rect 14976 14424 14982 14476
rect 15010 14424 15016 14476
rect 15068 14424 15074 14476
rect 15120 14464 15148 14504
rect 15197 14501 15209 14535
rect 15243 14532 15255 14535
rect 17126 14532 17132 14544
rect 15243 14504 15516 14532
rect 15243 14501 15255 14504
rect 15197 14495 15255 14501
rect 15488 14473 15516 14504
rect 15580 14504 17132 14532
rect 15580 14473 15608 14504
rect 17126 14492 17132 14504
rect 17184 14492 17190 14544
rect 22940 14532 22968 14563
rect 18524 14504 22968 14532
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 15120 14436 15301 14464
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15473 14467 15531 14473
rect 15473 14433 15485 14467
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 15654 14424 15660 14476
rect 15712 14424 15718 14476
rect 16298 14424 16304 14476
rect 16356 14424 16362 14476
rect 16574 14424 16580 14476
rect 16632 14424 16638 14476
rect 16758 14424 16764 14476
rect 16816 14424 16822 14476
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 17000 14436 18245 14464
rect 17000 14424 17006 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18233 14427 18291 14433
rect 18414 14424 18420 14476
rect 18472 14424 18478 14476
rect 18524 14473 18552 14504
rect 18509 14467 18567 14473
rect 18509 14433 18521 14467
rect 18555 14433 18567 14467
rect 18509 14427 18567 14433
rect 19010 14436 19472 14464
rect 16206 14396 16212 14408
rect 13004 14368 13584 14396
rect 13648 14368 16212 14396
rect 12802 14328 12808 14340
rect 12532 14300 12808 14328
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 13078 14288 13084 14340
rect 13136 14288 13142 14340
rect 13556 14328 13584 14368
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 19010 14396 19038 14436
rect 19444 14408 19472 14436
rect 19518 14424 19524 14476
rect 19576 14424 19582 14476
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 17552 14368 19038 14396
rect 17552 14356 17558 14368
rect 19334 14356 19340 14408
rect 19392 14356 19398 14408
rect 19426 14356 19432 14408
rect 19484 14356 19490 14408
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14396 19855 14399
rect 19904 14396 19932 14427
rect 19978 14424 19984 14476
rect 20036 14424 20042 14476
rect 22833 14467 22891 14473
rect 22572 14464 22784 14467
rect 22833 14464 22845 14467
rect 20640 14439 22845 14464
rect 20640 14436 22600 14439
rect 22756 14436 22845 14439
rect 20165 14399 20223 14405
rect 20165 14396 20177 14399
rect 19843 14368 19932 14396
rect 19996 14368 20177 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 15933 14331 15991 14337
rect 13556 14300 15884 14328
rect 8720 14232 11560 14260
rect 11609 14263 11667 14269
rect 8720 14220 8726 14232
rect 11609 14229 11621 14263
rect 11655 14260 11667 14263
rect 15654 14260 15660 14272
rect 11655 14232 15660 14260
rect 11655 14229 11667 14232
rect 11609 14223 11667 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 15856 14260 15884 14300
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16393 14331 16451 14337
rect 16393 14328 16405 14331
rect 15979 14300 16405 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16393 14297 16405 14300
rect 16439 14297 16451 14331
rect 16393 14291 16451 14297
rect 16485 14331 16543 14337
rect 16485 14297 16497 14331
rect 16531 14328 16543 14331
rect 16574 14328 16580 14340
rect 16531 14300 16580 14328
rect 16531 14297 16543 14300
rect 16485 14291 16543 14297
rect 16574 14288 16580 14300
rect 16632 14288 16638 14340
rect 16850 14288 16856 14340
rect 16908 14328 16914 14340
rect 16908 14300 17632 14328
rect 16908 14288 16914 14300
rect 17494 14260 17500 14272
rect 15856 14232 17500 14260
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 17604 14260 17632 14300
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19628 14328 19656 14359
rect 19886 14328 19892 14340
rect 19208 14300 19892 14328
rect 19208 14288 19214 14300
rect 19886 14288 19892 14300
rect 19944 14288 19950 14340
rect 19996 14260 20024 14368
rect 20165 14365 20177 14368
rect 20211 14365 20223 14399
rect 20165 14359 20223 14365
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20530 14396 20536 14408
rect 20404 14368 20536 14396
rect 20404 14356 20410 14368
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 20073 14331 20131 14337
rect 20073 14297 20085 14331
rect 20119 14328 20131 14331
rect 20640 14328 20668 14436
rect 22833 14433 22845 14436
rect 22879 14433 22891 14467
rect 22833 14427 22891 14433
rect 23014 14424 23020 14476
rect 23072 14464 23078 14476
rect 23492 14473 23520 14572
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 26418 14560 26424 14612
rect 26476 14600 26482 14612
rect 26476 14572 28396 14600
rect 26476 14560 26482 14572
rect 23584 14504 24164 14532
rect 23109 14467 23167 14473
rect 23109 14464 23121 14467
rect 23072 14436 23121 14464
rect 23072 14424 23078 14436
rect 23109 14433 23121 14436
rect 23155 14433 23167 14467
rect 23109 14427 23167 14433
rect 23477 14467 23535 14473
rect 23477 14433 23489 14467
rect 23523 14433 23535 14467
rect 23477 14427 23535 14433
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 20119 14300 20668 14328
rect 20119 14297 20131 14300
rect 20073 14291 20131 14297
rect 21174 14288 21180 14340
rect 21232 14328 21238 14340
rect 22278 14328 22284 14340
rect 21232 14300 22284 14328
rect 21232 14288 21238 14300
rect 22278 14288 22284 14300
rect 22336 14288 22342 14340
rect 22756 14328 22784 14359
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 23584 14396 23612 14504
rect 23658 14424 23664 14476
rect 23716 14464 23722 14476
rect 23845 14467 23903 14473
rect 23845 14464 23857 14467
rect 23716 14436 23857 14464
rect 23716 14424 23722 14436
rect 23845 14433 23857 14436
rect 23891 14433 23903 14467
rect 23845 14427 23903 14433
rect 24026 14424 24032 14476
rect 24084 14424 24090 14476
rect 24136 14473 24164 14504
rect 24210 14492 24216 14544
rect 24268 14532 24274 14544
rect 24268 14504 25268 14532
rect 24268 14492 24274 14504
rect 24121 14467 24179 14473
rect 24121 14433 24133 14467
rect 24167 14433 24179 14467
rect 24121 14427 24179 14433
rect 24302 14424 24308 14476
rect 24360 14424 24366 14476
rect 24397 14467 24455 14473
rect 24397 14433 24409 14467
rect 24443 14433 24455 14467
rect 24397 14427 24455 14433
rect 24489 14467 24547 14473
rect 24489 14433 24501 14467
rect 24535 14464 24547 14467
rect 24578 14464 24584 14476
rect 24535 14436 24584 14464
rect 24535 14433 24547 14436
rect 24489 14427 24547 14433
rect 23256 14368 23612 14396
rect 23937 14399 23995 14405
rect 23256 14356 23262 14368
rect 23937 14365 23949 14399
rect 23983 14396 23995 14399
rect 24412 14396 24440 14427
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 25240 14464 25268 14504
rect 25314 14492 25320 14544
rect 25372 14492 25378 14544
rect 27065 14535 27123 14541
rect 27065 14532 27077 14535
rect 25608 14504 27077 14532
rect 25608 14464 25636 14504
rect 27065 14501 27077 14504
rect 27111 14501 27123 14535
rect 28077 14535 28135 14541
rect 28077 14532 28089 14535
rect 27065 14495 27123 14501
rect 27172 14504 28089 14532
rect 25240 14436 25636 14464
rect 25685 14467 25743 14473
rect 25685 14433 25697 14467
rect 25731 14433 25743 14467
rect 25685 14427 25743 14433
rect 25869 14467 25927 14473
rect 25869 14433 25881 14467
rect 25915 14464 25927 14467
rect 25958 14464 25964 14476
rect 25915 14436 25964 14464
rect 25915 14433 25927 14436
rect 25869 14427 25927 14433
rect 25590 14396 25596 14408
rect 23983 14368 24440 14396
rect 24872 14368 25596 14396
rect 23983 14365 23995 14368
rect 23937 14359 23995 14365
rect 24872 14328 24900 14368
rect 25590 14356 25596 14368
rect 25648 14356 25654 14408
rect 25700 14396 25728 14427
rect 25958 14424 25964 14436
rect 26016 14464 26022 14476
rect 26234 14464 26240 14476
rect 26016 14436 26240 14464
rect 26016 14424 26022 14436
rect 26234 14424 26240 14436
rect 26292 14424 26298 14476
rect 26970 14424 26976 14476
rect 27028 14424 27034 14476
rect 27172 14473 27200 14504
rect 28077 14501 28089 14504
rect 28123 14501 28135 14535
rect 28077 14495 28135 14501
rect 28368 14476 28396 14572
rect 29086 14560 29092 14612
rect 29144 14600 29150 14612
rect 29365 14603 29423 14609
rect 29365 14600 29377 14603
rect 29144 14572 29377 14600
rect 29144 14560 29150 14572
rect 29365 14569 29377 14572
rect 29411 14569 29423 14603
rect 29365 14563 29423 14569
rect 30650 14560 30656 14612
rect 30708 14560 30714 14612
rect 29730 14532 29736 14544
rect 29380 14504 29736 14532
rect 27157 14467 27215 14473
rect 27157 14433 27169 14467
rect 27203 14433 27215 14467
rect 27157 14427 27215 14433
rect 27338 14424 27344 14476
rect 27396 14424 27402 14476
rect 27617 14467 27675 14473
rect 27617 14433 27629 14467
rect 27663 14464 27675 14467
rect 27893 14467 27951 14473
rect 27893 14464 27905 14467
rect 27663 14436 27905 14464
rect 27663 14433 27675 14436
rect 27617 14427 27675 14433
rect 27893 14433 27905 14436
rect 27939 14464 27951 14467
rect 27939 14436 28304 14464
rect 27939 14433 27951 14436
rect 27893 14427 27951 14433
rect 26050 14396 26056 14408
rect 25700 14368 26056 14396
rect 26050 14356 26056 14368
rect 26108 14356 26114 14408
rect 22756 14300 24900 14328
rect 24946 14288 24952 14340
rect 25004 14288 25010 14340
rect 26252 14328 26280 14424
rect 26988 14396 27016 14424
rect 27249 14399 27307 14405
rect 27249 14396 27261 14399
rect 26988 14368 27261 14396
rect 27249 14365 27261 14368
rect 27295 14365 27307 14399
rect 27249 14359 27307 14365
rect 28077 14399 28135 14405
rect 28077 14365 28089 14399
rect 28123 14396 28135 14399
rect 28166 14396 28172 14408
rect 28123 14368 28172 14396
rect 28123 14365 28135 14368
rect 28077 14359 28135 14365
rect 28166 14356 28172 14368
rect 28224 14356 28230 14408
rect 28276 14396 28304 14436
rect 28350 14424 28356 14476
rect 28408 14424 28414 14476
rect 28626 14424 28632 14476
rect 28684 14464 28690 14476
rect 28721 14467 28779 14473
rect 28721 14464 28733 14467
rect 28684 14436 28733 14464
rect 28684 14424 28690 14436
rect 28721 14433 28733 14436
rect 28767 14433 28779 14467
rect 28721 14427 28779 14433
rect 28902 14424 28908 14476
rect 28960 14424 28966 14476
rect 29380 14473 29408 14504
rect 29730 14492 29736 14504
rect 29788 14532 29794 14544
rect 31110 14532 31116 14544
rect 29788 14504 30236 14532
rect 29788 14492 29794 14504
rect 30208 14476 30236 14504
rect 30760 14504 31116 14532
rect 29365 14467 29423 14473
rect 29365 14433 29377 14467
rect 29411 14433 29423 14467
rect 29365 14427 29423 14433
rect 29549 14467 29607 14473
rect 29549 14433 29561 14467
rect 29595 14464 29607 14467
rect 29595 14436 29776 14464
rect 29595 14433 29607 14436
rect 29549 14427 29607 14433
rect 29641 14399 29699 14405
rect 29641 14396 29653 14399
rect 28276 14368 29653 14396
rect 29641 14365 29653 14368
rect 29687 14365 29699 14399
rect 29748 14396 29776 14436
rect 29822 14424 29828 14476
rect 29880 14424 29886 14476
rect 30006 14424 30012 14476
rect 30064 14424 30070 14476
rect 30190 14424 30196 14476
rect 30248 14424 30254 14476
rect 30466 14424 30472 14476
rect 30524 14424 30530 14476
rect 30760 14473 30788 14504
rect 31110 14492 31116 14504
rect 31168 14492 31174 14544
rect 30745 14467 30803 14473
rect 30745 14433 30757 14467
rect 30791 14433 30803 14467
rect 30745 14427 30803 14433
rect 30837 14467 30895 14473
rect 30837 14433 30849 14467
rect 30883 14464 30895 14467
rect 30926 14464 30932 14476
rect 30883 14436 30932 14464
rect 30883 14433 30895 14436
rect 30837 14427 30895 14433
rect 30926 14424 30932 14436
rect 30984 14424 30990 14476
rect 30484 14396 30512 14424
rect 31202 14396 31208 14408
rect 29748 14368 29868 14396
rect 30484 14368 31208 14396
rect 29641 14359 29699 14365
rect 27522 14328 27528 14340
rect 26252 14300 27528 14328
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 29656 14328 29684 14359
rect 29730 14328 29736 14340
rect 29656 14300 29736 14328
rect 29730 14288 29736 14300
rect 29788 14288 29794 14340
rect 29840 14328 29868 14368
rect 31202 14356 31208 14368
rect 31260 14356 31266 14408
rect 30834 14328 30840 14340
rect 29840 14300 30840 14328
rect 30834 14288 30840 14300
rect 30892 14288 30898 14340
rect 17604 14232 20024 14260
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 22462 14260 22468 14272
rect 20220 14232 22468 14260
rect 20220 14220 20226 14232
rect 22462 14220 22468 14232
rect 22520 14220 22526 14272
rect 22830 14220 22836 14272
rect 22888 14220 22894 14272
rect 23385 14263 23443 14269
rect 23385 14229 23397 14263
rect 23431 14260 23443 14263
rect 23474 14260 23480 14272
rect 23431 14232 23480 14260
rect 23431 14229 23443 14232
rect 23385 14223 23443 14229
rect 23474 14220 23480 14232
rect 23532 14220 23538 14272
rect 24210 14220 24216 14272
rect 24268 14260 24274 14272
rect 24578 14260 24584 14272
rect 24268 14232 24584 14260
rect 24268 14220 24274 14232
rect 24578 14220 24584 14232
rect 24636 14220 24642 14272
rect 24762 14220 24768 14272
rect 24820 14220 24826 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 25682 14220 25688 14272
rect 25740 14220 25746 14272
rect 27801 14263 27859 14269
rect 27801 14229 27813 14263
rect 27847 14260 27859 14263
rect 27982 14260 27988 14272
rect 27847 14232 27988 14260
rect 27847 14229 27859 14232
rect 27801 14223 27859 14229
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 28074 14220 28080 14272
rect 28132 14260 28138 14272
rect 28261 14263 28319 14269
rect 28261 14260 28273 14263
rect 28132 14232 28273 14260
rect 28132 14220 28138 14232
rect 28261 14229 28273 14232
rect 28307 14229 28319 14263
rect 28261 14223 28319 14229
rect 28442 14220 28448 14272
rect 28500 14260 28506 14272
rect 28813 14263 28871 14269
rect 28813 14260 28825 14263
rect 28500 14232 28825 14260
rect 28500 14220 28506 14232
rect 28813 14229 28825 14232
rect 28859 14229 28871 14263
rect 28813 14223 28871 14229
rect 30282 14220 30288 14272
rect 30340 14260 30346 14272
rect 31021 14263 31079 14269
rect 31021 14260 31033 14263
rect 30340 14232 31033 14260
rect 30340 14220 30346 14232
rect 31021 14229 31033 14232
rect 31067 14229 31079 14263
rect 31021 14223 31079 14229
rect 552 14170 31648 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 11436 14170
rect 11488 14118 11500 14170
rect 11552 14118 11564 14170
rect 11616 14118 11628 14170
rect 11680 14118 11692 14170
rect 11744 14118 19210 14170
rect 19262 14118 19274 14170
rect 19326 14118 19338 14170
rect 19390 14118 19402 14170
rect 19454 14118 19466 14170
rect 19518 14118 26984 14170
rect 27036 14118 27048 14170
rect 27100 14118 27112 14170
rect 27164 14118 27176 14170
rect 27228 14118 27240 14170
rect 27292 14118 31648 14170
rect 552 14096 31648 14118
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 5350 14056 5356 14068
rect 3835 14028 5356 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5994 14056 6000 14068
rect 5500 14028 6000 14056
rect 5500 14016 5506 14028
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6328 14028 6837 14056
rect 6328 14016 6334 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7064 14028 8156 14056
rect 7064 14016 7070 14028
rect 4525 13991 4583 13997
rect 4525 13988 4537 13991
rect 3620 13960 4537 13988
rect 2958 13880 2964 13932
rect 3016 13920 3022 13932
rect 3620 13929 3648 13960
rect 4525 13957 4537 13960
rect 4571 13957 4583 13991
rect 4525 13951 4583 13957
rect 4724 13960 6592 13988
rect 3605 13923 3663 13929
rect 3016 13892 3556 13920
rect 3016 13880 3022 13892
rect 3326 13812 3332 13864
rect 3384 13812 3390 13864
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 3528 13852 3556 13892
rect 3605 13889 3617 13923
rect 3651 13889 3663 13923
rect 4724 13920 4752 13960
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 3605 13883 3663 13889
rect 3804 13892 4752 13920
rect 4816 13892 5273 13920
rect 3528 13824 3648 13852
rect 3620 13784 3648 13824
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 3804 13784 3832 13892
rect 4706 13812 4712 13864
rect 4764 13812 4770 13864
rect 4816 13861 4844 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 3620 13756 3832 13784
rect 4246 13744 4252 13796
rect 4304 13784 4310 13796
rect 4893 13787 4951 13793
rect 4893 13784 4905 13787
rect 4304 13756 4905 13784
rect 4304 13744 4310 13756
rect 4893 13753 4905 13756
rect 4939 13753 4951 13787
rect 5092 13784 5120 13815
rect 5166 13812 5172 13864
rect 5224 13812 5230 13864
rect 5442 13812 5448 13864
rect 5500 13812 5506 13864
rect 5552 13852 5580 13960
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 5684 13892 6316 13920
rect 5684 13880 5690 13892
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 5552 13824 5733 13852
rect 5721 13821 5733 13824
rect 5767 13821 5779 13855
rect 5721 13815 5779 13821
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 6288 13861 6316 13892
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 6052 13824 6193 13852
rect 6052 13812 6058 13824
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 6273 13855 6331 13861
rect 6273 13821 6285 13855
rect 6319 13821 6331 13855
rect 6273 13815 6331 13821
rect 6454 13812 6460 13864
rect 6512 13812 6518 13864
rect 6564 13861 6592 13960
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 6972 13960 7788 13988
rect 6972 13948 6978 13960
rect 6656 13892 7328 13920
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 5534 13784 5540 13796
rect 5092 13756 5540 13784
rect 4893 13747 4951 13753
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13784 5687 13787
rect 6472 13784 6500 13812
rect 5675 13756 6500 13784
rect 5675 13753 5687 13756
rect 5629 13747 5687 13753
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 3970 13716 3976 13728
rect 2648 13688 3976 13716
rect 2648 13676 2654 13688
rect 3970 13676 3976 13688
rect 4028 13716 4034 13728
rect 5442 13716 5448 13728
rect 4028 13688 5448 13716
rect 4028 13676 4034 13688
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 6656 13716 6684 13892
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 6779 13824 7021 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 7009 13821 7021 13824
rect 7055 13821 7067 13855
rect 7009 13815 7067 13821
rect 7098 13812 7104 13864
rect 7156 13812 7162 13864
rect 7300 13861 7328 13892
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 7374 13812 7380 13864
rect 7432 13812 7438 13864
rect 7760 13861 7788 13960
rect 8128 13920 8156 14028
rect 8386 14016 8392 14068
rect 8444 14016 8450 14068
rect 9398 14016 9404 14068
rect 9456 14016 9462 14068
rect 10137 14059 10195 14065
rect 10137 14025 10149 14059
rect 10183 14056 10195 14059
rect 10502 14056 10508 14068
rect 10183 14028 10508 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 11606 14056 11612 14068
rect 10612 14028 11612 14056
rect 8662 13948 8668 14000
rect 8720 13988 8726 14000
rect 8846 13988 8852 14000
rect 8720 13960 8852 13988
rect 8720 13948 8726 13960
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 8938 13948 8944 14000
rect 8996 13988 9002 14000
rect 9490 13988 9496 14000
rect 8996 13960 9496 13988
rect 8996 13948 9002 13960
rect 9490 13948 9496 13960
rect 9548 13988 9554 14000
rect 10612 13988 10640 14028
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 12526 14056 12532 14068
rect 11848 14028 12532 14056
rect 11848 14016 11854 14028
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 13228 14028 13553 14056
rect 13228 14016 13234 14028
rect 13541 14025 13553 14028
rect 13587 14025 13599 14059
rect 13541 14019 13599 14025
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14090 14056 14096 14068
rect 13872 14028 14096 14056
rect 13872 14016 13878 14028
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15289 14059 15347 14065
rect 15289 14056 15301 14059
rect 14976 14028 15301 14056
rect 14976 14016 14982 14028
rect 15289 14025 15301 14028
rect 15335 14025 15347 14059
rect 15289 14019 15347 14025
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16264 14028 16865 14056
rect 16264 14016 16270 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 18414 14016 18420 14068
rect 18472 14056 18478 14068
rect 18693 14059 18751 14065
rect 18693 14056 18705 14059
rect 18472 14028 18705 14056
rect 18472 14016 18478 14028
rect 18693 14025 18705 14028
rect 18739 14025 18751 14059
rect 18693 14019 18751 14025
rect 18874 14016 18880 14068
rect 18932 14056 18938 14068
rect 19334 14056 19340 14068
rect 18932 14028 19340 14056
rect 18932 14016 18938 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19794 14056 19800 14068
rect 19484 14028 19800 14056
rect 19484 14016 19490 14028
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 19886 14016 19892 14068
rect 19944 14056 19950 14068
rect 20438 14056 20444 14068
rect 19944 14028 20444 14056
rect 19944 14016 19950 14028
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 20806 14016 20812 14068
rect 20864 14016 20870 14068
rect 21542 14056 21548 14068
rect 20917 14028 21548 14056
rect 9548 13960 9720 13988
rect 9548 13948 9554 13960
rect 8128 13892 9168 13920
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8294 13852 8300 13864
rect 8168 13824 8300 13852
rect 8168 13812 8174 13824
rect 8294 13812 8300 13824
rect 8352 13852 8358 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8352 13824 8401 13852
rect 8352 13812 8358 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8570 13812 8576 13864
rect 8628 13812 8634 13864
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 6840 13756 7573 13784
rect 6840 13728 6868 13756
rect 7561 13753 7573 13756
rect 7607 13784 7619 13787
rect 7834 13784 7840 13796
rect 7607 13756 7840 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 7834 13744 7840 13756
rect 7892 13744 7898 13796
rect 8772 13784 8800 13815
rect 8938 13812 8944 13864
rect 8996 13812 9002 13864
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9140 13861 9168 13892
rect 9416 13892 9628 13920
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 9416 13852 9444 13892
rect 9171 13824 9444 13852
rect 9493 13855 9551 13861
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 8846 13784 8852 13796
rect 8772 13756 8852 13784
rect 8846 13744 8852 13756
rect 8904 13784 8910 13796
rect 9508 13784 9536 13815
rect 8904 13756 9536 13784
rect 9600 13784 9628 13892
rect 9692 13861 9720 13960
rect 10244 13960 10640 13988
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9766 13812 9772 13864
rect 9824 13812 9830 13864
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10244 13852 10272 13960
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 12250 13988 12256 14000
rect 11112 13960 12256 13988
rect 11112 13948 11118 13960
rect 12250 13948 12256 13960
rect 12308 13948 12314 14000
rect 15102 13988 15108 14000
rect 12360 13960 15108 13988
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 12360 13920 12388 13960
rect 15102 13948 15108 13960
rect 15160 13948 15166 14000
rect 17218 13948 17224 14000
rect 17276 13948 17282 14000
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17678 13988 17684 14000
rect 17368 13960 17684 13988
rect 17368 13948 17374 13960
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 18046 13948 18052 14000
rect 18104 13988 18110 14000
rect 19058 13988 19064 14000
rect 18104 13960 19064 13988
rect 18104 13948 18110 13960
rect 19058 13948 19064 13960
rect 19116 13988 19122 14000
rect 20917 13988 20945 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 21634 14016 21640 14068
rect 21692 14056 21698 14068
rect 21692 14028 22140 14056
rect 21692 14016 21698 14028
rect 19116 13960 20945 13988
rect 20993 13991 21051 13997
rect 19116 13948 19122 13960
rect 20993 13957 21005 13991
rect 21039 13957 21051 13991
rect 20993 13951 21051 13957
rect 21821 13991 21879 13997
rect 21821 13957 21833 13991
rect 21867 13957 21879 13991
rect 21821 13951 21879 13957
rect 10652 13892 12388 13920
rect 10652 13880 10658 13892
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 13136 13892 14044 13920
rect 13136 13880 13142 13892
rect 9907 13824 10272 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 9876 13784 9904 13815
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 10376 13824 13768 13852
rect 10376 13812 10382 13824
rect 9600 13756 9904 13784
rect 8904 13744 8910 13756
rect 10502 13744 10508 13796
rect 10560 13784 10566 13796
rect 13740 13784 13768 13824
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 13906 13812 13912 13864
rect 13964 13812 13970 13864
rect 14016 13861 14044 13892
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 15930 13920 15936 13932
rect 14148 13892 15936 13920
rect 14148 13880 14154 13892
rect 15930 13880 15936 13892
rect 15988 13920 15994 13932
rect 16482 13920 16488 13932
rect 15988 13892 16488 13920
rect 15988 13880 15994 13892
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 17696 13920 17724 13948
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 16724 13892 17356 13920
rect 17696 13892 17785 13920
rect 16724 13880 16730 13892
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 14090 13784 14096 13796
rect 10560 13756 13518 13784
rect 13740 13756 14096 13784
rect 10560 13744 10566 13756
rect 5868 13688 6684 13716
rect 5868 13676 5874 13688
rect 6822 13676 6828 13728
rect 6880 13676 6886 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 11146 13716 11152 13728
rect 7524 13688 11152 13716
rect 7524 13676 7530 13688
rect 11146 13676 11152 13688
rect 11204 13716 11210 13728
rect 12618 13716 12624 13728
rect 11204 13688 12624 13716
rect 11204 13676 11210 13688
rect 12618 13676 12624 13688
rect 12676 13716 12682 13728
rect 13354 13716 13360 13728
rect 12676 13688 13360 13716
rect 12676 13676 12682 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13490 13716 13518 13756
rect 14090 13744 14096 13756
rect 14148 13744 14154 13796
rect 14200 13784 14228 13815
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 14734 13852 14740 13864
rect 14608 13824 14740 13852
rect 14608 13812 14614 13824
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15102 13812 15108 13864
rect 15160 13812 15166 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15378 13852 15384 13864
rect 15335 13824 15384 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 17034 13812 17040 13864
rect 17092 13812 17098 13864
rect 17126 13812 17132 13864
rect 17184 13812 17190 13864
rect 17328 13861 17356 13892
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13920 18015 13923
rect 18230 13920 18236 13932
rect 18003 13892 18236 13920
rect 18003 13889 18015 13892
rect 17957 13883 18015 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 18472 13892 18981 13920
rect 18472 13880 18478 13892
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 20441 13923 20499 13929
rect 20441 13920 20453 13923
rect 18969 13883 19027 13889
rect 19076 13892 20453 13920
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 15194 13784 15200 13796
rect 14200 13756 15200 13784
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 17696 13784 17724 13815
rect 17862 13812 17868 13864
rect 17920 13812 17926 13864
rect 19076 13784 19104 13892
rect 20441 13889 20453 13892
rect 20487 13920 20499 13923
rect 20898 13920 20904 13932
rect 20487 13892 20904 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 21008 13920 21036 13951
rect 21008 13892 21404 13920
rect 19150 13812 19156 13864
rect 19208 13812 19214 13864
rect 19242 13812 19248 13864
rect 19300 13812 19306 13864
rect 19426 13812 19432 13864
rect 19484 13812 19490 13864
rect 20530 13812 20536 13864
rect 20588 13852 20594 13864
rect 21376 13861 21404 13892
rect 21726 13880 21732 13932
rect 21784 13880 21790 13932
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20588 13824 21097 13852
rect 20588 13812 20594 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 21269 13815 21327 13821
rect 21361 13855 21419 13861
rect 21361 13821 21373 13855
rect 21407 13821 21419 13855
rect 21361 13815 21419 13821
rect 17696 13756 19104 13784
rect 19168 13784 19196 13812
rect 20162 13784 20168 13796
rect 19168 13756 20168 13784
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 20346 13744 20352 13796
rect 20404 13784 20410 13796
rect 21174 13784 21180 13796
rect 20404 13756 21180 13784
rect 20404 13744 20410 13756
rect 21174 13744 21180 13756
rect 21232 13744 21238 13796
rect 21284 13784 21312 13815
rect 21450 13812 21456 13864
rect 21508 13812 21514 13864
rect 21836 13852 21864 13951
rect 22112 13929 22140 14028
rect 22278 14016 22284 14068
rect 22336 14016 22342 14068
rect 22830 14016 22836 14068
rect 22888 14056 22894 14068
rect 22925 14059 22983 14065
rect 22925 14056 22937 14059
rect 22888 14028 22937 14056
rect 22888 14016 22894 14028
rect 22925 14025 22937 14028
rect 22971 14025 22983 14059
rect 22925 14019 22983 14025
rect 23934 14016 23940 14068
rect 23992 14056 23998 14068
rect 25314 14056 25320 14068
rect 23992 14028 25320 14056
rect 23992 14016 23998 14028
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 25590 14016 25596 14068
rect 25648 14016 25654 14068
rect 26694 14016 26700 14068
rect 26752 14056 26758 14068
rect 28626 14056 28632 14068
rect 26752 14028 28632 14056
rect 26752 14016 26758 14028
rect 28626 14016 28632 14028
rect 28684 14016 28690 14068
rect 28810 14016 28816 14068
rect 28868 14056 28874 14068
rect 30285 14059 30343 14065
rect 30285 14056 30297 14059
rect 28868 14028 30297 14056
rect 28868 14016 28874 14028
rect 30285 14025 30297 14028
rect 30331 14025 30343 14059
rect 30285 14019 30343 14025
rect 30742 14016 30748 14068
rect 30800 14056 30806 14068
rect 31113 14059 31171 14065
rect 31113 14056 31125 14059
rect 30800 14028 31125 14056
rect 30800 14016 30806 14028
rect 31113 14025 31125 14028
rect 31159 14025 31171 14059
rect 31113 14019 31171 14025
rect 24118 13948 24124 14000
rect 24176 13988 24182 14000
rect 24578 13988 24584 14000
rect 24176 13960 24584 13988
rect 24176 13948 24182 13960
rect 24578 13948 24584 13960
rect 24636 13988 24642 14000
rect 25682 13988 25688 14000
rect 24636 13960 25688 13988
rect 24636 13948 24642 13960
rect 25682 13948 25688 13960
rect 25740 13948 25746 14000
rect 25777 13991 25835 13997
rect 25777 13957 25789 13991
rect 25823 13988 25835 13991
rect 25958 13988 25964 14000
rect 25823 13960 25964 13988
rect 25823 13957 25835 13960
rect 25777 13951 25835 13957
rect 25958 13948 25964 13960
rect 26016 13988 26022 14000
rect 26602 13988 26608 14000
rect 26016 13960 26608 13988
rect 26016 13948 26022 13960
rect 26602 13948 26608 13960
rect 26660 13988 26666 14000
rect 26878 13988 26884 14000
rect 26660 13960 26884 13988
rect 26660 13948 26666 13960
rect 26878 13948 26884 13960
rect 26936 13948 26942 14000
rect 28166 13948 28172 14000
rect 28224 13988 28230 14000
rect 28442 13988 28448 14000
rect 28224 13960 28448 13988
rect 28224 13948 28230 13960
rect 28442 13948 28448 13960
rect 28500 13948 28506 14000
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22296 13892 24716 13920
rect 22296 13861 22324 13892
rect 21560 13824 21864 13852
rect 22005 13855 22063 13861
rect 21560 13784 21588 13824
rect 22005 13821 22017 13855
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 22281 13855 22339 13861
rect 22281 13821 22293 13855
rect 22327 13821 22339 13855
rect 22281 13815 22339 13821
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 22462 13852 22468 13864
rect 22419 13824 22468 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 21284 13756 21588 13784
rect 22020 13728 22048 13815
rect 22462 13812 22468 13824
rect 22520 13852 22526 13864
rect 23566 13852 23572 13864
rect 22520 13824 23572 13852
rect 22520 13812 22526 13824
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 24688 13852 24716 13892
rect 24762 13880 24768 13932
rect 24820 13920 24826 13932
rect 24820 13892 26096 13920
rect 24820 13880 24826 13892
rect 25406 13852 25412 13864
rect 24688 13824 25412 13852
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25682 13812 25688 13864
rect 25740 13812 25746 13864
rect 25958 13812 25964 13864
rect 26016 13812 26022 13864
rect 26068 13861 26096 13892
rect 28368 13892 29224 13920
rect 26053 13855 26111 13861
rect 26053 13821 26065 13855
rect 26099 13821 26111 13855
rect 26053 13815 26111 13821
rect 28258 13812 28264 13864
rect 28316 13812 28322 13864
rect 28368 13861 28396 13892
rect 28353 13855 28411 13861
rect 28353 13821 28365 13855
rect 28399 13821 28411 13855
rect 28353 13815 28411 13821
rect 28537 13855 28595 13861
rect 28537 13821 28549 13855
rect 28583 13821 28595 13855
rect 28537 13815 28595 13821
rect 28629 13855 28687 13861
rect 28629 13821 28641 13855
rect 28675 13821 28687 13855
rect 28629 13815 28687 13821
rect 28813 13855 28871 13861
rect 28813 13821 28825 13855
rect 28859 13852 28871 13855
rect 29086 13852 29092 13864
rect 28859 13824 29092 13852
rect 28859 13821 28871 13824
rect 28813 13815 28871 13821
rect 22557 13787 22615 13793
rect 22557 13753 22569 13787
rect 22603 13784 22615 13787
rect 23382 13784 23388 13796
rect 22603 13756 23388 13784
rect 22603 13753 22615 13756
rect 22557 13747 22615 13753
rect 23382 13744 23388 13756
rect 23440 13744 23446 13796
rect 23658 13744 23664 13796
rect 23716 13784 23722 13796
rect 25130 13784 25136 13796
rect 23716 13756 25136 13784
rect 23716 13744 23722 13756
rect 25130 13744 25136 13756
rect 25188 13744 25194 13796
rect 25424 13784 25452 13812
rect 28552 13784 28580 13815
rect 25424 13756 28580 13784
rect 28644 13784 28672 13815
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 29196 13852 29224 13892
rect 30650 13880 30656 13932
rect 30708 13920 30714 13932
rect 30708 13892 30972 13920
rect 30708 13880 30714 13892
rect 29917 13855 29975 13861
rect 29917 13852 29929 13855
rect 29196 13824 29929 13852
rect 29917 13821 29929 13824
rect 29963 13852 29975 13855
rect 30190 13852 30196 13864
rect 29963 13824 30196 13852
rect 29963 13821 29975 13824
rect 29917 13815 29975 13821
rect 30190 13812 30196 13824
rect 30248 13812 30254 13864
rect 30944 13861 30972 13892
rect 30377 13855 30435 13861
rect 30377 13821 30389 13855
rect 30423 13852 30435 13855
rect 30929 13855 30987 13861
rect 30423 13824 30880 13852
rect 30423 13821 30435 13824
rect 30377 13815 30435 13821
rect 29362 13784 29368 13796
rect 28644 13756 29368 13784
rect 15654 13716 15660 13728
rect 13490 13688 15660 13716
rect 15654 13676 15660 13688
rect 15712 13716 15718 13728
rect 19150 13716 19156 13728
rect 15712 13688 19156 13716
rect 15712 13676 15718 13688
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 19610 13676 19616 13728
rect 19668 13716 19674 13728
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 19668 13688 20821 13716
rect 19668 13676 19674 13688
rect 20809 13685 20821 13688
rect 20855 13716 20867 13719
rect 22002 13716 22008 13728
rect 20855 13688 22008 13716
rect 20855 13685 20867 13688
rect 20809 13679 20867 13685
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 22462 13676 22468 13728
rect 22520 13716 22526 13728
rect 22649 13719 22707 13725
rect 22649 13716 22661 13719
rect 22520 13688 22661 13716
rect 22520 13676 22526 13688
rect 22649 13685 22661 13688
rect 22695 13685 22707 13719
rect 22649 13679 22707 13685
rect 22738 13676 22744 13728
rect 22796 13676 22802 13728
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 25498 13716 25504 13728
rect 22888 13688 25504 13716
rect 22888 13676 22894 13688
rect 25498 13676 25504 13688
rect 25556 13676 25562 13728
rect 25590 13676 25596 13728
rect 25648 13716 25654 13728
rect 27890 13716 27896 13728
rect 25648 13688 27896 13716
rect 25648 13676 25654 13688
rect 27890 13676 27896 13688
rect 27948 13716 27954 13728
rect 28442 13716 28448 13728
rect 27948 13688 28448 13716
rect 27948 13676 27954 13688
rect 28442 13676 28448 13688
rect 28500 13676 28506 13728
rect 28552 13716 28580 13756
rect 29362 13744 29368 13756
rect 29420 13744 29426 13796
rect 30098 13744 30104 13796
rect 30156 13744 30162 13796
rect 30852 13784 30880 13824
rect 30929 13821 30941 13855
rect 30975 13821 30987 13855
rect 30929 13815 30987 13821
rect 31018 13812 31024 13864
rect 31076 13812 31082 13864
rect 31036 13784 31064 13812
rect 30852 13756 31064 13784
rect 28902 13716 28908 13728
rect 28552 13688 28908 13716
rect 28902 13676 28908 13688
rect 28960 13676 28966 13728
rect 29546 13676 29552 13728
rect 29604 13716 29610 13728
rect 29641 13719 29699 13725
rect 29641 13716 29653 13719
rect 29604 13688 29653 13716
rect 29604 13676 29610 13688
rect 29641 13685 29653 13688
rect 29687 13685 29699 13719
rect 29641 13679 29699 13685
rect 30009 13719 30067 13725
rect 30009 13685 30021 13719
rect 30055 13716 30067 13719
rect 30282 13716 30288 13728
rect 30055 13688 30288 13716
rect 30055 13685 30067 13688
rect 30009 13679 30067 13685
rect 30282 13676 30288 13688
rect 30340 13676 30346 13728
rect 552 13626 31648 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 12096 13626
rect 12148 13574 12160 13626
rect 12212 13574 12224 13626
rect 12276 13574 12288 13626
rect 12340 13574 12352 13626
rect 12404 13574 19870 13626
rect 19922 13574 19934 13626
rect 19986 13574 19998 13626
rect 20050 13574 20062 13626
rect 20114 13574 20126 13626
rect 20178 13574 27644 13626
rect 27696 13574 27708 13626
rect 27760 13574 27772 13626
rect 27824 13574 27836 13626
rect 27888 13574 27900 13626
rect 27952 13574 31648 13626
rect 552 13552 31648 13574
rect 845 13515 903 13521
rect 845 13481 857 13515
rect 891 13512 903 13515
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 891 13484 1869 13512
rect 891 13481 903 13484
rect 845 13475 903 13481
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 2041 13515 2099 13521
rect 2041 13481 2053 13515
rect 2087 13512 2099 13515
rect 3510 13512 3516 13524
rect 2087 13484 3516 13512
rect 2087 13481 2099 13484
rect 2041 13475 2099 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 5166 13512 5172 13524
rect 4580 13484 5172 13512
rect 4580 13472 4586 13484
rect 5166 13472 5172 13484
rect 5224 13512 5230 13524
rect 7558 13512 7564 13524
rect 5224 13484 7236 13512
rect 5224 13472 5230 13484
rect 7208 13456 7236 13484
rect 7392 13484 7564 13512
rect 1213 13447 1271 13453
rect 1213 13413 1225 13447
rect 1259 13444 1271 13447
rect 1259 13416 1440 13444
rect 1259 13413 1271 13416
rect 1213 13407 1271 13413
rect 1026 13336 1032 13388
rect 1084 13336 1090 13388
rect 1305 13379 1363 13385
rect 1305 13345 1317 13379
rect 1351 13345 1363 13379
rect 1412 13376 1440 13416
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 1544 13416 2912 13444
rect 1544 13404 1550 13416
rect 1762 13376 1768 13388
rect 1412 13348 1768 13376
rect 1305 13339 1363 13345
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1320 13308 1348 13339
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 1946 13385 1952 13388
rect 1916 13379 1952 13385
rect 1916 13345 1928 13379
rect 1916 13339 1952 13345
rect 1946 13336 1952 13339
rect 2004 13336 2010 13388
rect 2516 13385 2544 13416
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2648 13348 2697 13376
rect 2648 13336 2654 13348
rect 2685 13345 2697 13348
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 2884 13385 2912 13416
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 5534 13444 5540 13456
rect 3752 13416 5540 13444
rect 3752 13404 3758 13416
rect 5534 13404 5540 13416
rect 5592 13444 5598 13456
rect 5902 13444 5908 13456
rect 5592 13416 5908 13444
rect 5592 13404 5598 13416
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 5994 13404 6000 13456
rect 6052 13444 6058 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 6052 13416 6561 13444
rect 6052 13404 6058 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 7006 13444 7012 13456
rect 6549 13407 6607 13413
rect 6656 13416 7012 13444
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 3050 13336 3056 13388
rect 3108 13336 3114 13388
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 4982 13376 4988 13388
rect 4672 13348 4988 13376
rect 4672 13336 4678 13348
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 5224 13348 6469 13376
rect 5224 13336 5230 13348
rect 6457 13345 6469 13348
rect 6503 13376 6515 13379
rect 6656 13376 6684 13416
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 7190 13404 7196 13456
rect 7248 13404 7254 13456
rect 7392 13453 7420 13484
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 7708 13484 8805 13512
rect 7708 13472 7714 13484
rect 7377 13447 7435 13453
rect 7377 13413 7389 13447
rect 7423 13413 7435 13447
rect 8777 13444 8805 13484
rect 8846 13472 8852 13524
rect 8904 13472 8910 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 11238 13512 11244 13524
rect 9180 13484 10640 13512
rect 9180 13472 9186 13484
rect 8938 13444 8944 13456
rect 7377 13407 7435 13413
rect 7852 13416 8708 13444
rect 8777 13416 8944 13444
rect 6503 13348 6684 13376
rect 6733 13379 6791 13385
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6733 13345 6745 13379
rect 6779 13376 6791 13379
rect 6822 13376 6828 13388
rect 6779 13348 6828 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7558 13336 7564 13388
rect 7616 13336 7622 13388
rect 992 13280 1348 13308
rect 1397 13311 1455 13317
rect 992 13268 998 13280
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1443 13280 2360 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 2332 13184 2360 13280
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 7006 13308 7012 13320
rect 5960 13280 7012 13308
rect 5960 13268 5966 13280
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7852 13308 7880 13416
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 7984 13348 8309 13376
rect 7984 13336 7990 13348
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8478 13376 8484 13388
rect 8435 13348 8484 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 8570 13336 8576 13388
rect 8628 13336 8634 13388
rect 8680 13385 8708 13416
rect 8938 13404 8944 13416
rect 8996 13404 9002 13456
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 10502 13444 10508 13456
rect 9916 13416 10508 13444
rect 9916 13404 9922 13416
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 10612 13388 10640 13484
rect 11026 13484 11244 13512
rect 10778 13404 10784 13456
rect 10836 13444 10842 13456
rect 11026 13444 11054 13484
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 11974 13512 11980 13524
rect 11848 13484 11980 13512
rect 11848 13472 11854 13484
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12161 13515 12219 13521
rect 12161 13481 12173 13515
rect 12207 13512 12219 13515
rect 12250 13512 12256 13524
rect 12207 13484 12256 13512
rect 12207 13481 12219 13484
rect 12161 13475 12219 13481
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 12526 13512 12532 13524
rect 12360 13484 12532 13512
rect 10836 13416 11054 13444
rect 11256 13444 11284 13472
rect 11256 13416 11504 13444
rect 10836 13404 10842 13416
rect 8665 13379 8723 13385
rect 8665 13345 8677 13379
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 10042 13376 10048 13388
rect 8904 13348 10048 13376
rect 8904 13336 8910 13348
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10318 13385 10324 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10285 13379 10324 13385
rect 10285 13345 10297 13379
rect 10285 13339 10324 13345
rect 9950 13308 9956 13320
rect 7340 13280 7880 13308
rect 8319 13280 9956 13308
rect 7340 13268 7346 13280
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 4338 13240 4344 13252
rect 4028 13212 4344 13240
rect 4028 13200 4034 13212
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 7374 13240 7380 13252
rect 4488 13212 7380 13240
rect 4488 13200 4494 13212
rect 7374 13200 7380 13212
rect 7432 13240 7438 13252
rect 7432 13212 7604 13240
rect 7432 13200 7438 13212
rect 1486 13132 1492 13184
rect 1544 13132 1550 13184
rect 2314 13132 2320 13184
rect 2372 13132 2378 13184
rect 2866 13132 2872 13184
rect 2924 13132 2930 13184
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13172 3295 13175
rect 3326 13172 3332 13184
rect 3283 13144 3332 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 5902 13172 5908 13184
rect 4212 13144 5908 13172
rect 4212 13132 4218 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6270 13132 6276 13184
rect 6328 13172 6334 13184
rect 6546 13172 6552 13184
rect 6328 13144 6552 13172
rect 6328 13132 6334 13144
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7098 13172 7104 13184
rect 6963 13144 7104 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7576 13172 7604 13212
rect 7650 13200 7656 13252
rect 7708 13240 7714 13252
rect 7745 13243 7803 13249
rect 7745 13240 7757 13243
rect 7708 13212 7757 13240
rect 7708 13200 7714 13212
rect 7745 13209 7757 13212
rect 7791 13240 7803 13243
rect 8319 13240 8347 13280
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10152 13308 10180 13339
rect 10318 13336 10324 13339
rect 10376 13336 10382 13388
rect 10410 13336 10416 13388
rect 10468 13336 10474 13388
rect 10594 13336 10600 13388
rect 10652 13385 10658 13388
rect 10652 13376 10660 13385
rect 11144 13379 11202 13385
rect 11144 13376 11156 13379
rect 10652 13348 10697 13376
rect 10796 13348 11156 13376
rect 10652 13339 10660 13348
rect 10652 13336 10658 13339
rect 10502 13308 10508 13320
rect 10152 13280 10508 13308
rect 10502 13268 10508 13280
rect 10560 13268 10566 13320
rect 8478 13240 8484 13252
rect 7791 13212 8347 13240
rect 8405 13212 8484 13240
rect 7791 13209 7803 13212
rect 7745 13203 7803 13209
rect 7926 13172 7932 13184
rect 7576 13144 7932 13172
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8405 13172 8433 13212
rect 8478 13200 8484 13212
rect 8536 13200 8542 13252
rect 10796 13249 10824 13348
rect 11144 13345 11156 13348
rect 11190 13345 11202 13379
rect 11144 13339 11202 13345
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13345 11299 13379
rect 11241 13339 11299 13345
rect 10781 13243 10839 13249
rect 10781 13209 10793 13243
rect 10827 13209 10839 13243
rect 10781 13203 10839 13209
rect 10962 13200 10968 13252
rect 11020 13200 11026 13252
rect 11256 13240 11284 13339
rect 11330 13336 11336 13388
rect 11388 13336 11394 13388
rect 11476 13385 11504 13416
rect 11698 13404 11704 13456
rect 11756 13444 11762 13456
rect 12360 13444 12388 13484
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12952 13484 13001 13512
rect 12952 13472 12958 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13412 13484 15332 13512
rect 13412 13472 13418 13484
rect 13446 13444 13452 13456
rect 11756 13416 12388 13444
rect 12636 13416 13452 13444
rect 11756 13404 11762 13416
rect 11461 13379 11519 13385
rect 11461 13345 11473 13379
rect 11507 13345 11519 13379
rect 11461 13339 11519 13345
rect 11606 13336 11612 13388
rect 11664 13336 11670 13388
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12636 13385 12664 13416
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 14274 13404 14280 13456
rect 14332 13444 14338 13456
rect 15304 13444 15332 13484
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15528 13484 16129 13512
rect 15528 13472 15534 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 16117 13475 16175 13481
rect 18414 13472 18420 13524
rect 18472 13512 18478 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 18472 13484 18889 13512
rect 18472 13472 18478 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 18966 13472 18972 13524
rect 19024 13512 19030 13524
rect 22094 13512 22100 13524
rect 19024 13484 20576 13512
rect 19024 13472 19030 13484
rect 15930 13444 15936 13456
rect 14332 13416 15240 13444
rect 15304 13416 15936 13444
rect 14332 13404 14338 13416
rect 12621 13379 12679 13385
rect 11848 13348 12204 13376
rect 11848 13336 11854 13348
rect 11624 13308 11652 13336
rect 12066 13308 12072 13320
rect 11624 13280 12072 13308
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12176 13240 12204 13348
rect 12621 13345 12633 13379
rect 12667 13345 12679 13379
rect 12621 13339 12679 13345
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 13044 13348 13277 13376
rect 13044 13336 13050 13348
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 14642 13376 14648 13388
rect 13265 13339 13323 13345
rect 13556 13348 14648 13376
rect 13556 13320 13584 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 15013 13379 15071 13385
rect 15013 13345 15025 13379
rect 15059 13345 15071 13379
rect 15013 13339 15071 13345
rect 12250 13268 12256 13320
rect 12308 13308 12314 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12308 13280 12357 13308
rect 12308 13268 12314 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12434 13268 12440 13320
rect 12492 13268 12498 13320
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 13078 13308 13084 13320
rect 12768 13280 13084 13308
rect 12768 13268 12774 13280
rect 13078 13268 13084 13280
rect 13136 13308 13142 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13136 13280 13185 13308
rect 13136 13268 13142 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13538 13268 13544 13320
rect 13596 13268 13602 13320
rect 13633 13311 13691 13317
rect 13633 13277 13645 13311
rect 13679 13308 13691 13311
rect 13722 13308 13728 13320
rect 13679 13280 13728 13308
rect 13679 13277 13691 13280
rect 13633 13271 13691 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 14734 13268 14740 13320
rect 14792 13268 14798 13320
rect 15028 13308 15056 13339
rect 15102 13336 15108 13388
rect 15160 13336 15166 13388
rect 15212 13385 15240 13416
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 20070 13444 20076 13456
rect 16500 13416 20076 13444
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13376 15255 13379
rect 15286 13376 15292 13388
rect 15243 13348 15292 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13376 15439 13379
rect 15746 13376 15752 13388
rect 15427 13348 15752 13376
rect 15427 13345 15439 13348
rect 15381 13339 15439 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 15838 13336 15844 13388
rect 15896 13336 15902 13388
rect 16206 13336 16212 13388
rect 16264 13376 16270 13388
rect 16500 13385 16528 13416
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 16264 13348 16313 13376
rect 16264 13336 16270 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13345 16543 13379
rect 16485 13339 16543 13345
rect 17034 13336 17040 13388
rect 17092 13336 17098 13388
rect 17218 13336 17224 13388
rect 17276 13336 17282 13388
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13376 17555 13379
rect 17586 13376 17592 13388
rect 17543 13348 17592 13376
rect 17543 13345 17555 13348
rect 17497 13339 17555 13345
rect 17586 13336 17592 13348
rect 17644 13336 17650 13388
rect 18138 13336 18144 13388
rect 18196 13376 18202 13388
rect 18196 13348 18552 13376
rect 18196 13336 18202 13348
rect 15470 13308 15476 13320
rect 15028 13280 15476 13308
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 18414 13308 18420 13320
rect 16224 13280 18420 13308
rect 12802 13240 12808 13252
rect 11256 13212 12112 13240
rect 12176 13212 12808 13240
rect 11790 13172 11796 13184
rect 8076 13144 11796 13172
rect 8076 13132 8082 13144
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 12084 13172 12112 13212
rect 12802 13200 12808 13212
rect 12860 13240 12866 13252
rect 14274 13240 14280 13252
rect 12860 13212 14280 13240
rect 12860 13200 12866 13212
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 15286 13200 15292 13252
rect 15344 13240 15350 13252
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 15344 13212 15577 13240
rect 15344 13200 15350 13212
rect 15565 13209 15577 13212
rect 15611 13209 15623 13243
rect 15565 13203 15623 13209
rect 13814 13172 13820 13184
rect 12084 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 16224 13172 16252 13280
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 18524 13308 18552 13348
rect 18782 13336 18788 13388
rect 18840 13336 18846 13388
rect 19058 13336 19064 13388
rect 19116 13336 19122 13388
rect 19150 13336 19156 13388
rect 19208 13336 19214 13388
rect 19242 13336 19248 13388
rect 19300 13336 19306 13388
rect 19429 13379 19487 13385
rect 19429 13345 19441 13379
rect 19475 13376 19487 13379
rect 19886 13376 19892 13388
rect 19475 13348 19892 13376
rect 19475 13345 19487 13348
rect 19429 13339 19487 13345
rect 19886 13336 19892 13348
rect 19944 13376 19950 13388
rect 20346 13376 20352 13388
rect 19944 13348 20352 13376
rect 19944 13336 19950 13348
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 18969 13311 19027 13317
rect 18969 13308 18981 13311
rect 18524 13280 18981 13308
rect 18969 13277 18981 13280
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 20254 13308 20260 13320
rect 19392 13280 20260 13308
rect 19392 13268 19398 13280
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 20548 13308 20576 13484
rect 20824 13484 22100 13512
rect 20824 13385 20852 13484
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22244 13484 22416 13512
rect 22244 13472 22250 13484
rect 21174 13404 21180 13456
rect 21232 13444 21238 13456
rect 22281 13447 22339 13453
rect 22281 13444 22293 13447
rect 21232 13416 22293 13444
rect 21232 13404 21238 13416
rect 22281 13413 22293 13416
rect 22327 13413 22339 13447
rect 22388 13444 22416 13484
rect 22738 13472 22744 13524
rect 22796 13472 22802 13524
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 25314 13512 25320 13524
rect 23164 13484 25320 13512
rect 23164 13472 23170 13484
rect 25314 13472 25320 13484
rect 25372 13472 25378 13524
rect 25498 13472 25504 13524
rect 25556 13472 25562 13524
rect 25590 13472 25596 13524
rect 25648 13472 25654 13524
rect 28074 13512 28080 13524
rect 25792 13484 28080 13512
rect 25038 13444 25044 13456
rect 22388 13416 25044 13444
rect 22281 13407 22339 13413
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13345 20867 13379
rect 20809 13339 20867 13345
rect 20898 13336 20904 13388
rect 20956 13336 20962 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 21008 13348 21465 13376
rect 21008 13308 21036 13348
rect 21453 13345 21465 13348
rect 21499 13345 21511 13379
rect 21453 13339 21511 13345
rect 21634 13336 21640 13388
rect 21692 13336 21698 13388
rect 21729 13379 21787 13385
rect 21729 13345 21741 13379
rect 21775 13345 21787 13379
rect 21729 13339 21787 13345
rect 20548 13280 21036 13308
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 21174 13308 21180 13320
rect 21131 13280 21180 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 21174 13268 21180 13280
rect 21232 13268 21238 13320
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 21744 13308 21772 13339
rect 21910 13336 21916 13388
rect 21968 13376 21974 13388
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21968 13348 22017 13376
rect 21968 13336 21974 13348
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 22370 13376 22376 13388
rect 22152 13348 22376 13376
rect 22152 13336 22158 13348
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 22940 13385 22968 13416
rect 25038 13404 25044 13416
rect 25096 13404 25102 13456
rect 25608 13444 25636 13472
rect 25332 13416 25636 13444
rect 22925 13379 22983 13385
rect 22925 13345 22937 13379
rect 22971 13345 22983 13379
rect 22925 13339 22983 13345
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13376 23259 13379
rect 23658 13376 23664 13388
rect 23247 13348 23664 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 24026 13336 24032 13388
rect 24084 13336 24090 13388
rect 24397 13379 24455 13385
rect 24397 13345 24409 13379
rect 24443 13376 24455 13379
rect 24486 13376 24492 13388
rect 24443 13348 24492 13376
rect 24443 13345 24455 13348
rect 24397 13339 24455 13345
rect 24486 13336 24492 13348
rect 24544 13336 24550 13388
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13376 24915 13379
rect 24946 13376 24952 13388
rect 24903 13348 24952 13376
rect 24903 13345 24915 13348
rect 24857 13339 24915 13345
rect 24946 13336 24952 13348
rect 25004 13336 25010 13388
rect 25332 13385 25360 13416
rect 25317 13379 25375 13385
rect 25317 13345 25329 13379
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 25406 13336 25412 13388
rect 25464 13336 25470 13388
rect 25593 13379 25651 13385
rect 25593 13345 25605 13379
rect 25639 13376 25651 13379
rect 25792 13376 25820 13484
rect 28074 13472 28080 13484
rect 28132 13512 28138 13524
rect 28721 13515 28779 13521
rect 28132 13484 28672 13512
rect 28132 13472 28138 13484
rect 26053 13447 26111 13453
rect 26053 13413 26065 13447
rect 26099 13444 26111 13447
rect 26142 13444 26148 13456
rect 26099 13416 26148 13444
rect 26099 13413 26111 13416
rect 26053 13407 26111 13413
rect 26142 13404 26148 13416
rect 26200 13404 26206 13456
rect 26237 13447 26295 13453
rect 26237 13413 26249 13447
rect 26283 13444 26295 13447
rect 26326 13444 26332 13456
rect 26283 13416 26332 13444
rect 26283 13413 26295 13416
rect 26237 13407 26295 13413
rect 26326 13404 26332 13416
rect 26384 13444 26390 13456
rect 26510 13444 26516 13456
rect 26384 13416 26516 13444
rect 26384 13404 26390 13416
rect 26510 13404 26516 13416
rect 26568 13404 26574 13456
rect 27798 13444 27804 13456
rect 26712 13416 27804 13444
rect 25639 13348 25820 13376
rect 25639 13345 25651 13348
rect 25593 13339 25651 13345
rect 25866 13336 25872 13388
rect 25924 13376 25930 13388
rect 25961 13379 26019 13385
rect 25961 13376 25973 13379
rect 25924 13348 25973 13376
rect 25924 13336 25930 13348
rect 25961 13345 25973 13348
rect 26007 13345 26019 13379
rect 25961 13339 26019 13345
rect 26421 13379 26479 13385
rect 26421 13345 26433 13379
rect 26467 13345 26479 13379
rect 26421 13339 26479 13345
rect 21324 13280 21772 13308
rect 22189 13311 22247 13317
rect 21324 13268 21330 13280
rect 22189 13277 22201 13311
rect 22235 13308 22247 13311
rect 22830 13308 22836 13320
rect 22235 13280 22836 13308
rect 22235 13277 22247 13280
rect 22189 13271 22247 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 24210 13308 24216 13320
rect 24044 13280 24216 13308
rect 24044 13252 24072 13280
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 25041 13311 25099 13317
rect 25041 13308 25053 13311
rect 24320 13280 25053 13308
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17310 13240 17316 13252
rect 17092 13212 17316 13240
rect 17092 13200 17098 13212
rect 17310 13200 17316 13212
rect 17368 13200 17374 13252
rect 17402 13200 17408 13252
rect 17460 13200 17466 13252
rect 17954 13200 17960 13252
rect 18012 13240 18018 13252
rect 21821 13243 21879 13249
rect 21821 13240 21833 13243
rect 18012 13212 21833 13240
rect 18012 13200 18018 13212
rect 21821 13209 21833 13212
rect 21867 13209 21879 13243
rect 21821 13203 21879 13209
rect 24026 13200 24032 13252
rect 24084 13200 24090 13252
rect 24320 13240 24348 13280
rect 25041 13277 25053 13280
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 25130 13268 25136 13320
rect 25188 13268 25194 13320
rect 25774 13268 25780 13320
rect 25832 13308 25838 13320
rect 26436 13308 26464 13339
rect 26602 13336 26608 13388
rect 26660 13336 26666 13388
rect 26712 13385 26740 13416
rect 27798 13404 27804 13416
rect 27856 13404 27862 13456
rect 27890 13404 27896 13456
rect 27948 13444 27954 13456
rect 27948 13416 28396 13444
rect 27948 13404 27954 13416
rect 26697 13379 26755 13385
rect 26697 13345 26709 13379
rect 26743 13345 26755 13379
rect 26697 13339 26755 13345
rect 26970 13336 26976 13388
rect 27028 13376 27034 13388
rect 27614 13376 27620 13388
rect 27028 13348 27620 13376
rect 27028 13336 27034 13348
rect 27614 13336 27620 13348
rect 27672 13336 27678 13388
rect 27706 13336 27712 13388
rect 27764 13376 27770 13388
rect 28077 13379 28135 13385
rect 28077 13376 28089 13379
rect 27764 13348 28089 13376
rect 27764 13336 27770 13348
rect 28077 13345 28089 13348
rect 28123 13376 28135 13379
rect 28166 13376 28172 13388
rect 28123 13348 28172 13376
rect 28123 13345 28135 13348
rect 28077 13339 28135 13345
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 28368 13385 28396 13416
rect 28353 13379 28411 13385
rect 28353 13345 28365 13379
rect 28399 13345 28411 13379
rect 28353 13339 28411 13345
rect 28442 13336 28448 13388
rect 28500 13336 28506 13388
rect 28537 13379 28595 13385
rect 28537 13345 28549 13379
rect 28583 13345 28595 13379
rect 28644 13376 28672 13484
rect 28721 13481 28733 13515
rect 28767 13512 28779 13515
rect 28767 13484 29224 13512
rect 28767 13481 28779 13484
rect 28721 13475 28779 13481
rect 28994 13453 29000 13456
rect 28981 13447 29000 13453
rect 28981 13413 28993 13447
rect 28981 13407 29000 13413
rect 28994 13404 29000 13407
rect 29052 13404 29058 13456
rect 29196 13453 29224 13484
rect 29181 13447 29239 13453
rect 29181 13413 29193 13447
rect 29227 13413 29239 13447
rect 29181 13407 29239 13413
rect 29362 13404 29368 13456
rect 29420 13444 29426 13456
rect 30098 13444 30104 13456
rect 29420 13416 30104 13444
rect 29420 13404 29426 13416
rect 29638 13376 29644 13388
rect 28644 13348 29644 13376
rect 28537 13339 28595 13345
rect 25832 13280 26464 13308
rect 25832 13268 25838 13280
rect 26786 13268 26792 13320
rect 26844 13268 26850 13320
rect 28261 13311 28319 13317
rect 28261 13308 28273 13311
rect 26889 13280 28273 13308
rect 24136 13212 24348 13240
rect 14148 13144 16252 13172
rect 14148 13132 14154 13144
rect 16298 13132 16304 13184
rect 16356 13132 16362 13184
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 16448 13144 19257 13172
rect 16448 13132 16454 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19978 13172 19984 13184
rect 19576 13144 19984 13172
rect 19576 13132 19582 13144
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20070 13132 20076 13184
rect 20128 13172 20134 13184
rect 20438 13172 20444 13184
rect 20128 13144 20444 13172
rect 20128 13132 20134 13144
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 21269 13175 21327 13181
rect 21269 13172 21281 13175
rect 20680 13144 21281 13172
rect 20680 13132 20686 13144
rect 21269 13141 21281 13144
rect 21315 13141 21327 13175
rect 21269 13135 21327 13141
rect 22186 13132 22192 13184
rect 22244 13172 22250 13184
rect 24136 13172 24164 13212
rect 24670 13200 24676 13252
rect 24728 13200 24734 13252
rect 24949 13243 25007 13249
rect 24949 13209 24961 13243
rect 24995 13240 25007 13243
rect 24995 13212 26188 13240
rect 24995 13209 25007 13212
rect 24949 13203 25007 13209
rect 26160 13184 26188 13212
rect 26234 13200 26240 13252
rect 26292 13240 26298 13252
rect 26889 13240 26917 13280
rect 28261 13277 28273 13280
rect 28307 13277 28319 13311
rect 28552 13308 28580 13339
rect 29638 13336 29644 13348
rect 29696 13336 29702 13388
rect 29840 13385 29868 13416
rect 30098 13404 30104 13416
rect 30156 13404 30162 13456
rect 29825 13379 29883 13385
rect 29825 13345 29837 13379
rect 29871 13345 29883 13379
rect 29825 13339 29883 13345
rect 30009 13379 30067 13385
rect 30009 13345 30021 13379
rect 30055 13345 30067 13379
rect 30009 13339 30067 13345
rect 28718 13308 28724 13320
rect 28552 13280 28724 13308
rect 28261 13271 28319 13277
rect 27890 13240 27896 13252
rect 26292 13212 26917 13240
rect 26961 13212 27896 13240
rect 26292 13200 26298 13212
rect 22244 13144 24164 13172
rect 22244 13132 22250 13144
rect 24210 13132 24216 13184
rect 24268 13132 24274 13184
rect 24302 13132 24308 13184
rect 24360 13172 24366 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24360 13144 24593 13172
rect 24360 13132 24366 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 26142 13132 26148 13184
rect 26200 13132 26206 13184
rect 26326 13132 26332 13184
rect 26384 13172 26390 13184
rect 26961 13172 26989 13212
rect 27890 13200 27896 13212
rect 27948 13200 27954 13252
rect 28276 13240 28304 13271
rect 28718 13268 28724 13280
rect 28776 13268 28782 13320
rect 28902 13268 28908 13320
rect 28960 13308 28966 13320
rect 30024 13308 30052 13339
rect 30834 13308 30840 13320
rect 28960 13280 30840 13308
rect 28960 13268 28966 13280
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 29546 13240 29552 13252
rect 28276 13212 29552 13240
rect 29546 13200 29552 13212
rect 29604 13200 29610 13252
rect 26384 13144 26989 13172
rect 27157 13175 27215 13181
rect 26384 13132 26390 13144
rect 27157 13141 27169 13175
rect 27203 13172 27215 13175
rect 27430 13172 27436 13184
rect 27203 13144 27436 13172
rect 27203 13141 27215 13144
rect 27157 13135 27215 13141
rect 27430 13132 27436 13144
rect 27488 13132 27494 13184
rect 27982 13132 27988 13184
rect 28040 13172 28046 13184
rect 28813 13175 28871 13181
rect 28813 13172 28825 13175
rect 28040 13144 28825 13172
rect 28040 13132 28046 13144
rect 28813 13141 28825 13144
rect 28859 13141 28871 13175
rect 28813 13135 28871 13141
rect 28997 13175 29055 13181
rect 28997 13141 29009 13175
rect 29043 13172 29055 13175
rect 29086 13172 29092 13184
rect 29043 13144 29092 13172
rect 29043 13141 29055 13144
rect 28997 13135 29055 13141
rect 29086 13132 29092 13144
rect 29144 13132 29150 13184
rect 29914 13132 29920 13184
rect 29972 13132 29978 13184
rect 552 13082 31648 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 11436 13082
rect 11488 13030 11500 13082
rect 11552 13030 11564 13082
rect 11616 13030 11628 13082
rect 11680 13030 11692 13082
rect 11744 13030 19210 13082
rect 19262 13030 19274 13082
rect 19326 13030 19338 13082
rect 19390 13030 19402 13082
rect 19454 13030 19466 13082
rect 19518 13030 26984 13082
rect 27036 13030 27048 13082
rect 27100 13030 27112 13082
rect 27164 13030 27176 13082
rect 27228 13030 27240 13082
rect 27292 13030 31648 13082
rect 552 13008 31648 13030
rect 2498 12928 2504 12980
rect 2556 12968 2562 12980
rect 2866 12968 2872 12980
rect 2556 12940 2872 12968
rect 2556 12928 2562 12940
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 5166 12968 5172 12980
rect 4479 12940 5172 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3142 12900 3148 12912
rect 2832 12872 3148 12900
rect 2832 12860 2838 12872
rect 3142 12860 3148 12872
rect 3200 12900 3206 12912
rect 4448 12900 4476 12931
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12968 5687 12971
rect 6546 12968 6552 12980
rect 5675 12940 6552 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 6730 12928 6736 12980
rect 6788 12928 6794 12980
rect 6822 12928 6828 12980
rect 6880 12928 6886 12980
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7466 12968 7472 12980
rect 7248 12940 7472 12968
rect 7248 12928 7254 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 8021 12971 8079 12977
rect 8021 12968 8033 12971
rect 7800 12940 8033 12968
rect 7800 12928 7806 12940
rect 8021 12937 8033 12940
rect 8067 12937 8079 12971
rect 8021 12931 8079 12937
rect 8110 12928 8116 12980
rect 8168 12968 8174 12980
rect 8168 12940 8800 12968
rect 8168 12928 8174 12940
rect 3200 12872 4476 12900
rect 4617 12903 4675 12909
rect 3200 12860 3206 12872
rect 4617 12869 4629 12903
rect 4663 12869 4675 12903
rect 6840 12900 6868 12928
rect 8772 12912 8800 12940
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 11606 12968 11612 12980
rect 8996 12940 11612 12968
rect 8996 12928 9002 12940
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12158 12968 12164 12980
rect 11722 12940 12164 12968
rect 7006 12900 7012 12912
rect 4617 12863 4675 12869
rect 6748 12872 6868 12900
rect 6932 12872 7012 12900
rect 1946 12792 1952 12844
rect 2004 12832 2010 12844
rect 4154 12832 4160 12844
rect 2004 12804 4160 12832
rect 2004 12792 2010 12804
rect 4154 12792 4160 12804
rect 4212 12832 4218 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4212 12804 4353 12832
rect 4212 12792 4218 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4632 12832 4660 12863
rect 4632 12804 5672 12832
rect 4341 12795 4399 12801
rect 2130 12724 2136 12776
rect 2188 12764 2194 12776
rect 2590 12764 2596 12776
rect 2188 12736 2596 12764
rect 2188 12724 2194 12736
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 4522 12764 4528 12776
rect 4295 12736 4528 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 4614 12724 4620 12776
rect 4672 12764 4678 12776
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4672 12736 4721 12764
rect 4672 12724 4678 12736
rect 4709 12733 4721 12736
rect 4755 12764 4767 12767
rect 4798 12764 4804 12776
rect 4755 12736 4804 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5074 12764 5080 12776
rect 5031 12736 5080 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 5442 12764 5448 12776
rect 5316 12736 5448 12764
rect 5316 12724 5322 12736
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5644 12773 5672 12804
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 5960 12804 6224 12832
rect 5960 12792 5966 12804
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 3568 12600 4813 12628
rect 3568 12588 3574 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 5258 12588 5264 12640
rect 5316 12588 5322 12640
rect 5552 12628 5580 12727
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 6052 12736 6101 12764
rect 6052 12724 6058 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6196 12764 6224 12804
rect 6270 12792 6276 12844
rect 6328 12792 6334 12844
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 6748 12832 6776 12872
rect 6932 12841 6960 12872
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 7377 12903 7435 12909
rect 7377 12869 7389 12903
rect 7423 12900 7435 12903
rect 8202 12900 8208 12912
rect 7423 12872 8208 12900
rect 7423 12869 7435 12872
rect 7377 12863 7435 12869
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 8478 12860 8484 12912
rect 8536 12900 8542 12912
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 8536 12872 8677 12900
rect 8536 12860 8542 12872
rect 8665 12869 8677 12872
rect 8711 12869 8723 12903
rect 8665 12863 8723 12869
rect 8754 12860 8760 12912
rect 8812 12860 8818 12912
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12900 10195 12903
rect 10226 12900 10232 12912
rect 10183 12872 10232 12900
rect 10183 12869 10195 12872
rect 10137 12863 10195 12869
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10962 12860 10968 12912
rect 11020 12900 11026 12912
rect 11722 12900 11750 12940
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 13173 12971 13231 12977
rect 13173 12968 13185 12971
rect 12400 12940 13185 12968
rect 12400 12928 12406 12940
rect 13173 12937 13185 12940
rect 13219 12937 13231 12971
rect 13173 12931 13231 12937
rect 13722 12928 13728 12980
rect 13780 12928 13786 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 16390 12968 16396 12980
rect 13872 12940 16396 12968
rect 13872 12928 13878 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 16758 12968 16764 12980
rect 16715 12940 16764 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 16868 12940 17325 12968
rect 12529 12903 12587 12909
rect 11020 12872 11750 12900
rect 11896 12872 12480 12900
rect 11020 12860 11026 12872
rect 6503 12804 6776 12832
rect 6917 12835 6975 12841
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 6917 12801 6929 12835
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 7147 12804 8401 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 9306 12832 9312 12844
rect 8389 12795 8447 12801
rect 8588 12804 9312 12832
rect 6380 12764 6408 12795
rect 6196 12736 6408 12764
rect 6089 12727 6147 12733
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 6822 12724 6828 12776
rect 6880 12758 6886 12776
rect 7008 12767 7066 12773
rect 7008 12758 7020 12767
rect 6880 12733 7020 12758
rect 7054 12733 7066 12767
rect 6880 12730 7066 12733
rect 6880 12724 6886 12730
rect 7008 12727 7066 12730
rect 7193 12767 7251 12773
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 6178 12656 6184 12708
rect 6236 12696 6242 12708
rect 7208 12696 7236 12727
rect 7926 12724 7932 12776
rect 7984 12724 7990 12776
rect 8018 12724 8024 12776
rect 8076 12764 8082 12776
rect 8588 12773 8616 12804
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 8076 12736 8125 12764
rect 8076 12724 8082 12736
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 8573 12767 8631 12773
rect 8113 12727 8171 12733
rect 8266 12736 8524 12764
rect 6236 12668 7236 12696
rect 6236 12656 6242 12668
rect 8266 12628 8294 12736
rect 8496 12696 8524 12736
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 8573 12727 8631 12733
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 8849 12767 8907 12773
rect 8849 12764 8861 12767
rect 8812 12736 8861 12764
rect 8812 12724 8818 12736
rect 8849 12733 8861 12736
rect 8895 12733 8907 12767
rect 8849 12727 8907 12733
rect 9122 12696 9128 12708
rect 8496 12668 9128 12696
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 9232 12640 9260 12804
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10502 12832 10508 12844
rect 10367 12804 10508 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10502 12792 10508 12804
rect 10560 12832 10566 12844
rect 11896 12832 11924 12872
rect 10560 12804 11924 12832
rect 12452 12832 12480 12872
rect 12529 12869 12541 12903
rect 12575 12900 12587 12903
rect 12618 12900 12624 12912
rect 12575 12872 12624 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 12713 12903 12771 12909
rect 12713 12869 12725 12903
rect 12759 12900 12771 12903
rect 14829 12903 14887 12909
rect 14829 12900 14841 12903
rect 12759 12872 14841 12900
rect 12759 12869 12771 12872
rect 12713 12863 12771 12869
rect 14829 12869 14841 12872
rect 14875 12869 14887 12903
rect 15654 12900 15660 12912
rect 14829 12863 14887 12869
rect 15120 12872 15660 12900
rect 12452 12804 12560 12832
rect 10560 12792 10566 12804
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10410 12764 10416 12776
rect 10183 12736 10416 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 11431 12767 11489 12773
rect 11431 12733 11443 12767
rect 11477 12733 11489 12767
rect 11431 12727 11489 12733
rect 11609 12767 11667 12773
rect 11609 12733 11621 12767
rect 11655 12764 11667 12767
rect 12253 12767 12311 12773
rect 11655 12762 11750 12764
rect 11655 12736 11920 12762
rect 11655 12733 11667 12736
rect 11722 12734 11920 12736
rect 11609 12727 11667 12733
rect 9769 12699 9827 12705
rect 9769 12665 9781 12699
rect 9815 12696 9827 12699
rect 10686 12696 10692 12708
rect 9815 12668 10692 12696
rect 9815 12665 9827 12668
rect 9769 12659 9827 12665
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 11330 12656 11336 12708
rect 11388 12696 11394 12708
rect 11446 12696 11474 12727
rect 11892 12696 11920 12734
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12532 12764 12560 12804
rect 12820 12804 13400 12832
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 12532 12736 12633 12764
rect 12621 12733 12633 12736
rect 12667 12764 12679 12767
rect 12710 12764 12716 12776
rect 12667 12736 12716 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 12820 12773 12848 12804
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12989 12767 13047 12773
rect 12989 12733 13001 12767
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 12894 12696 12900 12708
rect 11388 12668 11652 12696
rect 11892 12668 12900 12696
rect 11388 12656 11394 12668
rect 5552 12600 8294 12628
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 11514 12588 11520 12640
rect 11572 12588 11578 12640
rect 11624 12628 11652 12668
rect 12894 12656 12900 12668
rect 12952 12696 12958 12708
rect 13004 12696 13032 12727
rect 12952 12668 13032 12696
rect 13096 12696 13124 12727
rect 13262 12724 13268 12776
rect 13320 12724 13326 12776
rect 13372 12764 13400 12804
rect 13630 12792 13636 12844
rect 13688 12792 13694 12844
rect 15120 12832 15148 12872
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 15028 12804 15148 12832
rect 15197 12835 15255 12841
rect 13722 12764 13728 12776
rect 13372 12736 13728 12764
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12764 13967 12767
rect 14274 12764 14280 12776
rect 13955 12736 14280 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 15028 12773 15056 12804
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15838 12832 15844 12844
rect 15243 12804 15844 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 15102 12724 15108 12776
rect 15160 12764 15166 12776
rect 15286 12764 15292 12776
rect 15160 12736 15292 12764
rect 15160 12724 15166 12736
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15381 12767 15439 12773
rect 15381 12733 15393 12767
rect 15427 12764 15439 12767
rect 15470 12764 15476 12776
rect 15427 12736 15476 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 15654 12764 15660 12776
rect 15611 12736 15660 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 13354 12696 13360 12708
rect 13096 12668 13360 12696
rect 12952 12656 12958 12668
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 11790 12628 11796 12640
rect 11624 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12628 11854 12640
rect 15580 12628 15608 12727
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 16868 12773 16896 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 17313 12931 17371 12937
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17552 12940 18184 12968
rect 17552 12928 17558 12940
rect 17218 12900 17224 12912
rect 16960 12872 17224 12900
rect 16960 12773 16988 12872
rect 17218 12860 17224 12872
rect 17276 12900 17282 12912
rect 17957 12903 18015 12909
rect 17957 12900 17969 12903
rect 17276 12872 17969 12900
rect 17276 12860 17282 12872
rect 17957 12869 17969 12872
rect 18003 12869 18015 12903
rect 17957 12863 18015 12869
rect 18156 12832 18184 12940
rect 18782 12928 18788 12980
rect 18840 12968 18846 12980
rect 20162 12968 20168 12980
rect 18840 12940 20168 12968
rect 18840 12928 18846 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20806 12928 20812 12980
rect 20864 12928 20870 12980
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 22646 12928 22652 12980
rect 22704 12928 22710 12980
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 23106 12968 23112 12980
rect 22787 12940 23112 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 23106 12928 23112 12940
rect 23164 12928 23170 12980
rect 24136 12940 28764 12968
rect 18230 12860 18236 12912
rect 18288 12900 18294 12912
rect 18969 12903 19027 12909
rect 18969 12900 18981 12903
rect 18288 12872 18981 12900
rect 18288 12860 18294 12872
rect 18969 12869 18981 12872
rect 19015 12869 19027 12903
rect 20824 12900 20852 12928
rect 18969 12863 19027 12869
rect 19720 12872 20852 12900
rect 22925 12903 22983 12909
rect 18325 12835 18383 12841
rect 17144 12804 17724 12832
rect 18156 12804 18276 12832
rect 17144 12773 17172 12804
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 17310 12764 17316 12776
rect 17267 12736 17316 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17497 12767 17555 12773
rect 17497 12733 17509 12767
rect 17543 12733 17555 12767
rect 17497 12727 17555 12733
rect 17034 12656 17040 12708
rect 17092 12696 17098 12708
rect 17512 12696 17540 12727
rect 17092 12668 17540 12696
rect 17092 12656 17098 12668
rect 11848 12600 15608 12628
rect 11848 12588 11854 12600
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 17218 12628 17224 12640
rect 15988 12600 17224 12628
rect 15988 12588 15994 12600
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17696 12628 17724 12804
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17828 12736 17877 12764
rect 17828 12724 17834 12736
rect 17865 12733 17877 12736
rect 17911 12733 17923 12767
rect 17865 12727 17923 12733
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18141 12767 18199 12773
rect 18141 12764 18153 12767
rect 18012 12736 18153 12764
rect 18012 12724 18018 12736
rect 18141 12733 18153 12736
rect 18187 12733 18199 12767
rect 18248 12764 18276 12804
rect 18325 12801 18337 12835
rect 18371 12832 18383 12835
rect 19337 12835 19395 12841
rect 19337 12832 19349 12835
rect 18371 12804 19349 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 19337 12801 19349 12804
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19720 12832 19748 12872
rect 22925 12869 22937 12903
rect 22971 12900 22983 12903
rect 24136 12900 24164 12940
rect 22971 12872 24164 12900
rect 24432 12872 27108 12900
rect 22971 12869 22983 12872
rect 22925 12863 22983 12869
rect 20714 12832 20720 12844
rect 19484 12804 19748 12832
rect 19484 12792 19490 12804
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 18248 12736 18429 12764
rect 18141 12727 18199 12733
rect 18417 12733 18429 12736
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12733 18935 12767
rect 18877 12727 18935 12733
rect 18892 12696 18920 12727
rect 19150 12724 19156 12776
rect 19208 12724 19214 12776
rect 19720 12773 19748 12804
rect 19996 12804 20720 12832
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19460 12736 19625 12764
rect 18432 12668 18920 12696
rect 19168 12696 19196 12724
rect 19334 12696 19340 12708
rect 19168 12668 19340 12696
rect 18432 12640 18460 12668
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 17770 12628 17776 12640
rect 17696 12600 17776 12628
rect 17770 12588 17776 12600
rect 17828 12588 17834 12640
rect 18414 12588 18420 12640
rect 18472 12588 18478 12640
rect 19460 12628 19488 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 19794 12724 19800 12776
rect 19852 12724 19858 12776
rect 19996 12773 20024 12804
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 22094 12832 22100 12844
rect 20855 12804 22100 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22646 12792 22652 12844
rect 22704 12832 22710 12844
rect 22741 12835 22799 12841
rect 22741 12832 22753 12835
rect 22704 12804 22753 12832
rect 22704 12792 22710 12804
rect 22741 12801 22753 12804
rect 22787 12801 22799 12835
rect 22741 12795 22799 12801
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 23198 12832 23204 12844
rect 22888 12804 23204 12832
rect 22888 12792 22894 12804
rect 23198 12792 23204 12804
rect 23256 12792 23262 12844
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20312 12736 20453 12764
rect 20312 12724 20318 12736
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 20441 12727 20499 12733
rect 20901 12767 20959 12773
rect 20901 12733 20913 12767
rect 20947 12764 20959 12767
rect 21910 12764 21916 12776
rect 20947 12736 21916 12764
rect 20947 12733 20959 12736
rect 20901 12727 20959 12733
rect 21910 12724 21916 12736
rect 21968 12764 21974 12776
rect 22557 12767 22615 12773
rect 22557 12764 22569 12767
rect 21968 12736 22569 12764
rect 21968 12724 21974 12736
rect 22557 12733 22569 12736
rect 22603 12733 22615 12767
rect 22557 12727 22615 12733
rect 24026 12724 24032 12776
rect 24084 12724 24090 12776
rect 24121 12767 24179 12773
rect 24121 12733 24133 12767
rect 24167 12764 24179 12767
rect 24432 12764 24460 12872
rect 24670 12792 24676 12844
rect 24728 12832 24734 12844
rect 24857 12835 24915 12841
rect 24857 12832 24869 12835
rect 24728 12804 24869 12832
rect 24728 12792 24734 12804
rect 24857 12801 24869 12804
rect 24903 12801 24915 12835
rect 26142 12832 26148 12844
rect 24857 12795 24915 12801
rect 24964 12804 26148 12832
rect 24167 12736 24460 12764
rect 24489 12767 24547 12773
rect 24167 12733 24179 12736
rect 24121 12727 24179 12733
rect 24489 12733 24501 12767
rect 24535 12764 24547 12767
rect 24578 12764 24584 12776
rect 24535 12736 24584 12764
rect 24535 12733 24547 12736
rect 24489 12727 24547 12733
rect 24578 12724 24584 12736
rect 24636 12724 24642 12776
rect 24964 12773 24992 12804
rect 26142 12792 26148 12804
rect 26200 12832 26206 12844
rect 26329 12835 26387 12841
rect 26329 12832 26341 12835
rect 26200 12804 26341 12832
rect 26200 12792 26206 12804
rect 26329 12801 26341 12804
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 26510 12792 26516 12844
rect 26568 12832 26574 12844
rect 26970 12832 26976 12844
rect 26568 12804 26976 12832
rect 26568 12792 26574 12804
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27080 12832 27108 12872
rect 27154 12860 27160 12912
rect 27212 12900 27218 12912
rect 27706 12900 27712 12912
rect 27212 12872 27712 12900
rect 27212 12860 27218 12872
rect 27706 12860 27712 12872
rect 27764 12860 27770 12912
rect 28736 12900 28764 12940
rect 28994 12928 29000 12980
rect 29052 12928 29058 12980
rect 29104 12940 29316 12968
rect 29104 12900 29132 12940
rect 28736 12872 29132 12900
rect 29288 12900 29316 12940
rect 29362 12928 29368 12980
rect 29420 12928 29426 12980
rect 29825 12903 29883 12909
rect 29825 12900 29837 12903
rect 29288 12872 29837 12900
rect 29825 12869 29837 12872
rect 29871 12869 29883 12903
rect 29825 12863 29883 12869
rect 29914 12860 29920 12912
rect 29972 12860 29978 12912
rect 30285 12835 30343 12841
rect 30285 12832 30297 12835
rect 27080 12804 30297 12832
rect 30285 12801 30297 12804
rect 30331 12832 30343 12835
rect 30377 12835 30435 12841
rect 30377 12832 30389 12835
rect 30331 12804 30389 12832
rect 30331 12801 30343 12804
rect 30285 12795 30343 12801
rect 30377 12801 30389 12804
rect 30423 12801 30435 12835
rect 30377 12795 30435 12801
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12733 24823 12767
rect 24765 12727 24823 12733
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12733 25007 12767
rect 26421 12767 26479 12773
rect 26421 12764 26433 12767
rect 24949 12727 25007 12733
rect 26344 12736 26433 12764
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19576 12668 20760 12696
rect 19576 12656 19582 12668
rect 19978 12628 19984 12640
rect 19460 12600 19984 12628
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 20732 12637 20760 12668
rect 22002 12656 22008 12708
rect 22060 12696 22066 12708
rect 22060 12668 24164 12696
rect 22060 12656 22066 12668
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 20404 12600 20545 12628
rect 20404 12588 20410 12600
rect 20533 12597 20545 12600
rect 20579 12597 20591 12631
rect 20533 12591 20591 12597
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 20898 12628 20904 12640
rect 20763 12600 20904 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 21818 12588 21824 12640
rect 21876 12628 21882 12640
rect 23845 12631 23903 12637
rect 23845 12628 23857 12631
rect 21876 12600 23857 12628
rect 21876 12588 21882 12600
rect 23845 12597 23857 12600
rect 23891 12597 23903 12631
rect 24136 12628 24164 12668
rect 24210 12656 24216 12708
rect 24268 12656 24274 12708
rect 24302 12656 24308 12708
rect 24360 12705 24366 12708
rect 24360 12699 24389 12705
rect 24377 12665 24389 12699
rect 24780 12696 24808 12727
rect 25130 12696 25136 12708
rect 24780 12668 25136 12696
rect 24360 12659 24389 12665
rect 24360 12656 24366 12659
rect 25130 12656 25136 12668
rect 25188 12696 25194 12708
rect 26142 12696 26148 12708
rect 25188 12668 26148 12696
rect 25188 12656 25194 12668
rect 26142 12656 26148 12668
rect 26200 12656 26206 12708
rect 26344 12628 26372 12736
rect 26421 12733 26433 12736
rect 26467 12764 26479 12767
rect 26467 12736 26917 12764
rect 26467 12733 26479 12736
rect 26421 12727 26479 12733
rect 26694 12656 26700 12708
rect 26752 12696 26758 12708
rect 26752 12668 26832 12696
rect 26752 12656 26758 12668
rect 26804 12637 26832 12668
rect 24136 12600 26372 12628
rect 26789 12631 26847 12637
rect 23845 12591 23903 12597
rect 26789 12597 26801 12631
rect 26835 12597 26847 12631
rect 26889 12628 26917 12736
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28626 12764 28632 12776
rect 27856 12736 28632 12764
rect 27856 12724 27862 12736
rect 28626 12724 28632 12736
rect 28684 12724 28690 12776
rect 28718 12724 28724 12776
rect 28776 12764 28782 12776
rect 28776 12736 29132 12764
rect 28776 12724 28782 12736
rect 29104 12696 29132 12736
rect 29178 12724 29184 12776
rect 29236 12724 29242 12776
rect 29273 12767 29331 12773
rect 29273 12733 29285 12767
rect 29319 12733 29331 12767
rect 29273 12727 29331 12733
rect 30561 12767 30619 12773
rect 30561 12733 30573 12767
rect 30607 12764 30619 12767
rect 30742 12764 30748 12776
rect 30607 12736 30748 12764
rect 30607 12733 30619 12736
rect 30561 12727 30619 12733
rect 29288 12696 29316 12727
rect 30742 12724 30748 12736
rect 30800 12724 30806 12776
rect 30834 12724 30840 12776
rect 30892 12724 30898 12776
rect 29104 12668 29316 12696
rect 29638 12656 29644 12708
rect 29696 12656 29702 12708
rect 30745 12631 30803 12637
rect 30745 12628 30757 12631
rect 26889 12600 30757 12628
rect 26789 12591 26847 12597
rect 30745 12597 30757 12600
rect 30791 12628 30803 12631
rect 31570 12628 31576 12640
rect 30791 12600 31576 12628
rect 30791 12597 30803 12600
rect 30745 12591 30803 12597
rect 31570 12588 31576 12600
rect 31628 12588 31634 12640
rect 552 12538 31648 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 12096 12538
rect 12148 12486 12160 12538
rect 12212 12486 12224 12538
rect 12276 12486 12288 12538
rect 12340 12486 12352 12538
rect 12404 12486 19870 12538
rect 19922 12486 19934 12538
rect 19986 12486 19998 12538
rect 20050 12486 20062 12538
rect 20114 12486 20126 12538
rect 20178 12486 27644 12538
rect 27696 12486 27708 12538
rect 27760 12486 27772 12538
rect 27824 12486 27836 12538
rect 27888 12486 27900 12538
rect 27952 12486 31648 12538
rect 552 12464 31648 12486
rect 1765 12427 1823 12433
rect 1765 12393 1777 12427
rect 1811 12424 1823 12427
rect 1854 12424 1860 12436
rect 1811 12396 1860 12424
rect 1811 12393 1823 12396
rect 1765 12387 1823 12393
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 3237 12427 3295 12433
rect 3237 12393 3249 12427
rect 3283 12424 3295 12427
rect 3418 12424 3424 12436
rect 3283 12396 3424 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4985 12427 5043 12433
rect 4985 12393 4997 12427
rect 5031 12424 5043 12427
rect 5166 12424 5172 12436
rect 5031 12396 5172 12424
rect 5031 12393 5043 12396
rect 4985 12387 5043 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 6178 12424 6184 12436
rect 5500 12396 6184 12424
rect 5500 12384 5506 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6822 12384 6828 12436
rect 6880 12384 6886 12436
rect 7558 12384 7564 12436
rect 7616 12384 7622 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 8570 12424 8576 12436
rect 7984 12396 8576 12424
rect 7984 12384 7990 12396
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 9088 12396 9137 12424
rect 9088 12384 9094 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9824 12396 9873 12424
rect 9824 12384 9830 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 9861 12387 9919 12393
rect 9968 12396 12204 12424
rect 1118 12316 1124 12368
rect 1176 12356 1182 12368
rect 1581 12359 1639 12365
rect 1581 12356 1593 12359
rect 1176 12328 1593 12356
rect 1176 12316 1182 12328
rect 1581 12325 1593 12328
rect 1627 12356 1639 12359
rect 1946 12356 1952 12368
rect 1627 12328 1952 12356
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 1946 12316 1952 12328
rect 2004 12316 2010 12368
rect 4706 12356 4712 12368
rect 3896 12328 4712 12356
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1544 12260 1869 12288
rect 1544 12248 1550 12260
rect 1857 12257 1869 12260
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 2038 12248 2044 12300
rect 2096 12288 2102 12300
rect 3418 12288 3424 12300
rect 2096 12260 3424 12288
rect 2096 12248 2102 12260
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 3510 12248 3516 12300
rect 3568 12248 3574 12300
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 3896 12297 3924 12328
rect 4706 12316 4712 12328
rect 4764 12356 4770 12368
rect 4801 12359 4859 12365
rect 4801 12356 4813 12359
rect 4764 12328 4813 12356
rect 4764 12316 4770 12328
rect 4801 12325 4813 12328
rect 4847 12356 4859 12359
rect 5626 12356 5632 12368
rect 4847 12328 5632 12356
rect 4847 12325 4859 12328
rect 4801 12319 4859 12325
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 7098 12316 7104 12368
rect 7156 12316 7162 12368
rect 7576 12356 7604 12384
rect 8478 12356 8484 12368
rect 7576 12328 8484 12356
rect 8478 12316 8484 12328
rect 8536 12356 8542 12368
rect 9968 12356 9996 12396
rect 10686 12356 10692 12368
rect 8536 12328 9996 12356
rect 10060 12328 10692 12356
rect 8536 12316 8542 12328
rect 3697 12291 3755 12297
rect 3697 12288 3709 12291
rect 3660 12260 3709 12288
rect 3660 12248 3666 12260
rect 3697 12257 3709 12260
rect 3743 12257 3755 12291
rect 3697 12251 3755 12257
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12257 3939 12291
rect 3881 12251 3939 12257
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5258 12288 5264 12300
rect 5123 12260 5264 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 7009 12291 7067 12297
rect 7009 12257 7021 12291
rect 7055 12288 7067 12291
rect 7116 12288 7144 12316
rect 7055 12260 7144 12288
rect 7055 12257 7067 12260
rect 7009 12251 7067 12257
rect 7190 12248 7196 12300
rect 7248 12248 7254 12300
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 3528 12152 3556 12248
rect 5994 12220 6000 12232
rect 3620 12192 6000 12220
rect 3620 12161 3648 12192
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 7098 12180 7104 12232
rect 7156 12180 7162 12232
rect 7300 12220 7328 12251
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 8754 12288 8760 12300
rect 8444 12260 8760 12288
rect 8444 12248 8450 12260
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9214 12248 9220 12300
rect 9272 12288 9278 12300
rect 10060 12297 10088 12328
rect 10686 12316 10692 12328
rect 10744 12316 10750 12368
rect 10962 12316 10968 12368
rect 11020 12356 11026 12368
rect 12066 12356 12072 12368
rect 11020 12328 12072 12356
rect 11020 12316 11026 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 9272 12260 9321 12288
rect 9272 12248 9278 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9309 12251 9367 12257
rect 9404 12260 9597 12288
rect 9404 12220 9432 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 7300 12192 7788 12220
rect 1627 12124 3556 12152
rect 3605 12155 3663 12161
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 3605 12121 3617 12155
rect 3651 12121 3663 12155
rect 3605 12115 3663 12121
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4522 12152 4528 12164
rect 4212 12124 4528 12152
rect 4212 12112 4218 12124
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 4798 12112 4804 12164
rect 4856 12112 4862 12164
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 6546 12152 6552 12164
rect 5132 12124 6552 12152
rect 5132 12112 5138 12124
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 7760 12096 7788 12192
rect 8496 12192 9432 12220
rect 2222 12044 2228 12096
rect 2280 12084 2286 12096
rect 4430 12084 4436 12096
rect 2280 12056 4436 12084
rect 2280 12044 2286 12056
rect 4430 12044 4436 12056
rect 4488 12084 4494 12096
rect 4890 12084 4896 12096
rect 4488 12056 4896 12084
rect 4488 12044 4494 12056
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 6454 12084 6460 12096
rect 5224 12056 6460 12084
rect 5224 12044 5230 12056
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 7742 12044 7748 12096
rect 7800 12044 7806 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8496 12084 8524 12192
rect 9490 12180 9496 12232
rect 9548 12180 9554 12232
rect 9784 12220 9812 12251
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10192 12260 10517 12288
rect 10192 12248 10198 12260
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 11514 12288 11520 12300
rect 10505 12251 10563 12257
rect 10980 12260 11520 12288
rect 10152 12220 10180 12248
rect 9784 12192 10180 12220
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10870 12220 10876 12232
rect 10367 12192 10876 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 9214 12152 9220 12164
rect 8628 12124 9220 12152
rect 8628 12112 8634 12124
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 9398 12112 9404 12164
rect 9456 12112 9462 12164
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10502 12152 10508 12164
rect 10192 12124 10508 12152
rect 10192 12112 10198 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 10980 12152 11008 12260
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 12176 12297 12204 12396
rect 12986 12384 12992 12436
rect 13044 12384 13050 12436
rect 13354 12384 13360 12436
rect 13412 12384 13418 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 12437 12359 12495 12365
rect 12437 12325 12449 12359
rect 12483 12356 12495 12359
rect 13372 12356 13400 12384
rect 12483 12328 13400 12356
rect 13475 12359 13533 12365
rect 12483 12325 12495 12328
rect 12437 12319 12495 12325
rect 13475 12325 13487 12359
rect 13521 12356 13533 12359
rect 13740 12356 13768 12387
rect 15010 12384 15016 12436
rect 15068 12384 15074 12436
rect 17402 12384 17408 12436
rect 17460 12424 17466 12436
rect 18138 12424 18144 12436
rect 17460 12396 18144 12424
rect 17460 12384 17466 12396
rect 18138 12384 18144 12396
rect 18196 12424 18202 12436
rect 18233 12427 18291 12433
rect 18233 12424 18245 12427
rect 18196 12396 18245 12424
rect 18196 12384 18202 12396
rect 18233 12393 18245 12396
rect 18279 12393 18291 12427
rect 18233 12387 18291 12393
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 18966 12424 18972 12436
rect 18656 12396 18972 12424
rect 18656 12384 18662 12396
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19242 12384 19248 12436
rect 19300 12424 19306 12436
rect 20346 12424 20352 12436
rect 19300 12396 20352 12424
rect 19300 12384 19306 12396
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 21542 12424 21548 12436
rect 20640 12396 21548 12424
rect 13521 12328 13768 12356
rect 13521 12325 13533 12328
rect 13475 12319 13533 12325
rect 14090 12316 14096 12368
rect 14148 12356 14154 12368
rect 16853 12359 16911 12365
rect 14148 12328 14504 12356
rect 14148 12316 14154 12328
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12894 12288 12900 12300
rect 12207 12260 12900 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13170 12248 13176 12300
rect 13228 12248 13234 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11882 12220 11888 12232
rect 11112 12192 11888 12220
rect 11112 12180 11118 12192
rect 11882 12180 11888 12192
rect 11940 12220 11946 12232
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 11940 12192 12265 12220
rect 11940 12180 11946 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 12437 12223 12495 12229
rect 12437 12220 12449 12223
rect 12400 12192 12449 12220
rect 12400 12180 12406 12192
rect 12437 12189 12449 12192
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13280 12220 13308 12251
rect 13044 12192 13308 12220
rect 13044 12180 13050 12192
rect 10704 12124 11008 12152
rect 7892 12056 8524 12084
rect 7892 12044 7898 12056
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 10226 12084 10232 12096
rect 9548 12056 10232 12084
rect 9548 12044 9554 12056
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 10704 12084 10732 12124
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 11204 12124 11652 12152
rect 11204 12112 11210 12124
rect 10376 12056 10732 12084
rect 10376 12044 10382 12056
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11330 12084 11336 12096
rect 10836 12056 11336 12084
rect 10836 12044 10842 12056
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 11624 12084 11652 12124
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 12894 12152 12900 12164
rect 11756 12124 12900 12152
rect 11756 12112 11762 12124
rect 12894 12112 12900 12124
rect 12952 12152 12958 12164
rect 13372 12152 13400 12251
rect 13630 12248 13636 12300
rect 13688 12248 13694 12300
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13780 12260 14013 12288
rect 13780 12248 13786 12260
rect 14001 12257 14013 12260
rect 14047 12257 14059 12291
rect 14001 12251 14059 12257
rect 14366 12248 14372 12300
rect 14424 12248 14430 12300
rect 14476 12288 14504 12328
rect 16853 12325 16865 12359
rect 16899 12356 16911 12359
rect 20530 12356 20536 12368
rect 16899 12328 20536 12356
rect 16899 12325 16911 12328
rect 16853 12319 16911 12325
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 14532 12291 14590 12297
rect 14532 12288 14544 12291
rect 14476 12260 14544 12288
rect 14532 12257 14544 12260
rect 14578 12257 14590 12291
rect 14532 12251 14590 12257
rect 14645 12291 14703 12297
rect 14645 12257 14657 12291
rect 14691 12257 14703 12291
rect 14645 12251 14703 12257
rect 13538 12180 13544 12232
rect 13596 12220 13602 12232
rect 13740 12220 13768 12248
rect 13596 12192 13768 12220
rect 13596 12180 13602 12192
rect 13906 12180 13912 12232
rect 13964 12180 13970 12232
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 12952 12124 13400 12152
rect 14108 12152 14136 12183
rect 14182 12180 14188 12232
rect 14240 12180 14246 12232
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 14660 12220 14688 12251
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14792 12260 15301 12288
rect 14792 12248 14798 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15488 12220 15516 12251
rect 16666 12248 16672 12300
rect 16724 12248 16730 12300
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 14332 12192 14688 12220
rect 15120 12192 15516 12220
rect 14332 12180 14338 12192
rect 14108 12124 14228 12152
rect 12952 12112 12958 12124
rect 14200 12096 14228 12124
rect 15120 12096 15148 12192
rect 15654 12180 15660 12232
rect 15712 12180 15718 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16960 12220 16988 12251
rect 17034 12248 17040 12300
rect 17092 12248 17098 12300
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17644 12260 17693 12288
rect 17644 12248 17650 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17828 12260 17877 12288
rect 17828 12248 17834 12260
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 18046 12248 18052 12300
rect 18104 12248 18110 12300
rect 18325 12291 18383 12297
rect 18325 12257 18337 12291
rect 18371 12257 18383 12291
rect 18325 12251 18383 12257
rect 15988 12192 16988 12220
rect 15988 12180 15994 12192
rect 15470 12112 15476 12164
rect 15528 12152 15534 12164
rect 15672 12152 15700 12180
rect 15528 12124 15700 12152
rect 15528 12112 15534 12124
rect 12434 12084 12440 12096
rect 11624 12056 12440 12084
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 14182 12044 14188 12096
rect 14240 12044 14246 12096
rect 15102 12044 15108 12096
rect 15160 12044 15166 12096
rect 16960 12084 16988 12192
rect 17402 12180 17408 12232
rect 17460 12220 17466 12232
rect 18340 12220 18368 12251
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 18748 12260 18981 12288
rect 18748 12248 18754 12260
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 19058 12248 19064 12300
rect 19116 12248 19122 12300
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 20640 12288 20668 12396
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 21634 12384 21640 12436
rect 21692 12424 21698 12436
rect 22097 12427 22155 12433
rect 22097 12424 22109 12427
rect 21692 12396 22109 12424
rect 21692 12384 21698 12396
rect 22097 12393 22109 12396
rect 22143 12393 22155 12427
rect 22097 12387 22155 12393
rect 22922 12384 22928 12436
rect 22980 12424 22986 12436
rect 23382 12424 23388 12436
rect 22980 12396 23388 12424
rect 22980 12384 22986 12396
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 23661 12427 23719 12433
rect 23661 12393 23673 12427
rect 23707 12424 23719 12427
rect 24026 12424 24032 12436
rect 23707 12396 24032 12424
rect 23707 12393 23719 12396
rect 23661 12387 23719 12393
rect 24026 12384 24032 12396
rect 24084 12384 24090 12436
rect 25958 12384 25964 12436
rect 26016 12424 26022 12436
rect 26421 12427 26479 12433
rect 26421 12424 26433 12427
rect 26016 12396 26433 12424
rect 26016 12384 26022 12396
rect 26421 12393 26433 12396
rect 26467 12393 26479 12427
rect 26421 12387 26479 12393
rect 26510 12384 26516 12436
rect 26568 12424 26574 12436
rect 26568 12396 26832 12424
rect 26568 12384 26574 12396
rect 22370 12316 22376 12368
rect 22428 12356 22434 12368
rect 22554 12356 22560 12368
rect 22428 12328 22560 12356
rect 22428 12316 22434 12328
rect 22554 12316 22560 12328
rect 22612 12356 22618 12368
rect 22612 12328 23428 12356
rect 22612 12316 22618 12328
rect 19760 12260 20668 12288
rect 19760 12248 19766 12260
rect 21174 12248 21180 12300
rect 21232 12288 21238 12300
rect 21910 12288 21916 12300
rect 21232 12260 21916 12288
rect 21232 12248 21238 12260
rect 21910 12248 21916 12260
rect 21968 12248 21974 12300
rect 22002 12248 22008 12300
rect 22060 12288 22066 12300
rect 22649 12291 22707 12297
rect 22649 12288 22661 12291
rect 22060 12260 22661 12288
rect 22060 12248 22066 12260
rect 22649 12257 22661 12260
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 22738 12248 22744 12300
rect 22796 12288 22802 12300
rect 22922 12288 22928 12300
rect 22796 12260 22928 12288
rect 22796 12248 22802 12260
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 23106 12248 23112 12300
rect 23164 12248 23170 12300
rect 23198 12248 23204 12300
rect 23256 12248 23262 12300
rect 23290 12248 23296 12300
rect 23348 12248 23354 12300
rect 23400 12297 23428 12328
rect 24210 12316 24216 12368
rect 24268 12356 24274 12368
rect 24268 12328 26096 12356
rect 24268 12316 24274 12328
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12257 23443 12291
rect 23385 12251 23443 12257
rect 23566 12248 23572 12300
rect 23624 12288 23630 12300
rect 24397 12291 24455 12297
rect 24397 12288 24409 12291
rect 23624 12260 24409 12288
rect 23624 12248 23630 12260
rect 24397 12257 24409 12260
rect 24443 12257 24455 12291
rect 24397 12251 24455 12257
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 24903 12260 25084 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 17460 12192 18368 12220
rect 17460 12180 17466 12192
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 18656 12192 18828 12220
rect 18656 12180 18662 12192
rect 17221 12155 17279 12161
rect 17221 12121 17233 12155
rect 17267 12152 17279 12155
rect 17494 12152 17500 12164
rect 17267 12124 17500 12152
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 17494 12112 17500 12124
rect 17552 12112 17558 12164
rect 18138 12112 18144 12164
rect 18196 12152 18202 12164
rect 18693 12155 18751 12161
rect 18693 12152 18705 12155
rect 18196 12124 18705 12152
rect 18196 12112 18202 12124
rect 18693 12121 18705 12124
rect 18739 12121 18751 12155
rect 18800 12152 18828 12192
rect 18874 12180 18880 12232
rect 18932 12180 18938 12232
rect 19153 12223 19211 12229
rect 19153 12189 19165 12223
rect 19199 12220 19211 12223
rect 20162 12220 20168 12232
rect 19199 12192 20168 12220
rect 19199 12189 19211 12192
rect 19153 12183 19211 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 20346 12180 20352 12232
rect 20404 12220 20410 12232
rect 22186 12220 22192 12232
rect 20404 12192 22192 12220
rect 20404 12180 20410 12192
rect 22186 12180 22192 12192
rect 22244 12180 22250 12232
rect 22373 12223 22431 12229
rect 22373 12189 22385 12223
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 19242 12152 19248 12164
rect 18800 12124 19248 12152
rect 18693 12115 18751 12121
rect 19242 12112 19248 12124
rect 19300 12112 19306 12164
rect 19334 12112 19340 12164
rect 19392 12152 19398 12164
rect 21450 12152 21456 12164
rect 19392 12124 21456 12152
rect 19392 12112 19398 12124
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 22388 12152 22416 12183
rect 24121 12155 24179 12161
rect 24121 12152 24133 12155
rect 22388 12124 24133 12152
rect 24121 12121 24133 12124
rect 24167 12121 24179 12155
rect 24121 12115 24179 12121
rect 24489 12155 24547 12161
rect 24489 12121 24501 12155
rect 24535 12152 24547 12155
rect 24949 12155 25007 12161
rect 24949 12152 24961 12155
rect 24535 12124 24961 12152
rect 24535 12121 24547 12124
rect 24489 12115 24547 12121
rect 24949 12121 24961 12124
rect 24995 12121 25007 12155
rect 25056 12152 25084 12260
rect 25130 12248 25136 12300
rect 25188 12248 25194 12300
rect 25498 12248 25504 12300
rect 25556 12248 25562 12300
rect 25685 12291 25743 12297
rect 25685 12257 25697 12291
rect 25731 12288 25743 12291
rect 25774 12288 25780 12300
rect 25731 12260 25780 12288
rect 25731 12257 25743 12260
rect 25685 12251 25743 12257
rect 25774 12248 25780 12260
rect 25832 12248 25838 12300
rect 26068 12297 26096 12328
rect 26694 12316 26700 12368
rect 26752 12316 26758 12368
rect 26804 12356 26832 12396
rect 27154 12384 27160 12436
rect 27212 12424 27218 12436
rect 27433 12427 27491 12433
rect 27433 12424 27445 12427
rect 27212 12396 27445 12424
rect 27212 12384 27218 12396
rect 27433 12393 27445 12396
rect 27479 12393 27491 12427
rect 27433 12387 27491 12393
rect 27525 12427 27583 12433
rect 27525 12393 27537 12427
rect 27571 12393 27583 12427
rect 27525 12387 27583 12393
rect 27540 12356 27568 12387
rect 26804 12328 27568 12356
rect 27614 12316 27620 12368
rect 27672 12356 27678 12368
rect 27709 12359 27767 12365
rect 27709 12356 27721 12359
rect 27672 12328 27721 12356
rect 27672 12316 27678 12328
rect 27709 12325 27721 12328
rect 27755 12325 27767 12359
rect 27709 12319 27767 12325
rect 28350 12316 28356 12368
rect 28408 12316 28414 12368
rect 29086 12316 29092 12368
rect 29144 12316 29150 12368
rect 29914 12316 29920 12368
rect 29972 12356 29978 12368
rect 29972 12328 30512 12356
rect 29972 12316 29978 12328
rect 26053 12291 26111 12297
rect 26053 12257 26065 12291
rect 26099 12257 26111 12291
rect 26053 12251 26111 12257
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12220 25467 12223
rect 25593 12223 25651 12229
rect 25593 12220 25605 12223
rect 25455 12192 25605 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 25593 12189 25605 12192
rect 25639 12189 25651 12223
rect 25593 12183 25651 12189
rect 26068 12152 26096 12251
rect 26234 12248 26240 12300
rect 26292 12248 26298 12300
rect 26418 12248 26424 12300
rect 26476 12288 26482 12300
rect 26605 12291 26663 12297
rect 26605 12288 26617 12291
rect 26476 12260 26617 12288
rect 26476 12248 26482 12260
rect 26605 12257 26617 12260
rect 26651 12257 26663 12291
rect 26605 12251 26663 12257
rect 26786 12248 26792 12300
rect 26844 12248 26850 12300
rect 26973 12291 27031 12297
rect 26973 12257 26985 12291
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 26145 12223 26203 12229
rect 26145 12189 26157 12223
rect 26191 12220 26203 12223
rect 26988 12220 27016 12251
rect 27062 12248 27068 12300
rect 27120 12248 27126 12300
rect 27246 12248 27252 12300
rect 27304 12288 27310 12300
rect 27341 12291 27399 12297
rect 27341 12288 27353 12291
rect 27304 12260 27353 12288
rect 27304 12248 27310 12260
rect 27341 12257 27353 12260
rect 27387 12288 27399 12291
rect 27985 12291 28043 12297
rect 27387 12260 27476 12288
rect 27387 12257 27399 12260
rect 27341 12251 27399 12257
rect 26191 12192 27016 12220
rect 26191 12189 26203 12192
rect 26145 12183 26203 12189
rect 27448 12164 27476 12260
rect 27985 12257 27997 12291
rect 28031 12288 28043 12291
rect 28074 12288 28080 12300
rect 28031 12260 28080 12288
rect 28031 12257 28043 12260
rect 27985 12251 28043 12257
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28169 12291 28227 12297
rect 28169 12257 28181 12291
rect 28215 12257 28227 12291
rect 28445 12291 28503 12297
rect 28445 12288 28457 12291
rect 28169 12251 28227 12257
rect 28368 12260 28457 12288
rect 26510 12152 26516 12164
rect 25056 12124 25728 12152
rect 26068 12124 26516 12152
rect 24949 12115 25007 12121
rect 17310 12084 17316 12096
rect 16960 12056 17316 12084
rect 17310 12044 17316 12056
rect 17368 12084 17374 12096
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 17368 12056 17417 12084
rect 17368 12044 17374 12056
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 22094 12084 22100 12096
rect 18564 12056 22100 12084
rect 18564 12044 18570 12056
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22557 12087 22615 12093
rect 22557 12053 22569 12087
rect 22603 12084 22615 12087
rect 22741 12087 22799 12093
rect 22741 12084 22753 12087
rect 22603 12056 22753 12084
rect 22603 12053 22615 12056
rect 22557 12047 22615 12053
rect 22741 12053 22753 12056
rect 22787 12053 22799 12087
rect 22741 12047 22799 12053
rect 23106 12044 23112 12096
rect 23164 12084 23170 12096
rect 23293 12087 23351 12093
rect 23293 12084 23305 12087
rect 23164 12056 23305 12084
rect 23164 12044 23170 12056
rect 23293 12053 23305 12056
rect 23339 12053 23351 12087
rect 23293 12047 23351 12053
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 24581 12087 24639 12093
rect 24581 12084 24593 12087
rect 23624 12056 24593 12084
rect 23624 12044 23630 12056
rect 24581 12053 24593 12056
rect 24627 12053 24639 12087
rect 24581 12047 24639 12053
rect 24673 12087 24731 12093
rect 24673 12053 24685 12087
rect 24719 12084 24731 12087
rect 24854 12084 24860 12096
rect 24719 12056 24860 12084
rect 24719 12053 24731 12056
rect 24673 12047 24731 12053
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 25317 12087 25375 12093
rect 25317 12053 25329 12087
rect 25363 12084 25375 12087
rect 25590 12084 25596 12096
rect 25363 12056 25596 12084
rect 25363 12053 25375 12056
rect 25317 12047 25375 12053
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 25700 12084 25728 12124
rect 26510 12112 26516 12124
rect 26568 12152 26574 12164
rect 27157 12155 27215 12161
rect 27157 12152 27169 12155
rect 26568 12124 27169 12152
rect 26568 12112 26574 12124
rect 27157 12121 27169 12124
rect 27203 12121 27215 12155
rect 27157 12115 27215 12121
rect 27430 12112 27436 12164
rect 27488 12112 27494 12164
rect 28184 12152 28212 12251
rect 28368 12232 28396 12260
rect 28445 12257 28457 12260
rect 28491 12257 28503 12291
rect 28445 12251 28503 12257
rect 28718 12248 28724 12300
rect 28776 12288 28782 12300
rect 30484 12297 30512 12328
rect 28905 12291 28963 12297
rect 28905 12288 28917 12291
rect 28776 12260 28917 12288
rect 28776 12248 28782 12260
rect 28905 12257 28917 12260
rect 28951 12257 28963 12291
rect 28905 12251 28963 12257
rect 29181 12291 29239 12297
rect 29181 12257 29193 12291
rect 29227 12288 29239 12291
rect 30469 12291 30527 12297
rect 29227 12260 29960 12288
rect 29227 12257 29239 12260
rect 29181 12251 29239 12257
rect 28350 12180 28356 12232
rect 28408 12180 28414 12232
rect 29362 12220 29368 12232
rect 28552 12192 29368 12220
rect 28552 12152 28580 12192
rect 29362 12180 29368 12192
rect 29420 12180 29426 12232
rect 28184 12124 28580 12152
rect 28626 12112 28632 12164
rect 28684 12152 28690 12164
rect 29932 12161 29960 12260
rect 30469 12257 30481 12291
rect 30515 12257 30527 12291
rect 30469 12251 30527 12257
rect 30193 12223 30251 12229
rect 30193 12189 30205 12223
rect 30239 12220 30251 12223
rect 30282 12220 30288 12232
rect 30239 12192 30288 12220
rect 30239 12189 30251 12192
rect 30193 12183 30251 12189
rect 30282 12180 30288 12192
rect 30340 12180 30346 12232
rect 29917 12155 29975 12161
rect 28684 12124 28856 12152
rect 28684 12112 28690 12124
rect 26418 12084 26424 12096
rect 25700 12056 26424 12084
rect 26418 12044 26424 12056
rect 26476 12044 26482 12096
rect 26694 12044 26700 12096
rect 26752 12084 26758 12096
rect 26878 12084 26884 12096
rect 26752 12056 26884 12084
rect 26752 12044 26758 12056
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 27798 12044 27804 12096
rect 27856 12084 27862 12096
rect 28721 12087 28779 12093
rect 28721 12084 28733 12087
rect 27856 12056 28733 12084
rect 27856 12044 27862 12056
rect 28721 12053 28733 12056
rect 28767 12053 28779 12087
rect 28828 12084 28856 12124
rect 29917 12121 29929 12155
rect 29963 12121 29975 12155
rect 29917 12115 29975 12121
rect 30101 12087 30159 12093
rect 30101 12084 30113 12087
rect 28828 12056 30113 12084
rect 28721 12047 28779 12053
rect 30101 12053 30113 12056
rect 30147 12053 30159 12087
rect 30101 12047 30159 12053
rect 552 11994 31648 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 11436 11994
rect 11488 11942 11500 11994
rect 11552 11942 11564 11994
rect 11616 11942 11628 11994
rect 11680 11942 11692 11994
rect 11744 11942 19210 11994
rect 19262 11942 19274 11994
rect 19326 11942 19338 11994
rect 19390 11942 19402 11994
rect 19454 11942 19466 11994
rect 19518 11942 26984 11994
rect 27036 11942 27048 11994
rect 27100 11942 27112 11994
rect 27164 11942 27176 11994
rect 27228 11942 27240 11994
rect 27292 11942 31648 11994
rect 552 11920 31648 11942
rect 1026 11840 1032 11892
rect 1084 11880 1090 11892
rect 1305 11883 1363 11889
rect 1305 11880 1317 11883
rect 1084 11852 1317 11880
rect 1084 11840 1090 11852
rect 1305 11849 1317 11852
rect 1351 11849 1363 11883
rect 1305 11843 1363 11849
rect 2225 11883 2283 11889
rect 2225 11849 2237 11883
rect 2271 11880 2283 11883
rect 2498 11880 2504 11892
rect 2271 11852 2504 11880
rect 2271 11849 2283 11852
rect 2225 11843 2283 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 2682 11880 2688 11892
rect 2639 11852 2688 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3329 11883 3387 11889
rect 3329 11880 3341 11883
rect 3200 11852 3341 11880
rect 3200 11840 3206 11852
rect 3329 11849 3341 11852
rect 3375 11849 3387 11883
rect 3329 11843 3387 11849
rect 3694 11840 3700 11892
rect 3752 11880 3758 11892
rect 5166 11880 5172 11892
rect 3752 11852 5172 11880
rect 3752 11840 3758 11852
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6638 11880 6644 11892
rect 5951 11852 6644 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 7006 11880 7012 11892
rect 6788 11852 7012 11880
rect 6788 11840 6794 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7561 11883 7619 11889
rect 7561 11849 7573 11883
rect 7607 11880 7619 11883
rect 7650 11880 7656 11892
rect 7607 11852 7656 11880
rect 7607 11849 7619 11852
rect 7561 11843 7619 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8849 11883 8907 11889
rect 7760 11852 8805 11880
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 5810 11812 5816 11824
rect 3476 11784 5816 11812
rect 3476 11772 3482 11784
rect 2222 11744 2228 11756
rect 1596 11716 2228 11744
rect 1596 11685 1624 11716
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2958 11704 2964 11756
rect 3016 11704 3022 11756
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3602 11744 3608 11756
rect 3099 11716 3608 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 3844 11716 4016 11744
rect 3844 11704 3850 11716
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 1670 11636 1676 11688
rect 1728 11636 1734 11688
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11645 1823 11679
rect 1765 11639 1823 11645
rect 1780 11608 1808 11639
rect 1946 11636 1952 11688
rect 2004 11636 2010 11688
rect 2038 11636 2044 11688
rect 2096 11636 2102 11688
rect 2130 11636 2136 11688
rect 2188 11636 2194 11688
rect 2866 11685 2872 11688
rect 2837 11679 2872 11685
rect 2837 11676 2849 11679
rect 2240 11648 2849 11676
rect 2240 11608 2268 11648
rect 2837 11645 2849 11648
rect 2837 11639 2872 11645
rect 2866 11636 2872 11639
rect 2924 11636 2930 11688
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 2976 11648 3525 11676
rect 2976 11608 3004 11648
rect 3513 11645 3525 11648
rect 3559 11676 3571 11679
rect 3694 11676 3700 11688
rect 3559 11648 3700 11676
rect 3559 11645 3571 11648
rect 3513 11639 3571 11645
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 3878 11636 3884 11688
rect 3936 11636 3942 11688
rect 3988 11676 4016 11716
rect 4062 11704 4068 11756
rect 4120 11753 4126 11756
rect 5000 11753 5028 11784
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 5994 11772 6000 11824
rect 6052 11812 6058 11824
rect 7760 11812 7788 11852
rect 6052 11784 7788 11812
rect 6052 11772 6058 11784
rect 7834 11772 7840 11824
rect 7892 11772 7898 11824
rect 8294 11772 8300 11824
rect 8352 11812 8358 11824
rect 8662 11812 8668 11824
rect 8352 11784 8668 11812
rect 8352 11772 8358 11784
rect 8662 11772 8668 11784
rect 8720 11772 8726 11824
rect 8777 11812 8805 11852
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 9122 11880 9128 11892
rect 8895 11852 9128 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 11790 11880 11796 11892
rect 9640 11852 11796 11880
rect 9640 11840 9646 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 11977 11883 12035 11889
rect 11977 11849 11989 11883
rect 12023 11880 12035 11883
rect 14274 11880 14280 11892
rect 12023 11852 14280 11880
rect 12023 11849 12035 11852
rect 11977 11843 12035 11849
rect 9490 11812 9496 11824
rect 8777 11784 9496 11812
rect 9490 11772 9496 11784
rect 9548 11812 9554 11824
rect 10042 11812 10048 11824
rect 9548 11784 10048 11812
rect 9548 11772 9554 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10134 11772 10140 11824
rect 10192 11812 10198 11824
rect 10318 11812 10324 11824
rect 10192 11784 10324 11812
rect 10192 11772 10198 11784
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 10594 11772 10600 11824
rect 10652 11812 10658 11824
rect 11054 11812 11060 11824
rect 10652 11784 11060 11812
rect 10652 11772 10658 11784
rect 4120 11747 4142 11753
rect 4130 11713 4142 11747
rect 4120 11707 4142 11713
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 4985 11707 5043 11713
rect 5828 11716 6377 11744
rect 4120 11704 4126 11707
rect 3988 11648 4200 11676
rect 1780 11580 2268 11608
rect 2884 11580 3004 11608
rect 1946 11500 1952 11552
rect 2004 11540 2010 11552
rect 2130 11540 2136 11552
rect 2004 11512 2136 11540
rect 2004 11500 2010 11512
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2406 11500 2412 11552
rect 2464 11500 2470 11552
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 2884 11540 2912 11580
rect 3142 11568 3148 11620
rect 3200 11608 3206 11620
rect 3418 11608 3424 11620
rect 3200 11580 3424 11608
rect 3200 11568 3206 11580
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 3789 11611 3847 11617
rect 3789 11577 3801 11611
rect 3835 11608 3847 11611
rect 4062 11608 4068 11620
rect 3835 11580 4068 11608
rect 3835 11577 3847 11580
rect 3789 11571 3847 11577
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 4172 11617 4200 11648
rect 4522 11636 4528 11688
rect 4580 11676 4586 11688
rect 5828 11685 5856 11716
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11744 6515 11747
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 6503 11716 10793 11744
rect 6503 11713 6515 11716
rect 6457 11707 6515 11713
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 4709 11679 4767 11685
rect 4709 11676 4721 11679
rect 4580 11648 4721 11676
rect 4580 11636 4586 11648
rect 4709 11645 4721 11648
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 5077 11679 5135 11685
rect 5077 11645 5089 11679
rect 5123 11676 5135 11679
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5123 11648 5825 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 5813 11645 5825 11648
rect 5859 11645 5871 11679
rect 5813 11639 5871 11645
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11676 6147 11679
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 6135 11648 6653 11676
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 6641 11645 6653 11648
rect 6687 11645 6699 11679
rect 6641 11639 6699 11645
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11577 4215 11611
rect 4157 11571 4215 11577
rect 4430 11568 4436 11620
rect 4488 11608 4494 11620
rect 4617 11611 4675 11617
rect 4617 11608 4629 11611
rect 4488 11580 4629 11608
rect 4488 11568 4494 11580
rect 4617 11577 4629 11580
rect 4663 11577 4675 11611
rect 4908 11608 4936 11639
rect 5166 11608 5172 11620
rect 4908 11580 5172 11608
rect 4617 11571 4675 11577
rect 5166 11568 5172 11580
rect 5224 11568 5230 11620
rect 5258 11568 5264 11620
rect 5316 11608 5322 11620
rect 6104 11608 6132 11639
rect 5316 11580 6132 11608
rect 6656 11608 6684 11639
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 7558 11676 7564 11688
rect 7248 11648 7564 11676
rect 7248 11636 7254 11648
rect 7558 11636 7564 11648
rect 7616 11676 7622 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7616 11648 7757 11676
rect 7616 11636 7622 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 7892 11648 7941 11676
rect 7892 11636 7898 11648
rect 7929 11645 7941 11648
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8573 11679 8631 11685
rect 8067 11648 8432 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8294 11608 8300 11620
rect 6656 11580 8300 11608
rect 5316 11568 5322 11580
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 2648 11512 2912 11540
rect 2648 11500 2654 11512
rect 3694 11500 3700 11552
rect 3752 11500 3758 11552
rect 3970 11500 3976 11552
rect 4028 11500 4034 11552
rect 6270 11500 6276 11552
rect 6328 11500 6334 11552
rect 6822 11500 6828 11552
rect 6880 11500 6886 11552
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7742 11540 7748 11552
rect 7156 11512 7748 11540
rect 7156 11500 7162 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 8404 11549 8432 11648
rect 8573 11645 8585 11679
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 9122 11676 9128 11688
rect 8711 11648 9128 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 8588 11608 8616 11639
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10410 11676 10416 11688
rect 10275 11648 10416 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 10870 11676 10876 11688
rect 10643 11648 10876 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 8588 11580 8708 11608
rect 8389 11543 8447 11549
rect 8389 11509 8401 11543
rect 8435 11509 8447 11543
rect 8680 11540 8708 11580
rect 8846 11568 8852 11620
rect 8904 11568 8910 11620
rect 10520 11608 10548 11639
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 10980 11676 11008 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 11992 11812 12020 11843
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 15105 11883 15163 11889
rect 15105 11880 15117 11883
rect 14424 11852 15117 11880
rect 14424 11840 14430 11852
rect 15105 11849 15117 11852
rect 15151 11849 15163 11883
rect 15105 11843 15163 11849
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15470 11880 15476 11892
rect 15252 11852 15476 11880
rect 15252 11840 15258 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 16298 11880 16304 11892
rect 15804 11852 16304 11880
rect 15804 11840 15810 11852
rect 16298 11840 16304 11852
rect 16356 11880 16362 11892
rect 16761 11883 16819 11889
rect 16761 11880 16773 11883
rect 16356 11852 16773 11880
rect 16356 11840 16362 11852
rect 16761 11849 16773 11852
rect 16807 11849 16819 11883
rect 16761 11843 16819 11849
rect 17129 11883 17187 11889
rect 17129 11849 17141 11883
rect 17175 11880 17187 11883
rect 17402 11880 17408 11892
rect 17175 11852 17408 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17773 11883 17831 11889
rect 17773 11849 17785 11883
rect 17819 11880 17831 11883
rect 19426 11880 19432 11892
rect 17819 11852 19432 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 19898 11883 19956 11889
rect 19898 11880 19910 11883
rect 19628 11852 19910 11880
rect 11532 11784 12020 11812
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11532 11744 11560 11784
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 12584 11784 16804 11812
rect 12584 11772 12590 11784
rect 11882 11744 11888 11756
rect 11388 11716 11560 11744
rect 11624 11716 11888 11744
rect 11388 11704 11394 11716
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10980 11648 11069 11676
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11146 11636 11152 11688
rect 11204 11636 11210 11688
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 11256 11608 11284 11639
rect 11422 11636 11428 11688
rect 11480 11636 11486 11688
rect 11514 11636 11520 11688
rect 11572 11636 11578 11688
rect 11624 11685 11652 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 12676 11716 15209 11744
rect 12676 11704 12682 11716
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 11974 11636 11980 11688
rect 12032 11636 12038 11688
rect 14458 11636 14464 11688
rect 14516 11636 14522 11688
rect 14752 11685 14780 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 14737 11679 14795 11685
rect 14737 11645 14749 11679
rect 14783 11645 14795 11679
rect 14737 11639 14795 11645
rect 14826 11636 14832 11688
rect 14884 11636 14890 11688
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11670 14979 11679
rect 15102 11676 15108 11688
rect 15100 11670 15108 11676
rect 14967 11645 15108 11670
rect 14921 11642 15108 11645
rect 14921 11639 14979 11642
rect 15102 11636 15108 11642
rect 15160 11636 15166 11688
rect 15381 11679 15439 11685
rect 15381 11645 15393 11679
rect 15427 11676 15439 11679
rect 15746 11676 15752 11688
rect 15427 11648 15752 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 16776 11685 16804 11784
rect 18230 11772 18236 11824
rect 18288 11812 18294 11824
rect 19628 11812 19656 11852
rect 19898 11849 19910 11852
rect 19944 11880 19956 11883
rect 20257 11883 20315 11889
rect 19944 11852 20209 11880
rect 19944 11849 19956 11852
rect 19898 11843 19956 11849
rect 18288 11784 19656 11812
rect 19705 11815 19763 11821
rect 18288 11772 18294 11784
rect 19705 11781 19717 11815
rect 19751 11812 19763 11815
rect 19751 11784 19932 11812
rect 19751 11781 19763 11784
rect 19705 11775 19763 11781
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 18322 11744 18328 11756
rect 17727 11716 18328 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 18690 11704 18696 11756
rect 18748 11704 18754 11756
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11744 18843 11747
rect 19518 11744 19524 11756
rect 18831 11716 19524 11744
rect 18831 11713 18843 11716
rect 18785 11707 18843 11713
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 19904 11744 19932 11784
rect 20070 11772 20076 11824
rect 20128 11772 20134 11824
rect 20181 11812 20209 11852
rect 20257 11849 20269 11883
rect 20303 11880 20315 11883
rect 20530 11880 20536 11892
rect 20303 11852 20536 11880
rect 20303 11849 20315 11852
rect 20257 11843 20315 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21358 11880 21364 11892
rect 21048 11852 21364 11880
rect 21048 11840 21054 11852
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 21726 11840 21732 11892
rect 21784 11840 21790 11892
rect 22002 11840 22008 11892
rect 22060 11840 22066 11892
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 22465 11883 22523 11889
rect 22465 11880 22477 11883
rect 22336 11852 22477 11880
rect 22336 11840 22342 11852
rect 22465 11849 22477 11852
rect 22511 11849 22523 11883
rect 22465 11843 22523 11849
rect 24394 11840 24400 11892
rect 24452 11880 24458 11892
rect 25866 11880 25872 11892
rect 24452 11852 25872 11880
rect 24452 11840 24458 11852
rect 25866 11840 25872 11852
rect 25924 11840 25930 11892
rect 26234 11840 26240 11892
rect 26292 11840 26298 11892
rect 26418 11840 26424 11892
rect 26476 11880 26482 11892
rect 27341 11883 27399 11889
rect 27341 11880 27353 11883
rect 26476 11852 27353 11880
rect 26476 11840 26482 11852
rect 27341 11849 27353 11852
rect 27387 11849 27399 11883
rect 27341 11843 27399 11849
rect 28074 11840 28080 11892
rect 28132 11840 28138 11892
rect 28258 11840 28264 11892
rect 28316 11880 28322 11892
rect 28442 11880 28448 11892
rect 28316 11852 28448 11880
rect 28316 11840 28322 11852
rect 28442 11840 28448 11852
rect 28500 11840 28506 11892
rect 28537 11883 28595 11889
rect 28537 11849 28549 11883
rect 28583 11880 28595 11883
rect 28718 11880 28724 11892
rect 28583 11852 28724 11880
rect 28583 11849 28595 11852
rect 28537 11843 28595 11849
rect 28718 11840 28724 11852
rect 28776 11840 28782 11892
rect 24210 11812 24216 11824
rect 20181 11784 24216 11812
rect 24210 11772 24216 11784
rect 24268 11772 24274 11824
rect 25498 11772 25504 11824
rect 25556 11812 25562 11824
rect 26252 11812 26280 11840
rect 25556 11784 26280 11812
rect 25556 11772 25562 11784
rect 26326 11772 26332 11824
rect 26384 11812 26390 11824
rect 28350 11812 28356 11824
rect 26384 11784 26924 11812
rect 26384 11772 26390 11784
rect 20088 11744 20116 11772
rect 20625 11747 20683 11753
rect 19904 11716 20484 11744
rect 16761 11679 16819 11685
rect 16761 11645 16773 11679
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 16853 11679 16911 11685
rect 16853 11645 16865 11679
rect 16899 11645 16911 11679
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 16853 11639 16911 11645
rect 17236 11648 17785 11676
rect 11992 11608 12020 11636
rect 10520 11580 11008 11608
rect 11256 11580 12020 11608
rect 8938 11540 8944 11552
rect 8680 11512 8944 11540
rect 8389 11503 8447 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 10410 11540 10416 11552
rect 9088 11512 10416 11540
rect 9088 11500 9094 11512
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10689 11543 10747 11549
rect 10689 11509 10701 11543
rect 10735 11540 10747 11543
rect 10870 11540 10876 11552
rect 10735 11512 10876 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 10980 11540 11008 11580
rect 12342 11568 12348 11620
rect 12400 11608 12406 11620
rect 13630 11608 13636 11620
rect 12400 11580 13636 11608
rect 12400 11568 12406 11580
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 14642 11617 14648 11620
rect 14599 11611 14648 11617
rect 14599 11608 14611 11611
rect 14108 11580 14611 11608
rect 11330 11540 11336 11552
rect 10980 11512 11336 11540
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12986 11540 12992 11552
rect 11756 11512 12992 11540
rect 11756 11500 11762 11512
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 14108 11540 14136 11580
rect 14599 11577 14611 11580
rect 14645 11577 14648 11611
rect 14599 11571 14648 11577
rect 14642 11568 14648 11571
rect 14700 11568 14706 11620
rect 15562 11608 15568 11620
rect 14936 11580 15568 11608
rect 13228 11512 14136 11540
rect 13228 11500 13234 11512
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 14936 11540 14964 11580
rect 15562 11568 15568 11580
rect 15620 11568 15626 11620
rect 16022 11568 16028 11620
rect 16080 11608 16086 11620
rect 16868 11608 16896 11639
rect 16080 11580 16896 11608
rect 16080 11568 16086 11580
rect 14240 11512 14964 11540
rect 14240 11500 14246 11512
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 17236 11549 17264 11648
rect 17773 11645 17785 11648
rect 17819 11645 17831 11679
rect 18340 11676 18368 11704
rect 18598 11676 18604 11688
rect 18340 11648 18604 11676
rect 17773 11639 17831 11645
rect 18598 11636 18604 11648
rect 18656 11676 18662 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18656 11648 18981 11676
rect 18656 11636 18662 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 20456 11685 20484 11716
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 21545 11747 21603 11753
rect 21545 11744 21557 11747
rect 20671 11716 21557 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 21545 11713 21557 11716
rect 21591 11713 21603 11747
rect 21545 11707 21603 11713
rect 21634 11704 21640 11756
rect 21692 11744 21698 11756
rect 23290 11744 23296 11756
rect 21692 11716 23296 11744
rect 21692 11704 21698 11716
rect 23290 11704 23296 11716
rect 23348 11704 23354 11756
rect 24118 11704 24124 11756
rect 24176 11744 24182 11756
rect 24176 11716 24624 11744
rect 24176 11704 24182 11716
rect 20165 11679 20223 11685
rect 19484 11648 20041 11676
rect 19484 11636 19490 11648
rect 18874 11568 18880 11620
rect 18932 11608 18938 11620
rect 18932 11580 19288 11608
rect 18932 11568 18938 11580
rect 17221 11543 17279 11549
rect 17221 11540 17233 11543
rect 15252 11512 17233 11540
rect 15252 11500 15258 11512
rect 17221 11509 17233 11512
rect 17267 11509 17279 11543
rect 17221 11503 17279 11509
rect 17402 11500 17408 11552
rect 17460 11500 17466 11552
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 19153 11543 19211 11549
rect 19153 11540 19165 11543
rect 18196 11512 19165 11540
rect 18196 11500 18202 11512
rect 19153 11509 19165 11512
rect 19199 11509 19211 11543
rect 19260 11540 19288 11580
rect 19518 11540 19524 11552
rect 19260 11512 19524 11540
rect 19153 11503 19211 11509
rect 19518 11500 19524 11512
rect 19576 11540 19582 11552
rect 19863 11543 19921 11549
rect 19863 11540 19875 11543
rect 19576 11512 19875 11540
rect 19576 11500 19582 11512
rect 19863 11509 19875 11512
rect 19909 11509 19921 11543
rect 20013 11540 20041 11648
rect 20165 11645 20177 11679
rect 20211 11645 20223 11679
rect 20165 11639 20223 11645
rect 20441 11679 20499 11685
rect 20441 11645 20453 11679
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 20070 11568 20076 11620
rect 20128 11568 20134 11620
rect 20180 11608 20208 11639
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 21453 11679 21511 11685
rect 21453 11676 21465 11679
rect 21416 11648 21465 11676
rect 21416 11636 21422 11648
rect 21453 11645 21465 11648
rect 21499 11645 21511 11679
rect 21453 11639 21511 11645
rect 21729 11679 21787 11685
rect 21729 11645 21741 11679
rect 21775 11676 21787 11679
rect 21818 11676 21824 11688
rect 21775 11648 21824 11676
rect 21775 11645 21787 11648
rect 21729 11639 21787 11645
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 22094 11636 22100 11688
rect 22152 11676 22158 11688
rect 22281 11679 22339 11685
rect 22281 11676 22293 11679
rect 22152 11648 22293 11676
rect 22152 11636 22158 11648
rect 22281 11645 22293 11648
rect 22327 11645 22339 11679
rect 22281 11639 22339 11645
rect 22370 11636 22376 11688
rect 22428 11636 22434 11688
rect 22554 11636 22560 11688
rect 22612 11636 22618 11688
rect 22738 11636 22744 11688
rect 22796 11676 22802 11688
rect 23014 11676 23020 11688
rect 22796 11648 23020 11676
rect 22796 11636 22802 11648
rect 23014 11636 23020 11648
rect 23072 11636 23078 11688
rect 23934 11636 23940 11688
rect 23992 11676 23998 11688
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 23992 11648 24225 11676
rect 23992 11636 23998 11648
rect 24213 11645 24225 11648
rect 24259 11645 24271 11679
rect 24213 11639 24271 11645
rect 24486 11636 24492 11688
rect 24544 11636 24550 11688
rect 24596 11685 24624 11716
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25004 11716 26556 11744
rect 25004 11704 25010 11716
rect 24581 11679 24639 11685
rect 24581 11645 24593 11679
rect 24627 11645 24639 11679
rect 24581 11639 24639 11645
rect 25314 11636 25320 11688
rect 25372 11636 25378 11688
rect 25498 11636 25504 11688
rect 25556 11676 25562 11688
rect 25593 11679 25651 11685
rect 25593 11676 25605 11679
rect 25556 11648 25605 11676
rect 25556 11636 25562 11648
rect 25593 11645 25605 11648
rect 25639 11645 25651 11679
rect 25593 11639 25651 11645
rect 25685 11679 25743 11685
rect 25685 11645 25697 11679
rect 25731 11676 25743 11679
rect 25866 11676 25872 11688
rect 25731 11648 25872 11676
rect 25731 11645 25743 11648
rect 25685 11639 25743 11645
rect 25866 11636 25872 11648
rect 25924 11636 25930 11688
rect 26142 11636 26148 11688
rect 26200 11676 26206 11688
rect 26396 11679 26454 11685
rect 26396 11676 26408 11679
rect 26200 11648 26408 11676
rect 26200 11636 26206 11648
rect 26396 11645 26408 11648
rect 26442 11645 26454 11679
rect 26528 11676 26556 11716
rect 26602 11704 26608 11756
rect 26660 11704 26666 11756
rect 26896 11753 26924 11784
rect 26988 11784 28356 11812
rect 26881 11747 26939 11753
rect 26881 11713 26893 11747
rect 26927 11713 26939 11747
rect 26881 11707 26939 11713
rect 26988 11676 27016 11784
rect 28350 11772 28356 11784
rect 28408 11812 28414 11824
rect 30466 11812 30472 11824
rect 28408 11784 30472 11812
rect 28408 11772 28414 11784
rect 27246 11704 27252 11756
rect 27304 11744 27310 11756
rect 27706 11744 27712 11756
rect 27304 11716 27712 11744
rect 27304 11704 27310 11716
rect 27706 11704 27712 11716
rect 27764 11704 27770 11756
rect 28534 11704 28540 11756
rect 28592 11744 28598 11756
rect 28592 11716 29592 11744
rect 28592 11704 28598 11716
rect 29564 11688 29592 11716
rect 26528 11648 27016 11676
rect 26396 11639 26454 11645
rect 27062 11636 27068 11688
rect 27120 11636 27126 11688
rect 27157 11679 27215 11685
rect 27157 11645 27169 11679
rect 27203 11676 27215 11679
rect 27890 11676 27896 11688
rect 27203 11648 27896 11676
rect 27203 11645 27215 11648
rect 27157 11639 27215 11645
rect 27890 11636 27896 11648
rect 27948 11636 27954 11688
rect 28350 11636 28356 11688
rect 28408 11636 28414 11688
rect 28629 11679 28687 11685
rect 28629 11645 28641 11679
rect 28675 11676 28687 11679
rect 28994 11676 29000 11688
rect 28675 11648 29000 11676
rect 28675 11645 28687 11648
rect 28629 11639 28687 11645
rect 28994 11636 29000 11648
rect 29052 11636 29058 11688
rect 29454 11636 29460 11688
rect 29512 11636 29518 11688
rect 29546 11636 29552 11688
rect 29604 11636 29610 11688
rect 29748 11685 29776 11784
rect 30466 11772 30472 11784
rect 30524 11812 30530 11824
rect 30561 11815 30619 11821
rect 30561 11812 30573 11815
rect 30524 11784 30573 11812
rect 30524 11772 30530 11784
rect 30561 11781 30573 11784
rect 30607 11781 30619 11815
rect 30561 11775 30619 11781
rect 29822 11704 29828 11756
rect 29880 11744 29886 11756
rect 30745 11747 30803 11753
rect 29880 11716 30236 11744
rect 29880 11704 29886 11716
rect 29733 11679 29791 11685
rect 29733 11645 29745 11679
rect 29779 11645 29791 11679
rect 29733 11639 29791 11645
rect 29917 11679 29975 11685
rect 29917 11645 29929 11679
rect 29963 11676 29975 11679
rect 30006 11676 30012 11688
rect 29963 11648 30012 11676
rect 29963 11645 29975 11648
rect 29917 11639 29975 11645
rect 20622 11608 20628 11620
rect 20180 11580 20628 11608
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 24302 11608 24308 11620
rect 21192 11580 24308 11608
rect 21192 11540 21220 11580
rect 24302 11568 24308 11580
rect 24360 11568 24366 11620
rect 24504 11608 24532 11636
rect 25409 11611 25467 11617
rect 25409 11608 25421 11611
rect 24504 11580 25421 11608
rect 25409 11577 25421 11580
rect 25455 11608 25467 11611
rect 25961 11611 26019 11617
rect 25961 11608 25973 11611
rect 25455 11580 25973 11608
rect 25455 11577 25467 11580
rect 25409 11571 25467 11577
rect 25961 11577 25973 11580
rect 26007 11577 26019 11611
rect 25961 11571 26019 11577
rect 27341 11611 27399 11617
rect 27341 11577 27353 11611
rect 27387 11608 27399 11611
rect 27522 11608 27528 11620
rect 27387 11580 27528 11608
rect 27387 11577 27399 11580
rect 27341 11571 27399 11577
rect 27522 11568 27528 11580
rect 27580 11568 27586 11620
rect 28258 11568 28264 11620
rect 28316 11608 28322 11620
rect 28534 11608 28540 11620
rect 28316 11580 28540 11608
rect 28316 11568 28322 11580
rect 28534 11568 28540 11580
rect 28592 11568 28598 11620
rect 28902 11568 28908 11620
rect 28960 11608 28966 11620
rect 29932 11608 29960 11639
rect 30006 11636 30012 11648
rect 30064 11636 30070 11688
rect 30208 11685 30236 11716
rect 30745 11713 30757 11747
rect 30791 11744 30803 11747
rect 31018 11744 31024 11756
rect 30791 11716 31024 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 31018 11704 31024 11716
rect 31076 11704 31082 11756
rect 30193 11679 30251 11685
rect 30193 11645 30205 11679
rect 30239 11645 30251 11679
rect 30193 11639 30251 11645
rect 30282 11636 30288 11688
rect 30340 11676 30346 11688
rect 30929 11679 30987 11685
rect 30929 11676 30941 11679
rect 30340 11648 30941 11676
rect 30340 11636 30346 11648
rect 30929 11645 30941 11648
rect 30975 11645 30987 11679
rect 30929 11639 30987 11645
rect 28960 11580 29960 11608
rect 28960 11568 28966 11580
rect 20013 11512 21220 11540
rect 21269 11543 21327 11549
rect 19863 11503 19921 11509
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21450 11540 21456 11552
rect 21315 11512 21456 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 22646 11500 22652 11552
rect 22704 11540 22710 11552
rect 24029 11543 24087 11549
rect 24029 11540 24041 11543
rect 22704 11512 24041 11540
rect 22704 11500 22710 11512
rect 24029 11509 24041 11512
rect 24075 11540 24087 11543
rect 24118 11540 24124 11552
rect 24075 11512 24124 11540
rect 24075 11509 24087 11512
rect 24029 11503 24087 11509
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 24486 11540 24492 11552
rect 24443 11512 24492 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 25498 11549 25504 11552
rect 25494 11503 25504 11549
rect 25498 11500 25504 11503
rect 25556 11500 25562 11552
rect 26513 11543 26571 11549
rect 26513 11509 26525 11543
rect 26559 11540 26571 11543
rect 27430 11540 27436 11552
rect 26559 11512 27436 11540
rect 26559 11509 26571 11512
rect 26513 11503 26571 11509
rect 27430 11500 27436 11512
rect 27488 11500 27494 11552
rect 27614 11500 27620 11552
rect 27672 11540 27678 11552
rect 29086 11540 29092 11552
rect 27672 11512 29092 11540
rect 27672 11500 27678 11512
rect 29086 11500 29092 11512
rect 29144 11500 29150 11552
rect 29178 11500 29184 11552
rect 29236 11540 29242 11552
rect 29273 11543 29331 11549
rect 29273 11540 29285 11543
rect 29236 11512 29285 11540
rect 29236 11500 29242 11512
rect 29273 11509 29285 11512
rect 29319 11509 29331 11543
rect 29273 11503 29331 11509
rect 29638 11500 29644 11552
rect 29696 11500 29702 11552
rect 552 11450 31648 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 12096 11450
rect 12148 11398 12160 11450
rect 12212 11398 12224 11450
rect 12276 11398 12288 11450
rect 12340 11398 12352 11450
rect 12404 11398 19870 11450
rect 19922 11398 19934 11450
rect 19986 11398 19998 11450
rect 20050 11398 20062 11450
rect 20114 11398 20126 11450
rect 20178 11398 27644 11450
rect 27696 11398 27708 11450
rect 27760 11398 27772 11450
rect 27824 11398 27836 11450
rect 27888 11398 27900 11450
rect 27952 11398 31648 11450
rect 552 11376 31648 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 2590 11336 2596 11348
rect 1452 11308 2596 11336
rect 1452 11296 1458 11308
rect 1302 11160 1308 11212
rect 1360 11200 1366 11212
rect 1504 11209 1532 11308
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 3970 11336 3976 11348
rect 3651 11308 3976 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5166 11336 5172 11348
rect 4672 11308 5172 11336
rect 4672 11296 4678 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 6086 11296 6092 11348
rect 6144 11336 6150 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6144 11308 6745 11336
rect 6144 11296 6150 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7708 11308 8033 11336
rect 7708 11296 7714 11308
rect 8021 11305 8033 11308
rect 8067 11305 8079 11339
rect 9582 11336 9588 11348
rect 8021 11299 8079 11305
rect 8128 11308 9588 11336
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 1820 11240 2268 11268
rect 1820 11228 1826 11240
rect 1397 11203 1455 11209
rect 1397 11200 1409 11203
rect 1360 11172 1409 11200
rect 1360 11160 1366 11172
rect 1397 11169 1409 11172
rect 1443 11169 1455 11203
rect 1397 11163 1455 11169
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11169 1547 11203
rect 1489 11163 1547 11169
rect 1412 11132 1440 11163
rect 2130 11160 2136 11212
rect 2188 11160 2194 11212
rect 2240 11200 2268 11240
rect 2314 11228 2320 11280
rect 2372 11268 2378 11280
rect 2372 11240 2544 11268
rect 2372 11228 2378 11240
rect 2516 11209 2544 11240
rect 2958 11228 2964 11280
rect 3016 11228 3022 11280
rect 3234 11228 3240 11280
rect 3292 11268 3298 11280
rect 4065 11271 4123 11277
rect 4065 11268 4077 11271
rect 3292 11240 4077 11268
rect 3292 11228 3298 11240
rect 4065 11237 4077 11240
rect 4111 11237 4123 11271
rect 4522 11268 4528 11280
rect 4065 11231 4123 11237
rect 4172 11240 4528 11268
rect 2501 11203 2559 11209
rect 2240 11172 2452 11200
rect 2424 11144 2452 11172
rect 2501 11169 2513 11203
rect 2547 11169 2559 11203
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2501 11163 2559 11169
rect 2793 11172 2881 11200
rect 2225 11135 2283 11141
rect 1412 11104 1532 11132
rect 1504 10996 1532 11104
rect 2225 11101 2237 11135
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2240 11064 2268 11095
rect 2406 11092 2412 11144
rect 2464 11132 2470 11144
rect 2793 11132 2821 11172
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 2976 11200 3004 11228
rect 3053 11203 3111 11209
rect 3053 11200 3065 11203
rect 2976 11172 3065 11200
rect 2869 11163 2927 11169
rect 3053 11169 3065 11172
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 3142 11160 3148 11212
rect 3200 11160 3206 11212
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11200 3479 11203
rect 3467 11172 3556 11200
rect 3467 11169 3479 11172
rect 3421 11163 3479 11169
rect 2464 11104 2821 11132
rect 2464 11092 2470 11104
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3344 11132 3372 11163
rect 3528 11144 3556 11172
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 4172 11200 4200 11240
rect 4522 11228 4528 11240
rect 4580 11228 4586 11280
rect 5092 11240 7972 11268
rect 3752 11172 4200 11200
rect 3752 11160 3758 11172
rect 4246 11160 4252 11212
rect 4304 11200 4310 11212
rect 4617 11203 4675 11209
rect 4617 11200 4629 11203
rect 4304 11172 4629 11200
rect 4304 11160 4310 11172
rect 4617 11169 4629 11172
rect 4663 11169 4675 11203
rect 4617 11163 4675 11169
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4764 11172 4997 11200
rect 4764 11160 4770 11172
rect 4985 11169 4997 11172
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 3016 11104 3372 11132
rect 3016 11092 3022 11104
rect 3510 11092 3516 11144
rect 3568 11132 3574 11144
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 3568 11104 4445 11132
rect 3568 11092 3574 11104
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 2866 11064 2872 11076
rect 2240 11036 2872 11064
rect 2866 11024 2872 11036
rect 2924 11064 2930 11076
rect 5092 11064 5120 11240
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 6730 11200 6736 11212
rect 5408 11172 6736 11200
rect 5408 11160 5414 11172
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 2924 11036 5120 11064
rect 2924 11024 2930 11036
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 6932 11064 6960 11163
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 7944 11209 7972 11240
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 7929 11163 7987 11169
rect 7098 11092 7104 11144
rect 7156 11092 7162 11144
rect 7944 11132 7972 11163
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 8128 11209 8156 11308
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11609 11339 11667 11345
rect 10928 11308 11560 11336
rect 10928 11296 10934 11308
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 8352 11240 11376 11268
rect 8352 11228 8358 11240
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 8076 11172 8125 11200
rect 8076 11160 8082 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8938 11160 8944 11212
rect 8996 11160 9002 11212
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11198 9183 11203
rect 9214 11198 9220 11212
rect 9171 11170 9220 11198
rect 9171 11169 9183 11170
rect 9125 11163 9183 11169
rect 9214 11160 9220 11170
rect 9272 11160 9278 11212
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9030 11132 9036 11144
rect 7944 11104 9036 11132
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9416 11132 9444 11163
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9548 11172 9597 11200
rect 9548 11160 9554 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 11348 11209 11376 11240
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 9824 11172 10977 11200
rect 9824 11160 9830 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 10686 11132 10692 11144
rect 9416 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 11164 11132 11192 11163
rect 10928 11104 11192 11132
rect 11348 11132 11376 11163
rect 11422 11160 11428 11212
rect 11480 11160 11486 11212
rect 11532 11209 11560 11308
rect 11609 11305 11621 11339
rect 11655 11336 11667 11339
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 11655 11308 12265 11336
rect 11655 11305 11667 11308
rect 11609 11299 11667 11305
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 13722 11336 13728 11348
rect 12253 11299 12311 11305
rect 12360 11308 13728 11336
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 12360 11268 12388 11308
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 14277 11339 14335 11345
rect 14277 11305 14289 11339
rect 14323 11336 14335 11339
rect 14458 11336 14464 11348
rect 14323 11308 14464 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 14642 11296 14648 11348
rect 14700 11336 14706 11348
rect 15197 11339 15255 11345
rect 15197 11336 15209 11339
rect 14700 11308 15209 11336
rect 14700 11296 14706 11308
rect 15197 11305 15209 11308
rect 15243 11305 15255 11339
rect 15197 11299 15255 11305
rect 11756 11240 12388 11268
rect 12452 11240 13216 11268
rect 11756 11228 11762 11240
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 11974 11200 11980 11212
rect 11839 11172 11980 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12342 11132 12348 11144
rect 11348 11104 12348 11132
rect 10928 11092 10934 11104
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12452 11141 12480 11240
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11200 12955 11203
rect 12986 11200 12992 11212
rect 12943 11172 12992 11200
rect 12943 11169 12955 11172
rect 12897 11163 12955 11169
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 13188 11209 13216 11240
rect 13262 11228 13268 11280
rect 13320 11268 13326 11280
rect 13320 11240 14780 11268
rect 13320 11228 13326 11240
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11169 13139 11203
rect 13081 11163 13139 11169
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12713 11135 12771 11141
rect 12575 11104 12664 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 6788 11036 11805 11064
rect 6788 11024 6794 11036
rect 11793 11033 11805 11036
rect 11839 11033 11851 11067
rect 12452 11064 12480 11095
rect 12636 11076 12664 11104
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 13096 11132 13124 11163
rect 13354 11160 13360 11212
rect 13412 11160 13418 11212
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13780 11172 14105 11200
rect 13780 11160 13786 11172
rect 14093 11169 14105 11172
rect 14139 11200 14151 11203
rect 14182 11200 14188 11212
rect 14139 11172 14188 11200
rect 14139 11169 14151 11172
rect 14093 11163 14151 11169
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11200 14335 11203
rect 14366 11200 14372 11212
rect 14323 11172 14372 11200
rect 14323 11169 14335 11172
rect 14277 11163 14335 11169
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 14752 11209 14780 11240
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 15013 11271 15071 11277
rect 15013 11268 15025 11271
rect 14976 11240 15025 11268
rect 14976 11228 14982 11240
rect 15013 11237 15025 11240
rect 15059 11237 15071 11271
rect 15212 11268 15240 11299
rect 16850 11296 16856 11348
rect 16908 11296 16914 11348
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 19702 11336 19708 11348
rect 17552 11308 19708 11336
rect 17552 11296 17558 11308
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 19886 11296 19892 11348
rect 19944 11336 19950 11348
rect 20438 11336 20444 11348
rect 19944 11308 20444 11336
rect 19944 11296 19950 11308
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 20732 11308 21772 11336
rect 20349 11271 20407 11277
rect 20349 11268 20361 11271
rect 15212 11240 20361 11268
rect 15013 11231 15071 11237
rect 20349 11237 20361 11240
rect 20395 11268 20407 11271
rect 20732 11268 20760 11308
rect 20395 11240 20760 11268
rect 20395 11237 20407 11240
rect 20349 11231 20407 11237
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 21634 11268 21640 11280
rect 21232 11240 21640 11268
rect 21232 11228 21238 11240
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 21744 11268 21772 11308
rect 22554 11296 22560 11348
rect 22612 11336 22618 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22612 11308 22937 11336
rect 22612 11296 22618 11308
rect 22925 11305 22937 11308
rect 22971 11336 22983 11339
rect 23014 11336 23020 11348
rect 22971 11308 23020 11336
rect 22971 11305 22983 11308
rect 22925 11299 22983 11305
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 23474 11296 23480 11348
rect 23532 11296 23538 11348
rect 24026 11336 24032 11348
rect 23584 11308 24032 11336
rect 21744 11240 22784 11268
rect 14737 11203 14795 11209
rect 14737 11169 14749 11203
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15378 11200 15384 11212
rect 15335 11172 15384 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 16347 11203 16405 11209
rect 16347 11200 16359 11203
rect 15620 11172 16359 11200
rect 15620 11160 15626 11172
rect 16347 11169 16359 11172
rect 16393 11169 16405 11203
rect 16347 11163 16405 11169
rect 16482 11160 16488 11212
rect 16540 11160 16546 11212
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 17402 11200 17408 11212
rect 16715 11172 17408 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 19150 11160 19156 11212
rect 19208 11200 19214 11212
rect 19610 11200 19616 11212
rect 19208 11172 19616 11200
rect 19208 11160 19214 11172
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 19978 11200 19984 11212
rect 19760 11172 19984 11200
rect 19760 11160 19766 11172
rect 19978 11160 19984 11172
rect 20036 11160 20042 11212
rect 20257 11203 20315 11209
rect 20257 11200 20269 11203
rect 20088 11172 20269 11200
rect 20088 11144 20116 11172
rect 20257 11169 20269 11172
rect 20303 11169 20315 11203
rect 20257 11163 20315 11169
rect 20438 11160 20444 11212
rect 20496 11200 20502 11212
rect 22186 11200 22192 11212
rect 20496 11172 22192 11200
rect 20496 11160 20502 11172
rect 22186 11160 22192 11172
rect 22244 11160 22250 11212
rect 13630 11132 13636 11144
rect 13096 11104 13636 11132
rect 12713 11095 12771 11101
rect 11793 11027 11851 11033
rect 12360 11036 12480 11064
rect 3694 10996 3700 11008
rect 1504 10968 3700 10996
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 3973 10999 4031 11005
rect 3973 10996 3985 10999
rect 3844 10968 3985 10996
rect 3844 10956 3850 10968
rect 3973 10965 3985 10968
rect 4019 10996 4031 10999
rect 4430 10996 4436 11008
rect 4019 10968 4436 10996
rect 4019 10965 4031 10968
rect 3973 10959 4031 10965
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 5810 10996 5816 11008
rect 4580 10968 5816 10996
rect 4580 10956 4586 10968
rect 5810 10956 5816 10968
rect 5868 10956 5874 11008
rect 6086 10956 6092 11008
rect 6144 10996 6150 11008
rect 6546 10996 6552 11008
rect 6144 10968 6552 10996
rect 6144 10956 6150 10968
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 6917 10999 6975 11005
rect 6917 10996 6929 10999
rect 6880 10968 6929 10996
rect 6880 10956 6886 10968
rect 6917 10965 6929 10968
rect 6963 10965 6975 10999
rect 6917 10959 6975 10965
rect 7742 10956 7748 11008
rect 7800 10996 7806 11008
rect 8754 10996 8760 11008
rect 7800 10968 8760 10996
rect 7800 10956 7806 10968
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 9125 10999 9183 11005
rect 9125 10996 9137 10999
rect 9088 10968 9137 10996
rect 9088 10956 9094 10968
rect 9125 10965 9137 10968
rect 9171 10965 9183 10999
rect 9125 10959 9183 10965
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 10226 10996 10232 11008
rect 9640 10968 10232 10996
rect 9640 10956 9646 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 12360 10996 12388 11036
rect 12618 11024 12624 11076
rect 12676 11024 12682 11076
rect 12728 11064 12756 11095
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 13786 11104 14565 11132
rect 12989 11067 13047 11073
rect 12989 11064 13001 11067
rect 12728 11036 13001 11064
rect 12989 11033 13001 11036
rect 13035 11033 13047 11067
rect 13786 11064 13814 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11132 14887 11135
rect 15085 11135 15143 11141
rect 15085 11132 15097 11135
rect 14875 11104 15097 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 15085 11101 15097 11104
rect 15131 11101 15143 11135
rect 16022 11132 16028 11144
rect 15085 11095 15143 11101
rect 15305 11104 16028 11132
rect 12989 11027 13047 11033
rect 13280 11036 13814 11064
rect 10468 10968 12388 10996
rect 10468 10956 10474 10968
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13280 11005 13308 11036
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14660 11064 14688 11095
rect 15305 11064 15333 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 16172 11104 16221 11132
rect 16172 11092 16178 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 16816 11104 20024 11132
rect 16816 11092 16822 11104
rect 14240 11036 14596 11064
rect 14660 11036 15333 11064
rect 14240 11024 14246 11036
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 12952 10968 13277 10996
rect 12952 10956 12958 10968
rect 13265 10965 13277 10968
rect 13311 10965 13323 10999
rect 13265 10959 13323 10965
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 13964 10968 14381 10996
rect 13964 10956 13970 10968
rect 14369 10965 14381 10968
rect 14415 10965 14427 10999
rect 14568 10996 14596 11036
rect 15378 11024 15384 11076
rect 15436 11064 15442 11076
rect 15562 11064 15568 11076
rect 15436 11036 15568 11064
rect 15436 11024 15442 11036
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 19886 11064 19892 11076
rect 15712 11036 19892 11064
rect 15712 11024 15718 11036
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 19996 11064 20024 11104
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 20180 11104 20714 11132
rect 20180 11064 20208 11104
rect 19996 11036 20208 11064
rect 20686 11064 20714 11104
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 22756 11132 22784 11240
rect 22830 11160 22836 11212
rect 22888 11160 22894 11212
rect 23017 11203 23075 11209
rect 23017 11169 23029 11203
rect 23063 11200 23075 11203
rect 23584 11200 23612 11308
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24302 11296 24308 11348
rect 24360 11336 24366 11348
rect 24578 11336 24584 11348
rect 24360 11308 24584 11336
rect 24360 11296 24366 11308
rect 24578 11296 24584 11308
rect 24636 11336 24642 11348
rect 24636 11308 25222 11336
rect 24636 11296 24642 11308
rect 23842 11268 23848 11280
rect 23768 11240 23848 11268
rect 23768 11209 23796 11240
rect 23842 11228 23848 11240
rect 23900 11228 23906 11280
rect 24118 11268 24124 11280
rect 23952 11240 24124 11268
rect 23952 11209 23980 11240
rect 24118 11228 24124 11240
rect 24176 11228 24182 11280
rect 24762 11228 24768 11280
rect 24820 11228 24826 11280
rect 25194 11277 25222 11308
rect 25590 11296 25596 11348
rect 25648 11336 25654 11348
rect 25685 11339 25743 11345
rect 25685 11336 25697 11339
rect 25648 11308 25697 11336
rect 25648 11296 25654 11308
rect 25685 11305 25697 11308
rect 25731 11305 25743 11339
rect 25685 11299 25743 11305
rect 27430 11296 27436 11348
rect 27488 11296 27494 11348
rect 27982 11336 27988 11348
rect 27632 11308 27988 11336
rect 25179 11271 25237 11277
rect 25179 11237 25191 11271
rect 25225 11237 25237 11271
rect 25179 11231 25237 11237
rect 25406 11228 25412 11280
rect 25464 11228 25470 11280
rect 27448 11268 27476 11296
rect 27632 11277 27660 11308
rect 27982 11296 27988 11308
rect 28040 11296 28046 11348
rect 28350 11296 28356 11348
rect 28408 11336 28414 11348
rect 29457 11339 29515 11345
rect 29457 11336 29469 11339
rect 28408 11308 29469 11336
rect 28408 11296 28414 11308
rect 29457 11305 29469 11308
rect 29503 11305 29515 11339
rect 29457 11299 29515 11305
rect 29546 11296 29552 11348
rect 29604 11336 29610 11348
rect 30285 11339 30343 11345
rect 30285 11336 30297 11339
rect 29604 11308 30297 11336
rect 29604 11296 29610 11308
rect 30285 11305 30297 11308
rect 30331 11305 30343 11339
rect 30285 11299 30343 11305
rect 27356 11240 27476 11268
rect 27617 11271 27675 11277
rect 23063 11172 23612 11200
rect 23661 11203 23719 11209
rect 23063 11169 23075 11172
rect 23017 11163 23075 11169
rect 23661 11169 23673 11203
rect 23707 11169 23719 11203
rect 23661 11163 23719 11169
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11169 23811 11203
rect 23753 11163 23811 11169
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11169 23995 11203
rect 23937 11163 23995 11169
rect 23676 11132 23704 11163
rect 24946 11160 24952 11212
rect 25004 11200 25010 11212
rect 25041 11203 25099 11209
rect 25041 11200 25053 11203
rect 25004 11172 25053 11200
rect 25004 11160 25010 11172
rect 25041 11169 25053 11172
rect 25087 11169 25099 11203
rect 25041 11163 25099 11169
rect 25317 11203 25375 11209
rect 25317 11169 25329 11203
rect 25363 11200 25375 11203
rect 25363 11172 25452 11200
rect 25363 11169 25375 11172
rect 25317 11163 25375 11169
rect 21600 11104 22692 11132
rect 22756 11104 23704 11132
rect 21600 11092 21606 11104
rect 21910 11064 21916 11076
rect 20686 11036 21916 11064
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 22664 11064 22692 11104
rect 23842 11092 23848 11144
rect 23900 11092 23906 11144
rect 24394 11092 24400 11144
rect 24452 11132 24458 11144
rect 25424 11132 25452 11172
rect 25498 11160 25504 11212
rect 25556 11160 25562 11212
rect 26234 11160 26240 11212
rect 26292 11200 26298 11212
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 26292 11172 27169 11200
rect 26292 11160 26298 11172
rect 27157 11169 27169 11172
rect 27203 11169 27215 11203
rect 27157 11163 27215 11169
rect 27246 11160 27252 11212
rect 27304 11160 27310 11212
rect 27356 11209 27384 11240
rect 27617 11237 27629 11271
rect 27663 11237 27675 11271
rect 27617 11231 27675 11237
rect 27798 11228 27804 11280
rect 27856 11268 27862 11280
rect 29638 11268 29644 11280
rect 27856 11240 28120 11268
rect 27856 11228 27862 11240
rect 27341 11203 27399 11209
rect 27341 11169 27353 11203
rect 27387 11169 27399 11203
rect 27341 11163 27399 11169
rect 27433 11203 27491 11209
rect 27433 11169 27445 11203
rect 27479 11200 27491 11203
rect 27522 11200 27528 11212
rect 27479 11172 27528 11200
rect 27479 11169 27491 11172
rect 27433 11163 27491 11169
rect 27522 11160 27528 11172
rect 27580 11160 27586 11212
rect 27706 11160 27712 11212
rect 27764 11200 27770 11212
rect 28092 11209 28120 11240
rect 29104 11240 29644 11268
rect 27893 11203 27951 11209
rect 27893 11200 27905 11203
rect 27764 11172 27905 11200
rect 27764 11160 27770 11172
rect 27893 11169 27905 11172
rect 27939 11169 27951 11203
rect 27893 11163 27951 11169
rect 27985 11203 28043 11209
rect 27985 11169 27997 11203
rect 28031 11169 28043 11203
rect 27985 11163 28043 11169
rect 28077 11203 28135 11209
rect 28077 11169 28089 11203
rect 28123 11169 28135 11203
rect 28077 11163 28135 11169
rect 27993 11132 28021 11163
rect 28258 11160 28264 11212
rect 28316 11160 28322 11212
rect 28445 11203 28503 11209
rect 28445 11169 28457 11203
rect 28491 11200 28503 11203
rect 28718 11200 28724 11212
rect 28491 11172 28724 11200
rect 28491 11169 28503 11172
rect 28445 11163 28503 11169
rect 28718 11160 28724 11172
rect 28776 11160 28782 11212
rect 29104 11209 29132 11240
rect 29638 11228 29644 11240
rect 29696 11268 29702 11280
rect 30837 11271 30895 11277
rect 29696 11240 29868 11268
rect 29696 11228 29702 11240
rect 29089 11203 29147 11209
rect 29089 11200 29101 11203
rect 29012 11172 29101 11200
rect 28905 11135 28963 11141
rect 28905 11132 28917 11135
rect 24452 11104 27844 11132
rect 27993 11104 28917 11132
rect 24452 11092 24458 11104
rect 24026 11064 24032 11076
rect 22664 11036 24032 11064
rect 24026 11024 24032 11036
rect 24084 11024 24090 11076
rect 26050 11064 26056 11076
rect 24136 11036 26056 11064
rect 18874 10996 18880 11008
rect 14568 10968 18880 10996
rect 14369 10959 14427 10965
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 20714 10996 20720 11008
rect 20036 10968 20720 10996
rect 20036 10956 20042 10968
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 20898 10956 20904 11008
rect 20956 10996 20962 11008
rect 22186 10996 22192 11008
rect 20956 10968 22192 10996
rect 20956 10956 20962 10968
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 22830 10956 22836 11008
rect 22888 10996 22894 11008
rect 24136 10996 24164 11036
rect 26050 11024 26056 11036
rect 26108 11064 26114 11076
rect 27706 11064 27712 11076
rect 26108 11036 27712 11064
rect 26108 11024 26114 11036
rect 27706 11024 27712 11036
rect 27764 11024 27770 11076
rect 27816 11064 27844 11104
rect 28905 11101 28917 11104
rect 28951 11101 28963 11135
rect 28905 11095 28963 11101
rect 29012 11064 29040 11172
rect 29089 11169 29101 11172
rect 29135 11169 29147 11203
rect 29089 11163 29147 11169
rect 29730 11160 29736 11212
rect 29788 11160 29794 11212
rect 29840 11209 29868 11240
rect 30837 11237 30849 11271
rect 30883 11268 30895 11271
rect 30926 11268 30932 11280
rect 30883 11240 30932 11268
rect 30883 11237 30895 11240
rect 30837 11231 30895 11237
rect 30926 11228 30932 11240
rect 30984 11228 30990 11280
rect 29825 11203 29883 11209
rect 29825 11169 29837 11203
rect 29871 11169 29883 11203
rect 29825 11163 29883 11169
rect 29914 11160 29920 11212
rect 29972 11160 29978 11212
rect 30101 11203 30159 11209
rect 30101 11169 30113 11203
rect 30147 11169 30159 11203
rect 30101 11163 30159 11169
rect 29365 11135 29423 11141
rect 29365 11132 29377 11135
rect 27816 11036 29040 11064
rect 29196 11104 29377 11132
rect 22888 10968 24164 10996
rect 22888 10956 22894 10968
rect 24302 10956 24308 11008
rect 24360 10996 24366 11008
rect 24489 10999 24547 11005
rect 24489 10996 24501 10999
rect 24360 10968 24501 10996
rect 24360 10956 24366 10968
rect 24489 10965 24501 10968
rect 24535 10965 24547 10999
rect 24489 10959 24547 10965
rect 25130 10956 25136 11008
rect 25188 10996 25194 11008
rect 26878 10996 26884 11008
rect 25188 10968 26884 10996
rect 25188 10956 25194 10968
rect 26878 10956 26884 10968
rect 26936 10956 26942 11008
rect 26973 10999 27031 11005
rect 26973 10965 26985 10999
rect 27019 10996 27031 10999
rect 27522 10996 27528 11008
rect 27019 10968 27528 10996
rect 27019 10965 27031 10968
rect 26973 10959 27031 10965
rect 27522 10956 27528 10968
rect 27580 10956 27586 11008
rect 27724 10996 27752 11024
rect 28537 10999 28595 11005
rect 28537 10996 28549 10999
rect 27724 10968 28549 10996
rect 28537 10965 28549 10968
rect 28583 10996 28595 10999
rect 28810 10996 28816 11008
rect 28583 10968 28816 10996
rect 28583 10965 28595 10968
rect 28537 10959 28595 10965
rect 28810 10956 28816 10968
rect 28868 10956 28874 11008
rect 29196 10996 29224 11104
rect 29365 11101 29377 11104
rect 29411 11101 29423 11135
rect 29365 11095 29423 11101
rect 29454 11092 29460 11144
rect 29512 11132 29518 11144
rect 30116 11132 30144 11163
rect 30558 11160 30564 11212
rect 30616 11160 30622 11212
rect 29512 11104 30144 11132
rect 29512 11092 29518 11104
rect 29273 11067 29331 11073
rect 29273 11033 29285 11067
rect 29319 11064 29331 11067
rect 29914 11064 29920 11076
rect 29319 11036 29920 11064
rect 29319 11033 29331 11036
rect 29273 11027 29331 11033
rect 29914 11024 29920 11036
rect 29972 11024 29978 11076
rect 31021 11067 31079 11073
rect 31021 11064 31033 11067
rect 30024 11036 31033 11064
rect 29730 10996 29736 11008
rect 29196 10968 29736 10996
rect 29730 10956 29736 10968
rect 29788 10996 29794 11008
rect 30024 10996 30052 11036
rect 31021 11033 31033 11036
rect 31067 11033 31079 11067
rect 31021 11027 31079 11033
rect 29788 10968 30052 10996
rect 29788 10956 29794 10968
rect 552 10906 31648 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 11436 10906
rect 11488 10854 11500 10906
rect 11552 10854 11564 10906
rect 11616 10854 11628 10906
rect 11680 10854 11692 10906
rect 11744 10854 19210 10906
rect 19262 10854 19274 10906
rect 19326 10854 19338 10906
rect 19390 10854 19402 10906
rect 19454 10854 19466 10906
rect 19518 10854 26984 10906
rect 27036 10854 27048 10906
rect 27100 10854 27112 10906
rect 27164 10854 27176 10906
rect 27228 10854 27240 10906
rect 27292 10854 31648 10906
rect 552 10832 31648 10854
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 3050 10792 3056 10804
rect 2924 10764 3056 10792
rect 2924 10752 2930 10764
rect 3050 10752 3056 10764
rect 3108 10792 3114 10804
rect 3786 10792 3792 10804
rect 3108 10764 3792 10792
rect 3108 10752 3114 10764
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 3881 10795 3939 10801
rect 3881 10761 3893 10795
rect 3927 10792 3939 10795
rect 4062 10792 4068 10804
rect 3927 10764 4068 10792
rect 3927 10761 3939 10764
rect 3881 10755 3939 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4798 10792 4804 10804
rect 4304 10764 4804 10792
rect 4304 10752 4310 10764
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5994 10792 6000 10804
rect 5000 10764 6000 10792
rect 1762 10684 1768 10736
rect 1820 10724 1826 10736
rect 1949 10727 2007 10733
rect 1949 10724 1961 10727
rect 1820 10696 1961 10724
rect 1820 10684 1826 10696
rect 1949 10693 1961 10696
rect 1995 10693 2007 10727
rect 5000 10724 5028 10764
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6086 10752 6092 10804
rect 6144 10752 6150 10804
rect 6825 10795 6883 10801
rect 6196 10764 6776 10792
rect 1949 10687 2007 10693
rect 2746 10696 5028 10724
rect 5077 10727 5135 10733
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2590 10656 2596 10668
rect 2087 10628 2596 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2590 10616 2596 10628
rect 2648 10656 2654 10668
rect 2746 10656 2774 10696
rect 5077 10693 5089 10727
rect 5123 10724 5135 10727
rect 5258 10724 5264 10736
rect 5123 10696 5264 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 2648 10628 2774 10656
rect 3160 10628 3985 10656
rect 2648 10616 2654 10628
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 2774 10588 2780 10600
rect 1811 10560 2780 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 2774 10548 2780 10560
rect 2832 10588 2838 10600
rect 3160 10588 3188 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 5166 10656 5172 10668
rect 3973 10619 4031 10625
rect 4099 10628 5028 10656
rect 2832 10560 3188 10588
rect 2832 10548 2838 10560
rect 3234 10548 3240 10600
rect 3292 10548 3298 10600
rect 3330 10591 3388 10597
rect 3330 10557 3342 10591
rect 3376 10588 3388 10591
rect 3376 10560 3464 10588
rect 3376 10557 3388 10560
rect 3330 10551 3388 10557
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3252 10452 3280 10548
rect 3436 10532 3464 10560
rect 3694 10548 3700 10600
rect 3752 10597 3758 10600
rect 3752 10588 3760 10597
rect 3752 10560 3797 10588
rect 3752 10551 3760 10560
rect 3752 10548 3758 10551
rect 3418 10480 3424 10532
rect 3476 10480 3482 10532
rect 3510 10480 3516 10532
rect 3568 10480 3574 10532
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 4099 10520 4127 10628
rect 4338 10548 4344 10600
rect 4396 10548 4402 10600
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 3651 10492 4127 10520
rect 4157 10523 4215 10529
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 4157 10489 4169 10523
rect 4203 10520 4215 10523
rect 5000 10520 5028 10628
rect 5092 10628 5172 10656
rect 5092 10597 5120 10628
rect 5166 10616 5172 10628
rect 5224 10656 5230 10668
rect 5442 10656 5448 10668
rect 5224 10628 5448 10656
rect 5224 10616 5230 10628
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 6196 10665 6224 10764
rect 6457 10727 6515 10733
rect 6457 10693 6469 10727
rect 6503 10724 6515 10727
rect 6503 10696 6684 10724
rect 6503 10693 6515 10696
rect 6457 10687 6515 10693
rect 6656 10665 6684 10696
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6748 10656 6776 10764
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 6871 10764 7144 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 7009 10727 7067 10733
rect 7009 10693 7021 10727
rect 7055 10693 7067 10727
rect 7116 10724 7144 10764
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7248 10764 7757 10792
rect 7248 10752 7254 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 8018 10752 8024 10804
rect 8076 10752 8082 10804
rect 8202 10752 8208 10804
rect 8260 10752 8266 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 8352 10764 11300 10792
rect 8352 10752 8358 10764
rect 8665 10727 8723 10733
rect 8665 10724 8677 10727
rect 7116 10696 8677 10724
rect 7009 10687 7067 10693
rect 8665 10693 8677 10696
rect 8711 10693 8723 10727
rect 9306 10724 9312 10736
rect 8665 10687 8723 10693
rect 8772 10696 9312 10724
rect 7024 10656 7052 10687
rect 6748 10628 6960 10656
rect 7024 10628 7972 10656
rect 6641 10619 6699 10625
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5626 10588 5632 10600
rect 5399 10560 5632 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 5276 10520 5304 10551
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 5718 10548 5724 10600
rect 5776 10548 5782 10600
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 6089 10591 6147 10597
rect 6089 10588 6101 10591
rect 6043 10560 6101 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 6089 10557 6101 10560
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6328 10560 6561 10588
rect 6328 10548 6334 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6788 10560 6837 10588
rect 6788 10548 6794 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6932 10588 6960 10628
rect 7006 10588 7012 10600
rect 6932 10560 7012 10588
rect 6825 10551 6883 10557
rect 7006 10548 7012 10560
rect 7064 10588 7070 10600
rect 7101 10591 7159 10597
rect 7101 10588 7113 10591
rect 7064 10560 7113 10588
rect 7064 10548 7070 10560
rect 7101 10557 7113 10560
rect 7147 10557 7159 10591
rect 7101 10551 7159 10557
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 5902 10520 5908 10532
rect 4203 10492 4292 10520
rect 5000 10492 5908 10520
rect 4203 10489 4215 10492
rect 4157 10483 4215 10489
rect 2832 10424 3280 10452
rect 4264 10452 4292 10492
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 7208 10520 7236 10551
rect 7466 10548 7472 10600
rect 7524 10548 7530 10600
rect 7558 10548 7564 10600
rect 7616 10548 7622 10600
rect 6564 10492 7236 10520
rect 7377 10523 7435 10529
rect 6564 10464 6592 10492
rect 7377 10489 7389 10523
rect 7423 10520 7435 10523
rect 7742 10520 7748 10532
rect 7423 10492 7748 10520
rect 7423 10489 7435 10492
rect 7377 10483 7435 10489
rect 7742 10480 7748 10492
rect 7800 10480 7806 10532
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10489 7895 10523
rect 7944 10520 7972 10628
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 8772 10656 8800 10696
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9582 10684 9588 10736
rect 9640 10724 9646 10736
rect 9769 10727 9827 10733
rect 9769 10724 9781 10727
rect 9640 10696 9781 10724
rect 9640 10684 9646 10696
rect 9769 10693 9781 10696
rect 9815 10693 9827 10727
rect 9769 10687 9827 10693
rect 9876 10696 10548 10724
rect 8260 10628 8800 10656
rect 8260 10616 8266 10628
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9490 10656 9496 10668
rect 9171 10628 9496 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9876 10656 9904 10696
rect 10410 10656 10416 10668
rect 9600 10628 9904 10656
rect 10060 10628 10416 10656
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 8037 10523 8095 10529
rect 8037 10520 8049 10523
rect 7944 10492 8049 10520
rect 7837 10483 7895 10489
rect 8037 10489 8049 10492
rect 8083 10489 8095 10523
rect 8037 10483 8095 10489
rect 4890 10452 4896 10464
rect 4264 10424 4896 10452
rect 2832 10412 2838 10424
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5534 10412 5540 10464
rect 5592 10412 5598 10464
rect 5629 10455 5687 10461
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 6178 10452 6184 10464
rect 5675 10424 6184 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6546 10412 6552 10464
rect 6604 10412 6610 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7852 10452 7880 10483
rect 8754 10480 8760 10532
rect 8812 10520 8818 10532
rect 8864 10520 8892 10551
rect 9214 10548 9220 10600
rect 9272 10548 9278 10600
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 9364 10560 9413 10588
rect 9364 10548 9370 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9493 10523 9551 10529
rect 9493 10520 9505 10523
rect 8812 10492 9505 10520
rect 8812 10480 8818 10492
rect 9493 10489 9505 10492
rect 9539 10489 9551 10523
rect 9493 10483 9551 10489
rect 9600 10452 9628 10628
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 9766 10588 9772 10600
rect 9723 10560 9772 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9858 10548 9864 10600
rect 9916 10548 9922 10600
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 9968 10520 9996 10551
rect 9692 10492 9996 10520
rect 9692 10464 9720 10492
rect 6972 10424 9628 10452
rect 6972 10412 6978 10424
rect 9674 10412 9680 10464
rect 9732 10412 9738 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10060 10452 10088 10628
rect 10410 10616 10416 10628
rect 10468 10616 10474 10668
rect 10134 10548 10140 10600
rect 10192 10548 10198 10600
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 10520 10597 10548 10696
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 10962 10724 10968 10736
rect 10744 10696 10968 10724
rect 10744 10684 10750 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 11272 10724 11300 10764
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11388 10764 17080 10792
rect 11388 10752 11394 10764
rect 11698 10724 11704 10736
rect 11272 10696 11704 10724
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 13170 10724 13176 10736
rect 12676 10696 13176 10724
rect 12676 10684 12682 10696
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 15286 10724 15292 10736
rect 13372 10696 15292 10724
rect 10612 10628 11468 10656
rect 10505 10591 10563 10597
rect 10505 10557 10517 10591
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 10244 10520 10272 10548
rect 10612 10520 10640 10628
rect 10781 10591 10839 10597
rect 10689 10585 10747 10591
rect 10689 10578 10701 10585
rect 10735 10578 10747 10585
rect 10686 10526 10692 10578
rect 10744 10526 10750 10578
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10244 10492 10640 10520
rect 9824 10424 10088 10452
rect 9824 10412 9830 10424
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10796 10452 10824 10551
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11330 10591 11388 10597
rect 11330 10588 11342 10591
rect 11287 10560 11342 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11330 10557 11342 10560
rect 11376 10557 11388 10591
rect 11440 10588 11468 10628
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 12526 10656 12532 10668
rect 11624 10628 12532 10656
rect 11624 10588 11652 10628
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 11440 10560 11652 10588
rect 11330 10551 11388 10557
rect 11072 10520 11100 10551
rect 11698 10548 11704 10600
rect 11756 10548 11762 10600
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10588 11851 10591
rect 13372 10588 13400 10696
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 15378 10684 15384 10736
rect 15436 10684 15442 10736
rect 15562 10733 15568 10736
rect 15519 10727 15568 10733
rect 15519 10693 15531 10727
rect 15565 10693 15568 10727
rect 15519 10687 15568 10693
rect 15562 10684 15568 10687
rect 15620 10684 15626 10736
rect 15657 10727 15715 10733
rect 15657 10693 15669 10727
rect 15703 10724 15715 10727
rect 15930 10724 15936 10736
rect 15703 10696 15936 10724
rect 15703 10693 15715 10696
rect 15657 10687 15715 10693
rect 15930 10684 15936 10696
rect 15988 10724 15994 10736
rect 16298 10724 16304 10736
rect 15988 10696 16304 10724
rect 15988 10684 15994 10696
rect 16298 10684 16304 10696
rect 16356 10684 16362 10736
rect 17052 10724 17080 10764
rect 17126 10752 17132 10804
rect 17184 10752 17190 10804
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 17770 10792 17776 10804
rect 17460 10764 17776 10792
rect 17460 10752 17466 10764
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 19429 10795 19487 10801
rect 19429 10761 19441 10795
rect 19475 10792 19487 10795
rect 19475 10764 22140 10792
rect 19475 10761 19487 10764
rect 19429 10755 19487 10761
rect 20162 10724 20168 10736
rect 17052 10696 20168 10724
rect 20162 10684 20168 10696
rect 20220 10684 20226 10736
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 20772 10696 20852 10724
rect 20772 10684 20778 10696
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 15194 10656 15200 10668
rect 14568 10628 15200 10656
rect 11839 10560 13400 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13633 10591 13691 10597
rect 13633 10588 13645 10591
rect 13504 10560 13645 10588
rect 13504 10548 13510 10560
rect 13633 10557 13645 10560
rect 13679 10557 13691 10591
rect 13633 10551 13691 10557
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 14182 10548 14188 10600
rect 14240 10548 14246 10600
rect 14458 10548 14464 10600
rect 14516 10548 14522 10600
rect 14568 10597 14596 10628
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15396 10656 15424 10684
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15396 10628 15761 10656
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 16482 10616 16488 10668
rect 16540 10656 16546 10668
rect 19702 10656 19708 10668
rect 16540 10628 19708 10656
rect 16540 10616 16546 10628
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14734 10548 14740 10600
rect 14792 10548 14798 10600
rect 15381 10591 15439 10597
rect 15381 10588 15393 10591
rect 15166 10560 15393 10588
rect 10888 10492 11100 10520
rect 10888 10464 10916 10492
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 13354 10520 13360 10532
rect 11940 10492 13360 10520
rect 11940 10480 11946 10492
rect 13354 10480 13360 10492
rect 13412 10520 13418 10532
rect 15166 10520 15194 10560
rect 15381 10557 15393 10560
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 15838 10548 15844 10600
rect 15896 10548 15902 10600
rect 16758 10588 16764 10600
rect 15948 10560 16764 10588
rect 13412 10492 15194 10520
rect 13412 10480 13418 10492
rect 15286 10480 15292 10532
rect 15344 10520 15350 10532
rect 15948 10520 15976 10560
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 16850 10548 16856 10600
rect 16908 10588 16914 10600
rect 17512 10597 17540 10628
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 20346 10656 20352 10668
rect 19996 10628 20352 10656
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 16908 10560 17417 10588
rect 16908 10548 16914 10560
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 17497 10591 17555 10597
rect 17497 10557 17509 10591
rect 17543 10557 17555 10591
rect 17497 10551 17555 10557
rect 17586 10548 17592 10600
rect 17644 10548 17650 10600
rect 17770 10548 17776 10600
rect 17828 10548 17834 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 15344 10492 15976 10520
rect 15344 10480 15350 10492
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 16080 10492 16804 10520
rect 16080 10480 16086 10492
rect 10284 10424 10824 10452
rect 10284 10412 10290 10424
rect 10870 10412 10876 10464
rect 10928 10412 10934 10464
rect 11514 10412 11520 10464
rect 11572 10412 11578 10464
rect 11606 10412 11612 10464
rect 11664 10412 11670 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12158 10452 12164 10464
rect 11756 10424 12164 10452
rect 11756 10412 11762 10424
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 12618 10412 12624 10464
rect 12676 10452 12682 10464
rect 12986 10452 12992 10464
rect 12676 10424 12992 10452
rect 12676 10412 12682 10424
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 13228 10424 14657 10452
rect 13228 10412 13234 10424
rect 14645 10421 14657 10424
rect 14691 10452 14703 10455
rect 16666 10452 16672 10464
rect 14691 10424 16672 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16776 10452 16804 10492
rect 17862 10480 17868 10532
rect 17920 10520 17926 10532
rect 18340 10520 18368 10551
rect 18506 10548 18512 10600
rect 18564 10548 18570 10600
rect 18874 10548 18880 10600
rect 18932 10548 18938 10600
rect 19150 10597 19156 10600
rect 19149 10588 19156 10597
rect 19111 10560 19156 10588
rect 19149 10551 19156 10560
rect 19150 10548 19156 10551
rect 19208 10548 19214 10600
rect 19996 10597 20024 10628
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20438 10616 20444 10668
rect 20496 10616 20502 10668
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 17920 10492 18368 10520
rect 18417 10523 18475 10529
rect 17920 10480 17926 10492
rect 18417 10489 18429 10523
rect 18463 10520 18475 10523
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 18463 10492 19073 10520
rect 18463 10489 18475 10492
rect 18417 10483 18475 10489
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19061 10483 19119 10489
rect 17957 10455 18015 10461
rect 17957 10452 17969 10455
rect 16776 10424 17969 10452
rect 17957 10421 17969 10424
rect 18003 10421 18015 10455
rect 17957 10415 18015 10421
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19260 10452 19288 10551
rect 19610 10480 19616 10532
rect 19668 10520 19674 10532
rect 20073 10523 20131 10529
rect 19668 10492 19840 10520
rect 19668 10480 19674 10492
rect 18748 10424 19288 10452
rect 18748 10412 18754 10424
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19702 10452 19708 10464
rect 19392 10424 19708 10452
rect 19392 10412 19398 10424
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 19812 10461 19840 10492
rect 20073 10489 20085 10523
rect 20119 10489 20131 10523
rect 20073 10483 20131 10489
rect 19797 10455 19855 10461
rect 19797 10421 19809 10455
rect 19843 10421 19855 10455
rect 19797 10415 19855 10421
rect 19886 10412 19892 10464
rect 19944 10452 19950 10464
rect 20088 10452 20116 10483
rect 20162 10480 20168 10532
rect 20220 10529 20226 10532
rect 20220 10523 20236 10529
rect 20224 10489 20236 10523
rect 20220 10483 20236 10489
rect 20283 10523 20341 10529
rect 20283 10489 20295 10523
rect 20329 10520 20341 10523
rect 20438 10520 20444 10566
rect 20329 10514 20444 10520
rect 20496 10514 20502 10566
rect 20824 10520 20852 10696
rect 21266 10684 21272 10736
rect 21324 10684 21330 10736
rect 22112 10724 22140 10764
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22336 10764 22385 10792
rect 22336 10752 22342 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 23014 10752 23020 10804
rect 23072 10752 23078 10804
rect 23290 10752 23296 10804
rect 23348 10792 23354 10804
rect 23937 10795 23995 10801
rect 23937 10792 23949 10795
rect 23348 10764 23949 10792
rect 23348 10752 23354 10764
rect 23937 10761 23949 10764
rect 23983 10761 23995 10795
rect 23937 10755 23995 10761
rect 24026 10752 24032 10804
rect 24084 10792 24090 10804
rect 24765 10795 24823 10801
rect 24765 10792 24777 10795
rect 24084 10764 24777 10792
rect 24084 10752 24090 10764
rect 24765 10761 24777 10764
rect 24811 10792 24823 10795
rect 24811 10764 25636 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25608 10724 25636 10764
rect 25682 10752 25688 10804
rect 25740 10792 25746 10804
rect 25777 10795 25835 10801
rect 25777 10792 25789 10795
rect 25740 10764 25789 10792
rect 25740 10752 25746 10764
rect 25777 10761 25789 10764
rect 25823 10761 25835 10795
rect 26418 10792 26424 10804
rect 25777 10755 25835 10761
rect 25976 10764 26424 10792
rect 25976 10724 26004 10764
rect 26418 10752 26424 10764
rect 26476 10752 26482 10804
rect 27617 10795 27675 10801
rect 27617 10761 27629 10795
rect 27663 10792 27675 10795
rect 28074 10792 28080 10804
rect 27663 10764 28080 10792
rect 27663 10761 27675 10764
rect 27617 10755 27675 10761
rect 28074 10752 28080 10764
rect 28132 10752 28138 10804
rect 22112 10696 24808 10724
rect 25608 10696 26004 10724
rect 20990 10616 20996 10668
rect 21048 10656 21054 10668
rect 21048 10628 21588 10656
rect 21048 10616 21054 10628
rect 21450 10548 21456 10600
rect 21508 10548 21514 10600
rect 21560 10597 21588 10628
rect 21910 10616 21916 10668
rect 21968 10656 21974 10668
rect 24673 10659 24731 10665
rect 24673 10656 24685 10659
rect 21968 10628 24685 10656
rect 21968 10616 21974 10628
rect 24673 10625 24685 10628
rect 24719 10625 24731 10659
rect 24780 10656 24808 10696
rect 26050 10684 26056 10736
rect 26108 10724 26114 10736
rect 26605 10727 26663 10733
rect 26605 10724 26617 10727
rect 26108 10696 26617 10724
rect 26108 10684 26114 10696
rect 26605 10693 26617 10696
rect 26651 10693 26663 10727
rect 26605 10687 26663 10693
rect 26694 10684 26700 10736
rect 26752 10684 26758 10736
rect 26786 10684 26792 10736
rect 26844 10724 26850 10736
rect 27157 10727 27215 10733
rect 27157 10724 27169 10727
rect 26844 10696 27169 10724
rect 26844 10684 26850 10696
rect 27157 10693 27169 10696
rect 27203 10693 27215 10727
rect 27157 10687 27215 10693
rect 27433 10727 27491 10733
rect 27433 10693 27445 10727
rect 27479 10724 27491 10727
rect 27706 10724 27712 10736
rect 27479 10696 27712 10724
rect 27479 10693 27491 10696
rect 27433 10687 27491 10693
rect 27706 10684 27712 10696
rect 27764 10684 27770 10736
rect 30374 10684 30380 10736
rect 30432 10684 30438 10736
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 24780 10628 26157 10656
rect 24673 10619 24731 10625
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26712 10656 26740 10684
rect 29178 10656 29184 10668
rect 26145 10619 26203 10625
rect 26620 10628 26740 10656
rect 27356 10628 29184 10656
rect 21545 10591 21603 10597
rect 21545 10557 21557 10591
rect 21591 10557 21603 10591
rect 21545 10551 21603 10557
rect 21634 10548 21640 10600
rect 21692 10588 21698 10600
rect 21729 10591 21787 10597
rect 21729 10588 21741 10591
rect 21692 10560 21741 10588
rect 21692 10548 21698 10560
rect 21729 10557 21741 10560
rect 21775 10557 21787 10591
rect 21729 10551 21787 10557
rect 21818 10548 21824 10600
rect 21876 10548 21882 10600
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22649 10591 22707 10597
rect 22649 10588 22661 10591
rect 22244 10560 22661 10588
rect 22244 10548 22250 10560
rect 22649 10557 22661 10560
rect 22695 10557 22707 10591
rect 22649 10551 22707 10557
rect 22830 10548 22836 10600
rect 22888 10588 22894 10600
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22888 10560 23121 10588
rect 22888 10548 22894 10560
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23109 10551 23167 10557
rect 24118 10548 24124 10600
rect 24176 10548 24182 10600
rect 24213 10591 24271 10597
rect 24213 10557 24225 10591
rect 24259 10588 24271 10591
rect 24394 10588 24400 10600
rect 24259 10560 24400 10588
rect 24259 10557 24271 10560
rect 24213 10551 24271 10557
rect 24394 10548 24400 10560
rect 24452 10548 24458 10600
rect 24489 10591 24547 10597
rect 24489 10557 24501 10591
rect 24535 10557 24547 10591
rect 24489 10551 24547 10557
rect 23290 10520 23296 10532
rect 20329 10492 20484 10514
rect 20824 10492 23296 10520
rect 20329 10489 20341 10492
rect 20283 10483 20341 10489
rect 20220 10480 20226 10483
rect 23290 10480 23296 10492
rect 23348 10480 23354 10532
rect 24302 10480 24308 10532
rect 24360 10480 24366 10532
rect 24504 10520 24532 10551
rect 24578 10548 24584 10600
rect 24636 10548 24642 10600
rect 24946 10548 24952 10600
rect 25004 10548 25010 10600
rect 25958 10548 25964 10600
rect 26016 10548 26022 10600
rect 26237 10591 26295 10597
rect 26237 10557 26249 10591
rect 26283 10557 26295 10591
rect 26237 10551 26295 10557
rect 25133 10523 25191 10529
rect 25133 10520 25145 10523
rect 24504 10492 25145 10520
rect 25133 10489 25145 10492
rect 25179 10489 25191 10523
rect 25133 10483 25191 10489
rect 26142 10480 26148 10532
rect 26200 10520 26206 10532
rect 26252 10520 26280 10551
rect 26326 10548 26332 10600
rect 26384 10548 26390 10600
rect 26418 10548 26424 10600
rect 26476 10548 26482 10600
rect 26620 10597 26648 10628
rect 26605 10591 26663 10597
rect 26605 10557 26617 10591
rect 26651 10557 26663 10591
rect 26605 10551 26663 10557
rect 26697 10591 26755 10597
rect 26697 10557 26709 10591
rect 26743 10557 26755 10591
rect 26697 10551 26755 10557
rect 26712 10520 26740 10551
rect 26878 10548 26884 10600
rect 26936 10588 26942 10600
rect 27356 10597 27384 10628
rect 29178 10616 29184 10628
rect 29236 10656 29242 10668
rect 29236 10628 30052 10656
rect 29236 10616 29242 10628
rect 27341 10591 27399 10597
rect 27341 10588 27353 10591
rect 26936 10560 27353 10588
rect 26936 10548 26942 10560
rect 27341 10557 27353 10560
rect 27387 10557 27399 10591
rect 27890 10588 27896 10600
rect 27341 10551 27399 10557
rect 27448 10560 27896 10588
rect 26200 10492 26280 10520
rect 26344 10492 26740 10520
rect 26200 10480 26206 10492
rect 19944 10424 20116 10452
rect 20181 10452 20209 10480
rect 22554 10452 22560 10464
rect 20181 10424 22560 10452
rect 19944 10412 19950 10424
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 22738 10412 22744 10464
rect 22796 10412 22802 10464
rect 22833 10455 22891 10461
rect 22833 10421 22845 10455
rect 22879 10452 22891 10455
rect 25498 10452 25504 10464
rect 22879 10424 25504 10452
rect 22879 10421 22891 10424
rect 22833 10415 22891 10421
rect 25498 10412 25504 10424
rect 25556 10412 25562 10464
rect 25590 10412 25596 10464
rect 25648 10452 25654 10464
rect 26344 10452 26372 10492
rect 27062 10480 27068 10532
rect 27120 10520 27126 10532
rect 27448 10520 27476 10560
rect 27890 10548 27896 10560
rect 27948 10548 27954 10600
rect 28629 10591 28687 10597
rect 28629 10557 28641 10591
rect 28675 10588 28687 10591
rect 28994 10588 29000 10600
rect 28675 10560 29000 10588
rect 28675 10557 28687 10560
rect 28629 10551 28687 10557
rect 28994 10548 29000 10560
rect 29052 10548 29058 10600
rect 29270 10548 29276 10600
rect 29328 10588 29334 10600
rect 30024 10597 30052 10628
rect 29457 10591 29515 10597
rect 29457 10588 29469 10591
rect 29328 10560 29469 10588
rect 29328 10548 29334 10560
rect 29457 10557 29469 10560
rect 29503 10557 29515 10591
rect 29457 10551 29515 10557
rect 30009 10591 30067 10597
rect 30009 10557 30021 10591
rect 30055 10588 30067 10591
rect 30190 10588 30196 10600
rect 30055 10560 30196 10588
rect 30055 10557 30067 10560
rect 30009 10551 30067 10557
rect 30190 10548 30196 10560
rect 30248 10548 30254 10600
rect 30282 10548 30288 10600
rect 30340 10588 30346 10600
rect 30377 10591 30435 10597
rect 30377 10588 30389 10591
rect 30340 10560 30389 10588
rect 30340 10548 30346 10560
rect 30377 10557 30389 10560
rect 30423 10557 30435 10591
rect 30377 10551 30435 10557
rect 30650 10548 30656 10600
rect 30708 10548 30714 10600
rect 31018 10548 31024 10600
rect 31076 10548 31082 10600
rect 27120 10492 27476 10520
rect 27120 10480 27126 10492
rect 27522 10480 27528 10532
rect 27580 10529 27586 10532
rect 27580 10523 27643 10529
rect 27580 10489 27597 10523
rect 27631 10489 27643 10523
rect 27580 10483 27643 10489
rect 27801 10523 27859 10529
rect 27801 10489 27813 10523
rect 27847 10520 27859 10523
rect 27908 10520 27936 10548
rect 27847 10492 27936 10520
rect 27847 10489 27859 10492
rect 27801 10483 27859 10489
rect 27580 10480 27586 10483
rect 28442 10480 28448 10532
rect 28500 10520 28506 10532
rect 29178 10520 29184 10532
rect 28500 10492 29184 10520
rect 28500 10480 28506 10492
rect 29178 10480 29184 10492
rect 29236 10480 29242 10532
rect 29733 10523 29791 10529
rect 29733 10489 29745 10523
rect 29779 10520 29791 10523
rect 31110 10520 31116 10532
rect 29779 10492 31116 10520
rect 29779 10489 29791 10492
rect 29733 10483 29791 10489
rect 31110 10480 31116 10492
rect 31168 10480 31174 10532
rect 25648 10424 26372 10452
rect 26881 10455 26939 10461
rect 25648 10412 25654 10424
rect 26881 10421 26893 10455
rect 26927 10452 26939 10455
rect 26970 10452 26976 10464
rect 26927 10424 26976 10452
rect 26927 10421 26939 10424
rect 26881 10415 26939 10421
rect 26970 10412 26976 10424
rect 27028 10412 27034 10464
rect 27154 10412 27160 10464
rect 27212 10452 27218 10464
rect 28074 10452 28080 10464
rect 27212 10424 28080 10452
rect 27212 10412 27218 10424
rect 28074 10412 28080 10424
rect 28132 10452 28138 10464
rect 28626 10452 28632 10464
rect 28132 10424 28632 10452
rect 28132 10412 28138 10424
rect 28626 10412 28632 10424
rect 28684 10412 28690 10464
rect 28810 10412 28816 10464
rect 28868 10412 28874 10464
rect 29273 10455 29331 10461
rect 29273 10421 29285 10455
rect 29319 10452 29331 10455
rect 30098 10452 30104 10464
rect 29319 10424 30104 10452
rect 29319 10421 29331 10424
rect 29273 10415 29331 10421
rect 30098 10412 30104 10424
rect 30156 10412 30162 10464
rect 552 10362 31648 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 12096 10362
rect 12148 10310 12160 10362
rect 12212 10310 12224 10362
rect 12276 10310 12288 10362
rect 12340 10310 12352 10362
rect 12404 10310 19870 10362
rect 19922 10310 19934 10362
rect 19986 10310 19998 10362
rect 20050 10310 20062 10362
rect 20114 10310 20126 10362
rect 20178 10310 27644 10362
rect 27696 10310 27708 10362
rect 27760 10310 27772 10362
rect 27824 10310 27836 10362
rect 27888 10310 27900 10362
rect 27952 10310 31648 10362
rect 552 10288 31648 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 1360 10220 3617 10248
rect 1360 10208 1366 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 3786 10208 3792 10260
rect 3844 10208 3850 10260
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 6273 10251 6331 10257
rect 6273 10248 6285 10251
rect 5960 10220 6285 10248
rect 5960 10208 5966 10220
rect 6273 10217 6285 10220
rect 6319 10217 6331 10251
rect 7006 10248 7012 10260
rect 6273 10211 6331 10217
rect 6380 10220 7012 10248
rect 3513 10183 3571 10189
rect 3513 10149 3525 10183
rect 3559 10180 3571 10183
rect 4798 10180 4804 10192
rect 3559 10152 4804 10180
rect 3559 10149 3571 10152
rect 3513 10143 3571 10149
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 6380 10180 6408 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 7156 10220 8309 10248
rect 7156 10208 7162 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9214 10248 9220 10260
rect 9079 10220 9220 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9674 10248 9680 10260
rect 9324 10220 9680 10248
rect 6104 10152 6408 10180
rect 3234 10072 3240 10124
rect 3292 10112 3298 10124
rect 3421 10115 3479 10121
rect 3421 10112 3433 10115
rect 3292 10084 3433 10112
rect 3292 10072 3298 10084
rect 3421 10081 3433 10084
rect 3467 10081 3479 10115
rect 3421 10075 3479 10081
rect 3878 10072 3884 10124
rect 3936 10072 3942 10124
rect 4157 10115 4215 10121
rect 4157 10081 4169 10115
rect 4203 10112 4215 10115
rect 4338 10112 4344 10124
rect 4203 10084 4344 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 1854 10004 1860 10056
rect 1912 10044 1918 10056
rect 2314 10044 2320 10056
rect 1912 10016 2320 10044
rect 1912 10004 1918 10016
rect 2314 10004 2320 10016
rect 2372 10044 2378 10056
rect 4172 10044 4200 10075
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 5258 10112 5264 10124
rect 4580 10084 5264 10112
rect 4580 10072 4586 10084
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 6104 10112 6132 10152
rect 6454 10140 6460 10192
rect 6512 10180 6518 10192
rect 6914 10180 6920 10192
rect 6512 10152 6920 10180
rect 6512 10140 6518 10152
rect 6914 10140 6920 10152
rect 6972 10180 6978 10192
rect 6972 10152 7321 10180
rect 6972 10140 6978 10152
rect 5552 10084 6132 10112
rect 2372 10016 4200 10044
rect 2372 10004 2378 10016
rect 4246 10004 4252 10056
rect 4304 10004 4310 10056
rect 5552 10044 5580 10084
rect 6178 10072 6184 10124
rect 6236 10072 6242 10124
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7190 10112 7196 10124
rect 7055 10084 7196 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7293 10112 7321 10152
rect 7558 10140 7564 10192
rect 7616 10180 7622 10192
rect 9324 10180 9352 10220
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10134 10248 10140 10260
rect 9784 10220 10140 10248
rect 7616 10152 9168 10180
rect 7616 10140 7622 10152
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 7293 10084 7665 10112
rect 7653 10081 7665 10084
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8665 10115 8723 10121
rect 8527 10084 8616 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 4816 10016 5580 10044
rect 3237 9979 3295 9985
rect 3237 9945 3249 9979
rect 3283 9976 3295 9979
rect 3418 9976 3424 9988
rect 3283 9948 3424 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 3418 9936 3424 9948
rect 3476 9976 3482 9988
rect 4816 9976 4844 10016
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 6641 10047 6699 10053
rect 6641 10044 6653 10047
rect 5684 10016 6653 10044
rect 5684 10004 5690 10016
rect 6641 10013 6653 10016
rect 6687 10044 6699 10047
rect 7374 10044 7380 10056
rect 6687 10016 7380 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 8202 10044 8208 10056
rect 7524 10016 8208 10044
rect 7524 10004 7530 10016
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 3476 9948 4844 9976
rect 3476 9936 3482 9948
rect 4890 9936 4896 9988
rect 4948 9976 4954 9988
rect 8588 9976 8616 10084
rect 8665 10081 8677 10115
rect 8711 10112 8723 10115
rect 9030 10112 9036 10124
rect 8711 10084 9036 10112
rect 8711 10081 8723 10084
rect 8665 10075 8723 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 8754 10004 8760 10056
rect 8812 10004 8818 10056
rect 9140 10044 9168 10152
rect 9232 10152 9352 10180
rect 9232 10121 9260 10152
rect 9398 10140 9404 10192
rect 9456 10180 9462 10192
rect 9456 10152 9536 10180
rect 9456 10140 9462 10152
rect 9508 10121 9536 10152
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9493 10115 9551 10121
rect 9355 10084 9444 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9416 10056 9444 10084
rect 9493 10081 9505 10115
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9784 10112 9812 10220
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 10226 10208 10232 10260
rect 10284 10208 10290 10260
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 10744 10220 10977 10248
rect 10744 10208 10750 10220
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13998 10248 14004 10260
rect 12492 10220 14004 10248
rect 12492 10208 12498 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14826 10248 14832 10260
rect 14476 10220 14832 10248
rect 9953 10183 10011 10189
rect 9953 10149 9965 10183
rect 9999 10180 10011 10183
rect 10594 10180 10600 10192
rect 9999 10152 10600 10180
rect 9999 10149 10011 10152
rect 9953 10143 10011 10149
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 12618 10180 12624 10192
rect 10704 10152 12624 10180
rect 10704 10124 10732 10152
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13078 10180 13084 10192
rect 12728 10152 13084 10180
rect 9723 10084 9812 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 9858 10072 9864 10124
rect 9916 10072 9922 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9968 10084 10057 10112
rect 9140 10016 9352 10044
rect 9214 9976 9220 9988
rect 4948 9948 8524 9976
rect 8588 9948 9220 9976
rect 4948 9936 4954 9948
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 6822 9908 6828 9920
rect 3660 9880 6828 9908
rect 3660 9868 3666 9880
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 7745 9911 7803 9917
rect 7745 9908 7757 9911
rect 7248 9880 7757 9908
rect 7248 9868 7254 9880
rect 7745 9877 7757 9880
rect 7791 9877 7803 9911
rect 8496 9908 8524 9948
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9324 9976 9352 10016
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 9968 9976 9996 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10502 10112 10508 10124
rect 10284 10084 10508 10112
rect 10284 10072 10290 10084
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10081 11115 10115
rect 11057 10075 11115 10081
rect 11425 10115 11483 10121
rect 11425 10081 11437 10115
rect 11471 10112 11483 10115
rect 12728 10112 12756 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 14476 10189 14504 10220
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 16666 10248 16672 10260
rect 14976 10220 16672 10248
rect 14976 10208 14982 10220
rect 16666 10208 16672 10220
rect 16724 10208 16730 10260
rect 17586 10248 17592 10260
rect 17052 10220 17592 10248
rect 14461 10183 14519 10189
rect 14461 10149 14473 10183
rect 14507 10149 14519 10183
rect 14461 10143 14519 10149
rect 14553 10183 14611 10189
rect 14553 10149 14565 10183
rect 14599 10180 14611 10183
rect 14734 10180 14740 10192
rect 14599 10152 14740 10180
rect 14599 10149 14611 10152
rect 14553 10143 14611 10149
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 15838 10180 15844 10192
rect 14936 10152 15844 10180
rect 11471 10084 12756 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10870 10044 10876 10056
rect 10376 10016 10876 10044
rect 10376 10004 10382 10016
rect 10870 10004 10876 10016
rect 10928 10044 10934 10056
rect 11072 10044 11100 10075
rect 12894 10072 12900 10124
rect 12952 10072 12958 10124
rect 12986 10072 12992 10124
rect 13044 10072 13050 10124
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13446 10112 13452 10124
rect 13311 10084 13452 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14323 10115 14381 10121
rect 14323 10112 14335 10115
rect 13872 10084 14335 10112
rect 13872 10072 13878 10084
rect 14323 10081 14335 10084
rect 14369 10081 14381 10115
rect 14323 10075 14381 10081
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10081 14703 10115
rect 14936 10112 14964 10152
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 16022 10140 16028 10192
rect 16080 10180 16086 10192
rect 16945 10183 17003 10189
rect 16080 10152 16530 10180
rect 16080 10140 16086 10152
rect 14645 10075 14703 10081
rect 14764 10084 14964 10112
rect 10928 10016 11100 10044
rect 11149 10047 11207 10053
rect 10928 10004 10934 10016
rect 11149 10013 11161 10047
rect 11195 10044 11207 10047
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 11195 10016 12725 10044
rect 11195 10013 11207 10016
rect 11149 10007 11207 10013
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 12820 10016 13814 10044
rect 11882 9976 11888 9988
rect 9324 9948 11888 9976
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 12342 9936 12348 9988
rect 12400 9976 12406 9988
rect 12820 9976 12848 10016
rect 12400 9948 12848 9976
rect 13786 9976 13814 10016
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13964 10016 14197 10044
rect 13964 10004 13970 10016
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14185 10007 14243 10013
rect 14550 10004 14556 10056
rect 14608 10044 14614 10056
rect 14660 10044 14688 10075
rect 14608 10016 14688 10044
rect 14608 10004 14614 10016
rect 14764 9976 14792 10084
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10044 14887 10047
rect 15010 10044 15016 10056
rect 14875 10016 15016 10044
rect 14875 10013 14887 10016
rect 14829 10007 14887 10013
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15856 10044 15884 10140
rect 16502 10121 16530 10152
rect 16945 10149 16957 10183
rect 16991 10180 17003 10183
rect 17052 10180 17080 10220
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 20990 10248 20996 10260
rect 18156 10220 20996 10248
rect 16991 10152 17080 10180
rect 17129 10183 17187 10189
rect 16991 10149 17003 10152
rect 16945 10143 17003 10149
rect 17129 10149 17141 10183
rect 17175 10180 17187 10183
rect 17770 10180 17776 10192
rect 17175 10152 17776 10180
rect 17175 10149 17187 10152
rect 17129 10143 17187 10149
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 16574 10072 16580 10124
rect 16632 10112 16638 10124
rect 17037 10115 17095 10121
rect 17037 10112 17049 10115
rect 16632 10084 17049 10112
rect 16632 10072 16638 10084
rect 17037 10081 17049 10084
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 17221 10115 17279 10121
rect 17221 10081 17233 10115
rect 17267 10112 17279 10115
rect 18156 10112 18184 10220
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 21082 10208 21088 10260
rect 21140 10208 21146 10260
rect 21634 10208 21640 10260
rect 21692 10208 21698 10260
rect 21836 10220 23704 10248
rect 18322 10140 18328 10192
rect 18380 10180 18386 10192
rect 20714 10180 20720 10192
rect 18380 10152 20720 10180
rect 18380 10140 18386 10152
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 21100 10180 21128 10208
rect 20824 10152 21128 10180
rect 17267 10084 18184 10112
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 15856 10016 16773 10044
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 16850 10004 16856 10056
rect 16908 10004 16914 10056
rect 13786 9948 14792 9976
rect 12400 9936 12406 9948
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 16577 9979 16635 9985
rect 16577 9976 16589 9979
rect 15344 9948 16589 9976
rect 15344 9936 15350 9948
rect 16577 9945 16589 9948
rect 16623 9945 16635 9979
rect 16577 9939 16635 9945
rect 17034 9936 17040 9988
rect 17092 9976 17098 9988
rect 17236 9976 17264 10075
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18506 10112 18512 10124
rect 18288 10084 18512 10112
rect 18288 10072 18294 10084
rect 18506 10072 18512 10084
rect 18564 10112 18570 10124
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18564 10084 18981 10112
rect 18564 10072 18570 10084
rect 18969 10081 18981 10084
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 19153 10115 19211 10121
rect 19153 10081 19165 10115
rect 19199 10112 19211 10115
rect 20622 10112 20628 10124
rect 19199 10084 20628 10112
rect 19199 10081 19211 10084
rect 19153 10075 19211 10081
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 20824 10121 20852 10152
rect 20809 10115 20867 10121
rect 20809 10081 20821 10115
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 20898 10072 20904 10124
rect 20956 10072 20962 10124
rect 21085 10115 21143 10121
rect 21085 10081 21097 10115
rect 21131 10112 21143 10115
rect 21634 10112 21640 10124
rect 21131 10084 21640 10112
rect 21131 10081 21143 10084
rect 21085 10075 21143 10081
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 21836 10121 21864 10220
rect 22186 10180 22192 10192
rect 22020 10152 22192 10180
rect 22020 10121 22048 10152
rect 22186 10140 22192 10152
rect 22244 10140 22250 10192
rect 22554 10140 22560 10192
rect 22612 10180 22618 10192
rect 22925 10183 22983 10189
rect 22925 10180 22937 10183
rect 22612 10152 22937 10180
rect 22612 10140 22618 10152
rect 22925 10149 22937 10152
rect 22971 10180 22983 10183
rect 23106 10180 23112 10192
rect 22971 10152 23112 10180
rect 22971 10149 22983 10152
rect 22925 10143 22983 10149
rect 23106 10140 23112 10152
rect 23164 10140 23170 10192
rect 21821 10115 21879 10121
rect 21821 10081 21833 10115
rect 21867 10081 21879 10115
rect 21821 10075 21879 10081
rect 22005 10115 22063 10121
rect 22005 10081 22017 10115
rect 22051 10081 22063 10115
rect 22005 10075 22063 10081
rect 22094 10072 22100 10124
rect 22152 10072 22158 10124
rect 23014 10072 23020 10124
rect 23072 10072 23078 10124
rect 23290 10072 23296 10124
rect 23348 10072 23354 10124
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19242 10044 19248 10056
rect 18380 10016 19248 10044
rect 18380 10004 18386 10016
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19334 10004 19340 10056
rect 19392 10004 19398 10056
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 20990 10044 20996 10056
rect 19484 10016 20996 10044
rect 19484 10004 19490 10016
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 21100 10016 21925 10044
rect 17092 9948 17264 9976
rect 17092 9936 17098 9948
rect 17770 9936 17776 9988
rect 17828 9976 17834 9988
rect 19150 9976 19156 9988
rect 17828 9948 19156 9976
rect 17828 9936 17834 9948
rect 19150 9936 19156 9948
rect 19208 9936 19214 9988
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9976 19763 9979
rect 21100 9976 21128 10016
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 21913 10007 21971 10013
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 23032 10044 23060 10072
rect 22612 10016 23060 10044
rect 22612 10004 22618 10016
rect 22830 9976 22836 9988
rect 19751 9948 21128 9976
rect 21560 9948 22836 9976
rect 19751 9945 19763 9948
rect 19705 9939 19763 9945
rect 8846 9908 8852 9920
rect 8496 9880 8852 9908
rect 7745 9871 7803 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9490 9908 9496 9920
rect 8996 9880 9496 9908
rect 8996 9868 9002 9880
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 11146 9908 11152 9920
rect 9916 9880 11152 9908
rect 9916 9868 9922 9880
rect 11146 9868 11152 9880
rect 11204 9908 11210 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 11204 9880 11345 9908
rect 11204 9868 11210 9880
rect 11333 9877 11345 9880
rect 11379 9877 11391 9911
rect 11333 9871 11391 9877
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 13722 9908 13728 9920
rect 11572 9880 13728 9908
rect 11572 9868 11578 9880
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 15378 9908 15384 9920
rect 14792 9880 15384 9908
rect 14792 9868 14798 9880
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 16666 9868 16672 9920
rect 16724 9908 16730 9920
rect 17310 9908 17316 9920
rect 16724 9880 17316 9908
rect 16724 9868 16730 9880
rect 17310 9868 17316 9880
rect 17368 9908 17374 9920
rect 21560 9908 21588 9948
rect 22830 9936 22836 9948
rect 22888 9936 22894 9988
rect 23676 9976 23704 10220
rect 23842 10208 23848 10260
rect 23900 10208 23906 10260
rect 24026 10257 24032 10260
rect 24013 10251 24032 10257
rect 24013 10217 24025 10251
rect 24013 10211 24032 10217
rect 24026 10208 24032 10211
rect 24084 10208 24090 10260
rect 24673 10251 24731 10257
rect 24673 10217 24685 10251
rect 24719 10248 24731 10251
rect 24719 10220 24992 10248
rect 24719 10217 24731 10220
rect 24673 10211 24731 10217
rect 24210 10140 24216 10192
rect 24268 10140 24274 10192
rect 24302 10140 24308 10192
rect 24360 10180 24366 10192
rect 24964 10180 24992 10220
rect 25038 10208 25044 10260
rect 25096 10248 25102 10260
rect 26237 10251 26295 10257
rect 25096 10220 26170 10248
rect 25096 10208 25102 10220
rect 25590 10180 25596 10192
rect 24360 10152 24900 10180
rect 24964 10152 25596 10180
rect 24360 10140 24366 10152
rect 23750 10072 23756 10124
rect 23808 10112 23814 10124
rect 24872 10121 24900 10152
rect 25056 10124 25084 10152
rect 25590 10140 25596 10152
rect 25648 10140 25654 10192
rect 25958 10180 25964 10192
rect 25792 10152 25964 10180
rect 24489 10115 24547 10121
rect 24489 10112 24501 10115
rect 23808 10084 24501 10112
rect 23808 10072 23814 10084
rect 24489 10081 24501 10084
rect 24535 10081 24547 10115
rect 24489 10075 24547 10081
rect 24857 10115 24915 10121
rect 24857 10081 24869 10115
rect 24903 10081 24915 10115
rect 24857 10075 24915 10081
rect 25038 10072 25044 10124
rect 25096 10072 25102 10124
rect 25792 10121 25820 10152
rect 25958 10140 25964 10152
rect 26016 10140 26022 10192
rect 25777 10115 25835 10121
rect 25777 10081 25789 10115
rect 25823 10081 25835 10115
rect 25777 10075 25835 10081
rect 26050 10072 26056 10124
rect 26108 10072 26114 10124
rect 26142 10112 26170 10220
rect 26237 10217 26249 10251
rect 26283 10217 26295 10251
rect 26237 10211 26295 10217
rect 26252 10180 26280 10211
rect 26418 10208 26424 10260
rect 26476 10248 26482 10260
rect 26476 10220 29868 10248
rect 26476 10208 26482 10220
rect 26252 10152 28488 10180
rect 26142 10084 27200 10112
rect 24394 10004 24400 10056
rect 24452 10004 24458 10056
rect 24762 10004 24768 10056
rect 24820 10004 24826 10056
rect 25869 10047 25927 10053
rect 25869 10013 25881 10047
rect 25915 10013 25927 10047
rect 25869 10007 25927 10013
rect 25590 9976 25596 9988
rect 23676 9948 25596 9976
rect 25590 9936 25596 9948
rect 25648 9936 25654 9988
rect 25884 9976 25912 10007
rect 25958 10004 25964 10056
rect 26016 10004 26022 10056
rect 26602 10004 26608 10056
rect 26660 10004 26666 10056
rect 26697 10047 26755 10053
rect 26697 10013 26709 10047
rect 26743 10013 26755 10047
rect 26697 10007 26755 10013
rect 26789 10047 26847 10053
rect 26789 10013 26801 10047
rect 26835 10013 26847 10047
rect 26789 10007 26847 10013
rect 26881 10047 26939 10053
rect 26881 10013 26893 10047
rect 26927 10044 26939 10047
rect 27065 10047 27123 10053
rect 27065 10044 27077 10047
rect 26927 10016 27077 10044
rect 26927 10013 26939 10016
rect 26881 10007 26939 10013
rect 27065 10013 27077 10016
rect 27111 10013 27123 10047
rect 27172 10044 27200 10084
rect 27246 10072 27252 10124
rect 27304 10072 27310 10124
rect 27522 10072 27528 10124
rect 27580 10072 27586 10124
rect 28166 10072 28172 10124
rect 28224 10072 28230 10124
rect 28460 10121 28488 10152
rect 29178 10140 29184 10192
rect 29236 10180 29242 10192
rect 29365 10183 29423 10189
rect 29365 10180 29377 10183
rect 29236 10152 29377 10180
rect 29236 10140 29242 10152
rect 29365 10149 29377 10152
rect 29411 10149 29423 10183
rect 29365 10143 29423 10149
rect 28445 10115 28503 10121
rect 28445 10081 28457 10115
rect 28491 10081 28503 10115
rect 28445 10075 28503 10081
rect 28721 10115 28779 10121
rect 28721 10081 28733 10115
rect 28767 10081 28779 10115
rect 28721 10075 28779 10081
rect 28997 10115 29055 10121
rect 28997 10081 29009 10115
rect 29043 10112 29055 10115
rect 29454 10112 29460 10124
rect 29043 10084 29460 10112
rect 29043 10081 29055 10084
rect 28997 10075 29055 10081
rect 27540 10044 27568 10072
rect 27172 10016 27568 10044
rect 27065 10007 27123 10013
rect 26421 9979 26479 9985
rect 26421 9976 26433 9979
rect 25884 9948 26433 9976
rect 26421 9945 26433 9948
rect 26467 9945 26479 9979
rect 26421 9939 26479 9945
rect 26510 9936 26516 9988
rect 26568 9976 26574 9988
rect 26712 9976 26740 10007
rect 26568 9948 26740 9976
rect 26804 9976 26832 10007
rect 27982 10004 27988 10056
rect 28040 10004 28046 10056
rect 28258 10004 28264 10056
rect 28316 10004 28322 10056
rect 28350 10004 28356 10056
rect 28408 10004 28414 10056
rect 26970 9976 26976 9988
rect 26804 9948 26976 9976
rect 26568 9936 26574 9948
rect 26970 9936 26976 9948
rect 27028 9936 27034 9988
rect 27154 9936 27160 9988
rect 27212 9976 27218 9988
rect 27341 9979 27399 9985
rect 27341 9976 27353 9979
rect 27212 9948 27353 9976
rect 27212 9936 27218 9948
rect 27341 9945 27353 9948
rect 27387 9945 27399 9979
rect 27341 9939 27399 9945
rect 27433 9979 27491 9985
rect 27433 9945 27445 9979
rect 27479 9945 27491 9979
rect 27433 9939 27491 9945
rect 17368 9880 21588 9908
rect 17368 9868 17374 9880
rect 21634 9868 21640 9920
rect 21692 9908 21698 9920
rect 23566 9908 23572 9920
rect 21692 9880 23572 9908
rect 21692 9868 21698 9880
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 23934 9868 23940 9920
rect 23992 9908 23998 9920
rect 24029 9911 24087 9917
rect 24029 9908 24041 9911
rect 23992 9880 24041 9908
rect 23992 9868 23998 9880
rect 24029 9877 24041 9880
rect 24075 9877 24087 9911
rect 24029 9871 24087 9877
rect 24762 9868 24768 9920
rect 24820 9908 24826 9920
rect 25041 9911 25099 9917
rect 25041 9908 25053 9911
rect 24820 9880 25053 9908
rect 24820 9868 24826 9880
rect 25041 9877 25053 9880
rect 25087 9877 25099 9911
rect 25041 9871 25099 9877
rect 25314 9868 25320 9920
rect 25372 9908 25378 9920
rect 25774 9908 25780 9920
rect 25372 9880 25780 9908
rect 25372 9868 25378 9880
rect 25774 9868 25780 9880
rect 25832 9868 25838 9920
rect 26326 9868 26332 9920
rect 26384 9908 26390 9920
rect 27448 9908 27476 9939
rect 26384 9880 27476 9908
rect 26384 9868 26390 9880
rect 28074 9868 28080 9920
rect 28132 9908 28138 9920
rect 28736 9908 28764 10075
rect 29454 10072 29460 10084
rect 29512 10072 29518 10124
rect 29546 10072 29552 10124
rect 29604 10072 29610 10124
rect 29641 10115 29699 10121
rect 29641 10081 29653 10115
rect 29687 10081 29699 10115
rect 29641 10075 29699 10081
rect 29270 10004 29276 10056
rect 29328 10044 29334 10056
rect 29656 10044 29684 10075
rect 29730 10072 29736 10124
rect 29788 10072 29794 10124
rect 29840 10121 29868 10220
rect 30190 10208 30196 10260
rect 30248 10248 30254 10260
rect 30248 10220 30972 10248
rect 30248 10208 30254 10220
rect 29914 10140 29920 10192
rect 29972 10180 29978 10192
rect 30282 10180 30288 10192
rect 29972 10152 30288 10180
rect 29972 10140 29978 10152
rect 30282 10140 30288 10152
rect 30340 10180 30346 10192
rect 30340 10152 30696 10180
rect 30340 10140 30346 10152
rect 29825 10115 29883 10121
rect 29825 10081 29837 10115
rect 29871 10081 29883 10115
rect 29825 10075 29883 10081
rect 30098 10072 30104 10124
rect 30156 10072 30162 10124
rect 30190 10072 30196 10124
rect 30248 10072 30254 10124
rect 30668 10121 30696 10152
rect 30377 10115 30435 10121
rect 30377 10112 30389 10115
rect 30300 10084 30389 10112
rect 29328 10016 29684 10044
rect 30300 10044 30328 10084
rect 30377 10081 30389 10084
rect 30423 10081 30435 10115
rect 30377 10075 30435 10081
rect 30653 10115 30711 10121
rect 30653 10081 30665 10115
rect 30699 10081 30711 10115
rect 30653 10075 30711 10081
rect 30834 10072 30840 10124
rect 30892 10072 30898 10124
rect 30944 10121 30972 10220
rect 30929 10115 30987 10121
rect 30929 10081 30941 10115
rect 30975 10081 30987 10115
rect 30929 10075 30987 10081
rect 31021 10115 31079 10121
rect 31021 10081 31033 10115
rect 31067 10081 31079 10115
rect 31021 10075 31079 10081
rect 31036 10044 31064 10075
rect 30300 10016 31064 10044
rect 29328 10004 29334 10016
rect 28810 9936 28816 9988
rect 28868 9976 28874 9988
rect 30300 9976 30328 10016
rect 28868 9948 30328 9976
rect 28868 9936 28874 9948
rect 30834 9936 30840 9988
rect 30892 9976 30898 9988
rect 31662 9976 31668 9988
rect 30892 9948 31668 9976
rect 30892 9936 30898 9948
rect 31662 9936 31668 9948
rect 31720 9936 31726 9988
rect 28132 9880 28764 9908
rect 29365 9911 29423 9917
rect 28132 9868 28138 9880
rect 29365 9877 29377 9911
rect 29411 9908 29423 9911
rect 29638 9908 29644 9920
rect 29411 9880 29644 9908
rect 29411 9877 29423 9880
rect 29365 9871 29423 9877
rect 29638 9868 29644 9880
rect 29696 9868 29702 9920
rect 30190 9868 30196 9920
rect 30248 9908 30254 9920
rect 31110 9908 31116 9920
rect 30248 9880 31116 9908
rect 30248 9868 30254 9880
rect 31110 9868 31116 9880
rect 31168 9868 31174 9920
rect 31294 9868 31300 9920
rect 31352 9868 31358 9920
rect 552 9818 31648 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 11436 9818
rect 11488 9766 11500 9818
rect 11552 9766 11564 9818
rect 11616 9766 11628 9818
rect 11680 9766 11692 9818
rect 11744 9766 19210 9818
rect 19262 9766 19274 9818
rect 19326 9766 19338 9818
rect 19390 9766 19402 9818
rect 19454 9766 19466 9818
rect 19518 9766 26984 9818
rect 27036 9766 27048 9818
rect 27100 9766 27112 9818
rect 27164 9766 27176 9818
rect 27228 9766 27240 9818
rect 27292 9766 31648 9818
rect 552 9744 31648 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 1765 9707 1823 9713
rect 1765 9704 1777 9707
rect 1636 9676 1777 9704
rect 1636 9664 1642 9676
rect 1765 9673 1777 9676
rect 1811 9673 1823 9707
rect 1765 9667 1823 9673
rect 3234 9664 3240 9716
rect 3292 9664 3298 9716
rect 4246 9704 4252 9716
rect 4080 9676 4252 9704
rect 1302 9596 1308 9648
rect 1360 9596 1366 9648
rect 1210 9528 1216 9580
rect 1268 9568 1274 9580
rect 4080 9568 4108 9676
rect 4246 9664 4252 9676
rect 4304 9664 4310 9716
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5442 9704 5448 9716
rect 4948 9676 5448 9704
rect 4948 9664 4954 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 5905 9707 5963 9713
rect 5776 9676 5856 9704
rect 5776 9664 5782 9676
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 4580 9608 4752 9636
rect 4580 9596 4586 9608
rect 1268 9540 1624 9568
rect 1268 9528 1274 9540
rect 1026 9460 1032 9512
rect 1084 9500 1090 9512
rect 1596 9509 1624 9540
rect 3528 9540 4108 9568
rect 1489 9503 1547 9509
rect 1489 9500 1501 9503
rect 1084 9472 1501 9500
rect 1084 9460 1090 9472
rect 1489 9469 1501 9472
rect 1535 9469 1547 9503
rect 1489 9463 1547 9469
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9469 1639 9503
rect 1581 9463 1639 9469
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2038 9500 2044 9512
rect 1903 9472 2044 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2038 9460 2044 9472
rect 2096 9500 2102 9512
rect 2682 9500 2688 9512
rect 2096 9472 2688 9500
rect 2096 9460 2102 9472
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3528 9509 3556 9540
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3108 9472 3433 9500
rect 3108 9460 3114 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 3694 9460 3700 9512
rect 3752 9460 3758 9512
rect 3786 9460 3792 9512
rect 3844 9460 3850 9512
rect 4724 9509 4752 9608
rect 4798 9596 4804 9648
rect 4856 9596 4862 9648
rect 5828 9636 5856 9676
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6454 9704 6460 9716
rect 5951 9676 6460 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 8021 9707 8079 9713
rect 8021 9673 8033 9707
rect 8067 9704 8079 9707
rect 8110 9704 8116 9716
rect 8067 9676 8116 9704
rect 8067 9673 8079 9676
rect 8021 9667 8079 9673
rect 7653 9639 7711 9645
rect 5828 9608 6316 9636
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5442 9568 5448 9580
rect 5399 9540 5448 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5776 9540 6193 9568
rect 5776 9528 5782 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9469 4767 9503
rect 4709 9463 4767 9469
rect 4798 9460 4804 9512
rect 4856 9500 4862 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4856 9472 4905 9500
rect 4856 9460 4862 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 5184 9432 5212 9463
rect 5626 9460 5632 9512
rect 5684 9460 5690 9512
rect 5994 9460 6000 9512
rect 6052 9460 6058 9512
rect 5258 9432 5264 9444
rect 3016 9404 5120 9432
rect 5184 9404 5264 9432
rect 3016 9392 3022 9404
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1854 9364 1860 9376
rect 1544 9336 1860 9364
rect 1544 9324 1550 9336
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 4430 9364 4436 9376
rect 3752 9336 4436 9364
rect 3752 9324 3758 9336
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4764 9336 4997 9364
rect 4764 9324 4770 9336
rect 4985 9333 4997 9336
rect 5031 9333 5043 9367
rect 5092 9364 5120 9404
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 5442 9392 5448 9444
rect 5500 9392 5506 9444
rect 5537 9435 5595 9441
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 5810 9432 5816 9444
rect 5583 9404 5816 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9401 5963 9435
rect 5905 9395 5963 9401
rect 5920 9364 5948 9395
rect 6288 9364 6316 9608
rect 7653 9605 7665 9639
rect 7699 9636 7711 9639
rect 8036 9636 8064 9667
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 9582 9704 9588 9716
rect 8777 9676 9588 9704
rect 8777 9636 8805 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 9824 9676 10732 9704
rect 9824 9664 9830 9676
rect 7699 9608 8064 9636
rect 8220 9608 8805 9636
rect 7699 9605 7711 9608
rect 7653 9599 7711 9605
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 6880 9540 7512 9568
rect 6880 9528 6886 9540
rect 7484 9512 7512 9540
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 8220 9577 8248 9608
rect 8846 9596 8852 9648
rect 8904 9596 8910 9648
rect 8941 9639 8999 9645
rect 8941 9605 8953 9639
rect 8987 9636 8999 9639
rect 9122 9636 9128 9648
rect 8987 9608 9128 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 9600 9636 9628 9664
rect 10704 9636 10732 9676
rect 11330 9664 11336 9716
rect 11388 9664 11394 9716
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11480 9676 12204 9704
rect 11480 9664 11486 9676
rect 12066 9636 12072 9648
rect 9600 9608 10640 9636
rect 10704 9608 12072 9636
rect 8205 9571 8263 9577
rect 7800 9540 8064 9568
rect 7800 9528 7806 9540
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6972 9472 7021 9500
rect 6972 9460 6978 9472
rect 7009 9469 7021 9472
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 7156 9472 7205 9500
rect 7156 9460 7162 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 7834 9500 7840 9512
rect 7524 9472 7840 9500
rect 7524 9460 7530 9472
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9469 7987 9503
rect 8036 9500 8064 9540
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 8205 9531 8263 9537
rect 8680 9540 9965 9568
rect 8680 9500 8708 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10502 9568 10508 9580
rect 10459 9540 10508 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 8036 9472 8708 9500
rect 7929 9463 7987 9469
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6733 9435 6791 9441
rect 6733 9432 6745 9435
rect 6420 9404 6745 9432
rect 6420 9392 6426 9404
rect 6733 9401 6745 9404
rect 6779 9401 6791 9435
rect 7944 9432 7972 9463
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 9030 9460 9036 9512
rect 9088 9460 9094 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9306 9500 9312 9512
rect 9263 9472 9312 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 10612 9509 10640 9608
rect 12066 9596 12072 9608
rect 12124 9596 12130 9648
rect 12176 9636 12204 9676
rect 12342 9664 12348 9716
rect 12400 9664 12406 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 13081 9707 13139 9713
rect 12492 9676 12756 9704
rect 12492 9664 12498 9676
rect 12621 9639 12679 9645
rect 12621 9636 12633 9639
rect 12176 9608 12633 9636
rect 12621 9605 12633 9608
rect 12667 9605 12679 9639
rect 12621 9599 12679 9605
rect 12728 9577 12756 9676
rect 13081 9673 13093 9707
rect 13127 9704 13139 9707
rect 13814 9704 13820 9716
rect 13127 9676 13820 9704
rect 13127 9673 13139 9676
rect 13081 9667 13139 9673
rect 13814 9664 13820 9676
rect 13872 9704 13878 9716
rect 13872 9676 17264 9704
rect 13872 9664 13878 9676
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13170 9636 13176 9648
rect 13044 9608 13176 9636
rect 13044 9596 13050 9608
rect 13170 9596 13176 9608
rect 13228 9596 13234 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 14001 9639 14059 9645
rect 14001 9636 14013 9639
rect 13964 9608 14013 9636
rect 13964 9596 13970 9608
rect 14001 9605 14013 9608
rect 14047 9605 14059 9639
rect 14001 9599 14059 9605
rect 14182 9596 14188 9648
rect 14240 9636 14246 9648
rect 14366 9636 14372 9648
rect 14240 9608 14372 9636
rect 14240 9596 14246 9608
rect 14366 9596 14372 9608
rect 14424 9596 14430 9648
rect 14550 9596 14556 9648
rect 14608 9636 14614 9648
rect 15010 9636 15016 9648
rect 14608 9608 15016 9636
rect 14608 9596 14614 9608
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15252 9608 15516 9636
rect 15252 9596 15258 9608
rect 12713 9571 12771 9577
rect 11272 9540 11920 9568
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9456 9472 9781 9500
rect 9456 9460 9462 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9500 10195 9503
rect 10597 9503 10655 9509
rect 10183 9472 10548 9500
rect 10183 9469 10195 9472
rect 10137 9463 10195 9469
rect 8110 9432 8116 9444
rect 7944 9404 8116 9432
rect 6733 9395 6791 9401
rect 8110 9392 8116 9404
rect 8168 9432 8174 9444
rect 9493 9435 9551 9441
rect 9493 9432 9505 9435
rect 8168 9404 9505 9432
rect 8168 9392 8174 9404
rect 9493 9401 9505 9404
rect 9539 9401 9551 9435
rect 9784 9432 9812 9463
rect 10520 9432 10548 9472
rect 10597 9469 10609 9503
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 11272 9432 11300 9540
rect 11514 9460 11520 9512
rect 11572 9460 11578 9512
rect 11790 9460 11796 9512
rect 11848 9460 11854 9512
rect 11892 9500 11920 9540
rect 12713 9537 12725 9571
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9537 12863 9571
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 12805 9531 12863 9537
rect 12912 9540 15301 9568
rect 12529 9503 12587 9509
rect 12529 9502 12541 9503
rect 12452 9500 12541 9502
rect 11892 9474 12541 9500
rect 11892 9472 12480 9474
rect 12529 9469 12541 9474
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12676 9494 12756 9500
rect 12820 9494 12848 9531
rect 12676 9472 12848 9494
rect 12676 9460 12682 9472
rect 12728 9466 12848 9472
rect 9784 9404 10272 9432
rect 10520 9404 11300 9432
rect 11624 9404 12020 9432
rect 9493 9395 9551 9401
rect 6822 9364 6828 9376
rect 5092 9336 6828 9364
rect 4985 9327 5043 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 7248 9336 7297 9364
rect 7248 9324 7254 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 7285 9327 7343 9333
rect 8202 9324 8208 9376
rect 8260 9324 8266 9376
rect 8386 9324 8392 9376
rect 8444 9364 8450 9376
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 8444 9336 8585 9364
rect 8444 9324 8450 9336
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8573 9327 8631 9333
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 9306 9364 9312 9376
rect 8812 9336 9312 9364
rect 8812 9324 8818 9336
rect 9306 9324 9312 9336
rect 9364 9364 9370 9376
rect 10134 9364 10140 9376
rect 9364 9336 10140 9364
rect 9364 9324 9370 9336
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10244 9364 10272 9404
rect 10612 9376 10640 9404
rect 10502 9364 10508 9376
rect 10244 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10594 9324 10600 9376
rect 10652 9324 10658 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 11624 9364 11652 9404
rect 10744 9336 11652 9364
rect 10744 9324 10750 9336
rect 11698 9324 11704 9376
rect 11756 9324 11762 9376
rect 11992 9364 12020 9404
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 12912 9432 12940 9540
rect 15289 9537 15301 9540
rect 15335 9568 15347 9571
rect 15378 9568 15384 9580
rect 15335 9540 15384 9568
rect 15335 9537 15347 9540
rect 15289 9531 15347 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 15488 9568 15516 9608
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 15896 9608 15945 9636
rect 15896 9596 15902 9608
rect 15933 9605 15945 9608
rect 15979 9605 15991 9639
rect 15933 9599 15991 9605
rect 16942 9596 16948 9648
rect 17000 9636 17006 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 17000 9608 17141 9636
rect 17000 9596 17006 9608
rect 17129 9605 17141 9608
rect 17175 9605 17187 9639
rect 17236 9636 17264 9676
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 18230 9704 18236 9716
rect 17828 9676 18236 9704
rect 17828 9664 17834 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 18782 9704 18788 9716
rect 18656 9676 18788 9704
rect 18656 9664 18662 9676
rect 18782 9664 18788 9676
rect 18840 9704 18846 9716
rect 18840 9676 19380 9704
rect 18840 9664 18846 9676
rect 19150 9636 19156 9648
rect 17236 9608 19156 9636
rect 17129 9599 17187 9605
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 19352 9636 19380 9676
rect 19426 9664 19432 9716
rect 19484 9704 19490 9716
rect 19484 9676 19932 9704
rect 19484 9664 19490 9676
rect 19904 9636 19932 9676
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20073 9707 20131 9713
rect 20073 9704 20085 9707
rect 20036 9676 20085 9704
rect 20036 9664 20042 9676
rect 20073 9673 20085 9676
rect 20119 9673 20131 9707
rect 20898 9704 20904 9716
rect 20073 9667 20131 9673
rect 20180 9676 20904 9704
rect 20180 9636 20208 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 21818 9664 21824 9716
rect 21876 9704 21882 9716
rect 22005 9707 22063 9713
rect 22005 9704 22017 9707
rect 21876 9676 22017 9704
rect 21876 9664 21882 9676
rect 22005 9673 22017 9676
rect 22051 9673 22063 9707
rect 22005 9667 22063 9673
rect 22738 9664 22744 9716
rect 22796 9704 22802 9716
rect 22833 9707 22891 9713
rect 22833 9704 22845 9707
rect 22796 9676 22845 9704
rect 22796 9664 22802 9676
rect 22833 9673 22845 9676
rect 22879 9673 22891 9707
rect 22833 9667 22891 9673
rect 23750 9664 23756 9716
rect 23808 9704 23814 9716
rect 25406 9704 25412 9716
rect 23808 9676 25412 9704
rect 23808 9664 23814 9676
rect 25406 9664 25412 9676
rect 25464 9664 25470 9716
rect 25498 9664 25504 9716
rect 25556 9704 25562 9716
rect 25556 9676 26648 9704
rect 25556 9664 25562 9676
rect 21450 9636 21456 9648
rect 19352 9608 19860 9636
rect 19904 9608 20208 9636
rect 20456 9608 21456 9636
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 15488 9540 16221 9568
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 17770 9568 17776 9580
rect 16724 9540 17080 9568
rect 16724 9528 16730 9540
rect 12986 9460 12992 9512
rect 13044 9460 13050 9512
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9500 13323 9503
rect 13311 9472 13492 9500
rect 13311 9469 13323 9472
rect 13265 9463 13323 9469
rect 12124 9404 12940 9432
rect 13096 9432 13124 9463
rect 13354 9432 13360 9444
rect 13096 9404 13360 9432
rect 12124 9392 12130 9404
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 13464 9364 13492 9472
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13780 9472 13921 9500
rect 13780 9460 13786 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9500 14151 9503
rect 14826 9500 14872 9502
rect 15194 9500 15200 9512
rect 14139 9472 15200 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 16390 9509 16396 9512
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15304 9472 15485 9500
rect 15304 9444 15332 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 16347 9503 16396 9509
rect 16347 9469 16359 9503
rect 16393 9469 16396 9503
rect 16347 9463 16396 9469
rect 16390 9460 16396 9463
rect 16448 9460 16454 9512
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 14277 9435 14335 9441
rect 14277 9432 14289 9435
rect 14240 9404 14289 9432
rect 14240 9392 14246 9404
rect 14277 9401 14289 9404
rect 14323 9401 14335 9435
rect 14550 9432 14556 9444
rect 14277 9395 14335 9401
rect 14384 9404 14556 9432
rect 14384 9373 14412 9404
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 14829 9435 14887 9441
rect 14829 9401 14841 9435
rect 14875 9401 14887 9435
rect 14829 9395 14887 9401
rect 14369 9367 14427 9373
rect 14369 9364 14381 9367
rect 11992 9336 14381 9364
rect 14369 9333 14381 9336
rect 14415 9333 14427 9367
rect 14369 9327 14427 9333
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 14844 9364 14872 9395
rect 15286 9392 15292 9444
rect 15344 9392 15350 9444
rect 17052 9432 17080 9540
rect 17604 9540 17776 9568
rect 17218 9460 17224 9512
rect 17276 9500 17282 9512
rect 17604 9509 17632 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17972 9540 18874 9568
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 17276 9472 17417 9500
rect 17276 9460 17282 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17405 9463 17463 9469
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 17589 9463 17647 9469
rect 17681 9503 17739 9509
rect 17681 9469 17693 9503
rect 17727 9500 17739 9503
rect 17862 9500 17868 9512
rect 17727 9472 17868 9500
rect 17727 9469 17739 9472
rect 17681 9463 17739 9469
rect 17696 9432 17724 9463
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 17052 9404 17724 9432
rect 17770 9392 17776 9444
rect 17828 9432 17834 9444
rect 17972 9441 18000 9540
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18230 9500 18236 9512
rect 18095 9472 18236 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18322 9460 18328 9512
rect 18380 9500 18386 9512
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 18380 9472 18705 9500
rect 18380 9460 18386 9472
rect 18693 9469 18705 9472
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 18846 9441 18874 9540
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19024 9540 19288 9568
rect 19024 9528 19030 9540
rect 19150 9460 19156 9512
rect 19208 9460 19214 9512
rect 19260 9500 19288 9540
rect 19334 9528 19340 9580
rect 19392 9528 19398 9580
rect 19832 9568 19860 9608
rect 19832 9540 19932 9568
rect 19429 9503 19487 9509
rect 19429 9500 19441 9503
rect 19260 9472 19441 9500
rect 19429 9469 19441 9472
rect 19475 9469 19487 9503
rect 19429 9463 19487 9469
rect 19518 9460 19524 9512
rect 19576 9500 19582 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19576 9472 19625 9500
rect 19576 9460 19582 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19702 9460 19708 9512
rect 19760 9460 19766 9512
rect 19817 9503 19875 9509
rect 19817 9469 19829 9503
rect 19863 9469 19875 9503
rect 19817 9463 19875 9469
rect 17957 9435 18015 9441
rect 17957 9432 17969 9435
rect 17828 9404 17969 9432
rect 17828 9392 17834 9404
rect 17957 9401 17969 9404
rect 18003 9401 18015 9435
rect 18846 9435 18909 9441
rect 18846 9404 18863 9435
rect 17957 9395 18015 9401
rect 18851 9401 18863 9404
rect 18897 9401 18909 9435
rect 18851 9395 18909 9401
rect 18966 9392 18972 9444
rect 19024 9392 19030 9444
rect 19058 9392 19064 9444
rect 19116 9392 19122 9444
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 19832 9432 19860 9463
rect 19392 9404 19860 9432
rect 19904 9432 19932 9540
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 20128 9540 20269 9568
rect 20128 9528 20134 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 20346 9460 20352 9512
rect 20404 9500 20410 9512
rect 20456 9509 20484 9608
rect 21450 9596 21456 9608
rect 21508 9596 21514 9648
rect 21729 9639 21787 9645
rect 21729 9605 21741 9639
rect 21775 9636 21787 9639
rect 22281 9639 22339 9645
rect 22281 9636 22293 9639
rect 21775 9608 22293 9636
rect 21775 9605 21787 9608
rect 21729 9599 21787 9605
rect 22281 9605 22293 9608
rect 22327 9605 22339 9639
rect 22281 9599 22339 9605
rect 23106 9596 23112 9648
rect 23164 9636 23170 9648
rect 23164 9608 25084 9636
rect 23164 9596 23170 9608
rect 20990 9568 20996 9580
rect 20640 9540 20996 9568
rect 20441 9503 20499 9509
rect 20441 9500 20453 9503
rect 20404 9472 20453 9500
rect 20404 9460 20410 9472
rect 20441 9469 20453 9472
rect 20487 9469 20499 9503
rect 20441 9463 20499 9469
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 20640 9500 20668 9540
rect 20990 9528 20996 9540
rect 21048 9568 21054 9580
rect 21634 9568 21640 9580
rect 21048 9540 21640 9568
rect 21048 9528 21054 9540
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 25056 9568 25084 9608
rect 25222 9596 25228 9648
rect 25280 9596 25286 9648
rect 26510 9596 26516 9648
rect 26568 9596 26574 9648
rect 26620 9636 26648 9676
rect 26786 9664 26792 9716
rect 26844 9664 26850 9716
rect 27249 9707 27307 9713
rect 27249 9704 27261 9707
rect 26889 9676 27261 9704
rect 26889 9636 26917 9676
rect 27249 9673 27261 9676
rect 27295 9673 27307 9707
rect 27614 9704 27620 9716
rect 27249 9667 27307 9673
rect 27540 9676 27620 9704
rect 26620 9608 26917 9636
rect 27065 9639 27123 9645
rect 27065 9605 27077 9639
rect 27111 9636 27123 9639
rect 27154 9636 27160 9648
rect 27111 9608 27160 9636
rect 27111 9605 27123 9608
rect 27065 9599 27123 9605
rect 27154 9596 27160 9608
rect 27212 9596 27218 9648
rect 27540 9636 27568 9676
rect 27614 9664 27620 9676
rect 27672 9664 27678 9716
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 28261 9707 28319 9713
rect 28261 9704 28273 9707
rect 27764 9676 28273 9704
rect 27764 9664 27770 9676
rect 28261 9673 28273 9676
rect 28307 9704 28319 9707
rect 28994 9704 29000 9716
rect 28307 9676 29000 9704
rect 28307 9673 28319 9676
rect 28261 9667 28319 9673
rect 28994 9664 29000 9676
rect 29052 9664 29058 9716
rect 29273 9639 29331 9645
rect 29273 9636 29285 9639
rect 27540 9608 29285 9636
rect 29273 9605 29285 9608
rect 29319 9605 29331 9639
rect 29273 9599 29331 9605
rect 26142 9568 26148 9580
rect 23308 9540 24992 9568
rect 25056 9540 26148 9568
rect 20717 9503 20775 9509
rect 20717 9500 20729 9503
rect 20640 9472 20729 9500
rect 20717 9469 20729 9472
rect 20763 9469 20775 9503
rect 20717 9463 20775 9469
rect 20809 9503 20867 9509
rect 20809 9469 20821 9503
rect 20855 9469 20867 9503
rect 20809 9463 20867 9469
rect 21729 9503 21787 9509
rect 21729 9469 21741 9503
rect 21775 9469 21787 9503
rect 21729 9463 21787 9469
rect 20824 9432 20852 9463
rect 20898 9432 20904 9444
rect 19904 9404 20904 9432
rect 19392 9392 19398 9404
rect 20898 9392 20904 9404
rect 20956 9392 20962 9444
rect 14516 9336 14872 9364
rect 15105 9367 15163 9373
rect 14516 9324 14522 9336
rect 15105 9333 15117 9367
rect 15151 9364 15163 9367
rect 15304 9364 15332 9392
rect 15151 9336 15332 9364
rect 15151 9333 15163 9336
rect 15105 9327 15163 9333
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 16758 9364 16764 9376
rect 15896 9336 16764 9364
rect 15896 9324 15902 9336
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17221 9367 17279 9373
rect 17221 9364 17233 9367
rect 17000 9336 17233 9364
rect 17000 9324 17006 9336
rect 17221 9333 17233 9336
rect 17267 9333 17279 9367
rect 17221 9327 17279 9333
rect 17402 9324 17408 9376
rect 17460 9364 17466 9376
rect 18598 9364 18604 9376
rect 17460 9336 18604 9364
rect 17460 9324 17466 9336
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 21744 9364 21772 9463
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 22186 9460 22192 9512
rect 22244 9460 22250 9512
rect 22373 9503 22431 9509
rect 22373 9469 22385 9503
rect 22419 9469 22431 9503
rect 22373 9463 22431 9469
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 22922 9500 22928 9512
rect 22511 9472 22928 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 19300 9336 21772 9364
rect 19300 9324 19306 9336
rect 21818 9324 21824 9376
rect 21876 9364 21882 9376
rect 22388 9364 22416 9463
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23014 9460 23020 9512
rect 23072 9460 23078 9512
rect 23308 9509 23336 9540
rect 23293 9503 23351 9509
rect 23293 9469 23305 9503
rect 23339 9469 23351 9503
rect 23293 9463 23351 9469
rect 22830 9392 22836 9444
rect 22888 9432 22894 9444
rect 23308 9432 23336 9463
rect 23566 9460 23572 9512
rect 23624 9500 23630 9512
rect 24121 9503 24179 9509
rect 24121 9500 24133 9503
rect 23624 9472 24133 9500
rect 23624 9460 23630 9472
rect 24121 9469 24133 9472
rect 24167 9469 24179 9503
rect 24121 9463 24179 9469
rect 24210 9460 24216 9512
rect 24268 9500 24274 9512
rect 24397 9503 24455 9509
rect 24397 9500 24409 9503
rect 24268 9472 24409 9500
rect 24268 9460 24274 9472
rect 24397 9469 24409 9472
rect 24443 9469 24455 9503
rect 24397 9463 24455 9469
rect 24486 9460 24492 9512
rect 24544 9460 24550 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 24964 9509 24992 9540
rect 26142 9528 26148 9540
rect 26200 9528 26206 9580
rect 26694 9528 26700 9580
rect 26752 9528 26758 9580
rect 26970 9568 26976 9580
rect 26896 9540 26976 9568
rect 24949 9503 25007 9509
rect 24949 9469 24961 9503
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 25222 9460 25228 9512
rect 25280 9460 25286 9512
rect 25501 9503 25559 9509
rect 25501 9469 25513 9503
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9500 25651 9503
rect 26050 9500 26056 9512
rect 25639 9472 26056 9500
rect 25639 9469 25651 9472
rect 25593 9463 25651 9469
rect 22888 9404 23336 9432
rect 22888 9392 22894 9404
rect 23658 9392 23664 9444
rect 23716 9432 23722 9444
rect 23716 9404 24808 9432
rect 23716 9392 23722 9404
rect 21876 9336 22416 9364
rect 21876 9324 21882 9336
rect 22922 9324 22928 9376
rect 22980 9364 22986 9376
rect 23201 9367 23259 9373
rect 23201 9364 23213 9367
rect 22980 9336 23213 9364
rect 22980 9324 22986 9336
rect 23201 9333 23213 9336
rect 23247 9364 23259 9367
rect 23842 9364 23848 9376
rect 23247 9336 23848 9364
rect 23247 9333 23259 9336
rect 23201 9327 23259 9333
rect 23842 9324 23848 9336
rect 23900 9324 23906 9376
rect 24780 9364 24808 9404
rect 24854 9392 24860 9444
rect 24912 9432 24918 9444
rect 25516 9432 25544 9463
rect 26050 9460 26056 9472
rect 26108 9460 26114 9512
rect 26237 9503 26295 9509
rect 26237 9469 26249 9503
rect 26283 9500 26295 9503
rect 26602 9500 26608 9512
rect 26283 9472 26608 9500
rect 26283 9469 26295 9472
rect 26237 9463 26295 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 26896 9509 26924 9540
rect 26970 9528 26976 9540
rect 27028 9568 27034 9580
rect 27028 9540 27476 9568
rect 27028 9528 27034 9540
rect 26881 9503 26939 9509
rect 26881 9469 26893 9503
rect 26927 9469 26939 9503
rect 26881 9463 26939 9469
rect 27154 9460 27160 9512
rect 27212 9460 27218 9512
rect 27338 9460 27344 9512
rect 27396 9460 27402 9512
rect 27448 9500 27476 9540
rect 27522 9528 27528 9580
rect 27580 9528 27586 9580
rect 27706 9568 27712 9580
rect 27632 9540 27712 9568
rect 27632 9500 27660 9540
rect 27706 9528 27712 9540
rect 27764 9528 27770 9580
rect 27982 9528 27988 9580
rect 28040 9568 28046 9580
rect 29178 9568 29184 9580
rect 28040 9540 29184 9568
rect 28040 9528 28046 9540
rect 29178 9528 29184 9540
rect 29236 9528 29242 9580
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 29917 9571 29975 9577
rect 29917 9568 29929 9571
rect 29595 9540 29929 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 29917 9537 29929 9540
rect 29963 9537 29975 9571
rect 31294 9568 31300 9580
rect 29917 9531 29975 9537
rect 30300 9540 31300 9568
rect 29270 9500 29276 9512
rect 27448 9472 27660 9500
rect 27724 9472 29276 9500
rect 25682 9432 25688 9444
rect 24912 9404 25688 9432
rect 24912 9392 24918 9404
rect 25682 9392 25688 9404
rect 25740 9392 25746 9444
rect 25774 9392 25780 9444
rect 25832 9432 25838 9444
rect 25869 9435 25927 9441
rect 25869 9432 25881 9435
rect 25832 9404 25881 9432
rect 25832 9392 25838 9404
rect 25869 9401 25881 9404
rect 25915 9401 25927 9435
rect 25869 9395 25927 9401
rect 26513 9435 26571 9441
rect 26513 9401 26525 9435
rect 26559 9432 26571 9435
rect 27724 9432 27752 9472
rect 29270 9460 29276 9472
rect 29328 9460 29334 9512
rect 29362 9460 29368 9512
rect 29420 9500 29426 9512
rect 29457 9503 29515 9509
rect 29457 9500 29469 9503
rect 29420 9472 29469 9500
rect 29420 9460 29426 9472
rect 29457 9469 29469 9472
rect 29503 9469 29515 9503
rect 29457 9463 29515 9469
rect 29638 9460 29644 9512
rect 29696 9460 29702 9512
rect 29730 9460 29736 9512
rect 29788 9460 29794 9512
rect 30190 9460 30196 9512
rect 30248 9460 30254 9512
rect 30300 9509 30328 9540
rect 31294 9528 31300 9540
rect 31352 9528 31358 9580
rect 30285 9503 30343 9509
rect 30285 9469 30297 9503
rect 30331 9469 30343 9503
rect 30285 9463 30343 9469
rect 30374 9460 30380 9512
rect 30432 9460 30438 9512
rect 30561 9503 30619 9509
rect 30561 9469 30573 9503
rect 30607 9500 30619 9503
rect 30742 9500 30748 9512
rect 30607 9472 30748 9500
rect 30607 9469 30619 9472
rect 30561 9463 30619 9469
rect 30742 9460 30748 9472
rect 30800 9460 30806 9512
rect 30837 9503 30895 9509
rect 30837 9469 30849 9503
rect 30883 9469 30895 9503
rect 30837 9463 30895 9469
rect 26559 9404 27752 9432
rect 27801 9435 27859 9441
rect 26559 9401 26571 9404
rect 26513 9395 26571 9401
rect 27801 9401 27813 9435
rect 27847 9401 27859 9435
rect 27801 9395 27859 9401
rect 28353 9435 28411 9441
rect 28353 9401 28365 9435
rect 28399 9432 28411 9435
rect 29288 9432 29316 9460
rect 30653 9435 30711 9441
rect 30653 9432 30665 9435
rect 28399 9404 29224 9432
rect 29288 9404 30665 9432
rect 28399 9401 28411 9404
rect 28353 9395 28411 9401
rect 24946 9364 24952 9376
rect 24780 9336 24952 9364
rect 24946 9324 24952 9336
rect 25004 9324 25010 9376
rect 25222 9324 25228 9376
rect 25280 9364 25286 9376
rect 25498 9364 25504 9376
rect 25280 9336 25504 9364
rect 25280 9324 25286 9336
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 26142 9324 26148 9376
rect 26200 9364 26206 9376
rect 26326 9364 26332 9376
rect 26200 9336 26332 9364
rect 26200 9324 26206 9336
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 27816 9364 27844 9395
rect 28442 9364 28448 9376
rect 27816 9336 28448 9364
rect 28442 9324 28448 9336
rect 28500 9324 28506 9376
rect 29196 9364 29224 9404
rect 30653 9401 30665 9404
rect 30699 9401 30711 9435
rect 30852 9432 30880 9463
rect 31018 9460 31024 9512
rect 31076 9460 31082 9512
rect 31110 9460 31116 9512
rect 31168 9500 31174 9512
rect 31754 9500 31760 9512
rect 31168 9472 31760 9500
rect 31168 9460 31174 9472
rect 31754 9460 31760 9472
rect 31812 9460 31818 9512
rect 31294 9432 31300 9444
rect 30852 9404 31300 9432
rect 30653 9395 30711 9401
rect 31294 9392 31300 9404
rect 31352 9392 31358 9444
rect 30834 9364 30840 9376
rect 29196 9336 30840 9364
rect 30834 9324 30840 9336
rect 30892 9324 30898 9376
rect 552 9274 31648 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 12096 9274
rect 12148 9222 12160 9274
rect 12212 9222 12224 9274
rect 12276 9222 12288 9274
rect 12340 9222 12352 9274
rect 12404 9222 19870 9274
rect 19922 9222 19934 9274
rect 19986 9222 19998 9274
rect 20050 9222 20062 9274
rect 20114 9222 20126 9274
rect 20178 9222 27644 9274
rect 27696 9222 27708 9274
rect 27760 9222 27772 9274
rect 27824 9222 27836 9274
rect 27888 9222 27900 9274
rect 27952 9222 31648 9274
rect 552 9200 31648 9222
rect 1026 9120 1032 9172
rect 1084 9120 1090 9172
rect 1762 9160 1768 9172
rect 1412 9132 1768 9160
rect 1210 8984 1216 9036
rect 1268 8984 1274 9036
rect 1412 9033 1440 9132
rect 1762 9120 1768 9132
rect 1820 9160 1826 9172
rect 2498 9160 2504 9172
rect 1820 9132 2504 9160
rect 1820 9120 1826 9132
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2590 9120 2596 9172
rect 2648 9120 2654 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 3786 9160 3792 9172
rect 3559 9132 3792 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4706 9160 4712 9172
rect 4120 9132 4712 9160
rect 4120 9120 4126 9132
rect 4706 9120 4712 9132
rect 4764 9160 4770 9172
rect 5994 9160 6000 9172
rect 4764 9132 6000 9160
rect 4764 9120 4770 9132
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 9398 9160 9404 9172
rect 6880 9132 9404 9160
rect 6880 9120 6886 9132
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 10226 9160 10232 9172
rect 9508 9132 10232 9160
rect 2608 9092 2636 9120
rect 1504 9064 2636 9092
rect 1504 9033 1532 9064
rect 2866 9052 2872 9104
rect 2924 9092 2930 9104
rect 2924 9064 5580 9092
rect 2924 9052 2930 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 8993 1547 9027
rect 1489 8987 1547 8993
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1636 8996 1961 9024
rect 1636 8984 1642 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 2958 9024 2964 9036
rect 2731 8996 2964 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3050 8984 3056 9036
rect 3108 8984 3114 9036
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 8993 3479 9027
rect 3421 8987 3479 8993
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 4062 9024 4068 9036
rect 3651 8996 4068 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 1857 8919 1915 8925
rect 1872 8820 1900 8919
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 3436 8956 3464 8987
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4522 8984 4528 9036
rect 4580 8984 4586 9036
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 4890 9024 4896 9036
rect 4755 8996 4896 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 4985 9027 5043 9033
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 5074 9024 5080 9036
rect 5031 8996 5080 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 2096 8928 3464 8956
rect 2096 8916 2102 8928
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4430 8956 4436 8968
rect 3752 8928 4436 8956
rect 3752 8916 3758 8928
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 5000 8956 5028 8987
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 9024 5227 9027
rect 5258 9024 5264 9036
rect 5215 8996 5264 9024
rect 5215 8993 5227 8996
rect 5169 8987 5227 8993
rect 4918 8928 5028 8956
rect 3237 8891 3295 8897
rect 3237 8857 3249 8891
rect 3283 8888 3295 8891
rect 4918 8888 4946 8928
rect 3283 8860 4946 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 1946 8820 1952 8832
rect 1872 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8820 2010 8832
rect 2866 8820 2872 8832
rect 2004 8792 2872 8820
rect 2004 8780 2010 8792
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 4617 8823 4675 8829
rect 4617 8789 4629 8823
rect 4663 8820 4675 8823
rect 4890 8820 4896 8832
rect 4663 8792 4896 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5074 8820 5080 8832
rect 5031 8792 5080 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5184 8820 5212 8987
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5552 8888 5580 9064
rect 5626 9052 5632 9104
rect 5684 9092 5690 9104
rect 6362 9092 6368 9104
rect 5684 9064 6368 9092
rect 5684 9052 5690 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 6549 9095 6607 9101
rect 6549 9061 6561 9095
rect 6595 9092 6607 9095
rect 6730 9092 6736 9104
rect 6595 9064 6736 9092
rect 6595 9061 6607 9064
rect 6549 9055 6607 9061
rect 6730 9052 6736 9064
rect 6788 9052 6794 9104
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 8260 9064 9168 9092
rect 8260 9052 8266 9064
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5868 8996 6285 9024
rect 5868 8984 5874 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 6288 8956 6316 8987
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6512 8996 6929 9024
rect 6512 8984 6518 8996
rect 6917 8993 6929 8996
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 8938 9024 8944 9036
rect 8720 8996 8944 9024
rect 8720 8984 8726 8996
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9140 9033 9168 9064
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 9214 8984 9220 9036
rect 9272 8984 9278 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9508 9033 9536 9132
rect 10226 9120 10232 9132
rect 10284 9160 10290 9172
rect 10410 9160 10416 9172
rect 10284 9132 10416 9160
rect 10284 9120 10290 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11698 9160 11704 9172
rect 11379 9132 11704 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 11940 9132 12173 9160
rect 11940 9120 11946 9132
rect 12161 9129 12173 9132
rect 12207 9160 12219 9163
rect 13906 9160 13912 9172
rect 12207 9132 13912 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 16117 9163 16175 9169
rect 16117 9160 16129 9163
rect 14016 9132 16129 9160
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 9640 9064 11008 9092
rect 9640 9052 9646 9064
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 10042 9024 10048 9036
rect 9723 8996 10048 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10980 9033 11008 9064
rect 11514 9052 11520 9104
rect 11572 9092 11578 9104
rect 13170 9092 13176 9104
rect 11572 9064 13176 9092
rect 11572 9052 11578 9064
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 9024 11207 9027
rect 11606 9024 11612 9036
rect 11195 8996 11612 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 11606 8984 11612 8996
rect 11664 8984 11670 9036
rect 12084 9033 12112 9064
rect 13170 9052 13176 9064
rect 13228 9052 13234 9104
rect 14016 9092 14044 9132
rect 16117 9129 16129 9132
rect 16163 9129 16175 9163
rect 16117 9123 16175 9129
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 18966 9160 18972 9172
rect 16448 9132 18972 9160
rect 16448 9120 16454 9132
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 19702 9120 19708 9172
rect 19760 9160 19766 9172
rect 19760 9132 20392 9160
rect 19760 9120 19766 9132
rect 15473 9095 15531 9101
rect 15473 9092 15485 9095
rect 13832 9064 14044 9092
rect 14476 9064 15485 9092
rect 12069 9027 12127 9033
rect 12069 8993 12081 9027
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 12894 9024 12900 9036
rect 12759 8996 12900 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 6362 8956 6368 8968
rect 6288 8928 6368 8956
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 8478 8956 8484 8968
rect 7432 8928 8484 8956
rect 7432 8916 7438 8928
rect 8478 8916 8484 8928
rect 8536 8956 8542 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8536 8928 8769 8956
rect 8536 8916 8542 8928
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 9232 8956 9260 8984
rect 11974 8956 11980 8968
rect 9232 8928 11980 8956
rect 8757 8919 8815 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12268 8956 12296 8987
rect 12894 8984 12900 8996
rect 12952 9024 12958 9036
rect 13832 9033 13860 9064
rect 13817 9027 13875 9033
rect 12952 8996 13768 9024
rect 12952 8984 12958 8996
rect 12618 8956 12624 8968
rect 12268 8928 12624 8956
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 12986 8916 12992 8968
rect 13044 8956 13050 8968
rect 13630 8956 13636 8968
rect 13044 8928 13636 8956
rect 13044 8916 13050 8928
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13740 8956 13768 8996
rect 13817 8993 13829 9027
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 14001 9027 14059 9033
rect 14001 9024 14013 9027
rect 13964 8996 14013 9024
rect 13964 8984 13970 8996
rect 14001 8993 14013 8996
rect 14047 8993 14059 9027
rect 14001 8987 14059 8993
rect 14274 8984 14280 9036
rect 14332 8984 14338 9036
rect 14476 9033 14504 9064
rect 15473 9061 15485 9064
rect 15519 9061 15531 9095
rect 15473 9055 15531 9061
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 20364 9092 20392 9132
rect 20438 9120 20444 9172
rect 20496 9120 20502 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 20898 9160 20904 9172
rect 20588 9132 20904 9160
rect 20588 9120 20594 9132
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 22830 9160 22836 9172
rect 21560 9132 22836 9160
rect 21560 9092 21588 9132
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 23014 9120 23020 9172
rect 23072 9120 23078 9172
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 25869 9163 25927 9169
rect 23532 9132 25176 9160
rect 23532 9120 23538 9132
rect 21726 9092 21732 9104
rect 17092 9064 20300 9092
rect 20364 9064 21588 9092
rect 21652 9064 21732 9092
rect 17092 9052 17098 9064
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 8993 14519 9027
rect 14461 8987 14519 8993
rect 14560 9002 14964 9030
rect 14560 8956 14588 9002
rect 13740 8928 14588 8956
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8925 14703 8959
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14645 8919 14703 8925
rect 14826 8925 14841 8956
rect 14875 8925 14887 8959
rect 14936 8956 14964 9002
rect 15010 8984 15016 9036
rect 15068 8984 15074 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15120 8996 15669 9024
rect 15120 8956 15148 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 8993 15991 9027
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 15933 8987 15991 8993
rect 16040 8996 16497 9024
rect 14936 8928 15148 8956
rect 14826 8919 14887 8925
rect 7006 8888 7012 8900
rect 5552 8860 7012 8888
rect 7006 8848 7012 8860
rect 7064 8848 7070 8900
rect 7101 8891 7159 8897
rect 7101 8857 7113 8891
rect 7147 8888 7159 8891
rect 9766 8888 9772 8900
rect 7147 8860 9772 8888
rect 7147 8857 7159 8860
rect 7101 8851 7159 8857
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 12434 8888 12440 8900
rect 10192 8860 12440 8888
rect 10192 8848 10198 8860
rect 12434 8848 12440 8860
rect 12492 8888 12498 8900
rect 12897 8891 12955 8897
rect 12897 8888 12909 8891
rect 12492 8860 12909 8888
rect 12492 8848 12498 8860
rect 12897 8857 12909 8860
rect 12943 8857 12955 8891
rect 12897 8851 12955 8857
rect 13722 8848 13728 8900
rect 13780 8888 13786 8900
rect 14660 8888 14688 8919
rect 13780 8860 14688 8888
rect 14826 8888 14854 8919
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15565 8959 15623 8965
rect 15565 8956 15577 8959
rect 15436 8928 15577 8956
rect 15436 8916 15442 8928
rect 15565 8925 15577 8928
rect 15611 8925 15623 8959
rect 15764 8956 15792 8987
rect 15565 8919 15623 8925
rect 15672 8928 15792 8956
rect 14918 8888 14924 8900
rect 14826 8860 14924 8888
rect 13780 8848 13786 8860
rect 14918 8848 14924 8860
rect 14976 8848 14982 8900
rect 15289 8891 15347 8897
rect 15289 8857 15301 8891
rect 15335 8888 15347 8891
rect 15672 8888 15700 8928
rect 15948 8900 15976 8987
rect 15335 8860 15700 8888
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 6270 8820 6276 8832
rect 5184 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 8202 8820 8208 8832
rect 7432 8792 8208 8820
rect 7432 8780 7438 8792
rect 8202 8780 8208 8792
rect 8260 8820 8266 8832
rect 8386 8820 8392 8832
rect 8260 8792 8392 8820
rect 8260 8780 8266 8792
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 8665 8823 8723 8829
rect 8665 8820 8677 8823
rect 8536 8792 8677 8820
rect 8536 8780 8542 8792
rect 8665 8789 8677 8792
rect 8711 8789 8723 8823
rect 8665 8783 8723 8789
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9401 8823 9459 8829
rect 9401 8820 9413 8823
rect 9180 8792 9413 8820
rect 9180 8780 9186 8792
rect 9401 8789 9413 8792
rect 9447 8789 9459 8823
rect 9401 8783 9459 8789
rect 10318 8780 10324 8832
rect 10376 8820 10382 8832
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 10376 8792 11161 8820
rect 10376 8780 10382 8792
rect 11149 8789 11161 8792
rect 11195 8820 11207 8823
rect 12342 8820 12348 8832
rect 11195 8792 12348 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12526 8780 12532 8832
rect 12584 8780 12590 8832
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 15304 8820 15332 8851
rect 15930 8848 15936 8900
rect 15988 8848 15994 8900
rect 13228 8792 15332 8820
rect 13228 8780 13234 8792
rect 15378 8780 15384 8832
rect 15436 8820 15442 8832
rect 16040 8820 16068 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16758 8984 16764 9036
rect 16816 9024 16822 9036
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 16816 8996 17325 9024
rect 16816 8984 16822 8996
rect 17313 8993 17325 8996
rect 17359 9024 17371 9027
rect 17359 8996 17724 9024
rect 17359 8993 17371 8996
rect 17313 8987 17371 8993
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 16776 8956 16804 8984
rect 16439 8928 16804 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8925 17647 8959
rect 17696 8956 17724 8996
rect 17769 8984 17775 9036
rect 17827 9024 17833 9036
rect 18616 9033 18644 9064
rect 18417 9027 18475 9033
rect 17827 8996 17872 9024
rect 17827 8984 17833 8996
rect 18417 8993 18429 9027
rect 18463 8993 18475 9027
rect 18417 8987 18475 8993
rect 18601 9027 18659 9033
rect 18601 8993 18613 9027
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 18046 8956 18052 8968
rect 17696 8928 18052 8956
rect 17589 8919 17647 8925
rect 16758 8848 16764 8900
rect 16816 8888 16822 8900
rect 17405 8891 17463 8897
rect 17405 8888 17417 8891
rect 16816 8860 17417 8888
rect 16816 8848 16822 8860
rect 17405 8857 17417 8860
rect 17451 8857 17463 8891
rect 17405 8851 17463 8857
rect 15436 8792 16068 8820
rect 16485 8823 16543 8829
rect 15436 8780 15442 8792
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 17034 8820 17040 8832
rect 16531 8792 17040 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8820 17187 8823
rect 17218 8820 17224 8832
rect 17175 8792 17224 8820
rect 17175 8789 17187 8792
rect 17129 8783 17187 8789
rect 17218 8780 17224 8792
rect 17276 8780 17282 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17604 8820 17632 8919
rect 18046 8916 18052 8928
rect 18104 8956 18110 8968
rect 18432 8956 18460 8987
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 18969 9027 19027 9033
rect 18969 9024 18981 9027
rect 18840 8996 18981 9024
rect 18840 8984 18846 8996
rect 18969 8993 18981 8996
rect 19015 8993 19027 9027
rect 18969 8987 19027 8993
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 19702 9024 19708 9036
rect 19208 8996 19708 9024
rect 19208 8984 19214 8996
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 19981 9027 20039 9033
rect 19981 8993 19993 9027
rect 20027 9024 20039 9027
rect 20027 8996 20116 9024
rect 20027 8993 20039 8996
rect 19981 8987 20039 8993
rect 18104 8928 18460 8956
rect 18104 8916 18110 8928
rect 17368 8792 17632 8820
rect 17368 8780 17374 8792
rect 17678 8780 17684 8832
rect 17736 8820 17742 8832
rect 17862 8820 17868 8832
rect 17736 8792 17868 8820
rect 17736 8780 17742 8792
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18432 8820 18460 8928
rect 18506 8848 18512 8900
rect 18564 8888 18570 8900
rect 19518 8888 19524 8900
rect 18564 8860 19524 8888
rect 18564 8848 18570 8860
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 19978 8848 19984 8900
rect 20036 8888 20042 8900
rect 20088 8888 20116 8996
rect 20162 8984 20168 9036
rect 20220 8984 20226 9036
rect 20272 9024 20300 9064
rect 20990 9024 20996 9036
rect 20272 8996 20996 9024
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 21100 8996 21281 9024
rect 20441 8959 20499 8965
rect 20441 8925 20453 8959
rect 20487 8956 20499 8959
rect 21100 8956 21128 8996
rect 21269 8993 21281 8996
rect 21315 9024 21327 9027
rect 21315 8996 21496 9024
rect 21315 8993 21327 8996
rect 21269 8987 21327 8993
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 20487 8928 21128 8956
rect 21192 8928 21373 8956
rect 20487 8925 20499 8928
rect 20441 8919 20499 8925
rect 20530 8888 20536 8900
rect 20036 8860 20536 8888
rect 20036 8848 20042 8860
rect 20530 8848 20536 8860
rect 20588 8848 20594 8900
rect 21082 8848 21088 8900
rect 21140 8888 21146 8900
rect 21192 8888 21220 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21468 8956 21496 8996
rect 21542 8984 21548 9036
rect 21600 8984 21606 9036
rect 21652 9033 21680 9064
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 22094 9052 22100 9104
rect 22152 9092 22158 9104
rect 23658 9092 23664 9104
rect 22152 9064 23664 9092
rect 22152 9052 22158 9064
rect 21637 9027 21695 9033
rect 21637 8993 21649 9027
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 21818 8984 21824 9036
rect 21876 8984 21882 9036
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 23014 9024 23020 9036
rect 22060 8996 23020 9024
rect 22060 8984 22066 8996
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 23290 8984 23296 9036
rect 23348 8984 23354 9036
rect 23400 9033 23428 9064
rect 23658 9052 23664 9064
rect 23716 9052 23722 9104
rect 23842 9052 23848 9104
rect 23900 9092 23906 9104
rect 24765 9095 24823 9101
rect 23900 9064 24608 9092
rect 23900 9052 23906 9064
rect 23385 9027 23443 9033
rect 23385 8993 23397 9027
rect 23431 8993 23443 9027
rect 23385 8987 23443 8993
rect 23566 8984 23572 9036
rect 23624 9024 23630 9036
rect 23624 8996 23796 9024
rect 23624 8984 23630 8996
rect 22922 8956 22928 8968
rect 21468 8928 22928 8956
rect 21361 8919 21419 8925
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 23106 8916 23112 8968
rect 23164 8956 23170 8968
rect 23201 8959 23259 8965
rect 23201 8956 23213 8959
rect 23164 8928 23213 8956
rect 23164 8916 23170 8928
rect 23201 8925 23213 8928
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8956 23535 8959
rect 23658 8956 23664 8968
rect 23523 8928 23664 8956
rect 23523 8925 23535 8928
rect 23477 8919 23535 8925
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 23768 8956 23796 8996
rect 24026 8984 24032 9036
rect 24084 8984 24090 9036
rect 24210 8984 24216 9036
rect 24268 8984 24274 9036
rect 24486 8984 24492 9036
rect 24544 8984 24550 9036
rect 24580 9024 24608 9064
rect 24765 9061 24777 9095
rect 24811 9092 24823 9095
rect 25148 9092 25176 9132
rect 25869 9129 25881 9163
rect 25915 9160 25927 9163
rect 25958 9160 25964 9172
rect 25915 9132 25964 9160
rect 25915 9129 25927 9132
rect 25869 9123 25927 9129
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 26050 9120 26056 9172
rect 26108 9160 26114 9172
rect 27522 9160 27528 9172
rect 26108 9132 27528 9160
rect 26108 9120 26114 9132
rect 27522 9120 27528 9132
rect 27580 9120 27586 9172
rect 27617 9163 27675 9169
rect 27617 9129 27629 9163
rect 27663 9160 27675 9163
rect 28258 9160 28264 9172
rect 27663 9132 28264 9160
rect 27663 9129 27675 9132
rect 27617 9123 27675 9129
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 28408 9132 28457 9160
rect 28408 9120 28414 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 28445 9123 28503 9129
rect 29086 9120 29092 9172
rect 29144 9160 29150 9172
rect 29362 9160 29368 9172
rect 29144 9132 29368 9160
rect 29144 9120 29150 9132
rect 29362 9120 29368 9132
rect 29420 9120 29426 9172
rect 29638 9120 29644 9172
rect 29696 9160 29702 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 29696 9132 29837 9160
rect 29696 9120 29702 9132
rect 29825 9129 29837 9132
rect 29871 9129 29883 9163
rect 29825 9123 29883 9129
rect 30282 9120 30288 9172
rect 30340 9120 30346 9172
rect 30300 9092 30328 9120
rect 30653 9095 30711 9101
rect 30653 9092 30665 9095
rect 24811 9064 25084 9092
rect 25148 9064 30665 9092
rect 24811 9061 24823 9064
rect 24765 9055 24823 9061
rect 24857 9027 24915 9033
rect 24857 9024 24869 9027
rect 24580 8996 24869 9024
rect 24857 8993 24869 8996
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 24504 8956 24532 8984
rect 23768 8928 24532 8956
rect 24394 8888 24400 8900
rect 21140 8860 21220 8888
rect 21651 8860 24400 8888
rect 21140 8848 21146 8860
rect 19153 8823 19211 8829
rect 19153 8820 19165 8823
rect 18432 8792 19165 8820
rect 19153 8789 19165 8792
rect 19199 8820 19211 8823
rect 19334 8820 19340 8832
rect 19199 8792 19340 8820
rect 19199 8789 19211 8792
rect 19153 8783 19211 8789
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19794 8780 19800 8832
rect 19852 8780 19858 8832
rect 19886 8780 19892 8832
rect 19944 8820 19950 8832
rect 20254 8820 20260 8832
rect 19944 8792 20260 8820
rect 19944 8780 19950 8792
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 20622 8780 20628 8832
rect 20680 8820 20686 8832
rect 21651 8820 21679 8860
rect 24394 8848 24400 8860
rect 24452 8848 24458 8900
rect 25056 8888 25084 9064
rect 30653 9061 30665 9064
rect 30699 9061 30711 9095
rect 30653 9055 30711 9061
rect 30834 9052 30840 9104
rect 30892 9092 30898 9104
rect 31202 9092 31208 9104
rect 30892 9064 31208 9092
rect 30892 9052 30898 9064
rect 31202 9052 31208 9064
rect 31260 9052 31266 9104
rect 25406 8984 25412 9036
rect 25464 8984 25470 9036
rect 25685 9027 25743 9033
rect 25685 8993 25697 9027
rect 25731 9024 25743 9027
rect 26878 9024 26884 9036
rect 25731 8996 26884 9024
rect 25731 8993 25743 8996
rect 25685 8987 25743 8993
rect 26878 8984 26884 8996
rect 26936 9024 26942 9036
rect 27157 9027 27215 9033
rect 26936 8996 27108 9024
rect 26936 8984 26942 8996
rect 25222 8916 25228 8968
rect 25280 8956 25286 8968
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25280 8928 25513 8956
rect 25280 8916 25286 8928
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 26786 8956 26792 8968
rect 25501 8919 25559 8925
rect 25608 8928 26792 8956
rect 25608 8888 25636 8928
rect 26786 8916 26792 8928
rect 26844 8916 26850 8968
rect 27080 8956 27108 8996
rect 27157 8993 27169 9027
rect 27203 9024 27215 9027
rect 27338 9024 27344 9036
rect 27203 8996 27344 9024
rect 27203 8993 27215 8996
rect 27157 8987 27215 8993
rect 27338 8984 27344 8996
rect 27396 8984 27402 9036
rect 27433 9027 27491 9033
rect 27433 8993 27445 9027
rect 27479 9024 27491 9027
rect 27479 8996 27568 9024
rect 27479 8993 27491 8996
rect 27433 8987 27491 8993
rect 27080 8928 27476 8956
rect 27448 8900 27476 8928
rect 25056 8860 25636 8888
rect 26694 8848 26700 8900
rect 26752 8888 26758 8900
rect 27249 8891 27307 8897
rect 27249 8888 27261 8891
rect 26752 8860 27261 8888
rect 26752 8848 26758 8860
rect 27249 8857 27261 8860
rect 27295 8857 27307 8891
rect 27249 8851 27307 8857
rect 27341 8891 27399 8897
rect 27341 8857 27353 8891
rect 27387 8857 27399 8891
rect 27341 8851 27399 8857
rect 20680 8792 21679 8820
rect 20680 8780 20686 8792
rect 22002 8780 22008 8832
rect 22060 8820 22066 8832
rect 23474 8820 23480 8832
rect 22060 8792 23480 8820
rect 22060 8780 22066 8792
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 25038 8780 25044 8832
rect 25096 8780 25102 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 25958 8780 25964 8832
rect 26016 8820 26022 8832
rect 26418 8820 26424 8832
rect 26016 8792 26424 8820
rect 26016 8780 26022 8792
rect 26418 8780 26424 8792
rect 26476 8780 26482 8832
rect 26510 8780 26516 8832
rect 26568 8820 26574 8832
rect 26881 8823 26939 8829
rect 26881 8820 26893 8823
rect 26568 8792 26893 8820
rect 26568 8780 26574 8792
rect 26881 8789 26893 8792
rect 26927 8820 26939 8823
rect 27356 8820 27384 8851
rect 27430 8848 27436 8900
rect 27488 8848 27494 8900
rect 27540 8832 27568 8996
rect 27614 8984 27620 9036
rect 27672 9024 27678 9036
rect 28077 9027 28135 9033
rect 28077 9024 28089 9027
rect 27672 8996 28089 9024
rect 27672 8984 27678 8996
rect 28077 8993 28089 8996
rect 28123 8993 28135 9027
rect 28077 8987 28135 8993
rect 28261 9027 28319 9033
rect 28261 8993 28273 9027
rect 28307 9024 28319 9027
rect 28350 9024 28356 9036
rect 28307 8996 28356 9024
rect 28307 8993 28319 8996
rect 28261 8987 28319 8993
rect 28350 8984 28356 8996
rect 28408 8984 28414 9036
rect 28902 9024 28908 9036
rect 28552 8996 28908 9024
rect 27706 8916 27712 8968
rect 27764 8956 27770 8968
rect 28552 8956 28580 8996
rect 28902 8984 28908 8996
rect 28960 8984 28966 9036
rect 29089 9027 29147 9033
rect 29089 8993 29101 9027
rect 29135 8993 29147 9027
rect 29089 8987 29147 8993
rect 29365 9027 29423 9033
rect 29365 8993 29377 9027
rect 29411 9024 29423 9027
rect 29454 9024 29460 9036
rect 29411 8996 29460 9024
rect 29411 8993 29423 8996
rect 29365 8987 29423 8993
rect 29104 8956 29132 8987
rect 29454 8984 29460 8996
rect 29512 9024 29518 9036
rect 29914 9024 29920 9036
rect 29512 8996 29920 9024
rect 29512 8984 29518 8996
rect 29914 8984 29920 8996
rect 29972 8984 29978 9036
rect 30098 8984 30104 9036
rect 30156 8984 30162 9036
rect 30190 8984 30196 9036
rect 30248 8984 30254 9036
rect 30285 9027 30343 9033
rect 30285 8993 30297 9027
rect 30331 9024 30343 9027
rect 30469 9027 30527 9033
rect 30331 8996 30420 9024
rect 30331 8993 30343 8996
rect 30285 8987 30343 8993
rect 30392 8968 30420 8996
rect 30469 8993 30481 9027
rect 30515 9024 30527 9027
rect 30558 9024 30564 9036
rect 30515 8996 30564 9024
rect 30515 8993 30527 8996
rect 30469 8987 30527 8993
rect 30558 8984 30564 8996
rect 30616 8984 30622 9036
rect 30926 8984 30932 9036
rect 30984 9024 30990 9036
rect 31478 9024 31484 9036
rect 30984 8996 31484 9024
rect 30984 8984 30990 8996
rect 31478 8984 31484 8996
rect 31536 8984 31542 9036
rect 27764 8928 28580 8956
rect 28644 8928 30144 8956
rect 27764 8916 27770 8928
rect 26927 8792 27384 8820
rect 26927 8789 26939 8792
rect 26881 8783 26939 8789
rect 27522 8780 27528 8832
rect 27580 8780 27586 8832
rect 28074 8780 28080 8832
rect 28132 8820 28138 8832
rect 28644 8829 28672 8928
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 29362 8888 29368 8900
rect 29052 8860 29368 8888
rect 29052 8848 29058 8860
rect 29362 8848 29368 8860
rect 29420 8848 29426 8900
rect 30116 8888 30144 8928
rect 30374 8916 30380 8968
rect 30432 8916 30438 8968
rect 30190 8888 30196 8900
rect 30116 8860 30196 8888
rect 30190 8848 30196 8860
rect 30248 8848 30254 8900
rect 30466 8848 30472 8900
rect 30524 8888 30530 8900
rect 30837 8891 30895 8897
rect 30837 8888 30849 8891
rect 30524 8860 30849 8888
rect 30524 8848 30530 8860
rect 30837 8857 30849 8860
rect 30883 8888 30895 8891
rect 31294 8888 31300 8900
rect 30883 8860 31300 8888
rect 30883 8857 30895 8860
rect 30837 8851 30895 8857
rect 31294 8848 31300 8860
rect 31352 8848 31358 8900
rect 28629 8823 28687 8829
rect 28629 8820 28641 8823
rect 28132 8792 28641 8820
rect 28132 8780 28138 8792
rect 28629 8789 28641 8792
rect 28675 8789 28687 8823
rect 28629 8783 28687 8789
rect 552 8730 31648 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 11436 8730
rect 11488 8678 11500 8730
rect 11552 8678 11564 8730
rect 11616 8678 11628 8730
rect 11680 8678 11692 8730
rect 11744 8678 19210 8730
rect 19262 8678 19274 8730
rect 19326 8678 19338 8730
rect 19390 8678 19402 8730
rect 19454 8678 19466 8730
rect 19518 8678 26984 8730
rect 27036 8678 27048 8730
rect 27100 8678 27112 8730
rect 27164 8678 27176 8730
rect 27228 8678 27240 8730
rect 27292 8678 31648 8730
rect 552 8656 31648 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2041 8619 2099 8625
rect 2041 8616 2053 8619
rect 1811 8588 2053 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2041 8585 2053 8588
rect 2087 8616 2099 8619
rect 3050 8616 3056 8628
rect 2087 8588 3056 8616
rect 2087 8585 2099 8588
rect 2041 8579 2099 8585
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3970 8576 3976 8628
rect 4028 8616 4034 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4028 8588 4261 8616
rect 4028 8576 4034 8588
rect 4249 8585 4261 8588
rect 4295 8616 4307 8619
rect 4338 8616 4344 8628
rect 4295 8588 4344 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5074 8616 5080 8628
rect 4856 8588 5080 8616
rect 4856 8576 4862 8588
rect 5074 8576 5080 8588
rect 5132 8616 5138 8628
rect 5258 8616 5264 8628
rect 5132 8588 5264 8616
rect 5132 8576 5138 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 6454 8576 6460 8628
rect 6512 8576 6518 8628
rect 7466 8576 7472 8628
rect 7524 8576 7530 8628
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 9398 8616 9404 8628
rect 8352 8588 9404 8616
rect 8352 8576 8358 8588
rect 9398 8576 9404 8588
rect 9456 8616 9462 8628
rect 10686 8616 10692 8628
rect 9456 8588 10692 8616
rect 9456 8576 9462 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11514 8616 11520 8628
rect 11204 8588 11520 8616
rect 11204 8576 11210 8588
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11848 8588 12081 8616
rect 11848 8576 11854 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 12250 8576 12256 8628
rect 12308 8616 12314 8628
rect 12802 8616 12808 8628
rect 12308 8588 12808 8616
rect 12308 8576 12314 8588
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 14182 8616 14188 8628
rect 13219 8588 14188 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 1581 8551 1639 8557
rect 1581 8517 1593 8551
rect 1627 8548 1639 8551
rect 1670 8548 1676 8560
rect 1627 8520 1676 8548
rect 1627 8517 1639 8520
rect 1581 8511 1639 8517
rect 1670 8508 1676 8520
rect 1728 8508 1734 8560
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8517 2283 8551
rect 2225 8511 2283 8517
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 1673 8415 1731 8421
rect 1673 8412 1685 8415
rect 1636 8384 1685 8412
rect 1636 8372 1642 8384
rect 1673 8381 1685 8384
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8381 1915 8415
rect 1857 8375 1915 8381
rect 1305 8347 1363 8353
rect 1305 8313 1317 8347
rect 1351 8344 1363 8347
rect 1486 8344 1492 8356
rect 1351 8316 1492 8344
rect 1351 8313 1363 8316
rect 1305 8307 1363 8313
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 1872 8344 1900 8375
rect 2038 8372 2044 8424
rect 2096 8372 2102 8424
rect 2240 8412 2268 8511
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 5537 8551 5595 8557
rect 5537 8548 5549 8551
rect 2464 8520 5549 8548
rect 2464 8508 2470 8520
rect 5537 8517 5549 8520
rect 5583 8517 5595 8551
rect 5537 8511 5595 8517
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 6730 8548 6736 8560
rect 5868 8520 6736 8548
rect 5868 8508 5874 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 6825 8551 6883 8557
rect 6825 8517 6837 8551
rect 6871 8517 6883 8551
rect 6825 8511 6883 8517
rect 7193 8551 7251 8557
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 7374 8548 7380 8560
rect 7239 8520 7380 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 5353 8483 5411 8489
rect 4212 8452 5028 8480
rect 4212 8440 4218 8452
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2240 8384 3249 8412
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 3384 8384 3433 8412
rect 3384 8372 3390 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 3510 8372 3516 8424
rect 3568 8372 3574 8424
rect 3602 8372 3608 8424
rect 3660 8372 3666 8424
rect 3694 8372 3700 8424
rect 3752 8372 3758 8424
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4304 8384 4353 8412
rect 4304 8372 4310 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 4672 8384 4721 8412
rect 4672 8372 4678 8384
rect 4709 8381 4721 8384
rect 4755 8381 4767 8415
rect 4709 8375 4767 8381
rect 4890 8372 4896 8424
rect 4948 8372 4954 8424
rect 5000 8421 5028 8452
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 6086 8480 6092 8492
rect 5399 8452 6092 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 6454 8412 6460 8424
rect 5276 8384 6460 8412
rect 2222 8344 2228 8356
rect 1872 8316 2228 8344
rect 2222 8304 2228 8316
rect 2280 8304 2286 8356
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 2924 8316 3893 8344
rect 2924 8304 2930 8316
rect 3881 8313 3893 8316
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8344 4583 8347
rect 5166 8344 5172 8356
rect 4571 8316 5172 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 1394 8236 1400 8288
rect 1452 8276 1458 8288
rect 2406 8276 2412 8288
rect 1452 8248 2412 8276
rect 1452 8236 1458 8248
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3234 8276 3240 8288
rect 3016 8248 3240 8276
rect 3016 8236 3022 8248
rect 3234 8236 3240 8248
rect 3292 8276 3298 8288
rect 3694 8276 3700 8288
rect 3292 8248 3700 8276
rect 3292 8236 3298 8248
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 5276 8276 5304 8384
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 6546 8372 6552 8424
rect 6604 8412 6610 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6604 8384 6653 8412
rect 6604 8372 6610 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6840 8412 6868 8511
rect 7374 8508 7380 8520
rect 7432 8508 7438 8560
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7147 8452 7573 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7852 8480 7880 8576
rect 8389 8551 8447 8557
rect 8389 8517 8401 8551
rect 8435 8548 8447 8551
rect 13722 8548 13728 8560
rect 8435 8520 11376 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 7561 8443 7619 8449
rect 7760 8452 8156 8480
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6840 8384 7021 8412
rect 6641 8375 6699 8381
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7650 8412 7656 8424
rect 7331 8384 7656 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5684 8316 5917 8344
rect 5684 8304 5690 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 6656 8344 6684 8375
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 7760 8421 7788 8452
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8381 7803 8415
rect 7745 8375 7803 8381
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7892 8384 8033 8412
rect 7892 8372 7898 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8128 8412 8156 8452
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8665 8483 8723 8489
rect 8665 8480 8677 8483
rect 8260 8452 8677 8480
rect 8260 8440 8266 8452
rect 8665 8449 8677 8452
rect 8711 8449 8723 8483
rect 8665 8443 8723 8449
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 10686 8480 10692 8492
rect 8864 8452 10692 8480
rect 8864 8424 8892 8452
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11348 8489 11376 8520
rect 11532 8520 13728 8548
rect 11532 8489 11560 8520
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 11020 8452 11161 8480
rect 11020 8440 11026 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 13832 8480 13860 8588
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14553 8619 14611 8625
rect 14553 8616 14565 8619
rect 14415 8588 14565 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14553 8585 14565 8588
rect 14599 8585 14611 8619
rect 14553 8579 14611 8585
rect 14936 8588 15243 8616
rect 14936 8548 14964 8588
rect 12728 8452 13860 8480
rect 14016 8520 14964 8548
rect 8294 8412 8300 8424
rect 8128 8384 8300 8412
rect 8021 8375 8079 8381
rect 8294 8372 8300 8384
rect 8352 8412 8358 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8352 8384 8585 8412
rect 8352 8372 8358 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8846 8372 8852 8424
rect 8904 8372 8910 8424
rect 9030 8372 9036 8424
rect 9088 8372 9094 8424
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 10008 8384 10333 8412
rect 10008 8372 10014 8384
rect 10321 8381 10333 8384
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 10560 8384 10640 8412
rect 10560 8372 10566 8384
rect 10612 8344 10640 8384
rect 11422 8372 11428 8424
rect 11480 8372 11486 8424
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8412 11667 8415
rect 11790 8412 11796 8424
rect 11655 8384 11796 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12250 8372 12256 8424
rect 12308 8372 12314 8424
rect 12342 8372 12348 8424
rect 12400 8372 12406 8424
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 11974 8344 11980 8356
rect 6656 8316 10548 8344
rect 10612 8316 11980 8344
rect 5905 8307 5963 8313
rect 4488 8248 5304 8276
rect 4488 8236 4494 8248
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8662 8276 8668 8288
rect 7984 8248 8668 8276
rect 7984 8236 7990 8248
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 9858 8276 9864 8288
rect 8904 8248 9864 8276
rect 8904 8236 8910 8248
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10410 8236 10416 8288
rect 10468 8236 10474 8288
rect 10520 8276 10548 8316
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12452 8344 12480 8375
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12728 8421 12756 8452
rect 12713 8415 12771 8421
rect 12713 8412 12725 8415
rect 12676 8384 12725 8412
rect 12676 8372 12682 8384
rect 12713 8381 12725 8384
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12802 8372 12808 8424
rect 12860 8372 12866 8424
rect 12989 8415 13047 8421
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13170 8412 13176 8424
rect 13035 8384 13176 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 13906 8372 13912 8424
rect 13964 8372 13970 8424
rect 14016 8421 14044 8520
rect 15010 8508 15016 8560
rect 15068 8508 15074 8560
rect 15215 8548 15243 8588
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 18230 8616 18236 8628
rect 15436 8588 18236 8616
rect 15436 8576 15442 8588
rect 18230 8576 18236 8588
rect 18288 8616 18294 8628
rect 18966 8616 18972 8628
rect 18288 8588 18972 8616
rect 18288 8576 18294 8588
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 20346 8616 20352 8628
rect 19484 8588 20352 8616
rect 19484 8576 19490 8588
rect 20346 8576 20352 8588
rect 20404 8576 20410 8628
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 21634 8616 21640 8628
rect 20864 8588 21640 8616
rect 20864 8576 20870 8588
rect 21634 8576 21640 8588
rect 21692 8616 21698 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21692 8588 22017 8616
rect 21692 8576 21698 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 22370 8576 22376 8628
rect 22428 8576 22434 8628
rect 23106 8576 23112 8628
rect 23164 8576 23170 8628
rect 24397 8619 24455 8625
rect 24397 8585 24409 8619
rect 24443 8616 24455 8619
rect 24578 8616 24584 8628
rect 24443 8588 24584 8616
rect 24443 8585 24455 8588
rect 24397 8579 24455 8585
rect 24578 8576 24584 8588
rect 24636 8576 24642 8628
rect 25590 8576 25596 8628
rect 25648 8576 25654 8628
rect 25774 8576 25780 8628
rect 25832 8616 25838 8628
rect 25832 8588 26280 8616
rect 25832 8576 25838 8588
rect 19061 8551 19119 8557
rect 19061 8548 19073 8551
rect 15215 8520 19073 8548
rect 19061 8517 19073 8520
rect 19107 8517 19119 8551
rect 19061 8511 19119 8517
rect 19242 8508 19248 8560
rect 19300 8548 19306 8560
rect 19978 8548 19984 8560
rect 19300 8520 19984 8548
rect 19300 8508 19306 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 20165 8551 20223 8557
rect 20165 8517 20177 8551
rect 20211 8548 20223 8551
rect 20211 8520 21496 8548
rect 20211 8517 20223 8520
rect 20165 8511 20223 8517
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 16758 8480 16764 8492
rect 14240 8452 16764 8480
rect 14240 8440 14246 8452
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17310 8440 17316 8492
rect 17368 8440 17374 8492
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17586 8480 17592 8492
rect 17451 8452 17592 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 13354 8344 13360 8356
rect 12452 8316 13360 8344
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 14108 8344 14136 8375
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 14700 8384 14749 8412
rect 14700 8372 14706 8384
rect 14737 8381 14749 8384
rect 14783 8381 14795 8415
rect 15289 8415 15347 8421
rect 15289 8412 15301 8415
rect 14737 8375 14795 8381
rect 14826 8384 15301 8412
rect 13504 8316 14136 8344
rect 13504 8304 13510 8316
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 14826 8344 14854 8384
rect 15289 8381 15301 8384
rect 15335 8381 15347 8415
rect 15289 8375 15347 8381
rect 16298 8372 16304 8424
rect 16356 8412 16362 8424
rect 17420 8412 17448 8443
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 18690 8480 18696 8492
rect 17727 8452 18696 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 21468 8480 21496 8520
rect 21542 8508 21548 8560
rect 21600 8508 21606 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 22738 8548 22744 8560
rect 21784 8520 22744 8548
rect 21784 8508 21790 8520
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 23014 8508 23020 8560
rect 23072 8548 23078 8560
rect 24596 8548 24624 8576
rect 25225 8551 25283 8557
rect 23072 8520 23428 8548
rect 24596 8520 25176 8548
rect 23072 8508 23078 8520
rect 18800 8452 21036 8480
rect 21468 8452 22784 8480
rect 16356 8384 17448 8412
rect 17497 8415 17555 8421
rect 16356 8372 16362 8384
rect 17497 8381 17509 8415
rect 17543 8412 17555 8415
rect 17543 8384 17816 8412
rect 17543 8381 17555 8384
rect 17497 8375 17555 8381
rect 14608 8316 14854 8344
rect 14608 8304 14614 8316
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 15105 8347 15163 8353
rect 15105 8344 15117 8347
rect 15068 8316 15117 8344
rect 15068 8304 15074 8316
rect 15105 8313 15117 8316
rect 15151 8313 15163 8347
rect 15105 8307 15163 8313
rect 15654 8304 15660 8356
rect 15712 8344 15718 8356
rect 16482 8344 16488 8356
rect 15712 8316 16488 8344
rect 15712 8304 15718 8316
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 16758 8304 16764 8356
rect 16816 8344 16822 8356
rect 16816 8316 17172 8344
rect 16816 8304 16822 8316
rect 11330 8276 11336 8288
rect 10520 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11514 8236 11520 8288
rect 11572 8276 11578 8288
rect 13722 8276 13728 8288
rect 11572 8248 13728 8276
rect 11572 8236 11578 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 14734 8276 14740 8288
rect 13872 8248 14740 8276
rect 13872 8236 13878 8248
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 14918 8236 14924 8288
rect 14976 8276 14982 8288
rect 16298 8276 16304 8288
rect 14976 8248 16304 8276
rect 14976 8236 14982 8248
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 17034 8236 17040 8288
rect 17092 8236 17098 8288
rect 17144 8276 17172 8316
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 17681 8347 17739 8353
rect 17681 8344 17693 8347
rect 17368 8316 17693 8344
rect 17368 8304 17374 8316
rect 17681 8313 17693 8316
rect 17727 8313 17739 8347
rect 17681 8307 17739 8313
rect 17788 8276 17816 8384
rect 17862 8372 17868 8424
rect 17920 8372 17926 8424
rect 17957 8415 18015 8421
rect 17957 8381 17969 8415
rect 18003 8412 18015 8415
rect 18046 8412 18052 8424
rect 18003 8384 18052 8412
rect 18003 8381 18015 8384
rect 17957 8375 18015 8381
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18230 8372 18236 8424
rect 18288 8412 18294 8424
rect 18800 8412 18828 8452
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 18288 8384 18828 8412
rect 19878 8409 19901 8412
rect 18288 8372 18294 8384
rect 19812 8381 19901 8409
rect 19935 8381 19947 8415
rect 18690 8304 18696 8356
rect 18748 8304 18754 8356
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 18877 8347 18935 8353
rect 18877 8344 18889 8347
rect 18840 8316 18889 8344
rect 18840 8304 18846 8316
rect 18877 8313 18889 8316
rect 18923 8313 18935 8347
rect 18877 8307 18935 8313
rect 18966 8304 18972 8356
rect 19024 8344 19030 8356
rect 19812 8344 19840 8381
rect 19889 8375 19947 8381
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 20714 8412 20720 8424
rect 20579 8384 20720 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 20806 8372 20812 8424
rect 20864 8372 20870 8424
rect 20901 8418 20959 8421
rect 20898 8366 20904 8418
rect 20956 8366 20962 8418
rect 21008 8412 21036 8452
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 21008 8384 21189 8412
rect 21177 8381 21189 8384
rect 21223 8381 21235 8415
rect 21177 8375 21235 8381
rect 21266 8372 21272 8424
rect 21324 8412 21330 8424
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 21324 8384 21465 8412
rect 21324 8372 21330 8384
rect 21453 8381 21465 8384
rect 21499 8412 21511 8415
rect 21726 8412 21732 8424
rect 21499 8384 21732 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 21818 8372 21824 8424
rect 21876 8372 21882 8424
rect 21913 8415 21971 8421
rect 21913 8381 21925 8415
rect 21959 8412 21971 8415
rect 22002 8412 22008 8424
rect 21959 8384 22008 8412
rect 21959 8381 21971 8384
rect 21913 8375 21971 8381
rect 20070 8344 20076 8356
rect 19024 8316 19840 8344
rect 19904 8316 20076 8344
rect 19024 8304 19030 8316
rect 17954 8276 17960 8288
rect 17144 8248 17960 8276
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 19150 8276 19156 8288
rect 18564 8248 19156 8276
rect 18564 8236 18570 8248
rect 19150 8236 19156 8248
rect 19208 8276 19214 8288
rect 19904 8276 19932 8316
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 20165 8347 20223 8353
rect 20165 8313 20177 8347
rect 20211 8344 20223 8347
rect 20346 8344 20352 8356
rect 20211 8316 20352 8344
rect 20211 8313 20223 8316
rect 20165 8307 20223 8313
rect 20346 8304 20352 8316
rect 20404 8304 20410 8356
rect 21361 8347 21419 8353
rect 21361 8313 21373 8347
rect 21407 8344 21419 8347
rect 21634 8344 21640 8356
rect 21407 8316 21640 8344
rect 21407 8313 21419 8316
rect 21361 8307 21419 8313
rect 21634 8304 21640 8316
rect 21692 8304 21698 8356
rect 19208 8248 19932 8276
rect 19981 8279 20039 8285
rect 19208 8236 19214 8248
rect 19981 8245 19993 8279
rect 20027 8276 20039 8279
rect 20714 8276 20720 8288
rect 20027 8248 20720 8276
rect 20027 8245 20039 8248
rect 19981 8239 20039 8245
rect 20714 8236 20720 8248
rect 20772 8276 20778 8288
rect 21928 8276 21956 8375
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 22097 8415 22155 8421
rect 22097 8381 22109 8415
rect 22143 8381 22155 8415
rect 22097 8375 22155 8381
rect 22281 8415 22339 8421
rect 22281 8381 22293 8415
rect 22327 8412 22339 8415
rect 22370 8412 22376 8424
rect 22327 8384 22376 8412
rect 22327 8381 22339 8384
rect 22281 8375 22339 8381
rect 22112 8344 22140 8375
rect 22370 8372 22376 8384
rect 22428 8372 22434 8424
rect 22646 8372 22652 8424
rect 22704 8372 22710 8424
rect 22756 8421 22784 8452
rect 22940 8452 23152 8480
rect 22741 8415 22799 8421
rect 22741 8381 22753 8415
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 22830 8372 22836 8424
rect 22888 8372 22894 8424
rect 22940 8344 22968 8452
rect 23017 8415 23075 8421
rect 23017 8381 23029 8415
rect 23063 8381 23075 8415
rect 23124 8412 23152 8452
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 23400 8489 23428 8520
rect 23385 8483 23443 8489
rect 23385 8449 23397 8483
rect 23431 8449 23443 8483
rect 25148 8480 25176 8520
rect 25225 8517 25237 8551
rect 25271 8548 25283 8551
rect 26053 8551 26111 8557
rect 26053 8548 26065 8551
rect 25271 8520 26065 8548
rect 25271 8517 25283 8520
rect 25225 8511 25283 8517
rect 26053 8517 26065 8520
rect 26099 8517 26111 8551
rect 26252 8548 26280 8588
rect 26326 8576 26332 8628
rect 26384 8616 26390 8628
rect 26384 8588 27292 8616
rect 26384 8576 26390 8588
rect 26053 8511 26111 8517
rect 26142 8520 26372 8548
rect 23385 8443 23443 8449
rect 24228 8452 24624 8480
rect 25148 8452 25452 8480
rect 23474 8412 23480 8424
rect 23124 8384 23480 8412
rect 23017 8375 23075 8381
rect 22112 8316 22968 8344
rect 20772 8248 21956 8276
rect 20772 8236 20778 8248
rect 22002 8236 22008 8288
rect 22060 8276 22066 8288
rect 22278 8276 22284 8288
rect 22060 8248 22284 8276
rect 22060 8236 22066 8248
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 23032 8276 23060 8375
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 24228 8421 24256 8452
rect 24596 8424 24624 8452
rect 23569 8415 23627 8421
rect 23569 8381 23581 8415
rect 23615 8412 23627 8415
rect 23937 8415 23995 8421
rect 23937 8412 23949 8415
rect 23615 8384 23949 8412
rect 23615 8381 23627 8384
rect 23569 8375 23627 8381
rect 23937 8381 23949 8384
rect 23983 8381 23995 8415
rect 23937 8375 23995 8381
rect 24213 8415 24271 8421
rect 24213 8381 24225 8415
rect 24259 8381 24271 8415
rect 24213 8375 24271 8381
rect 23106 8304 23112 8356
rect 23164 8344 23170 8356
rect 23584 8344 23612 8375
rect 24394 8372 24400 8424
rect 24452 8372 24458 8424
rect 24578 8372 24584 8424
rect 24636 8412 24642 8424
rect 24762 8412 24768 8424
rect 24636 8384 24768 8412
rect 24636 8372 24642 8384
rect 24762 8372 24768 8384
rect 24820 8372 24826 8424
rect 25130 8372 25136 8424
rect 25188 8412 25194 8424
rect 25424 8421 25452 8452
rect 25590 8440 25596 8492
rect 25648 8480 25654 8492
rect 26142 8480 26170 8520
rect 25648 8452 26170 8480
rect 25648 8440 25654 8452
rect 26234 8440 26240 8492
rect 26292 8440 26298 8492
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 25188 8384 25237 8412
rect 25188 8372 25194 8384
rect 25225 8381 25237 8384
rect 25271 8381 25283 8415
rect 25225 8375 25283 8381
rect 25409 8415 25467 8421
rect 25409 8381 25421 8415
rect 25455 8381 25467 8415
rect 25409 8375 25467 8381
rect 25501 8415 25559 8421
rect 25501 8381 25513 8415
rect 25547 8381 25559 8415
rect 25501 8375 25559 8381
rect 23164 8316 23612 8344
rect 23164 8304 23170 8316
rect 23842 8304 23848 8356
rect 23900 8304 23906 8356
rect 25148 8344 25176 8372
rect 23952 8316 25176 8344
rect 25516 8344 25544 8375
rect 25774 8372 25780 8424
rect 25832 8372 25838 8424
rect 25869 8415 25927 8421
rect 25869 8381 25881 8415
rect 25915 8412 25927 8415
rect 25958 8412 25964 8424
rect 25915 8384 25964 8412
rect 25915 8381 25927 8384
rect 25869 8375 25927 8381
rect 25958 8372 25964 8384
rect 26016 8372 26022 8424
rect 26142 8372 26148 8424
rect 26200 8372 26206 8424
rect 26344 8412 26372 8520
rect 26418 8508 26424 8560
rect 26476 8508 26482 8560
rect 27264 8548 27292 8588
rect 27338 8576 27344 8628
rect 27396 8616 27402 8628
rect 27890 8616 27896 8628
rect 27396 8588 27896 8616
rect 27396 8576 27402 8588
rect 27890 8576 27896 8588
rect 27948 8576 27954 8628
rect 29917 8619 29975 8625
rect 29917 8585 29929 8619
rect 29963 8616 29975 8619
rect 30098 8616 30104 8628
rect 29963 8588 30104 8616
rect 29963 8585 29975 8588
rect 29917 8579 29975 8585
rect 27522 8548 27528 8560
rect 27264 8520 27528 8548
rect 27522 8508 27528 8520
rect 27580 8508 27586 8560
rect 28445 8551 28503 8557
rect 28445 8517 28457 8551
rect 28491 8548 28503 8551
rect 29273 8551 29331 8557
rect 29273 8548 29285 8551
rect 28491 8520 29285 8548
rect 28491 8517 28503 8520
rect 28445 8511 28503 8517
rect 29273 8517 29285 8520
rect 29319 8548 29331 8551
rect 29932 8548 29960 8579
rect 30098 8576 30104 8588
rect 30156 8576 30162 8628
rect 30558 8576 30564 8628
rect 30616 8616 30622 8628
rect 30653 8619 30711 8625
rect 30653 8616 30665 8619
rect 30616 8588 30665 8616
rect 30616 8576 30622 8588
rect 30653 8585 30665 8588
rect 30699 8585 30711 8619
rect 30653 8579 30711 8585
rect 29319 8520 29960 8548
rect 29319 8517 29331 8520
rect 29273 8511 29331 8517
rect 27982 8440 27988 8492
rect 28040 8480 28046 8492
rect 28040 8452 29132 8480
rect 28040 8440 28046 8452
rect 26513 8415 26571 8421
rect 26513 8412 26525 8415
rect 26344 8384 26525 8412
rect 26513 8381 26525 8384
rect 26559 8381 26571 8415
rect 27522 8412 27528 8424
rect 26513 8375 26571 8381
rect 26620 8384 27528 8412
rect 26237 8347 26295 8353
rect 26237 8344 26249 8347
rect 25516 8316 26249 8344
rect 23952 8276 23980 8316
rect 26237 8313 26249 8316
rect 26283 8313 26295 8347
rect 26237 8307 26295 8313
rect 23032 8248 23980 8276
rect 24762 8236 24768 8288
rect 24820 8276 24826 8288
rect 25038 8276 25044 8288
rect 24820 8248 25044 8276
rect 24820 8236 24826 8248
rect 25038 8236 25044 8248
rect 25096 8236 25102 8288
rect 25498 8236 25504 8288
rect 25556 8276 25562 8288
rect 26620 8276 26648 8384
rect 27522 8372 27528 8384
rect 27580 8412 27586 8424
rect 28368 8421 28396 8452
rect 28169 8415 28227 8421
rect 28169 8412 28181 8415
rect 27580 8384 28181 8412
rect 27580 8372 27586 8384
rect 28169 8381 28181 8384
rect 28215 8381 28227 8415
rect 28169 8375 28227 8381
rect 28353 8415 28411 8421
rect 28353 8381 28365 8415
rect 28399 8381 28411 8415
rect 28353 8375 28411 8381
rect 28537 8415 28595 8421
rect 28537 8381 28549 8415
rect 28583 8381 28595 8415
rect 28537 8375 28595 8381
rect 28629 8415 28687 8421
rect 28629 8381 28641 8415
rect 28675 8412 28687 8415
rect 29104 8412 29132 8452
rect 29362 8440 29368 8492
rect 29420 8440 29426 8492
rect 29914 8440 29920 8492
rect 29972 8480 29978 8492
rect 29972 8452 30144 8480
rect 29972 8440 29978 8452
rect 30116 8424 30144 8452
rect 29181 8415 29239 8421
rect 29181 8412 29193 8415
rect 28675 8384 28856 8412
rect 29104 8384 29193 8412
rect 28675 8381 28687 8384
rect 28629 8375 28687 8381
rect 27062 8304 27068 8356
rect 27120 8304 27126 8356
rect 27246 8353 27252 8356
rect 27241 8307 27252 8353
rect 27304 8344 27310 8356
rect 27304 8316 27341 8344
rect 27246 8304 27252 8307
rect 27304 8304 27310 8316
rect 27430 8304 27436 8356
rect 27488 8304 27494 8356
rect 27709 8347 27767 8353
rect 27709 8313 27721 8347
rect 27755 8344 27767 8347
rect 28258 8344 28264 8356
rect 27755 8316 28264 8344
rect 27755 8313 27767 8316
rect 27709 8307 27767 8313
rect 28258 8304 28264 8316
rect 28316 8304 28322 8356
rect 28552 8344 28580 8375
rect 28828 8344 28856 8384
rect 29181 8381 29193 8384
rect 29227 8412 29239 8415
rect 29270 8412 29276 8424
rect 29227 8384 29276 8412
rect 29227 8381 29239 8384
rect 29181 8375 29239 8381
rect 29270 8372 29276 8384
rect 29328 8372 29334 8424
rect 29457 8415 29515 8421
rect 29457 8381 29469 8415
rect 29503 8412 29515 8415
rect 30006 8412 30012 8424
rect 29503 8384 30012 8412
rect 29503 8381 29515 8384
rect 29457 8375 29515 8381
rect 30006 8372 30012 8384
rect 30064 8372 30070 8424
rect 30098 8372 30104 8424
rect 30156 8372 30162 8424
rect 30282 8372 30288 8424
rect 30340 8372 30346 8424
rect 30834 8372 30840 8424
rect 30892 8372 30898 8424
rect 30300 8344 30328 8372
rect 31662 8344 31668 8356
rect 28552 8316 28764 8344
rect 28828 8316 29316 8344
rect 30300 8316 31668 8344
rect 25556 8248 26648 8276
rect 25556 8236 25562 8248
rect 26786 8236 26792 8288
rect 26844 8276 26850 8288
rect 27264 8276 27292 8304
rect 26844 8248 27292 8276
rect 26844 8236 26850 8248
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 28626 8276 28632 8288
rect 27856 8248 28632 8276
rect 27856 8236 27862 8248
rect 28626 8236 28632 8248
rect 28684 8236 28690 8288
rect 28736 8276 28764 8316
rect 28902 8276 28908 8288
rect 28736 8248 28908 8276
rect 28902 8236 28908 8248
rect 28960 8236 28966 8288
rect 28994 8236 29000 8288
rect 29052 8236 29058 8288
rect 29288 8276 29316 8316
rect 31662 8304 31668 8316
rect 31720 8304 31726 8356
rect 29546 8276 29552 8288
rect 29288 8248 29552 8276
rect 29546 8236 29552 8248
rect 29604 8236 29610 8288
rect 552 8186 31648 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 12096 8186
rect 12148 8134 12160 8186
rect 12212 8134 12224 8186
rect 12276 8134 12288 8186
rect 12340 8134 12352 8186
rect 12404 8134 19870 8186
rect 19922 8134 19934 8186
rect 19986 8134 19998 8186
rect 20050 8134 20062 8186
rect 20114 8134 20126 8186
rect 20178 8134 27644 8186
rect 27696 8134 27708 8186
rect 27760 8134 27772 8186
rect 27824 8134 27836 8186
rect 27888 8134 27900 8186
rect 27952 8134 31648 8186
rect 552 8112 31648 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 9398 8072 9404 8084
rect 1912 8044 9404 8072
rect 1912 8032 1918 8044
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 11422 8032 11428 8084
rect 11480 8032 11486 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 11563 8044 12756 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 1302 7964 1308 8016
rect 1360 8004 1366 8016
rect 1581 8007 1639 8013
rect 1581 8004 1593 8007
rect 1360 7976 1593 8004
rect 1360 7964 1366 7976
rect 1581 7973 1593 7976
rect 1627 7973 1639 8007
rect 1581 7967 1639 7973
rect 1946 7964 1952 8016
rect 2004 7964 2010 8016
rect 4338 7964 4344 8016
rect 4396 8004 4402 8016
rect 5350 8004 5356 8016
rect 4396 7976 5356 8004
rect 4396 7964 4402 7976
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 8754 8004 8760 8016
rect 7432 7976 8760 8004
rect 7432 7964 7438 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 8849 8007 8907 8013
rect 8849 7973 8861 8007
rect 8895 7973 8907 8007
rect 8849 7967 8907 7973
rect 8941 8007 8999 8013
rect 8941 7973 8953 8007
rect 8987 8004 8999 8007
rect 9030 8004 9036 8016
rect 8987 7976 9036 8004
rect 8987 7973 8999 7976
rect 8941 7967 8999 7973
rect 1213 7939 1271 7945
rect 1213 7905 1225 7939
rect 1259 7936 1271 7939
rect 1397 7939 1455 7945
rect 1259 7908 1348 7936
rect 1259 7905 1271 7908
rect 1213 7899 1271 7905
rect 1320 7732 1348 7908
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 1412 7868 1440 7899
rect 1486 7896 1492 7948
rect 1544 7896 1550 7948
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 1765 7939 1823 7945
rect 1765 7936 1777 7939
rect 1728 7908 1777 7936
rect 1728 7896 1734 7908
rect 1765 7905 1777 7908
rect 1811 7905 1823 7939
rect 1765 7899 1823 7905
rect 2406 7896 2412 7948
rect 2464 7896 2470 7948
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4614 7936 4620 7948
rect 4120 7908 4620 7936
rect 4120 7896 4126 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7936 4951 7939
rect 5166 7936 5172 7948
rect 4939 7908 5172 7936
rect 4939 7905 4951 7908
rect 4893 7899 4951 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5258 7896 5264 7948
rect 5316 7896 5322 7948
rect 5442 7896 5448 7948
rect 5500 7896 5506 7948
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8864 7936 8892 7967
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9600 7976 10088 8004
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 8619 7908 8653 7936
rect 8864 7908 9229 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 2222 7868 2228 7880
rect 1412 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7868 8539 7871
rect 8588 7868 8616 7899
rect 9398 7896 9404 7948
rect 9456 7896 9462 7948
rect 8754 7868 8760 7880
rect 8527 7840 8760 7868
rect 8527 7837 8539 7840
rect 8481 7831 8539 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 8846 7828 8852 7880
rect 8904 7828 8910 7880
rect 9306 7828 9312 7880
rect 9364 7868 9370 7880
rect 9600 7868 9628 7976
rect 10060 7948 10088 7976
rect 10226 7964 10232 8016
rect 10284 8004 10290 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 10284 7976 11897 8004
rect 10284 7964 10290 7976
rect 11885 7973 11897 7976
rect 11931 7973 11943 8007
rect 12618 8004 12624 8016
rect 11885 7967 11943 7973
rect 12084 7976 12624 8004
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 9950 7936 9956 7948
rect 9723 7908 9956 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10042 7896 10048 7948
rect 10100 7896 10106 7948
rect 10962 7896 10968 7948
rect 11020 7896 11026 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11330 7936 11336 7948
rect 11287 7908 11336 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 9364 7840 9628 7868
rect 9364 7828 9370 7840
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 11146 7868 11152 7880
rect 9916 7840 11152 7868
rect 9916 7828 9922 7840
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 1397 7803 1455 7809
rect 1397 7769 1409 7803
rect 1443 7800 1455 7803
rect 4154 7800 4160 7812
rect 1443 7772 4160 7800
rect 1443 7769 1455 7772
rect 1397 7763 1455 7769
rect 4154 7760 4160 7772
rect 4212 7760 4218 7812
rect 4890 7760 4896 7812
rect 4948 7760 4954 7812
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 5491 7772 9352 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 2038 7732 2044 7744
rect 1320 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7732 2102 7744
rect 2225 7735 2283 7741
rect 2225 7732 2237 7735
rect 2096 7704 2237 7732
rect 2096 7692 2102 7704
rect 2225 7701 2237 7704
rect 2271 7701 2283 7735
rect 2225 7695 2283 7701
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4246 7732 4252 7744
rect 4028 7704 4252 7732
rect 4028 7692 4034 7704
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 6638 7732 6644 7744
rect 4672 7704 6644 7732
rect 4672 7692 4678 7704
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 9122 7732 9128 7744
rect 8711 7704 9128 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9324 7732 9352 7772
rect 9490 7760 9496 7812
rect 9548 7760 9554 7812
rect 11716 7800 11744 7899
rect 9600 7772 11744 7800
rect 9600 7732 9628 7772
rect 9324 7704 9628 7732
rect 10410 7692 10416 7744
rect 10468 7732 10474 7744
rect 10965 7735 11023 7741
rect 10965 7732 10977 7735
rect 10468 7704 10977 7732
rect 10468 7692 10474 7704
rect 10965 7701 10977 7704
rect 11011 7701 11023 7735
rect 11808 7732 11836 7899
rect 11900 7800 11928 7967
rect 12084 7945 12112 7976
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 12728 8004 12756 8044
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 13262 8072 13268 8084
rect 12860 8044 13268 8072
rect 12860 8032 12866 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 13688 8044 13768 8072
rect 13688 8032 13694 8044
rect 13740 8013 13768 8044
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 15102 8072 15108 8084
rect 14700 8044 15108 8072
rect 14700 8032 14706 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15286 8032 15292 8084
rect 15344 8032 15350 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 15436 8044 15577 8072
rect 15436 8032 15442 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 15838 8032 15844 8084
rect 15896 8072 15902 8084
rect 16482 8072 16488 8084
rect 15896 8044 16488 8072
rect 15896 8032 15902 8044
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 17092 8044 17141 8072
rect 17092 8032 17098 8044
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 18509 8075 18567 8081
rect 18509 8041 18521 8075
rect 18555 8072 18567 8075
rect 18690 8072 18696 8084
rect 18555 8044 18696 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 20625 8075 20683 8081
rect 19024 8044 20576 8072
rect 19024 8032 19030 8044
rect 13541 8007 13599 8013
rect 12728 7976 13308 8004
rect 13280 7948 13308 7976
rect 13541 7973 13553 8007
rect 13587 7973 13599 8007
rect 13541 7967 13599 7973
rect 13725 8007 13783 8013
rect 13725 7973 13737 8007
rect 13771 8004 13783 8007
rect 13771 7976 15056 8004
rect 13771 7973 13783 7976
rect 13725 7967 13783 7973
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7905 12127 7939
rect 12069 7899 12127 7905
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7905 12219 7939
rect 12161 7899 12219 7905
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12434 7936 12440 7948
rect 12391 7908 12440 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 12176 7868 12204 7899
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 12618 7868 12624 7880
rect 12176 7840 12624 7868
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 13188 7868 13216 7899
rect 13262 7896 13268 7948
rect 13320 7896 13326 7948
rect 13556 7936 13584 7967
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 13556 7908 13645 7936
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 13998 7936 14004 7948
rect 13863 7908 14004 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13538 7868 13544 7880
rect 13188 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13170 7800 13176 7812
rect 11900 7772 13176 7800
rect 13170 7760 13176 7772
rect 13228 7760 13234 7812
rect 13648 7800 13676 7899
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 14090 7896 14096 7948
rect 14148 7896 14154 7948
rect 14182 7896 14188 7948
rect 14240 7896 14246 7948
rect 14366 7896 14372 7948
rect 14424 7896 14430 7948
rect 14458 7896 14464 7948
rect 14516 7896 14522 7948
rect 14734 7896 14740 7948
rect 14792 7896 14798 7948
rect 14918 7896 14924 7948
rect 14976 7896 14982 7948
rect 15028 7945 15056 7976
rect 15304 7955 15332 8032
rect 15285 7949 15343 7955
rect 15013 7939 15071 7945
rect 15013 7905 15025 7939
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7905 15163 7939
rect 15285 7915 15297 7949
rect 15331 7915 15343 7949
rect 15378 7930 15384 7982
rect 15436 7930 15442 7982
rect 16390 7964 16396 8016
rect 16448 8004 16454 8016
rect 16850 8004 16856 8016
rect 16448 7976 16856 8004
rect 16448 7964 16454 7976
rect 16850 7964 16856 7976
rect 16908 8004 16914 8016
rect 16908 7976 17172 8004
rect 16908 7964 16914 7976
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15285 7909 15343 7915
rect 15105 7899 15163 7905
rect 15488 7908 15669 7936
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14826 7868 14832 7880
rect 13964 7840 14832 7868
rect 13964 7828 13970 7840
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 15132 7868 15160 7899
rect 15488 7868 15516 7908
rect 15657 7905 15669 7908
rect 15703 7936 15715 7939
rect 15703 7908 16972 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 16577 7871 16635 7877
rect 16577 7868 16589 7871
rect 15132 7840 15516 7868
rect 15672 7840 16589 7868
rect 13280 7772 13676 7800
rect 12158 7732 12164 7744
rect 11808 7704 12164 7732
rect 10965 7695 11023 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12618 7692 12624 7744
rect 12676 7692 12682 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 13280 7732 13308 7772
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 14424 7772 15393 7800
rect 14424 7760 14430 7772
rect 15381 7769 15393 7772
rect 15427 7769 15439 7803
rect 15381 7763 15439 7769
rect 12768 7704 13308 7732
rect 12768 7692 12774 7704
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13504 7704 13921 7732
rect 13504 7692 13510 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14553 7735 14611 7741
rect 14553 7732 14565 7735
rect 14148 7704 14565 7732
rect 14148 7692 14154 7704
rect 14553 7701 14565 7704
rect 14599 7701 14611 7735
rect 14553 7695 14611 7701
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 15672 7732 15700 7840
rect 16577 7837 16589 7840
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16666 7828 16672 7880
rect 16724 7828 16730 7880
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 16944 7800 16972 7908
rect 17034 7896 17040 7948
rect 17092 7896 17098 7948
rect 17144 7936 17172 7976
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 18598 8004 18604 8016
rect 17276 7976 18604 8004
rect 17276 7964 17282 7976
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 19337 8007 19395 8013
rect 19337 8004 19349 8007
rect 18708 7976 19349 8004
rect 18708 7945 18736 7976
rect 19337 7973 19349 7976
rect 19383 8004 19395 8007
rect 19383 7976 19564 8004
rect 19383 7973 19395 7976
rect 19337 7967 19395 7973
rect 17313 7939 17371 7945
rect 17313 7936 17325 7939
rect 17144 7908 17325 7936
rect 17313 7905 17325 7908
rect 17359 7905 17371 7939
rect 17313 7899 17371 7905
rect 18693 7939 18751 7945
rect 18693 7905 18705 7939
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 18782 7896 18788 7948
rect 18840 7896 18846 7948
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 18892 7868 18920 7899
rect 18966 7896 18972 7948
rect 19024 7945 19030 7948
rect 19024 7939 19053 7945
rect 19041 7905 19053 7939
rect 19024 7899 19053 7905
rect 19024 7896 19030 7899
rect 19150 7896 19156 7948
rect 19208 7896 19214 7948
rect 19242 7896 19248 7948
rect 19300 7896 19306 7948
rect 19426 7896 19432 7948
rect 19484 7896 19490 7948
rect 19536 7945 19564 7976
rect 20438 7964 20444 8016
rect 20496 7964 20502 8016
rect 20548 8004 20576 8044
rect 20625 8041 20637 8075
rect 20671 8072 20683 8075
rect 20898 8072 20904 8084
rect 20671 8044 20904 8072
rect 20671 8041 20683 8044
rect 20625 8035 20683 8041
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 21634 8032 21640 8084
rect 21692 8072 21698 8084
rect 22094 8072 22100 8084
rect 21692 8044 22100 8072
rect 21692 8032 21698 8044
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 23017 8075 23075 8081
rect 23017 8041 23029 8075
rect 23063 8072 23075 8075
rect 23198 8072 23204 8084
rect 23063 8044 23204 8072
rect 23063 8041 23075 8044
rect 23017 8035 23075 8041
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 23382 8032 23388 8084
rect 23440 8072 23446 8084
rect 24026 8072 24032 8084
rect 23440 8044 24032 8072
rect 23440 8032 23446 8044
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 24578 8072 24584 8084
rect 24360 8044 24584 8072
rect 24360 8032 24366 8044
rect 24578 8032 24584 8044
rect 24636 8032 24642 8084
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 25004 8044 25452 8072
rect 25004 8032 25010 8044
rect 21266 8004 21272 8016
rect 20548 7976 21272 8004
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 21821 8007 21879 8013
rect 21821 7973 21833 8007
rect 21867 8004 21879 8007
rect 22370 8004 22376 8016
rect 21867 7976 22376 8004
rect 21867 7973 21879 7976
rect 21821 7967 21879 7973
rect 22370 7964 22376 7976
rect 22428 8004 22434 8016
rect 25038 8004 25044 8016
rect 22428 7976 25044 8004
rect 22428 7964 22434 7976
rect 25038 7964 25044 7976
rect 25096 7964 25102 8016
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7905 19579 7939
rect 19521 7899 19579 7905
rect 19705 7939 19763 7945
rect 19705 7905 19717 7939
rect 19751 7936 19763 7939
rect 19794 7936 19800 7948
rect 19751 7908 19800 7936
rect 19751 7905 19763 7908
rect 19705 7899 19763 7905
rect 19794 7896 19800 7908
rect 19852 7896 19858 7948
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20346 7936 20352 7948
rect 19944 7908 20352 7936
rect 19944 7896 19950 7908
rect 20346 7896 20352 7908
rect 20404 7896 20410 7948
rect 20456 7936 20484 7964
rect 20533 7939 20591 7945
rect 20533 7936 20545 7939
rect 20456 7908 20545 7936
rect 20533 7905 20545 7908
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 20622 7896 20628 7948
rect 20680 7896 20686 7948
rect 20990 7896 20996 7948
rect 21048 7936 21054 7948
rect 22002 7936 22008 7948
rect 21048 7908 22008 7936
rect 21048 7896 21054 7908
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 22094 7896 22100 7948
rect 22152 7896 22158 7948
rect 22646 7896 22652 7948
rect 22704 7896 22710 7948
rect 23201 7939 23259 7945
rect 23201 7905 23213 7939
rect 23247 7936 23259 7939
rect 23382 7936 23388 7948
rect 23247 7908 23388 7936
rect 23247 7905 23259 7908
rect 23201 7899 23259 7905
rect 23382 7896 23388 7908
rect 23440 7896 23446 7948
rect 23474 7896 23480 7948
rect 23532 7896 23538 7948
rect 23658 7896 23664 7948
rect 23716 7936 23722 7948
rect 24026 7936 24032 7948
rect 23716 7908 24032 7936
rect 23716 7896 23722 7908
rect 24026 7896 24032 7908
rect 24084 7936 24090 7948
rect 24084 7908 24440 7936
rect 24084 7896 24090 7908
rect 19334 7868 19340 7880
rect 18288 7840 19340 7868
rect 18288 7828 18294 7840
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 20438 7828 20444 7880
rect 20496 7868 20502 7880
rect 23293 7871 23351 7877
rect 23293 7868 23305 7871
rect 20496 7840 23305 7868
rect 20496 7828 20502 7840
rect 23293 7837 23305 7840
rect 23339 7837 23351 7871
rect 23293 7831 23351 7837
rect 19613 7803 19671 7809
rect 19613 7800 19625 7803
rect 16944 7772 19625 7800
rect 19613 7769 19625 7772
rect 19659 7769 19671 7803
rect 19613 7763 19671 7769
rect 20070 7760 20076 7812
rect 20128 7800 20134 7812
rect 20128 7772 20392 7800
rect 20128 7760 20134 7772
rect 14884 7704 15700 7732
rect 14884 7692 14890 7704
rect 16298 7692 16304 7744
rect 16356 7732 16362 7744
rect 16393 7735 16451 7741
rect 16393 7732 16405 7735
rect 16356 7704 16405 7732
rect 16356 7692 16362 7704
rect 16393 7701 16405 7704
rect 16439 7701 16451 7735
rect 16393 7695 16451 7701
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 16724 7704 17325 7732
rect 16724 7692 16730 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17313 7695 17371 7701
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 19242 7732 19248 7744
rect 18748 7704 19248 7732
rect 18748 7692 18754 7704
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 20254 7732 20260 7744
rect 19392 7704 20260 7732
rect 19392 7692 19398 7704
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 20364 7732 20392 7772
rect 20530 7760 20536 7812
rect 20588 7800 20594 7812
rect 21634 7800 21640 7812
rect 20588 7772 21640 7800
rect 20588 7760 20594 7772
rect 21634 7760 21640 7772
rect 21692 7760 21698 7812
rect 22830 7800 22836 7812
rect 22388 7772 22836 7800
rect 20714 7732 20720 7744
rect 20364 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 21821 7735 21879 7741
rect 21821 7732 21833 7735
rect 21140 7704 21833 7732
rect 21140 7692 21146 7704
rect 21821 7701 21833 7704
rect 21867 7701 21879 7735
rect 21821 7695 21879 7701
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7732 22339 7735
rect 22388 7732 22416 7772
rect 22830 7760 22836 7772
rect 22888 7760 22894 7812
rect 23385 7803 23443 7809
rect 23385 7769 23397 7803
rect 23431 7800 23443 7803
rect 23842 7800 23848 7812
rect 23431 7772 23848 7800
rect 23431 7769 23443 7772
rect 23385 7763 23443 7769
rect 23842 7760 23848 7772
rect 23900 7760 23906 7812
rect 22327 7704 22416 7732
rect 22465 7735 22523 7741
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 22465 7701 22477 7735
rect 22511 7732 22523 7735
rect 22646 7732 22652 7744
rect 22511 7704 22652 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 24305 7735 24363 7741
rect 24305 7732 24317 7735
rect 23808 7704 24317 7732
rect 23808 7692 23814 7704
rect 24305 7701 24317 7704
rect 24351 7701 24363 7735
rect 24412 7732 24440 7908
rect 24486 7896 24492 7948
rect 24544 7896 24550 7948
rect 24581 7939 24639 7945
rect 24581 7905 24593 7939
rect 24627 7936 24639 7939
rect 24670 7936 24676 7948
rect 24627 7908 24676 7936
rect 24627 7905 24639 7908
rect 24581 7899 24639 7905
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 24765 7939 24823 7945
rect 24765 7905 24777 7939
rect 24811 7905 24823 7939
rect 24765 7899 24823 7905
rect 24780 7868 24808 7899
rect 24854 7896 24860 7948
rect 24912 7936 24918 7948
rect 24912 7908 25084 7936
rect 24912 7896 24918 7908
rect 24949 7871 25007 7877
rect 24949 7868 24961 7871
rect 24780 7840 24961 7868
rect 24949 7837 24961 7840
rect 24995 7837 25007 7871
rect 25056 7868 25084 7908
rect 25130 7896 25136 7948
rect 25188 7896 25194 7948
rect 25314 7896 25320 7948
rect 25372 7896 25378 7948
rect 25424 7945 25452 8044
rect 25774 8032 25780 8084
rect 25832 8072 25838 8084
rect 28077 8075 28135 8081
rect 28077 8072 28089 8075
rect 25832 8044 28089 8072
rect 25832 8032 25838 8044
rect 28077 8041 28089 8044
rect 28123 8041 28135 8075
rect 28077 8035 28135 8041
rect 28718 8032 28724 8084
rect 28776 8032 28782 8084
rect 29546 8032 29552 8084
rect 29604 8032 29610 8084
rect 29638 8032 29644 8084
rect 29696 8072 29702 8084
rect 29914 8072 29920 8084
rect 29696 8044 29920 8072
rect 29696 8032 29702 8044
rect 29914 8032 29920 8044
rect 29972 8032 29978 8084
rect 30006 8032 30012 8084
rect 30064 8072 30070 8084
rect 30745 8075 30803 8081
rect 30745 8072 30757 8075
rect 30064 8044 30757 8072
rect 30064 8032 30070 8044
rect 30745 8041 30757 8044
rect 30791 8072 30803 8075
rect 31570 8072 31576 8084
rect 30791 8044 31576 8072
rect 30791 8041 30803 8044
rect 30745 8035 30803 8041
rect 31570 8032 31576 8044
rect 31628 8032 31634 8084
rect 25516 7976 25912 8004
rect 25409 7939 25467 7945
rect 25409 7905 25421 7939
rect 25455 7905 25467 7939
rect 25409 7899 25467 7905
rect 25225 7871 25283 7877
rect 25225 7868 25237 7871
rect 25056 7840 25237 7868
rect 24949 7831 25007 7837
rect 25225 7837 25237 7840
rect 25271 7868 25283 7871
rect 25516 7868 25544 7976
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 25271 7840 25544 7868
rect 25608 7908 25697 7936
rect 25271 7837 25283 7840
rect 25225 7831 25283 7837
rect 24673 7803 24731 7809
rect 24673 7769 24685 7803
rect 24719 7800 24731 7803
rect 25498 7800 25504 7812
rect 24719 7772 25504 7800
rect 24719 7769 24731 7772
rect 24673 7763 24731 7769
rect 25498 7760 25504 7772
rect 25556 7760 25562 7812
rect 25608 7800 25636 7908
rect 25685 7905 25697 7908
rect 25731 7905 25743 7939
rect 25884 7936 25912 7976
rect 25958 7964 25964 8016
rect 26016 8004 26022 8016
rect 27249 8007 27307 8013
rect 27249 8004 27261 8007
rect 26016 7976 27261 8004
rect 26016 7964 26022 7976
rect 27249 7973 27261 7976
rect 27295 7973 27307 8007
rect 29270 8004 29276 8016
rect 27249 7967 27307 7973
rect 27540 7976 29276 8004
rect 26053 7939 26111 7945
rect 26053 7936 26065 7939
rect 25884 7908 26065 7936
rect 25685 7899 25743 7905
rect 26053 7905 26065 7908
rect 26099 7936 26111 7939
rect 26326 7936 26332 7948
rect 26099 7908 26332 7936
rect 26099 7905 26111 7908
rect 26053 7899 26111 7905
rect 26326 7896 26332 7908
rect 26384 7896 26390 7948
rect 26697 7939 26755 7945
rect 26697 7905 26709 7939
rect 26743 7936 26755 7939
rect 26878 7936 26884 7948
rect 26743 7908 26884 7936
rect 26743 7905 26755 7908
rect 26697 7899 26755 7905
rect 26878 7896 26884 7908
rect 26936 7896 26942 7948
rect 26970 7896 26976 7948
rect 27028 7896 27034 7948
rect 27540 7945 27568 7976
rect 29270 7964 29276 7976
rect 29328 8004 29334 8016
rect 29564 8004 29592 8032
rect 29328 7976 30880 8004
rect 29328 7964 29334 7976
rect 27157 7939 27215 7945
rect 27157 7905 27169 7939
rect 27203 7905 27215 7939
rect 27157 7899 27215 7905
rect 27525 7939 27583 7945
rect 27525 7905 27537 7939
rect 27571 7905 27583 7939
rect 27525 7899 27583 7905
rect 25958 7828 25964 7880
rect 26016 7868 26022 7880
rect 26988 7868 27016 7896
rect 26016 7840 27016 7868
rect 27172 7868 27200 7899
rect 27890 7896 27896 7948
rect 27948 7896 27954 7948
rect 27982 7896 27988 7948
rect 28040 7936 28046 7948
rect 28261 7939 28319 7945
rect 28261 7936 28273 7939
rect 28040 7908 28273 7936
rect 28040 7896 28046 7908
rect 28261 7905 28273 7908
rect 28307 7905 28319 7939
rect 28261 7899 28319 7905
rect 28350 7896 28356 7948
rect 28408 7936 28414 7948
rect 28537 7939 28595 7945
rect 28537 7936 28549 7939
rect 28408 7908 28549 7936
rect 28408 7896 28414 7908
rect 28537 7905 28549 7908
rect 28583 7905 28595 7939
rect 28537 7899 28595 7905
rect 28626 7896 28632 7948
rect 28684 7936 28690 7948
rect 29380 7945 29408 7976
rect 28935 7939 28993 7945
rect 28935 7936 28947 7939
rect 28684 7908 28947 7936
rect 28684 7896 28690 7908
rect 28935 7905 28947 7908
rect 28981 7905 28993 7939
rect 28935 7899 28993 7905
rect 29089 7939 29147 7945
rect 29089 7905 29101 7939
rect 29135 7905 29147 7939
rect 29089 7899 29147 7905
rect 29365 7939 29423 7945
rect 29365 7905 29377 7939
rect 29411 7905 29423 7939
rect 29365 7899 29423 7905
rect 28074 7868 28080 7880
rect 27172 7840 28080 7868
rect 26016 7828 26022 7840
rect 25682 7800 25688 7812
rect 25608 7772 25688 7800
rect 25682 7760 25688 7772
rect 25740 7760 25746 7812
rect 25774 7760 25780 7812
rect 25832 7800 25838 7812
rect 26988 7800 27016 7840
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28368 7868 28396 7896
rect 28276 7840 28396 7868
rect 28166 7800 28172 7812
rect 25832 7772 26648 7800
rect 26988 7772 28172 7800
rect 25832 7760 25838 7772
rect 25976 7741 26004 7772
rect 25961 7735 26019 7741
rect 25961 7732 25973 7735
rect 24412 7704 25973 7732
rect 24305 7695 24363 7701
rect 25961 7701 25973 7704
rect 26007 7701 26019 7735
rect 25961 7695 26019 7701
rect 26050 7692 26056 7744
rect 26108 7732 26114 7744
rect 26237 7735 26295 7741
rect 26237 7732 26249 7735
rect 26108 7704 26249 7732
rect 26108 7692 26114 7704
rect 26237 7701 26249 7704
rect 26283 7701 26295 7735
rect 26237 7695 26295 7701
rect 26510 7692 26516 7744
rect 26568 7692 26574 7744
rect 26620 7732 26648 7772
rect 28166 7760 28172 7772
rect 28224 7760 28230 7812
rect 28276 7732 28304 7840
rect 28350 7760 28356 7812
rect 28408 7760 28414 7812
rect 28445 7803 28503 7809
rect 28445 7769 28457 7803
rect 28491 7800 28503 7803
rect 28994 7800 29000 7812
rect 28491 7772 29000 7800
rect 28491 7769 28503 7772
rect 28445 7763 28503 7769
rect 28994 7760 29000 7772
rect 29052 7760 29058 7812
rect 29104 7800 29132 7899
rect 29546 7896 29552 7948
rect 29604 7896 29610 7948
rect 29914 7896 29920 7948
rect 29972 7896 29978 7948
rect 30466 7896 30472 7948
rect 30524 7896 30530 7948
rect 30852 7945 30880 7976
rect 30837 7939 30895 7945
rect 30837 7905 30849 7939
rect 30883 7936 30895 7939
rect 31754 7936 31760 7948
rect 30883 7908 31760 7936
rect 30883 7905 30895 7908
rect 30837 7899 30895 7905
rect 31754 7896 31760 7908
rect 31812 7896 31818 7948
rect 29178 7828 29184 7880
rect 29236 7868 29242 7880
rect 29564 7868 29592 7896
rect 30484 7868 30512 7896
rect 29236 7840 30512 7868
rect 29236 7828 29242 7840
rect 30006 7800 30012 7812
rect 29104 7772 30012 7800
rect 30006 7760 30012 7772
rect 30064 7760 30070 7812
rect 30282 7760 30288 7812
rect 30340 7760 30346 7812
rect 26620 7704 28304 7732
rect 29457 7735 29515 7741
rect 29457 7701 29469 7735
rect 29503 7732 29515 7735
rect 29638 7732 29644 7744
rect 29503 7704 29644 7732
rect 29503 7701 29515 7704
rect 29457 7695 29515 7701
rect 29638 7692 29644 7704
rect 29696 7692 29702 7744
rect 552 7642 31648 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 11436 7642
rect 11488 7590 11500 7642
rect 11552 7590 11564 7642
rect 11616 7590 11628 7642
rect 11680 7590 11692 7642
rect 11744 7590 19210 7642
rect 19262 7590 19274 7642
rect 19326 7590 19338 7642
rect 19390 7590 19402 7642
rect 19454 7590 19466 7642
rect 19518 7590 26984 7642
rect 27036 7590 27048 7642
rect 27100 7590 27112 7642
rect 27164 7590 27176 7642
rect 27228 7590 27240 7642
rect 27292 7590 31648 7642
rect 552 7568 31648 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 1946 7528 1952 7540
rect 1636 7500 1952 7528
rect 1636 7488 1642 7500
rect 1946 7488 1952 7500
rect 2004 7488 2010 7540
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 4246 7528 4252 7540
rect 3752 7500 4252 7528
rect 3752 7488 3758 7500
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4798 7488 4804 7540
rect 4856 7488 4862 7540
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 5040 7500 5089 7528
rect 5040 7488 5046 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7282 7528 7288 7540
rect 7055 7500 7288 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 9582 7528 9588 7540
rect 9456 7500 9588 7528
rect 9456 7488 9462 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7528 10287 7531
rect 10962 7528 10968 7540
rect 10275 7500 10968 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11514 7528 11520 7540
rect 11112 7500 11520 7528
rect 11112 7488 11118 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 11848 7500 14473 7528
rect 11848 7488 11854 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14461 7491 14519 7497
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 14826 7528 14832 7540
rect 14608 7500 14832 7528
rect 14608 7488 14614 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15197 7531 15255 7537
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15286 7528 15292 7540
rect 15243 7500 15292 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15528 7500 16129 7528
rect 15528 7488 15534 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 16761 7531 16819 7537
rect 16761 7497 16773 7531
rect 16807 7528 16819 7531
rect 16850 7528 16856 7540
rect 16807 7500 16856 7528
rect 16807 7497 16819 7500
rect 16761 7491 16819 7497
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 16942 7488 16948 7540
rect 17000 7488 17006 7540
rect 17494 7488 17500 7540
rect 17552 7528 17558 7540
rect 18138 7528 18144 7540
rect 17552 7500 18144 7528
rect 17552 7488 17558 7500
rect 18138 7488 18144 7500
rect 18196 7528 18202 7540
rect 20438 7528 20444 7540
rect 18196 7500 20444 7528
rect 18196 7488 18202 7500
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 20864 7500 21465 7528
rect 20864 7488 20870 7500
rect 21453 7497 21465 7500
rect 21499 7528 21511 7531
rect 21818 7528 21824 7540
rect 21499 7500 21824 7528
rect 21499 7497 21511 7500
rect 21453 7491 21511 7497
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 23198 7528 23204 7540
rect 22204 7500 23204 7528
rect 1670 7420 1676 7472
rect 1728 7420 1734 7472
rect 2222 7420 2228 7472
rect 2280 7420 2286 7472
rect 1688 7392 1716 7420
rect 2240 7392 2268 7420
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 1688 7364 2084 7392
rect 2240 7364 2789 7392
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7324 1547 7327
rect 1578 7324 1584 7336
rect 1535 7296 1584 7324
rect 1535 7293 1547 7296
rect 1489 7287 1547 7293
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 1854 7324 1860 7336
rect 1811 7296 1860 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 1394 7216 1400 7268
rect 1452 7256 1458 7268
rect 1780 7256 1808 7287
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 1946 7284 1952 7336
rect 2004 7284 2010 7336
rect 2056 7333 2084 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 4304 7364 4537 7392
rect 4304 7352 4310 7364
rect 4525 7361 4537 7364
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 4816 7336 4844 7488
rect 4908 7392 4936 7488
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10321 7463 10379 7469
rect 10008 7432 10272 7460
rect 10008 7420 10014 7432
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 4908 7364 5549 7392
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 7190 7392 7196 7404
rect 5537 7355 5595 7361
rect 6472 7364 7196 7392
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 2130 7284 2136 7336
rect 2188 7324 2194 7336
rect 2225 7327 2283 7333
rect 2225 7324 2237 7327
rect 2188 7296 2237 7324
rect 2188 7284 2194 7296
rect 2225 7293 2237 7296
rect 2271 7293 2283 7327
rect 2225 7287 2283 7293
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3568 7296 3893 7324
rect 3568 7284 3574 7296
rect 3881 7293 3893 7296
rect 3927 7324 3939 7327
rect 3970 7324 3976 7336
rect 3927 7296 3976 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 1452 7228 1808 7256
rect 1452 7216 1458 7228
rect 3602 7216 3608 7268
rect 3660 7256 3666 7268
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3660 7228 4077 7256
rect 3660 7216 3666 7228
rect 4065 7225 4077 7228
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4172 7188 4200 7287
rect 4338 7284 4344 7336
rect 4396 7284 4402 7336
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 4706 7324 4712 7336
rect 4663 7296 4712 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 4448 7256 4476 7287
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4798 7284 4804 7336
rect 4856 7284 4862 7336
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 4948 7296 5273 7324
rect 4948 7284 4954 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 5350 7284 5356 7336
rect 5408 7284 5414 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 6472 7324 6500 7364
rect 7190 7352 7196 7364
rect 7248 7392 7254 7404
rect 8202 7392 8208 7404
rect 7248 7364 8208 7392
rect 7248 7352 7254 7364
rect 8202 7352 8208 7364
rect 8260 7392 8266 7404
rect 8260 7364 8616 7392
rect 8260 7352 8266 7364
rect 5491 7296 6500 7324
rect 6549 7327 6607 7333
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 6730 7324 6736 7336
rect 6595 7296 6736 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 8588 7333 8616 7364
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 10244 7401 10272 7432
rect 10321 7429 10333 7463
rect 10367 7460 10379 7463
rect 12158 7460 12164 7472
rect 10367 7432 12164 7460
rect 10367 7429 10379 7432
rect 10321 7423 10379 7429
rect 12158 7420 12164 7432
rect 12216 7460 12222 7472
rect 12216 7432 15056 7460
rect 12216 7420 12222 7432
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9140 7364 10057 7392
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 7064 7296 8401 7324
rect 7064 7284 7070 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 8294 7256 8300 7268
rect 4448 7228 8300 7256
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 8404 7256 8432 7287
rect 8846 7284 8852 7336
rect 8904 7284 8910 7336
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9140 7256 9168 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7361 10287 7395
rect 14734 7392 14740 7404
rect 10229 7355 10287 7361
rect 10336 7364 14740 7392
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 10336 7324 10364 7364
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15028 7392 15056 7432
rect 15215 7432 20209 7460
rect 15215 7392 15243 7432
rect 15028 7364 15243 7392
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 15896 7364 16620 7392
rect 15896 7352 15902 7364
rect 9263 7296 10364 7324
rect 10413 7327 10471 7333
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 10413 7293 10425 7327
rect 10459 7324 10471 7327
rect 10502 7324 10508 7336
rect 10459 7296 10508 7324
rect 10459 7293 10471 7296
rect 10413 7287 10471 7293
rect 8404 7228 9168 7256
rect 4028 7160 4200 7188
rect 4801 7191 4859 7197
rect 4028 7148 4034 7160
rect 4801 7157 4813 7191
rect 4847 7188 4859 7191
rect 5534 7188 5540 7200
rect 4847 7160 5540 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 6638 7148 6644 7200
rect 6696 7148 6702 7200
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 9232 7188 9260 7287
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 11974 7324 11980 7336
rect 11204 7296 11980 7324
rect 11204 7284 11210 7296
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12897 7327 12955 7333
rect 12124 7296 12848 7324
rect 12124 7284 12130 7296
rect 10134 7216 10140 7268
rect 10192 7256 10198 7268
rect 12710 7256 12716 7268
rect 10192 7228 12716 7256
rect 10192 7216 10198 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 12820 7256 12848 7296
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 12986 7324 12992 7336
rect 12943 7296 12992 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 14550 7324 14556 7336
rect 13320 7296 14556 7324
rect 13320 7284 13326 7296
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 14642 7284 14648 7336
rect 14700 7284 14706 7336
rect 14918 7284 14924 7336
rect 14976 7284 14982 7336
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15286 7324 15292 7336
rect 15151 7296 15292 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15120 7256 15148 7287
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15381 7327 15439 7333
rect 15381 7302 15393 7327
rect 15427 7302 15439 7327
rect 12820 7228 15148 7256
rect 15378 7250 15384 7302
rect 15436 7250 15442 7302
rect 15470 7284 15476 7336
rect 15528 7284 15534 7336
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 15565 7287 15623 7293
rect 7892 7160 9260 7188
rect 7892 7148 7898 7160
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10226 7188 10232 7200
rect 9824 7160 10232 7188
rect 9824 7148 9830 7160
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 12526 7188 12532 7200
rect 11204 7160 12532 7188
rect 11204 7148 11210 7160
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12802 7148 12808 7200
rect 12860 7148 12866 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 15580 7188 15608 7287
rect 15654 7284 15660 7336
rect 15712 7284 15718 7336
rect 16298 7284 16304 7336
rect 16356 7284 16362 7336
rect 16390 7284 16396 7336
rect 16448 7284 16454 7336
rect 16592 7333 16620 7364
rect 16850 7352 16856 7404
rect 16908 7392 16914 7404
rect 17402 7392 17408 7404
rect 16908 7364 17408 7392
rect 16908 7352 16914 7364
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 18046 7352 18052 7404
rect 18104 7392 18110 7404
rect 18782 7392 18788 7404
rect 18104 7364 18788 7392
rect 18104 7352 18110 7364
rect 18782 7352 18788 7364
rect 18840 7392 18846 7404
rect 19518 7392 19524 7404
rect 18840 7364 19524 7392
rect 18840 7352 18846 7364
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 20181 7392 20209 7432
rect 20254 7420 20260 7472
rect 20312 7460 20318 7472
rect 20622 7460 20628 7472
rect 20312 7432 20628 7460
rect 20312 7420 20318 7432
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 21232 7432 21526 7460
rect 21232 7420 21238 7432
rect 20717 7395 20775 7401
rect 20181 7364 20668 7392
rect 16577 7327 16635 7333
rect 16577 7293 16589 7327
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 19794 7324 19800 7336
rect 16816 7296 19800 7324
rect 16816 7284 16822 7296
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 20070 7284 20076 7336
rect 20128 7324 20134 7336
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 20128 7296 20177 7324
rect 20128 7284 20134 7296
rect 20165 7293 20177 7296
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 20254 7284 20260 7336
rect 20312 7284 20318 7336
rect 20456 7333 20484 7364
rect 20441 7327 20499 7333
rect 20441 7293 20453 7327
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7293 20591 7327
rect 20640 7324 20668 7364
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 20898 7392 20904 7404
rect 20763 7364 20904 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 20806 7324 20812 7336
rect 20640 7296 20812 7324
rect 20533 7287 20591 7293
rect 17129 7259 17187 7265
rect 17129 7256 17141 7259
rect 16592 7228 17141 7256
rect 16592 7200 16620 7228
rect 17129 7225 17141 7228
rect 17175 7225 17187 7259
rect 17129 7219 17187 7225
rect 17678 7216 17684 7268
rect 17736 7256 17742 7268
rect 17954 7256 17960 7268
rect 17736 7228 17960 7256
rect 17736 7216 17742 7228
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 13228 7160 15608 7188
rect 13228 7148 13234 7160
rect 16574 7148 16580 7200
rect 16632 7148 16638 7200
rect 16929 7191 16987 7197
rect 16929 7157 16941 7191
rect 16975 7188 16987 7191
rect 17218 7188 17224 7200
rect 16975 7160 17224 7188
rect 16975 7157 16987 7160
rect 16929 7151 16987 7157
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 20548 7188 20576 7287
rect 20806 7284 20812 7296
rect 20864 7284 20870 7336
rect 20990 7284 20996 7336
rect 21048 7284 21054 7336
rect 21174 7284 21180 7336
rect 21232 7284 21238 7336
rect 21498 7333 21526 7432
rect 22204 7392 22232 7500
rect 23198 7488 23204 7500
rect 23256 7488 23262 7540
rect 23842 7488 23848 7540
rect 23900 7488 23906 7540
rect 24762 7528 24768 7540
rect 23952 7500 24768 7528
rect 22281 7463 22339 7469
rect 22281 7429 22293 7463
rect 22327 7429 22339 7463
rect 23952 7460 23980 7500
rect 24762 7488 24768 7500
rect 24820 7488 24826 7540
rect 24946 7488 24952 7540
rect 25004 7528 25010 7540
rect 25961 7531 26019 7537
rect 25961 7528 25973 7531
rect 25004 7500 25973 7528
rect 25004 7488 25010 7500
rect 25961 7497 25973 7500
rect 26007 7497 26019 7531
rect 25961 7491 26019 7497
rect 26142 7488 26148 7540
rect 26200 7488 26206 7540
rect 27433 7531 27491 7537
rect 27433 7497 27445 7531
rect 27479 7528 27491 7531
rect 28350 7528 28356 7540
rect 27479 7500 28356 7528
rect 27479 7497 27491 7500
rect 27433 7491 27491 7497
rect 28350 7488 28356 7500
rect 28408 7488 28414 7540
rect 28534 7488 28540 7540
rect 28592 7528 28598 7540
rect 29273 7531 29331 7537
rect 29273 7528 29285 7531
rect 28592 7500 29285 7528
rect 28592 7488 28598 7500
rect 29273 7497 29285 7500
rect 29319 7497 29331 7531
rect 29273 7491 29331 7497
rect 30098 7488 30104 7540
rect 30156 7528 30162 7540
rect 30377 7531 30435 7537
rect 30377 7528 30389 7531
rect 30156 7500 30389 7528
rect 30156 7488 30162 7500
rect 30377 7497 30389 7500
rect 30423 7497 30435 7531
rect 30377 7491 30435 7497
rect 30745 7531 30803 7537
rect 30745 7497 30757 7531
rect 30791 7528 30803 7531
rect 30834 7528 30840 7540
rect 30791 7500 30840 7528
rect 30791 7497 30803 7500
rect 30745 7491 30803 7497
rect 30834 7488 30840 7500
rect 30892 7488 30898 7540
rect 22281 7423 22339 7429
rect 22664 7432 23980 7460
rect 21652 7364 22232 7392
rect 22296 7392 22324 7423
rect 22296 7364 22600 7392
rect 21652 7333 21680 7364
rect 21483 7327 21541 7333
rect 21483 7293 21495 7327
rect 21529 7293 21541 7327
rect 21483 7287 21541 7293
rect 21637 7327 21695 7333
rect 21637 7293 21649 7327
rect 21683 7293 21695 7327
rect 21637 7287 21695 7293
rect 21726 7284 21732 7336
rect 21784 7284 21790 7336
rect 21818 7284 21824 7336
rect 21876 7324 21882 7336
rect 22097 7327 22155 7333
rect 22097 7324 22109 7327
rect 21876 7296 22109 7324
rect 21876 7284 21882 7296
rect 22097 7293 22109 7296
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 22278 7284 22284 7336
rect 22336 7324 22342 7336
rect 22572 7333 22600 7364
rect 22664 7333 22692 7432
rect 24118 7420 24124 7472
rect 24176 7460 24182 7472
rect 24394 7460 24400 7472
rect 24176 7432 24400 7460
rect 24176 7420 24182 7432
rect 24394 7420 24400 7432
rect 24452 7420 24458 7472
rect 24578 7420 24584 7472
rect 24636 7460 24642 7472
rect 24673 7463 24731 7469
rect 24673 7460 24685 7463
rect 24636 7432 24685 7460
rect 24636 7420 24642 7432
rect 24673 7429 24685 7432
rect 24719 7429 24731 7463
rect 24673 7423 24731 7429
rect 25038 7420 25044 7472
rect 25096 7460 25102 7472
rect 28552 7460 28580 7488
rect 30650 7460 30656 7472
rect 25096 7432 28580 7460
rect 30116 7432 30656 7460
rect 25096 7420 25102 7432
rect 23198 7352 23204 7404
rect 23256 7392 23262 7404
rect 25406 7392 25412 7404
rect 23256 7364 25412 7392
rect 23256 7352 23262 7364
rect 25406 7352 25412 7364
rect 25464 7352 25470 7404
rect 22373 7327 22431 7333
rect 22373 7324 22385 7327
rect 22336 7296 22385 7324
rect 22336 7284 22342 7296
rect 22373 7293 22385 7296
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 22557 7327 22615 7333
rect 22557 7293 22569 7327
rect 22603 7293 22615 7327
rect 22557 7287 22615 7293
rect 22649 7327 22707 7333
rect 22649 7293 22661 7327
rect 22695 7293 22707 7327
rect 22649 7287 22707 7293
rect 21085 7259 21143 7265
rect 21085 7225 21097 7259
rect 21131 7256 21143 7259
rect 21913 7259 21971 7265
rect 21913 7256 21925 7259
rect 21131 7228 21925 7256
rect 21131 7225 21143 7228
rect 21085 7219 21143 7225
rect 21913 7225 21925 7228
rect 21959 7225 21971 7259
rect 21913 7219 21971 7225
rect 22005 7259 22063 7265
rect 22005 7225 22017 7259
rect 22051 7256 22063 7259
rect 22462 7256 22468 7268
rect 22051 7228 22468 7256
rect 22051 7225 22063 7228
rect 22005 7219 22063 7225
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 17368 7160 20576 7188
rect 17368 7148 17374 7160
rect 20622 7148 20628 7200
rect 20680 7188 20686 7200
rect 22664 7188 22692 7287
rect 22830 7284 22836 7336
rect 22888 7284 22894 7336
rect 22925 7327 22983 7333
rect 22925 7293 22937 7327
rect 22971 7324 22983 7327
rect 24026 7324 24032 7336
rect 22971 7296 24032 7324
rect 22971 7293 22983 7296
rect 22925 7287 22983 7293
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 24121 7327 24179 7333
rect 24121 7293 24133 7327
rect 24167 7324 24179 7327
rect 24394 7324 24400 7336
rect 24167 7296 24400 7324
rect 24167 7293 24179 7296
rect 24121 7287 24179 7293
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 24489 7327 24547 7333
rect 24489 7293 24501 7327
rect 24535 7293 24547 7327
rect 24489 7287 24547 7293
rect 22738 7216 22744 7268
rect 22796 7256 22802 7268
rect 24305 7259 24363 7265
rect 24305 7256 24317 7259
rect 22796 7228 24317 7256
rect 22796 7216 22802 7228
rect 24305 7225 24317 7228
rect 24351 7225 24363 7259
rect 24504 7256 24532 7287
rect 24578 7284 24584 7336
rect 24636 7284 24642 7336
rect 25038 7324 25044 7336
rect 24688 7296 25044 7324
rect 24688 7256 24716 7296
rect 25038 7284 25044 7296
rect 25096 7284 25102 7336
rect 25225 7293 25283 7299
rect 25225 7268 25237 7293
rect 25271 7268 25283 7293
rect 25498 7284 25504 7336
rect 25556 7284 25562 7336
rect 25608 7333 25636 7432
rect 26050 7352 26056 7404
rect 26108 7352 26114 7404
rect 26510 7392 26516 7404
rect 26142 7364 26516 7392
rect 25593 7327 25651 7333
rect 25593 7293 25605 7327
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 25685 7327 25743 7333
rect 25685 7293 25697 7327
rect 25731 7324 25743 7327
rect 26142 7324 26170 7364
rect 26510 7352 26516 7364
rect 26568 7352 26574 7404
rect 28077 7395 28135 7401
rect 28077 7392 28089 7395
rect 27448 7364 28089 7392
rect 27448 7336 27476 7364
rect 28077 7361 28089 7364
rect 28123 7361 28135 7395
rect 28810 7392 28816 7404
rect 28077 7355 28135 7361
rect 28276 7364 28816 7392
rect 25731 7296 26170 7324
rect 25731 7293 25743 7296
rect 25685 7287 25743 7293
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26292 7296 26985 7324
rect 26292 7284 26298 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 27062 7284 27068 7336
rect 27120 7284 27126 7336
rect 27249 7327 27307 7333
rect 27249 7293 27261 7327
rect 27295 7324 27307 7327
rect 27338 7324 27344 7336
rect 27295 7296 27344 7324
rect 27295 7293 27307 7296
rect 27249 7287 27307 7293
rect 27338 7284 27344 7296
rect 27396 7284 27402 7336
rect 27430 7284 27436 7336
rect 27488 7284 27494 7336
rect 28276 7333 28304 7364
rect 28810 7352 28816 7364
rect 28868 7392 28874 7404
rect 29917 7395 29975 7401
rect 29917 7392 29929 7395
rect 28868 7364 29929 7392
rect 28868 7352 28874 7364
rect 29917 7361 29929 7364
rect 29963 7392 29975 7395
rect 30009 7395 30067 7401
rect 30009 7392 30021 7395
rect 29963 7364 30021 7392
rect 29963 7361 29975 7364
rect 29917 7355 29975 7361
rect 30009 7361 30021 7364
rect 30055 7361 30067 7395
rect 30009 7355 30067 7361
rect 27525 7327 27583 7333
rect 27525 7293 27537 7327
rect 27571 7293 27583 7327
rect 27525 7287 27583 7293
rect 28261 7327 28319 7333
rect 28261 7293 28273 7327
rect 28307 7293 28319 7327
rect 28537 7327 28595 7333
rect 28537 7324 28549 7327
rect 28261 7287 28319 7293
rect 28368 7296 28549 7324
rect 24504 7228 24716 7256
rect 24305 7219 24363 7225
rect 24854 7216 24860 7268
rect 24912 7216 24918 7268
rect 25222 7216 25228 7268
rect 25280 7216 25286 7268
rect 25516 7256 25544 7284
rect 25516 7228 26741 7256
rect 20680 7160 22692 7188
rect 24213 7191 24271 7197
rect 20680 7148 20686 7160
rect 24213 7157 24225 7191
rect 24259 7188 24271 7191
rect 24762 7188 24768 7200
rect 24259 7160 24768 7188
rect 24259 7157 24271 7160
rect 24213 7151 24271 7157
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 24946 7148 24952 7200
rect 25004 7188 25010 7200
rect 25317 7191 25375 7197
rect 25317 7188 25329 7191
rect 25004 7160 25329 7188
rect 25004 7148 25010 7160
rect 25317 7157 25329 7160
rect 25363 7157 25375 7191
rect 25317 7151 25375 7157
rect 25777 7191 25835 7197
rect 25777 7157 25789 7191
rect 25823 7188 25835 7191
rect 26050 7188 26056 7200
rect 25823 7160 26056 7188
rect 25823 7157 25835 7160
rect 25777 7151 25835 7157
rect 26050 7148 26056 7160
rect 26108 7148 26114 7200
rect 26713 7188 26741 7228
rect 26786 7216 26792 7268
rect 26844 7256 26850 7268
rect 27540 7256 27568 7287
rect 26844 7228 27568 7256
rect 27801 7259 27859 7265
rect 26844 7216 26850 7228
rect 27801 7225 27813 7259
rect 27847 7256 27859 7259
rect 27982 7256 27988 7268
rect 27847 7228 27988 7256
rect 27847 7225 27859 7228
rect 27801 7219 27859 7225
rect 27982 7216 27988 7228
rect 28040 7216 28046 7268
rect 28166 7216 28172 7268
rect 28224 7256 28230 7268
rect 28368 7256 28396 7296
rect 28537 7293 28549 7296
rect 28583 7293 28595 7327
rect 28537 7287 28595 7293
rect 28718 7284 28724 7336
rect 28776 7324 28782 7336
rect 29178 7324 29184 7336
rect 28776 7296 29184 7324
rect 28776 7284 28782 7296
rect 29178 7284 29184 7296
rect 29236 7284 29242 7336
rect 29454 7284 29460 7336
rect 29512 7284 29518 7336
rect 29549 7327 29607 7333
rect 29549 7293 29561 7327
rect 29595 7324 29607 7327
rect 30116 7324 30144 7432
rect 30650 7420 30656 7432
rect 30708 7420 30714 7472
rect 30282 7352 30288 7404
rect 30340 7392 30346 7404
rect 30340 7364 30696 7392
rect 30340 7352 30346 7364
rect 29595 7296 30144 7324
rect 29595 7293 29607 7296
rect 29549 7287 29607 7293
rect 30374 7284 30380 7336
rect 30432 7284 30438 7336
rect 30668 7333 30696 7364
rect 30653 7327 30711 7333
rect 30653 7293 30665 7327
rect 30699 7293 30711 7327
rect 30653 7287 30711 7293
rect 28224 7228 28396 7256
rect 28445 7259 28503 7265
rect 28224 7216 28230 7228
rect 28445 7225 28457 7259
rect 28491 7256 28503 7259
rect 29086 7256 29092 7268
rect 28491 7228 29092 7256
rect 28491 7225 28503 7228
rect 28445 7219 28503 7225
rect 29086 7216 29092 7228
rect 29144 7256 29150 7268
rect 30098 7256 30104 7268
rect 29144 7228 30104 7256
rect 29144 7216 29150 7228
rect 30098 7216 30104 7228
rect 30156 7216 30162 7268
rect 28626 7188 28632 7200
rect 26713 7160 28632 7188
rect 28626 7148 28632 7160
rect 28684 7148 28690 7200
rect 28721 7191 28779 7197
rect 28721 7157 28733 7191
rect 28767 7188 28779 7191
rect 28994 7188 29000 7200
rect 28767 7160 29000 7188
rect 28767 7157 28779 7160
rect 28721 7151 28779 7157
rect 28994 7148 29000 7160
rect 29052 7148 29058 7200
rect 29178 7148 29184 7200
rect 29236 7188 29242 7200
rect 30190 7188 30196 7200
rect 29236 7160 30196 7188
rect 29236 7148 29242 7160
rect 30190 7148 30196 7160
rect 30248 7148 30254 7200
rect 552 7098 31648 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 12096 7098
rect 12148 7046 12160 7098
rect 12212 7046 12224 7098
rect 12276 7046 12288 7098
rect 12340 7046 12352 7098
rect 12404 7046 19870 7098
rect 19922 7046 19934 7098
rect 19986 7046 19998 7098
rect 20050 7046 20062 7098
rect 20114 7046 20126 7098
rect 20178 7046 27644 7098
rect 27696 7046 27708 7098
rect 27760 7046 27772 7098
rect 27824 7046 27836 7098
rect 27888 7046 27900 7098
rect 27952 7046 31648 7098
rect 552 7024 31648 7046
rect 1578 6944 1584 6996
rect 1636 6944 1642 6996
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 2041 6987 2099 6993
rect 2041 6984 2053 6987
rect 1912 6956 2053 6984
rect 1912 6944 1918 6956
rect 2041 6953 2053 6956
rect 2087 6984 2099 6987
rect 2222 6984 2228 6996
rect 2087 6956 2228 6984
rect 2087 6953 2099 6956
rect 2041 6947 2099 6953
rect 2222 6944 2228 6956
rect 2280 6944 2286 6996
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 4614 6984 4620 6996
rect 2740 6956 4620 6984
rect 2740 6944 2746 6956
rect 1596 6916 1624 6944
rect 3988 6925 4016 6956
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 5258 6944 5264 6996
rect 5316 6984 5322 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 5316 6956 5457 6984
rect 5316 6944 5322 6956
rect 5445 6953 5457 6956
rect 5491 6953 5503 6987
rect 5445 6947 5503 6953
rect 2133 6919 2191 6925
rect 2133 6916 2145 6919
rect 1596 6888 2145 6916
rect 2133 6885 2145 6888
rect 2179 6885 2191 6919
rect 2133 6879 2191 6885
rect 3973 6919 4031 6925
rect 3973 6885 3985 6919
rect 4019 6885 4031 6919
rect 5166 6916 5172 6928
rect 3973 6879 4031 6885
rect 4356 6888 5172 6916
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 1581 6851 1639 6857
rect 1581 6848 1593 6851
rect 1268 6820 1593 6848
rect 1268 6808 1274 6820
rect 1581 6817 1593 6820
rect 1627 6817 1639 6851
rect 1581 6811 1639 6817
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 2409 6851 2467 6857
rect 2409 6848 2421 6851
rect 2096 6820 2421 6848
rect 2096 6808 2102 6820
rect 2409 6817 2421 6820
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3326 6848 3332 6860
rect 3283 6820 3332 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 3602 6808 3608 6860
rect 3660 6808 3666 6860
rect 3694 6808 3700 6860
rect 3752 6808 3758 6860
rect 4062 6808 4068 6860
rect 4120 6808 4126 6860
rect 4154 6808 4160 6860
rect 4212 6808 4218 6860
rect 4356 6857 4384 6888
rect 5166 6876 5172 6888
rect 5224 6876 5230 6928
rect 5460 6916 5488 6947
rect 7650 6944 7656 6996
rect 7708 6944 7714 6996
rect 8938 6944 8944 6996
rect 8996 6944 9002 6996
rect 9490 6984 9496 6996
rect 9324 6956 9496 6984
rect 6638 6916 6644 6928
rect 5460 6888 6644 6916
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4709 6851 4767 6857
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 4798 6848 4804 6860
rect 4755 6820 4804 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 1780 6712 1808 6743
rect 1854 6740 1860 6792
rect 1912 6740 1918 6792
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2314 6780 2320 6792
rect 2271 6752 2320 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3712 6780 3740 6808
rect 4172 6780 4200 6808
rect 2832 6752 3740 6780
rect 3804 6752 4200 6780
rect 5000 6780 5028 6811
rect 5350 6808 5356 6860
rect 5408 6808 5414 6860
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6288 6857 6316 6888
rect 6638 6876 6644 6888
rect 6696 6876 6702 6928
rect 7668 6916 7696 6944
rect 8956 6916 8984 6944
rect 9214 6916 9220 6928
rect 6840 6888 7696 6916
rect 8312 6888 9220 6916
rect 6181 6851 6239 6857
rect 6181 6848 6193 6851
rect 6144 6820 6193 6848
rect 6144 6808 6150 6820
rect 6181 6817 6193 6820
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 5810 6780 5816 6792
rect 5000 6752 5816 6780
rect 2832 6740 2838 6752
rect 2593 6715 2651 6721
rect 2593 6712 2605 6715
rect 1780 6684 2605 6712
rect 2593 6681 2605 6684
rect 2639 6712 2651 6715
rect 2958 6712 2964 6724
rect 2639 6684 2964 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 2958 6672 2964 6684
rect 3016 6712 3022 6724
rect 3602 6712 3608 6724
rect 3016 6684 3608 6712
rect 3016 6672 3022 6684
rect 3602 6672 3608 6684
rect 3660 6672 3666 6724
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3418 6644 3424 6656
rect 3108 6616 3424 6644
rect 3108 6604 3114 6616
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3697 6647 3755 6653
rect 3697 6613 3709 6647
rect 3743 6644 3755 6647
rect 3804 6644 3832 6752
rect 3881 6715 3939 6721
rect 3881 6681 3893 6715
rect 3927 6712 3939 6715
rect 4154 6712 4160 6724
rect 3927 6684 4160 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 3743 6616 3832 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5000 6644 5028 6752
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 6472 6780 6500 6811
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 6840 6848 6868 6888
rect 8312 6857 8340 6888
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 6604 6820 6868 6848
rect 7009 6851 7067 6857
rect 6604 6808 6610 6820
rect 7009 6817 7021 6851
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6848 7803 6851
rect 8297 6851 8355 6857
rect 7791 6820 8064 6848
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 6730 6780 6736 6792
rect 6472 6752 6736 6780
rect 6730 6740 6736 6752
rect 6788 6780 6794 6792
rect 6914 6780 6920 6792
rect 6788 6752 6920 6780
rect 6788 6740 6794 6752
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 7024 6712 7052 6811
rect 6696 6684 7052 6712
rect 6696 6672 6702 6684
rect 4120 6616 5028 6644
rect 4120 6604 4126 6616
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 8036 6644 8064 6820
rect 8297 6817 8309 6851
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 8846 6808 8852 6860
rect 8904 6808 8910 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9324 6848 9352 6956
rect 9490 6944 9496 6956
rect 9548 6984 9554 6996
rect 9548 6956 12848 6984
rect 9548 6944 9554 6956
rect 9766 6916 9772 6928
rect 9416 6888 9772 6916
rect 9416 6857 9444 6888
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 10321 6919 10379 6925
rect 10321 6885 10333 6919
rect 10367 6916 10379 6919
rect 10594 6916 10600 6928
rect 10367 6888 10600 6916
rect 10367 6885 10379 6888
rect 10321 6879 10379 6885
rect 10594 6876 10600 6888
rect 10652 6916 10658 6928
rect 11977 6919 12035 6925
rect 11977 6916 11989 6919
rect 10652 6888 11989 6916
rect 10652 6876 10658 6888
rect 11977 6885 11989 6888
rect 12023 6885 12035 6919
rect 11977 6879 12035 6885
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 12308 6888 12756 6916
rect 12308 6876 12314 6888
rect 8987 6820 9352 6848
rect 9401 6851 9459 6857
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9401 6817 9413 6851
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9582 6808 9588 6860
rect 9640 6808 9646 6860
rect 10134 6808 10140 6860
rect 10192 6848 10198 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 10192 6820 10241 6848
rect 10192 6808 10198 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10229 6811 10287 6817
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 10502 6848 10508 6860
rect 10459 6820 10508 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 10502 6808 10508 6820
rect 10560 6848 10566 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10560 6820 10977 6848
rect 10560 6808 10566 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11241 6851 11299 6857
rect 11241 6848 11253 6851
rect 11204 6820 11253 6848
rect 11204 6808 11210 6820
rect 11241 6817 11253 6820
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 11379 6820 11744 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8435 6752 8769 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 9232 6712 9260 6743
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 11164 6780 11192 6808
rect 9364 6752 11192 6780
rect 9364 6740 9370 6752
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 8168 6684 9260 6712
rect 8168 6672 8174 6684
rect 10226 6672 10232 6724
rect 10284 6712 10290 6724
rect 10284 6684 11192 6712
rect 10284 6672 10290 6684
rect 8294 6644 8300 6656
rect 6328 6616 8300 6644
rect 6328 6604 6334 6616
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8812 6616 9137 6644
rect 8812 6604 8818 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 10042 6604 10048 6656
rect 10100 6644 10106 6656
rect 11054 6644 11060 6656
rect 10100 6616 11060 6644
rect 10100 6604 10106 6616
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11164 6644 11192 6684
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 11609 6715 11667 6721
rect 11609 6712 11621 6715
rect 11296 6684 11621 6712
rect 11296 6672 11302 6684
rect 11609 6681 11621 6684
rect 11655 6681 11667 6715
rect 11609 6675 11667 6681
rect 11716 6644 11744 6820
rect 11790 6808 11796 6860
rect 11848 6808 11854 6860
rect 12069 6851 12127 6857
rect 12069 6817 12081 6851
rect 12115 6848 12127 6851
rect 12342 6848 12348 6860
rect 12115 6820 12348 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 12728 6857 12756 6888
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12400 6820 12633 6848
rect 12400 6808 12406 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 12820 6780 12848 6956
rect 12894 6944 12900 6996
rect 12952 6944 12958 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 14458 6984 14464 6996
rect 13044 6956 14464 6984
rect 13044 6944 13050 6956
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 15381 6987 15439 6993
rect 15381 6984 15393 6987
rect 14700 6956 15393 6984
rect 14700 6944 14706 6956
rect 15381 6953 15393 6956
rect 15427 6953 15439 6987
rect 15381 6947 15439 6953
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 15528 6956 20760 6984
rect 15528 6944 15534 6956
rect 12912 6916 12940 6944
rect 13446 6916 13452 6928
rect 12912 6888 13452 6916
rect 12912 6857 12940 6888
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 13722 6876 13728 6928
rect 13780 6916 13786 6928
rect 13780 6888 15194 6916
rect 13780 6876 13786 6888
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 12986 6808 12992 6860
rect 13044 6808 13050 6860
rect 13262 6808 13268 6860
rect 13320 6808 13326 6860
rect 13372 6820 13676 6848
rect 13078 6780 13084 6792
rect 12820 6752 13084 6780
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 13372 6712 13400 6820
rect 13538 6740 13544 6792
rect 13596 6740 13602 6792
rect 13648 6780 13676 6820
rect 14550 6808 14556 6860
rect 14608 6808 14614 6860
rect 15013 6851 15071 6857
rect 15013 6817 15025 6851
rect 15059 6817 15071 6851
rect 15166 6848 15194 6888
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 16172 6888 16896 6916
rect 16172 6876 16178 6888
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 15166 6820 16313 6848
rect 15013 6811 15071 6817
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 15028 6780 15056 6811
rect 13648 6752 15056 6780
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 15286 6740 15292 6792
rect 15344 6740 15350 6792
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6780 15439 6783
rect 16114 6780 16120 6792
rect 15427 6752 16120 6780
rect 15427 6749 15439 6752
rect 15381 6743 15439 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16316 6780 16344 6811
rect 16482 6808 16488 6860
rect 16540 6808 16546 6860
rect 16868 6857 16896 6888
rect 17770 6876 17776 6928
rect 17828 6916 17834 6928
rect 18385 6919 18443 6925
rect 18385 6916 18397 6919
rect 17828 6888 18397 6916
rect 17828 6876 17834 6888
rect 18385 6885 18397 6888
rect 18431 6885 18443 6919
rect 18385 6879 18443 6885
rect 18601 6919 18659 6925
rect 18601 6885 18613 6919
rect 18647 6916 18659 6919
rect 18690 6916 18696 6928
rect 18647 6888 18696 6916
rect 18647 6885 18659 6888
rect 18601 6879 18659 6885
rect 18690 6876 18696 6888
rect 18748 6876 18754 6928
rect 19518 6876 19524 6928
rect 19576 6916 19582 6928
rect 20732 6916 20760 6956
rect 21174 6944 21180 6996
rect 21232 6984 21238 6996
rect 23014 6984 23020 6996
rect 21232 6956 23020 6984
rect 21232 6944 21238 6956
rect 23014 6944 23020 6956
rect 23072 6944 23078 6996
rect 23382 6984 23388 6996
rect 23124 6956 23388 6984
rect 21450 6916 21456 6928
rect 19576 6888 20300 6916
rect 19576 6876 19582 6888
rect 16761 6851 16819 6857
rect 16761 6848 16773 6851
rect 16592 6820 16773 6848
rect 16592 6780 16620 6820
rect 16761 6817 16773 6820
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6817 16911 6851
rect 16853 6811 16911 6817
rect 17037 6851 17095 6857
rect 17037 6817 17049 6851
rect 17083 6848 17095 6851
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 17083 6820 17141 6848
rect 17083 6817 17095 6820
rect 17037 6811 17095 6817
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17313 6851 17371 6857
rect 17313 6817 17325 6851
rect 17359 6848 17371 6851
rect 17402 6848 17408 6860
rect 17359 6820 17408 6848
rect 17359 6817 17371 6820
rect 17313 6811 17371 6817
rect 16316 6752 16620 6780
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6780 16727 6783
rect 17328 6780 17356 6811
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17494 6808 17500 6860
rect 17552 6808 17558 6860
rect 17678 6808 17684 6860
rect 17736 6808 17742 6860
rect 17862 6808 17868 6860
rect 17920 6808 17926 6860
rect 17954 6808 17960 6860
rect 18012 6848 18018 6860
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 18012 6820 18061 6848
rect 18012 6808 18018 6820
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 16715 6752 17356 6780
rect 17589 6783 17647 6789
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 18156 6780 18184 6811
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 18288 6820 18797 6848
rect 18288 6808 18294 6820
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 18969 6851 19027 6857
rect 18969 6848 18981 6851
rect 18932 6820 18981 6848
rect 18932 6808 18938 6820
rect 18969 6817 18981 6820
rect 19015 6817 19027 6851
rect 19610 6848 19616 6860
rect 18969 6811 19027 6817
rect 19352 6820 19616 6848
rect 19242 6780 19248 6792
rect 17635 6752 19248 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 12032 6684 13400 6712
rect 13449 6715 13507 6721
rect 12032 6672 12038 6684
rect 13449 6681 13461 6715
rect 13495 6712 13507 6715
rect 13495 6684 15884 6712
rect 13495 6681 13507 6684
rect 13449 6675 13507 6681
rect 11164 6616 11744 6644
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 13081 6647 13139 6653
rect 13081 6644 13093 6647
rect 12860 6616 13093 6644
rect 12860 6604 12866 6616
rect 13081 6613 13093 6616
rect 13127 6613 13139 6647
rect 13081 6607 13139 6613
rect 14090 6604 14096 6656
rect 14148 6644 14154 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 14148 6616 14657 6644
rect 14148 6604 14154 6616
rect 14645 6613 14657 6616
rect 14691 6644 14703 6647
rect 15654 6644 15660 6656
rect 14691 6616 15660 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 15856 6644 15884 6684
rect 17034 6672 17040 6724
rect 17092 6672 17098 6724
rect 17494 6672 17500 6724
rect 17552 6712 17558 6724
rect 18969 6715 19027 6721
rect 18969 6712 18981 6715
rect 17552 6684 18981 6712
rect 17552 6672 17558 6684
rect 18969 6681 18981 6684
rect 19015 6681 19027 6715
rect 19352 6712 19380 6820
rect 19610 6808 19616 6820
rect 19668 6848 19674 6860
rect 20272 6857 20300 6888
rect 20732 6888 21456 6916
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 19668 6820 19809 6848
rect 19668 6808 19674 6820
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 20257 6851 20315 6857
rect 19797 6811 19855 6817
rect 19883 6820 20116 6848
rect 19702 6740 19708 6792
rect 19760 6780 19766 6792
rect 19883 6780 19911 6820
rect 20088 6792 20116 6820
rect 20257 6817 20269 6851
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 19760 6752 19911 6780
rect 19981 6783 20039 6789
rect 19760 6740 19766 6752
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 18969 6675 19027 6681
rect 19076 6684 19380 6712
rect 18233 6647 18291 6653
rect 18233 6644 18245 6647
rect 15856 6616 18245 6644
rect 18233 6613 18245 6616
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 18414 6604 18420 6656
rect 18472 6604 18478 6656
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 19076 6644 19104 6684
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 19996 6712 20024 6743
rect 20070 6740 20076 6792
rect 20128 6740 20134 6792
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 20272 6780 20300 6811
rect 20438 6808 20444 6860
rect 20496 6848 20502 6860
rect 20533 6851 20591 6857
rect 20533 6848 20545 6851
rect 20496 6820 20545 6848
rect 20496 6808 20502 6820
rect 20533 6817 20545 6820
rect 20579 6848 20591 6851
rect 20622 6848 20628 6860
rect 20579 6820 20628 6848
rect 20579 6817 20591 6820
rect 20533 6811 20591 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 20732 6857 20760 6888
rect 21450 6876 21456 6888
rect 21508 6876 21514 6928
rect 21634 6916 21640 6928
rect 21560 6888 21640 6916
rect 21560 6857 21588 6888
rect 21634 6876 21640 6888
rect 21692 6916 21698 6928
rect 22646 6916 22652 6928
rect 21692 6888 22652 6916
rect 21692 6876 21698 6888
rect 22646 6876 22652 6888
rect 22704 6876 22710 6928
rect 20717 6851 20775 6857
rect 20717 6817 20729 6851
rect 20763 6817 20775 6851
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 20717 6811 20775 6817
rect 20824 6820 21373 6848
rect 20824 6780 20852 6820
rect 21361 6817 21373 6820
rect 21407 6817 21419 6851
rect 21361 6811 21419 6817
rect 21545 6851 21603 6857
rect 21545 6817 21557 6851
rect 21591 6817 21603 6851
rect 21545 6811 21603 6817
rect 20272 6752 20852 6780
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 21560 6780 21588 6811
rect 21726 6808 21732 6860
rect 21784 6848 21790 6860
rect 22189 6851 22247 6857
rect 22189 6848 22201 6851
rect 21784 6820 22201 6848
rect 21784 6808 21790 6820
rect 22189 6817 22201 6820
rect 22235 6817 22247 6851
rect 22189 6811 22247 6817
rect 22278 6808 22284 6860
rect 22336 6808 22342 6860
rect 22370 6808 22376 6860
rect 22428 6808 22434 6860
rect 22557 6851 22615 6857
rect 22557 6817 22569 6851
rect 22603 6848 22615 6851
rect 23124 6848 23152 6956
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 23474 6944 23480 6996
rect 23532 6984 23538 6996
rect 24578 6993 24584 6996
rect 23661 6987 23719 6993
rect 23661 6984 23673 6987
rect 23532 6956 23673 6984
rect 23532 6944 23538 6956
rect 23661 6953 23673 6956
rect 23707 6953 23719 6987
rect 24555 6987 24584 6993
rect 23661 6947 23719 6953
rect 23952 6956 24348 6984
rect 23952 6916 23980 6956
rect 22603 6820 23152 6848
rect 23216 6888 23980 6916
rect 24029 6919 24087 6925
rect 22603 6817 22615 6820
rect 22557 6811 22615 6817
rect 21232 6752 21588 6780
rect 21232 6740 21238 6752
rect 21910 6740 21916 6792
rect 21968 6740 21974 6792
rect 22738 6740 22744 6792
rect 22796 6780 22802 6792
rect 23216 6780 23244 6888
rect 24029 6885 24041 6919
rect 24075 6916 24087 6919
rect 24118 6916 24124 6928
rect 24075 6888 24124 6916
rect 24075 6885 24087 6888
rect 24029 6879 24087 6885
rect 24118 6876 24124 6888
rect 24176 6876 24182 6928
rect 23293 6851 23351 6857
rect 23293 6817 23305 6851
rect 23339 6817 23351 6851
rect 23293 6811 23351 6817
rect 23477 6851 23535 6857
rect 23477 6817 23489 6851
rect 23523 6817 23535 6851
rect 23477 6811 23535 6817
rect 23569 6851 23627 6857
rect 23569 6817 23581 6851
rect 23615 6817 23627 6851
rect 23569 6811 23627 6817
rect 22796 6752 23244 6780
rect 23308 6780 23336 6811
rect 23382 6780 23388 6792
rect 23308 6752 23388 6780
rect 22796 6740 22802 6752
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 19668 6684 20024 6712
rect 20441 6715 20499 6721
rect 19668 6672 19674 6684
rect 20441 6681 20453 6715
rect 20487 6712 20499 6715
rect 22830 6712 22836 6724
rect 20487 6684 22836 6712
rect 20487 6681 20499 6684
rect 20441 6675 20499 6681
rect 22830 6672 22836 6684
rect 22888 6672 22894 6724
rect 23014 6672 23020 6724
rect 23072 6712 23078 6724
rect 23492 6712 23520 6811
rect 23584 6780 23612 6811
rect 23658 6808 23664 6860
rect 23716 6848 23722 6860
rect 24320 6857 24348 6956
rect 24555 6953 24567 6987
rect 24555 6947 24584 6953
rect 24578 6944 24584 6947
rect 24636 6944 24642 6996
rect 25406 6944 25412 6996
rect 25464 6984 25470 6996
rect 25501 6987 25559 6993
rect 25501 6984 25513 6987
rect 25464 6956 25513 6984
rect 25464 6944 25470 6956
rect 25501 6953 25513 6956
rect 25547 6953 25559 6987
rect 25501 6947 25559 6953
rect 25774 6944 25780 6996
rect 25832 6984 25838 6996
rect 29822 6984 29828 6996
rect 25832 6956 29828 6984
rect 25832 6944 25838 6956
rect 29822 6944 29828 6956
rect 29880 6944 29886 6996
rect 24762 6876 24768 6928
rect 24820 6876 24826 6928
rect 25424 6916 25452 6944
rect 25240 6888 25452 6916
rect 25685 6919 25743 6925
rect 23845 6851 23903 6857
rect 23845 6848 23857 6851
rect 23716 6820 23857 6848
rect 23716 6808 23722 6820
rect 23845 6817 23857 6820
rect 23891 6817 23903 6851
rect 23845 6811 23903 6817
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6817 23995 6851
rect 23937 6811 23995 6817
rect 24213 6851 24271 6857
rect 24213 6817 24225 6851
rect 24259 6817 24271 6851
rect 24213 6811 24271 6817
rect 24305 6851 24363 6857
rect 24305 6817 24317 6851
rect 24351 6817 24363 6851
rect 24305 6811 24363 6817
rect 23584 6752 23704 6780
rect 23676 6724 23704 6752
rect 23072 6684 23520 6712
rect 23072 6672 23078 6684
rect 23658 6672 23664 6724
rect 23716 6672 23722 6724
rect 23952 6712 23980 6811
rect 24228 6780 24256 6811
rect 24670 6808 24676 6860
rect 24728 6848 24734 6860
rect 25133 6851 25191 6857
rect 25133 6848 25145 6851
rect 24728 6820 25145 6848
rect 24728 6808 24734 6820
rect 25133 6817 25145 6820
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 24946 6780 24952 6792
rect 24228 6752 24952 6780
rect 24946 6740 24952 6752
rect 25004 6740 25010 6792
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6780 25099 6783
rect 25240 6780 25268 6888
rect 25685 6885 25697 6919
rect 25731 6916 25743 6919
rect 26878 6916 26884 6928
rect 25731 6888 26884 6916
rect 25731 6885 25743 6888
rect 25685 6879 25743 6885
rect 25792 6860 25820 6888
rect 26878 6876 26884 6888
rect 26936 6876 26942 6928
rect 27801 6919 27859 6925
rect 27801 6885 27813 6919
rect 27847 6916 27859 6919
rect 28350 6916 28356 6928
rect 27847 6888 28356 6916
rect 27847 6885 27859 6888
rect 27801 6879 27859 6885
rect 28350 6876 28356 6888
rect 28408 6876 28414 6928
rect 28994 6916 29000 6928
rect 28460 6888 29000 6916
rect 25314 6808 25320 6860
rect 25372 6848 25378 6860
rect 25409 6851 25467 6857
rect 25409 6848 25421 6851
rect 25372 6820 25421 6848
rect 25372 6808 25378 6820
rect 25409 6817 25421 6820
rect 25455 6817 25467 6851
rect 25409 6811 25467 6817
rect 25774 6808 25780 6860
rect 25832 6808 25838 6860
rect 25869 6851 25927 6857
rect 25869 6817 25881 6851
rect 25915 6817 25927 6851
rect 25869 6811 25927 6817
rect 25087 6752 25268 6780
rect 25087 6749 25099 6752
rect 25041 6743 25099 6749
rect 25590 6740 25596 6792
rect 25648 6780 25654 6792
rect 25884 6780 25912 6811
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 27525 6851 27583 6857
rect 27525 6848 27537 6851
rect 26384 6820 27537 6848
rect 26384 6808 26390 6820
rect 27525 6817 27537 6820
rect 27571 6848 27583 6851
rect 28460 6848 28488 6888
rect 27571 6820 28488 6848
rect 27571 6817 27583 6820
rect 27525 6811 27583 6817
rect 28534 6808 28540 6860
rect 28592 6808 28598 6860
rect 28626 6808 28632 6860
rect 28684 6808 28690 6860
rect 28828 6857 28856 6888
rect 28994 6876 29000 6888
rect 29052 6876 29058 6928
rect 28813 6851 28871 6857
rect 28813 6817 28825 6851
rect 28859 6817 28871 6851
rect 28813 6811 28871 6817
rect 29454 6808 29460 6860
rect 29512 6808 29518 6860
rect 30098 6808 30104 6860
rect 30156 6808 30162 6860
rect 30561 6851 30619 6857
rect 30561 6817 30573 6851
rect 30607 6848 30619 6851
rect 30650 6848 30656 6860
rect 30607 6820 30656 6848
rect 30607 6817 30619 6820
rect 30561 6811 30619 6817
rect 30650 6808 30656 6820
rect 30708 6808 30714 6860
rect 30834 6808 30840 6860
rect 30892 6848 30898 6860
rect 31018 6848 31024 6860
rect 30892 6820 31024 6848
rect 30892 6808 30898 6820
rect 31018 6808 31024 6820
rect 31076 6848 31082 6860
rect 31113 6851 31171 6857
rect 31113 6848 31125 6851
rect 31076 6820 31125 6848
rect 31076 6808 31082 6820
rect 31113 6817 31125 6820
rect 31159 6817 31171 6851
rect 31113 6811 31171 6817
rect 26142 6780 26148 6792
rect 25648 6752 26148 6780
rect 25648 6740 25654 6752
rect 26142 6740 26148 6752
rect 26200 6740 26206 6792
rect 27338 6740 27344 6792
rect 27396 6780 27402 6792
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 27396 6752 27629 6780
rect 27396 6740 27402 6752
rect 27617 6749 27629 6752
rect 27663 6749 27675 6783
rect 28644 6780 28672 6808
rect 30009 6783 30067 6789
rect 30009 6780 30021 6783
rect 28644 6752 30021 6780
rect 27617 6743 27675 6749
rect 30009 6749 30021 6752
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 24302 6712 24308 6724
rect 23952 6684 24308 6712
rect 24302 6672 24308 6684
rect 24360 6672 24366 6724
rect 24394 6672 24400 6724
rect 24452 6672 24458 6724
rect 27062 6672 27068 6724
rect 27120 6712 27126 6724
rect 27120 6684 27660 6712
rect 27120 6672 27126 6684
rect 18748 6616 19104 6644
rect 18748 6604 18754 6616
rect 19242 6604 19248 6656
rect 19300 6644 19306 6656
rect 20622 6644 20628 6656
rect 19300 6616 20628 6644
rect 19300 6604 19306 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 21361 6647 21419 6653
rect 21361 6644 21373 6647
rect 20772 6616 21373 6644
rect 20772 6604 20778 6616
rect 21361 6613 21373 6616
rect 21407 6613 21419 6647
rect 21361 6607 21419 6613
rect 21726 6604 21732 6656
rect 21784 6604 21790 6656
rect 21910 6604 21916 6656
rect 21968 6644 21974 6656
rect 22094 6644 22100 6656
rect 21968 6616 22100 6644
rect 21968 6604 21974 6616
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 23198 6604 23204 6656
rect 23256 6644 23262 6656
rect 23293 6647 23351 6653
rect 23293 6644 23305 6647
rect 23256 6616 23305 6644
rect 23256 6604 23262 6616
rect 23293 6613 23305 6616
rect 23339 6613 23351 6647
rect 23293 6607 23351 6613
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 24578 6644 24584 6656
rect 23440 6616 24584 6644
rect 23440 6604 23446 6616
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 24949 6647 25007 6653
rect 24949 6644 24961 6647
rect 24912 6616 24961 6644
rect 24912 6604 24918 6616
rect 24949 6613 24961 6616
rect 24995 6613 25007 6647
rect 24949 6607 25007 6613
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 25280 6616 25329 6644
rect 25280 6604 25286 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 25317 6607 25375 6613
rect 25590 6604 25596 6656
rect 25648 6644 25654 6656
rect 27632 6653 27660 6684
rect 28166 6672 28172 6724
rect 28224 6712 28230 6724
rect 28902 6712 28908 6724
rect 28224 6684 28908 6712
rect 28224 6672 28230 6684
rect 28902 6672 28908 6684
rect 28960 6712 28966 6724
rect 29181 6715 29239 6721
rect 29181 6712 29193 6715
rect 28960 6684 29193 6712
rect 28960 6672 28966 6684
rect 29181 6681 29193 6684
rect 29227 6681 29239 6715
rect 29181 6675 29239 6681
rect 27341 6647 27399 6653
rect 27341 6644 27353 6647
rect 25648 6616 27353 6644
rect 25648 6604 25654 6616
rect 27341 6613 27353 6616
rect 27387 6613 27399 6647
rect 27341 6607 27399 6613
rect 27617 6647 27675 6653
rect 27617 6613 27629 6647
rect 27663 6613 27675 6647
rect 27617 6607 27675 6613
rect 28994 6604 29000 6656
rect 29052 6604 29058 6656
rect 552 6554 31648 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 11436 6554
rect 11488 6502 11500 6554
rect 11552 6502 11564 6554
rect 11616 6502 11628 6554
rect 11680 6502 11692 6554
rect 11744 6502 19210 6554
rect 19262 6502 19274 6554
rect 19326 6502 19338 6554
rect 19390 6502 19402 6554
rect 19454 6502 19466 6554
rect 19518 6502 26984 6554
rect 27036 6502 27048 6554
rect 27100 6502 27112 6554
rect 27164 6502 27176 6554
rect 27228 6502 27240 6554
rect 27292 6502 31648 6554
rect 552 6480 31648 6502
rect 1762 6400 1768 6452
rect 1820 6400 1826 6452
rect 2866 6400 2872 6452
rect 2924 6400 2930 6452
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 6641 6443 6699 6449
rect 6641 6440 6653 6443
rect 3007 6412 6653 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 6641 6409 6653 6412
rect 6687 6409 6699 6443
rect 6641 6403 6699 6409
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 8018 6440 8024 6452
rect 7147 6412 8024 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 10134 6440 10140 6452
rect 8352 6412 10140 6440
rect 8352 6400 8358 6412
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 1946 6332 1952 6384
rect 2004 6372 2010 6384
rect 4249 6375 4307 6381
rect 2004 6344 3372 6372
rect 2004 6332 2010 6344
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1670 6304 1676 6316
rect 1443 6276 1676 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1670 6264 1676 6276
rect 1728 6304 1734 6316
rect 1728 6276 3004 6304
rect 1728 6264 1734 6276
rect 1578 6196 1584 6248
rect 1636 6196 1642 6248
rect 2774 6196 2780 6248
rect 2832 6196 2838 6248
rect 2976 6236 3004 6276
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 3344 6304 3372 6344
rect 4249 6341 4261 6375
rect 4295 6372 4307 6375
rect 10612 6372 10640 6403
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11698 6440 11704 6452
rect 11112 6412 11704 6440
rect 11112 6400 11118 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 14369 6443 14427 6449
rect 11848 6412 13952 6440
rect 11848 6400 11854 6412
rect 13722 6372 13728 6384
rect 4295 6344 13728 6372
rect 4295 6341 4307 6344
rect 4249 6335 4307 6341
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 13924 6372 13952 6412
rect 14369 6409 14381 6443
rect 14415 6440 14427 6443
rect 15286 6440 15292 6452
rect 14415 6412 15292 6440
rect 14415 6409 14427 6412
rect 14369 6403 14427 6409
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 15436 6412 15485 6440
rect 15436 6400 15442 6412
rect 15473 6409 15485 6412
rect 15519 6409 15531 6443
rect 15473 6403 15531 6409
rect 16114 6400 16120 6452
rect 16172 6400 16178 6452
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17954 6440 17960 6452
rect 17460 6412 17960 6440
rect 17460 6400 17466 6412
rect 17954 6400 17960 6412
rect 18012 6440 18018 6452
rect 18322 6440 18328 6452
rect 18012 6412 18328 6440
rect 18012 6400 18018 6412
rect 18322 6400 18328 6412
rect 18380 6440 18386 6452
rect 19794 6440 19800 6452
rect 18380 6412 19800 6440
rect 18380 6400 18386 6412
rect 19794 6400 19800 6412
rect 19852 6440 19858 6452
rect 20438 6440 20444 6452
rect 19852 6412 20444 6440
rect 19852 6400 19858 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 22002 6440 22008 6452
rect 20680 6412 22008 6440
rect 20680 6400 20686 6412
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 22097 6443 22155 6449
rect 22097 6409 22109 6443
rect 22143 6440 22155 6443
rect 22278 6440 22284 6452
rect 22143 6412 22284 6440
rect 22143 6409 22155 6412
rect 22097 6403 22155 6409
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 24026 6400 24032 6452
rect 24084 6400 24090 6452
rect 24397 6443 24455 6449
rect 24397 6409 24409 6443
rect 24443 6440 24455 6443
rect 24578 6440 24584 6452
rect 24443 6412 24584 6440
rect 24443 6409 24455 6412
rect 24397 6403 24455 6409
rect 24578 6400 24584 6412
rect 24636 6400 24642 6452
rect 24854 6400 24860 6452
rect 24912 6440 24918 6452
rect 25133 6443 25191 6449
rect 25133 6440 25145 6443
rect 24912 6412 25145 6440
rect 24912 6400 24918 6412
rect 25133 6409 25145 6412
rect 25179 6409 25191 6443
rect 25133 6403 25191 6409
rect 25501 6443 25559 6449
rect 25501 6409 25513 6443
rect 25547 6440 25559 6443
rect 25866 6440 25872 6452
rect 25547 6412 25872 6440
rect 25547 6409 25559 6412
rect 25501 6403 25559 6409
rect 25866 6400 25872 6412
rect 25924 6400 25930 6452
rect 27338 6400 27344 6452
rect 27396 6400 27402 6452
rect 28258 6400 28264 6452
rect 28316 6440 28322 6452
rect 30377 6443 30435 6449
rect 30377 6440 30389 6443
rect 28316 6412 30389 6440
rect 28316 6400 28322 6412
rect 30377 6409 30389 6412
rect 30423 6409 30435 6443
rect 30377 6403 30435 6409
rect 13924 6344 15056 6372
rect 5350 6304 5356 6316
rect 3344 6276 5356 6304
rect 3344 6248 3372 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 6638 6304 6644 6316
rect 5460 6276 6644 6304
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 2976 6208 3249 6236
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3252 6168 3280 6199
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 3384 6208 3525 6236
rect 3384 6196 3390 6208
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3660 6208 3709 6236
rect 3660 6196 3666 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 3927 6208 4108 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 3970 6168 3976 6180
rect 3252 6140 3976 6168
rect 3970 6128 3976 6140
rect 4028 6128 4034 6180
rect 4080 6177 4108 6208
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 4672 6208 5273 6236
rect 4672 6196 4678 6208
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 5460 6236 5488 6276
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6779 6276 7205 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 8720 6276 12434 6304
rect 8720 6264 8726 6276
rect 5307 6208 5488 6236
rect 5537 6239 5595 6245
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 6546 6236 6552 6248
rect 5583 6208 6552 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6228 6975 6239
rect 7024 6228 7236 6230
rect 6963 6205 7236 6228
rect 6917 6202 7236 6205
rect 6917 6200 7052 6202
rect 6917 6199 6975 6200
rect 4065 6171 4123 6177
rect 4065 6137 4077 6171
rect 4111 6168 4123 6171
rect 4982 6168 4988 6180
rect 4111 6140 4988 6168
rect 4111 6137 4123 6140
rect 4065 6131 4123 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 5491 6140 5948 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6100 5135 6103
rect 5166 6100 5172 6112
rect 5123 6072 5172 6100
rect 5123 6069 5135 6072
rect 5077 6063 5135 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 5810 6100 5816 6112
rect 5767 6072 5816 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 5920 6100 5948 6140
rect 5994 6128 6000 6180
rect 6052 6128 6058 6180
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 6641 6171 6699 6177
rect 6641 6168 6653 6171
rect 6328 6140 6653 6168
rect 6328 6128 6334 6140
rect 6641 6137 6653 6140
rect 6687 6137 6699 6171
rect 7208 6168 7236 6202
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7340 6208 7389 6236
rect 7340 6196 7346 6208
rect 7377 6205 7389 6208
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 7650 6196 7656 6248
rect 7708 6196 7714 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8018 6236 8024 6248
rect 7883 6208 8024 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 10226 6196 10232 6248
rect 10284 6196 10290 6248
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 10502 6236 10508 6248
rect 10367 6208 10508 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 11974 6236 11980 6248
rect 10744 6208 11980 6236
rect 10744 6196 10750 6208
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12406 6236 12434 6276
rect 12802 6264 12808 6316
rect 12860 6264 12866 6316
rect 12894 6264 12900 6316
rect 12952 6264 12958 6316
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12406 6208 12633 6236
rect 12621 6205 12633 6208
rect 12667 6236 12679 6239
rect 12986 6236 12992 6248
rect 12667 6208 12992 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 13078 6196 13084 6248
rect 13136 6196 13142 6248
rect 13265 6239 13323 6245
rect 13265 6205 13277 6239
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 12437 6171 12495 6177
rect 12437 6168 12449 6171
rect 7208 6140 12449 6168
rect 6641 6131 6699 6137
rect 12437 6137 12449 6140
rect 12483 6137 12495 6171
rect 12437 6131 12495 6137
rect 12710 6128 12716 6180
rect 12768 6168 12774 6180
rect 13280 6168 13308 6199
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13924 6245 13952 6344
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14200 6276 14473 6304
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13504 6208 13829 6236
rect 13504 6196 13510 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 14090 6196 14096 6248
rect 14148 6196 14154 6248
rect 14200 6245 14228 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14826 6304 14832 6316
rect 14461 6267 14519 6273
rect 14560 6276 14832 6304
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 14560 6236 14588 6276
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 15028 6304 15056 6344
rect 18230 6332 18236 6384
rect 18288 6372 18294 6384
rect 22554 6372 22560 6384
rect 18288 6344 22560 6372
rect 18288 6332 18294 6344
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 23474 6332 23480 6384
rect 23532 6372 23538 6384
rect 24762 6372 24768 6384
rect 23532 6344 24768 6372
rect 23532 6332 23538 6344
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 25774 6372 25780 6384
rect 24872 6344 25780 6372
rect 24394 6304 24400 6316
rect 15028 6276 24400 6304
rect 24394 6264 24400 6276
rect 24452 6264 24458 6316
rect 14332 6208 14588 6236
rect 14332 6196 14338 6208
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 14734 6196 14740 6248
rect 14792 6196 14798 6248
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6236 14979 6239
rect 15010 6236 15016 6248
rect 14967 6208 15016 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15010 6196 15016 6208
rect 15068 6196 15074 6248
rect 15194 6196 15200 6248
rect 15252 6236 15258 6248
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 15252 6208 15301 6236
rect 15252 6196 15258 6208
rect 15289 6205 15301 6208
rect 15335 6236 15347 6239
rect 16114 6236 16120 6248
rect 15335 6208 16120 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 16390 6236 16396 6248
rect 16347 6208 16396 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16482 6196 16488 6248
rect 16540 6196 16546 6248
rect 16574 6196 16580 6248
rect 16632 6196 16638 6248
rect 19150 6236 19156 6248
rect 18432 6208 19156 6236
rect 12768 6140 13308 6168
rect 14660 6168 14688 6196
rect 15105 6171 15163 6177
rect 15105 6168 15117 6171
rect 14660 6140 15117 6168
rect 12768 6128 12774 6140
rect 15105 6137 15117 6140
rect 15151 6137 15163 6171
rect 15105 6131 15163 6137
rect 15378 6128 15384 6180
rect 15436 6168 15442 6180
rect 16758 6168 16764 6180
rect 15436 6140 16764 6168
rect 15436 6128 15442 6140
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 10318 6100 10324 6112
rect 5920 6072 10324 6100
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6100 10471 6103
rect 10594 6100 10600 6112
rect 10459 6072 10600 6100
rect 10459 6069 10471 6072
rect 10413 6063 10471 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 11146 6100 11152 6112
rect 10735 6072 11152 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11514 6100 11520 6112
rect 11296 6072 11520 6100
rect 11296 6060 11302 6072
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12986 6100 12992 6112
rect 11848 6072 12992 6100
rect 11848 6060 11854 6072
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13262 6060 13268 6112
rect 13320 6060 13326 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 18432 6100 18460 6208
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19245 6239 19303 6245
rect 19245 6205 19257 6239
rect 19291 6205 19303 6239
rect 19245 6199 19303 6205
rect 18506 6128 18512 6180
rect 18564 6168 18570 6180
rect 18782 6168 18788 6180
rect 18564 6140 18788 6168
rect 18564 6128 18570 6140
rect 18782 6128 18788 6140
rect 18840 6168 18846 6180
rect 19260 6168 19288 6199
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19484 6208 19533 6236
rect 19484 6196 19490 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 21266 6196 21272 6248
rect 21324 6236 21330 6248
rect 21910 6236 21916 6248
rect 21324 6208 21916 6236
rect 21324 6196 21330 6208
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6205 22155 6239
rect 22097 6199 22155 6205
rect 20070 6168 20076 6180
rect 18840 6140 19288 6168
rect 19352 6140 20076 6168
rect 18840 6128 18846 6140
rect 13780 6072 18460 6100
rect 13780 6060 13786 6072
rect 18874 6060 18880 6112
rect 18932 6100 18938 6112
rect 19061 6103 19119 6109
rect 19061 6100 19073 6103
rect 18932 6072 19073 6100
rect 18932 6060 18938 6072
rect 19061 6069 19073 6072
rect 19107 6069 19119 6103
rect 19061 6063 19119 6069
rect 19150 6060 19156 6112
rect 19208 6100 19214 6112
rect 19352 6100 19380 6140
rect 20070 6128 20076 6140
rect 20128 6128 20134 6180
rect 21082 6128 21088 6180
rect 21140 6168 21146 6180
rect 22112 6168 22140 6199
rect 23750 6196 23756 6248
rect 23808 6236 23814 6248
rect 24305 6239 24363 6245
rect 24305 6236 24317 6239
rect 23808 6208 24317 6236
rect 23808 6196 23814 6208
rect 24305 6205 24317 6208
rect 24351 6205 24363 6239
rect 24305 6199 24363 6205
rect 24489 6239 24547 6245
rect 24489 6205 24501 6239
rect 24535 6236 24547 6239
rect 24872 6236 24900 6344
rect 25774 6332 25780 6344
rect 25832 6332 25838 6384
rect 26142 6332 26148 6384
rect 26200 6372 26206 6384
rect 30650 6372 30656 6384
rect 26200 6344 30656 6372
rect 26200 6332 26206 6344
rect 30650 6332 30656 6344
rect 30708 6332 30714 6384
rect 26602 6304 26608 6316
rect 25240 6276 26608 6304
rect 25240 6245 25268 6276
rect 26602 6264 26608 6276
rect 26660 6304 26666 6316
rect 26660 6276 27384 6304
rect 26660 6264 26666 6276
rect 24535 6208 24900 6236
rect 25041 6239 25099 6245
rect 24535 6205 24547 6208
rect 24489 6199 24547 6205
rect 25041 6205 25053 6239
rect 25087 6205 25099 6239
rect 25041 6199 25099 6205
rect 25225 6239 25283 6245
rect 25225 6205 25237 6239
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 21140 6140 22140 6168
rect 21140 6128 21146 6140
rect 24210 6128 24216 6180
rect 24268 6128 24274 6180
rect 24320 6168 24348 6199
rect 24670 6168 24676 6180
rect 24320 6140 24676 6168
rect 24670 6128 24676 6140
rect 24728 6128 24734 6180
rect 25056 6168 25084 6199
rect 25314 6196 25320 6248
rect 25372 6236 25378 6248
rect 25685 6239 25743 6245
rect 25685 6236 25697 6239
rect 25372 6208 25697 6236
rect 25372 6196 25378 6208
rect 25685 6205 25697 6208
rect 25731 6205 25743 6239
rect 25685 6199 25743 6205
rect 25774 6196 25780 6248
rect 25832 6196 25838 6248
rect 26878 6196 26884 6248
rect 26936 6236 26942 6248
rect 27356 6245 27384 6276
rect 28994 6264 29000 6316
rect 29052 6264 29058 6316
rect 29549 6307 29607 6313
rect 29104 6276 29316 6304
rect 27157 6239 27215 6245
rect 27157 6236 27169 6239
rect 26936 6208 27169 6236
rect 26936 6196 26942 6208
rect 27157 6205 27169 6208
rect 27203 6205 27215 6239
rect 27157 6199 27215 6205
rect 27341 6239 27399 6245
rect 27341 6205 27353 6239
rect 27387 6205 27399 6239
rect 27341 6199 27399 6205
rect 28442 6196 28448 6248
rect 28500 6236 28506 6248
rect 29104 6236 29132 6276
rect 28500 6208 29132 6236
rect 28500 6196 28506 6208
rect 29178 6196 29184 6248
rect 29236 6196 29242 6248
rect 29288 6236 29316 6276
rect 29549 6273 29561 6307
rect 29595 6304 29607 6307
rect 29641 6307 29699 6313
rect 29641 6304 29653 6307
rect 29595 6276 29653 6304
rect 29595 6273 29607 6276
rect 29549 6267 29607 6273
rect 29641 6273 29653 6276
rect 29687 6273 29699 6307
rect 29641 6267 29699 6273
rect 29822 6264 29828 6316
rect 29880 6264 29886 6316
rect 30006 6264 30012 6316
rect 30064 6264 30070 6316
rect 30098 6264 30104 6316
rect 30156 6264 30162 6316
rect 29917 6239 29975 6245
rect 29917 6236 29929 6239
rect 29288 6208 29929 6236
rect 29917 6205 29929 6208
rect 29963 6205 29975 6239
rect 29917 6199 29975 6205
rect 25406 6168 25412 6180
rect 25056 6140 25412 6168
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 26970 6128 26976 6180
rect 27028 6168 27034 6180
rect 30116 6168 30144 6264
rect 30282 6196 30288 6248
rect 30340 6196 30346 6248
rect 30469 6239 30527 6245
rect 30469 6236 30481 6239
rect 30392 6208 30481 6236
rect 27028 6140 30144 6168
rect 27028 6128 27034 6140
rect 19208 6072 19380 6100
rect 19429 6103 19487 6109
rect 19208 6060 19214 6072
rect 19429 6069 19441 6103
rect 19475 6100 19487 6103
rect 20162 6100 20168 6112
rect 19475 6072 20168 6100
rect 19475 6069 19487 6072
rect 19429 6063 19487 6069
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 22738 6100 22744 6112
rect 20312 6072 22744 6100
rect 20312 6060 20318 6072
rect 22738 6060 22744 6072
rect 22796 6060 22802 6112
rect 23842 6060 23848 6112
rect 23900 6060 23906 6112
rect 24026 6109 24032 6112
rect 24013 6103 24032 6109
rect 24013 6069 24025 6103
rect 24013 6063 24032 6069
rect 24026 6060 24032 6063
rect 24084 6060 24090 6112
rect 28994 6060 29000 6112
rect 29052 6100 29058 6112
rect 29181 6103 29239 6109
rect 29181 6100 29193 6103
rect 29052 6072 29193 6100
rect 29052 6060 29058 6072
rect 29181 6069 29193 6072
rect 29227 6069 29239 6103
rect 29181 6063 29239 6069
rect 30006 6060 30012 6112
rect 30064 6100 30070 6112
rect 30392 6100 30420 6208
rect 30469 6205 30481 6208
rect 30515 6205 30527 6239
rect 30469 6199 30527 6205
rect 30064 6072 30420 6100
rect 30064 6060 30070 6072
rect 552 6010 31648 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 12096 6010
rect 12148 5958 12160 6010
rect 12212 5958 12224 6010
rect 12276 5958 12288 6010
rect 12340 5958 12352 6010
rect 12404 5958 19870 6010
rect 19922 5958 19934 6010
rect 19986 5958 19998 6010
rect 20050 5958 20062 6010
rect 20114 5958 20126 6010
rect 20178 5958 27644 6010
rect 27696 5958 27708 6010
rect 27760 5958 27772 6010
rect 27824 5958 27836 6010
rect 27888 5958 27900 6010
rect 27952 5958 31648 6010
rect 552 5936 31648 5958
rect 934 5856 940 5908
rect 992 5896 998 5908
rect 1397 5899 1455 5905
rect 1397 5896 1409 5899
rect 992 5868 1409 5896
rect 992 5856 998 5868
rect 1397 5865 1409 5868
rect 1443 5896 1455 5899
rect 4617 5899 4675 5905
rect 1443 5868 4384 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 1946 5788 1952 5840
rect 2004 5788 2010 5840
rect 2130 5788 2136 5840
rect 2188 5828 2194 5840
rect 2317 5831 2375 5837
rect 2317 5828 2329 5831
rect 2188 5800 2329 5828
rect 2188 5788 2194 5800
rect 2317 5797 2329 5800
rect 2363 5828 2375 5831
rect 3510 5828 3516 5840
rect 2363 5800 3516 5828
rect 2363 5797 2375 5800
rect 2317 5791 2375 5797
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 4062 5828 4068 5840
rect 3988 5800 4068 5828
rect 1302 5720 1308 5772
rect 1360 5720 1366 5772
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5729 1547 5763
rect 1489 5723 1547 5729
rect 1504 5624 1532 5723
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1728 5732 1869 5760
rect 1728 5720 1734 5732
rect 1857 5729 1869 5732
rect 1903 5729 1915 5763
rect 3050 5760 3056 5772
rect 1857 5723 1915 5729
rect 2056 5732 3056 5760
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 2056 5701 2084 5732
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 3988 5769 4016 5800
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 3292 5732 3341 5760
rect 3292 5720 3298 5732
rect 3329 5729 3341 5732
rect 3375 5729 3387 5763
rect 3329 5723 3387 5729
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5729 4031 5763
rect 3973 5723 4031 5729
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1636 5664 2053 5692
rect 1636 5652 1642 5664
rect 2041 5661 2053 5664
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 3252 5692 3280 5720
rect 2280 5664 3280 5692
rect 2280 5652 2286 5664
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3476 5664 4077 5692
rect 3476 5652 3482 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4356 5692 4384 5868
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 4706 5896 4712 5908
rect 4663 5868 4712 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5865 4859 5899
rect 4801 5859 4859 5865
rect 4816 5828 4844 5859
rect 6270 5856 6276 5908
rect 6328 5856 6334 5908
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 7282 5896 7288 5908
rect 6696 5868 7288 5896
rect 6696 5856 6702 5868
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7558 5896 7564 5908
rect 7432 5868 7564 5896
rect 7432 5856 7438 5868
rect 7558 5856 7564 5868
rect 7616 5896 7622 5908
rect 7616 5868 8294 5896
rect 7616 5856 7622 5868
rect 5810 5828 5816 5840
rect 4816 5800 5816 5828
rect 5810 5788 5816 5800
rect 5868 5828 5874 5840
rect 5868 5800 6408 5828
rect 5868 5788 5874 5800
rect 4798 5760 4804 5772
rect 4759 5732 4804 5760
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 5166 5720 5172 5772
rect 5224 5720 5230 5772
rect 5258 5720 5264 5772
rect 5316 5720 5322 5772
rect 6270 5720 6276 5772
rect 6328 5720 6334 5772
rect 6380 5769 6408 5800
rect 6546 5788 6552 5840
rect 6604 5788 6610 5840
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 7742 5828 7748 5840
rect 7064 5800 7748 5828
rect 7064 5788 7070 5800
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 8266 5828 8294 5868
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8628 5868 8861 5896
rect 8628 5856 8634 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 9456 5868 9689 5896
rect 9456 5856 9462 5868
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 11882 5896 11888 5908
rect 9677 5859 9735 5865
rect 11256 5868 11888 5896
rect 8757 5831 8815 5837
rect 8757 5828 8769 5831
rect 8266 5800 8769 5828
rect 8757 5797 8769 5800
rect 8803 5828 8815 5831
rect 9125 5831 9183 5837
rect 9125 5828 9137 5831
rect 8803 5800 9137 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9125 5797 9137 5800
rect 9171 5797 9183 5831
rect 9125 5791 9183 5797
rect 9214 5788 9220 5840
rect 9272 5828 9278 5840
rect 10134 5828 10140 5840
rect 9272 5800 10140 5828
rect 9272 5788 9278 5800
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 10318 5788 10324 5840
rect 10376 5828 10382 5840
rect 11256 5828 11284 5868
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 13446 5896 13452 5908
rect 12032 5868 13452 5896
rect 12032 5856 12038 5868
rect 13446 5856 13452 5868
rect 13504 5856 13510 5908
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 13722 5896 13728 5908
rect 13596 5868 13728 5896
rect 13596 5856 13602 5868
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 15286 5896 15292 5908
rect 13964 5868 15292 5896
rect 13964 5856 13970 5868
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 17405 5899 17463 5905
rect 17405 5896 17417 5899
rect 16540 5868 17417 5896
rect 16540 5856 16546 5868
rect 17405 5865 17417 5868
rect 17451 5865 17463 5899
rect 17405 5859 17463 5865
rect 18230 5856 18236 5908
rect 18288 5856 18294 5908
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 19058 5896 19064 5908
rect 18371 5868 19064 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5865 19303 5899
rect 20257 5899 20315 5905
rect 20257 5896 20269 5899
rect 19245 5859 19303 5865
rect 19444 5868 20269 5896
rect 10376 5800 11284 5828
rect 10376 5788 10382 5800
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 7558 5720 7564 5772
rect 7616 5720 7622 5772
rect 7760 5760 7788 5788
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 7760 5732 8493 5760
rect 8481 5729 8493 5732
rect 8527 5729 8539 5763
rect 8481 5723 8539 5729
rect 8570 5720 8576 5772
rect 8628 5720 8634 5772
rect 9028 5763 9086 5769
rect 9028 5729 9040 5763
rect 9074 5760 9086 5763
rect 9306 5760 9312 5772
rect 9074 5732 9312 5760
rect 9074 5729 9086 5732
rect 9028 5723 9086 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9398 5720 9404 5772
rect 9456 5720 9462 5772
rect 9490 5720 9496 5772
rect 9548 5720 9554 5772
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5760 9643 5763
rect 9766 5760 9772 5772
rect 9631 5732 9772 5760
rect 9631 5729 9643 5732
rect 9585 5723 9643 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5760 10011 5763
rect 10594 5760 10600 5772
rect 9999 5732 10600 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 11146 5760 11152 5772
rect 11072 5732 11152 5760
rect 6638 5692 6644 5704
rect 4356 5664 6644 5692
rect 4065 5655 4123 5661
rect 6638 5652 6644 5664
rect 6696 5692 6702 5704
rect 7098 5692 7104 5704
rect 6696 5664 7104 5692
rect 6696 5652 6702 5664
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7800 5664 7849 5692
rect 7800 5652 7806 5664
rect 7837 5661 7849 5664
rect 7883 5692 7895 5695
rect 7883 5664 9628 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 2498 5624 2504 5636
rect 1504 5596 2504 5624
rect 2498 5584 2504 5596
rect 2556 5584 2562 5636
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 8757 5627 8815 5633
rect 4387 5596 8616 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 8588 5568 8616 5596
rect 8757 5593 8769 5627
rect 8803 5624 8815 5627
rect 9214 5624 9220 5636
rect 8803 5596 9220 5624
rect 8803 5593 8815 5596
rect 8757 5587 8815 5593
rect 9214 5584 9220 5596
rect 9272 5584 9278 5636
rect 9600 5624 9628 5664
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9732 5664 10149 5692
rect 9732 5652 9738 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10778 5692 10784 5704
rect 10137 5655 10195 5661
rect 10612 5664 10784 5692
rect 10612 5624 10640 5664
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 11072 5692 11100 5732
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11256 5769 11284 5800
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 11609 5831 11667 5837
rect 11609 5828 11621 5831
rect 11388 5800 11621 5828
rect 11388 5788 11394 5800
rect 11609 5797 11621 5800
rect 11655 5797 11667 5831
rect 11609 5791 11667 5797
rect 11793 5831 11851 5837
rect 11793 5797 11805 5831
rect 11839 5828 11851 5831
rect 12066 5828 12072 5840
rect 11839 5800 12072 5828
rect 11839 5797 11851 5800
rect 11793 5791 11851 5797
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 13262 5828 13268 5840
rect 12492 5800 13268 5828
rect 12492 5788 12498 5800
rect 13262 5788 13268 5800
rect 13320 5828 13326 5840
rect 15378 5828 15384 5840
rect 13320 5800 15384 5828
rect 13320 5788 13326 5800
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 18248 5828 18276 5856
rect 16408 5800 18276 5828
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 11422 5720 11428 5772
rect 11480 5720 11486 5772
rect 11514 5720 11520 5772
rect 11572 5720 11578 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 16408 5760 16436 5800
rect 18598 5788 18604 5840
rect 18656 5828 18662 5840
rect 19260 5828 19288 5859
rect 18656 5800 19288 5828
rect 18656 5788 18662 5800
rect 11756 5732 16436 5760
rect 11756 5720 11762 5732
rect 16482 5720 16488 5772
rect 16540 5720 16546 5772
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 16761 5763 16819 5769
rect 16761 5729 16773 5763
rect 16807 5760 16819 5763
rect 16850 5760 16856 5772
rect 16807 5732 16856 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11072 5664 11989 5692
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 15746 5692 15752 5704
rect 12124 5664 15752 5692
rect 12124 5652 12130 5664
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 11790 5624 11796 5636
rect 9600 5596 10640 5624
rect 10704 5596 11796 5624
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9030 5556 9036 5568
rect 8628 5528 9036 5556
rect 8628 5516 8634 5528
rect 9030 5516 9036 5528
rect 9088 5556 9094 5568
rect 10704 5556 10732 5596
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 14550 5624 14556 5636
rect 12268 5596 14556 5624
rect 9088 5528 10732 5556
rect 9088 5516 9094 5528
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 12268 5556 12296 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 15654 5584 15660 5636
rect 15712 5624 15718 5636
rect 16684 5624 16712 5723
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 17604 5692 17632 5723
rect 17678 5720 17684 5772
rect 17736 5720 17742 5772
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 18012 5732 18245 5760
rect 18012 5720 18018 5732
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5729 18475 5763
rect 18417 5723 18475 5729
rect 17770 5692 17776 5704
rect 17604 5664 17776 5692
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5692 17923 5695
rect 18432 5692 18460 5723
rect 18506 5720 18512 5772
rect 18564 5720 18570 5772
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 18966 5760 18972 5772
rect 18739 5732 18972 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 18966 5720 18972 5732
rect 19024 5760 19030 5772
rect 19444 5760 19472 5868
rect 20257 5865 20269 5868
rect 20303 5896 20315 5899
rect 21174 5896 21180 5908
rect 20303 5868 21180 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 21174 5856 21180 5868
rect 21232 5856 21238 5908
rect 21358 5856 21364 5908
rect 21416 5856 21422 5908
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 23753 5899 23811 5905
rect 23753 5896 23765 5899
rect 21692 5868 23765 5896
rect 21692 5856 21698 5868
rect 23753 5865 23765 5868
rect 23799 5896 23811 5899
rect 24486 5896 24492 5908
rect 23799 5868 24492 5896
rect 23799 5865 23811 5868
rect 23753 5859 23811 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 25314 5856 25320 5908
rect 25372 5896 25378 5908
rect 27065 5899 27123 5905
rect 27065 5896 27077 5899
rect 25372 5868 27077 5896
rect 25372 5856 25378 5868
rect 27065 5865 27077 5868
rect 27111 5896 27123 5899
rect 27430 5896 27436 5908
rect 27111 5868 27436 5896
rect 27111 5865 27123 5868
rect 27065 5859 27123 5865
rect 27430 5856 27436 5868
rect 27488 5856 27494 5908
rect 28442 5856 28448 5908
rect 28500 5896 28506 5908
rect 28905 5899 28963 5905
rect 28905 5896 28917 5899
rect 28500 5868 28917 5896
rect 28500 5856 28506 5868
rect 28905 5865 28917 5868
rect 28951 5865 28963 5899
rect 28905 5859 28963 5865
rect 29178 5856 29184 5908
rect 29236 5896 29242 5908
rect 29641 5899 29699 5905
rect 29641 5896 29653 5899
rect 29236 5868 29653 5896
rect 29236 5856 29242 5868
rect 29641 5865 29653 5868
rect 29687 5865 29699 5899
rect 29641 5859 29699 5865
rect 26605 5831 26663 5837
rect 26605 5828 26617 5831
rect 19536 5800 26617 5828
rect 19536 5769 19564 5800
rect 26605 5797 26617 5800
rect 26651 5797 26663 5831
rect 26970 5828 26976 5840
rect 26605 5791 26663 5797
rect 26712 5800 26976 5828
rect 19024 5732 19472 5760
rect 19521 5763 19579 5769
rect 19024 5720 19030 5732
rect 19521 5729 19533 5763
rect 19567 5729 19579 5763
rect 19521 5723 19579 5729
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 19889 5763 19947 5769
rect 19889 5760 19901 5763
rect 19843 5732 19901 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 19889 5729 19901 5732
rect 19935 5729 19947 5763
rect 19889 5723 19947 5729
rect 20070 5720 20076 5772
rect 20128 5720 20134 5772
rect 20346 5720 20352 5772
rect 20404 5720 20410 5772
rect 21542 5720 21548 5772
rect 21600 5720 21606 5772
rect 21818 5720 21824 5772
rect 21876 5720 21882 5772
rect 22002 5720 22008 5772
rect 22060 5720 22066 5772
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 18601 5695 18659 5701
rect 18601 5692 18613 5695
rect 17911 5664 18613 5692
rect 17911 5661 17923 5664
rect 17865 5655 17923 5661
rect 18601 5661 18613 5664
rect 18647 5661 18659 5695
rect 19334 5692 19340 5704
rect 18601 5655 18659 5661
rect 18708 5664 19340 5692
rect 15712 5596 16712 5624
rect 17788 5624 17816 5652
rect 18708 5624 18736 5664
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 21266 5692 21272 5704
rect 19484 5664 21272 5692
rect 19484 5652 19490 5664
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21637 5695 21695 5701
rect 21637 5661 21649 5695
rect 21683 5692 21695 5695
rect 22097 5695 22155 5701
rect 22097 5692 22109 5695
rect 21683 5664 22109 5692
rect 21683 5661 21695 5664
rect 21637 5655 21695 5661
rect 22097 5661 22109 5664
rect 22143 5661 22155 5695
rect 22204 5692 22232 5723
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 22373 5763 22431 5769
rect 22373 5760 22385 5763
rect 22336 5732 22385 5760
rect 22336 5720 22342 5732
rect 22373 5729 22385 5732
rect 22419 5729 22431 5763
rect 22373 5723 22431 5729
rect 22557 5763 22615 5769
rect 22557 5729 22569 5763
rect 22603 5729 22615 5763
rect 22557 5723 22615 5729
rect 24121 5763 24179 5769
rect 24121 5729 24133 5763
rect 24167 5760 24179 5763
rect 24762 5760 24768 5772
rect 24167 5732 24768 5760
rect 24167 5729 24179 5732
rect 24121 5723 24179 5729
rect 22204 5664 22508 5692
rect 22097 5655 22155 5661
rect 17788 5596 18736 5624
rect 15712 5584 15718 5596
rect 19058 5584 19064 5636
rect 19116 5624 19122 5636
rect 19116 5596 19472 5624
rect 19116 5584 19122 5596
rect 10836 5528 12296 5556
rect 10836 5516 10842 5528
rect 12342 5516 12348 5568
rect 12400 5556 12406 5568
rect 19444 5565 19472 5596
rect 21726 5584 21732 5636
rect 21784 5584 21790 5636
rect 22480 5568 22508 5664
rect 22572 5624 22600 5723
rect 24762 5720 24768 5732
rect 24820 5720 24826 5772
rect 25501 5763 25559 5769
rect 25501 5729 25513 5763
rect 25547 5729 25559 5763
rect 25501 5723 25559 5729
rect 24026 5652 24032 5704
rect 24084 5692 24090 5704
rect 25314 5692 25320 5704
rect 24084 5664 25320 5692
rect 24084 5652 24090 5664
rect 25314 5652 25320 5664
rect 25372 5652 25378 5704
rect 25406 5652 25412 5704
rect 25464 5652 25470 5704
rect 25516 5692 25544 5723
rect 25590 5720 25596 5772
rect 25648 5760 25654 5772
rect 25777 5763 25835 5769
rect 25777 5760 25789 5763
rect 25648 5732 25789 5760
rect 25648 5720 25654 5732
rect 25777 5729 25789 5732
rect 25823 5760 25835 5763
rect 25866 5760 25872 5772
rect 25823 5732 25872 5760
rect 25823 5729 25835 5732
rect 25777 5723 25835 5729
rect 25866 5720 25872 5732
rect 25924 5720 25930 5772
rect 25958 5720 25964 5772
rect 26016 5720 26022 5772
rect 26326 5720 26332 5772
rect 26384 5760 26390 5772
rect 26712 5760 26740 5800
rect 26970 5788 26976 5800
rect 27028 5788 27034 5840
rect 27338 5828 27344 5840
rect 27264 5800 27344 5828
rect 26384 5732 26740 5760
rect 26384 5720 26390 5732
rect 26878 5720 26884 5772
rect 26936 5720 26942 5772
rect 27264 5769 27292 5800
rect 27338 5788 27344 5800
rect 27396 5788 27402 5840
rect 27448 5828 27476 5856
rect 30282 5828 30288 5840
rect 27448 5800 30288 5828
rect 30282 5788 30288 5800
rect 30340 5788 30346 5840
rect 27249 5763 27307 5769
rect 27249 5729 27261 5763
rect 27295 5729 27307 5763
rect 27249 5723 27307 5729
rect 27706 5720 27712 5772
rect 27764 5760 27770 5772
rect 27982 5760 27988 5772
rect 27764 5732 27988 5760
rect 27764 5720 27770 5732
rect 27982 5720 27988 5732
rect 28040 5760 28046 5772
rect 28445 5763 28503 5769
rect 28445 5760 28457 5763
rect 28040 5732 28457 5760
rect 28040 5720 28046 5732
rect 28445 5729 28457 5732
rect 28491 5729 28503 5763
rect 28445 5723 28503 5729
rect 28721 5763 28779 5769
rect 28721 5729 28733 5763
rect 28767 5760 28779 5763
rect 29086 5760 29092 5772
rect 28767 5732 29092 5760
rect 28767 5729 28779 5732
rect 28721 5723 28779 5729
rect 26786 5692 26792 5704
rect 25516 5664 26792 5692
rect 25516 5636 25544 5664
rect 26786 5652 26792 5664
rect 26844 5652 26850 5704
rect 27341 5695 27399 5701
rect 27341 5661 27353 5695
rect 27387 5692 27399 5695
rect 27522 5692 27528 5704
rect 27387 5664 27528 5692
rect 27387 5661 27399 5664
rect 27341 5655 27399 5661
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 28077 5695 28135 5701
rect 28077 5661 28089 5695
rect 28123 5661 28135 5695
rect 28460 5692 28488 5723
rect 29086 5720 29092 5732
rect 29144 5760 29150 5772
rect 29454 5769 29460 5772
rect 29402 5763 29460 5769
rect 29402 5760 29414 5763
rect 29144 5732 29414 5760
rect 29144 5720 29150 5732
rect 29402 5729 29414 5732
rect 29448 5729 29460 5763
rect 29402 5723 29460 5729
rect 29454 5720 29460 5723
rect 29512 5720 29518 5772
rect 29546 5720 29552 5772
rect 29604 5720 29610 5772
rect 29641 5763 29699 5769
rect 29641 5729 29653 5763
rect 29687 5729 29699 5763
rect 29641 5723 29699 5729
rect 29181 5695 29239 5701
rect 29181 5692 29193 5695
rect 28460 5664 29193 5692
rect 28077 5655 28135 5661
rect 29181 5661 29193 5664
rect 29227 5661 29239 5695
rect 29656 5692 29684 5723
rect 29822 5720 29828 5772
rect 29880 5720 29886 5772
rect 29181 5655 29239 5661
rect 29564 5664 29684 5692
rect 23566 5624 23572 5636
rect 22572 5596 23572 5624
rect 23566 5584 23572 5596
rect 23624 5624 23630 5636
rect 23624 5596 24056 5624
rect 23624 5584 23630 5596
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 12400 5528 16313 5556
rect 12400 5516 12406 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 19429 5559 19487 5565
rect 19429 5525 19441 5559
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 21634 5556 21640 5568
rect 20128 5528 21640 5556
rect 20128 5516 20134 5528
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 22462 5516 22468 5568
rect 22520 5516 22526 5568
rect 23750 5516 23756 5568
rect 23808 5556 23814 5568
rect 23937 5559 23995 5565
rect 23937 5556 23949 5559
rect 23808 5528 23949 5556
rect 23808 5516 23814 5528
rect 23937 5525 23949 5528
rect 23983 5525 23995 5559
rect 24028 5556 24056 5596
rect 25498 5584 25504 5636
rect 25556 5584 25562 5636
rect 26878 5584 26884 5636
rect 26936 5624 26942 5636
rect 28092 5624 28120 5655
rect 26936 5596 28120 5624
rect 28629 5627 28687 5633
rect 26936 5584 26942 5596
rect 28629 5593 28641 5627
rect 28675 5624 28687 5627
rect 29270 5624 29276 5636
rect 28675 5596 29276 5624
rect 28675 5593 28687 5596
rect 28629 5587 28687 5593
rect 29270 5584 29276 5596
rect 29328 5584 29334 5636
rect 25961 5559 26019 5565
rect 25961 5556 25973 5559
rect 24028 5528 25973 5556
rect 23937 5519 23995 5525
rect 25961 5525 25973 5528
rect 26007 5556 26019 5559
rect 26050 5556 26056 5568
rect 26007 5528 26056 5556
rect 26007 5525 26019 5528
rect 25961 5519 26019 5525
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 28442 5516 28448 5568
rect 28500 5556 28506 5568
rect 29564 5556 29592 5664
rect 28500 5528 29592 5556
rect 28500 5516 28506 5528
rect 552 5466 31648 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 11436 5466
rect 11488 5414 11500 5466
rect 11552 5414 11564 5466
rect 11616 5414 11628 5466
rect 11680 5414 11692 5466
rect 11744 5414 19210 5466
rect 19262 5414 19274 5466
rect 19326 5414 19338 5466
rect 19390 5414 19402 5466
rect 19454 5414 19466 5466
rect 19518 5414 26984 5466
rect 27036 5414 27048 5466
rect 27100 5414 27112 5466
rect 27164 5414 27176 5466
rect 27228 5414 27240 5466
rect 27292 5414 31648 5466
rect 552 5392 31648 5414
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6270 5352 6276 5364
rect 5951 5324 6276 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 10410 5352 10416 5364
rect 6380 5324 10416 5352
rect 2498 5244 2504 5296
rect 2556 5244 2562 5296
rect 4982 5244 4988 5296
rect 5040 5284 5046 5296
rect 6380 5284 6408 5324
rect 10410 5312 10416 5324
rect 10468 5352 10474 5364
rect 12434 5352 12440 5364
rect 10468 5324 12440 5352
rect 10468 5312 10474 5324
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 12526 5312 12532 5364
rect 12584 5312 12590 5364
rect 12894 5312 12900 5364
rect 12952 5352 12958 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 12952 5324 13553 5352
rect 12952 5312 12958 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 14826 5312 14832 5364
rect 14884 5352 14890 5364
rect 17313 5355 17371 5361
rect 14884 5324 17264 5352
rect 14884 5312 14890 5324
rect 5040 5256 6408 5284
rect 5040 5244 5046 5256
rect 7834 5244 7840 5296
rect 7892 5244 7898 5296
rect 11238 5244 11244 5296
rect 11296 5284 11302 5296
rect 11698 5284 11704 5296
rect 11296 5256 11704 5284
rect 11296 5244 11302 5256
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 11900 5256 13308 5284
rect 3605 5219 3663 5225
rect 1872 5188 3556 5216
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 1872 5157 1900 5188
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1360 5120 1869 5148
rect 1360 5108 1366 5120
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 2774 5108 2780 5160
rect 2832 5108 2838 5160
rect 3528 5157 3556 5188
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 7006 5216 7012 5228
rect 3651 5188 7012 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 9674 5216 9680 5228
rect 7668 5188 9680 5216
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 4154 5148 4160 5160
rect 3559 5120 4160 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3344 5080 3372 5111
rect 4154 5108 4160 5120
rect 4212 5148 4218 5160
rect 5074 5148 5080 5160
rect 4212 5120 5080 5148
rect 4212 5108 4218 5120
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 6052 5120 6101 5148
rect 6052 5108 6058 5120
rect 6089 5117 6101 5120
rect 6135 5117 6147 5151
rect 6089 5111 6147 5117
rect 6178 5108 6184 5160
rect 6236 5148 6242 5160
rect 6273 5151 6331 5157
rect 6273 5148 6285 5151
rect 6236 5120 6285 5148
rect 6236 5108 6242 5120
rect 6273 5117 6285 5120
rect 6319 5117 6331 5151
rect 6273 5111 6331 5117
rect 6365 5151 6423 5157
rect 6365 5117 6377 5151
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 6457 5151 6515 5157
rect 6457 5117 6469 5151
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 3602 5080 3608 5092
rect 3344 5052 3608 5080
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 6380 5080 6408 5111
rect 6288 5052 6408 5080
rect 6288 5024 6316 5052
rect 6472 5024 6500 5111
rect 6638 5108 6644 5160
rect 6696 5108 6702 5160
rect 7374 5108 7380 5160
rect 7432 5108 7438 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7668 5157 7696 5188
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11900 5225 11928 5256
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 11204 5188 11805 5216
rect 11204 5176 11210 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12526 5216 12532 5228
rect 12023 5188 12532 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 12894 5176 12900 5228
rect 12952 5176 12958 5228
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13170 5216 13176 5228
rect 13035 5188 13176 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13280 5216 13308 5256
rect 14918 5244 14924 5296
rect 14976 5244 14982 5296
rect 15930 5244 15936 5296
rect 15988 5244 15994 5296
rect 17236 5284 17264 5324
rect 17313 5321 17325 5355
rect 17359 5352 17371 5355
rect 17494 5352 17500 5364
rect 17359 5324 17500 5352
rect 17359 5321 17371 5324
rect 17313 5315 17371 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 19058 5312 19064 5364
rect 19116 5312 19122 5364
rect 21453 5355 21511 5361
rect 21453 5321 21465 5355
rect 21499 5352 21511 5355
rect 21542 5352 21548 5364
rect 21499 5324 21548 5352
rect 21499 5321 21511 5324
rect 21453 5315 21511 5321
rect 21542 5312 21548 5324
rect 21600 5312 21606 5364
rect 23934 5312 23940 5364
rect 23992 5312 23998 5364
rect 25314 5352 25320 5364
rect 24044 5324 25320 5352
rect 20346 5284 20352 5296
rect 17236 5256 20352 5284
rect 20346 5244 20352 5256
rect 20404 5284 20410 5296
rect 21082 5284 21088 5296
rect 20404 5256 21088 5284
rect 20404 5244 20410 5256
rect 21082 5244 21088 5256
rect 21140 5244 21146 5296
rect 23750 5244 23756 5296
rect 23808 5284 23814 5296
rect 24044 5284 24072 5324
rect 25314 5312 25320 5324
rect 25372 5312 25378 5364
rect 25593 5355 25651 5361
rect 25593 5321 25605 5355
rect 25639 5352 25651 5355
rect 25774 5352 25780 5364
rect 25639 5324 25780 5352
rect 25639 5321 25651 5324
rect 25593 5315 25651 5321
rect 25774 5312 25780 5324
rect 25832 5312 25838 5364
rect 25866 5312 25872 5364
rect 25924 5352 25930 5364
rect 25924 5324 26464 5352
rect 25924 5312 25930 5324
rect 23808 5256 24072 5284
rect 23808 5244 23814 5256
rect 24118 5244 24124 5296
rect 24176 5244 24182 5296
rect 24394 5244 24400 5296
rect 24452 5284 24458 5296
rect 24762 5284 24768 5296
rect 24452 5256 24768 5284
rect 24452 5244 24458 5256
rect 24762 5244 24768 5256
rect 24820 5284 24826 5296
rect 26326 5284 26332 5296
rect 24820 5256 26332 5284
rect 24820 5244 24826 5256
rect 26326 5244 26332 5256
rect 26384 5244 26390 5296
rect 26436 5293 26464 5324
rect 26602 5312 26608 5364
rect 26660 5312 26666 5364
rect 28997 5355 29055 5361
rect 28997 5321 29009 5355
rect 29043 5352 29055 5355
rect 29822 5352 29828 5364
rect 29043 5324 29828 5352
rect 29043 5321 29055 5324
rect 28997 5315 29055 5321
rect 29822 5312 29828 5324
rect 29880 5312 29886 5364
rect 26421 5287 26479 5293
rect 26421 5253 26433 5287
rect 26467 5253 26479 5287
rect 28074 5284 28080 5296
rect 26421 5247 26479 5253
rect 27356 5256 28080 5284
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13280 5188 14105 5216
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 15102 5216 15108 5228
rect 14139 5188 15108 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 23106 5216 23112 5228
rect 15212 5188 20392 5216
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7524 5120 7573 5148
rect 7524 5108 7530 5120
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 7926 5108 7932 5160
rect 7984 5108 7990 5160
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 11330 5148 11336 5160
rect 9640 5120 11336 5148
rect 9640 5108 9646 5120
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 11698 5108 11704 5160
rect 11756 5148 11762 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11756 5120 12081 5148
rect 11756 5108 11762 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 7392 5080 7420 5108
rect 7392 5052 8294 5080
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 6270 5012 6276 5024
rect 4304 4984 6276 5012
rect 4304 4972 4310 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 6604 4984 7389 5012
rect 6604 4972 6610 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 8266 5012 8294 5052
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 12820 5086 13032 5114
rect 13630 5108 13636 5160
rect 13688 5157 13694 5160
rect 13688 5151 13724 5157
rect 13712 5117 13724 5151
rect 13688 5111 13724 5117
rect 13688 5108 13694 5111
rect 14182 5108 14188 5160
rect 14240 5108 14246 5160
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 14826 5108 14832 5160
rect 14884 5108 14890 5160
rect 15212 5157 15240 5188
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5117 15255 5151
rect 15197 5111 15255 5117
rect 15286 5108 15292 5160
rect 15344 5108 15350 5160
rect 15378 5108 15384 5160
rect 15436 5108 15442 5160
rect 15764 5157 15792 5188
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5117 15807 5151
rect 15749 5111 15807 5117
rect 16022 5108 16028 5160
rect 16080 5108 16086 5160
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 17052 5157 17080 5188
rect 20364 5160 20392 5188
rect 20732 5188 23112 5216
rect 16209 5151 16267 5157
rect 16209 5148 16221 5151
rect 16172 5120 16221 5148
rect 16172 5108 16178 5120
rect 16209 5117 16221 5120
rect 16255 5117 16267 5151
rect 16209 5111 16267 5117
rect 17037 5151 17095 5157
rect 17037 5117 17049 5151
rect 17083 5117 17095 5151
rect 17037 5111 17095 5117
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 18414 5148 18420 5160
rect 17175 5120 18420 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 18414 5108 18420 5120
rect 18472 5108 18478 5160
rect 18690 5108 18696 5160
rect 18748 5108 18754 5160
rect 18782 5108 18788 5160
rect 18840 5108 18846 5160
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18932 5120 18981 5148
rect 18932 5108 18938 5120
rect 18969 5117 18981 5120
rect 19015 5117 19027 5151
rect 18969 5111 19027 5117
rect 19058 5108 19064 5160
rect 19116 5148 19122 5160
rect 20254 5148 20260 5160
rect 19116 5120 20260 5148
rect 19116 5108 19122 5120
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 20732 5157 20760 5188
rect 23106 5176 23112 5188
rect 23164 5216 23170 5228
rect 23201 5219 23259 5225
rect 23201 5216 23213 5219
rect 23164 5188 23213 5216
rect 23164 5176 23170 5188
rect 23201 5185 23213 5188
rect 23247 5185 23259 5219
rect 23201 5179 23259 5185
rect 23569 5219 23627 5225
rect 23569 5185 23581 5219
rect 23615 5216 23627 5219
rect 24670 5216 24676 5228
rect 23615 5188 24676 5216
rect 23615 5185 23627 5188
rect 23569 5179 23627 5185
rect 24670 5176 24676 5188
rect 24728 5216 24734 5228
rect 25958 5216 25964 5228
rect 24728 5188 25964 5216
rect 24728 5176 24734 5188
rect 25958 5176 25964 5188
rect 26016 5216 26022 5228
rect 26145 5219 26203 5225
rect 26145 5216 26157 5219
rect 26016 5188 26157 5216
rect 26016 5176 26022 5188
rect 26145 5185 26157 5188
rect 26191 5216 26203 5219
rect 26191 5188 26740 5216
rect 26191 5185 26203 5188
rect 26145 5179 26203 5185
rect 20625 5151 20683 5157
rect 20625 5148 20637 5151
rect 20404 5120 20637 5148
rect 20404 5108 20410 5120
rect 20625 5117 20637 5120
rect 20671 5117 20683 5151
rect 20625 5111 20683 5117
rect 20717 5151 20775 5157
rect 20717 5117 20729 5151
rect 20763 5117 20775 5151
rect 20717 5111 20775 5117
rect 20898 5108 20904 5160
rect 20956 5108 20962 5160
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5148 21143 5151
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 21131 5120 21189 5148
rect 21131 5117 21143 5120
rect 21085 5111 21143 5117
rect 21177 5117 21189 5120
rect 21223 5117 21235 5151
rect 21177 5111 21235 5117
rect 21450 5108 21456 5160
rect 21508 5108 21514 5160
rect 22646 5108 22652 5160
rect 22704 5148 22710 5160
rect 23385 5151 23443 5157
rect 23385 5148 23397 5151
rect 22704 5120 23397 5148
rect 22704 5108 22710 5120
rect 23385 5117 23397 5120
rect 23431 5117 23443 5151
rect 23385 5111 23443 5117
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 24210 5148 24216 5160
rect 23707 5120 24216 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24210 5108 24216 5120
rect 24268 5108 24274 5160
rect 24394 5108 24400 5160
rect 24452 5108 24458 5160
rect 24486 5108 24492 5160
rect 24544 5148 24550 5160
rect 24765 5151 24823 5157
rect 24765 5148 24777 5151
rect 24544 5120 24777 5148
rect 24544 5108 24550 5120
rect 24765 5117 24777 5120
rect 24811 5117 24823 5151
rect 24765 5111 24823 5117
rect 25041 5151 25099 5157
rect 25041 5117 25053 5151
rect 25087 5148 25099 5151
rect 25087 5120 25268 5148
rect 25087 5117 25099 5120
rect 25041 5111 25099 5117
rect 12820 5080 12848 5086
rect 9456 5052 12848 5080
rect 13004 5080 13032 5086
rect 14461 5083 14519 5089
rect 14461 5080 14473 5083
rect 13004 5052 14473 5080
rect 9456 5040 9462 5052
rect 14461 5049 14473 5052
rect 14507 5049 14519 5083
rect 14461 5043 14519 5049
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5049 15623 5083
rect 15565 5043 15623 5049
rect 11146 5012 11152 5024
rect 8266 4984 11152 5012
rect 7377 4975 7435 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 11388 4984 11621 5012
rect 11388 4972 11394 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 11609 4975 11667 4981
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 11882 5012 11888 5024
rect 11756 4984 11888 5012
rect 11756 4972 11762 4984
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12894 4972 12900 5024
rect 12952 5012 12958 5024
rect 13725 5015 13783 5021
rect 13725 5012 13737 5015
rect 12952 4984 13737 5012
rect 12952 4972 12958 4984
rect 13725 4981 13737 4984
rect 13771 4981 13783 5015
rect 13725 4975 13783 4981
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 15105 5015 15163 5021
rect 15105 5012 15117 5015
rect 14332 4984 15117 5012
rect 14332 4972 14338 4984
rect 15105 4981 15117 4984
rect 15151 5012 15163 5015
rect 15580 5012 15608 5043
rect 15654 5040 15660 5092
rect 15712 5040 15718 5092
rect 17313 5083 17371 5089
rect 17313 5049 17325 5083
rect 17359 5080 17371 5083
rect 17954 5080 17960 5092
rect 17359 5052 17960 5080
rect 17359 5049 17371 5052
rect 17313 5043 17371 5049
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 15151 4984 15608 5012
rect 15151 4981 15163 4984
rect 15105 4975 15163 4981
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 16117 5015 16175 5021
rect 16117 5012 16129 5015
rect 15804 4984 16129 5012
rect 15804 4972 15810 4984
rect 16117 4981 16129 4984
rect 16163 4981 16175 5015
rect 16117 4975 16175 4981
rect 16390 4972 16396 5024
rect 16448 5012 16454 5024
rect 20916 5012 20944 5108
rect 16448 4984 20944 5012
rect 16448 4972 16454 4984
rect 21266 4972 21272 5024
rect 21324 4972 21330 5024
rect 24578 4972 24584 5024
rect 24636 4972 24642 5024
rect 24949 5015 25007 5021
rect 24949 4981 24961 5015
rect 24995 5012 25007 5015
rect 25038 5012 25044 5024
rect 24995 4984 25044 5012
rect 24995 4981 25007 4984
rect 24949 4975 25007 4981
rect 25038 4972 25044 4984
rect 25096 4972 25102 5024
rect 25240 5021 25268 5120
rect 25406 5108 25412 5160
rect 25464 5108 25470 5160
rect 25593 5151 25651 5157
rect 25593 5117 25605 5151
rect 25639 5148 25651 5151
rect 26602 5148 26608 5160
rect 25639 5120 26608 5148
rect 25639 5117 25651 5120
rect 25593 5111 25651 5117
rect 26602 5108 26608 5120
rect 26660 5108 26666 5160
rect 26712 5157 26740 5188
rect 27356 5157 27384 5256
rect 28074 5244 28080 5256
rect 28132 5284 28138 5296
rect 28132 5256 29868 5284
rect 28132 5244 28138 5256
rect 27985 5219 28043 5225
rect 27985 5185 27997 5219
rect 28031 5216 28043 5219
rect 29546 5216 29552 5228
rect 28031 5188 29552 5216
rect 28031 5185 28043 5188
rect 27985 5179 28043 5185
rect 29546 5176 29552 5188
rect 29604 5176 29610 5228
rect 26697 5151 26755 5157
rect 26697 5117 26709 5151
rect 26743 5117 26755 5151
rect 26697 5111 26755 5117
rect 27341 5151 27399 5157
rect 27341 5117 27353 5151
rect 27387 5117 27399 5151
rect 27341 5111 27399 5117
rect 27706 5108 27712 5160
rect 27764 5108 27770 5160
rect 28537 5151 28595 5157
rect 28537 5117 28549 5151
rect 28583 5148 28595 5151
rect 29270 5148 29276 5160
rect 28583 5120 29276 5148
rect 28583 5117 28595 5120
rect 28537 5111 28595 5117
rect 29270 5108 29276 5120
rect 29328 5108 29334 5160
rect 29365 5151 29423 5157
rect 29365 5117 29377 5151
rect 29411 5117 29423 5151
rect 29365 5111 29423 5117
rect 29380 5080 29408 5111
rect 29454 5108 29460 5160
rect 29512 5148 29518 5160
rect 29733 5151 29791 5157
rect 29733 5148 29745 5151
rect 29512 5120 29745 5148
rect 29512 5108 29518 5120
rect 29733 5117 29745 5120
rect 29779 5117 29791 5151
rect 29840 5148 29868 5256
rect 30193 5151 30251 5157
rect 30193 5148 30205 5151
rect 29840 5120 30205 5148
rect 29733 5111 29791 5117
rect 30193 5117 30205 5120
rect 30239 5117 30251 5151
rect 30193 5111 30251 5117
rect 30834 5108 30840 5160
rect 30892 5108 30898 5160
rect 30282 5080 30288 5092
rect 29380 5052 30288 5080
rect 30282 5040 30288 5052
rect 30340 5040 30346 5092
rect 25225 5015 25283 5021
rect 25225 4981 25237 5015
rect 25271 4981 25283 5015
rect 25225 4975 25283 4981
rect 28534 4972 28540 5024
rect 28592 4972 28598 5024
rect 552 4922 31648 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 12096 4922
rect 12148 4870 12160 4922
rect 12212 4870 12224 4922
rect 12276 4870 12288 4922
rect 12340 4870 12352 4922
rect 12404 4870 19870 4922
rect 19922 4870 19934 4922
rect 19986 4870 19998 4922
rect 20050 4870 20062 4922
rect 20114 4870 20126 4922
rect 20178 4870 27644 4922
rect 27696 4870 27708 4922
rect 27760 4870 27772 4922
rect 27824 4870 27836 4922
rect 27888 4870 27900 4922
rect 27952 4870 31648 4922
rect 552 4848 31648 4870
rect 2406 4768 2412 4820
rect 2464 4768 2470 4820
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 3200 4780 3249 4808
rect 3200 4768 3206 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 3973 4811 4031 4817
rect 3973 4777 3985 4811
rect 4019 4808 4031 4811
rect 4246 4808 4252 4820
rect 4019 4780 4252 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 4982 4768 4988 4820
rect 5040 4768 5046 4820
rect 5810 4768 5816 4820
rect 5868 4768 5874 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 6972 4780 12434 4808
rect 6972 4768 6978 4780
rect 2038 4700 2044 4752
rect 2096 4700 2102 4752
rect 3605 4743 3663 4749
rect 2792 4712 3556 4740
rect 2792 4684 2820 4712
rect 3528 4684 3556 4712
rect 3605 4709 3617 4743
rect 3651 4740 3663 4743
rect 7558 4740 7564 4752
rect 3651 4712 7564 4740
rect 3651 4709 3663 4712
rect 3605 4703 3663 4709
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 9674 4740 9680 4752
rect 9508 4712 9680 4740
rect 9508 4684 9536 4712
rect 9674 4700 9680 4712
rect 9732 4700 9738 4752
rect 10410 4700 10416 4752
rect 10468 4740 10474 4752
rect 12406 4740 12434 4780
rect 12526 4768 12532 4820
rect 12584 4808 12590 4820
rect 13078 4808 13084 4820
rect 12584 4780 13084 4808
rect 12584 4768 12590 4780
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 16390 4808 16396 4820
rect 15436 4780 16396 4808
rect 15436 4768 15442 4780
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 17218 4768 17224 4820
rect 17276 4768 17282 4820
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 18598 4808 18604 4820
rect 17460 4780 18604 4808
rect 17460 4768 17466 4780
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 18693 4811 18751 4817
rect 18693 4777 18705 4811
rect 18739 4808 18751 4811
rect 18782 4808 18788 4820
rect 18739 4780 18788 4808
rect 18739 4777 18751 4780
rect 18693 4771 18751 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 19429 4811 19487 4817
rect 19429 4777 19441 4811
rect 19475 4808 19487 4811
rect 21726 4808 21732 4820
rect 19475 4780 21732 4808
rect 19475 4777 19487 4780
rect 19429 4771 19487 4777
rect 21726 4768 21732 4780
rect 21784 4768 21790 4820
rect 22186 4768 22192 4820
rect 22244 4808 22250 4820
rect 22373 4811 22431 4817
rect 22373 4808 22385 4811
rect 22244 4780 22385 4808
rect 22244 4768 22250 4780
rect 22373 4777 22385 4780
rect 22419 4777 22431 4811
rect 22373 4771 22431 4777
rect 25038 4768 25044 4820
rect 25096 4768 25102 4820
rect 29362 4768 29368 4820
rect 29420 4768 29426 4820
rect 17310 4740 17316 4752
rect 10468 4712 11100 4740
rect 12406 4712 17316 4740
rect 10468 4700 10474 4712
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 1857 4675 1915 4681
rect 1857 4672 1869 4675
rect 1360 4644 1869 4672
rect 1360 4632 1366 4644
rect 1857 4641 1869 4644
rect 1903 4672 1915 4675
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 1903 4644 2421 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 2409 4641 2421 4644
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4672 2651 4675
rect 2774 4672 2780 4684
rect 2639 4644 2780 4672
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 2608 4604 2636 4635
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3418 4632 3424 4684
rect 3476 4632 3482 4684
rect 3510 4632 3516 4684
rect 3568 4672 3574 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3568 4644 3801 4672
rect 3568 4632 3574 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 3789 4635 3847 4641
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 4212 4644 4353 4672
rect 4212 4632 4218 4644
rect 4341 4641 4353 4644
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 4939 4644 5028 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 2179 4576 2636 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 4246 4604 4252 4616
rect 3660 4576 4252 4604
rect 3660 4564 3666 4576
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 5000 4468 5028 4644
rect 5074 4632 5080 4684
rect 5132 4632 5138 4684
rect 5994 4632 6000 4684
rect 6052 4632 6058 4684
rect 6086 4632 6092 4684
rect 6144 4672 6150 4684
rect 6365 4675 6423 4681
rect 6365 4672 6377 4675
rect 6144 4644 6377 4672
rect 6144 4632 6150 4644
rect 6365 4641 6377 4644
rect 6411 4672 6423 4675
rect 6454 4672 6460 4684
rect 6411 4644 6460 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6546 4632 6552 4684
rect 6604 4632 6610 4684
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 7742 4632 7748 4684
rect 7800 4632 7806 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 8205 4675 8263 4681
rect 8205 4672 8217 4675
rect 7892 4644 8217 4672
rect 7892 4632 7898 4644
rect 8205 4641 8217 4644
rect 8251 4672 8263 4675
rect 9398 4672 9404 4684
rect 8251 4644 9404 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9490 4632 9496 4684
rect 9548 4632 9554 4684
rect 9582 4632 9588 4684
rect 9640 4632 9646 4684
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 10321 4675 10379 4681
rect 9815 4644 10180 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 6270 4564 6276 4616
rect 6328 4564 6334 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 6472 4576 7941 4604
rect 6196 4536 6224 4564
rect 6472 4536 6500 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8386 4604 8392 4616
rect 8159 4576 8392 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 10152 4536 10180 4644
rect 10321 4641 10333 4675
rect 10367 4672 10379 4675
rect 10962 4672 10968 4684
rect 10367 4644 10968 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 10226 4564 10232 4616
rect 10284 4564 10290 4616
rect 10410 4564 10416 4616
rect 10468 4564 10474 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10551 4576 11008 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 10980 4548 11008 4576
rect 6196 4508 6500 4536
rect 6564 4508 10088 4536
rect 10152 4508 10456 4536
rect 5166 4468 5172 4480
rect 5000 4440 5172 4468
rect 5166 4428 5172 4440
rect 5224 4468 5230 4480
rect 6564 4468 6592 4508
rect 5224 4440 6592 4468
rect 5224 4428 5230 4440
rect 8018 4428 8024 4480
rect 8076 4428 8082 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 9953 4471 10011 4477
rect 9953 4468 9965 4471
rect 9824 4440 9965 4468
rect 9824 4428 9830 4440
rect 9953 4437 9965 4440
rect 9999 4437 10011 4471
rect 10060 4468 10088 4508
rect 10428 4480 10456 4508
rect 10962 4496 10968 4548
rect 11020 4496 11026 4548
rect 11072 4536 11100 4712
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4672 11759 4675
rect 11747 4644 12434 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11204 4576 11805 4604
rect 11204 4564 11210 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 11882 4564 11888 4616
rect 11940 4564 11946 4616
rect 11974 4564 11980 4616
rect 12032 4564 12038 4616
rect 12406 4604 12434 4644
rect 12526 4632 12532 4684
rect 12584 4672 12590 4684
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 12584 4644 15577 4672
rect 12584 4632 12590 4644
rect 15565 4641 15577 4644
rect 15611 4641 15623 4675
rect 15565 4635 15623 4641
rect 15746 4632 15752 4684
rect 15804 4632 15810 4684
rect 16684 4681 16712 4712
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 18414 4700 18420 4752
rect 18472 4740 18478 4752
rect 18509 4743 18567 4749
rect 18509 4740 18521 4743
rect 18472 4712 18521 4740
rect 18472 4700 18478 4712
rect 18509 4709 18521 4712
rect 18555 4709 18567 4743
rect 18800 4740 18828 4768
rect 18800 4712 19012 4740
rect 18509 4703 18567 4709
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 16132 4644 16497 4672
rect 12406 4576 13308 4604
rect 12802 4536 12808 4548
rect 11072 4508 12808 4536
rect 12802 4496 12808 4508
rect 12860 4496 12866 4548
rect 13280 4536 13308 4576
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 16132 4604 16160 4644
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 16669 4675 16727 4681
rect 16669 4641 16681 4675
rect 16715 4641 16727 4675
rect 16669 4635 16727 4641
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 18049 4675 18107 4681
rect 18049 4672 18061 4675
rect 17184 4644 18061 4672
rect 17184 4632 17190 4644
rect 18049 4641 18061 4644
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 18230 4632 18236 4684
rect 18288 4632 18294 4684
rect 18322 4632 18328 4684
rect 18380 4632 18386 4684
rect 18598 4632 18604 4684
rect 18656 4672 18662 4684
rect 18984 4681 19012 4712
rect 19702 4700 19708 4752
rect 19760 4740 19766 4752
rect 19978 4740 19984 4752
rect 19760 4712 19984 4740
rect 19760 4700 19766 4712
rect 19978 4700 19984 4712
rect 20036 4700 20042 4752
rect 20346 4700 20352 4752
rect 20404 4700 20410 4752
rect 21082 4700 21088 4752
rect 21140 4740 21146 4752
rect 25774 4740 25780 4752
rect 21140 4712 24532 4740
rect 21140 4700 21146 4712
rect 18785 4675 18843 4681
rect 18785 4672 18797 4675
rect 18656 4644 18797 4672
rect 18656 4632 18662 4644
rect 18785 4641 18797 4644
rect 18831 4641 18843 4675
rect 18785 4635 18843 4641
rect 18969 4675 19027 4681
rect 18969 4641 18981 4675
rect 19015 4641 19027 4675
rect 18969 4635 19027 4641
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4672 19211 4675
rect 19199 4644 19288 4672
rect 19199 4641 19211 4644
rect 19153 4635 19211 4641
rect 13412 4576 16160 4604
rect 13412 4564 13418 4576
rect 16132 4536 16160 4576
rect 16206 4564 16212 4616
rect 16264 4604 16270 4616
rect 16761 4607 16819 4613
rect 16761 4604 16773 4607
rect 16264 4576 16773 4604
rect 16264 4564 16270 4576
rect 16761 4573 16773 4576
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 17402 4604 17408 4616
rect 16899 4576 17408 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4604 18199 4607
rect 19076 4604 19104 4635
rect 18187 4576 19104 4604
rect 18187 4573 18199 4576
rect 18141 4567 18199 4573
rect 19260 4536 19288 4644
rect 20530 4632 20536 4684
rect 20588 4681 20594 4684
rect 20588 4675 20621 4681
rect 20609 4641 20621 4675
rect 20588 4635 20621 4641
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4672 20775 4675
rect 20806 4672 20812 4684
rect 20763 4644 20812 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 20588 4632 20606 4635
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 22649 4675 22707 4681
rect 22649 4641 22661 4675
rect 22695 4641 22707 4675
rect 22649 4635 22707 4641
rect 20578 4604 20606 4632
rect 21542 4604 21548 4616
rect 20578 4576 21548 4604
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 20714 4536 20720 4548
rect 13280 4508 16068 4536
rect 16132 4508 19012 4536
rect 19260 4508 20720 4536
rect 10318 4468 10324 4480
rect 10060 4440 10324 4468
rect 9953 4431 10011 4437
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 10410 4428 10416 4480
rect 10468 4468 10474 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 10468 4440 11529 4468
rect 10468 4428 10474 4440
rect 11517 4437 11529 4440
rect 11563 4437 11575 4471
rect 11517 4431 11575 4437
rect 11790 4428 11796 4480
rect 11848 4468 11854 4480
rect 15378 4468 15384 4480
rect 11848 4440 15384 4468
rect 11848 4428 11854 4440
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 16040 4468 16068 4508
rect 16850 4468 16856 4480
rect 16040 4440 16856 4468
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 16942 4428 16948 4480
rect 17000 4468 17006 4480
rect 18874 4468 18880 4480
rect 17000 4440 18880 4468
rect 17000 4428 17006 4440
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 18984 4468 19012 4508
rect 20714 4496 20720 4508
rect 20772 4496 20778 4548
rect 22664 4536 22692 4635
rect 22738 4632 22744 4684
rect 22796 4632 22802 4684
rect 22830 4632 22836 4684
rect 22888 4632 22894 4684
rect 23017 4675 23075 4681
rect 23017 4641 23029 4675
rect 23063 4672 23075 4675
rect 23934 4672 23940 4684
rect 23063 4644 23940 4672
rect 23063 4641 23075 4644
rect 23017 4635 23075 4641
rect 23934 4632 23940 4644
rect 23992 4632 23998 4684
rect 24504 4604 24532 4712
rect 25056 4712 25780 4740
rect 25056 4684 25084 4712
rect 25774 4700 25780 4712
rect 25832 4700 25838 4752
rect 25038 4632 25044 4684
rect 25096 4632 25102 4684
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 25188 4644 25237 4672
rect 25188 4632 25194 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 25314 4632 25320 4684
rect 25372 4672 25378 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 25372 4644 26801 4672
rect 25372 4632 25378 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 26789 4635 26847 4641
rect 25148 4604 25176 4632
rect 24504 4576 25176 4604
rect 26694 4564 26700 4616
rect 26752 4564 26758 4616
rect 26804 4604 26832 4635
rect 27430 4632 27436 4684
rect 27488 4632 27494 4684
rect 29457 4675 29515 4681
rect 29457 4641 29469 4675
rect 29503 4672 29515 4675
rect 30006 4672 30012 4684
rect 29503 4644 30012 4672
rect 29503 4641 29515 4644
rect 29457 4635 29515 4641
rect 29472 4604 29500 4635
rect 30006 4632 30012 4644
rect 30064 4632 30070 4684
rect 26804 4576 29500 4604
rect 28902 4536 28908 4548
rect 22664 4508 28908 4536
rect 28902 4496 28908 4508
rect 28960 4496 28966 4548
rect 19518 4468 19524 4480
rect 18984 4440 19524 4468
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 28534 4468 28540 4480
rect 19668 4440 28540 4468
rect 19668 4428 19674 4440
rect 28534 4428 28540 4440
rect 28592 4428 28598 4480
rect 552 4378 31648 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 11436 4378
rect 11488 4326 11500 4378
rect 11552 4326 11564 4378
rect 11616 4326 11628 4378
rect 11680 4326 11692 4378
rect 11744 4326 19210 4378
rect 19262 4326 19274 4378
rect 19326 4326 19338 4378
rect 19390 4326 19402 4378
rect 19454 4326 19466 4378
rect 19518 4326 26984 4378
rect 27036 4326 27048 4378
rect 27100 4326 27112 4378
rect 27164 4326 27176 4378
rect 27228 4326 27240 4378
rect 27292 4326 31648 4378
rect 552 4304 31648 4326
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 4246 4264 4252 4276
rect 3752 4236 4252 4264
rect 3752 4224 3758 4236
rect 4246 4224 4252 4236
rect 4304 4264 4310 4276
rect 7650 4264 7656 4276
rect 4304 4236 7656 4264
rect 4304 4224 4310 4236
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 7834 4224 7840 4276
rect 7892 4264 7898 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7892 4236 7941 4264
rect 7892 4224 7898 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 8018 4224 8024 4276
rect 8076 4264 8082 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 8076 4236 8493 4264
rect 8076 4224 8082 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 9953 4267 10011 4273
rect 9953 4233 9965 4267
rect 9999 4264 10011 4267
rect 10134 4264 10140 4276
rect 9999 4236 10140 4264
rect 9999 4233 10011 4236
rect 9953 4227 10011 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10226 4224 10232 4276
rect 10284 4224 10290 4276
rect 12618 4224 12624 4276
rect 12676 4224 12682 4276
rect 15933 4267 15991 4273
rect 15933 4233 15945 4267
rect 15979 4264 15991 4267
rect 16206 4264 16212 4276
rect 15979 4236 16212 4264
rect 15979 4233 15991 4236
rect 15933 4227 15991 4233
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 19978 4264 19984 4276
rect 16908 4236 19984 4264
rect 16908 4224 16914 4236
rect 19978 4224 19984 4236
rect 20036 4264 20042 4276
rect 20441 4267 20499 4273
rect 20441 4264 20453 4267
rect 20036 4236 20453 4264
rect 20036 4224 20042 4236
rect 20441 4233 20453 4236
rect 20487 4233 20499 4267
rect 20441 4227 20499 4233
rect 20622 4224 20628 4276
rect 20680 4264 20686 4276
rect 22649 4267 22707 4273
rect 20680 4236 22048 4264
rect 20680 4224 20686 4236
rect 5994 4156 6000 4208
rect 6052 4196 6058 4208
rect 8941 4199 8999 4205
rect 8941 4196 8953 4199
rect 6052 4168 8953 4196
rect 6052 4156 6058 4168
rect 8941 4165 8953 4168
rect 8987 4196 8999 4199
rect 12894 4196 12900 4208
rect 8987 4168 12900 4196
rect 8987 4165 8999 4168
rect 8941 4159 8999 4165
rect 12894 4156 12900 4168
rect 12952 4196 12958 4208
rect 12952 4168 13584 4196
rect 12952 4156 12958 4168
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 6178 4128 6184 4140
rect 5399 4100 6184 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6420 4100 6868 4128
rect 6420 4088 6426 4100
rect 6840 4072 6868 4100
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 8202 4128 8208 4140
rect 7576 4100 8208 4128
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3568 4032 3801 4060
rect 3568 4020 3574 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 3789 4023 3847 4029
rect 4154 4020 4160 4072
rect 4212 4020 4218 4072
rect 5166 4020 5172 4072
rect 5224 4020 5230 4072
rect 6546 4020 6552 4072
rect 6604 4020 6610 4072
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7576 4069 7604 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8754 4128 8760 4140
rect 8711 4100 8760 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9674 4128 9680 4140
rect 8956 4100 9680 4128
rect 7101 4063 7159 4069
rect 7101 4060 7113 4063
rect 6880 4032 7113 4060
rect 6880 4020 6886 4032
rect 7101 4029 7113 4032
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7708 4032 8033 4060
rect 7708 4020 7714 4032
rect 8021 4029 8033 4032
rect 8067 4060 8079 4063
rect 8110 4060 8116 4072
rect 8067 4032 8116 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8266 4032 8401 4060
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 4985 3995 5043 4001
rect 4985 3992 4997 3995
rect 3476 3964 4997 3992
rect 3476 3952 3482 3964
rect 4985 3961 4997 3964
rect 5031 3992 5043 3995
rect 5074 3992 5080 4004
rect 5031 3964 5080 3992
rect 5031 3961 5043 3964
rect 4985 3955 5043 3961
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 8266 3992 8294 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8956 4060 8984 4100
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 11241 4131 11299 4137
rect 11241 4128 11253 4131
rect 10060 4100 11253 4128
rect 8389 4023 8447 4029
rect 8680 4032 8984 4060
rect 9033 4063 9091 4069
rect 8680 4001 8708 4032
rect 9033 4029 9045 4063
rect 9079 4060 9091 4063
rect 9490 4060 9496 4072
rect 9079 4032 9496 4060
rect 9079 4029 9091 4032
rect 9033 4023 9091 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 7432 3964 8294 3992
rect 8665 3995 8723 4001
rect 7432 3952 7438 3964
rect 8665 3961 8677 3995
rect 8711 3961 8723 3995
rect 8665 3955 8723 3961
rect 8757 3995 8815 4001
rect 8757 3961 8769 3995
rect 8803 3992 8815 3995
rect 10060 3992 10088 4100
rect 11241 4097 11253 4100
rect 11287 4097 11299 4131
rect 11241 4091 11299 4097
rect 11330 4088 11336 4140
rect 11388 4088 11394 4140
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13446 4128 13452 4140
rect 13127 4100 13452 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13556 4137 13584 4168
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17497 4199 17555 4205
rect 17497 4196 17509 4199
rect 17184 4168 17509 4196
rect 17184 4156 17190 4168
rect 17497 4165 17509 4168
rect 17543 4165 17555 4199
rect 17497 4159 17555 4165
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 20806 4196 20812 4208
rect 18288 4168 20812 4196
rect 18288 4156 18294 4168
rect 20806 4156 20812 4168
rect 20864 4196 20870 4208
rect 21177 4199 21235 4205
rect 21177 4196 21189 4199
rect 20864 4168 21189 4196
rect 20864 4156 20870 4168
rect 21177 4165 21189 4168
rect 21223 4165 21235 4199
rect 21177 4159 21235 4165
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4097 13599 4131
rect 13541 4091 13599 4097
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 19610 4128 19616 4140
rect 14240 4100 19616 4128
rect 14240 4088 14246 4100
rect 19610 4088 19616 4100
rect 19668 4088 19674 4140
rect 19794 4088 19800 4140
rect 19852 4088 19858 4140
rect 20622 4128 20628 4140
rect 20180 4100 20628 4128
rect 10410 4020 10416 4072
rect 10468 4020 10474 4072
rect 10502 4020 10508 4072
rect 10560 4020 10566 4072
rect 10594 4020 10600 4072
rect 10652 4020 10658 4072
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 10704 3992 10732 4023
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 11112 4032 11161 4060
rect 11112 4020 11118 4032
rect 11149 4029 11161 4032
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 11425 4063 11483 4069
rect 11425 4029 11437 4063
rect 11471 4029 11483 4063
rect 11425 4023 11483 4029
rect 11440 3992 11468 4023
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12492 4032 12817 4060
rect 12492 4020 12498 4032
rect 12805 4029 12817 4032
rect 12851 4029 12863 4063
rect 12805 4023 12863 4029
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 13004 3992 13032 4023
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13228 4032 13645 4060
rect 13228 4020 13234 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 13832 3992 13860 4023
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 13964 4032 14565 4060
rect 13964 4020 13970 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14826 4060 14832 4072
rect 14783 4032 14832 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 14458 3992 14464 4004
rect 8803 3964 10088 3992
rect 10152 3964 11468 3992
rect 11532 3964 12952 3992
rect 13004 3964 14464 3992
rect 8803 3961 8815 3964
rect 8757 3955 8815 3961
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3660 3896 4077 3924
rect 3660 3884 3666 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 10042 3924 10048 3936
rect 6328 3896 10048 3924
rect 6328 3884 6334 3896
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10152 3933 10180 3964
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3893 10195 3927
rect 10137 3887 10195 3893
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 11532 3924 11560 3964
rect 10284 3896 11560 3924
rect 10284 3884 10290 3896
rect 11606 3884 11612 3936
rect 11664 3884 11670 3936
rect 12924 3924 12952 3964
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 14936 3992 14964 4023
rect 15286 4020 15292 4072
rect 15344 4020 15350 4072
rect 15470 4020 15476 4072
rect 15528 4020 15534 4072
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4060 15807 4063
rect 15795 4032 15829 4060
rect 15795 4029 15807 4032
rect 15749 4023 15807 4029
rect 15657 3995 15715 4001
rect 15657 3992 15669 3995
rect 14936 3964 15669 3992
rect 15657 3961 15669 3964
rect 15703 3992 15715 3995
rect 15764 3992 15792 4023
rect 15930 4020 15936 4072
rect 15988 4020 15994 4072
rect 17772 4063 17830 4069
rect 17772 4029 17784 4063
rect 17818 4029 17830 4063
rect 17772 4023 17830 4029
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 17954 4060 17960 4072
rect 17911 4032 17960 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 16114 3992 16120 4004
rect 15703 3964 16120 3992
rect 15703 3961 15715 3964
rect 15657 3955 15715 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 17788 3992 17816 4023
rect 17954 4020 17960 4032
rect 18012 4060 18018 4072
rect 18966 4060 18972 4072
rect 18012 4032 18972 4060
rect 18012 4020 18018 4032
rect 18966 4020 18972 4032
rect 19024 4060 19030 4072
rect 19024 4032 19656 4060
rect 19024 4020 19030 4032
rect 17788 3964 17908 3992
rect 17678 3924 17684 3936
rect 12924 3896 17684 3924
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17880 3924 17908 3964
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 19153 3995 19211 4001
rect 19153 3992 19165 3995
rect 18472 3964 19165 3992
rect 18472 3952 18478 3964
rect 19153 3961 19165 3964
rect 19199 3961 19211 3995
rect 19334 3992 19340 4004
rect 19153 3955 19211 3961
rect 19306 3952 19340 3992
rect 19392 3952 19398 4004
rect 19521 3995 19579 4001
rect 19521 3961 19533 3995
rect 19567 3961 19579 3995
rect 19628 3992 19656 4032
rect 19702 4020 19708 4072
rect 19760 4020 19766 4072
rect 20180 4069 20208 4100
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 21192 4128 21220 4159
rect 21192 4100 21772 4128
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4060 19947 4063
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19935 4032 19993 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4029 20223 4063
rect 20714 4060 20720 4072
rect 20165 4023 20223 4029
rect 20364 4032 20720 4060
rect 20180 3992 20208 4023
rect 20364 4001 20392 4032
rect 20714 4020 20720 4032
rect 20772 4060 20778 4072
rect 20772 4032 21220 4060
rect 20772 4020 20778 4032
rect 21192 4001 21220 4032
rect 21542 4020 21548 4072
rect 21600 4060 21606 4072
rect 21744 4069 21772 4100
rect 21636 4063 21694 4069
rect 21636 4060 21648 4063
rect 21600 4032 21648 4060
rect 21600 4020 21606 4032
rect 21636 4029 21648 4032
rect 21682 4029 21694 4063
rect 21636 4023 21694 4029
rect 21729 4063 21787 4069
rect 21729 4029 21741 4063
rect 21775 4029 21787 4063
rect 21729 4023 21787 4029
rect 21818 4020 21824 4072
rect 21876 4020 21882 4072
rect 22020 4069 22048 4236
rect 22649 4233 22661 4267
rect 22695 4264 22707 4267
rect 22738 4264 22744 4276
rect 22695 4236 22744 4264
rect 22695 4233 22707 4236
rect 22649 4227 22707 4233
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 24670 4224 24676 4276
rect 24728 4264 24734 4276
rect 24765 4267 24823 4273
rect 24765 4264 24777 4267
rect 24728 4236 24777 4264
rect 24728 4224 24734 4236
rect 24765 4233 24777 4236
rect 24811 4233 24823 4267
rect 24765 4227 24823 4233
rect 22830 4196 22836 4208
rect 22756 4168 22836 4196
rect 22756 4137 22784 4168
rect 22830 4156 22836 4168
rect 22888 4156 22894 4208
rect 22922 4156 22928 4208
rect 22980 4156 22986 4208
rect 25130 4156 25136 4208
rect 25188 4196 25194 4208
rect 25225 4199 25283 4205
rect 25225 4196 25237 4199
rect 25188 4168 25237 4196
rect 25188 4156 25194 4168
rect 25225 4165 25237 4168
rect 25271 4165 25283 4199
rect 25225 4159 25283 4165
rect 22741 4131 22799 4137
rect 22741 4097 22753 4131
rect 22787 4097 22799 4131
rect 22940 4128 22968 4156
rect 24121 4131 24179 4137
rect 24121 4128 24133 4131
rect 22940 4100 24133 4128
rect 22741 4091 22799 4097
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4029 22063 4063
rect 22005 4023 22063 4029
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 22462 4060 22468 4072
rect 22419 4032 22468 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 22462 4020 22468 4032
rect 22520 4060 22526 4072
rect 22925 4063 22983 4069
rect 22925 4060 22937 4063
rect 22520 4032 22937 4060
rect 22520 4020 22526 4032
rect 22925 4029 22937 4032
rect 22971 4029 22983 4063
rect 22925 4023 22983 4029
rect 23017 4063 23075 4069
rect 23017 4029 23029 4063
rect 23063 4029 23075 4063
rect 23017 4023 23075 4029
rect 19628 3964 20208 3992
rect 20349 3995 20407 4001
rect 19521 3955 19579 3961
rect 20349 3961 20361 3995
rect 20395 3961 20407 3995
rect 20349 3955 20407 3961
rect 21177 3995 21235 4001
rect 21177 3961 21189 3995
rect 21223 3961 21235 3995
rect 21177 3955 21235 3961
rect 19306 3924 19334 3952
rect 17880 3896 19334 3924
rect 19536 3924 19564 3955
rect 21358 3952 21364 4004
rect 21416 3992 21422 4004
rect 22278 3992 22284 4004
rect 21416 3964 22284 3992
rect 21416 3952 21422 3964
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 22649 3995 22707 4001
rect 22649 3961 22661 3995
rect 22695 3992 22707 3995
rect 22830 3992 22836 4004
rect 22695 3964 22836 3992
rect 22695 3961 22707 3964
rect 22649 3955 22707 3961
rect 22830 3952 22836 3964
rect 22888 3952 22894 4004
rect 20530 3924 20536 3936
rect 19536 3896 20536 3924
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 21818 3924 21824 3936
rect 20772 3896 21824 3924
rect 20772 3884 20778 3896
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22462 3884 22468 3936
rect 22520 3924 22526 3936
rect 23032 3924 23060 4023
rect 23198 4020 23204 4072
rect 23256 4020 23262 4072
rect 23308 4069 23336 4100
rect 24121 4097 24133 4100
rect 24167 4097 24179 4131
rect 24121 4091 24179 4097
rect 24210 4088 24216 4140
rect 24268 4128 24274 4140
rect 24268 4100 25360 4128
rect 24268 4088 24274 4100
rect 24412 4069 24440 4100
rect 25332 4069 25360 4100
rect 25958 4088 25964 4140
rect 26016 4088 26022 4140
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 24397 4063 24455 4069
rect 24397 4029 24409 4063
rect 24443 4029 24455 4063
rect 24397 4023 24455 4029
rect 24857 4063 24915 4069
rect 24857 4029 24869 4063
rect 24903 4060 24915 4063
rect 25317 4063 25375 4069
rect 24903 4032 25268 4060
rect 24903 4029 24915 4032
rect 24857 4023 24915 4029
rect 24489 3995 24547 4001
rect 24489 3961 24501 3995
rect 24535 3992 24547 3995
rect 25038 3992 25044 4004
rect 24535 3964 25044 3992
rect 24535 3961 24547 3964
rect 24489 3955 24547 3961
rect 25038 3952 25044 3964
rect 25096 3952 25102 4004
rect 25240 3992 25268 4032
rect 25317 4029 25329 4063
rect 25363 4060 25375 4063
rect 25498 4060 25504 4072
rect 25363 4032 25504 4060
rect 25363 4029 25375 4032
rect 25317 4023 25375 4029
rect 25498 4020 25504 4032
rect 25556 4020 25562 4072
rect 25866 4020 25872 4072
rect 25924 4020 25930 4072
rect 25884 3992 25912 4020
rect 25240 3964 25912 3992
rect 22520 3896 23060 3924
rect 22520 3884 22526 3896
rect 24026 3884 24032 3936
rect 24084 3924 24090 3936
rect 24581 3927 24639 3933
rect 24581 3924 24593 3927
rect 24084 3896 24593 3924
rect 24084 3884 24090 3896
rect 24581 3893 24593 3896
rect 24627 3893 24639 3927
rect 24581 3887 24639 3893
rect 552 3834 31648 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 12096 3834
rect 12148 3782 12160 3834
rect 12212 3782 12224 3834
rect 12276 3782 12288 3834
rect 12340 3782 12352 3834
rect 12404 3782 19870 3834
rect 19922 3782 19934 3834
rect 19986 3782 19998 3834
rect 20050 3782 20062 3834
rect 20114 3782 20126 3834
rect 20178 3782 27644 3834
rect 27696 3782 27708 3834
rect 27760 3782 27772 3834
rect 27824 3782 27836 3834
rect 27888 3782 27900 3834
rect 27952 3782 31648 3834
rect 552 3760 31648 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3513 3723 3571 3729
rect 3513 3720 3525 3723
rect 3476 3692 3525 3720
rect 3476 3680 3482 3692
rect 3513 3689 3525 3692
rect 3559 3689 3571 3723
rect 3513 3683 3571 3689
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 4948 3692 14228 3720
rect 4948 3680 4954 3692
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 3145 3655 3203 3661
rect 3145 3652 3157 3655
rect 3108 3624 3157 3652
rect 3108 3612 3114 3624
rect 3145 3621 3157 3624
rect 3191 3652 3203 3655
rect 5718 3652 5724 3664
rect 3191 3624 5724 3652
rect 3191 3621 3203 3624
rect 3145 3615 3203 3621
rect 5718 3612 5724 3624
rect 5776 3652 5782 3664
rect 5776 3624 6684 3652
rect 5776 3612 5782 3624
rect 3234 3544 3240 3596
rect 3292 3544 3298 3596
rect 3326 3544 3332 3596
rect 3384 3584 3390 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3384 3556 3433 3584
rect 3384 3544 3390 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 4062 3584 4068 3596
rect 3559 3556 4068 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 6656 3593 6684 3624
rect 8386 3612 8392 3664
rect 8444 3652 8450 3664
rect 8481 3655 8539 3661
rect 8481 3652 8493 3655
rect 8444 3624 8493 3652
rect 8444 3612 8450 3624
rect 8481 3621 8493 3624
rect 8527 3621 8539 3655
rect 8481 3615 8539 3621
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 10827 3624 13768 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 6641 3587 6699 3593
rect 6641 3553 6653 3587
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6880 3556 7021 3584
rect 6880 3544 6886 3556
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 7009 3547 7067 3553
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 10643 3556 12848 3584
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 3252 3516 3280 3544
rect 6546 3516 6552 3528
rect 3252 3488 6552 3516
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 10520 3516 10548 3547
rect 12820 3516 12848 3556
rect 12894 3544 12900 3596
rect 12952 3544 12958 3596
rect 13740 3593 13768 3624
rect 12989 3587 13047 3593
rect 12989 3553 13001 3587
rect 13035 3553 13047 3587
rect 12989 3547 13047 3553
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3553 13783 3587
rect 13725 3547 13783 3553
rect 13004 3516 13032 3547
rect 10520 3488 12480 3516
rect 12820 3488 13032 3516
rect 13740 3516 13768 3547
rect 13906 3544 13912 3596
rect 13964 3544 13970 3596
rect 13998 3516 14004 3528
rect 13740 3488 14004 3516
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 12342 3448 12348 3460
rect 2464 3420 12348 3448
rect 2464 3408 2470 3420
rect 12342 3408 12348 3420
rect 12400 3408 12406 3460
rect 12452 3448 12480 3488
rect 12894 3448 12900 3460
rect 12452 3420 12900 3448
rect 12894 3408 12900 3420
rect 12952 3408 12958 3460
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 3694 3380 3700 3392
rect 3375 3352 3700 3380
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 10502 3340 10508 3392
rect 10560 3340 10566 3392
rect 13004 3380 13032 3488
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14200 3516 14228 3692
rect 14642 3680 14648 3732
rect 14700 3680 14706 3732
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 20714 3720 20720 3732
rect 19392 3692 20720 3720
rect 19392 3680 19398 3692
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 21266 3680 21272 3732
rect 21324 3720 21330 3732
rect 31386 3720 31392 3732
rect 21324 3692 31392 3720
rect 21324 3680 21330 3692
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 14458 3612 14464 3664
rect 14516 3652 14522 3664
rect 22462 3652 22468 3664
rect 14516 3624 22468 3652
rect 14516 3612 14522 3624
rect 22462 3612 22468 3624
rect 22520 3612 22526 3664
rect 14274 3544 14280 3596
rect 14332 3544 14338 3596
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 14424 3556 14469 3584
rect 14424 3544 14430 3556
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 21358 3584 21364 3596
rect 16540 3556 21364 3584
rect 16540 3544 16546 3556
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 24854 3516 24860 3528
rect 14200 3488 24860 3516
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 14093 3451 14151 3457
rect 14093 3417 14105 3451
rect 14139 3448 14151 3451
rect 14458 3448 14464 3460
rect 14139 3420 14464 3448
rect 14139 3417 14151 3420
rect 14093 3411 14151 3417
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14734 3380 14740 3392
rect 13004 3352 14740 3380
rect 14734 3340 14740 3352
rect 14792 3380 14798 3392
rect 15470 3380 15476 3392
rect 14792 3352 15476 3380
rect 14792 3340 14798 3352
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 552 3290 31648 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 11436 3290
rect 11488 3238 11500 3290
rect 11552 3238 11564 3290
rect 11616 3238 11628 3290
rect 11680 3238 11692 3290
rect 11744 3238 19210 3290
rect 19262 3238 19274 3290
rect 19326 3238 19338 3290
rect 19390 3238 19402 3290
rect 19454 3238 19466 3290
rect 19518 3238 26984 3290
rect 27036 3238 27048 3290
rect 27100 3238 27112 3290
rect 27164 3238 27176 3290
rect 27228 3238 27240 3290
rect 27292 3238 31648 3290
rect 552 3216 31648 3238
rect 552 2746 31648 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 12096 2746
rect 12148 2694 12160 2746
rect 12212 2694 12224 2746
rect 12276 2694 12288 2746
rect 12340 2694 12352 2746
rect 12404 2694 19870 2746
rect 19922 2694 19934 2746
rect 19986 2694 19998 2746
rect 20050 2694 20062 2746
rect 20114 2694 20126 2746
rect 20178 2694 27644 2746
rect 27696 2694 27708 2746
rect 27760 2694 27772 2746
rect 27824 2694 27836 2746
rect 27888 2694 27900 2746
rect 27952 2694 31648 2746
rect 552 2672 31648 2694
rect 1026 2592 1032 2644
rect 1084 2632 1090 2644
rect 24578 2632 24584 2644
rect 1084 2604 24584 2632
rect 1084 2592 1090 2604
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 2222 2524 2228 2576
rect 2280 2564 2286 2576
rect 24854 2564 24860 2576
rect 2280 2536 24860 2564
rect 2280 2524 2286 2536
rect 24854 2524 24860 2536
rect 24912 2524 24918 2576
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 23382 2496 23388 2508
rect 8352 2468 23388 2496
rect 8352 2456 8358 2468
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 566 2388 572 2440
rect 624 2428 630 2440
rect 11882 2428 11888 2440
rect 624 2400 11888 2428
rect 624 2388 630 2400
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 552 2202 31648 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 11436 2202
rect 11488 2150 11500 2202
rect 11552 2150 11564 2202
rect 11616 2150 11628 2202
rect 11680 2150 11692 2202
rect 11744 2150 19210 2202
rect 19262 2150 19274 2202
rect 19326 2150 19338 2202
rect 19390 2150 19402 2202
rect 19454 2150 19466 2202
rect 19518 2150 26984 2202
rect 27036 2150 27048 2202
rect 27100 2150 27112 2202
rect 27164 2150 27176 2202
rect 27228 2150 27240 2202
rect 27292 2150 31648 2202
rect 552 2128 31648 2150
rect 552 1658 31648 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 12096 1658
rect 12148 1606 12160 1658
rect 12212 1606 12224 1658
rect 12276 1606 12288 1658
rect 12340 1606 12352 1658
rect 12404 1606 19870 1658
rect 19922 1606 19934 1658
rect 19986 1606 19998 1658
rect 20050 1606 20062 1658
rect 20114 1606 20126 1658
rect 20178 1606 27644 1658
rect 27696 1606 27708 1658
rect 27760 1606 27772 1658
rect 27824 1606 27836 1658
rect 27888 1606 27900 1658
rect 27952 1606 31648 1658
rect 552 1584 31648 1606
rect 552 1114 31648 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 11436 1114
rect 11488 1062 11500 1114
rect 11552 1062 11564 1114
rect 11616 1062 11628 1114
rect 11680 1062 11692 1114
rect 11744 1062 19210 1114
rect 19262 1062 19274 1114
rect 19326 1062 19338 1114
rect 19390 1062 19402 1114
rect 19454 1062 19466 1114
rect 19518 1062 26984 1114
rect 27036 1062 27048 1114
rect 27100 1062 27112 1114
rect 27164 1062 27176 1114
rect 27228 1062 27240 1114
rect 27292 1062 31648 1114
rect 552 1040 31648 1062
rect 552 570 31648 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 12096 570
rect 12148 518 12160 570
rect 12212 518 12224 570
rect 12276 518 12288 570
rect 12340 518 12352 570
rect 12404 518 19870 570
rect 19922 518 19934 570
rect 19986 518 19998 570
rect 20050 518 20062 570
rect 20114 518 20126 570
rect 20178 518 27644 570
rect 27696 518 27708 570
rect 27760 518 27772 570
rect 27824 518 27836 570
rect 27888 518 27900 570
rect 27952 518 31648 570
rect 552 496 31648 518
<< via1 >>
rect 11980 21972 12032 22024
rect 26884 21972 26936 22024
rect 13820 21904 13872 21956
rect 26240 21904 26292 21956
rect 27988 21904 28040 21956
rect 30932 21904 30984 21956
rect 9128 21836 9180 21888
rect 18788 21836 18840 21888
rect 24768 21836 24820 21888
rect 27528 21836 27580 21888
rect 30288 21836 30340 21888
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 11436 21734 11488 21786
rect 11500 21734 11552 21786
rect 11564 21734 11616 21786
rect 11628 21734 11680 21786
rect 11692 21734 11744 21786
rect 19210 21734 19262 21786
rect 19274 21734 19326 21786
rect 19338 21734 19390 21786
rect 19402 21734 19454 21786
rect 19466 21734 19518 21786
rect 26984 21734 27036 21786
rect 27048 21734 27100 21786
rect 27112 21734 27164 21786
rect 27176 21734 27228 21786
rect 27240 21734 27292 21786
rect 6184 21675 6236 21684
rect 6184 21641 6193 21675
rect 6193 21641 6227 21675
rect 6227 21641 6236 21675
rect 6184 21632 6236 21641
rect 6736 21675 6788 21684
rect 6736 21641 6745 21675
rect 6745 21641 6779 21675
rect 6779 21641 6788 21675
rect 6736 21632 6788 21641
rect 7288 21675 7340 21684
rect 7288 21641 7297 21675
rect 7297 21641 7331 21675
rect 7331 21641 7340 21675
rect 7288 21632 7340 21641
rect 7840 21675 7892 21684
rect 7840 21641 7849 21675
rect 7849 21641 7883 21675
rect 7883 21641 7892 21675
rect 7840 21632 7892 21641
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 9588 21632 9640 21684
rect 10048 21675 10100 21684
rect 10048 21641 10057 21675
rect 10057 21641 10091 21675
rect 10091 21641 10100 21675
rect 10048 21632 10100 21641
rect 10600 21675 10652 21684
rect 10600 21641 10609 21675
rect 10609 21641 10643 21675
rect 10643 21641 10652 21675
rect 10600 21632 10652 21641
rect 11152 21675 11204 21684
rect 11152 21641 11161 21675
rect 11161 21641 11195 21675
rect 11195 21641 11204 21675
rect 11152 21632 11204 21641
rect 11428 21632 11480 21684
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 13360 21675 13412 21684
rect 13360 21641 13369 21675
rect 13369 21641 13403 21675
rect 13403 21641 13412 21675
rect 13360 21632 13412 21641
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 16672 21632 16724 21684
rect 22284 21632 22336 21684
rect 23112 21675 23164 21684
rect 23112 21641 23121 21675
rect 23121 21641 23155 21675
rect 23155 21641 23164 21675
rect 23112 21632 23164 21641
rect 26424 21632 26476 21684
rect 10784 21564 10836 21616
rect 13820 21564 13872 21616
rect 21180 21564 21232 21616
rect 25228 21564 25280 21616
rect 28356 21564 28408 21616
rect 11336 21496 11388 21548
rect 14648 21496 14700 21548
rect 14740 21496 14792 21548
rect 17224 21496 17276 21548
rect 9956 21428 10008 21480
rect 16396 21471 16448 21480
rect 16396 21437 16405 21471
rect 16405 21437 16439 21471
rect 16439 21437 16448 21471
rect 16396 21428 16448 21437
rect 18420 21539 18472 21548
rect 18420 21505 18429 21539
rect 18429 21505 18463 21539
rect 18463 21505 18472 21539
rect 18420 21496 18472 21505
rect 19432 21496 19484 21548
rect 7840 21292 7892 21344
rect 9036 21292 9088 21344
rect 10600 21292 10652 21344
rect 11796 21335 11848 21344
rect 11796 21301 11805 21335
rect 11805 21301 11839 21335
rect 11839 21301 11848 21335
rect 11796 21292 11848 21301
rect 14280 21403 14332 21412
rect 14280 21369 14289 21403
rect 14289 21369 14323 21403
rect 14323 21369 14332 21403
rect 14280 21360 14332 21369
rect 14740 21360 14792 21412
rect 16120 21292 16172 21344
rect 16764 21360 16816 21412
rect 18972 21403 19024 21412
rect 18972 21369 18981 21403
rect 18981 21369 19015 21403
rect 19015 21369 19024 21403
rect 18972 21360 19024 21369
rect 20260 21360 20312 21412
rect 17316 21292 17368 21344
rect 18328 21292 18380 21344
rect 20628 21360 20680 21412
rect 20904 21335 20956 21344
rect 20904 21301 20931 21335
rect 20931 21301 20956 21335
rect 20904 21292 20956 21301
rect 21088 21403 21140 21412
rect 21088 21369 21097 21403
rect 21097 21369 21131 21403
rect 21131 21369 21140 21403
rect 21088 21360 21140 21369
rect 22928 21428 22980 21480
rect 23020 21428 23072 21480
rect 24860 21496 24912 21548
rect 26332 21496 26384 21548
rect 26056 21428 26108 21480
rect 24124 21360 24176 21412
rect 24216 21403 24268 21412
rect 24216 21369 24225 21403
rect 24225 21369 24259 21403
rect 24259 21369 24268 21403
rect 24216 21360 24268 21369
rect 23112 21292 23164 21344
rect 24032 21292 24084 21344
rect 24308 21292 24360 21344
rect 26148 21403 26200 21412
rect 26148 21369 26157 21403
rect 26157 21369 26191 21403
rect 26191 21369 26200 21403
rect 26148 21360 26200 21369
rect 26608 21292 26660 21344
rect 27988 21360 28040 21412
rect 28264 21403 28316 21412
rect 28264 21369 28273 21403
rect 28273 21369 28307 21403
rect 28307 21369 28316 21403
rect 28264 21360 28316 21369
rect 28080 21292 28132 21344
rect 28172 21292 28224 21344
rect 28540 21335 28592 21344
rect 28540 21301 28549 21335
rect 28549 21301 28583 21335
rect 28583 21301 28592 21335
rect 28540 21292 28592 21301
rect 28632 21335 28684 21344
rect 28632 21301 28641 21335
rect 28641 21301 28675 21335
rect 28675 21301 28684 21335
rect 28632 21292 28684 21301
rect 31208 21428 31260 21480
rect 31392 21428 31444 21480
rect 29368 21360 29420 21412
rect 30564 21360 30616 21412
rect 29000 21292 29052 21344
rect 30196 21292 30248 21344
rect 30840 21335 30892 21344
rect 30840 21301 30849 21335
rect 30849 21301 30883 21335
rect 30883 21301 30892 21335
rect 30840 21292 30892 21301
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 12096 21190 12148 21242
rect 12160 21190 12212 21242
rect 12224 21190 12276 21242
rect 12288 21190 12340 21242
rect 12352 21190 12404 21242
rect 19870 21190 19922 21242
rect 19934 21190 19986 21242
rect 19998 21190 20050 21242
rect 20062 21190 20114 21242
rect 20126 21190 20178 21242
rect 27644 21190 27696 21242
rect 27708 21190 27760 21242
rect 27772 21190 27824 21242
rect 27836 21190 27888 21242
rect 27900 21190 27952 21242
rect 10600 21131 10652 21140
rect 10600 21097 10609 21131
rect 10609 21097 10643 21131
rect 10643 21097 10652 21131
rect 10600 21088 10652 21097
rect 9588 21020 9640 21072
rect 11244 21088 11296 21140
rect 11428 21131 11480 21140
rect 11428 21097 11437 21131
rect 11437 21097 11471 21131
rect 11471 21097 11480 21131
rect 11428 21088 11480 21097
rect 7656 20995 7708 21004
rect 7656 20961 7665 20995
rect 7665 20961 7699 20995
rect 7699 20961 7708 20995
rect 7656 20952 7708 20961
rect 7840 20995 7892 21004
rect 7840 20961 7849 20995
rect 7849 20961 7883 20995
rect 7883 20961 7892 20995
rect 7840 20952 7892 20961
rect 7196 20884 7248 20936
rect 9956 20884 10008 20936
rect 10600 20995 10652 21004
rect 10600 20961 10609 20995
rect 10609 20961 10643 20995
rect 10643 20961 10652 20995
rect 10600 20952 10652 20961
rect 11796 21063 11848 21072
rect 11796 21029 11805 21063
rect 11805 21029 11839 21063
rect 11839 21029 11848 21063
rect 11796 21020 11848 21029
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 16764 21131 16816 21140
rect 16764 21097 16773 21131
rect 16773 21097 16807 21131
rect 16807 21097 16816 21131
rect 16764 21088 16816 21097
rect 17316 21088 17368 21140
rect 21916 21088 21968 21140
rect 14740 21020 14792 21072
rect 10968 20995 11020 21004
rect 10968 20961 10977 20995
rect 10977 20961 11011 20995
rect 11011 20961 11020 20995
rect 10968 20952 11020 20961
rect 13084 20952 13136 21004
rect 11152 20816 11204 20868
rect 10600 20748 10652 20800
rect 10968 20748 11020 20800
rect 11336 20884 11388 20936
rect 12440 20884 12492 20936
rect 14096 20995 14148 21004
rect 14096 20961 14105 20995
rect 14105 20961 14139 20995
rect 14139 20961 14148 20995
rect 14096 20952 14148 20961
rect 16488 21020 16540 21072
rect 17224 21020 17276 21072
rect 18144 21020 18196 21072
rect 19064 21063 19116 21072
rect 19064 21029 19073 21063
rect 19073 21029 19107 21063
rect 19107 21029 19116 21063
rect 19064 21020 19116 21029
rect 23112 21088 23164 21140
rect 24216 21088 24268 21140
rect 28080 21088 28132 21140
rect 28816 21088 28868 21140
rect 29276 21088 29328 21140
rect 29368 21131 29420 21140
rect 29368 21097 29377 21131
rect 29377 21097 29411 21131
rect 29411 21097 29420 21131
rect 29368 21088 29420 21097
rect 30564 21088 30616 21140
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 16028 20952 16080 21004
rect 16120 20995 16172 21004
rect 16120 20961 16129 20995
rect 16129 20961 16163 20995
rect 16163 20961 16172 20995
rect 16120 20952 16172 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 20628 20995 20680 21004
rect 20628 20961 20637 20995
rect 20637 20961 20671 20995
rect 20671 20961 20680 20995
rect 20628 20952 20680 20961
rect 20996 20952 21048 21004
rect 21272 20995 21324 21004
rect 21272 20961 21281 20995
rect 21281 20961 21315 20995
rect 21315 20961 21324 20995
rect 21272 20952 21324 20961
rect 21548 20995 21600 21004
rect 21548 20961 21557 20995
rect 21557 20961 21591 20995
rect 21591 20961 21600 20995
rect 21548 20952 21600 20961
rect 22928 20952 22980 21004
rect 23480 20995 23532 21004
rect 23480 20961 23489 20995
rect 23489 20961 23523 20995
rect 23523 20961 23532 20995
rect 23480 20952 23532 20961
rect 15476 20884 15528 20936
rect 17040 20884 17092 20936
rect 18052 20884 18104 20936
rect 19616 20884 19668 20936
rect 21456 20884 21508 20936
rect 15384 20816 15436 20868
rect 16488 20816 16540 20868
rect 19432 20816 19484 20868
rect 19800 20816 19852 20868
rect 23664 20816 23716 20868
rect 24032 20995 24084 21004
rect 24032 20961 24041 20995
rect 24041 20961 24075 20995
rect 24075 20961 24084 20995
rect 24032 20952 24084 20961
rect 26424 20952 26476 21004
rect 28724 21020 28776 21072
rect 28908 21063 28960 21072
rect 28908 21029 28917 21063
rect 28917 21029 28951 21063
rect 28951 21029 28960 21063
rect 28908 21020 28960 21029
rect 29828 21063 29880 21072
rect 29828 21029 29863 21063
rect 29863 21029 29880 21063
rect 29828 21020 29880 21029
rect 30932 21063 30984 21072
rect 30932 21029 30941 21063
rect 30941 21029 30975 21063
rect 30975 21029 30984 21063
rect 30932 21020 30984 21029
rect 27344 20995 27396 21004
rect 27344 20961 27353 20995
rect 27353 20961 27387 20995
rect 27387 20961 27396 20995
rect 27344 20952 27396 20961
rect 27528 20995 27580 21004
rect 27528 20961 27537 20995
rect 27537 20961 27571 20995
rect 27571 20961 27580 20995
rect 27528 20952 27580 20961
rect 27620 20995 27672 21004
rect 27620 20961 27655 20995
rect 27655 20961 27672 20995
rect 27620 20952 27672 20961
rect 28816 20995 28868 21004
rect 28816 20961 28825 20995
rect 28825 20961 28859 20995
rect 28859 20961 28868 20995
rect 28816 20952 28868 20961
rect 24216 20927 24268 20936
rect 24216 20893 24225 20927
rect 24225 20893 24259 20927
rect 24259 20893 24268 20927
rect 24216 20884 24268 20893
rect 24768 20884 24820 20936
rect 25780 20884 25832 20936
rect 28448 20927 28500 20936
rect 28448 20893 28457 20927
rect 28457 20893 28491 20927
rect 28491 20893 28500 20927
rect 28448 20884 28500 20893
rect 29552 20995 29604 21004
rect 29552 20961 29561 20995
rect 29561 20961 29595 20995
rect 29595 20961 29604 20995
rect 29552 20952 29604 20961
rect 29644 20995 29696 21004
rect 29644 20961 29653 20995
rect 29653 20961 29687 20995
rect 29687 20961 29696 20995
rect 29644 20952 29696 20961
rect 29736 20995 29788 21004
rect 29736 20961 29745 20995
rect 29745 20961 29779 20995
rect 29779 20961 29788 20995
rect 29736 20952 29788 20961
rect 25964 20816 26016 20868
rect 29460 20816 29512 20868
rect 30196 20884 30248 20936
rect 31208 20884 31260 20936
rect 12900 20748 12952 20800
rect 15200 20748 15252 20800
rect 16764 20748 16816 20800
rect 19708 20748 19760 20800
rect 20168 20748 20220 20800
rect 20720 20748 20772 20800
rect 24124 20748 24176 20800
rect 26332 20748 26384 20800
rect 26608 20748 26660 20800
rect 27344 20748 27396 20800
rect 29092 20748 29144 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 11436 20646 11488 20698
rect 11500 20646 11552 20698
rect 11564 20646 11616 20698
rect 11628 20646 11680 20698
rect 11692 20646 11744 20698
rect 19210 20646 19262 20698
rect 19274 20646 19326 20698
rect 19338 20646 19390 20698
rect 19402 20646 19454 20698
rect 19466 20646 19518 20698
rect 26984 20646 27036 20698
rect 27048 20646 27100 20698
rect 27112 20646 27164 20698
rect 27176 20646 27228 20698
rect 27240 20646 27292 20698
rect 13728 20544 13780 20596
rect 8484 20476 8536 20528
rect 9220 20519 9272 20528
rect 9220 20485 9229 20519
rect 9229 20485 9263 20519
rect 9263 20485 9272 20519
rect 9220 20476 9272 20485
rect 14096 20544 14148 20596
rect 14464 20587 14516 20596
rect 14464 20553 14473 20587
rect 14473 20553 14507 20587
rect 14507 20553 14516 20587
rect 14464 20544 14516 20553
rect 16396 20544 16448 20596
rect 7656 20408 7708 20460
rect 8852 20340 8904 20392
rect 8944 20383 8996 20392
rect 8944 20349 8953 20383
rect 8953 20349 8987 20383
rect 8987 20349 8996 20383
rect 8944 20340 8996 20349
rect 9036 20383 9088 20392
rect 9036 20349 9045 20383
rect 9045 20349 9079 20383
rect 9079 20349 9088 20383
rect 9036 20340 9088 20349
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 10508 20340 10560 20392
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 13452 20408 13504 20460
rect 13728 20383 13780 20392
rect 13728 20349 13737 20383
rect 13737 20349 13771 20383
rect 13771 20349 13780 20383
rect 13728 20340 13780 20349
rect 14096 20408 14148 20460
rect 15384 20408 15436 20460
rect 16488 20451 16540 20460
rect 16488 20417 16497 20451
rect 16497 20417 16531 20451
rect 16531 20417 16540 20451
rect 16488 20408 16540 20417
rect 16764 20451 16816 20460
rect 16764 20417 16773 20451
rect 16773 20417 16807 20451
rect 16807 20417 16816 20451
rect 16764 20408 16816 20417
rect 17960 20544 18012 20596
rect 18972 20587 19024 20596
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 20076 20544 20128 20596
rect 20352 20544 20404 20596
rect 21272 20544 21324 20596
rect 22928 20544 22980 20596
rect 23940 20587 23992 20596
rect 23940 20553 23949 20587
rect 23949 20553 23983 20587
rect 23983 20553 23992 20587
rect 23940 20544 23992 20553
rect 25964 20587 26016 20596
rect 25964 20553 25973 20587
rect 25973 20553 26007 20587
rect 26007 20553 26016 20587
rect 25964 20544 26016 20553
rect 26516 20544 26568 20596
rect 18880 20476 18932 20528
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 14740 20340 14792 20392
rect 19156 20383 19208 20392
rect 19156 20349 19165 20383
rect 19165 20349 19199 20383
rect 19199 20349 19208 20383
rect 19156 20340 19208 20349
rect 19708 20408 19760 20460
rect 11060 20315 11112 20324
rect 11060 20281 11069 20315
rect 11069 20281 11103 20315
rect 11103 20281 11112 20315
rect 11060 20272 11112 20281
rect 11336 20272 11388 20324
rect 9312 20247 9364 20256
rect 9312 20213 9321 20247
rect 9321 20213 9355 20247
rect 9355 20213 9364 20247
rect 9312 20204 9364 20213
rect 11888 20204 11940 20256
rect 12808 20204 12860 20256
rect 14740 20204 14792 20256
rect 16120 20315 16172 20324
rect 16120 20281 16129 20315
rect 16129 20281 16163 20315
rect 16163 20281 16172 20315
rect 16120 20272 16172 20281
rect 17224 20272 17276 20324
rect 18236 20272 18288 20324
rect 18696 20272 18748 20324
rect 18604 20204 18656 20256
rect 19524 20340 19576 20392
rect 21364 20408 21416 20460
rect 21640 20408 21692 20460
rect 23480 20408 23532 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 25412 20408 25464 20460
rect 19984 20383 20036 20392
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 20076 20272 20128 20324
rect 21272 20272 21324 20324
rect 21732 20315 21784 20324
rect 21732 20281 21741 20315
rect 21741 20281 21775 20315
rect 21775 20281 21784 20315
rect 21732 20272 21784 20281
rect 21824 20272 21876 20324
rect 24032 20383 24084 20392
rect 24032 20349 24041 20383
rect 24041 20349 24075 20383
rect 24075 20349 24084 20383
rect 24032 20340 24084 20349
rect 26240 20383 26292 20392
rect 26240 20349 26249 20383
rect 26249 20349 26283 20383
rect 26283 20349 26292 20383
rect 26240 20340 26292 20349
rect 24676 20272 24728 20324
rect 26056 20272 26108 20324
rect 26516 20340 26568 20392
rect 27160 20408 27212 20460
rect 26884 20383 26936 20392
rect 26884 20349 26893 20383
rect 26893 20349 26927 20383
rect 26927 20349 26936 20383
rect 26884 20340 26936 20349
rect 26976 20272 27028 20324
rect 27344 20383 27396 20392
rect 27344 20349 27353 20383
rect 27353 20349 27387 20383
rect 27387 20349 27396 20383
rect 27344 20340 27396 20349
rect 28448 20544 28500 20596
rect 28724 20587 28776 20596
rect 28724 20553 28733 20587
rect 28733 20553 28767 20587
rect 28767 20553 28776 20587
rect 28724 20544 28776 20553
rect 28816 20544 28868 20596
rect 30288 20544 30340 20596
rect 27620 20383 27672 20392
rect 27620 20349 27655 20383
rect 27655 20349 27672 20383
rect 27620 20340 27672 20349
rect 28264 20340 28316 20392
rect 28448 20340 28500 20392
rect 28908 20408 28960 20460
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 30380 20476 30432 20528
rect 28724 20340 28776 20392
rect 30564 20340 30616 20392
rect 30840 20383 30892 20392
rect 30840 20349 30849 20383
rect 30849 20349 30883 20383
rect 30883 20349 30892 20383
rect 30840 20340 30892 20349
rect 19984 20204 20036 20256
rect 22744 20204 22796 20256
rect 26792 20204 26844 20256
rect 27344 20204 27396 20256
rect 29276 20315 29328 20324
rect 29276 20281 29285 20315
rect 29285 20281 29319 20315
rect 29319 20281 29328 20315
rect 29276 20272 29328 20281
rect 27528 20204 27580 20256
rect 29000 20204 29052 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 12096 20102 12148 20154
rect 12160 20102 12212 20154
rect 12224 20102 12276 20154
rect 12288 20102 12340 20154
rect 12352 20102 12404 20154
rect 19870 20102 19922 20154
rect 19934 20102 19986 20154
rect 19998 20102 20050 20154
rect 20062 20102 20114 20154
rect 20126 20102 20178 20154
rect 27644 20102 27696 20154
rect 27708 20102 27760 20154
rect 27772 20102 27824 20154
rect 27836 20102 27888 20154
rect 27900 20102 27952 20154
rect 7196 20000 7248 20052
rect 7196 19907 7248 19916
rect 7196 19873 7205 19907
rect 7205 19873 7239 19907
rect 7239 19873 7248 19907
rect 7196 19864 7248 19873
rect 11060 20000 11112 20052
rect 9220 19932 9272 19984
rect 9588 19932 9640 19984
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 8944 19796 8996 19848
rect 10968 19932 11020 19984
rect 12348 20000 12400 20052
rect 12440 20043 12492 20052
rect 12440 20009 12449 20043
rect 12449 20009 12483 20043
rect 12483 20009 12492 20043
rect 12440 20000 12492 20009
rect 12532 20000 12584 20052
rect 11060 19864 11112 19916
rect 12256 19932 12308 19984
rect 14004 20000 14056 20052
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 12072 19907 12124 19916
rect 12072 19873 12081 19907
rect 12081 19873 12115 19907
rect 12115 19873 12124 19907
rect 12072 19864 12124 19873
rect 12624 19913 12676 19916
rect 12624 19879 12655 19913
rect 12655 19879 12676 19913
rect 11244 19796 11296 19848
rect 11336 19771 11388 19780
rect 8944 19703 8996 19712
rect 8944 19669 8953 19703
rect 8953 19669 8987 19703
rect 8987 19669 8996 19703
rect 8944 19660 8996 19669
rect 11336 19737 11345 19771
rect 11345 19737 11379 19771
rect 11379 19737 11388 19771
rect 11336 19728 11388 19737
rect 12624 19864 12676 19879
rect 12808 19907 12860 19916
rect 12808 19873 12817 19907
rect 12817 19873 12851 19907
rect 12851 19873 12860 19907
rect 12808 19864 12860 19873
rect 13544 19864 13596 19916
rect 13176 19796 13228 19848
rect 15568 19975 15620 19984
rect 15568 19941 15577 19975
rect 15577 19941 15611 19975
rect 15611 19941 15620 19975
rect 15568 19932 15620 19941
rect 16304 19932 16356 19984
rect 17040 20043 17092 20052
rect 17040 20009 17049 20043
rect 17049 20009 17083 20043
rect 17083 20009 17092 20043
rect 17040 20000 17092 20009
rect 17132 20000 17184 20052
rect 19432 20000 19484 20052
rect 14740 19864 14792 19916
rect 15016 19907 15068 19916
rect 15016 19873 15025 19907
rect 15025 19873 15059 19907
rect 15059 19873 15068 19907
rect 15016 19864 15068 19873
rect 18236 19932 18288 19984
rect 18420 19975 18472 19984
rect 18420 19941 18429 19975
rect 18429 19941 18463 19975
rect 18463 19941 18472 19975
rect 18420 19932 18472 19941
rect 18880 19975 18932 19984
rect 18880 19941 18889 19975
rect 18889 19941 18923 19975
rect 18923 19941 18932 19975
rect 18880 19932 18932 19941
rect 18972 19932 19024 19984
rect 17500 19907 17552 19916
rect 17500 19873 17509 19907
rect 17509 19873 17543 19907
rect 17543 19873 17552 19907
rect 17500 19864 17552 19873
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 13452 19728 13504 19780
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 16580 19839 16632 19848
rect 16580 19805 16589 19839
rect 16589 19805 16623 19839
rect 16623 19805 16632 19839
rect 16580 19796 16632 19805
rect 16672 19796 16724 19848
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 18052 19907 18104 19916
rect 18052 19873 18061 19907
rect 18061 19873 18095 19907
rect 18095 19873 18104 19907
rect 18052 19864 18104 19873
rect 19524 19932 19576 19984
rect 20260 20000 20312 20052
rect 21180 20000 21232 20052
rect 23480 20000 23532 20052
rect 23940 20000 23992 20052
rect 26884 20000 26936 20052
rect 26976 20000 27028 20052
rect 28540 20000 28592 20052
rect 28816 20000 28868 20052
rect 28908 20000 28960 20052
rect 21272 19932 21324 19984
rect 21640 19975 21692 19984
rect 21640 19941 21649 19975
rect 21649 19941 21683 19975
rect 21683 19941 21692 19975
rect 21640 19932 21692 19941
rect 22928 19932 22980 19984
rect 23296 19932 23348 19984
rect 23756 19932 23808 19984
rect 24124 19932 24176 19984
rect 24860 19932 24912 19984
rect 29276 20000 29328 20052
rect 29828 20000 29880 20052
rect 29460 19932 29512 19984
rect 31760 20000 31812 20052
rect 30288 19932 30340 19984
rect 26332 19864 26384 19916
rect 27988 19864 28040 19916
rect 28540 19907 28592 19916
rect 28540 19873 28549 19907
rect 28549 19873 28583 19907
rect 28583 19873 28592 19907
rect 28540 19864 28592 19873
rect 18328 19771 18380 19780
rect 18328 19737 18337 19771
rect 18337 19737 18371 19771
rect 18371 19737 18380 19771
rect 18328 19728 18380 19737
rect 9496 19660 9548 19712
rect 12900 19660 12952 19712
rect 13360 19660 13412 19712
rect 13912 19703 13964 19712
rect 13912 19669 13921 19703
rect 13921 19669 13955 19703
rect 13955 19669 13964 19703
rect 13912 19660 13964 19669
rect 15752 19703 15804 19712
rect 15752 19669 15761 19703
rect 15761 19669 15795 19703
rect 15795 19669 15804 19703
rect 15752 19660 15804 19669
rect 16028 19660 16080 19712
rect 16396 19660 16448 19712
rect 18696 19660 18748 19712
rect 19064 19703 19116 19712
rect 19064 19669 19073 19703
rect 19073 19669 19107 19703
rect 19107 19669 19116 19703
rect 19064 19660 19116 19669
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24400 19796 24452 19848
rect 19340 19728 19392 19780
rect 20812 19728 20864 19780
rect 20996 19660 21048 19712
rect 21824 19728 21876 19780
rect 23572 19728 23624 19780
rect 25044 19728 25096 19780
rect 26700 19839 26752 19848
rect 26700 19805 26709 19839
rect 26709 19805 26743 19839
rect 26743 19805 26752 19839
rect 26700 19796 26752 19805
rect 26792 19796 26844 19848
rect 28172 19796 28224 19848
rect 28356 19796 28408 19848
rect 21548 19660 21600 19712
rect 22100 19660 22152 19712
rect 24216 19660 24268 19712
rect 25688 19660 25740 19712
rect 26240 19660 26292 19712
rect 28448 19728 28500 19780
rect 28540 19728 28592 19780
rect 29368 19907 29420 19916
rect 29368 19873 29377 19907
rect 29377 19873 29411 19907
rect 29411 19873 29420 19907
rect 29368 19864 29420 19873
rect 29644 19796 29696 19848
rect 29460 19728 29512 19780
rect 29920 19907 29972 19916
rect 29920 19873 29929 19907
rect 29929 19873 29963 19907
rect 29963 19873 29972 19907
rect 29920 19864 29972 19873
rect 30472 19796 30524 19848
rect 31300 19907 31352 19916
rect 31300 19873 31309 19907
rect 31309 19873 31343 19907
rect 31343 19873 31352 19907
rect 31300 19864 31352 19873
rect 30656 19728 30708 19780
rect 27804 19660 27856 19712
rect 28264 19660 28316 19712
rect 28632 19660 28684 19712
rect 28816 19703 28868 19712
rect 28816 19669 28825 19703
rect 28825 19669 28859 19703
rect 28859 19669 28868 19703
rect 28816 19660 28868 19669
rect 29276 19660 29328 19712
rect 29736 19660 29788 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 11436 19558 11488 19610
rect 11500 19558 11552 19610
rect 11564 19558 11616 19610
rect 11628 19558 11680 19610
rect 11692 19558 11744 19610
rect 19210 19558 19262 19610
rect 19274 19558 19326 19610
rect 19338 19558 19390 19610
rect 19402 19558 19454 19610
rect 19466 19558 19518 19610
rect 26984 19558 27036 19610
rect 27048 19558 27100 19610
rect 27112 19558 27164 19610
rect 27176 19558 27228 19610
rect 27240 19558 27292 19610
rect 7472 19456 7524 19508
rect 8944 19456 8996 19508
rect 10600 19456 10652 19508
rect 11060 19456 11112 19508
rect 12072 19456 12124 19508
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 12808 19388 12860 19440
rect 9312 19320 9364 19372
rect 11336 19320 11388 19372
rect 5448 19252 5500 19304
rect 8484 19252 8536 19304
rect 3884 19184 3936 19236
rect 9036 19184 9088 19236
rect 10048 19184 10100 19236
rect 12072 19184 12124 19236
rect 12440 19295 12492 19304
rect 12440 19261 12449 19295
rect 12449 19261 12483 19295
rect 12483 19261 12492 19295
rect 12440 19252 12492 19261
rect 13268 19320 13320 19372
rect 12992 19184 13044 19236
rect 3424 19116 3476 19168
rect 6276 19116 6328 19168
rect 6368 19159 6420 19168
rect 6368 19125 6377 19159
rect 6377 19125 6411 19159
rect 6411 19125 6420 19159
rect 6368 19116 6420 19125
rect 6828 19116 6880 19168
rect 9220 19116 9272 19168
rect 14096 19456 14148 19508
rect 16580 19456 16632 19508
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 17500 19499 17552 19508
rect 17500 19465 17509 19499
rect 17509 19465 17543 19499
rect 17543 19465 17552 19499
rect 17500 19456 17552 19465
rect 18604 19456 18656 19508
rect 20444 19456 20496 19508
rect 21732 19456 21784 19508
rect 23848 19499 23900 19508
rect 23848 19465 23857 19499
rect 23857 19465 23891 19499
rect 23891 19465 23900 19499
rect 23848 19456 23900 19465
rect 24032 19456 24084 19508
rect 13636 19388 13688 19440
rect 18328 19388 18380 19440
rect 20352 19388 20404 19440
rect 21640 19388 21692 19440
rect 25412 19499 25464 19508
rect 25412 19465 25421 19499
rect 25421 19465 25455 19499
rect 25455 19465 25464 19499
rect 25412 19456 25464 19465
rect 26700 19456 26752 19508
rect 28724 19456 28776 19508
rect 28816 19456 28868 19508
rect 30012 19456 30064 19508
rect 13728 19320 13780 19372
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 13636 19295 13688 19304
rect 13636 19261 13646 19295
rect 13646 19261 13680 19295
rect 13680 19261 13688 19295
rect 13636 19252 13688 19261
rect 14096 19252 14148 19304
rect 14740 19320 14792 19372
rect 18420 19320 18472 19372
rect 21916 19320 21968 19372
rect 13452 19184 13504 19236
rect 13728 19184 13780 19236
rect 15568 19184 15620 19236
rect 16396 19252 16448 19304
rect 16672 19252 16724 19304
rect 17592 19295 17644 19304
rect 17592 19261 17601 19295
rect 17601 19261 17635 19295
rect 17635 19261 17644 19295
rect 17592 19252 17644 19261
rect 20352 19252 20404 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 20720 19295 20772 19304
rect 20720 19261 20729 19295
rect 20729 19261 20763 19295
rect 20763 19261 20772 19295
rect 20720 19252 20772 19261
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 20904 19295 20956 19304
rect 20904 19261 20913 19295
rect 20913 19261 20947 19295
rect 20947 19261 20956 19295
rect 20904 19252 20956 19261
rect 21456 19252 21508 19304
rect 23756 19252 23808 19304
rect 23848 19252 23900 19304
rect 24216 19252 24268 19304
rect 24400 19295 24452 19304
rect 24400 19261 24418 19295
rect 24418 19261 24452 19295
rect 24400 19252 24452 19261
rect 24860 19295 24912 19304
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 25044 19295 25096 19304
rect 25044 19261 25053 19295
rect 25053 19261 25087 19295
rect 25087 19261 25096 19295
rect 25044 19252 25096 19261
rect 25228 19252 25280 19304
rect 25412 19252 25464 19304
rect 28264 19388 28316 19440
rect 28908 19388 28960 19440
rect 27804 19320 27856 19372
rect 27988 19320 28040 19372
rect 25688 19295 25740 19304
rect 25688 19261 25697 19295
rect 25697 19261 25731 19295
rect 25731 19261 25740 19295
rect 25688 19252 25740 19261
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 25964 19252 26016 19304
rect 26332 19295 26384 19304
rect 26332 19261 26341 19295
rect 26341 19261 26375 19295
rect 26375 19261 26384 19295
rect 26332 19252 26384 19261
rect 18052 19227 18104 19236
rect 18052 19193 18061 19227
rect 18061 19193 18095 19227
rect 18095 19193 18104 19227
rect 18052 19184 18104 19193
rect 18512 19184 18564 19236
rect 18788 19184 18840 19236
rect 19800 19184 19852 19236
rect 21364 19184 21416 19236
rect 21640 19227 21692 19236
rect 21640 19193 21649 19227
rect 21649 19193 21683 19227
rect 21683 19193 21692 19227
rect 21640 19184 21692 19193
rect 22836 19184 22888 19236
rect 23112 19184 23164 19236
rect 24124 19184 24176 19236
rect 24768 19184 24820 19236
rect 26240 19184 26292 19236
rect 26792 19184 26844 19236
rect 29000 19295 29052 19304
rect 29000 19261 29009 19295
rect 29009 19261 29043 19295
rect 29043 19261 29052 19295
rect 29000 19252 29052 19261
rect 30564 19252 30616 19304
rect 15108 19116 15160 19168
rect 19616 19116 19668 19168
rect 20260 19116 20312 19168
rect 21088 19116 21140 19168
rect 22100 19116 22152 19168
rect 24952 19116 25004 19168
rect 25320 19159 25372 19168
rect 25320 19125 25329 19159
rect 25329 19125 25363 19159
rect 25363 19125 25372 19159
rect 25320 19116 25372 19125
rect 27344 19184 27396 19236
rect 27528 19116 27580 19168
rect 27620 19116 27672 19168
rect 28816 19116 28868 19168
rect 29276 19227 29328 19236
rect 29276 19193 29285 19227
rect 29285 19193 29319 19227
rect 29319 19193 29328 19227
rect 29276 19184 29328 19193
rect 31024 19227 31076 19236
rect 31024 19193 31033 19227
rect 31033 19193 31067 19227
rect 31067 19193 31076 19227
rect 31024 19184 31076 19193
rect 31116 19184 31168 19236
rect 30748 19159 30800 19168
rect 30748 19125 30757 19159
rect 30757 19125 30791 19159
rect 30791 19125 30800 19159
rect 30748 19116 30800 19125
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 12096 19014 12148 19066
rect 12160 19014 12212 19066
rect 12224 19014 12276 19066
rect 12288 19014 12340 19066
rect 12352 19014 12404 19066
rect 19870 19014 19922 19066
rect 19934 19014 19986 19066
rect 19998 19014 20050 19066
rect 20062 19014 20114 19066
rect 20126 19014 20178 19066
rect 27644 19014 27696 19066
rect 27708 19014 27760 19066
rect 27772 19014 27824 19066
rect 27836 19014 27888 19066
rect 27900 19014 27952 19066
rect 5448 18912 5500 18964
rect 3424 18776 3476 18828
rect 3240 18683 3292 18692
rect 3240 18649 3249 18683
rect 3249 18649 3283 18683
rect 3283 18649 3292 18683
rect 3240 18640 3292 18649
rect 3884 18819 3936 18828
rect 3884 18785 3893 18819
rect 3893 18785 3927 18819
rect 3927 18785 3936 18819
rect 3884 18776 3936 18785
rect 4068 18844 4120 18896
rect 4896 18776 4948 18828
rect 6092 18844 6144 18896
rect 5264 18819 5316 18828
rect 5264 18785 5273 18819
rect 5273 18785 5307 18819
rect 5307 18785 5316 18819
rect 5264 18776 5316 18785
rect 5356 18776 5408 18828
rect 6000 18708 6052 18760
rect 6184 18819 6236 18828
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 6460 18708 6512 18760
rect 7012 18776 7064 18828
rect 11244 18844 11296 18896
rect 12440 18912 12492 18964
rect 13636 18912 13688 18964
rect 16672 18955 16724 18964
rect 7104 18708 7156 18760
rect 7380 18708 7432 18760
rect 3516 18572 3568 18624
rect 5908 18683 5960 18692
rect 5908 18649 5917 18683
rect 5917 18649 5951 18683
rect 5951 18649 5960 18683
rect 5908 18640 5960 18649
rect 6828 18640 6880 18692
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 8576 18819 8628 18828
rect 8576 18785 8585 18819
rect 8585 18785 8619 18819
rect 8619 18785 8628 18819
rect 8576 18776 8628 18785
rect 8944 18776 8996 18828
rect 9220 18819 9272 18828
rect 9220 18785 9229 18819
rect 9229 18785 9263 18819
rect 9263 18785 9272 18819
rect 9220 18776 9272 18785
rect 9312 18819 9364 18828
rect 9312 18785 9321 18819
rect 9321 18785 9355 18819
rect 9355 18785 9364 18819
rect 9312 18776 9364 18785
rect 9864 18819 9916 18828
rect 9864 18785 9873 18819
rect 9873 18785 9907 18819
rect 9907 18785 9916 18819
rect 9864 18776 9916 18785
rect 9956 18819 10008 18828
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 11060 18776 11112 18828
rect 11152 18776 11204 18828
rect 12164 18776 12216 18828
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 13452 18844 13504 18896
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 16304 18887 16356 18896
rect 16304 18853 16331 18887
rect 16331 18853 16356 18887
rect 16304 18844 16356 18853
rect 18052 18912 18104 18964
rect 18420 18912 18472 18964
rect 19616 18912 19668 18964
rect 19892 18912 19944 18964
rect 20536 18912 20588 18964
rect 20904 18912 20956 18964
rect 23112 18912 23164 18964
rect 23756 18912 23808 18964
rect 17132 18887 17184 18896
rect 17132 18853 17141 18887
rect 17141 18853 17175 18887
rect 17175 18853 17184 18887
rect 17132 18844 17184 18853
rect 18144 18844 18196 18896
rect 18788 18844 18840 18896
rect 19064 18844 19116 18896
rect 14096 18776 14148 18828
rect 14280 18776 14332 18828
rect 16580 18819 16632 18828
rect 16580 18785 16589 18819
rect 16589 18785 16623 18819
rect 16623 18785 16632 18819
rect 16580 18776 16632 18785
rect 16764 18819 16816 18828
rect 16764 18785 16773 18819
rect 16773 18785 16807 18819
rect 16807 18785 16816 18819
rect 16764 18776 16816 18785
rect 11060 18640 11112 18692
rect 11336 18640 11388 18692
rect 11796 18708 11848 18760
rect 11980 18708 12032 18760
rect 12072 18708 12124 18760
rect 14464 18708 14516 18760
rect 14556 18708 14608 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16488 18708 16540 18760
rect 18604 18708 18656 18760
rect 19248 18708 19300 18760
rect 16396 18640 16448 18692
rect 6644 18615 6696 18624
rect 6644 18581 6653 18615
rect 6653 18581 6687 18615
rect 6687 18581 6696 18615
rect 6644 18572 6696 18581
rect 7472 18572 7524 18624
rect 8944 18572 8996 18624
rect 11152 18572 11204 18624
rect 11796 18572 11848 18624
rect 12164 18572 12216 18624
rect 14740 18572 14792 18624
rect 14924 18572 14976 18624
rect 16212 18572 16264 18624
rect 16580 18572 16632 18624
rect 18512 18572 18564 18624
rect 18880 18640 18932 18692
rect 20260 18819 20312 18828
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 20352 18776 20404 18828
rect 19524 18708 19576 18760
rect 20076 18708 20128 18760
rect 19616 18640 19668 18692
rect 19984 18640 20036 18692
rect 20812 18776 20864 18828
rect 21088 18776 21140 18828
rect 21180 18708 21232 18760
rect 23296 18844 23348 18896
rect 24032 18844 24084 18896
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 25872 18912 25924 18964
rect 25228 18844 25280 18896
rect 27712 18912 27764 18964
rect 29184 18912 29236 18964
rect 29920 18912 29972 18964
rect 30012 18912 30064 18964
rect 26424 18887 26476 18896
rect 26424 18853 26433 18887
rect 26433 18853 26467 18887
rect 26467 18853 26476 18887
rect 26424 18844 26476 18853
rect 20352 18683 20404 18692
rect 20352 18649 20361 18683
rect 20361 18649 20395 18683
rect 20395 18649 20404 18683
rect 20352 18640 20404 18649
rect 21640 18640 21692 18692
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 23388 18708 23440 18760
rect 24032 18708 24084 18760
rect 24492 18708 24544 18760
rect 25044 18776 25096 18828
rect 27896 18776 27948 18828
rect 25412 18708 25464 18760
rect 25504 18751 25556 18760
rect 25504 18717 25513 18751
rect 25513 18717 25547 18751
rect 25547 18717 25556 18751
rect 25504 18708 25556 18717
rect 26424 18708 26476 18760
rect 27344 18708 27396 18760
rect 29092 18844 29144 18896
rect 29644 18844 29696 18896
rect 28080 18776 28132 18828
rect 29276 18776 29328 18828
rect 29736 18819 29788 18828
rect 29736 18785 29745 18819
rect 29745 18785 29779 18819
rect 29779 18785 29788 18819
rect 29736 18776 29788 18785
rect 30288 18819 30340 18828
rect 30288 18785 30297 18819
rect 30297 18785 30331 18819
rect 30331 18785 30340 18819
rect 30288 18776 30340 18785
rect 30748 18912 30800 18964
rect 30840 18912 30892 18964
rect 31024 18844 31076 18896
rect 20904 18572 20956 18624
rect 21456 18572 21508 18624
rect 21548 18572 21600 18624
rect 23112 18615 23164 18624
rect 23112 18581 23121 18615
rect 23121 18581 23155 18615
rect 23155 18581 23164 18615
rect 23112 18572 23164 18581
rect 24860 18640 24912 18692
rect 24952 18640 25004 18692
rect 25136 18572 25188 18624
rect 26148 18615 26200 18624
rect 26148 18581 26157 18615
rect 26157 18581 26191 18615
rect 26191 18581 26200 18615
rect 26148 18572 26200 18581
rect 27528 18572 27580 18624
rect 28172 18572 28224 18624
rect 29644 18640 29696 18692
rect 29920 18708 29972 18760
rect 30104 18751 30156 18760
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 30196 18751 30248 18760
rect 30196 18717 30205 18751
rect 30205 18717 30239 18751
rect 30239 18717 30248 18751
rect 31116 18776 31168 18828
rect 30196 18708 30248 18717
rect 31024 18751 31076 18760
rect 31024 18717 31033 18751
rect 31033 18717 31067 18751
rect 31067 18717 31076 18751
rect 31024 18708 31076 18717
rect 30840 18640 30892 18692
rect 31484 18776 31536 18828
rect 31024 18572 31076 18624
rect 31300 18572 31352 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 11436 18470 11488 18522
rect 11500 18470 11552 18522
rect 11564 18470 11616 18522
rect 11628 18470 11680 18522
rect 11692 18470 11744 18522
rect 19210 18470 19262 18522
rect 19274 18470 19326 18522
rect 19338 18470 19390 18522
rect 19402 18470 19454 18522
rect 19466 18470 19518 18522
rect 26984 18470 27036 18522
rect 27048 18470 27100 18522
rect 27112 18470 27164 18522
rect 27176 18470 27228 18522
rect 27240 18470 27292 18522
rect 2504 18368 2556 18420
rect 5816 18368 5868 18420
rect 7472 18368 7524 18420
rect 8024 18368 8076 18420
rect 8668 18368 8720 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 6828 18300 6880 18352
rect 15384 18368 15436 18420
rect 16764 18368 16816 18420
rect 17224 18368 17276 18420
rect 17868 18368 17920 18420
rect 2412 18232 2464 18284
rect 4068 18232 4120 18284
rect 5172 18232 5224 18284
rect 6276 18232 6328 18284
rect 1952 18164 2004 18216
rect 2136 18164 2188 18216
rect 1768 18139 1820 18148
rect 1768 18105 1777 18139
rect 1777 18105 1811 18139
rect 1811 18105 1820 18139
rect 1768 18096 1820 18105
rect 2412 18139 2464 18148
rect 2412 18105 2421 18139
rect 2421 18105 2455 18139
rect 2455 18105 2464 18139
rect 2412 18096 2464 18105
rect 2044 18028 2096 18080
rect 3976 18164 4028 18216
rect 4712 18164 4764 18216
rect 3792 18096 3844 18148
rect 5264 18096 5316 18148
rect 6184 18207 6236 18216
rect 6184 18173 6193 18207
rect 6193 18173 6227 18207
rect 6227 18173 6236 18207
rect 6184 18164 6236 18173
rect 12072 18232 12124 18284
rect 12624 18300 12676 18352
rect 14372 18300 14424 18352
rect 6644 18207 6696 18216
rect 6644 18173 6653 18207
rect 6653 18173 6687 18207
rect 6687 18173 6696 18207
rect 6644 18164 6696 18173
rect 8484 18164 8536 18216
rect 8852 18164 8904 18216
rect 4252 18028 4304 18080
rect 5356 18028 5408 18080
rect 6276 18028 6328 18080
rect 7012 18096 7064 18148
rect 7288 18139 7340 18148
rect 7288 18105 7297 18139
rect 7297 18105 7331 18139
rect 7331 18105 7340 18139
rect 7288 18096 7340 18105
rect 7380 18139 7432 18148
rect 7380 18105 7389 18139
rect 7389 18105 7423 18139
rect 7423 18105 7432 18139
rect 7380 18096 7432 18105
rect 7564 18139 7616 18148
rect 7564 18105 7573 18139
rect 7573 18105 7607 18139
rect 7607 18105 7616 18139
rect 7564 18096 7616 18105
rect 8300 18096 8352 18148
rect 10140 18207 10192 18216
rect 10140 18173 10149 18207
rect 10149 18173 10183 18207
rect 10183 18173 10192 18207
rect 10140 18164 10192 18173
rect 10324 18164 10376 18216
rect 11796 18164 11848 18216
rect 10508 18096 10560 18148
rect 10600 18139 10652 18148
rect 10600 18105 10609 18139
rect 10609 18105 10643 18139
rect 10643 18105 10652 18139
rect 10600 18096 10652 18105
rect 11060 18139 11112 18148
rect 11060 18105 11069 18139
rect 11069 18105 11103 18139
rect 11103 18105 11112 18139
rect 11060 18096 11112 18105
rect 11152 18096 11204 18148
rect 7104 18028 7156 18080
rect 8392 18028 8444 18080
rect 9220 18028 9272 18080
rect 11244 18071 11296 18080
rect 12624 18096 12676 18148
rect 12808 18096 12860 18148
rect 13636 18164 13688 18216
rect 13820 18164 13872 18216
rect 14096 18232 14148 18284
rect 14648 18275 14700 18284
rect 14648 18241 14657 18275
rect 14657 18241 14691 18275
rect 14691 18241 14700 18275
rect 14648 18232 14700 18241
rect 14924 18275 14976 18284
rect 14924 18241 14933 18275
rect 14933 18241 14967 18275
rect 14967 18241 14976 18275
rect 14924 18232 14976 18241
rect 14004 18207 14056 18216
rect 14004 18173 14013 18207
rect 14013 18173 14047 18207
rect 14047 18173 14056 18207
rect 14004 18164 14056 18173
rect 14372 18164 14424 18216
rect 18144 18300 18196 18352
rect 18696 18300 18748 18352
rect 19616 18368 19668 18420
rect 20260 18300 20312 18352
rect 20444 18300 20496 18352
rect 20628 18300 20680 18352
rect 16304 18232 16356 18284
rect 16396 18164 16448 18216
rect 11244 18037 11269 18071
rect 11269 18037 11296 18071
rect 11244 18028 11296 18037
rect 12256 18028 12308 18080
rect 13452 18028 13504 18080
rect 14280 18071 14332 18080
rect 14280 18037 14289 18071
rect 14289 18037 14323 18071
rect 14323 18037 14332 18071
rect 14280 18028 14332 18037
rect 15844 18028 15896 18080
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 18972 18164 19024 18216
rect 19156 18164 19208 18216
rect 19984 18164 20036 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 20812 18164 20864 18216
rect 22376 18368 22428 18420
rect 23204 18368 23256 18420
rect 23388 18368 23440 18420
rect 28448 18368 28500 18420
rect 21180 18300 21232 18352
rect 21548 18300 21600 18352
rect 21088 18232 21140 18284
rect 21824 18232 21876 18284
rect 22744 18300 22796 18352
rect 23572 18300 23624 18352
rect 24492 18300 24544 18352
rect 28264 18300 28316 18352
rect 29092 18368 29144 18420
rect 29276 18368 29328 18420
rect 29460 18368 29512 18420
rect 29736 18368 29788 18420
rect 30932 18368 30984 18420
rect 28908 18300 28960 18352
rect 17592 18096 17644 18148
rect 19524 18096 19576 18148
rect 16304 18028 16356 18080
rect 17776 18028 17828 18080
rect 19616 18028 19668 18080
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 19984 18028 20036 18080
rect 20444 18139 20496 18148
rect 20444 18105 20453 18139
rect 20453 18105 20487 18139
rect 20487 18105 20496 18139
rect 20444 18096 20496 18105
rect 20720 18028 20772 18080
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 21364 18071 21416 18080
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 21916 18096 21968 18148
rect 23296 18164 23348 18216
rect 23848 18164 23900 18216
rect 23940 18207 23992 18216
rect 23940 18173 23949 18207
rect 23949 18173 23983 18207
rect 23983 18173 23992 18207
rect 23940 18164 23992 18173
rect 24676 18275 24728 18284
rect 24676 18241 24685 18275
rect 24685 18241 24719 18275
rect 24719 18241 24728 18275
rect 24676 18232 24728 18241
rect 24400 18164 24452 18216
rect 24584 18164 24636 18216
rect 23480 18139 23532 18148
rect 23480 18105 23489 18139
rect 23489 18105 23523 18139
rect 23523 18105 23532 18139
rect 23480 18096 23532 18105
rect 24124 18096 24176 18148
rect 27528 18232 27580 18284
rect 28724 18232 28776 18284
rect 29000 18275 29052 18284
rect 29000 18241 29009 18275
rect 29009 18241 29043 18275
rect 29043 18241 29052 18275
rect 29000 18232 29052 18241
rect 30748 18343 30800 18352
rect 30748 18309 30757 18343
rect 30757 18309 30791 18343
rect 30791 18309 30800 18343
rect 30748 18300 30800 18309
rect 30012 18232 30064 18284
rect 31116 18232 31168 18284
rect 27712 18207 27764 18216
rect 27712 18173 27721 18207
rect 27721 18173 27755 18207
rect 27755 18173 27764 18207
rect 27712 18164 27764 18173
rect 27896 18164 27948 18216
rect 28264 18164 28316 18216
rect 28448 18207 28500 18216
rect 28448 18173 28457 18207
rect 28457 18173 28491 18207
rect 28491 18173 28500 18207
rect 28448 18164 28500 18173
rect 28632 18207 28684 18216
rect 28632 18173 28641 18207
rect 28641 18173 28675 18207
rect 28675 18173 28684 18207
rect 28632 18164 28684 18173
rect 25136 18096 25188 18148
rect 22100 18071 22152 18080
rect 22100 18037 22109 18071
rect 22109 18037 22143 18071
rect 22143 18037 22152 18071
rect 22100 18028 22152 18037
rect 22836 18028 22888 18080
rect 24952 18028 25004 18080
rect 25228 18028 25280 18080
rect 26332 18096 26384 18148
rect 26516 18096 26568 18148
rect 26884 18096 26936 18148
rect 29184 18096 29236 18148
rect 29276 18139 29328 18148
rect 29276 18105 29285 18139
rect 29285 18105 29319 18139
rect 29319 18105 29328 18139
rect 29276 18096 29328 18105
rect 29736 18096 29788 18148
rect 31208 18139 31260 18148
rect 31208 18105 31217 18139
rect 31217 18105 31251 18139
rect 31251 18105 31260 18139
rect 31208 18096 31260 18105
rect 25872 18028 25924 18080
rect 28540 18028 28592 18080
rect 30196 18028 30248 18080
rect 31392 18028 31444 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 12096 17926 12148 17978
rect 12160 17926 12212 17978
rect 12224 17926 12276 17978
rect 12288 17926 12340 17978
rect 12352 17926 12404 17978
rect 19870 17926 19922 17978
rect 19934 17926 19986 17978
rect 19998 17926 20050 17978
rect 20062 17926 20114 17978
rect 20126 17926 20178 17978
rect 27644 17926 27696 17978
rect 27708 17926 27760 17978
rect 27772 17926 27824 17978
rect 27836 17926 27888 17978
rect 27900 17926 27952 17978
rect 2964 17824 3016 17876
rect 2228 17799 2280 17808
rect 2228 17765 2237 17799
rect 2237 17765 2271 17799
rect 2271 17765 2280 17799
rect 2228 17756 2280 17765
rect 3792 17756 3844 17808
rect 1768 17688 1820 17740
rect 1860 17688 1912 17740
rect 2596 17731 2648 17740
rect 2596 17697 2605 17731
rect 2605 17697 2639 17731
rect 2639 17697 2648 17731
rect 2596 17688 2648 17697
rect 4068 17756 4120 17808
rect 4712 17824 4764 17876
rect 5632 17824 5684 17876
rect 6644 17824 6696 17876
rect 7472 17824 7524 17876
rect 8208 17824 8260 17876
rect 8116 17756 8168 17808
rect 9220 17824 9272 17876
rect 9128 17756 9180 17808
rect 1308 17663 1360 17672
rect 1308 17629 1317 17663
rect 1317 17629 1351 17663
rect 1351 17629 1360 17663
rect 1308 17620 1360 17629
rect 2228 17620 2280 17672
rect 2964 17552 3016 17604
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 2228 17484 2280 17536
rect 3976 17688 4028 17740
rect 4068 17620 4120 17672
rect 4252 17663 4304 17672
rect 4252 17629 4261 17663
rect 4261 17629 4295 17663
rect 4295 17629 4304 17663
rect 4252 17620 4304 17629
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 5816 17731 5868 17740
rect 5816 17697 5825 17731
rect 5825 17697 5859 17731
rect 5859 17697 5868 17731
rect 5816 17688 5868 17697
rect 6000 17688 6052 17740
rect 6828 17688 6880 17740
rect 7104 17731 7156 17740
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 6552 17620 6604 17672
rect 6920 17663 6972 17672
rect 6920 17629 6929 17663
rect 6929 17629 6963 17663
rect 6963 17629 6972 17663
rect 6920 17620 6972 17629
rect 7012 17663 7064 17672
rect 7012 17629 7021 17663
rect 7021 17629 7055 17663
rect 7055 17629 7064 17663
rect 7012 17620 7064 17629
rect 7380 17688 7432 17740
rect 7840 17688 7892 17740
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 5908 17484 5960 17536
rect 6000 17484 6052 17536
rect 6276 17527 6328 17536
rect 6276 17493 6285 17527
rect 6285 17493 6319 17527
rect 6319 17493 6328 17527
rect 6276 17484 6328 17493
rect 6460 17484 6512 17536
rect 7932 17552 7984 17604
rect 8392 17731 8444 17740
rect 8392 17697 8429 17731
rect 8429 17697 8444 17731
rect 8392 17688 8444 17697
rect 8852 17688 8904 17740
rect 10232 17824 10284 17876
rect 10416 17824 10468 17876
rect 10600 17824 10652 17876
rect 9404 17756 9456 17808
rect 9864 17756 9916 17808
rect 9588 17731 9640 17740
rect 9588 17697 9597 17731
rect 9597 17697 9631 17731
rect 9631 17697 9640 17731
rect 9588 17688 9640 17697
rect 10140 17688 10192 17740
rect 10416 17688 10468 17740
rect 11244 17688 11296 17740
rect 11796 17688 11848 17740
rect 16396 17756 16448 17808
rect 12716 17731 12768 17740
rect 12716 17697 12725 17731
rect 12725 17697 12759 17731
rect 12759 17697 12768 17731
rect 12716 17688 12768 17697
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 13084 17688 13136 17740
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 14188 17731 14240 17740
rect 14188 17697 14197 17731
rect 14197 17697 14231 17731
rect 14231 17697 14240 17731
rect 14188 17688 14240 17697
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 14648 17688 14700 17740
rect 16580 17688 16632 17740
rect 8944 17620 8996 17672
rect 10232 17620 10284 17672
rect 9220 17552 9272 17604
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 10140 17552 10192 17604
rect 12440 17552 12492 17604
rect 12624 17620 12676 17672
rect 14004 17620 14056 17672
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 15844 17620 15896 17672
rect 17684 17824 17736 17876
rect 17040 17799 17092 17808
rect 17040 17765 17049 17799
rect 17049 17765 17083 17799
rect 17083 17765 17092 17799
rect 17040 17756 17092 17765
rect 17224 17799 17276 17808
rect 17224 17765 17249 17799
rect 17249 17765 17276 17799
rect 17224 17756 17276 17765
rect 17684 17731 17736 17740
rect 17684 17697 17693 17731
rect 17693 17697 17727 17731
rect 17727 17697 17736 17731
rect 17684 17688 17736 17697
rect 19524 17824 19576 17876
rect 19892 17824 19944 17876
rect 18052 17731 18104 17740
rect 18052 17697 18061 17731
rect 18061 17697 18095 17731
rect 18095 17697 18104 17731
rect 18052 17688 18104 17697
rect 18328 17731 18380 17740
rect 18328 17697 18337 17731
rect 18337 17697 18371 17731
rect 18371 17697 18380 17731
rect 18328 17688 18380 17697
rect 18604 17688 18656 17740
rect 19616 17756 19668 17808
rect 20076 17688 20128 17740
rect 21088 17824 21140 17876
rect 21916 17824 21968 17876
rect 21456 17756 21508 17808
rect 23480 17756 23532 17808
rect 24032 17824 24084 17876
rect 24216 17824 24268 17876
rect 24400 17824 24452 17876
rect 19892 17620 19944 17672
rect 20444 17731 20496 17740
rect 20444 17697 20453 17731
rect 20453 17697 20487 17731
rect 20487 17697 20496 17731
rect 20444 17688 20496 17697
rect 20628 17731 20680 17740
rect 20628 17697 20645 17731
rect 20645 17697 20680 17731
rect 20628 17688 20680 17697
rect 20720 17731 20772 17740
rect 20720 17697 20729 17731
rect 20729 17697 20763 17731
rect 20763 17697 20772 17731
rect 20720 17688 20772 17697
rect 20352 17620 20404 17672
rect 21180 17688 21232 17740
rect 25872 17799 25924 17808
rect 25872 17765 25881 17799
rect 25881 17765 25915 17799
rect 25915 17765 25924 17799
rect 25872 17756 25924 17765
rect 14188 17552 14240 17604
rect 16212 17552 16264 17604
rect 17684 17552 17736 17604
rect 18052 17552 18104 17604
rect 7380 17484 7432 17536
rect 8116 17484 8168 17536
rect 9404 17484 9456 17536
rect 9680 17484 9732 17536
rect 10324 17484 10376 17536
rect 10600 17484 10652 17536
rect 10692 17484 10744 17536
rect 11980 17484 12032 17536
rect 12164 17484 12216 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 13084 17484 13136 17536
rect 13728 17484 13780 17536
rect 14004 17527 14056 17536
rect 14004 17493 14013 17527
rect 14013 17493 14047 17527
rect 14047 17493 14056 17527
rect 14004 17484 14056 17493
rect 14740 17484 14792 17536
rect 15752 17484 15804 17536
rect 16764 17484 16816 17536
rect 20260 17552 20312 17604
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 18972 17484 19024 17536
rect 19708 17484 19760 17536
rect 19800 17484 19852 17536
rect 23940 17620 23992 17672
rect 24400 17620 24452 17672
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 26516 17824 26568 17876
rect 26332 17756 26384 17808
rect 27988 17824 28040 17876
rect 27620 17756 27672 17808
rect 29000 17824 29052 17876
rect 25044 17620 25096 17672
rect 25136 17552 25188 17604
rect 21640 17484 21692 17536
rect 23848 17484 23900 17536
rect 24124 17484 24176 17536
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 25504 17552 25556 17604
rect 26424 17688 26476 17740
rect 28356 17756 28408 17808
rect 29644 17756 29696 17808
rect 30012 17731 30064 17740
rect 30012 17697 30021 17731
rect 30021 17697 30055 17731
rect 30055 17697 30064 17731
rect 30012 17688 30064 17697
rect 30196 17688 30248 17740
rect 25872 17620 25924 17672
rect 26148 17620 26200 17672
rect 29644 17620 29696 17672
rect 30104 17620 30156 17672
rect 26884 17552 26936 17604
rect 26424 17527 26476 17536
rect 26424 17493 26433 17527
rect 26433 17493 26467 17527
rect 26467 17493 26476 17527
rect 26424 17484 26476 17493
rect 26608 17484 26660 17536
rect 28356 17552 28408 17604
rect 28264 17527 28316 17536
rect 28264 17493 28273 17527
rect 28273 17493 28307 17527
rect 28307 17493 28316 17527
rect 28264 17484 28316 17493
rect 28632 17484 28684 17536
rect 30288 17484 30340 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 11436 17382 11488 17434
rect 11500 17382 11552 17434
rect 11564 17382 11616 17434
rect 11628 17382 11680 17434
rect 11692 17382 11744 17434
rect 19210 17382 19262 17434
rect 19274 17382 19326 17434
rect 19338 17382 19390 17434
rect 19402 17382 19454 17434
rect 19466 17382 19518 17434
rect 26984 17382 27036 17434
rect 27048 17382 27100 17434
rect 27112 17382 27164 17434
rect 27176 17382 27228 17434
rect 27240 17382 27292 17434
rect 2412 17280 2464 17332
rect 2504 17280 2556 17332
rect 3056 17212 3108 17264
rect 5264 17280 5316 17332
rect 6092 17280 6144 17332
rect 6644 17280 6696 17332
rect 6828 17280 6880 17332
rect 7012 17280 7064 17332
rect 7288 17280 7340 17332
rect 8300 17280 8352 17332
rect 8392 17280 8444 17332
rect 8760 17323 8812 17332
rect 8760 17289 8769 17323
rect 8769 17289 8803 17323
rect 8803 17289 8812 17323
rect 8760 17280 8812 17289
rect 11336 17280 11388 17332
rect 11796 17280 11848 17332
rect 14556 17280 14608 17332
rect 15568 17280 15620 17332
rect 17224 17280 17276 17332
rect 18420 17280 18472 17332
rect 19800 17280 19852 17332
rect 20628 17280 20680 17332
rect 1584 17076 1636 17128
rect 2044 17119 2096 17128
rect 2044 17085 2054 17119
rect 2054 17085 2088 17119
rect 2088 17085 2096 17119
rect 2320 17144 2372 17196
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 5448 17212 5500 17264
rect 5908 17212 5960 17264
rect 12716 17212 12768 17264
rect 13084 17212 13136 17264
rect 14188 17255 14240 17264
rect 14188 17221 14197 17255
rect 14197 17221 14231 17255
rect 14231 17221 14240 17255
rect 14188 17212 14240 17221
rect 2044 17076 2096 17085
rect 2412 17119 2464 17128
rect 2412 17085 2426 17119
rect 2426 17085 2460 17119
rect 2460 17085 2464 17119
rect 2412 17076 2464 17085
rect 3240 17076 3292 17128
rect 4160 17076 4212 17128
rect 4344 17119 4396 17128
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 5080 17076 5132 17085
rect 5632 17076 5684 17128
rect 6092 17076 6144 17128
rect 1216 16940 1268 16992
rect 2136 17008 2188 17060
rect 4712 17008 4764 17060
rect 5172 17051 5224 17060
rect 5172 17017 5181 17051
rect 5181 17017 5215 17051
rect 5215 17017 5224 17051
rect 5172 17008 5224 17017
rect 5540 17008 5592 17060
rect 6460 17008 6512 17060
rect 7196 17076 7248 17128
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 7472 17076 7524 17128
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 8760 17076 8812 17128
rect 10048 17119 10100 17128
rect 10048 17085 10057 17119
rect 10057 17085 10091 17119
rect 10091 17085 10100 17119
rect 10048 17076 10100 17085
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 8484 17008 8536 17060
rect 9588 17008 9640 17060
rect 2872 16940 2924 16992
rect 3148 16940 3200 16992
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 4988 16940 5040 16992
rect 5264 16940 5316 16992
rect 7288 16940 7340 16992
rect 7472 16940 7524 16992
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 10876 17076 10928 17128
rect 11336 17076 11388 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 11980 17144 12032 17196
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 11060 16940 11112 16992
rect 11520 16940 11572 16992
rect 12440 17008 12492 17060
rect 12716 16940 12768 16992
rect 13544 17008 13596 17060
rect 14280 17119 14332 17128
rect 14280 17085 14289 17119
rect 14289 17085 14323 17119
rect 14323 17085 14332 17119
rect 14280 17076 14332 17085
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 14556 17119 14608 17128
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 14832 17144 14884 17196
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 16764 17144 16816 17196
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15752 17076 15804 17128
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 16580 17076 16632 17128
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 18144 17255 18196 17264
rect 18144 17221 18153 17255
rect 18153 17221 18187 17255
rect 18187 17221 18196 17255
rect 18144 17212 18196 17221
rect 18052 17144 18104 17196
rect 18972 17076 19024 17128
rect 20996 17212 21048 17264
rect 19340 17076 19392 17128
rect 21640 17144 21692 17196
rect 13728 16940 13780 16992
rect 15108 17008 15160 17060
rect 15384 17008 15436 17060
rect 16764 17008 16816 17060
rect 16856 17008 16908 17060
rect 16948 16940 17000 16992
rect 17500 17008 17552 17060
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 18604 17008 18656 17060
rect 19616 17076 19668 17128
rect 19800 17076 19852 17128
rect 19984 17119 20036 17128
rect 19984 17085 19993 17119
rect 19993 17085 20027 17119
rect 20027 17085 20036 17119
rect 19984 17076 20036 17085
rect 20076 17076 20128 17128
rect 20260 17119 20312 17128
rect 20260 17085 20269 17119
rect 20269 17085 20303 17119
rect 20303 17085 20312 17119
rect 20260 17076 20312 17085
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 21732 17076 21784 17128
rect 21824 17076 21876 17128
rect 22192 17212 22244 17264
rect 23388 17280 23440 17332
rect 24032 17280 24084 17332
rect 22468 17076 22520 17128
rect 22744 17255 22796 17264
rect 22744 17221 22753 17255
rect 22753 17221 22787 17255
rect 22787 17221 22796 17255
rect 22744 17212 22796 17221
rect 23848 17212 23900 17264
rect 24768 17280 24820 17332
rect 25964 17280 26016 17332
rect 27160 17280 27212 17332
rect 27528 17280 27580 17332
rect 29276 17280 29328 17332
rect 26240 17212 26292 17264
rect 29460 17280 29512 17332
rect 30748 17280 30800 17332
rect 31116 17323 31168 17332
rect 31116 17289 31125 17323
rect 31125 17289 31159 17323
rect 31159 17289 31168 17323
rect 31116 17280 31168 17289
rect 23480 17144 23532 17196
rect 23940 17144 23992 17196
rect 24952 17144 25004 17196
rect 22744 17076 22796 17128
rect 23020 17119 23072 17128
rect 23020 17085 23029 17119
rect 23029 17085 23063 17119
rect 23063 17085 23072 17119
rect 23020 17076 23072 17085
rect 18788 16940 18840 16992
rect 19616 16940 19668 16992
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 22284 17008 22336 17060
rect 23848 17119 23900 17128
rect 23848 17085 23857 17119
rect 23857 17085 23891 17119
rect 23891 17085 23900 17119
rect 23848 17076 23900 17085
rect 24032 17119 24084 17128
rect 24032 17085 24041 17119
rect 24041 17085 24075 17119
rect 24075 17085 24084 17119
rect 24032 17076 24084 17085
rect 26056 17076 26108 17128
rect 27344 17144 27396 17196
rect 27528 17144 27580 17196
rect 27988 17144 28040 17196
rect 28448 17144 28500 17196
rect 30012 17144 30064 17196
rect 21088 16940 21140 16992
rect 21364 16940 21416 16992
rect 22008 16940 22060 16992
rect 22928 16940 22980 16992
rect 23388 17008 23440 17060
rect 23572 17051 23624 17060
rect 23572 17017 23581 17051
rect 23581 17017 23615 17051
rect 23615 17017 23624 17051
rect 23572 17008 23624 17017
rect 24676 16940 24728 16992
rect 25596 16940 25648 16992
rect 26976 17076 27028 17128
rect 26056 16940 26108 16992
rect 27344 17008 27396 17060
rect 26608 16940 26660 16992
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 27804 16940 27856 16992
rect 28448 17008 28500 17060
rect 28908 17008 28960 17060
rect 28816 16940 28868 16992
rect 29276 17119 29328 17128
rect 29276 17085 29285 17119
rect 29285 17085 29319 17119
rect 29319 17085 29328 17119
rect 29276 17076 29328 17085
rect 29184 17008 29236 17060
rect 29736 17008 29788 17060
rect 30104 17008 30156 17060
rect 30472 16940 30524 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 12096 16838 12148 16890
rect 12160 16838 12212 16890
rect 12224 16838 12276 16890
rect 12288 16838 12340 16890
rect 12352 16838 12404 16890
rect 19870 16838 19922 16890
rect 19934 16838 19986 16890
rect 19998 16838 20050 16890
rect 20062 16838 20114 16890
rect 20126 16838 20178 16890
rect 27644 16838 27696 16890
rect 27708 16838 27760 16890
rect 27772 16838 27824 16890
rect 27836 16838 27888 16890
rect 27900 16838 27952 16890
rect 1676 16736 1728 16788
rect 4988 16736 5040 16788
rect 5080 16736 5132 16788
rect 6184 16736 6236 16788
rect 6644 16736 6696 16788
rect 664 16668 716 16720
rect 4160 16668 4212 16720
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 5172 16668 5224 16720
rect 8668 16736 8720 16788
rect 11612 16736 11664 16788
rect 11980 16736 12032 16788
rect 12440 16736 12492 16788
rect 12900 16736 12952 16788
rect 13360 16779 13412 16788
rect 13360 16745 13369 16779
rect 13369 16745 13403 16779
rect 13403 16745 13412 16779
rect 13360 16736 13412 16745
rect 4988 16643 5040 16652
rect 4988 16609 4997 16643
rect 4997 16609 5031 16643
rect 5031 16609 5040 16643
rect 4988 16600 5040 16609
rect 6000 16600 6052 16652
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 6368 16643 6420 16652
rect 6368 16609 6377 16643
rect 6377 16609 6411 16643
rect 6411 16609 6420 16643
rect 6368 16600 6420 16609
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 4896 16532 4948 16584
rect 2872 16464 2924 16516
rect 3148 16464 3200 16516
rect 5540 16532 5592 16584
rect 6552 16600 6604 16652
rect 7196 16668 7248 16720
rect 8208 16711 8260 16720
rect 8208 16677 8217 16711
rect 8217 16677 8251 16711
rect 8251 16677 8260 16711
rect 8208 16668 8260 16677
rect 8024 16643 8076 16652
rect 8024 16609 8033 16643
rect 8033 16609 8067 16643
rect 8067 16609 8076 16643
rect 8024 16600 8076 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8484 16600 8536 16652
rect 10140 16668 10192 16720
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 7564 16532 7616 16584
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 11152 16600 11204 16652
rect 14924 16668 14976 16720
rect 16120 16736 16172 16788
rect 16764 16736 16816 16788
rect 18236 16736 18288 16788
rect 18420 16736 18472 16788
rect 16028 16668 16080 16720
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 13084 16600 13136 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 16396 16643 16448 16652
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 10048 16532 10100 16584
rect 11060 16532 11112 16584
rect 11336 16532 11388 16584
rect 12072 16575 12124 16584
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 4804 16396 4856 16448
rect 4988 16396 5040 16448
rect 7472 16464 7524 16516
rect 8300 16464 8352 16516
rect 10324 16464 10376 16516
rect 11704 16464 11756 16516
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 13728 16575 13780 16584
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 14372 16532 14424 16584
rect 16028 16532 16080 16584
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 17040 16600 17092 16652
rect 17500 16643 17552 16652
rect 17500 16609 17509 16643
rect 17509 16609 17543 16643
rect 17543 16609 17552 16643
rect 17500 16600 17552 16609
rect 18328 16668 18380 16720
rect 18604 16736 18656 16788
rect 19708 16736 19760 16788
rect 21088 16736 21140 16788
rect 20812 16668 20864 16720
rect 19340 16600 19392 16652
rect 19800 16600 19852 16652
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 20628 16600 20680 16652
rect 20904 16643 20956 16652
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 12348 16464 12400 16516
rect 14648 16464 14700 16516
rect 15660 16464 15712 16516
rect 18052 16532 18104 16584
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 21916 16600 21968 16652
rect 22100 16643 22152 16652
rect 22100 16609 22109 16643
rect 22109 16609 22143 16643
rect 22143 16609 22152 16643
rect 22100 16600 22152 16609
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 22560 16600 22612 16652
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 23756 16668 23808 16720
rect 24308 16668 24360 16720
rect 21732 16532 21784 16584
rect 22928 16575 22980 16584
rect 22928 16541 22937 16575
rect 22937 16541 22971 16575
rect 22971 16541 22980 16575
rect 22928 16532 22980 16541
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 23940 16600 23992 16652
rect 24492 16643 24544 16652
rect 24492 16609 24501 16643
rect 24501 16609 24535 16643
rect 24535 16609 24544 16643
rect 24492 16600 24544 16609
rect 24860 16736 24912 16788
rect 25780 16736 25832 16788
rect 25872 16779 25924 16788
rect 25872 16745 25881 16779
rect 25881 16745 25915 16779
rect 25915 16745 25924 16779
rect 25872 16736 25924 16745
rect 26792 16736 26844 16788
rect 26976 16736 27028 16788
rect 27804 16779 27856 16788
rect 27804 16745 27813 16779
rect 27813 16745 27847 16779
rect 27847 16745 27856 16779
rect 27804 16736 27856 16745
rect 24400 16532 24452 16584
rect 24952 16643 25004 16652
rect 24952 16609 24961 16643
rect 24961 16609 24995 16643
rect 24995 16609 25004 16643
rect 24952 16600 25004 16609
rect 25320 16600 25372 16652
rect 25136 16532 25188 16584
rect 17132 16464 17184 16516
rect 17960 16464 18012 16516
rect 19800 16464 19852 16516
rect 20628 16464 20680 16516
rect 22560 16464 22612 16516
rect 22836 16464 22888 16516
rect 23848 16464 23900 16516
rect 24216 16464 24268 16516
rect 6828 16396 6880 16448
rect 10232 16396 10284 16448
rect 11060 16396 11112 16448
rect 11888 16396 11940 16448
rect 11980 16396 12032 16448
rect 14280 16396 14332 16448
rect 15936 16396 15988 16448
rect 16396 16396 16448 16448
rect 20904 16396 20956 16448
rect 21364 16396 21416 16448
rect 22468 16396 22520 16448
rect 23112 16396 23164 16448
rect 23388 16396 23440 16448
rect 23480 16396 23532 16448
rect 25596 16464 25648 16516
rect 26424 16600 26476 16652
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 26516 16600 26568 16609
rect 26332 16532 26384 16584
rect 26792 16643 26844 16652
rect 26792 16609 26801 16643
rect 26801 16609 26835 16643
rect 26835 16609 26844 16643
rect 26792 16600 26844 16609
rect 28724 16736 28776 16788
rect 28816 16779 28868 16788
rect 28816 16745 28825 16779
rect 28825 16745 28859 16779
rect 28859 16745 28868 16779
rect 28816 16736 28868 16745
rect 28908 16736 28960 16788
rect 31024 16736 31076 16788
rect 28080 16668 28132 16720
rect 29552 16668 29604 16720
rect 28172 16600 28224 16652
rect 28356 16600 28408 16652
rect 27160 16532 27212 16584
rect 27804 16532 27856 16584
rect 27988 16532 28040 16584
rect 26976 16464 27028 16516
rect 28080 16464 28132 16516
rect 29736 16643 29788 16652
rect 29736 16609 29745 16643
rect 29745 16609 29779 16643
rect 29779 16609 29788 16643
rect 29736 16600 29788 16609
rect 29460 16532 29512 16584
rect 30288 16600 30340 16652
rect 30472 16600 30524 16652
rect 31116 16643 31168 16652
rect 31116 16609 31125 16643
rect 31125 16609 31159 16643
rect 31159 16609 31168 16643
rect 31116 16600 31168 16609
rect 30012 16532 30064 16584
rect 26332 16396 26384 16448
rect 26792 16396 26844 16448
rect 27068 16396 27120 16448
rect 27896 16396 27948 16448
rect 29000 16464 29052 16516
rect 28448 16396 28500 16448
rect 29184 16396 29236 16448
rect 29552 16396 29604 16448
rect 31300 16464 31352 16516
rect 31208 16439 31260 16448
rect 31208 16405 31217 16439
rect 31217 16405 31251 16439
rect 31251 16405 31260 16439
rect 31208 16396 31260 16405
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 11436 16294 11488 16346
rect 11500 16294 11552 16346
rect 11564 16294 11616 16346
rect 11628 16294 11680 16346
rect 11692 16294 11744 16346
rect 19210 16294 19262 16346
rect 19274 16294 19326 16346
rect 19338 16294 19390 16346
rect 19402 16294 19454 16346
rect 19466 16294 19518 16346
rect 26984 16294 27036 16346
rect 27048 16294 27100 16346
rect 27112 16294 27164 16346
rect 27176 16294 27228 16346
rect 27240 16294 27292 16346
rect 2136 16192 2188 16244
rect 2412 16192 2464 16244
rect 3516 16192 3568 16244
rect 5264 16192 5316 16244
rect 6368 16192 6420 16244
rect 7104 16192 7156 16244
rect 10048 16192 10100 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 11336 16192 11388 16244
rect 11612 16192 11664 16244
rect 11888 16192 11940 16244
rect 572 16124 624 16176
rect 1952 16124 2004 16176
rect 1308 15988 1360 16040
rect 1492 15988 1544 16040
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 2228 16124 2280 16176
rect 2320 15988 2372 16040
rect 3516 16056 3568 16108
rect 2596 15988 2648 16040
rect 4252 16031 4304 16040
rect 4252 15997 4261 16031
rect 4261 15997 4295 16031
rect 4295 15997 4304 16031
rect 4252 15988 4304 15997
rect 4988 16031 5040 16040
rect 4988 15997 4997 16031
rect 4997 15997 5031 16031
rect 5031 15997 5040 16031
rect 4988 15988 5040 15997
rect 6000 15988 6052 16040
rect 6920 16056 6972 16108
rect 7012 16056 7064 16108
rect 7196 15988 7248 16040
rect 8116 16056 8168 16108
rect 1492 15852 1544 15904
rect 1768 15852 1820 15904
rect 2228 15852 2280 15904
rect 2596 15852 2648 15904
rect 5632 15920 5684 15972
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 8208 15988 8260 16040
rect 8300 15988 8352 16040
rect 7932 15920 7984 15972
rect 8576 15920 8628 15972
rect 12072 16167 12124 16176
rect 12072 16133 12081 16167
rect 12081 16133 12115 16167
rect 12115 16133 12124 16167
rect 12072 16124 12124 16133
rect 9312 16056 9364 16108
rect 8944 15988 8996 16040
rect 9496 15963 9548 15972
rect 9496 15929 9505 15963
rect 9505 15929 9539 15963
rect 9539 15929 9548 15963
rect 9496 15920 9548 15929
rect 10048 15988 10100 16040
rect 11336 15988 11388 16040
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 12440 16056 12492 16108
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 14280 16235 14332 16244
rect 14280 16201 14289 16235
rect 14289 16201 14323 16235
rect 14323 16201 14332 16235
rect 14280 16192 14332 16201
rect 14464 16235 14516 16244
rect 14464 16201 14473 16235
rect 14473 16201 14507 16235
rect 14507 16201 14516 16235
rect 14464 16192 14516 16201
rect 15016 16192 15068 16244
rect 12532 15988 12584 16040
rect 12624 16031 12676 16040
rect 12624 15997 12633 16031
rect 12633 15997 12667 16031
rect 12667 15997 12676 16031
rect 12624 15988 12676 15997
rect 5540 15852 5592 15904
rect 6000 15852 6052 15904
rect 7472 15852 7524 15904
rect 7656 15852 7708 15904
rect 9036 15852 9088 15904
rect 10140 15852 10192 15904
rect 10876 15920 10928 15972
rect 12072 15920 12124 15972
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 16028 16124 16080 16176
rect 19800 16192 19852 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 20260 16192 20312 16244
rect 22100 16235 22152 16244
rect 22100 16201 22109 16235
rect 22109 16201 22143 16235
rect 22143 16201 22152 16235
rect 22100 16192 22152 16201
rect 22192 16192 22244 16244
rect 22560 16192 22612 16244
rect 23020 16192 23072 16244
rect 23204 16192 23256 16244
rect 23388 16192 23440 16244
rect 25044 16192 25096 16244
rect 26240 16235 26292 16244
rect 26240 16201 26249 16235
rect 26249 16201 26283 16235
rect 26283 16201 26292 16235
rect 26240 16192 26292 16201
rect 26516 16192 26568 16244
rect 28724 16192 28776 16244
rect 29828 16192 29880 16244
rect 15936 16056 15988 16108
rect 12164 15852 12216 15904
rect 12992 15963 13044 15972
rect 12992 15929 13001 15963
rect 13001 15929 13035 15963
rect 13035 15929 13044 15963
rect 12992 15920 13044 15929
rect 13636 15920 13688 15972
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 16488 15988 16540 16040
rect 18696 16056 18748 16108
rect 19248 16056 19300 16108
rect 19800 16056 19852 16108
rect 12440 15852 12492 15904
rect 13820 15852 13872 15904
rect 14004 15852 14056 15904
rect 16120 15920 16172 15972
rect 17040 15920 17092 15972
rect 18604 15920 18656 15972
rect 19248 15963 19300 15972
rect 19248 15929 19257 15963
rect 19257 15929 19291 15963
rect 19291 15929 19300 15963
rect 19248 15920 19300 15929
rect 19432 15963 19484 15972
rect 19432 15929 19457 15963
rect 19457 15929 19484 15963
rect 19432 15920 19484 15929
rect 21180 15988 21232 16040
rect 21456 16031 21508 16040
rect 21456 15997 21465 16031
rect 21465 15997 21499 16031
rect 21499 15997 21508 16031
rect 21456 15988 21508 15997
rect 21548 16031 21600 16040
rect 21548 15997 21557 16031
rect 21557 15997 21591 16031
rect 21591 15997 21600 16031
rect 21548 15988 21600 15997
rect 21732 16031 21784 16040
rect 21732 15997 21741 16031
rect 21741 15997 21775 16031
rect 21775 15997 21784 16031
rect 21732 15988 21784 15997
rect 22468 16056 22520 16108
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 15384 15852 15436 15904
rect 15568 15852 15620 15904
rect 19340 15852 19392 15904
rect 22008 15920 22060 15972
rect 22100 15920 22152 15972
rect 23020 16056 23072 16108
rect 23572 16056 23624 16108
rect 23664 15988 23716 16040
rect 23756 15988 23808 16040
rect 24308 16099 24360 16108
rect 24308 16065 24317 16099
rect 24317 16065 24351 16099
rect 24351 16065 24360 16099
rect 24308 16056 24360 16065
rect 24860 16056 24912 16108
rect 25044 16056 25096 16108
rect 25688 16124 25740 16176
rect 25872 16124 25924 16176
rect 26884 16124 26936 16176
rect 27068 16124 27120 16176
rect 25964 16056 26016 16108
rect 26424 16056 26476 16108
rect 26700 16056 26752 16108
rect 27160 16056 27212 16108
rect 27528 16124 27580 16176
rect 27620 16124 27672 16176
rect 27988 16124 28040 16176
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 24216 15988 24268 16040
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 22928 15920 22980 15972
rect 20812 15852 20864 15904
rect 21640 15852 21692 15904
rect 22560 15852 22612 15904
rect 23204 15852 23256 15904
rect 23480 15852 23532 15904
rect 23572 15895 23624 15904
rect 23572 15861 23581 15895
rect 23581 15861 23615 15895
rect 23615 15861 23624 15895
rect 23572 15852 23624 15861
rect 23940 15920 23992 15972
rect 25044 15920 25096 15972
rect 26056 15988 26108 16040
rect 25688 15920 25740 15972
rect 26332 16031 26384 16040
rect 26332 15997 26341 16031
rect 26341 15997 26375 16031
rect 26375 15997 26384 16031
rect 26332 15988 26384 15997
rect 26884 15988 26936 16040
rect 27804 15988 27856 16040
rect 28264 16056 28316 16108
rect 29184 16124 29236 16176
rect 29552 16099 29604 16108
rect 28632 16031 28684 16040
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 28632 15997 28671 16031
rect 28671 15997 28684 16031
rect 28632 15988 28684 15997
rect 28908 15988 28960 16040
rect 30380 16031 30432 16040
rect 30380 15997 30389 16031
rect 30389 15997 30423 16031
rect 30423 15997 30432 16031
rect 30380 15988 30432 15997
rect 30932 16031 30984 16040
rect 30932 15997 30941 16031
rect 30941 15997 30975 16031
rect 30975 15997 30984 16031
rect 30932 15988 30984 15997
rect 31116 16031 31168 16040
rect 31116 15997 31125 16031
rect 31125 15997 31159 16031
rect 31159 15997 31168 16031
rect 31116 15988 31168 15997
rect 31392 15988 31444 16040
rect 26884 15895 26936 15904
rect 26884 15861 26893 15895
rect 26893 15861 26927 15895
rect 26927 15861 26936 15895
rect 26884 15852 26936 15861
rect 27160 15852 27212 15904
rect 29460 15920 29512 15972
rect 30196 15963 30248 15972
rect 30196 15929 30205 15963
rect 30205 15929 30239 15963
rect 30239 15929 30248 15963
rect 30196 15920 30248 15929
rect 28632 15852 28684 15904
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 12096 15750 12148 15802
rect 12160 15750 12212 15802
rect 12224 15750 12276 15802
rect 12288 15750 12340 15802
rect 12352 15750 12404 15802
rect 19870 15750 19922 15802
rect 19934 15750 19986 15802
rect 19998 15750 20050 15802
rect 20062 15750 20114 15802
rect 20126 15750 20178 15802
rect 27644 15750 27696 15802
rect 27708 15750 27760 15802
rect 27772 15750 27824 15802
rect 27836 15750 27888 15802
rect 27900 15750 27952 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 4068 15648 4120 15700
rect 5448 15648 5500 15700
rect 1216 15512 1268 15564
rect 1584 15512 1636 15564
rect 3148 15555 3200 15564
rect 3148 15521 3157 15555
rect 3157 15521 3191 15555
rect 3191 15521 3200 15555
rect 3148 15512 3200 15521
rect 3240 15512 3292 15564
rect 4712 15580 4764 15632
rect 3424 15512 3476 15564
rect 2688 15444 2740 15496
rect 4068 15512 4120 15564
rect 3332 15308 3384 15360
rect 5080 15444 5132 15496
rect 5632 15555 5684 15564
rect 5632 15521 5641 15555
rect 5641 15521 5675 15555
rect 5675 15521 5684 15555
rect 5632 15512 5684 15521
rect 7472 15648 7524 15700
rect 9588 15648 9640 15700
rect 9956 15648 10008 15700
rect 11888 15648 11940 15700
rect 13544 15648 13596 15700
rect 13820 15648 13872 15700
rect 15200 15648 15252 15700
rect 15752 15648 15804 15700
rect 16488 15648 16540 15700
rect 20168 15648 20220 15700
rect 20260 15648 20312 15700
rect 20812 15648 20864 15700
rect 20904 15648 20956 15700
rect 22652 15648 22704 15700
rect 22928 15691 22980 15700
rect 22928 15657 22937 15691
rect 22937 15657 22971 15691
rect 22971 15657 22980 15691
rect 22928 15648 22980 15657
rect 7012 15580 7064 15632
rect 8484 15580 8536 15632
rect 9036 15580 9088 15632
rect 5540 15444 5592 15496
rect 6000 15444 6052 15496
rect 6828 15512 6880 15564
rect 7472 15555 7524 15564
rect 7472 15521 7481 15555
rect 7481 15521 7515 15555
rect 7515 15521 7524 15555
rect 7472 15512 7524 15521
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 8944 15444 8996 15496
rect 10876 15580 10928 15632
rect 11612 15580 11664 15632
rect 11980 15580 12032 15632
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 10232 15555 10284 15564
rect 10232 15521 10241 15555
rect 10241 15521 10275 15555
rect 10275 15521 10284 15555
rect 10232 15512 10284 15521
rect 10324 15512 10376 15564
rect 11244 15512 11296 15564
rect 12440 15580 12492 15632
rect 12532 15512 12584 15564
rect 12900 15512 12952 15564
rect 12992 15512 13044 15564
rect 13636 15512 13688 15564
rect 14556 15580 14608 15632
rect 14648 15580 14700 15632
rect 14832 15555 14884 15564
rect 14832 15521 14841 15555
rect 14841 15521 14875 15555
rect 14875 15521 14884 15555
rect 14832 15512 14884 15521
rect 15016 15623 15068 15632
rect 15016 15589 15025 15623
rect 15025 15589 15059 15623
rect 15059 15589 15068 15623
rect 15016 15580 15068 15589
rect 15568 15512 15620 15564
rect 15660 15555 15712 15564
rect 15660 15521 15669 15555
rect 15669 15521 15703 15555
rect 15703 15521 15712 15555
rect 15660 15512 15712 15521
rect 15752 15512 15804 15564
rect 10784 15444 10836 15496
rect 10876 15444 10928 15496
rect 13084 15444 13136 15496
rect 10324 15419 10376 15428
rect 10324 15385 10333 15419
rect 10333 15385 10367 15419
rect 10367 15385 10376 15419
rect 10324 15376 10376 15385
rect 10968 15376 11020 15428
rect 11060 15376 11112 15428
rect 16396 15376 16448 15428
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 16948 15555 17000 15564
rect 16948 15521 16957 15555
rect 16957 15521 16991 15555
rect 16991 15521 17000 15555
rect 16948 15512 17000 15521
rect 17776 15580 17828 15632
rect 18144 15580 18196 15632
rect 20720 15580 20772 15632
rect 17316 15444 17368 15496
rect 17684 15444 17736 15496
rect 17960 15555 18012 15564
rect 17960 15521 17969 15555
rect 17969 15521 18003 15555
rect 18003 15521 18012 15555
rect 17960 15512 18012 15521
rect 19524 15512 19576 15564
rect 20076 15512 20128 15564
rect 22376 15580 22428 15632
rect 24584 15648 24636 15700
rect 24768 15648 24820 15700
rect 21180 15512 21232 15564
rect 23480 15580 23532 15632
rect 19708 15444 19760 15496
rect 20168 15444 20220 15496
rect 23204 15512 23256 15564
rect 23756 15623 23808 15632
rect 23756 15589 23765 15623
rect 23765 15589 23799 15623
rect 23799 15589 23808 15623
rect 23756 15580 23808 15589
rect 26516 15648 26568 15700
rect 20812 15376 20864 15428
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 23940 15555 23992 15564
rect 23940 15521 23949 15555
rect 23949 15521 23983 15555
rect 23983 15521 23992 15555
rect 23940 15512 23992 15521
rect 6552 15308 6604 15360
rect 8024 15308 8076 15360
rect 8852 15308 8904 15360
rect 9588 15308 9640 15360
rect 11612 15308 11664 15360
rect 13360 15308 13412 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 13820 15308 13872 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 15752 15308 15804 15360
rect 17776 15308 17828 15360
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 19340 15308 19392 15360
rect 22836 15419 22888 15428
rect 22836 15385 22845 15419
rect 22845 15385 22879 15419
rect 22879 15385 22888 15419
rect 22836 15376 22888 15385
rect 24124 15512 24176 15564
rect 24400 15555 24452 15564
rect 24400 15521 24409 15555
rect 24409 15521 24443 15555
rect 24443 15521 24452 15555
rect 24400 15512 24452 15521
rect 24584 15512 24636 15564
rect 25596 15512 25648 15564
rect 26148 15580 26200 15632
rect 26424 15580 26476 15632
rect 27620 15648 27672 15700
rect 27896 15648 27948 15700
rect 28080 15648 28132 15700
rect 28448 15691 28500 15700
rect 28448 15657 28457 15691
rect 28457 15657 28491 15691
rect 28491 15657 28500 15691
rect 28448 15648 28500 15657
rect 29276 15648 29328 15700
rect 29552 15648 29604 15700
rect 30104 15648 30156 15700
rect 30196 15648 30248 15700
rect 26332 15512 26384 15564
rect 27160 15555 27212 15564
rect 27160 15521 27169 15555
rect 27169 15521 27203 15555
rect 27203 15521 27212 15555
rect 27160 15512 27212 15521
rect 24676 15444 24728 15496
rect 24860 15444 24912 15496
rect 25320 15444 25372 15496
rect 27620 15512 27672 15564
rect 28356 15512 28408 15564
rect 28448 15512 28500 15564
rect 31208 15580 31260 15632
rect 29184 15512 29236 15564
rect 29552 15555 29604 15564
rect 29552 15521 29561 15555
rect 29561 15521 29595 15555
rect 29595 15521 29604 15555
rect 29552 15512 29604 15521
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 30380 15512 30432 15564
rect 30840 15512 30892 15564
rect 31300 15555 31352 15564
rect 31300 15521 31309 15555
rect 31309 15521 31343 15555
rect 31343 15521 31352 15555
rect 31300 15512 31352 15521
rect 20996 15308 21048 15360
rect 23848 15308 23900 15360
rect 24308 15308 24360 15360
rect 24584 15376 24636 15428
rect 28172 15444 28224 15496
rect 28264 15444 28316 15496
rect 28632 15444 28684 15496
rect 30012 15487 30064 15496
rect 30012 15453 30018 15487
rect 30018 15453 30064 15487
rect 30012 15444 30064 15453
rect 24952 15308 25004 15360
rect 25320 15308 25372 15360
rect 28908 15376 28960 15428
rect 29552 15376 29604 15428
rect 31668 15444 31720 15496
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 26700 15308 26752 15360
rect 27160 15308 27212 15360
rect 28356 15308 28408 15360
rect 29000 15308 29052 15360
rect 29276 15308 29328 15360
rect 29736 15308 29788 15360
rect 30472 15376 30524 15428
rect 30288 15351 30340 15360
rect 30288 15317 30297 15351
rect 30297 15317 30331 15351
rect 30331 15317 30340 15351
rect 30288 15308 30340 15317
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11436 15206 11488 15258
rect 11500 15206 11552 15258
rect 11564 15206 11616 15258
rect 11628 15206 11680 15258
rect 11692 15206 11744 15258
rect 19210 15206 19262 15258
rect 19274 15206 19326 15258
rect 19338 15206 19390 15258
rect 19402 15206 19454 15258
rect 19466 15206 19518 15258
rect 26984 15206 27036 15258
rect 27048 15206 27100 15258
rect 27112 15206 27164 15258
rect 27176 15206 27228 15258
rect 27240 15206 27292 15258
rect 5448 15104 5500 15156
rect 6092 15104 6144 15156
rect 6368 15104 6420 15156
rect 3516 15036 3568 15088
rect 1216 14968 1268 15020
rect 1492 14943 1544 14952
rect 1492 14909 1501 14943
rect 1501 14909 1535 14943
rect 1535 14909 1544 14943
rect 1492 14900 1544 14909
rect 1860 14764 1912 14816
rect 3332 14943 3384 14952
rect 3332 14909 3341 14943
rect 3341 14909 3375 14943
rect 3375 14909 3384 14943
rect 3332 14900 3384 14909
rect 3608 14943 3660 14952
rect 3608 14909 3617 14943
rect 3617 14909 3651 14943
rect 3651 14909 3660 14943
rect 3608 14900 3660 14909
rect 5080 15011 5132 15020
rect 5080 14977 5089 15011
rect 5089 14977 5123 15011
rect 5123 14977 5132 15011
rect 5080 14968 5132 14977
rect 7656 15104 7708 15156
rect 8024 15079 8076 15088
rect 8024 15045 8033 15079
rect 8033 15045 8067 15079
rect 8067 15045 8076 15079
rect 8024 15036 8076 15045
rect 8576 15036 8628 15088
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 4896 14943 4948 14952
rect 4896 14909 4905 14943
rect 4905 14909 4939 14943
rect 4939 14909 4948 14943
rect 4896 14900 4948 14909
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 6920 14968 6972 15020
rect 3976 14764 4028 14816
rect 5172 14764 5224 14816
rect 5724 14900 5776 14952
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 6828 14900 6880 14952
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7012 14900 7064 14909
rect 5540 14764 5592 14816
rect 6828 14764 6880 14816
rect 7288 14968 7340 15020
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 7288 14875 7340 14884
rect 7288 14841 7297 14875
rect 7297 14841 7331 14875
rect 7331 14841 7340 14875
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 8484 14943 8536 14952
rect 8484 14909 8493 14943
rect 8493 14909 8527 14943
rect 8527 14909 8536 14943
rect 8484 14900 8536 14909
rect 8576 14900 8628 14952
rect 9220 15079 9272 15088
rect 9220 15045 9229 15079
rect 9229 15045 9263 15079
rect 9263 15045 9272 15079
rect 9220 15036 9272 15045
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 10232 15036 10284 15088
rect 11060 15036 11112 15088
rect 11244 15036 11296 15088
rect 11336 15036 11388 15088
rect 14188 15104 14240 15156
rect 14280 15104 14332 15156
rect 9956 14968 10008 15020
rect 12992 14968 13044 15020
rect 9588 14900 9640 14952
rect 10508 14900 10560 14952
rect 7288 14832 7340 14841
rect 8852 14832 8904 14884
rect 9036 14832 9088 14884
rect 9956 14832 10008 14884
rect 10876 14832 10928 14884
rect 11428 14943 11480 14952
rect 11428 14909 11437 14943
rect 11437 14909 11471 14943
rect 11471 14909 11480 14943
rect 11428 14900 11480 14909
rect 11520 14900 11572 14952
rect 12072 14900 12124 14952
rect 12164 14900 12216 14952
rect 12716 14900 12768 14952
rect 12900 14832 12952 14884
rect 13268 15036 13320 15088
rect 13452 14968 13504 15020
rect 14372 15036 14424 15088
rect 15016 15104 15068 15156
rect 21180 15104 21232 15156
rect 21640 15104 21692 15156
rect 22744 15104 22796 15156
rect 23756 15104 23808 15156
rect 24032 15104 24084 15156
rect 25320 15104 25372 15156
rect 26056 15104 26108 15156
rect 15200 15036 15252 15088
rect 14648 14968 14700 15020
rect 15292 14968 15344 15020
rect 15752 14968 15804 15020
rect 16212 14968 16264 15020
rect 16948 14968 17000 15020
rect 13268 14900 13320 14952
rect 13728 14943 13780 14952
rect 13728 14909 13737 14943
rect 13737 14909 13771 14943
rect 13771 14909 13780 14943
rect 13728 14900 13780 14909
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 14096 14943 14148 14952
rect 14096 14909 14105 14943
rect 14105 14909 14139 14943
rect 14139 14909 14148 14943
rect 14096 14900 14148 14909
rect 7656 14764 7708 14816
rect 8116 14764 8168 14816
rect 13544 14764 13596 14816
rect 14648 14832 14700 14884
rect 14924 14832 14976 14884
rect 15108 14832 15160 14884
rect 15660 14900 15712 14952
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 17408 14968 17460 15020
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 19340 14968 19392 15020
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 17592 14900 17644 14952
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 20260 14900 20312 14952
rect 14188 14764 14240 14816
rect 14280 14764 14332 14816
rect 16764 14764 16816 14816
rect 17224 14764 17276 14816
rect 19340 14764 19392 14816
rect 19892 14832 19944 14884
rect 20168 14875 20220 14884
rect 20168 14841 20177 14875
rect 20177 14841 20211 14875
rect 20211 14841 20220 14875
rect 20168 14832 20220 14841
rect 20720 14832 20772 14884
rect 21456 14968 21508 15020
rect 21824 14968 21876 15020
rect 21640 14943 21692 14952
rect 21640 14909 21649 14943
rect 21649 14909 21683 14943
rect 21683 14909 21692 14943
rect 21640 14900 21692 14909
rect 21732 14900 21784 14952
rect 22376 14900 22428 14952
rect 22652 14968 22704 15020
rect 22744 14900 22796 14952
rect 23112 14943 23164 14952
rect 23112 14909 23121 14943
rect 23121 14909 23155 14943
rect 23155 14909 23164 14943
rect 23112 14900 23164 14909
rect 21088 14832 21140 14884
rect 21456 14832 21508 14884
rect 22192 14875 22244 14884
rect 22192 14841 22201 14875
rect 22201 14841 22235 14875
rect 22235 14841 22244 14875
rect 22192 14832 22244 14841
rect 21640 14764 21692 14816
rect 21824 14764 21876 14816
rect 23020 14875 23072 14884
rect 23020 14841 23029 14875
rect 23029 14841 23063 14875
rect 23063 14841 23072 14875
rect 23020 14832 23072 14841
rect 23572 15036 23624 15088
rect 24952 14968 25004 15020
rect 25136 14968 25188 15020
rect 23388 14943 23440 14952
rect 23388 14909 23397 14943
rect 23397 14909 23431 14943
rect 23431 14909 23440 14943
rect 23388 14900 23440 14909
rect 24308 14943 24360 14952
rect 24308 14909 24317 14943
rect 24317 14909 24351 14943
rect 24351 14909 24360 14943
rect 24308 14900 24360 14909
rect 24492 14943 24544 14952
rect 24492 14909 24501 14943
rect 24501 14909 24535 14943
rect 24535 14909 24544 14943
rect 24492 14900 24544 14909
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24860 14832 24912 14884
rect 25136 14832 25188 14884
rect 25596 14832 25648 14884
rect 26332 14968 26384 15020
rect 22468 14764 22520 14816
rect 23940 14764 23992 14816
rect 25320 14764 25372 14816
rect 25412 14764 25464 14816
rect 25872 14807 25924 14816
rect 25872 14773 25881 14807
rect 25881 14773 25915 14807
rect 25915 14773 25924 14807
rect 25872 14764 25924 14773
rect 27620 15104 27672 15156
rect 29368 15104 29420 15156
rect 27436 15036 27488 15088
rect 28448 15036 28500 15088
rect 30932 15104 30984 15156
rect 31760 15104 31812 15156
rect 30288 15036 30340 15088
rect 27344 14900 27396 14952
rect 28540 14968 28592 15020
rect 26148 14764 26200 14816
rect 26240 14807 26292 14816
rect 26240 14773 26249 14807
rect 26249 14773 26283 14807
rect 26283 14773 26292 14807
rect 26240 14764 26292 14773
rect 27344 14764 27396 14816
rect 27712 14764 27764 14816
rect 28172 14900 28224 14952
rect 29276 14943 29328 14952
rect 29276 14909 29285 14943
rect 29285 14909 29319 14943
rect 29319 14909 29328 14943
rect 29276 14900 29328 14909
rect 29552 14968 29604 15020
rect 29920 14900 29972 14952
rect 30380 14900 30432 14952
rect 28356 14832 28408 14884
rect 29644 14832 29696 14884
rect 29184 14807 29236 14816
rect 29184 14773 29193 14807
rect 29193 14773 29227 14807
rect 29227 14773 29236 14807
rect 29184 14764 29236 14773
rect 29920 14764 29972 14816
rect 30380 14807 30432 14816
rect 30380 14773 30389 14807
rect 30389 14773 30423 14807
rect 30423 14773 30432 14807
rect 30380 14764 30432 14773
rect 30564 14943 30616 14952
rect 30564 14909 30573 14943
rect 30573 14909 30607 14943
rect 30607 14909 30616 14943
rect 30564 14900 30616 14909
rect 31576 14900 31628 14952
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 12096 14662 12148 14714
rect 12160 14662 12212 14714
rect 12224 14662 12276 14714
rect 12288 14662 12340 14714
rect 12352 14662 12404 14714
rect 19870 14662 19922 14714
rect 19934 14662 19986 14714
rect 19998 14662 20050 14714
rect 20062 14662 20114 14714
rect 20126 14662 20178 14714
rect 27644 14662 27696 14714
rect 27708 14662 27760 14714
rect 27772 14662 27824 14714
rect 27836 14662 27888 14714
rect 27900 14662 27952 14714
rect 3240 14560 3292 14612
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 3148 14535 3200 14544
rect 3148 14501 3157 14535
rect 3157 14501 3191 14535
rect 3191 14501 3200 14535
rect 3148 14492 3200 14501
rect 2872 14424 2924 14476
rect 3240 14424 3292 14476
rect 4160 14424 4212 14476
rect 5356 14492 5408 14544
rect 6000 14492 6052 14544
rect 6552 14560 6604 14612
rect 7012 14560 7064 14612
rect 7288 14603 7340 14612
rect 7288 14569 7290 14603
rect 7290 14569 7324 14603
rect 7324 14569 7340 14603
rect 7288 14560 7340 14569
rect 7380 14560 7432 14612
rect 8116 14492 8168 14544
rect 8760 14560 8812 14612
rect 5448 14467 5500 14476
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 1032 14288 1084 14340
rect 4068 14356 4120 14408
rect 3240 14288 3292 14340
rect 3424 14288 3476 14340
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5724 14424 5776 14476
rect 5356 14356 5408 14365
rect 5540 14288 5592 14340
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6920 14467 6972 14476
rect 6920 14433 6929 14467
rect 6929 14433 6963 14467
rect 6963 14433 6972 14467
rect 6920 14424 6972 14433
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 7104 14424 7156 14433
rect 7288 14424 7340 14476
rect 7472 14424 7524 14476
rect 8576 14424 8628 14476
rect 8760 14424 8812 14476
rect 8944 14492 8996 14544
rect 9220 14560 9272 14612
rect 10232 14560 10284 14612
rect 10784 14560 10836 14612
rect 9036 14424 9088 14476
rect 9588 14492 9640 14544
rect 10508 14492 10560 14544
rect 8116 14356 8168 14408
rect 10416 14424 10468 14476
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 10784 14467 10836 14476
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 6828 14288 6880 14340
rect 6920 14288 6972 14340
rect 7380 14288 7432 14340
rect 9588 14356 9640 14408
rect 13728 14560 13780 14612
rect 13912 14560 13964 14612
rect 14832 14603 14884 14612
rect 14832 14569 14841 14603
rect 14841 14569 14875 14603
rect 14875 14569 14884 14603
rect 14832 14560 14884 14569
rect 15292 14560 15344 14612
rect 16396 14560 16448 14612
rect 17776 14560 17828 14612
rect 17868 14560 17920 14612
rect 18236 14560 18288 14612
rect 19432 14560 19484 14612
rect 19708 14560 19760 14612
rect 19984 14560 20036 14612
rect 20812 14560 20864 14612
rect 22192 14560 22244 14612
rect 22468 14603 22520 14612
rect 22468 14569 22477 14603
rect 22477 14569 22511 14603
rect 22511 14569 22520 14603
rect 22468 14560 22520 14569
rect 11612 14424 11664 14476
rect 14280 14492 14332 14544
rect 14648 14492 14700 14544
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 9036 14331 9088 14340
rect 9036 14297 9045 14331
rect 9045 14297 9079 14331
rect 9079 14297 9088 14331
rect 9036 14288 9088 14297
rect 9496 14288 9548 14340
rect 11520 14356 11572 14408
rect 12072 14424 12124 14476
rect 12624 14424 12676 14476
rect 12256 14356 12308 14408
rect 3976 14220 4028 14272
rect 5724 14220 5776 14272
rect 6460 14220 6512 14272
rect 7472 14220 7524 14272
rect 8392 14220 8444 14272
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 12440 14288 12492 14340
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 13268 14424 13320 14476
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 14096 14424 14148 14476
rect 14924 14424 14976 14476
rect 15016 14467 15068 14476
rect 15016 14433 15025 14467
rect 15025 14433 15059 14467
rect 15059 14433 15068 14467
rect 15016 14424 15068 14433
rect 17132 14492 17184 14544
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 16304 14467 16356 14476
rect 16304 14433 16313 14467
rect 16313 14433 16347 14467
rect 16347 14433 16356 14467
rect 16304 14424 16356 14433
rect 16580 14467 16632 14476
rect 16580 14433 16589 14467
rect 16589 14433 16623 14467
rect 16623 14433 16632 14467
rect 16580 14424 16632 14433
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 16948 14424 17000 14476
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 12808 14288 12860 14340
rect 13084 14331 13136 14340
rect 13084 14297 13093 14331
rect 13093 14297 13127 14331
rect 13127 14297 13136 14331
rect 13084 14288 13136 14297
rect 16212 14356 16264 14408
rect 17500 14356 17552 14408
rect 19524 14467 19576 14476
rect 19524 14433 19533 14467
rect 19533 14433 19567 14467
rect 19567 14433 19576 14467
rect 19524 14424 19576 14433
rect 19340 14399 19392 14408
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 19984 14467 20036 14476
rect 19984 14433 19993 14467
rect 19993 14433 20027 14467
rect 20027 14433 20036 14467
rect 19984 14424 20036 14433
rect 8668 14220 8720 14229
rect 15660 14220 15712 14272
rect 16580 14288 16632 14340
rect 16856 14288 16908 14340
rect 17500 14220 17552 14272
rect 19156 14288 19208 14340
rect 19892 14288 19944 14340
rect 20352 14356 20404 14408
rect 20536 14356 20588 14408
rect 23020 14424 23072 14476
rect 25964 14560 26016 14612
rect 26424 14560 26476 14612
rect 21180 14288 21232 14340
rect 22284 14288 22336 14340
rect 23204 14356 23256 14408
rect 23664 14424 23716 14476
rect 24032 14467 24084 14476
rect 24032 14433 24041 14467
rect 24041 14433 24075 14467
rect 24075 14433 24084 14467
rect 24032 14424 24084 14433
rect 24216 14492 24268 14544
rect 24308 14467 24360 14476
rect 24308 14433 24317 14467
rect 24317 14433 24351 14467
rect 24351 14433 24360 14467
rect 24308 14424 24360 14433
rect 24584 14424 24636 14476
rect 25320 14535 25372 14544
rect 25320 14501 25329 14535
rect 25329 14501 25363 14535
rect 25363 14501 25372 14535
rect 25320 14492 25372 14501
rect 25596 14356 25648 14408
rect 25964 14424 26016 14476
rect 26240 14424 26292 14476
rect 26976 14467 27028 14476
rect 26976 14433 26985 14467
rect 26985 14433 27019 14467
rect 27019 14433 27028 14467
rect 26976 14424 27028 14433
rect 29092 14560 29144 14612
rect 30656 14603 30708 14612
rect 30656 14569 30665 14603
rect 30665 14569 30699 14603
rect 30699 14569 30708 14603
rect 30656 14560 30708 14569
rect 27344 14467 27396 14476
rect 27344 14433 27353 14467
rect 27353 14433 27387 14467
rect 27387 14433 27396 14467
rect 27344 14424 27396 14433
rect 26056 14356 26108 14408
rect 24952 14331 25004 14340
rect 24952 14297 24961 14331
rect 24961 14297 24995 14331
rect 24995 14297 25004 14331
rect 24952 14288 25004 14297
rect 28172 14356 28224 14408
rect 28356 14467 28408 14476
rect 28356 14433 28365 14467
rect 28365 14433 28399 14467
rect 28399 14433 28408 14467
rect 28356 14424 28408 14433
rect 28632 14424 28684 14476
rect 28908 14467 28960 14476
rect 28908 14433 28917 14467
rect 28917 14433 28951 14467
rect 28951 14433 28960 14467
rect 28908 14424 28960 14433
rect 29736 14492 29788 14544
rect 29828 14467 29880 14476
rect 29828 14433 29837 14467
rect 29837 14433 29871 14467
rect 29871 14433 29880 14467
rect 29828 14424 29880 14433
rect 30012 14467 30064 14476
rect 30012 14433 30021 14467
rect 30021 14433 30055 14467
rect 30055 14433 30064 14467
rect 30012 14424 30064 14433
rect 30196 14467 30248 14476
rect 30196 14433 30205 14467
rect 30205 14433 30239 14467
rect 30239 14433 30248 14467
rect 30196 14424 30248 14433
rect 30472 14467 30524 14476
rect 30472 14433 30481 14467
rect 30481 14433 30515 14467
rect 30515 14433 30524 14467
rect 30472 14424 30524 14433
rect 31116 14492 31168 14544
rect 30932 14424 30984 14476
rect 27528 14288 27580 14340
rect 29736 14288 29788 14340
rect 31208 14356 31260 14408
rect 30840 14288 30892 14340
rect 20168 14220 20220 14272
rect 22468 14220 22520 14272
rect 22836 14263 22888 14272
rect 22836 14229 22845 14263
rect 22845 14229 22879 14263
rect 22879 14229 22888 14263
rect 22836 14220 22888 14229
rect 23480 14220 23532 14272
rect 24216 14220 24268 14272
rect 24584 14220 24636 14272
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 25688 14263 25740 14272
rect 25688 14229 25697 14263
rect 25697 14229 25731 14263
rect 25731 14229 25740 14263
rect 25688 14220 25740 14229
rect 27988 14220 28040 14272
rect 28080 14220 28132 14272
rect 28448 14220 28500 14272
rect 30288 14220 30340 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 11436 14118 11488 14170
rect 11500 14118 11552 14170
rect 11564 14118 11616 14170
rect 11628 14118 11680 14170
rect 11692 14118 11744 14170
rect 19210 14118 19262 14170
rect 19274 14118 19326 14170
rect 19338 14118 19390 14170
rect 19402 14118 19454 14170
rect 19466 14118 19518 14170
rect 26984 14118 27036 14170
rect 27048 14118 27100 14170
rect 27112 14118 27164 14170
rect 27176 14118 27228 14170
rect 27240 14118 27292 14170
rect 5356 14016 5408 14068
rect 5448 14016 5500 14068
rect 6000 14016 6052 14068
rect 6276 14016 6328 14068
rect 7012 14016 7064 14068
rect 2964 13880 3016 13932
rect 3332 13855 3384 13864
rect 3332 13821 3341 13855
rect 3341 13821 3375 13855
rect 3375 13821 3384 13855
rect 3332 13812 3384 13821
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 4712 13855 4764 13864
rect 4712 13821 4721 13855
rect 4721 13821 4755 13855
rect 4755 13821 4764 13855
rect 4712 13812 4764 13821
rect 4252 13744 4304 13796
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 5632 13880 5684 13932
rect 6000 13812 6052 13864
rect 6460 13855 6512 13864
rect 6460 13821 6469 13855
rect 6469 13821 6503 13855
rect 6503 13821 6512 13855
rect 6460 13812 6512 13821
rect 6920 13948 6972 14000
rect 5540 13744 5592 13796
rect 2596 13676 2648 13728
rect 3976 13676 4028 13728
rect 5448 13676 5500 13728
rect 5816 13676 5868 13728
rect 7104 13855 7156 13864
rect 7104 13821 7113 13855
rect 7113 13821 7147 13855
rect 7147 13821 7156 13855
rect 7104 13812 7156 13821
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 8392 14059 8444 14068
rect 8392 14025 8401 14059
rect 8401 14025 8435 14059
rect 8435 14025 8444 14059
rect 8392 14016 8444 14025
rect 9404 14059 9456 14068
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 10508 14016 10560 14068
rect 8668 13948 8720 14000
rect 8852 13948 8904 14000
rect 8944 13948 8996 14000
rect 9496 13948 9548 14000
rect 11612 14016 11664 14068
rect 11796 14016 11848 14068
rect 12532 14016 12584 14068
rect 13176 14016 13228 14068
rect 13820 14016 13872 14068
rect 14096 14016 14148 14068
rect 14924 14016 14976 14068
rect 16212 14016 16264 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 18420 14016 18472 14068
rect 18880 14016 18932 14068
rect 19340 14016 19392 14068
rect 19432 14016 19484 14068
rect 19800 14016 19852 14068
rect 19892 14016 19944 14068
rect 20444 14016 20496 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 8116 13855 8168 13864
rect 8116 13821 8125 13855
rect 8125 13821 8159 13855
rect 8159 13821 8168 13855
rect 8116 13812 8168 13821
rect 8300 13812 8352 13864
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 7840 13744 7892 13796
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 8852 13744 8904 13796
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 11060 13948 11112 14000
rect 12256 13948 12308 14000
rect 10600 13880 10652 13932
rect 15108 13948 15160 14000
rect 17224 13991 17276 14000
rect 17224 13957 17233 13991
rect 17233 13957 17267 13991
rect 17267 13957 17276 13991
rect 17224 13948 17276 13957
rect 17316 13948 17368 14000
rect 17684 13948 17736 14000
rect 18052 13948 18104 14000
rect 19064 13991 19116 14000
rect 19064 13957 19073 13991
rect 19073 13957 19107 13991
rect 19107 13957 19116 13991
rect 21548 14016 21600 14068
rect 21640 14016 21692 14068
rect 19064 13948 19116 13957
rect 13084 13880 13136 13932
rect 10324 13812 10376 13864
rect 10508 13744 10560 13796
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 14096 13880 14148 13932
rect 15936 13880 15988 13932
rect 16488 13880 16540 13932
rect 16672 13880 16724 13932
rect 6828 13676 6880 13728
rect 7472 13676 7524 13728
rect 11152 13676 11204 13728
rect 12624 13676 12676 13728
rect 13360 13676 13412 13728
rect 14096 13744 14148 13796
rect 14556 13812 14608 13864
rect 14740 13812 14792 13864
rect 15108 13855 15160 13864
rect 15108 13821 15117 13855
rect 15117 13821 15151 13855
rect 15151 13821 15160 13855
rect 15108 13812 15160 13821
rect 15384 13812 15436 13864
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 18236 13880 18288 13932
rect 18420 13880 18472 13932
rect 15200 13744 15252 13796
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 20904 13880 20956 13932
rect 19156 13855 19208 13864
rect 19156 13821 19165 13855
rect 19165 13821 19199 13855
rect 19199 13821 19208 13855
rect 19156 13812 19208 13821
rect 19248 13855 19300 13864
rect 19248 13821 19257 13855
rect 19257 13821 19291 13855
rect 19291 13821 19300 13855
rect 19248 13812 19300 13821
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 20536 13812 20588 13864
rect 21732 13923 21784 13932
rect 21732 13889 21741 13923
rect 21741 13889 21775 13923
rect 21775 13889 21784 13923
rect 21732 13880 21784 13889
rect 20168 13744 20220 13796
rect 20352 13744 20404 13796
rect 21180 13744 21232 13796
rect 21456 13855 21508 13864
rect 21456 13821 21465 13855
rect 21465 13821 21499 13855
rect 21499 13821 21508 13855
rect 21456 13812 21508 13821
rect 22284 14059 22336 14068
rect 22284 14025 22293 14059
rect 22293 14025 22327 14059
rect 22327 14025 22336 14059
rect 22284 14016 22336 14025
rect 22836 14016 22888 14068
rect 23940 14016 23992 14068
rect 25320 14016 25372 14068
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 26700 14016 26752 14068
rect 28632 14016 28684 14068
rect 28816 14016 28868 14068
rect 30748 14016 30800 14068
rect 24124 13948 24176 14000
rect 24584 13948 24636 14000
rect 25688 13948 25740 14000
rect 25964 13948 26016 14000
rect 26608 13948 26660 14000
rect 26884 13948 26936 14000
rect 28172 13948 28224 14000
rect 28448 13948 28500 14000
rect 22468 13812 22520 13864
rect 23572 13812 23624 13864
rect 24768 13880 24820 13932
rect 25412 13812 25464 13864
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 25964 13855 26016 13864
rect 25964 13821 25973 13855
rect 25973 13821 26007 13855
rect 26007 13821 26016 13855
rect 25964 13812 26016 13821
rect 28264 13855 28316 13864
rect 28264 13821 28273 13855
rect 28273 13821 28307 13855
rect 28307 13821 28316 13855
rect 28264 13812 28316 13821
rect 23388 13744 23440 13796
rect 23664 13744 23716 13796
rect 25136 13744 25188 13796
rect 29092 13812 29144 13864
rect 30656 13880 30708 13932
rect 30196 13812 30248 13864
rect 15660 13676 15712 13728
rect 19156 13676 19208 13728
rect 19616 13676 19668 13728
rect 22008 13676 22060 13728
rect 22468 13676 22520 13728
rect 22744 13719 22796 13728
rect 22744 13685 22753 13719
rect 22753 13685 22787 13719
rect 22787 13685 22796 13719
rect 22744 13676 22796 13685
rect 22836 13676 22888 13728
rect 25504 13676 25556 13728
rect 25596 13676 25648 13728
rect 27896 13676 27948 13728
rect 28448 13676 28500 13728
rect 29368 13744 29420 13796
rect 30104 13787 30156 13796
rect 30104 13753 30113 13787
rect 30113 13753 30147 13787
rect 30147 13753 30156 13787
rect 30104 13744 30156 13753
rect 31024 13812 31076 13864
rect 28908 13676 28960 13728
rect 29552 13676 29604 13728
rect 30288 13676 30340 13728
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 12096 13574 12148 13626
rect 12160 13574 12212 13626
rect 12224 13574 12276 13626
rect 12288 13574 12340 13626
rect 12352 13574 12404 13626
rect 19870 13574 19922 13626
rect 19934 13574 19986 13626
rect 19998 13574 20050 13626
rect 20062 13574 20114 13626
rect 20126 13574 20178 13626
rect 27644 13574 27696 13626
rect 27708 13574 27760 13626
rect 27772 13574 27824 13626
rect 27836 13574 27888 13626
rect 27900 13574 27952 13626
rect 3516 13472 3568 13524
rect 4528 13472 4580 13524
rect 5172 13472 5224 13524
rect 1032 13379 1084 13388
rect 1032 13345 1041 13379
rect 1041 13345 1075 13379
rect 1075 13345 1084 13379
rect 1032 13336 1084 13345
rect 1492 13404 1544 13456
rect 940 13268 992 13320
rect 1768 13336 1820 13388
rect 1952 13379 2004 13388
rect 1952 13345 1962 13379
rect 1962 13345 2004 13379
rect 1952 13336 2004 13345
rect 2596 13336 2648 13388
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3700 13404 3752 13456
rect 5540 13404 5592 13456
rect 5908 13404 5960 13456
rect 6000 13404 6052 13456
rect 3056 13379 3108 13388
rect 3056 13345 3065 13379
rect 3065 13345 3099 13379
rect 3099 13345 3108 13379
rect 3056 13336 3108 13345
rect 4620 13336 4672 13388
rect 4988 13336 5040 13388
rect 5172 13336 5224 13388
rect 7012 13404 7064 13456
rect 7196 13404 7248 13456
rect 7564 13472 7616 13524
rect 7656 13472 7708 13524
rect 8852 13515 8904 13524
rect 8852 13481 8861 13515
rect 8861 13481 8895 13515
rect 8895 13481 8904 13515
rect 8852 13472 8904 13481
rect 9128 13472 9180 13524
rect 6828 13336 6880 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 5908 13268 5960 13320
rect 7012 13268 7064 13320
rect 7288 13268 7340 13320
rect 7932 13336 7984 13388
rect 8484 13336 8536 13388
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 8944 13404 8996 13456
rect 9864 13404 9916 13456
rect 10508 13447 10560 13456
rect 10508 13413 10517 13447
rect 10517 13413 10551 13447
rect 10551 13413 10560 13447
rect 10508 13404 10560 13413
rect 10784 13404 10836 13456
rect 11244 13472 11296 13524
rect 11796 13472 11848 13524
rect 11980 13472 12032 13524
rect 12256 13472 12308 13524
rect 8852 13336 8904 13388
rect 10048 13336 10100 13388
rect 10324 13379 10376 13388
rect 10324 13345 10331 13379
rect 10331 13345 10376 13379
rect 3976 13200 4028 13252
rect 4344 13200 4396 13252
rect 4436 13200 4488 13252
rect 7380 13200 7432 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 3332 13132 3384 13184
rect 4160 13132 4212 13184
rect 5908 13132 5960 13184
rect 6276 13132 6328 13184
rect 6552 13132 6604 13184
rect 7104 13132 7156 13184
rect 7656 13200 7708 13252
rect 9956 13268 10008 13320
rect 10324 13336 10376 13345
rect 10416 13379 10468 13388
rect 10416 13345 10425 13379
rect 10425 13345 10459 13379
rect 10459 13345 10468 13379
rect 10416 13336 10468 13345
rect 10600 13379 10652 13388
rect 10600 13345 10614 13379
rect 10614 13345 10648 13379
rect 10648 13345 10652 13379
rect 10600 13336 10652 13345
rect 10508 13268 10560 13320
rect 7932 13132 7984 13184
rect 8024 13132 8076 13184
rect 8484 13200 8536 13252
rect 10968 13243 11020 13252
rect 10968 13209 10977 13243
rect 10977 13209 11011 13243
rect 11011 13209 11020 13243
rect 10968 13200 11020 13209
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 11704 13404 11756 13456
rect 12532 13472 12584 13524
rect 12900 13472 12952 13524
rect 13360 13472 13412 13524
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 11796 13336 11848 13388
rect 13452 13404 13504 13456
rect 14280 13404 14332 13456
rect 15476 13472 15528 13524
rect 18420 13472 18472 13524
rect 18972 13472 19024 13524
rect 12072 13268 12124 13320
rect 12992 13336 13044 13388
rect 14648 13336 14700 13388
rect 12256 13268 12308 13320
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 12716 13268 12768 13320
rect 13084 13268 13136 13320
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 13728 13268 13780 13320
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 15936 13404 15988 13456
rect 15292 13336 15344 13388
rect 15752 13336 15804 13388
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 16212 13336 16264 13388
rect 20076 13404 20128 13456
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 17224 13379 17276 13388
rect 17224 13345 17233 13379
rect 17233 13345 17267 13379
rect 17267 13345 17276 13379
rect 17224 13336 17276 13345
rect 17592 13336 17644 13388
rect 18144 13336 18196 13388
rect 15476 13268 15528 13320
rect 11796 13132 11848 13184
rect 12808 13200 12860 13252
rect 14280 13200 14332 13252
rect 15292 13200 15344 13252
rect 13820 13132 13872 13184
rect 14096 13132 14148 13184
rect 18420 13268 18472 13320
rect 18788 13379 18840 13388
rect 18788 13345 18797 13379
rect 18797 13345 18831 13379
rect 18831 13345 18840 13379
rect 18788 13336 18840 13345
rect 19064 13379 19116 13388
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 19156 13379 19208 13388
rect 19156 13345 19165 13379
rect 19165 13345 19199 13379
rect 19199 13345 19208 13379
rect 19156 13336 19208 13345
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 19892 13336 19944 13388
rect 20352 13336 20404 13388
rect 19340 13268 19392 13320
rect 20260 13268 20312 13320
rect 22100 13472 22152 13524
rect 22192 13472 22244 13524
rect 21180 13404 21232 13456
rect 22744 13515 22796 13524
rect 22744 13481 22753 13515
rect 22753 13481 22787 13515
rect 22787 13481 22796 13515
rect 22744 13472 22796 13481
rect 23112 13515 23164 13524
rect 23112 13481 23121 13515
rect 23121 13481 23155 13515
rect 23155 13481 23164 13515
rect 23112 13472 23164 13481
rect 25320 13472 25372 13524
rect 25504 13515 25556 13524
rect 25504 13481 25513 13515
rect 25513 13481 25547 13515
rect 25547 13481 25556 13515
rect 25504 13472 25556 13481
rect 25596 13472 25648 13524
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 21640 13379 21692 13388
rect 21640 13345 21649 13379
rect 21649 13345 21683 13379
rect 21683 13345 21692 13379
rect 21640 13336 21692 13345
rect 21180 13268 21232 13320
rect 21272 13268 21324 13320
rect 21916 13336 21968 13388
rect 22100 13336 22152 13388
rect 22376 13336 22428 13388
rect 25044 13404 25096 13456
rect 23664 13336 23716 13388
rect 24032 13379 24084 13388
rect 24032 13345 24041 13379
rect 24041 13345 24075 13379
rect 24075 13345 24084 13379
rect 24032 13336 24084 13345
rect 24492 13336 24544 13388
rect 24952 13336 25004 13388
rect 25412 13379 25464 13388
rect 25412 13345 25421 13379
rect 25421 13345 25455 13379
rect 25455 13345 25464 13379
rect 25412 13336 25464 13345
rect 28080 13472 28132 13524
rect 26148 13404 26200 13456
rect 26332 13404 26384 13456
rect 26516 13404 26568 13456
rect 25872 13336 25924 13388
rect 22836 13268 22888 13320
rect 24216 13268 24268 13320
rect 17040 13200 17092 13252
rect 17316 13243 17368 13252
rect 17316 13209 17325 13243
rect 17325 13209 17359 13243
rect 17359 13209 17368 13243
rect 17316 13200 17368 13209
rect 17408 13243 17460 13252
rect 17408 13209 17417 13243
rect 17417 13209 17451 13243
rect 17451 13209 17460 13243
rect 17408 13200 17460 13209
rect 17960 13200 18012 13252
rect 24032 13200 24084 13252
rect 25136 13311 25188 13320
rect 25136 13277 25145 13311
rect 25145 13277 25179 13311
rect 25179 13277 25188 13311
rect 25136 13268 25188 13277
rect 25780 13268 25832 13320
rect 26608 13379 26660 13388
rect 26608 13345 26617 13379
rect 26617 13345 26651 13379
rect 26651 13345 26660 13379
rect 26608 13336 26660 13345
rect 27804 13404 27856 13456
rect 27896 13404 27948 13456
rect 26976 13379 27028 13388
rect 26976 13345 26985 13379
rect 26985 13345 27019 13379
rect 27019 13345 27028 13379
rect 26976 13336 27028 13345
rect 27620 13336 27672 13388
rect 27712 13336 27764 13388
rect 28172 13336 28224 13388
rect 28448 13379 28500 13388
rect 28448 13345 28457 13379
rect 28457 13345 28491 13379
rect 28491 13345 28500 13379
rect 28448 13336 28500 13345
rect 29000 13447 29052 13456
rect 29000 13413 29027 13447
rect 29027 13413 29052 13447
rect 29000 13404 29052 13413
rect 29368 13404 29420 13456
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 16396 13132 16448 13184
rect 19524 13132 19576 13184
rect 19984 13132 20036 13184
rect 20076 13132 20128 13184
rect 20444 13132 20496 13184
rect 20628 13132 20680 13184
rect 22192 13175 22244 13184
rect 22192 13141 22201 13175
rect 22201 13141 22235 13175
rect 22235 13141 22244 13175
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 24676 13200 24728 13209
rect 26240 13200 26292 13252
rect 29644 13336 29696 13388
rect 30104 13404 30156 13456
rect 22192 13132 22244 13141
rect 24216 13175 24268 13184
rect 24216 13141 24225 13175
rect 24225 13141 24259 13175
rect 24259 13141 24268 13175
rect 24216 13132 24268 13141
rect 24308 13132 24360 13184
rect 26148 13175 26200 13184
rect 26148 13141 26157 13175
rect 26157 13141 26191 13175
rect 26191 13141 26200 13175
rect 26148 13132 26200 13141
rect 26332 13132 26384 13184
rect 27896 13200 27948 13252
rect 28724 13268 28776 13320
rect 28908 13268 28960 13320
rect 30840 13268 30892 13320
rect 29552 13200 29604 13252
rect 27436 13132 27488 13184
rect 27988 13132 28040 13184
rect 29092 13132 29144 13184
rect 29920 13175 29972 13184
rect 29920 13141 29929 13175
rect 29929 13141 29963 13175
rect 29963 13141 29972 13175
rect 29920 13132 29972 13141
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 11436 13030 11488 13082
rect 11500 13030 11552 13082
rect 11564 13030 11616 13082
rect 11628 13030 11680 13082
rect 11692 13030 11744 13082
rect 19210 13030 19262 13082
rect 19274 13030 19326 13082
rect 19338 13030 19390 13082
rect 19402 13030 19454 13082
rect 19466 13030 19518 13082
rect 26984 13030 27036 13082
rect 27048 13030 27100 13082
rect 27112 13030 27164 13082
rect 27176 13030 27228 13082
rect 27240 13030 27292 13082
rect 2504 12928 2556 12980
rect 2872 12928 2924 12980
rect 2780 12860 2832 12912
rect 3148 12860 3200 12912
rect 5172 12928 5224 12980
rect 6552 12928 6604 12980
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 6828 12928 6880 12980
rect 7196 12928 7248 12980
rect 7472 12928 7524 12980
rect 7748 12928 7800 12980
rect 8116 12928 8168 12980
rect 8944 12928 8996 12980
rect 11612 12928 11664 12980
rect 1952 12792 2004 12844
rect 4160 12792 4212 12844
rect 2136 12724 2188 12776
rect 2596 12724 2648 12776
rect 4528 12724 4580 12776
rect 4620 12724 4672 12776
rect 4804 12724 4856 12776
rect 5080 12724 5132 12776
rect 5264 12724 5316 12776
rect 5448 12724 5500 12776
rect 5908 12792 5960 12844
rect 3516 12588 3568 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 6000 12724 6052 12776
rect 6276 12835 6328 12844
rect 6276 12801 6285 12835
rect 6285 12801 6319 12835
rect 6319 12801 6328 12835
rect 6276 12792 6328 12801
rect 7012 12860 7064 12912
rect 8208 12860 8260 12912
rect 8484 12860 8536 12912
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 8760 12860 8812 12869
rect 10232 12860 10284 12912
rect 10968 12860 11020 12912
rect 12164 12928 12216 12980
rect 12348 12928 12400 12980
rect 13728 12971 13780 12980
rect 13728 12937 13737 12971
rect 13737 12937 13771 12971
rect 13771 12937 13780 12971
rect 13728 12928 13780 12937
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 16396 12928 16448 12980
rect 16764 12928 16816 12980
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 6828 12724 6880 12776
rect 6184 12656 6236 12708
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8024 12724 8076 12776
rect 8760 12724 8812 12776
rect 9128 12656 9180 12708
rect 9312 12792 9364 12844
rect 10508 12792 10560 12844
rect 12624 12860 12676 12912
rect 10416 12724 10468 12776
rect 10692 12656 10744 12708
rect 11336 12656 11388 12708
rect 12440 12724 12492 12776
rect 12716 12724 12768 12776
rect 9220 12588 9272 12640
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 12900 12656 12952 12708
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 15660 12860 15712 12912
rect 13728 12724 13780 12776
rect 14280 12724 14332 12776
rect 15844 12792 15896 12844
rect 15108 12724 15160 12776
rect 15292 12767 15344 12776
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 15476 12724 15528 12776
rect 13360 12656 13412 12708
rect 11796 12588 11848 12640
rect 15660 12724 15712 12776
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 17224 12860 17276 12912
rect 18788 12928 18840 12980
rect 20168 12928 20220 12980
rect 20812 12928 20864 12980
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 22652 12971 22704 12980
rect 22652 12937 22661 12971
rect 22661 12937 22695 12971
rect 22695 12937 22704 12971
rect 22652 12928 22704 12937
rect 23112 12928 23164 12980
rect 18236 12860 18288 12912
rect 17316 12724 17368 12776
rect 17040 12656 17092 12708
rect 15936 12588 15988 12640
rect 17224 12588 17276 12640
rect 17776 12724 17828 12776
rect 17960 12724 18012 12776
rect 19432 12792 19484 12844
rect 19156 12767 19208 12776
rect 19156 12733 19165 12767
rect 19165 12733 19199 12767
rect 19199 12733 19208 12767
rect 19156 12724 19208 12733
rect 19340 12656 19392 12708
rect 17776 12588 17828 12640
rect 18420 12588 18472 12640
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 20720 12792 20772 12844
rect 22100 12792 22152 12844
rect 22652 12792 22704 12844
rect 22836 12792 22888 12844
rect 23204 12792 23256 12844
rect 20260 12724 20312 12776
rect 21916 12724 21968 12776
rect 24032 12767 24084 12776
rect 24032 12733 24041 12767
rect 24041 12733 24075 12767
rect 24075 12733 24084 12767
rect 24032 12724 24084 12733
rect 24676 12792 24728 12844
rect 24584 12724 24636 12776
rect 26148 12792 26200 12844
rect 26516 12792 26568 12844
rect 26976 12792 27028 12844
rect 27160 12860 27212 12912
rect 27712 12860 27764 12912
rect 29000 12971 29052 12980
rect 29000 12937 29009 12971
rect 29009 12937 29043 12971
rect 29043 12937 29052 12971
rect 29000 12928 29052 12937
rect 29368 12971 29420 12980
rect 29368 12937 29377 12971
rect 29377 12937 29411 12971
rect 29411 12937 29420 12971
rect 29368 12928 29420 12937
rect 29920 12903 29972 12912
rect 29920 12869 29929 12903
rect 29929 12869 29963 12903
rect 29963 12869 29972 12903
rect 29920 12860 29972 12869
rect 19524 12656 19576 12708
rect 19984 12588 20036 12640
rect 20352 12588 20404 12640
rect 22008 12656 22060 12708
rect 20904 12588 20956 12640
rect 21824 12588 21876 12640
rect 24216 12699 24268 12708
rect 24216 12665 24225 12699
rect 24225 12665 24259 12699
rect 24259 12665 24268 12699
rect 24216 12656 24268 12665
rect 24308 12699 24360 12708
rect 24308 12665 24343 12699
rect 24343 12665 24360 12699
rect 24308 12656 24360 12665
rect 25136 12656 25188 12708
rect 26148 12656 26200 12708
rect 26700 12656 26752 12708
rect 27804 12724 27856 12776
rect 28632 12724 28684 12776
rect 28724 12724 28776 12776
rect 29184 12767 29236 12776
rect 29184 12733 29196 12767
rect 29196 12733 29230 12767
rect 29230 12733 29236 12767
rect 29184 12724 29236 12733
rect 30748 12724 30800 12776
rect 30840 12767 30892 12776
rect 30840 12733 30849 12767
rect 30849 12733 30883 12767
rect 30883 12733 30892 12767
rect 30840 12724 30892 12733
rect 29644 12699 29696 12708
rect 29644 12665 29653 12699
rect 29653 12665 29687 12699
rect 29687 12665 29696 12699
rect 29644 12656 29696 12665
rect 31576 12588 31628 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 12096 12486 12148 12538
rect 12160 12486 12212 12538
rect 12224 12486 12276 12538
rect 12288 12486 12340 12538
rect 12352 12486 12404 12538
rect 19870 12486 19922 12538
rect 19934 12486 19986 12538
rect 19998 12486 20050 12538
rect 20062 12486 20114 12538
rect 20126 12486 20178 12538
rect 27644 12486 27696 12538
rect 27708 12486 27760 12538
rect 27772 12486 27824 12538
rect 27836 12486 27888 12538
rect 27900 12486 27952 12538
rect 1860 12384 1912 12436
rect 3424 12384 3476 12436
rect 5172 12384 5224 12436
rect 5448 12384 5500 12436
rect 6184 12384 6236 12436
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 7564 12384 7616 12436
rect 7932 12384 7984 12436
rect 8576 12384 8628 12436
rect 9036 12384 9088 12436
rect 9772 12384 9824 12436
rect 1124 12316 1176 12368
rect 1952 12316 2004 12368
rect 1492 12248 1544 12300
rect 2044 12248 2096 12300
rect 3424 12291 3476 12300
rect 3424 12257 3433 12291
rect 3433 12257 3467 12291
rect 3467 12257 3476 12291
rect 3424 12248 3476 12257
rect 3516 12291 3568 12300
rect 3516 12257 3525 12291
rect 3525 12257 3559 12291
rect 3559 12257 3568 12291
rect 3516 12248 3568 12257
rect 3608 12248 3660 12300
rect 4712 12316 4764 12368
rect 5632 12316 5684 12368
rect 7104 12316 7156 12368
rect 8484 12316 8536 12368
rect 5264 12248 5316 12300
rect 7196 12291 7248 12300
rect 7196 12257 7205 12291
rect 7205 12257 7239 12291
rect 7239 12257 7248 12291
rect 7196 12248 7248 12257
rect 6000 12180 6052 12232
rect 7104 12223 7156 12232
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 7104 12180 7156 12189
rect 8392 12248 8444 12300
rect 8760 12248 8812 12300
rect 9220 12248 9272 12300
rect 10692 12316 10744 12368
rect 10968 12316 11020 12368
rect 12072 12316 12124 12368
rect 4160 12112 4212 12164
rect 4528 12112 4580 12164
rect 4804 12155 4856 12164
rect 4804 12121 4813 12155
rect 4813 12121 4847 12155
rect 4847 12121 4856 12155
rect 4804 12112 4856 12121
rect 5080 12112 5132 12164
rect 6552 12112 6604 12164
rect 2228 12044 2280 12096
rect 4436 12044 4488 12096
rect 4896 12044 4948 12096
rect 5172 12044 5224 12096
rect 6460 12044 6512 12096
rect 7748 12044 7800 12096
rect 7840 12044 7892 12096
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 10140 12248 10192 12300
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10876 12180 10928 12232
rect 8576 12112 8628 12164
rect 9220 12112 9272 12164
rect 9404 12155 9456 12164
rect 9404 12121 9413 12155
rect 9413 12121 9447 12155
rect 9447 12121 9456 12155
rect 9404 12112 9456 12121
rect 10140 12155 10192 12164
rect 10140 12121 10149 12155
rect 10149 12121 10183 12155
rect 10183 12121 10192 12155
rect 10140 12112 10192 12121
rect 10508 12112 10560 12164
rect 11520 12248 11572 12300
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 13360 12384 13412 12436
rect 15016 12427 15068 12436
rect 15016 12393 15025 12427
rect 15025 12393 15059 12427
rect 15059 12393 15068 12427
rect 15016 12384 15068 12393
rect 17408 12384 17460 12436
rect 18144 12384 18196 12436
rect 18604 12384 18656 12436
rect 18972 12384 19024 12436
rect 19248 12384 19300 12436
rect 20352 12384 20404 12436
rect 14096 12316 14148 12368
rect 12900 12248 12952 12300
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 11060 12180 11112 12232
rect 11888 12180 11940 12232
rect 12348 12180 12400 12232
rect 12992 12180 13044 12232
rect 9496 12044 9548 12096
rect 10232 12044 10284 12096
rect 10324 12044 10376 12096
rect 11152 12112 11204 12164
rect 10784 12044 10836 12096
rect 11336 12044 11388 12096
rect 11704 12112 11756 12164
rect 12900 12112 12952 12164
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 13728 12248 13780 12300
rect 14372 12291 14424 12300
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 20536 12316 20588 12368
rect 13544 12180 13596 12232
rect 13912 12223 13964 12232
rect 13912 12189 13921 12223
rect 13921 12189 13955 12223
rect 13955 12189 13964 12223
rect 13912 12180 13964 12189
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 14280 12180 14332 12232
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 15660 12223 15712 12232
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 15936 12180 15988 12232
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 17592 12248 17644 12300
rect 17776 12248 17828 12300
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 15476 12112 15528 12164
rect 12440 12044 12492 12096
rect 14188 12044 14240 12096
rect 15108 12087 15160 12096
rect 15108 12053 15117 12087
rect 15117 12053 15151 12087
rect 15151 12053 15160 12087
rect 15108 12044 15160 12053
rect 17408 12180 17460 12232
rect 18696 12248 18748 12300
rect 19064 12291 19116 12300
rect 19064 12257 19073 12291
rect 19073 12257 19107 12291
rect 19107 12257 19116 12291
rect 19064 12248 19116 12257
rect 19708 12248 19760 12300
rect 21548 12384 21600 12436
rect 21640 12384 21692 12436
rect 22928 12384 22980 12436
rect 23388 12384 23440 12436
rect 24032 12384 24084 12436
rect 25964 12384 26016 12436
rect 26516 12384 26568 12436
rect 22376 12316 22428 12368
rect 22560 12316 22612 12368
rect 21180 12248 21232 12300
rect 21916 12248 21968 12300
rect 22008 12248 22060 12300
rect 22744 12248 22796 12300
rect 22928 12291 22980 12300
rect 22928 12257 22937 12291
rect 22937 12257 22971 12291
rect 22971 12257 22980 12291
rect 22928 12248 22980 12257
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 23204 12291 23256 12300
rect 23204 12257 23213 12291
rect 23213 12257 23247 12291
rect 23247 12257 23256 12291
rect 23204 12248 23256 12257
rect 23296 12291 23348 12300
rect 23296 12257 23305 12291
rect 23305 12257 23339 12291
rect 23339 12257 23348 12291
rect 23296 12248 23348 12257
rect 24216 12316 24268 12368
rect 23572 12248 23624 12300
rect 18604 12180 18656 12232
rect 17500 12112 17552 12164
rect 18144 12112 18196 12164
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 20168 12180 20220 12232
rect 20352 12180 20404 12232
rect 22192 12180 22244 12232
rect 19248 12112 19300 12164
rect 19340 12112 19392 12164
rect 21456 12112 21508 12164
rect 25136 12291 25188 12300
rect 25136 12257 25145 12291
rect 25145 12257 25179 12291
rect 25179 12257 25188 12291
rect 25136 12248 25188 12257
rect 25504 12291 25556 12300
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 25780 12248 25832 12300
rect 26700 12359 26752 12368
rect 26700 12325 26709 12359
rect 26709 12325 26743 12359
rect 26743 12325 26752 12359
rect 26700 12316 26752 12325
rect 27160 12384 27212 12436
rect 27620 12316 27672 12368
rect 28356 12359 28408 12368
rect 28356 12325 28365 12359
rect 28365 12325 28399 12359
rect 28399 12325 28408 12359
rect 28356 12316 28408 12325
rect 29092 12359 29144 12368
rect 29092 12325 29101 12359
rect 29101 12325 29135 12359
rect 29135 12325 29144 12359
rect 29092 12316 29144 12325
rect 29920 12316 29972 12368
rect 26240 12291 26292 12300
rect 26240 12257 26249 12291
rect 26249 12257 26283 12291
rect 26283 12257 26292 12291
rect 26240 12248 26292 12257
rect 26424 12248 26476 12300
rect 26792 12291 26844 12300
rect 26792 12257 26801 12291
rect 26801 12257 26835 12291
rect 26835 12257 26844 12291
rect 26792 12248 26844 12257
rect 27068 12291 27120 12300
rect 27068 12257 27077 12291
rect 27077 12257 27111 12291
rect 27111 12257 27120 12291
rect 27068 12248 27120 12257
rect 27252 12248 27304 12300
rect 28080 12248 28132 12300
rect 17316 12044 17368 12096
rect 18512 12044 18564 12096
rect 22100 12044 22152 12096
rect 23112 12044 23164 12096
rect 23572 12044 23624 12096
rect 24860 12044 24912 12096
rect 25596 12044 25648 12096
rect 26516 12112 26568 12164
rect 27436 12112 27488 12164
rect 28724 12248 28776 12300
rect 28356 12180 28408 12232
rect 29368 12180 29420 12232
rect 28632 12112 28684 12164
rect 30288 12180 30340 12232
rect 26424 12044 26476 12096
rect 26700 12044 26752 12096
rect 26884 12044 26936 12096
rect 27804 12044 27856 12096
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 11436 11942 11488 11994
rect 11500 11942 11552 11994
rect 11564 11942 11616 11994
rect 11628 11942 11680 11994
rect 11692 11942 11744 11994
rect 19210 11942 19262 11994
rect 19274 11942 19326 11994
rect 19338 11942 19390 11994
rect 19402 11942 19454 11994
rect 19466 11942 19518 11994
rect 26984 11942 27036 11994
rect 27048 11942 27100 11994
rect 27112 11942 27164 11994
rect 27176 11942 27228 11994
rect 27240 11942 27292 11994
rect 1032 11840 1084 11892
rect 2504 11840 2556 11892
rect 2688 11840 2740 11892
rect 3148 11840 3200 11892
rect 3700 11840 3752 11892
rect 5172 11840 5224 11892
rect 6644 11840 6696 11892
rect 6736 11840 6788 11892
rect 7012 11840 7064 11892
rect 7656 11840 7708 11892
rect 3424 11772 3476 11824
rect 2228 11704 2280 11756
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 3608 11704 3660 11756
rect 3792 11704 3844 11756
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 1952 11679 2004 11688
rect 1952 11645 1961 11679
rect 1961 11645 1995 11679
rect 1995 11645 2004 11679
rect 1952 11636 2004 11645
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 2872 11679 2924 11688
rect 2872 11645 2883 11679
rect 2883 11645 2924 11679
rect 2872 11636 2924 11645
rect 3700 11636 3752 11688
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4068 11747 4120 11756
rect 5816 11772 5868 11824
rect 6000 11772 6052 11824
rect 7840 11815 7892 11824
rect 7840 11781 7849 11815
rect 7849 11781 7883 11815
rect 7883 11781 7892 11815
rect 7840 11772 7892 11781
rect 8300 11772 8352 11824
rect 8668 11772 8720 11824
rect 9128 11840 9180 11892
rect 9588 11840 9640 11892
rect 11796 11840 11848 11892
rect 9496 11772 9548 11824
rect 10048 11772 10100 11824
rect 10140 11772 10192 11824
rect 10324 11815 10376 11824
rect 10324 11781 10333 11815
rect 10333 11781 10367 11815
rect 10367 11781 10376 11815
rect 10324 11772 10376 11781
rect 10600 11772 10652 11824
rect 4068 11713 4096 11747
rect 4096 11713 4120 11747
rect 4068 11704 4120 11713
rect 1952 11500 2004 11552
rect 2136 11500 2188 11552
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 2596 11500 2648 11552
rect 3148 11568 3200 11620
rect 3424 11568 3476 11620
rect 4068 11568 4120 11620
rect 4528 11636 4580 11688
rect 4436 11568 4488 11620
rect 5172 11568 5224 11620
rect 5264 11568 5316 11620
rect 7196 11636 7248 11688
rect 7564 11636 7616 11688
rect 7840 11636 7892 11688
rect 8300 11568 8352 11620
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7104 11500 7156 11552
rect 7748 11500 7800 11552
rect 9128 11636 9180 11688
rect 10416 11636 10468 11688
rect 8852 11611 8904 11620
rect 8852 11577 8861 11611
rect 8861 11577 8895 11611
rect 8895 11577 8904 11611
rect 8852 11568 8904 11577
rect 10876 11636 10928 11688
rect 11060 11772 11112 11824
rect 14280 11840 14332 11892
rect 14372 11840 14424 11892
rect 15200 11840 15252 11892
rect 15476 11840 15528 11892
rect 15752 11840 15804 11892
rect 16304 11840 16356 11892
rect 17408 11840 17460 11892
rect 19432 11840 19484 11892
rect 11336 11704 11388 11756
rect 12532 11772 12584 11824
rect 11152 11679 11204 11688
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 11428 11679 11480 11688
rect 11428 11645 11437 11679
rect 11437 11645 11471 11679
rect 11471 11645 11480 11679
rect 11428 11636 11480 11645
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 11888 11704 11940 11756
rect 12624 11704 12676 11756
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 11980 11636 12032 11688
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 14832 11679 14884 11688
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 15108 11636 15160 11688
rect 15752 11636 15804 11688
rect 18236 11772 18288 11824
rect 18328 11704 18380 11756
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 19524 11704 19576 11756
rect 20076 11772 20128 11824
rect 20536 11840 20588 11892
rect 20996 11840 21048 11892
rect 21364 11840 21416 11892
rect 21732 11883 21784 11892
rect 21732 11849 21741 11883
rect 21741 11849 21775 11883
rect 21775 11849 21784 11883
rect 21732 11840 21784 11849
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 22284 11840 22336 11892
rect 24400 11840 24452 11892
rect 25872 11840 25924 11892
rect 26240 11883 26292 11892
rect 26240 11849 26249 11883
rect 26249 11849 26283 11883
rect 26283 11849 26292 11883
rect 26240 11840 26292 11849
rect 26424 11840 26476 11892
rect 28080 11883 28132 11892
rect 28080 11849 28089 11883
rect 28089 11849 28123 11883
rect 28123 11849 28132 11883
rect 28080 11840 28132 11849
rect 28264 11840 28316 11892
rect 28448 11840 28500 11892
rect 28724 11840 28776 11892
rect 24216 11772 24268 11824
rect 25504 11772 25556 11824
rect 26332 11772 26384 11824
rect 8944 11500 8996 11552
rect 9036 11500 9088 11552
rect 10416 11500 10468 11552
rect 10876 11500 10928 11552
rect 12348 11568 12400 11620
rect 13636 11568 13688 11620
rect 11336 11500 11388 11552
rect 11704 11500 11756 11552
rect 12992 11500 13044 11552
rect 13176 11500 13228 11552
rect 14648 11568 14700 11620
rect 14188 11500 14240 11552
rect 15568 11568 15620 11620
rect 16028 11568 16080 11620
rect 15200 11500 15252 11552
rect 18604 11636 18656 11688
rect 19432 11636 19484 11688
rect 21640 11704 21692 11756
rect 23296 11704 23348 11756
rect 24124 11704 24176 11756
rect 18880 11568 18932 11620
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 18144 11500 18196 11552
rect 19524 11500 19576 11552
rect 20076 11611 20128 11620
rect 20076 11577 20085 11611
rect 20085 11577 20119 11611
rect 20119 11577 20128 11611
rect 20076 11568 20128 11577
rect 21364 11636 21416 11688
rect 21824 11636 21876 11688
rect 22100 11636 22152 11688
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 22560 11679 22612 11688
rect 22560 11645 22569 11679
rect 22569 11645 22603 11679
rect 22603 11645 22612 11679
rect 22560 11636 22612 11645
rect 22744 11679 22796 11688
rect 22744 11645 22753 11679
rect 22753 11645 22787 11679
rect 22787 11645 22796 11679
rect 22744 11636 22796 11645
rect 23020 11636 23072 11688
rect 23940 11636 23992 11688
rect 24492 11636 24544 11688
rect 24952 11704 25004 11756
rect 25320 11679 25372 11688
rect 25320 11645 25329 11679
rect 25329 11645 25363 11679
rect 25363 11645 25372 11679
rect 25320 11636 25372 11645
rect 25504 11636 25556 11688
rect 25872 11636 25924 11688
rect 26148 11636 26200 11688
rect 26608 11747 26660 11756
rect 26608 11713 26617 11747
rect 26617 11713 26651 11747
rect 26651 11713 26660 11747
rect 26608 11704 26660 11713
rect 28356 11772 28408 11824
rect 27252 11704 27304 11756
rect 27712 11704 27764 11756
rect 28540 11704 28592 11756
rect 27068 11679 27120 11688
rect 27068 11645 27077 11679
rect 27077 11645 27111 11679
rect 27111 11645 27120 11679
rect 27068 11636 27120 11645
rect 27896 11636 27948 11688
rect 28356 11679 28408 11688
rect 28356 11645 28365 11679
rect 28365 11645 28399 11679
rect 28399 11645 28408 11679
rect 28356 11636 28408 11645
rect 29000 11636 29052 11688
rect 29460 11679 29512 11688
rect 29460 11645 29469 11679
rect 29469 11645 29503 11679
rect 29503 11645 29512 11679
rect 29460 11636 29512 11645
rect 29552 11679 29604 11688
rect 29552 11645 29561 11679
rect 29561 11645 29595 11679
rect 29595 11645 29604 11679
rect 29552 11636 29604 11645
rect 30472 11772 30524 11824
rect 29828 11704 29880 11756
rect 20628 11568 20680 11620
rect 24308 11568 24360 11620
rect 27528 11568 27580 11620
rect 28264 11568 28316 11620
rect 28540 11568 28592 11620
rect 28908 11568 28960 11620
rect 30012 11636 30064 11688
rect 31024 11704 31076 11756
rect 30288 11636 30340 11688
rect 21456 11500 21508 11552
rect 22652 11500 22704 11552
rect 24124 11500 24176 11552
rect 24492 11500 24544 11552
rect 25504 11543 25556 11552
rect 25504 11509 25506 11543
rect 25506 11509 25540 11543
rect 25540 11509 25556 11543
rect 25504 11500 25556 11509
rect 27436 11500 27488 11552
rect 27620 11500 27672 11552
rect 29092 11500 29144 11552
rect 29184 11500 29236 11552
rect 29644 11543 29696 11552
rect 29644 11509 29653 11543
rect 29653 11509 29687 11543
rect 29687 11509 29696 11543
rect 29644 11500 29696 11509
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 12096 11398 12148 11450
rect 12160 11398 12212 11450
rect 12224 11398 12276 11450
rect 12288 11398 12340 11450
rect 12352 11398 12404 11450
rect 19870 11398 19922 11450
rect 19934 11398 19986 11450
rect 19998 11398 20050 11450
rect 20062 11398 20114 11450
rect 20126 11398 20178 11450
rect 27644 11398 27696 11450
rect 27708 11398 27760 11450
rect 27772 11398 27824 11450
rect 27836 11398 27888 11450
rect 27900 11398 27952 11450
rect 1400 11296 1452 11348
rect 1308 11160 1360 11212
rect 2596 11296 2648 11348
rect 3976 11296 4028 11348
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 5172 11296 5224 11348
rect 6092 11296 6144 11348
rect 7656 11296 7708 11348
rect 1768 11228 1820 11280
rect 2136 11203 2188 11212
rect 2136 11169 2145 11203
rect 2145 11169 2179 11203
rect 2179 11169 2188 11203
rect 2136 11160 2188 11169
rect 2320 11228 2372 11280
rect 2964 11228 3016 11280
rect 3240 11228 3292 11280
rect 2412 11092 2464 11144
rect 3148 11203 3200 11212
rect 3148 11169 3157 11203
rect 3157 11169 3191 11203
rect 3191 11169 3200 11203
rect 3148 11160 3200 11169
rect 2964 11092 3016 11144
rect 3700 11160 3752 11212
rect 4528 11228 4580 11280
rect 4252 11160 4304 11212
rect 4712 11160 4764 11212
rect 3516 11092 3568 11144
rect 2872 11024 2924 11076
rect 5356 11160 5408 11212
rect 6736 11160 6788 11212
rect 6736 11024 6788 11076
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 8024 11160 8076 11212
rect 9588 11296 9640 11348
rect 10876 11296 10928 11348
rect 8300 11228 8352 11280
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9220 11160 9272 11212
rect 9036 11092 9088 11144
rect 9496 11160 9548 11212
rect 9772 11160 9824 11212
rect 10692 11092 10744 11144
rect 10876 11092 10928 11144
rect 11428 11203 11480 11212
rect 11428 11169 11437 11203
rect 11437 11169 11471 11203
rect 11471 11169 11480 11203
rect 11428 11160 11480 11169
rect 11704 11228 11756 11280
rect 13728 11296 13780 11348
rect 14464 11296 14516 11348
rect 14648 11296 14700 11348
rect 11980 11160 12032 11212
rect 12348 11092 12400 11144
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 12992 11160 13044 11212
rect 13268 11228 13320 11280
rect 13360 11203 13412 11212
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 13728 11160 13780 11212
rect 14188 11160 14240 11212
rect 14372 11160 14424 11212
rect 14924 11228 14976 11280
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 17500 11296 17552 11348
rect 19708 11296 19760 11348
rect 19892 11296 19944 11348
rect 20444 11296 20496 11348
rect 21180 11228 21232 11280
rect 21640 11228 21692 11280
rect 22560 11296 22612 11348
rect 23020 11296 23072 11348
rect 23480 11339 23532 11348
rect 23480 11305 23489 11339
rect 23489 11305 23523 11339
rect 23523 11305 23532 11339
rect 23480 11296 23532 11305
rect 15384 11160 15436 11212
rect 15568 11160 15620 11212
rect 16488 11203 16540 11212
rect 16488 11169 16497 11203
rect 16497 11169 16531 11203
rect 16531 11169 16540 11203
rect 16488 11160 16540 11169
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 17408 11160 17460 11212
rect 19156 11160 19208 11212
rect 19616 11160 19668 11212
rect 19708 11160 19760 11212
rect 19984 11160 20036 11212
rect 20444 11203 20496 11212
rect 20444 11169 20453 11203
rect 20453 11169 20487 11203
rect 20487 11169 20496 11203
rect 20444 11160 20496 11169
rect 22192 11160 22244 11212
rect 3700 10956 3752 11008
rect 3792 10956 3844 11008
rect 4436 10956 4488 11008
rect 4528 10956 4580 11008
rect 5816 10956 5868 11008
rect 6092 10956 6144 11008
rect 6552 10956 6604 11008
rect 6828 10956 6880 11008
rect 7748 10956 7800 11008
rect 8760 10956 8812 11008
rect 9036 10956 9088 11008
rect 9588 10999 9640 11008
rect 9588 10965 9597 10999
rect 9597 10965 9631 10999
rect 9631 10965 9640 10999
rect 9588 10956 9640 10965
rect 10232 10956 10284 11008
rect 10416 10956 10468 11008
rect 12624 11024 12676 11076
rect 13636 11092 13688 11144
rect 12900 10956 12952 11008
rect 14188 11024 14240 11076
rect 16028 11092 16080 11144
rect 16120 11092 16172 11144
rect 16764 11092 16816 11144
rect 13912 10956 13964 11008
rect 15384 11024 15436 11076
rect 15568 11024 15620 11076
rect 15660 11024 15712 11076
rect 19892 11024 19944 11076
rect 20076 11092 20128 11144
rect 21548 11092 21600 11144
rect 22836 11203 22888 11212
rect 22836 11169 22845 11203
rect 22845 11169 22879 11203
rect 22879 11169 22888 11203
rect 22836 11160 22888 11169
rect 24032 11296 24084 11348
rect 24308 11296 24360 11348
rect 24584 11296 24636 11348
rect 23848 11228 23900 11280
rect 24124 11228 24176 11280
rect 24768 11271 24820 11280
rect 24768 11237 24777 11271
rect 24777 11237 24811 11271
rect 24811 11237 24820 11271
rect 24768 11228 24820 11237
rect 25596 11296 25648 11348
rect 27436 11296 27488 11348
rect 25412 11271 25464 11280
rect 25412 11237 25421 11271
rect 25421 11237 25455 11271
rect 25455 11237 25464 11271
rect 25412 11228 25464 11237
rect 27988 11296 28040 11348
rect 28356 11296 28408 11348
rect 29552 11296 29604 11348
rect 24952 11160 25004 11212
rect 21916 11024 21968 11076
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 24400 11092 24452 11144
rect 25504 11203 25556 11212
rect 25504 11169 25513 11203
rect 25513 11169 25547 11203
rect 25547 11169 25556 11203
rect 25504 11160 25556 11169
rect 26240 11160 26292 11212
rect 27252 11203 27304 11212
rect 27252 11169 27261 11203
rect 27261 11169 27295 11203
rect 27295 11169 27304 11203
rect 27252 11160 27304 11169
rect 27804 11228 27856 11280
rect 27528 11160 27580 11212
rect 27712 11160 27764 11212
rect 28264 11203 28316 11212
rect 28264 11169 28273 11203
rect 28273 11169 28307 11203
rect 28307 11169 28316 11203
rect 28264 11160 28316 11169
rect 28724 11160 28776 11212
rect 29644 11228 29696 11280
rect 24032 11024 24084 11076
rect 18880 10956 18932 11008
rect 19984 10956 20036 11008
rect 20720 10956 20772 11008
rect 20904 10956 20956 11008
rect 22192 10956 22244 11008
rect 22836 10956 22888 11008
rect 26056 11024 26108 11076
rect 27712 11024 27764 11076
rect 29736 11203 29788 11212
rect 29736 11169 29745 11203
rect 29745 11169 29779 11203
rect 29779 11169 29788 11203
rect 29736 11160 29788 11169
rect 30932 11228 30984 11280
rect 29920 11203 29972 11212
rect 29920 11169 29929 11203
rect 29929 11169 29963 11203
rect 29963 11169 29972 11203
rect 29920 11160 29972 11169
rect 24308 10956 24360 11008
rect 25136 10956 25188 11008
rect 26884 10956 26936 11008
rect 27528 10956 27580 11008
rect 28816 10956 28868 11008
rect 29460 11092 29512 11144
rect 30564 11203 30616 11212
rect 30564 11169 30573 11203
rect 30573 11169 30607 11203
rect 30607 11169 30616 11203
rect 30564 11160 30616 11169
rect 29920 11024 29972 11076
rect 29736 10956 29788 11008
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 11436 10854 11488 10906
rect 11500 10854 11552 10906
rect 11564 10854 11616 10906
rect 11628 10854 11680 10906
rect 11692 10854 11744 10906
rect 19210 10854 19262 10906
rect 19274 10854 19326 10906
rect 19338 10854 19390 10906
rect 19402 10854 19454 10906
rect 19466 10854 19518 10906
rect 26984 10854 27036 10906
rect 27048 10854 27100 10906
rect 27112 10854 27164 10906
rect 27176 10854 27228 10906
rect 27240 10854 27292 10906
rect 2872 10752 2924 10804
rect 3056 10752 3108 10804
rect 3792 10752 3844 10804
rect 4068 10752 4120 10804
rect 4252 10752 4304 10804
rect 4804 10752 4856 10804
rect 1768 10684 1820 10736
rect 6000 10752 6052 10804
rect 6092 10795 6144 10804
rect 6092 10761 6101 10795
rect 6101 10761 6135 10795
rect 6135 10761 6144 10795
rect 6092 10752 6144 10761
rect 2596 10616 2648 10668
rect 5264 10684 5316 10736
rect 2780 10548 2832 10600
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 2780 10412 2832 10464
rect 3700 10591 3752 10600
rect 3700 10557 3714 10591
rect 3714 10557 3748 10591
rect 3748 10557 3752 10591
rect 3700 10548 3752 10557
rect 3424 10480 3476 10532
rect 3516 10523 3568 10532
rect 3516 10489 3525 10523
rect 3525 10489 3559 10523
rect 3559 10489 3568 10523
rect 3516 10480 3568 10489
rect 4344 10591 4396 10600
rect 4344 10557 4353 10591
rect 4353 10557 4387 10591
rect 4387 10557 4396 10591
rect 4344 10548 4396 10557
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 5172 10616 5224 10668
rect 5448 10616 5500 10668
rect 7196 10752 7248 10804
rect 8024 10795 8076 10804
rect 8024 10761 8033 10795
rect 8033 10761 8067 10795
rect 8067 10761 8076 10795
rect 8024 10752 8076 10761
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 8300 10752 8352 10804
rect 5632 10548 5684 10600
rect 5724 10591 5776 10600
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 6276 10548 6328 10600
rect 6736 10548 6788 10600
rect 7012 10548 7064 10600
rect 5908 10480 5960 10532
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 7564 10591 7616 10600
rect 7564 10557 7573 10591
rect 7573 10557 7607 10591
rect 7607 10557 7616 10591
rect 7564 10548 7616 10557
rect 7748 10480 7800 10532
rect 8208 10616 8260 10668
rect 9312 10684 9364 10736
rect 9588 10684 9640 10736
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9496 10616 9548 10668
rect 4896 10412 4948 10464
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6184 10412 6236 10464
rect 6552 10412 6604 10464
rect 6920 10412 6972 10464
rect 8760 10480 8812 10532
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9312 10548 9364 10600
rect 9772 10548 9824 10600
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 9680 10412 9732 10464
rect 9772 10412 9824 10464
rect 10416 10616 10468 10668
rect 10140 10591 10192 10600
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 10232 10548 10284 10600
rect 10692 10684 10744 10736
rect 10968 10684 11020 10736
rect 11336 10752 11388 10804
rect 11704 10684 11756 10736
rect 12624 10684 12676 10736
rect 13176 10684 13228 10736
rect 10692 10551 10701 10578
rect 10701 10551 10735 10578
rect 10735 10551 10744 10578
rect 10692 10526 10744 10551
rect 10232 10412 10284 10464
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12532 10616 12584 10668
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 15292 10684 15344 10736
rect 15384 10684 15436 10736
rect 15568 10684 15620 10736
rect 15936 10684 15988 10736
rect 16304 10684 16356 10736
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 17408 10752 17460 10804
rect 17776 10752 17828 10804
rect 20168 10684 20220 10736
rect 20720 10684 20772 10736
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 13452 10548 13504 10600
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 15200 10616 15252 10668
rect 16488 10616 16540 10668
rect 14740 10591 14792 10600
rect 14740 10557 14749 10591
rect 14749 10557 14783 10591
rect 14783 10557 14792 10591
rect 14740 10548 14792 10557
rect 11888 10480 11940 10532
rect 13360 10480 13412 10532
rect 15844 10591 15896 10600
rect 15844 10557 15853 10591
rect 15853 10557 15887 10591
rect 15887 10557 15896 10591
rect 15844 10548 15896 10557
rect 15292 10480 15344 10532
rect 16764 10548 16816 10600
rect 16856 10548 16908 10600
rect 19708 10616 19760 10668
rect 17592 10591 17644 10600
rect 17592 10557 17601 10591
rect 17601 10557 17635 10591
rect 17635 10557 17644 10591
rect 17592 10548 17644 10557
rect 17776 10591 17828 10600
rect 17776 10557 17785 10591
rect 17785 10557 17819 10591
rect 17819 10557 17828 10591
rect 17776 10548 17828 10557
rect 18144 10548 18196 10600
rect 16028 10480 16080 10532
rect 10876 10412 10928 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 11612 10455 11664 10464
rect 11612 10421 11621 10455
rect 11621 10421 11655 10455
rect 11655 10421 11664 10455
rect 11612 10412 11664 10421
rect 11704 10412 11756 10464
rect 12164 10412 12216 10464
rect 12624 10412 12676 10464
rect 12992 10412 13044 10464
rect 13176 10412 13228 10464
rect 16672 10412 16724 10464
rect 17868 10480 17920 10532
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 18880 10591 18932 10600
rect 18880 10557 18889 10591
rect 18889 10557 18923 10591
rect 18923 10557 18932 10591
rect 18880 10548 18932 10557
rect 19156 10591 19208 10600
rect 19156 10557 19161 10591
rect 19161 10557 19195 10591
rect 19195 10557 19208 10591
rect 19156 10548 19208 10557
rect 20352 10616 20404 10668
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 19616 10480 19668 10532
rect 18696 10412 18748 10421
rect 19340 10412 19392 10464
rect 19708 10412 19760 10464
rect 19892 10412 19944 10464
rect 20168 10523 20220 10532
rect 20168 10489 20190 10523
rect 20190 10489 20220 10523
rect 20168 10480 20220 10489
rect 20444 10514 20496 10566
rect 21272 10727 21324 10736
rect 21272 10693 21281 10727
rect 21281 10693 21315 10727
rect 21315 10693 21324 10727
rect 21272 10684 21324 10693
rect 22284 10752 22336 10804
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 23296 10752 23348 10804
rect 24032 10752 24084 10804
rect 25688 10752 25740 10804
rect 26424 10752 26476 10804
rect 28080 10752 28132 10804
rect 20996 10616 21048 10668
rect 21456 10591 21508 10600
rect 21456 10557 21465 10591
rect 21465 10557 21499 10591
rect 21499 10557 21508 10591
rect 21456 10548 21508 10557
rect 21916 10616 21968 10668
rect 26056 10684 26108 10736
rect 26700 10684 26752 10736
rect 26792 10684 26844 10736
rect 27712 10684 27764 10736
rect 30380 10727 30432 10736
rect 30380 10693 30389 10727
rect 30389 10693 30423 10727
rect 30423 10693 30432 10727
rect 30380 10684 30432 10693
rect 21640 10548 21692 10600
rect 21824 10591 21876 10600
rect 21824 10557 21833 10591
rect 21833 10557 21867 10591
rect 21867 10557 21876 10591
rect 21824 10548 21876 10557
rect 22192 10548 22244 10600
rect 22836 10548 22888 10600
rect 24124 10591 24176 10600
rect 24124 10557 24133 10591
rect 24133 10557 24167 10591
rect 24167 10557 24176 10591
rect 24124 10548 24176 10557
rect 24400 10548 24452 10600
rect 23296 10480 23348 10532
rect 24308 10523 24360 10532
rect 24308 10489 24317 10523
rect 24317 10489 24351 10523
rect 24351 10489 24360 10523
rect 24308 10480 24360 10489
rect 24584 10591 24636 10600
rect 24584 10557 24593 10591
rect 24593 10557 24627 10591
rect 24627 10557 24636 10591
rect 24584 10548 24636 10557
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 26148 10480 26200 10532
rect 26332 10591 26384 10600
rect 26332 10557 26341 10591
rect 26341 10557 26375 10591
rect 26375 10557 26384 10591
rect 26332 10548 26384 10557
rect 26424 10591 26476 10600
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 26884 10548 26936 10600
rect 29184 10616 29236 10668
rect 22560 10412 22612 10464
rect 22744 10455 22796 10464
rect 22744 10421 22753 10455
rect 22753 10421 22787 10455
rect 22787 10421 22796 10455
rect 22744 10412 22796 10421
rect 25504 10412 25556 10464
rect 25596 10412 25648 10464
rect 27068 10480 27120 10532
rect 27896 10548 27948 10600
rect 29000 10548 29052 10600
rect 29276 10548 29328 10600
rect 30196 10548 30248 10600
rect 30288 10548 30340 10600
rect 30656 10591 30708 10600
rect 30656 10557 30665 10591
rect 30665 10557 30699 10591
rect 30699 10557 30708 10591
rect 30656 10548 30708 10557
rect 31024 10591 31076 10600
rect 31024 10557 31033 10591
rect 31033 10557 31067 10591
rect 31067 10557 31076 10591
rect 31024 10548 31076 10557
rect 27528 10480 27580 10532
rect 28448 10480 28500 10532
rect 29184 10480 29236 10532
rect 31116 10480 31168 10532
rect 26976 10412 27028 10464
rect 27160 10412 27212 10464
rect 28080 10412 28132 10464
rect 28632 10412 28684 10464
rect 28816 10455 28868 10464
rect 28816 10421 28825 10455
rect 28825 10421 28859 10455
rect 28859 10421 28868 10455
rect 28816 10412 28868 10421
rect 30104 10412 30156 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 12096 10310 12148 10362
rect 12160 10310 12212 10362
rect 12224 10310 12276 10362
rect 12288 10310 12340 10362
rect 12352 10310 12404 10362
rect 19870 10310 19922 10362
rect 19934 10310 19986 10362
rect 19998 10310 20050 10362
rect 20062 10310 20114 10362
rect 20126 10310 20178 10362
rect 27644 10310 27696 10362
rect 27708 10310 27760 10362
rect 27772 10310 27824 10362
rect 27836 10310 27888 10362
rect 27900 10310 27952 10362
rect 1308 10208 1360 10260
rect 3792 10251 3844 10260
rect 3792 10217 3801 10251
rect 3801 10217 3835 10251
rect 3835 10217 3844 10251
rect 3792 10208 3844 10217
rect 5908 10208 5960 10260
rect 4804 10140 4856 10192
rect 7012 10208 7064 10260
rect 7104 10208 7156 10260
rect 9220 10208 9272 10260
rect 3240 10072 3292 10124
rect 3884 10115 3936 10124
rect 3884 10081 3893 10115
rect 3893 10081 3927 10115
rect 3927 10081 3936 10115
rect 3884 10072 3936 10081
rect 1860 10004 1912 10056
rect 2320 10004 2372 10056
rect 4344 10072 4396 10124
rect 4528 10072 4580 10124
rect 5264 10072 5316 10124
rect 6460 10140 6512 10192
rect 6920 10140 6972 10192
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 7196 10072 7248 10124
rect 7564 10140 7616 10192
rect 9680 10208 9732 10260
rect 3424 9936 3476 9988
rect 5632 10004 5684 10056
rect 7380 10004 7432 10056
rect 7472 10004 7524 10056
rect 8208 10004 8260 10056
rect 4896 9936 4948 9988
rect 9036 10072 9088 10124
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 9404 10140 9456 10192
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 10140 10208 10192 10260
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 10692 10208 10744 10260
rect 12440 10208 12492 10260
rect 14004 10208 14056 10260
rect 10600 10140 10652 10192
rect 12624 10140 12676 10192
rect 9864 10115 9916 10124
rect 9864 10081 9873 10115
rect 9873 10081 9907 10115
rect 9907 10081 9916 10115
rect 9864 10072 9916 10081
rect 3608 9868 3660 9920
rect 6828 9868 6880 9920
rect 7196 9868 7248 9920
rect 9220 9936 9272 9988
rect 9404 10004 9456 10056
rect 10232 10072 10284 10124
rect 10508 10072 10560 10124
rect 10692 10072 10744 10124
rect 13084 10140 13136 10192
rect 14832 10208 14884 10260
rect 14924 10208 14976 10260
rect 16672 10208 16724 10260
rect 14740 10140 14792 10192
rect 10324 10004 10376 10056
rect 10876 10004 10928 10056
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 13452 10072 13504 10124
rect 13820 10072 13872 10124
rect 15844 10140 15896 10192
rect 16028 10140 16080 10192
rect 11888 9936 11940 9988
rect 12348 9936 12400 9988
rect 13912 10004 13964 10056
rect 14556 10004 14608 10056
rect 15016 10004 15068 10056
rect 17592 10208 17644 10260
rect 17776 10140 17828 10192
rect 16580 10072 16632 10124
rect 20996 10208 21048 10260
rect 21088 10208 21140 10260
rect 21640 10251 21692 10260
rect 21640 10217 21649 10251
rect 21649 10217 21683 10251
rect 21683 10217 21692 10251
rect 21640 10208 21692 10217
rect 18328 10140 18380 10192
rect 20720 10140 20772 10192
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 15292 9936 15344 9988
rect 17040 9936 17092 9988
rect 18236 10072 18288 10124
rect 18512 10072 18564 10124
rect 20628 10072 20680 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 21640 10072 21692 10124
rect 22192 10140 22244 10192
rect 22560 10140 22612 10192
rect 23112 10140 23164 10192
rect 22100 10115 22152 10124
rect 22100 10081 22109 10115
rect 22109 10081 22143 10115
rect 22143 10081 22152 10115
rect 22100 10072 22152 10081
rect 23020 10115 23072 10124
rect 23020 10081 23029 10115
rect 23029 10081 23063 10115
rect 23063 10081 23072 10115
rect 23020 10072 23072 10081
rect 23296 10115 23348 10124
rect 23296 10081 23305 10115
rect 23305 10081 23339 10115
rect 23339 10081 23348 10115
rect 23296 10072 23348 10081
rect 18328 10004 18380 10056
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 20996 10004 21048 10056
rect 17776 9936 17828 9988
rect 19156 9936 19208 9988
rect 22560 10004 22612 10056
rect 8852 9868 8904 9920
rect 8944 9868 8996 9920
rect 9496 9868 9548 9920
rect 9864 9868 9916 9920
rect 11152 9868 11204 9920
rect 11520 9868 11572 9920
rect 13728 9868 13780 9920
rect 14740 9868 14792 9920
rect 15384 9868 15436 9920
rect 16672 9868 16724 9920
rect 17316 9868 17368 9920
rect 22836 9936 22888 9988
rect 23848 10251 23900 10260
rect 23848 10217 23857 10251
rect 23857 10217 23891 10251
rect 23891 10217 23900 10251
rect 23848 10208 23900 10217
rect 24032 10251 24084 10260
rect 24032 10217 24059 10251
rect 24059 10217 24084 10251
rect 24032 10208 24084 10217
rect 24216 10183 24268 10192
rect 24216 10149 24225 10183
rect 24225 10149 24259 10183
rect 24259 10149 24268 10183
rect 24216 10140 24268 10149
rect 24308 10140 24360 10192
rect 25044 10208 25096 10260
rect 23756 10072 23808 10124
rect 25596 10140 25648 10192
rect 25044 10072 25096 10124
rect 25964 10140 26016 10192
rect 26056 10115 26108 10124
rect 26056 10081 26065 10115
rect 26065 10081 26099 10115
rect 26099 10081 26108 10115
rect 26056 10072 26108 10081
rect 26424 10208 26476 10260
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 24768 10047 24820 10056
rect 24768 10013 24777 10047
rect 24777 10013 24811 10047
rect 24811 10013 24820 10047
rect 24768 10004 24820 10013
rect 25596 9936 25648 9988
rect 25964 10047 26016 10056
rect 25964 10013 25973 10047
rect 25973 10013 26007 10047
rect 26007 10013 26016 10047
rect 25964 10004 26016 10013
rect 26608 10047 26660 10056
rect 26608 10013 26617 10047
rect 26617 10013 26651 10047
rect 26651 10013 26660 10047
rect 26608 10004 26660 10013
rect 27252 10115 27304 10124
rect 27252 10081 27261 10115
rect 27261 10081 27295 10115
rect 27295 10081 27304 10115
rect 27252 10072 27304 10081
rect 27528 10115 27580 10124
rect 27528 10081 27537 10115
rect 27537 10081 27571 10115
rect 27571 10081 27580 10115
rect 27528 10072 27580 10081
rect 28172 10115 28224 10124
rect 28172 10081 28181 10115
rect 28181 10081 28215 10115
rect 28215 10081 28224 10115
rect 28172 10072 28224 10081
rect 29184 10140 29236 10192
rect 26516 9936 26568 9988
rect 27988 10047 28040 10056
rect 27988 10013 27997 10047
rect 27997 10013 28031 10047
rect 28031 10013 28040 10047
rect 27988 10004 28040 10013
rect 28264 10047 28316 10056
rect 28264 10013 28273 10047
rect 28273 10013 28307 10047
rect 28307 10013 28316 10047
rect 28264 10004 28316 10013
rect 28356 10047 28408 10056
rect 28356 10013 28365 10047
rect 28365 10013 28399 10047
rect 28399 10013 28408 10047
rect 28356 10004 28408 10013
rect 26976 9936 27028 9988
rect 27160 9936 27212 9988
rect 21640 9868 21692 9920
rect 23572 9868 23624 9920
rect 23940 9868 23992 9920
rect 24768 9868 24820 9920
rect 25320 9868 25372 9920
rect 25780 9868 25832 9920
rect 26332 9868 26384 9920
rect 28080 9868 28132 9920
rect 29460 10072 29512 10124
rect 29552 10115 29604 10124
rect 29552 10081 29561 10115
rect 29561 10081 29595 10115
rect 29595 10081 29604 10115
rect 29552 10072 29604 10081
rect 29276 10004 29328 10056
rect 29736 10115 29788 10124
rect 29736 10081 29745 10115
rect 29745 10081 29779 10115
rect 29779 10081 29788 10115
rect 29736 10072 29788 10081
rect 30196 10208 30248 10260
rect 29920 10140 29972 10192
rect 30288 10140 30340 10192
rect 30104 10115 30156 10124
rect 30104 10081 30113 10115
rect 30113 10081 30147 10115
rect 30147 10081 30156 10115
rect 30104 10072 30156 10081
rect 30196 10115 30248 10124
rect 30196 10081 30205 10115
rect 30205 10081 30239 10115
rect 30239 10081 30248 10115
rect 30196 10072 30248 10081
rect 30840 10115 30892 10124
rect 30840 10081 30849 10115
rect 30849 10081 30883 10115
rect 30883 10081 30892 10115
rect 30840 10072 30892 10081
rect 28816 9936 28868 9988
rect 30840 9936 30892 9988
rect 31668 9936 31720 9988
rect 29644 9868 29696 9920
rect 30196 9868 30248 9920
rect 31116 9868 31168 9920
rect 31300 9911 31352 9920
rect 31300 9877 31309 9911
rect 31309 9877 31343 9911
rect 31343 9877 31352 9911
rect 31300 9868 31352 9877
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 11436 9766 11488 9818
rect 11500 9766 11552 9818
rect 11564 9766 11616 9818
rect 11628 9766 11680 9818
rect 11692 9766 11744 9818
rect 19210 9766 19262 9818
rect 19274 9766 19326 9818
rect 19338 9766 19390 9818
rect 19402 9766 19454 9818
rect 19466 9766 19518 9818
rect 26984 9766 27036 9818
rect 27048 9766 27100 9818
rect 27112 9766 27164 9818
rect 27176 9766 27228 9818
rect 27240 9766 27292 9818
rect 1584 9664 1636 9716
rect 3240 9707 3292 9716
rect 3240 9673 3249 9707
rect 3249 9673 3283 9707
rect 3283 9673 3292 9707
rect 3240 9664 3292 9673
rect 1308 9639 1360 9648
rect 1308 9605 1317 9639
rect 1317 9605 1351 9639
rect 1351 9605 1360 9639
rect 1308 9596 1360 9605
rect 1216 9528 1268 9580
rect 4252 9664 4304 9716
rect 4896 9664 4948 9716
rect 5448 9707 5500 9716
rect 5448 9673 5457 9707
rect 5457 9673 5491 9707
rect 5491 9673 5500 9707
rect 5448 9664 5500 9673
rect 5724 9664 5776 9716
rect 4528 9596 4580 9648
rect 1032 9460 1084 9512
rect 2044 9460 2096 9512
rect 2688 9460 2740 9512
rect 3056 9460 3108 9512
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 3792 9503 3844 9512
rect 3792 9469 3801 9503
rect 3801 9469 3835 9503
rect 3835 9469 3844 9503
rect 3792 9460 3844 9469
rect 4804 9639 4856 9648
rect 4804 9605 4813 9639
rect 4813 9605 4847 9639
rect 4847 9605 4856 9639
rect 4804 9596 4856 9605
rect 6460 9664 6512 9716
rect 5448 9528 5500 9580
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 4804 9460 4856 9512
rect 2964 9392 3016 9444
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 6000 9503 6052 9512
rect 6000 9469 6009 9503
rect 6009 9469 6043 9503
rect 6043 9469 6052 9503
rect 6000 9460 6052 9469
rect 1492 9324 1544 9376
rect 1860 9324 1912 9376
rect 3700 9324 3752 9376
rect 4436 9324 4488 9376
rect 4712 9324 4764 9376
rect 5264 9392 5316 9444
rect 5448 9435 5500 9444
rect 5448 9401 5457 9435
rect 5457 9401 5491 9435
rect 5491 9401 5500 9435
rect 5448 9392 5500 9401
rect 5816 9392 5868 9444
rect 8116 9664 8168 9716
rect 9588 9664 9640 9716
rect 9772 9664 9824 9716
rect 6828 9528 6880 9580
rect 7748 9528 7800 9580
rect 8852 9639 8904 9648
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 9128 9596 9180 9648
rect 11336 9707 11388 9716
rect 11336 9673 11345 9707
rect 11345 9673 11379 9707
rect 11379 9673 11388 9707
rect 11336 9664 11388 9673
rect 11428 9664 11480 9716
rect 6920 9460 6972 9512
rect 7104 9460 7156 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7840 9460 7892 9512
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10508 9528 10560 9580
rect 6368 9392 6420 9444
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9036 9503 9088 9512
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 9312 9460 9364 9512
rect 9404 9460 9456 9512
rect 12072 9596 12124 9648
rect 12348 9707 12400 9716
rect 12348 9673 12357 9707
rect 12357 9673 12391 9707
rect 12391 9673 12400 9707
rect 12348 9664 12400 9673
rect 12440 9664 12492 9716
rect 13820 9664 13872 9716
rect 12992 9596 13044 9648
rect 13176 9596 13228 9648
rect 13912 9596 13964 9648
rect 14188 9596 14240 9648
rect 14372 9596 14424 9648
rect 14556 9596 14608 9648
rect 15016 9596 15068 9648
rect 15200 9596 15252 9648
rect 8116 9392 8168 9444
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 12624 9460 12676 9512
rect 6828 9324 6880 9376
rect 7196 9324 7248 9376
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 8392 9324 8444 9376
rect 8760 9324 8812 9376
rect 9312 9324 9364 9376
rect 10140 9324 10192 9376
rect 10508 9324 10560 9376
rect 10600 9324 10652 9376
rect 10692 9324 10744 9376
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 12072 9392 12124 9444
rect 15384 9528 15436 9580
rect 15844 9596 15896 9648
rect 16948 9596 17000 9648
rect 17776 9664 17828 9716
rect 18236 9664 18288 9716
rect 18604 9664 18656 9716
rect 18788 9664 18840 9716
rect 19156 9596 19208 9648
rect 19432 9664 19484 9716
rect 19984 9664 20036 9716
rect 20904 9664 20956 9716
rect 21824 9664 21876 9716
rect 22744 9664 22796 9716
rect 23756 9664 23808 9716
rect 25412 9664 25464 9716
rect 25504 9664 25556 9716
rect 16488 9571 16540 9580
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 16672 9528 16724 9580
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 13360 9392 13412 9444
rect 13728 9460 13780 9512
rect 15200 9460 15252 9512
rect 16396 9460 16448 9512
rect 14188 9392 14240 9444
rect 14556 9392 14608 9444
rect 14464 9324 14516 9376
rect 15292 9392 15344 9444
rect 17224 9460 17276 9512
rect 17776 9528 17828 9580
rect 17868 9503 17920 9512
rect 17868 9469 17877 9503
rect 17877 9469 17911 9503
rect 17911 9469 17920 9503
rect 17868 9460 17920 9469
rect 17776 9392 17828 9444
rect 18236 9460 18288 9512
rect 18328 9460 18380 9512
rect 18972 9528 19024 9580
rect 19156 9503 19208 9512
rect 19156 9469 19165 9503
rect 19165 9469 19199 9503
rect 19199 9469 19208 9503
rect 19156 9460 19208 9469
rect 19340 9571 19392 9580
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 19524 9460 19576 9512
rect 19708 9503 19760 9512
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 19708 9460 19760 9469
rect 18972 9435 19024 9444
rect 18972 9401 18981 9435
rect 18981 9401 19015 9435
rect 19015 9401 19024 9435
rect 18972 9392 19024 9401
rect 19064 9435 19116 9444
rect 19064 9401 19073 9435
rect 19073 9401 19107 9435
rect 19107 9401 19116 9435
rect 19064 9392 19116 9401
rect 19340 9392 19392 9444
rect 20076 9528 20128 9580
rect 20352 9460 20404 9512
rect 21456 9596 21508 9648
rect 23112 9596 23164 9648
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 20996 9528 21048 9580
rect 21640 9528 21692 9580
rect 25228 9639 25280 9648
rect 25228 9605 25237 9639
rect 25237 9605 25271 9639
rect 25271 9605 25280 9639
rect 25228 9596 25280 9605
rect 26516 9639 26568 9648
rect 26516 9605 26525 9639
rect 26525 9605 26559 9639
rect 26559 9605 26568 9639
rect 26516 9596 26568 9605
rect 26792 9707 26844 9716
rect 26792 9673 26801 9707
rect 26801 9673 26835 9707
rect 26835 9673 26844 9707
rect 26792 9664 26844 9673
rect 27160 9596 27212 9648
rect 27620 9664 27672 9716
rect 27712 9664 27764 9716
rect 29000 9664 29052 9716
rect 20904 9392 20956 9444
rect 15844 9324 15896 9376
rect 16764 9324 16816 9376
rect 16948 9324 17000 9376
rect 17408 9324 17460 9376
rect 18604 9324 18656 9376
rect 19248 9324 19300 9376
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 22192 9503 22244 9512
rect 22192 9469 22201 9503
rect 22201 9469 22235 9503
rect 22235 9469 22244 9503
rect 22192 9460 22244 9469
rect 21824 9324 21876 9376
rect 22928 9460 22980 9512
rect 23020 9503 23072 9512
rect 23020 9469 23029 9503
rect 23029 9469 23063 9503
rect 23063 9469 23072 9503
rect 23020 9460 23072 9469
rect 22836 9392 22888 9444
rect 23572 9460 23624 9512
rect 24216 9460 24268 9512
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 26148 9528 26200 9580
rect 26700 9571 26752 9580
rect 26700 9537 26709 9571
rect 26709 9537 26743 9571
rect 26743 9537 26752 9571
rect 26700 9528 26752 9537
rect 25228 9503 25280 9512
rect 25228 9469 25237 9503
rect 25237 9469 25271 9503
rect 25271 9469 25280 9503
rect 25228 9460 25280 9469
rect 23664 9392 23716 9444
rect 22928 9324 22980 9376
rect 23848 9324 23900 9376
rect 24860 9392 24912 9444
rect 26056 9460 26108 9512
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 26976 9528 27028 9580
rect 27160 9503 27212 9512
rect 27160 9469 27169 9503
rect 27169 9469 27203 9503
rect 27203 9469 27212 9503
rect 27160 9460 27212 9469
rect 27344 9503 27396 9512
rect 27344 9469 27353 9503
rect 27353 9469 27387 9503
rect 27387 9469 27396 9503
rect 27344 9460 27396 9469
rect 27528 9571 27580 9580
rect 27528 9537 27537 9571
rect 27537 9537 27571 9571
rect 27571 9537 27580 9571
rect 27528 9528 27580 9537
rect 27712 9528 27764 9580
rect 27988 9528 28040 9580
rect 29184 9528 29236 9580
rect 25688 9392 25740 9444
rect 25780 9392 25832 9444
rect 29276 9460 29328 9512
rect 29368 9460 29420 9512
rect 29644 9503 29696 9512
rect 29644 9469 29653 9503
rect 29653 9469 29687 9503
rect 29687 9469 29696 9503
rect 29644 9460 29696 9469
rect 29736 9503 29788 9512
rect 29736 9469 29745 9503
rect 29745 9469 29779 9503
rect 29779 9469 29788 9503
rect 29736 9460 29788 9469
rect 30196 9503 30248 9512
rect 30196 9469 30205 9503
rect 30205 9469 30239 9503
rect 30239 9469 30248 9503
rect 30196 9460 30248 9469
rect 31300 9528 31352 9580
rect 30380 9503 30432 9512
rect 30380 9469 30389 9503
rect 30389 9469 30423 9503
rect 30423 9469 30432 9503
rect 30380 9460 30432 9469
rect 30748 9460 30800 9512
rect 24952 9324 25004 9376
rect 25228 9324 25280 9376
rect 25504 9324 25556 9376
rect 26148 9324 26200 9376
rect 26332 9367 26384 9376
rect 26332 9333 26341 9367
rect 26341 9333 26375 9367
rect 26375 9333 26384 9367
rect 26332 9324 26384 9333
rect 28448 9324 28500 9376
rect 31024 9503 31076 9512
rect 31024 9469 31033 9503
rect 31033 9469 31067 9503
rect 31067 9469 31076 9503
rect 31024 9460 31076 9469
rect 31116 9503 31168 9512
rect 31116 9469 31125 9503
rect 31125 9469 31159 9503
rect 31159 9469 31168 9503
rect 31116 9460 31168 9469
rect 31760 9460 31812 9512
rect 31300 9392 31352 9444
rect 30840 9324 30892 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 12096 9222 12148 9274
rect 12160 9222 12212 9274
rect 12224 9222 12276 9274
rect 12288 9222 12340 9274
rect 12352 9222 12404 9274
rect 19870 9222 19922 9274
rect 19934 9222 19986 9274
rect 19998 9222 20050 9274
rect 20062 9222 20114 9274
rect 20126 9222 20178 9274
rect 27644 9222 27696 9274
rect 27708 9222 27760 9274
rect 27772 9222 27824 9274
rect 27836 9222 27888 9274
rect 27900 9222 27952 9274
rect 1032 9163 1084 9172
rect 1032 9129 1041 9163
rect 1041 9129 1075 9163
rect 1075 9129 1084 9163
rect 1032 9120 1084 9129
rect 1216 9027 1268 9036
rect 1216 8993 1225 9027
rect 1225 8993 1259 9027
rect 1259 8993 1268 9027
rect 1216 8984 1268 8993
rect 1768 9120 1820 9172
rect 2504 9120 2556 9172
rect 2596 9163 2648 9172
rect 2596 9129 2605 9163
rect 2605 9129 2639 9163
rect 2639 9129 2648 9163
rect 2596 9120 2648 9129
rect 3792 9120 3844 9172
rect 4068 9120 4120 9172
rect 4712 9120 4764 9172
rect 6000 9120 6052 9172
rect 6828 9120 6880 9172
rect 9404 9120 9456 9172
rect 2872 9052 2924 9104
rect 1584 8984 1636 9036
rect 2964 8984 3016 9036
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 3056 8984 3108 8993
rect 2044 8916 2096 8968
rect 4068 8984 4120 9036
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 4896 8984 4948 9036
rect 3700 8916 3752 8968
rect 4436 8916 4488 8968
rect 5080 8984 5132 9036
rect 1952 8780 2004 8832
rect 2872 8780 2924 8832
rect 4896 8780 4948 8832
rect 5080 8780 5132 8832
rect 5264 8984 5316 9036
rect 5632 9052 5684 9104
rect 6368 9052 6420 9104
rect 6736 9052 6788 9104
rect 8208 9052 8260 9104
rect 5816 8984 5868 9036
rect 6460 8984 6512 9036
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 8668 8984 8720 8993
rect 8944 8984 8996 9036
rect 9220 9027 9272 9036
rect 9220 8993 9229 9027
rect 9229 8993 9263 9027
rect 9263 8993 9272 9027
rect 9220 8984 9272 8993
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 10232 9120 10284 9172
rect 10416 9120 10468 9172
rect 11704 9120 11756 9172
rect 11888 9120 11940 9172
rect 13912 9120 13964 9172
rect 9588 9095 9640 9104
rect 9588 9061 9597 9095
rect 9597 9061 9631 9095
rect 9631 9061 9640 9095
rect 9588 9052 9640 9061
rect 10048 8984 10100 9036
rect 11520 9052 11572 9104
rect 11612 8984 11664 9036
rect 13176 9052 13228 9104
rect 16396 9120 16448 9172
rect 18972 9120 19024 9172
rect 19708 9120 19760 9172
rect 6368 8916 6420 8968
rect 7380 8916 7432 8968
rect 8484 8916 8536 8968
rect 11980 8916 12032 8968
rect 12900 8984 12952 9036
rect 12624 8916 12676 8968
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 13636 8916 13688 8968
rect 13912 8984 13964 9036
rect 14280 9027 14332 9036
rect 14280 8993 14289 9027
rect 14289 8993 14323 9027
rect 14323 8993 14332 9027
rect 14280 8984 14332 8993
rect 17040 9052 17092 9104
rect 20444 9163 20496 9172
rect 20444 9129 20453 9163
rect 20453 9129 20487 9163
rect 20487 9129 20496 9163
rect 20444 9120 20496 9129
rect 20536 9120 20588 9172
rect 20904 9120 20956 9172
rect 22836 9120 22888 9172
rect 23020 9163 23072 9172
rect 23020 9129 23029 9163
rect 23029 9129 23063 9163
rect 23063 9129 23072 9163
rect 23020 9120 23072 9129
rect 23480 9120 23532 9172
rect 15016 9027 15068 9036
rect 15016 8993 15025 9027
rect 15025 8993 15059 9027
rect 15059 8993 15068 9027
rect 15016 8984 15068 8993
rect 7012 8848 7064 8900
rect 9772 8848 9824 8900
rect 10140 8848 10192 8900
rect 12440 8848 12492 8900
rect 13728 8848 13780 8900
rect 15384 8916 15436 8968
rect 14924 8848 14976 8900
rect 6276 8780 6328 8832
rect 7380 8780 7432 8832
rect 8208 8780 8260 8832
rect 8392 8780 8444 8832
rect 8484 8780 8536 8832
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 9128 8780 9180 8832
rect 10324 8780 10376 8832
rect 12348 8780 12400 8832
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 13176 8780 13228 8832
rect 15936 8848 15988 8900
rect 15384 8780 15436 8832
rect 16764 8984 16816 9036
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 17775 9027 17827 9036
rect 17775 8993 17785 9027
rect 17785 8993 17819 9027
rect 17819 8993 17827 9027
rect 17775 8984 17827 8993
rect 16764 8848 16816 8900
rect 17040 8780 17092 8832
rect 17224 8780 17276 8832
rect 17316 8780 17368 8832
rect 18052 8916 18104 8968
rect 18788 8984 18840 9036
rect 19156 8984 19208 9036
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 17684 8780 17736 8832
rect 17868 8780 17920 8832
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 19524 8848 19576 8900
rect 19984 8848 20036 8900
rect 20168 9027 20220 9036
rect 20168 8993 20177 9027
rect 20177 8993 20211 9027
rect 20211 8993 20220 9027
rect 20168 8984 20220 8993
rect 20996 8984 21048 9036
rect 20536 8848 20588 8900
rect 21088 8848 21140 8900
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 21732 9052 21784 9104
rect 22100 9052 22152 9104
rect 21824 9027 21876 9036
rect 21824 8993 21833 9027
rect 21833 8993 21867 9027
rect 21867 8993 21876 9027
rect 21824 8984 21876 8993
rect 22008 8984 22060 9036
rect 23020 8984 23072 9036
rect 23296 9027 23348 9036
rect 23296 8993 23305 9027
rect 23305 8993 23339 9027
rect 23339 8993 23348 9027
rect 23296 8984 23348 8993
rect 23664 9052 23716 9104
rect 23848 9052 23900 9104
rect 23572 8984 23624 9036
rect 22928 8916 22980 8968
rect 23112 8916 23164 8968
rect 23664 8916 23716 8968
rect 24032 9027 24084 9036
rect 24032 8993 24041 9027
rect 24041 8993 24075 9027
rect 24075 8993 24084 9027
rect 24032 8984 24084 8993
rect 24216 9027 24268 9036
rect 24216 8993 24225 9027
rect 24225 8993 24259 9027
rect 24259 8993 24268 9027
rect 24216 8984 24268 8993
rect 24492 9027 24544 9036
rect 24492 8993 24501 9027
rect 24501 8993 24535 9027
rect 24535 8993 24544 9027
rect 24492 8984 24544 8993
rect 25964 9120 26016 9172
rect 26056 9120 26108 9172
rect 27528 9120 27580 9172
rect 28264 9120 28316 9172
rect 28356 9120 28408 9172
rect 29092 9120 29144 9172
rect 29368 9120 29420 9172
rect 29644 9120 29696 9172
rect 30288 9120 30340 9172
rect 24400 8891 24452 8900
rect 19340 8780 19392 8832
rect 19800 8823 19852 8832
rect 19800 8789 19809 8823
rect 19809 8789 19843 8823
rect 19843 8789 19852 8823
rect 19800 8780 19852 8789
rect 19892 8780 19944 8832
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 20260 8780 20312 8789
rect 20628 8780 20680 8832
rect 24400 8857 24409 8891
rect 24409 8857 24443 8891
rect 24443 8857 24452 8891
rect 24400 8848 24452 8857
rect 30840 9052 30892 9104
rect 31208 9052 31260 9104
rect 25412 9027 25464 9036
rect 25412 8993 25421 9027
rect 25421 8993 25455 9027
rect 25455 8993 25464 9027
rect 25412 8984 25464 8993
rect 26884 8984 26936 9036
rect 25228 8916 25280 8968
rect 26792 8916 26844 8968
rect 27344 8984 27396 9036
rect 26700 8848 26752 8900
rect 22008 8780 22060 8832
rect 23480 8780 23532 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 25964 8780 26016 8832
rect 26424 8780 26476 8832
rect 26516 8780 26568 8832
rect 27436 8848 27488 8900
rect 27620 8984 27672 9036
rect 28356 8984 28408 9036
rect 28908 9027 28960 9036
rect 27712 8916 27764 8968
rect 28908 8993 28917 9027
rect 28917 8993 28951 9027
rect 28951 8993 28960 9027
rect 28908 8984 28960 8993
rect 29460 8984 29512 9036
rect 29920 8984 29972 9036
rect 30104 9027 30156 9036
rect 30104 8993 30113 9027
rect 30113 8993 30147 9027
rect 30147 8993 30156 9027
rect 30104 8984 30156 8993
rect 30196 9027 30248 9036
rect 30196 8993 30205 9027
rect 30205 8993 30239 9027
rect 30239 8993 30248 9027
rect 30196 8984 30248 8993
rect 30564 8984 30616 9036
rect 30932 8984 30984 9036
rect 31484 8984 31536 9036
rect 27528 8780 27580 8832
rect 28080 8780 28132 8832
rect 29000 8848 29052 8900
rect 29368 8891 29420 8900
rect 29368 8857 29377 8891
rect 29377 8857 29411 8891
rect 29411 8857 29420 8891
rect 29368 8848 29420 8857
rect 30380 8916 30432 8968
rect 30196 8848 30248 8900
rect 30472 8848 30524 8900
rect 31300 8848 31352 8900
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 11436 8678 11488 8730
rect 11500 8678 11552 8730
rect 11564 8678 11616 8730
rect 11628 8678 11680 8730
rect 11692 8678 11744 8730
rect 19210 8678 19262 8730
rect 19274 8678 19326 8730
rect 19338 8678 19390 8730
rect 19402 8678 19454 8730
rect 19466 8678 19518 8730
rect 26984 8678 27036 8730
rect 27048 8678 27100 8730
rect 27112 8678 27164 8730
rect 27176 8678 27228 8730
rect 27240 8678 27292 8730
rect 3056 8576 3108 8628
rect 3976 8576 4028 8628
rect 4344 8576 4396 8628
rect 4804 8576 4856 8628
rect 5080 8576 5132 8628
rect 5264 8576 5316 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 7840 8576 7892 8628
rect 8300 8576 8352 8628
rect 9404 8576 9456 8628
rect 10692 8576 10744 8628
rect 11152 8576 11204 8628
rect 11520 8576 11572 8628
rect 11796 8576 11848 8628
rect 12256 8576 12308 8628
rect 12808 8576 12860 8628
rect 1676 8508 1728 8560
rect 1584 8372 1636 8424
rect 1492 8304 1544 8356
rect 2044 8415 2096 8424
rect 2044 8381 2053 8415
rect 2053 8381 2087 8415
rect 2087 8381 2096 8415
rect 2044 8372 2096 8381
rect 2412 8508 2464 8560
rect 5816 8508 5868 8560
rect 6736 8508 6788 8560
rect 4160 8440 4212 8492
rect 3332 8372 3384 8424
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 4252 8372 4304 8424
rect 4620 8372 4672 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 6092 8440 6144 8492
rect 5080 8415 5132 8424
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 6460 8415 6512 8424
rect 2228 8304 2280 8356
rect 2872 8304 2924 8356
rect 5172 8304 5224 8356
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 2412 8236 2464 8288
rect 2964 8236 3016 8288
rect 3240 8236 3292 8288
rect 3700 8236 3752 8288
rect 4436 8236 4488 8288
rect 6460 8381 6469 8415
rect 6469 8381 6503 8415
rect 6503 8381 6512 8415
rect 6460 8372 6512 8381
rect 6552 8372 6604 8424
rect 7380 8508 7432 8560
rect 5632 8304 5684 8356
rect 7656 8372 7708 8424
rect 7840 8372 7892 8424
rect 8208 8440 8260 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 10692 8440 10744 8492
rect 10968 8440 11020 8492
rect 13728 8508 13780 8560
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 14188 8576 14240 8628
rect 8300 8372 8352 8424
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 9956 8372 10008 8424
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11428 8415 11480 8424
rect 11428 8381 11437 8415
rect 11437 8381 11471 8415
rect 11471 8381 11480 8415
rect 11428 8372 11480 8381
rect 11796 8372 11848 8424
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 12348 8415 12400 8424
rect 12348 8381 12357 8415
rect 12357 8381 12391 8415
rect 12391 8381 12400 8415
rect 12348 8372 12400 8381
rect 7932 8279 7984 8288
rect 7932 8245 7941 8279
rect 7941 8245 7975 8279
rect 7975 8245 7984 8279
rect 7932 8236 7984 8245
rect 8668 8236 8720 8288
rect 8852 8236 8904 8288
rect 9864 8236 9916 8288
rect 10416 8279 10468 8288
rect 10416 8245 10425 8279
rect 10425 8245 10459 8279
rect 10459 8245 10468 8279
rect 10416 8236 10468 8245
rect 11980 8304 12032 8356
rect 12624 8372 12676 8424
rect 12808 8415 12860 8424
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 13176 8372 13228 8424
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 13912 8415 13964 8424
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 15016 8551 15068 8560
rect 15016 8517 15025 8551
rect 15025 8517 15059 8551
rect 15059 8517 15068 8551
rect 15016 8508 15068 8517
rect 15384 8576 15436 8628
rect 18236 8576 18288 8628
rect 18972 8576 19024 8628
rect 19432 8576 19484 8628
rect 20352 8576 20404 8628
rect 20812 8576 20864 8628
rect 21640 8576 21692 8628
rect 22376 8619 22428 8628
rect 22376 8585 22385 8619
rect 22385 8585 22419 8619
rect 22419 8585 22428 8619
rect 22376 8576 22428 8585
rect 23112 8619 23164 8628
rect 23112 8585 23121 8619
rect 23121 8585 23155 8619
rect 23155 8585 23164 8619
rect 23112 8576 23164 8585
rect 24584 8576 24636 8628
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 25780 8576 25832 8628
rect 19248 8508 19300 8560
rect 19984 8508 20036 8560
rect 14188 8440 14240 8492
rect 16764 8440 16816 8492
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 13360 8304 13412 8356
rect 13452 8304 13504 8356
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14648 8372 14700 8424
rect 14556 8304 14608 8356
rect 16304 8372 16356 8424
rect 17592 8440 17644 8492
rect 18696 8440 18748 8492
rect 21548 8551 21600 8560
rect 21548 8517 21557 8551
rect 21557 8517 21591 8551
rect 21591 8517 21600 8551
rect 21548 8508 21600 8517
rect 21732 8508 21784 8560
rect 22744 8508 22796 8560
rect 23020 8508 23072 8560
rect 15016 8304 15068 8356
rect 15660 8304 15712 8356
rect 16488 8304 16540 8356
rect 16764 8304 16816 8356
rect 11336 8236 11388 8288
rect 11520 8236 11572 8288
rect 13728 8236 13780 8288
rect 13820 8236 13872 8288
rect 14740 8236 14792 8288
rect 14924 8236 14976 8288
rect 16304 8236 16356 8288
rect 17040 8279 17092 8288
rect 17040 8245 17049 8279
rect 17049 8245 17083 8279
rect 17083 8245 17092 8279
rect 17040 8236 17092 8245
rect 17316 8304 17368 8356
rect 17868 8415 17920 8424
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 18052 8372 18104 8424
rect 18236 8372 18288 8424
rect 18696 8347 18748 8356
rect 18696 8313 18705 8347
rect 18705 8313 18739 8347
rect 18739 8313 18748 8347
rect 18696 8304 18748 8313
rect 18788 8304 18840 8356
rect 18972 8304 19024 8356
rect 20720 8372 20772 8424
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 20904 8415 20956 8418
rect 20904 8381 20913 8415
rect 20913 8381 20947 8415
rect 20947 8381 20956 8415
rect 20904 8366 20956 8381
rect 21272 8372 21324 8424
rect 21732 8372 21784 8424
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 17960 8236 18012 8288
rect 18512 8236 18564 8288
rect 19156 8236 19208 8288
rect 20076 8304 20128 8356
rect 20352 8304 20404 8356
rect 21640 8304 21692 8356
rect 20720 8236 20772 8288
rect 22008 8372 22060 8424
rect 22376 8372 22428 8424
rect 22652 8415 22704 8424
rect 22652 8381 22661 8415
rect 22661 8381 22695 8415
rect 22695 8381 22704 8415
rect 22652 8372 22704 8381
rect 22836 8415 22888 8424
rect 22836 8381 22845 8415
rect 22845 8381 22879 8415
rect 22879 8381 22888 8415
rect 22836 8372 22888 8381
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 26332 8576 26384 8628
rect 23480 8415 23532 8424
rect 22008 8236 22060 8288
rect 22284 8236 22336 8288
rect 23480 8381 23489 8415
rect 23489 8381 23523 8415
rect 23523 8381 23532 8415
rect 23480 8372 23532 8381
rect 23112 8304 23164 8356
rect 24400 8415 24452 8424
rect 24400 8381 24409 8415
rect 24409 8381 24443 8415
rect 24443 8381 24452 8415
rect 24400 8372 24452 8381
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 24584 8372 24636 8381
rect 24768 8372 24820 8424
rect 25136 8372 25188 8424
rect 25596 8440 25648 8492
rect 26240 8483 26292 8492
rect 26240 8449 26249 8483
rect 26249 8449 26283 8483
rect 26283 8449 26292 8483
rect 26240 8440 26292 8449
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 25780 8415 25832 8424
rect 25780 8381 25789 8415
rect 25789 8381 25823 8415
rect 25823 8381 25832 8415
rect 25780 8372 25832 8381
rect 25964 8372 26016 8424
rect 26148 8415 26200 8424
rect 26148 8381 26157 8415
rect 26157 8381 26191 8415
rect 26191 8381 26200 8415
rect 26148 8372 26200 8381
rect 26424 8551 26476 8560
rect 26424 8517 26433 8551
rect 26433 8517 26467 8551
rect 26467 8517 26476 8551
rect 26424 8508 26476 8517
rect 27344 8576 27396 8628
rect 27896 8576 27948 8628
rect 27528 8508 27580 8560
rect 30104 8576 30156 8628
rect 30564 8576 30616 8628
rect 27988 8440 28040 8492
rect 24768 8236 24820 8288
rect 25044 8236 25096 8288
rect 25504 8236 25556 8288
rect 27528 8372 27580 8424
rect 29368 8483 29420 8492
rect 29368 8449 29377 8483
rect 29377 8449 29411 8483
rect 29411 8449 29420 8483
rect 29368 8440 29420 8449
rect 29920 8440 29972 8492
rect 27068 8347 27120 8356
rect 27068 8313 27077 8347
rect 27077 8313 27111 8347
rect 27111 8313 27120 8347
rect 27068 8304 27120 8313
rect 27252 8347 27304 8356
rect 27252 8313 27253 8347
rect 27253 8313 27287 8347
rect 27287 8313 27304 8347
rect 27252 8304 27304 8313
rect 27436 8347 27488 8356
rect 27436 8313 27445 8347
rect 27445 8313 27479 8347
rect 27479 8313 27488 8347
rect 27436 8304 27488 8313
rect 28264 8304 28316 8356
rect 29276 8372 29328 8424
rect 30012 8372 30064 8424
rect 30104 8415 30156 8424
rect 30104 8381 30113 8415
rect 30113 8381 30147 8415
rect 30147 8381 30156 8415
rect 30104 8372 30156 8381
rect 30288 8415 30340 8424
rect 30288 8381 30297 8415
rect 30297 8381 30331 8415
rect 30331 8381 30340 8415
rect 30288 8372 30340 8381
rect 30840 8415 30892 8424
rect 30840 8381 30849 8415
rect 30849 8381 30883 8415
rect 30883 8381 30892 8415
rect 30840 8372 30892 8381
rect 26792 8236 26844 8288
rect 27804 8279 27856 8288
rect 27804 8245 27813 8279
rect 27813 8245 27847 8279
rect 27847 8245 27856 8279
rect 27804 8236 27856 8245
rect 28632 8236 28684 8288
rect 28908 8236 28960 8288
rect 29000 8279 29052 8288
rect 29000 8245 29009 8279
rect 29009 8245 29043 8279
rect 29043 8245 29052 8279
rect 29000 8236 29052 8245
rect 31668 8304 31720 8356
rect 29552 8236 29604 8288
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 12096 8134 12148 8186
rect 12160 8134 12212 8186
rect 12224 8134 12276 8186
rect 12288 8134 12340 8186
rect 12352 8134 12404 8186
rect 19870 8134 19922 8186
rect 19934 8134 19986 8186
rect 19998 8134 20050 8186
rect 20062 8134 20114 8186
rect 20126 8134 20178 8186
rect 27644 8134 27696 8186
rect 27708 8134 27760 8186
rect 27772 8134 27824 8186
rect 27836 8134 27888 8186
rect 27900 8134 27952 8186
rect 1860 8032 1912 8084
rect 9404 8032 9456 8084
rect 11428 8075 11480 8084
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 1308 7964 1360 8016
rect 1952 8007 2004 8016
rect 1952 7973 1961 8007
rect 1961 7973 1995 8007
rect 1995 7973 2004 8007
rect 1952 7964 2004 7973
rect 4344 7964 4396 8016
rect 5356 7964 5408 8016
rect 7380 7964 7432 8016
rect 8760 7964 8812 8016
rect 1492 7939 1544 7948
rect 1492 7905 1501 7939
rect 1501 7905 1535 7939
rect 1535 7905 1544 7939
rect 1492 7896 1544 7905
rect 1676 7896 1728 7948
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 4068 7896 4120 7948
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 5172 7896 5224 7948
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 9036 7964 9088 8016
rect 2228 7828 2280 7880
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 8760 7828 8812 7880
rect 8852 7871 8904 7880
rect 8852 7837 8861 7871
rect 8861 7837 8895 7871
rect 8895 7837 8904 7871
rect 8852 7828 8904 7837
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 10232 7964 10284 8016
rect 9956 7896 10008 7948
rect 10048 7896 10100 7948
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 11336 7896 11388 7948
rect 9312 7828 9364 7837
rect 9864 7828 9916 7880
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 4160 7760 4212 7812
rect 4896 7803 4948 7812
rect 4896 7769 4905 7803
rect 4905 7769 4939 7803
rect 4939 7769 4948 7803
rect 4896 7760 4948 7769
rect 2044 7692 2096 7744
rect 3976 7692 4028 7744
rect 4252 7692 4304 7744
rect 4620 7692 4672 7744
rect 6644 7692 6696 7744
rect 9128 7692 9180 7744
rect 9496 7803 9548 7812
rect 9496 7769 9505 7803
rect 9505 7769 9539 7803
rect 9539 7769 9548 7803
rect 9496 7760 9548 7769
rect 10416 7692 10468 7744
rect 12624 7964 12676 8016
rect 12808 8032 12860 8084
rect 13268 8032 13320 8084
rect 13636 8032 13688 8084
rect 14648 8032 14700 8084
rect 15108 8032 15160 8084
rect 15292 8032 15344 8084
rect 15384 8032 15436 8084
rect 15844 8032 15896 8084
rect 16488 8032 16540 8084
rect 17040 8032 17092 8084
rect 18696 8032 18748 8084
rect 18972 8032 19024 8084
rect 12440 7896 12492 7948
rect 12624 7828 12676 7880
rect 13268 7896 13320 7948
rect 13544 7828 13596 7880
rect 13176 7760 13228 7812
rect 14004 7896 14056 7948
rect 14096 7939 14148 7948
rect 14096 7905 14105 7939
rect 14105 7905 14139 7939
rect 14139 7905 14148 7939
rect 14096 7896 14148 7905
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 14372 7939 14424 7948
rect 14372 7905 14381 7939
rect 14381 7905 14415 7939
rect 14415 7905 14424 7939
rect 14372 7896 14424 7905
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 14924 7939 14976 7948
rect 14924 7905 14933 7939
rect 14933 7905 14967 7939
rect 14967 7905 14976 7939
rect 14924 7896 14976 7905
rect 15384 7973 15436 7982
rect 15384 7939 15393 7973
rect 15393 7939 15427 7973
rect 15427 7939 15436 7973
rect 15384 7930 15436 7939
rect 16396 7964 16448 8016
rect 16856 7964 16908 8016
rect 13912 7828 13964 7880
rect 14832 7828 14884 7880
rect 12164 7692 12216 7744
rect 12624 7735 12676 7744
rect 12624 7701 12633 7735
rect 12633 7701 12667 7735
rect 12667 7701 12676 7735
rect 12624 7692 12676 7701
rect 12716 7692 12768 7744
rect 14372 7760 14424 7812
rect 13452 7692 13504 7744
rect 14096 7692 14148 7744
rect 14832 7692 14884 7744
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 17040 7939 17092 7948
rect 17040 7905 17049 7939
rect 17049 7905 17083 7939
rect 17083 7905 17092 7939
rect 17040 7896 17092 7905
rect 17224 7964 17276 8016
rect 18604 7964 18656 8016
rect 18788 7939 18840 7948
rect 18788 7905 18797 7939
rect 18797 7905 18831 7939
rect 18831 7905 18840 7939
rect 18788 7896 18840 7905
rect 18236 7828 18288 7880
rect 18972 7939 19024 7948
rect 18972 7905 19007 7939
rect 19007 7905 19024 7939
rect 18972 7896 19024 7905
rect 19156 7939 19208 7948
rect 19156 7905 19165 7939
rect 19165 7905 19199 7939
rect 19199 7905 19208 7939
rect 19156 7896 19208 7905
rect 19248 7939 19300 7948
rect 19248 7905 19257 7939
rect 19257 7905 19291 7939
rect 19291 7905 19300 7939
rect 19248 7896 19300 7905
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 20444 7964 20496 8016
rect 20904 8032 20956 8084
rect 21640 8032 21692 8084
rect 22100 8032 22152 8084
rect 23204 8032 23256 8084
rect 23388 8032 23440 8084
rect 24032 8032 24084 8084
rect 24308 8032 24360 8084
rect 24584 8032 24636 8084
rect 24952 8032 25004 8084
rect 21272 7964 21324 8016
rect 22376 7964 22428 8016
rect 25044 7964 25096 8016
rect 19800 7896 19852 7948
rect 19892 7896 19944 7948
rect 20352 7939 20404 7948
rect 20352 7905 20361 7939
rect 20361 7905 20395 7939
rect 20395 7905 20404 7939
rect 20352 7896 20404 7905
rect 20628 7939 20680 7948
rect 20628 7905 20637 7939
rect 20637 7905 20671 7939
rect 20671 7905 20680 7939
rect 20628 7896 20680 7905
rect 20996 7896 21048 7948
rect 22008 7939 22060 7948
rect 22008 7905 22017 7939
rect 22017 7905 22051 7939
rect 22051 7905 22060 7939
rect 22008 7896 22060 7905
rect 22100 7939 22152 7948
rect 22100 7905 22109 7939
rect 22109 7905 22143 7939
rect 22143 7905 22152 7939
rect 22100 7896 22152 7905
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 23388 7896 23440 7948
rect 23480 7939 23532 7948
rect 23480 7905 23489 7939
rect 23489 7905 23523 7939
rect 23523 7905 23532 7939
rect 23480 7896 23532 7905
rect 23664 7939 23716 7948
rect 23664 7905 23673 7939
rect 23673 7905 23707 7939
rect 23707 7905 23716 7939
rect 23664 7896 23716 7905
rect 24032 7896 24084 7948
rect 19340 7828 19392 7880
rect 20444 7828 20496 7880
rect 20076 7760 20128 7812
rect 16304 7692 16356 7744
rect 16672 7692 16724 7744
rect 18696 7692 18748 7744
rect 19248 7692 19300 7744
rect 19340 7692 19392 7744
rect 20260 7692 20312 7744
rect 20536 7760 20588 7812
rect 21640 7760 21692 7812
rect 20720 7692 20772 7744
rect 21088 7692 21140 7744
rect 22836 7760 22888 7812
rect 23848 7760 23900 7812
rect 22652 7692 22704 7744
rect 23756 7692 23808 7744
rect 24492 7939 24544 7948
rect 24492 7905 24501 7939
rect 24501 7905 24535 7939
rect 24535 7905 24544 7939
rect 24492 7896 24544 7905
rect 24676 7896 24728 7948
rect 24860 7896 24912 7948
rect 25136 7939 25188 7948
rect 25136 7905 25145 7939
rect 25145 7905 25179 7939
rect 25179 7905 25188 7939
rect 25136 7896 25188 7905
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 25780 8032 25832 8084
rect 28724 8075 28776 8084
rect 28724 8041 28733 8075
rect 28733 8041 28767 8075
rect 28767 8041 28776 8075
rect 28724 8032 28776 8041
rect 29552 8032 29604 8084
rect 29644 8032 29696 8084
rect 29920 8032 29972 8084
rect 30012 8032 30064 8084
rect 31576 8032 31628 8084
rect 25504 7760 25556 7812
rect 25964 7964 26016 8016
rect 26332 7896 26384 7948
rect 26884 7896 26936 7948
rect 26976 7939 27028 7948
rect 26976 7905 26985 7939
rect 26985 7905 27019 7939
rect 27019 7905 27028 7939
rect 26976 7896 27028 7905
rect 29276 7964 29328 8016
rect 25964 7828 26016 7880
rect 27896 7939 27948 7948
rect 27896 7905 27905 7939
rect 27905 7905 27939 7939
rect 27939 7905 27948 7939
rect 27896 7896 27948 7905
rect 27988 7896 28040 7948
rect 28356 7896 28408 7948
rect 28632 7896 28684 7948
rect 25688 7760 25740 7812
rect 25780 7760 25832 7812
rect 28080 7828 28132 7880
rect 26056 7692 26108 7744
rect 26516 7735 26568 7744
rect 26516 7701 26525 7735
rect 26525 7701 26559 7735
rect 26559 7701 26568 7735
rect 26516 7692 26568 7701
rect 28172 7760 28224 7812
rect 28356 7803 28408 7812
rect 28356 7769 28365 7803
rect 28365 7769 28399 7803
rect 28399 7769 28408 7803
rect 28356 7760 28408 7769
rect 29000 7760 29052 7812
rect 29552 7939 29604 7948
rect 29552 7905 29561 7939
rect 29561 7905 29595 7939
rect 29595 7905 29604 7939
rect 29552 7896 29604 7905
rect 29920 7939 29972 7948
rect 29920 7905 29929 7939
rect 29929 7905 29963 7939
rect 29963 7905 29972 7939
rect 29920 7896 29972 7905
rect 30472 7939 30524 7948
rect 30472 7905 30481 7939
rect 30481 7905 30515 7939
rect 30515 7905 30524 7939
rect 30472 7896 30524 7905
rect 31760 7896 31812 7948
rect 29184 7828 29236 7880
rect 30012 7760 30064 7812
rect 30288 7803 30340 7812
rect 30288 7769 30297 7803
rect 30297 7769 30331 7803
rect 30331 7769 30340 7803
rect 30288 7760 30340 7769
rect 29644 7692 29696 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 11436 7590 11488 7642
rect 11500 7590 11552 7642
rect 11564 7590 11616 7642
rect 11628 7590 11680 7642
rect 11692 7590 11744 7642
rect 19210 7590 19262 7642
rect 19274 7590 19326 7642
rect 19338 7590 19390 7642
rect 19402 7590 19454 7642
rect 19466 7590 19518 7642
rect 26984 7590 27036 7642
rect 27048 7590 27100 7642
rect 27112 7590 27164 7642
rect 27176 7590 27228 7642
rect 27240 7590 27292 7642
rect 1584 7488 1636 7540
rect 1952 7488 2004 7540
rect 3700 7488 3752 7540
rect 4252 7488 4304 7540
rect 4804 7488 4856 7540
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 4988 7488 5040 7540
rect 7288 7488 7340 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 9404 7488 9456 7540
rect 9588 7488 9640 7540
rect 10968 7488 11020 7540
rect 11060 7488 11112 7540
rect 11520 7488 11572 7540
rect 11796 7488 11848 7540
rect 14556 7488 14608 7540
rect 14832 7488 14884 7540
rect 15292 7488 15344 7540
rect 15476 7488 15528 7540
rect 16856 7488 16908 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 17500 7488 17552 7540
rect 18144 7488 18196 7540
rect 20444 7488 20496 7540
rect 20812 7488 20864 7540
rect 21824 7488 21876 7540
rect 1676 7420 1728 7472
rect 2228 7420 2280 7472
rect 1584 7284 1636 7336
rect 1400 7216 1452 7268
rect 1860 7284 1912 7336
rect 1952 7327 2004 7336
rect 1952 7293 1961 7327
rect 1961 7293 1995 7327
rect 1995 7293 2004 7327
rect 1952 7284 2004 7293
rect 4252 7352 4304 7404
rect 9956 7420 10008 7472
rect 2136 7284 2188 7336
rect 3516 7284 3568 7336
rect 3976 7327 4028 7336
rect 3976 7293 3985 7327
rect 3985 7293 4019 7327
rect 4019 7293 4028 7327
rect 3976 7284 4028 7293
rect 3608 7216 3660 7268
rect 3976 7148 4028 7200
rect 4344 7327 4396 7336
rect 4344 7293 4353 7327
rect 4353 7293 4387 7327
rect 4387 7293 4396 7327
rect 4344 7284 4396 7293
rect 4712 7284 4764 7336
rect 4804 7284 4856 7336
rect 4896 7284 4948 7336
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 7196 7352 7248 7404
rect 8208 7352 8260 7404
rect 6736 7284 6788 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 7012 7284 7064 7336
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 12164 7420 12216 7472
rect 8300 7216 8352 7268
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 14740 7352 14792 7404
rect 15844 7352 15896 7404
rect 5540 7148 5592 7200
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 7840 7148 7892 7200
rect 10508 7284 10560 7336
rect 11152 7284 11204 7336
rect 11980 7284 12032 7336
rect 12072 7284 12124 7336
rect 10140 7216 10192 7268
rect 12716 7216 12768 7268
rect 12992 7284 13044 7336
rect 13268 7284 13320 7336
rect 14556 7284 14608 7336
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 14924 7327 14976 7336
rect 14924 7293 14933 7327
rect 14933 7293 14967 7327
rect 14967 7293 14976 7327
rect 14924 7284 14976 7293
rect 15292 7284 15344 7336
rect 15384 7293 15393 7302
rect 15393 7293 15427 7302
rect 15427 7293 15436 7302
rect 15384 7250 15436 7293
rect 15476 7327 15528 7336
rect 15476 7293 15485 7327
rect 15485 7293 15519 7327
rect 15519 7293 15528 7327
rect 15476 7284 15528 7293
rect 9772 7148 9824 7200
rect 10232 7148 10284 7200
rect 11152 7148 11204 7200
rect 12532 7148 12584 7200
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 13176 7148 13228 7200
rect 15660 7327 15712 7336
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 15660 7284 15712 7293
rect 16304 7327 16356 7336
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 16396 7327 16448 7336
rect 16396 7293 16405 7327
rect 16405 7293 16439 7327
rect 16439 7293 16448 7327
rect 16396 7284 16448 7293
rect 16856 7352 16908 7404
rect 17408 7352 17460 7404
rect 18052 7352 18104 7404
rect 18788 7352 18840 7404
rect 19524 7352 19576 7404
rect 20260 7420 20312 7472
rect 20628 7420 20680 7472
rect 21180 7420 21232 7472
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 16764 7284 16816 7336
rect 19800 7284 19852 7336
rect 20076 7284 20128 7336
rect 20260 7327 20312 7336
rect 20260 7293 20269 7327
rect 20269 7293 20303 7327
rect 20303 7293 20312 7327
rect 20260 7284 20312 7293
rect 20904 7352 20956 7404
rect 17684 7216 17736 7268
rect 17960 7216 18012 7268
rect 16580 7148 16632 7200
rect 17224 7148 17276 7200
rect 17316 7148 17368 7200
rect 20812 7284 20864 7336
rect 20996 7327 21048 7336
rect 20996 7293 21005 7327
rect 21005 7293 21039 7327
rect 21039 7293 21048 7327
rect 20996 7284 21048 7293
rect 21180 7327 21232 7336
rect 21180 7293 21189 7327
rect 21189 7293 21223 7327
rect 21223 7293 21232 7327
rect 21180 7284 21232 7293
rect 23204 7488 23256 7540
rect 23848 7531 23900 7540
rect 23848 7497 23857 7531
rect 23857 7497 23891 7531
rect 23891 7497 23900 7531
rect 23848 7488 23900 7497
rect 24768 7488 24820 7540
rect 24952 7488 25004 7540
rect 26148 7531 26200 7540
rect 26148 7497 26157 7531
rect 26157 7497 26191 7531
rect 26191 7497 26200 7531
rect 26148 7488 26200 7497
rect 28356 7488 28408 7540
rect 28540 7488 28592 7540
rect 30104 7488 30156 7540
rect 30840 7488 30892 7540
rect 21732 7327 21784 7336
rect 21732 7293 21741 7327
rect 21741 7293 21775 7327
rect 21775 7293 21784 7327
rect 21732 7284 21784 7293
rect 21824 7284 21876 7336
rect 22284 7284 22336 7336
rect 24124 7420 24176 7472
rect 24400 7420 24452 7472
rect 24584 7420 24636 7472
rect 25044 7420 25096 7472
rect 23204 7352 23256 7404
rect 25412 7395 25464 7404
rect 25412 7361 25421 7395
rect 25421 7361 25455 7395
rect 25455 7361 25464 7395
rect 25412 7352 25464 7361
rect 22468 7216 22520 7268
rect 20628 7148 20680 7200
rect 22836 7327 22888 7336
rect 22836 7293 22845 7327
rect 22845 7293 22879 7327
rect 22879 7293 22888 7327
rect 22836 7284 22888 7293
rect 24032 7284 24084 7336
rect 24400 7284 24452 7336
rect 22744 7216 22796 7268
rect 24584 7327 24636 7336
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 25044 7284 25096 7336
rect 25504 7327 25556 7336
rect 25504 7293 25513 7327
rect 25513 7293 25547 7327
rect 25547 7293 25556 7327
rect 25504 7284 25556 7293
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 26516 7352 26568 7404
rect 26240 7284 26292 7336
rect 27068 7327 27120 7336
rect 27068 7293 27077 7327
rect 27077 7293 27111 7327
rect 27111 7293 27120 7327
rect 27068 7284 27120 7293
rect 27344 7284 27396 7336
rect 27436 7327 27488 7336
rect 27436 7293 27445 7327
rect 27445 7293 27479 7327
rect 27479 7293 27488 7327
rect 27436 7284 27488 7293
rect 28816 7352 28868 7404
rect 24860 7259 24912 7268
rect 24860 7225 24869 7259
rect 24869 7225 24903 7259
rect 24903 7225 24912 7259
rect 24860 7216 24912 7225
rect 25228 7259 25237 7268
rect 25237 7259 25271 7268
rect 25271 7259 25280 7268
rect 25228 7216 25280 7259
rect 24768 7148 24820 7200
rect 24952 7148 25004 7200
rect 26056 7148 26108 7200
rect 26792 7216 26844 7268
rect 27988 7216 28040 7268
rect 28172 7216 28224 7268
rect 28724 7284 28776 7336
rect 29184 7284 29236 7336
rect 29460 7327 29512 7336
rect 29460 7293 29469 7327
rect 29469 7293 29503 7327
rect 29503 7293 29512 7327
rect 29460 7284 29512 7293
rect 30656 7420 30708 7472
rect 30288 7352 30340 7404
rect 30380 7327 30432 7336
rect 30380 7293 30389 7327
rect 30389 7293 30423 7327
rect 30423 7293 30432 7327
rect 30380 7284 30432 7293
rect 29092 7216 29144 7268
rect 30104 7216 30156 7268
rect 28632 7148 28684 7200
rect 29000 7148 29052 7200
rect 29184 7148 29236 7200
rect 30196 7191 30248 7200
rect 30196 7157 30205 7191
rect 30205 7157 30239 7191
rect 30239 7157 30248 7191
rect 30196 7148 30248 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 12096 7046 12148 7098
rect 12160 7046 12212 7098
rect 12224 7046 12276 7098
rect 12288 7046 12340 7098
rect 12352 7046 12404 7098
rect 19870 7046 19922 7098
rect 19934 7046 19986 7098
rect 19998 7046 20050 7098
rect 20062 7046 20114 7098
rect 20126 7046 20178 7098
rect 27644 7046 27696 7098
rect 27708 7046 27760 7098
rect 27772 7046 27824 7098
rect 27836 7046 27888 7098
rect 27900 7046 27952 7098
rect 1584 6944 1636 6996
rect 1860 6944 1912 6996
rect 2228 6944 2280 6996
rect 2688 6944 2740 6996
rect 4620 6944 4672 6996
rect 5264 6944 5316 6996
rect 1216 6808 1268 6860
rect 2044 6808 2096 6860
rect 3332 6808 3384 6860
rect 3608 6851 3660 6860
rect 3608 6817 3617 6851
rect 3617 6817 3651 6851
rect 3651 6817 3660 6851
rect 3608 6808 3660 6817
rect 3700 6851 3752 6860
rect 3700 6817 3709 6851
rect 3709 6817 3743 6851
rect 3743 6817 3752 6851
rect 3700 6808 3752 6817
rect 4068 6851 4120 6860
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4160 6808 4212 6860
rect 5172 6876 5224 6928
rect 7656 6987 7708 6996
rect 7656 6953 7665 6987
rect 7665 6953 7699 6987
rect 7699 6953 7708 6987
rect 7656 6944 7708 6953
rect 8944 6944 8996 6996
rect 4804 6808 4856 6860
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 2320 6740 2372 6792
rect 2780 6740 2832 6792
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 6092 6808 6144 6860
rect 6644 6876 6696 6928
rect 2964 6672 3016 6724
rect 3608 6672 3660 6724
rect 3056 6604 3108 6656
rect 3424 6604 3476 6656
rect 4160 6672 4212 6724
rect 4068 6604 4120 6656
rect 5816 6740 5868 6792
rect 6552 6808 6604 6860
rect 9220 6876 9272 6928
rect 6736 6740 6788 6792
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 6644 6672 6696 6724
rect 6276 6604 6328 6656
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 9496 6944 9548 6996
rect 9772 6876 9824 6928
rect 10600 6876 10652 6928
rect 12256 6876 12308 6928
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 10140 6808 10192 6860
rect 10508 6808 10560 6860
rect 11152 6808 11204 6860
rect 8116 6672 8168 6724
rect 9312 6740 9364 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 10232 6672 10284 6724
rect 8300 6604 8352 6656
rect 8760 6604 8812 6656
rect 10048 6604 10100 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11244 6672 11296 6724
rect 11796 6851 11848 6860
rect 11796 6817 11805 6851
rect 11805 6817 11839 6851
rect 11839 6817 11848 6851
rect 11796 6808 11848 6817
rect 12348 6808 12400 6860
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 12900 6944 12952 6996
rect 12992 6944 13044 6996
rect 14464 6944 14516 6996
rect 14648 6944 14700 6996
rect 15476 6944 15528 6996
rect 13452 6876 13504 6928
rect 13728 6876 13780 6928
rect 12992 6851 13044 6860
rect 12992 6817 13001 6851
rect 13001 6817 13035 6851
rect 13035 6817 13044 6851
rect 12992 6808 13044 6817
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 13084 6740 13136 6792
rect 11980 6672 12032 6724
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 16120 6876 16172 6928
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 16120 6740 16172 6792
rect 16488 6851 16540 6860
rect 16488 6817 16497 6851
rect 16497 6817 16531 6851
rect 16531 6817 16540 6851
rect 16488 6808 16540 6817
rect 17776 6876 17828 6928
rect 18696 6876 18748 6928
rect 19524 6876 19576 6928
rect 21180 6944 21232 6996
rect 23020 6944 23072 6996
rect 17408 6808 17460 6860
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 17684 6851 17736 6860
rect 17684 6817 17693 6851
rect 17693 6817 17727 6851
rect 17727 6817 17736 6851
rect 17684 6808 17736 6817
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 17960 6808 18012 6860
rect 18236 6808 18288 6860
rect 18880 6808 18932 6860
rect 19248 6740 19300 6792
rect 12808 6604 12860 6656
rect 14096 6604 14148 6656
rect 15660 6604 15712 6656
rect 17040 6715 17092 6724
rect 17040 6681 17049 6715
rect 17049 6681 17083 6715
rect 17083 6681 17092 6715
rect 17040 6672 17092 6681
rect 17500 6672 17552 6724
rect 19616 6808 19668 6860
rect 19708 6740 19760 6792
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 18696 6604 18748 6656
rect 19616 6672 19668 6724
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20444 6808 20496 6860
rect 20628 6808 20680 6860
rect 21456 6876 21508 6928
rect 21640 6876 21692 6928
rect 22652 6876 22704 6928
rect 21180 6740 21232 6792
rect 21732 6808 21784 6860
rect 22284 6851 22336 6860
rect 22284 6817 22293 6851
rect 22293 6817 22327 6851
rect 22327 6817 22336 6851
rect 22284 6808 22336 6817
rect 22376 6851 22428 6860
rect 22376 6817 22385 6851
rect 22385 6817 22419 6851
rect 22419 6817 22428 6851
rect 22376 6808 22428 6817
rect 23388 6944 23440 6996
rect 23480 6944 23532 6996
rect 24584 6987 24636 6996
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 22744 6740 22796 6792
rect 24124 6876 24176 6928
rect 23388 6740 23440 6792
rect 22836 6672 22888 6724
rect 23020 6672 23072 6724
rect 23664 6808 23716 6860
rect 24584 6953 24601 6987
rect 24601 6953 24636 6987
rect 24584 6944 24636 6953
rect 25412 6944 25464 6996
rect 25780 6944 25832 6996
rect 29828 6944 29880 6996
rect 24768 6919 24820 6928
rect 24768 6885 24777 6919
rect 24777 6885 24811 6919
rect 24811 6885 24820 6919
rect 24768 6876 24820 6885
rect 23664 6672 23716 6724
rect 24676 6808 24728 6860
rect 24952 6740 25004 6792
rect 26884 6876 26936 6928
rect 28356 6876 28408 6928
rect 25320 6808 25372 6860
rect 25780 6808 25832 6860
rect 25596 6740 25648 6792
rect 26332 6808 26384 6860
rect 28540 6851 28592 6860
rect 28540 6817 28549 6851
rect 28549 6817 28583 6851
rect 28583 6817 28592 6851
rect 28540 6808 28592 6817
rect 28632 6851 28684 6860
rect 28632 6817 28641 6851
rect 28641 6817 28675 6851
rect 28675 6817 28684 6851
rect 28632 6808 28684 6817
rect 29000 6876 29052 6928
rect 29460 6851 29512 6860
rect 29460 6817 29469 6851
rect 29469 6817 29503 6851
rect 29503 6817 29512 6851
rect 29460 6808 29512 6817
rect 30104 6851 30156 6860
rect 30104 6817 30113 6851
rect 30113 6817 30147 6851
rect 30147 6817 30156 6851
rect 30104 6808 30156 6817
rect 30656 6808 30708 6860
rect 30840 6808 30892 6860
rect 31024 6808 31076 6860
rect 26148 6740 26200 6792
rect 27344 6740 27396 6792
rect 24308 6672 24360 6724
rect 24400 6715 24452 6724
rect 24400 6681 24409 6715
rect 24409 6681 24443 6715
rect 24443 6681 24452 6715
rect 24400 6672 24452 6681
rect 27068 6672 27120 6724
rect 19248 6604 19300 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 20720 6604 20772 6656
rect 21732 6647 21784 6656
rect 21732 6613 21741 6647
rect 21741 6613 21775 6647
rect 21775 6613 21784 6647
rect 21732 6604 21784 6613
rect 21916 6604 21968 6656
rect 22100 6604 22152 6656
rect 23204 6604 23256 6656
rect 23388 6604 23440 6656
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 24860 6604 24912 6656
rect 25228 6604 25280 6656
rect 25596 6604 25648 6656
rect 28172 6672 28224 6724
rect 28908 6672 28960 6724
rect 29000 6647 29052 6656
rect 29000 6613 29009 6647
rect 29009 6613 29043 6647
rect 29043 6613 29052 6647
rect 29000 6604 29052 6613
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 11436 6502 11488 6554
rect 11500 6502 11552 6554
rect 11564 6502 11616 6554
rect 11628 6502 11680 6554
rect 11692 6502 11744 6554
rect 19210 6502 19262 6554
rect 19274 6502 19326 6554
rect 19338 6502 19390 6554
rect 19402 6502 19454 6554
rect 19466 6502 19518 6554
rect 26984 6502 27036 6554
rect 27048 6502 27100 6554
rect 27112 6502 27164 6554
rect 27176 6502 27228 6554
rect 27240 6502 27292 6554
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 2872 6443 2924 6452
rect 2872 6409 2881 6443
rect 2881 6409 2915 6443
rect 2915 6409 2924 6443
rect 2872 6400 2924 6409
rect 8024 6400 8076 6452
rect 8300 6400 8352 6452
rect 10140 6400 10192 6452
rect 1952 6332 2004 6384
rect 1676 6264 1728 6316
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 11060 6400 11112 6452
rect 11704 6400 11756 6452
rect 11796 6400 11848 6452
rect 13728 6332 13780 6384
rect 15292 6400 15344 6452
rect 15384 6400 15436 6452
rect 16120 6443 16172 6452
rect 16120 6409 16129 6443
rect 16129 6409 16163 6443
rect 16163 6409 16172 6443
rect 16120 6400 16172 6409
rect 17408 6400 17460 6452
rect 17960 6400 18012 6452
rect 18328 6400 18380 6452
rect 19800 6400 19852 6452
rect 20444 6400 20496 6452
rect 20628 6400 20680 6452
rect 22008 6400 22060 6452
rect 22284 6400 22336 6452
rect 24032 6443 24084 6452
rect 24032 6409 24041 6443
rect 24041 6409 24075 6443
rect 24075 6409 24084 6443
rect 24032 6400 24084 6409
rect 24584 6400 24636 6452
rect 24860 6400 24912 6452
rect 25872 6400 25924 6452
rect 27344 6443 27396 6452
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 28264 6400 28316 6452
rect 5356 6264 5408 6316
rect 3332 6196 3384 6248
rect 3608 6196 3660 6248
rect 3976 6128 4028 6180
rect 4620 6196 4672 6248
rect 6644 6264 6696 6316
rect 8668 6264 8720 6316
rect 6552 6196 6604 6248
rect 4988 6128 5040 6180
rect 5172 6060 5224 6112
rect 5816 6060 5868 6112
rect 6000 6171 6052 6180
rect 6000 6137 6009 6171
rect 6009 6137 6043 6171
rect 6043 6137 6052 6171
rect 6000 6128 6052 6137
rect 6276 6128 6328 6180
rect 7288 6196 7340 6248
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 8024 6196 8076 6248
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 10508 6196 10560 6248
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 11980 6196 12032 6248
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 12900 6264 12952 6273
rect 12992 6196 13044 6248
rect 13084 6239 13136 6248
rect 13084 6205 13093 6239
rect 13093 6205 13127 6239
rect 13127 6205 13136 6239
rect 13084 6196 13136 6205
rect 12716 6128 12768 6180
rect 13452 6196 13504 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14832 6307 14884 6316
rect 14280 6196 14332 6248
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 18236 6332 18288 6384
rect 22560 6332 22612 6384
rect 23480 6332 23532 6384
rect 24768 6332 24820 6384
rect 24400 6264 24452 6316
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 15016 6196 15068 6248
rect 15200 6196 15252 6248
rect 16120 6196 16172 6248
rect 16396 6196 16448 6248
rect 16488 6239 16540 6248
rect 16488 6205 16497 6239
rect 16497 6205 16531 6239
rect 16531 6205 16540 6239
rect 16488 6196 16540 6205
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 15384 6128 15436 6180
rect 16764 6128 16816 6180
rect 10324 6060 10376 6112
rect 10600 6060 10652 6112
rect 11152 6060 11204 6112
rect 11244 6060 11296 6112
rect 11520 6060 11572 6112
rect 11796 6060 11848 6112
rect 12992 6060 13044 6112
rect 13268 6103 13320 6112
rect 13268 6069 13277 6103
rect 13277 6069 13311 6103
rect 13311 6069 13320 6103
rect 13268 6060 13320 6069
rect 13728 6060 13780 6112
rect 19156 6196 19208 6248
rect 18512 6128 18564 6180
rect 18788 6128 18840 6180
rect 19432 6196 19484 6248
rect 21272 6196 21324 6248
rect 21916 6239 21968 6248
rect 21916 6205 21925 6239
rect 21925 6205 21959 6239
rect 21959 6205 21968 6239
rect 21916 6196 21968 6205
rect 18880 6060 18932 6112
rect 19156 6060 19208 6112
rect 20076 6128 20128 6180
rect 21088 6128 21140 6180
rect 23756 6196 23808 6248
rect 25780 6332 25832 6384
rect 26148 6332 26200 6384
rect 30656 6332 30708 6384
rect 26608 6264 26660 6316
rect 24216 6171 24268 6180
rect 24216 6137 24225 6171
rect 24225 6137 24259 6171
rect 24259 6137 24268 6171
rect 24216 6128 24268 6137
rect 24676 6128 24728 6180
rect 25320 6196 25372 6248
rect 25780 6239 25832 6248
rect 25780 6205 25789 6239
rect 25789 6205 25823 6239
rect 25823 6205 25832 6239
rect 25780 6196 25832 6205
rect 26884 6196 26936 6248
rect 29000 6307 29052 6316
rect 29000 6273 29009 6307
rect 29009 6273 29043 6307
rect 29043 6273 29052 6307
rect 29000 6264 29052 6273
rect 28448 6196 28500 6248
rect 29184 6239 29236 6248
rect 29184 6205 29193 6239
rect 29193 6205 29227 6239
rect 29227 6205 29236 6239
rect 29184 6196 29236 6205
rect 29828 6307 29880 6316
rect 29828 6273 29837 6307
rect 29837 6273 29871 6307
rect 29871 6273 29880 6307
rect 29828 6264 29880 6273
rect 30012 6307 30064 6316
rect 30012 6273 30021 6307
rect 30021 6273 30055 6307
rect 30055 6273 30064 6307
rect 30012 6264 30064 6273
rect 30104 6307 30156 6316
rect 30104 6273 30113 6307
rect 30113 6273 30147 6307
rect 30147 6273 30156 6307
rect 30104 6264 30156 6273
rect 25412 6128 25464 6180
rect 26976 6128 27028 6180
rect 30288 6239 30340 6248
rect 30288 6205 30297 6239
rect 30297 6205 30331 6239
rect 30331 6205 30340 6239
rect 30288 6196 30340 6205
rect 20168 6060 20220 6112
rect 20260 6060 20312 6112
rect 22744 6060 22796 6112
rect 23848 6103 23900 6112
rect 23848 6069 23857 6103
rect 23857 6069 23891 6103
rect 23891 6069 23900 6103
rect 23848 6060 23900 6069
rect 24032 6103 24084 6112
rect 24032 6069 24059 6103
rect 24059 6069 24084 6103
rect 24032 6060 24084 6069
rect 29000 6060 29052 6112
rect 30012 6060 30064 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 12096 5958 12148 6010
rect 12160 5958 12212 6010
rect 12224 5958 12276 6010
rect 12288 5958 12340 6010
rect 12352 5958 12404 6010
rect 19870 5958 19922 6010
rect 19934 5958 19986 6010
rect 19998 5958 20050 6010
rect 20062 5958 20114 6010
rect 20126 5958 20178 6010
rect 27644 5958 27696 6010
rect 27708 5958 27760 6010
rect 27772 5958 27824 6010
rect 27836 5958 27888 6010
rect 27900 5958 27952 6010
rect 940 5856 992 5908
rect 1952 5831 2004 5840
rect 1952 5797 1961 5831
rect 1961 5797 1995 5831
rect 1995 5797 2004 5831
rect 1952 5788 2004 5797
rect 2136 5788 2188 5840
rect 3516 5788 3568 5840
rect 1308 5763 1360 5772
rect 1308 5729 1317 5763
rect 1317 5729 1351 5763
rect 1351 5729 1360 5763
rect 1308 5720 1360 5729
rect 1676 5720 1728 5772
rect 3056 5763 3108 5772
rect 1584 5652 1636 5704
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 3056 5720 3108 5729
rect 3240 5720 3292 5772
rect 4068 5788 4120 5840
rect 2228 5652 2280 5704
rect 3424 5652 3476 5704
rect 4712 5856 4764 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 6644 5856 6696 5908
rect 7288 5856 7340 5908
rect 7380 5856 7432 5908
rect 7564 5856 7616 5908
rect 5816 5788 5868 5840
rect 4804 5763 4856 5772
rect 4804 5729 4810 5763
rect 4810 5729 4844 5763
rect 4844 5729 4856 5763
rect 4804 5720 4856 5729
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 5264 5763 5316 5772
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 6552 5831 6604 5840
rect 6552 5797 6561 5831
rect 6561 5797 6595 5831
rect 6595 5797 6604 5831
rect 6552 5788 6604 5797
rect 7012 5788 7064 5840
rect 7748 5788 7800 5840
rect 8576 5856 8628 5908
rect 9404 5856 9456 5908
rect 9220 5831 9272 5840
rect 9220 5797 9229 5831
rect 9229 5797 9263 5831
rect 9263 5797 9272 5831
rect 9220 5788 9272 5797
rect 10140 5788 10192 5840
rect 10324 5788 10376 5840
rect 11888 5856 11940 5908
rect 11980 5856 12032 5908
rect 13452 5856 13504 5908
rect 13544 5856 13596 5908
rect 13728 5856 13780 5908
rect 13912 5856 13964 5908
rect 15292 5856 15344 5908
rect 16488 5856 16540 5908
rect 18236 5856 18288 5908
rect 19064 5856 19116 5908
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9312 5720 9364 5772
rect 9404 5763 9456 5772
rect 9404 5729 9412 5763
rect 9412 5729 9446 5763
rect 9446 5729 9456 5763
rect 9404 5720 9456 5729
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 9772 5720 9824 5772
rect 10600 5720 10652 5772
rect 11152 5763 11204 5772
rect 6644 5652 6696 5704
rect 7104 5652 7156 5704
rect 7748 5652 7800 5704
rect 2504 5627 2556 5636
rect 2504 5593 2513 5627
rect 2513 5593 2547 5627
rect 2547 5593 2556 5627
rect 2504 5584 2556 5593
rect 9220 5584 9272 5636
rect 9680 5652 9732 5704
rect 10784 5652 10836 5704
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11152 5729 11161 5763
rect 11161 5729 11195 5763
rect 11195 5729 11204 5763
rect 11152 5720 11204 5729
rect 11336 5788 11388 5840
rect 12072 5788 12124 5840
rect 12440 5788 12492 5840
rect 13268 5788 13320 5840
rect 15384 5788 15436 5840
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11704 5720 11756 5772
rect 18604 5788 18656 5840
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 12072 5652 12124 5704
rect 15752 5652 15804 5704
rect 8576 5516 8628 5568
rect 9036 5516 9088 5568
rect 11796 5584 11848 5636
rect 10784 5516 10836 5568
rect 14556 5584 14608 5636
rect 15660 5584 15712 5636
rect 16856 5720 16908 5772
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 17960 5763 18012 5772
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 17776 5652 17828 5704
rect 18512 5763 18564 5772
rect 18512 5729 18521 5763
rect 18521 5729 18555 5763
rect 18555 5729 18564 5763
rect 18512 5720 18564 5729
rect 18972 5720 19024 5772
rect 21180 5856 21232 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 21640 5856 21692 5908
rect 24492 5856 24544 5908
rect 25320 5856 25372 5908
rect 27436 5856 27488 5908
rect 28448 5856 28500 5908
rect 29184 5856 29236 5908
rect 26976 5831 27028 5840
rect 20076 5763 20128 5772
rect 20076 5729 20085 5763
rect 20085 5729 20119 5763
rect 20119 5729 20128 5763
rect 20076 5720 20128 5729
rect 20352 5763 20404 5772
rect 20352 5729 20361 5763
rect 20361 5729 20395 5763
rect 20395 5729 20404 5763
rect 20352 5720 20404 5729
rect 21548 5763 21600 5772
rect 21548 5729 21557 5763
rect 21557 5729 21591 5763
rect 21591 5729 21600 5763
rect 21548 5720 21600 5729
rect 21824 5763 21876 5772
rect 21824 5729 21833 5763
rect 21833 5729 21867 5763
rect 21867 5729 21876 5763
rect 21824 5720 21876 5729
rect 22008 5763 22060 5772
rect 22008 5729 22017 5763
rect 22017 5729 22051 5763
rect 22051 5729 22060 5763
rect 22008 5720 22060 5729
rect 19340 5652 19392 5704
rect 19432 5652 19484 5704
rect 21272 5652 21324 5704
rect 22284 5720 22336 5772
rect 19064 5584 19116 5636
rect 12348 5516 12400 5568
rect 21732 5627 21784 5636
rect 21732 5593 21741 5627
rect 21741 5593 21775 5627
rect 21775 5593 21784 5627
rect 21732 5584 21784 5593
rect 24768 5720 24820 5772
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 25320 5652 25372 5704
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25412 5652 25464 5661
rect 25596 5720 25648 5772
rect 25872 5720 25924 5772
rect 25964 5763 26016 5772
rect 25964 5729 25973 5763
rect 25973 5729 26007 5763
rect 26007 5729 26016 5763
rect 25964 5720 26016 5729
rect 26332 5720 26384 5772
rect 26976 5797 26985 5831
rect 26985 5797 27019 5831
rect 27019 5797 27028 5831
rect 26976 5788 27028 5797
rect 26884 5763 26936 5772
rect 26884 5729 26893 5763
rect 26893 5729 26927 5763
rect 26927 5729 26936 5763
rect 26884 5720 26936 5729
rect 27344 5788 27396 5840
rect 30288 5788 30340 5840
rect 27712 5720 27764 5772
rect 27988 5720 28040 5772
rect 26792 5652 26844 5704
rect 27528 5652 27580 5704
rect 29092 5720 29144 5772
rect 29460 5720 29512 5772
rect 29552 5763 29604 5772
rect 29552 5729 29561 5763
rect 29561 5729 29595 5763
rect 29595 5729 29604 5763
rect 29552 5720 29604 5729
rect 29828 5763 29880 5772
rect 29828 5729 29837 5763
rect 29837 5729 29871 5763
rect 29871 5729 29880 5763
rect 29828 5720 29880 5729
rect 23572 5584 23624 5636
rect 20076 5516 20128 5568
rect 21640 5516 21692 5568
rect 22468 5559 22520 5568
rect 22468 5525 22477 5559
rect 22477 5525 22511 5559
rect 22511 5525 22520 5559
rect 22468 5516 22520 5525
rect 23756 5516 23808 5568
rect 25504 5584 25556 5636
rect 26884 5584 26936 5636
rect 29276 5627 29328 5636
rect 29276 5593 29285 5627
rect 29285 5593 29319 5627
rect 29319 5593 29328 5627
rect 29276 5584 29328 5593
rect 26056 5516 26108 5568
rect 28448 5516 28500 5568
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 11436 5414 11488 5466
rect 11500 5414 11552 5466
rect 11564 5414 11616 5466
rect 11628 5414 11680 5466
rect 11692 5414 11744 5466
rect 19210 5414 19262 5466
rect 19274 5414 19326 5466
rect 19338 5414 19390 5466
rect 19402 5414 19454 5466
rect 19466 5414 19518 5466
rect 26984 5414 27036 5466
rect 27048 5414 27100 5466
rect 27112 5414 27164 5466
rect 27176 5414 27228 5466
rect 27240 5414 27292 5466
rect 6276 5312 6328 5364
rect 2504 5287 2556 5296
rect 2504 5253 2513 5287
rect 2513 5253 2547 5287
rect 2547 5253 2556 5287
rect 2504 5244 2556 5253
rect 4988 5244 5040 5296
rect 10416 5312 10468 5364
rect 12440 5312 12492 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 12900 5312 12952 5364
rect 14832 5312 14884 5364
rect 7840 5287 7892 5296
rect 7840 5253 7849 5287
rect 7849 5253 7883 5287
rect 7883 5253 7892 5287
rect 7840 5244 7892 5253
rect 11244 5244 11296 5296
rect 11704 5244 11756 5296
rect 1308 5108 1360 5160
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 7012 5176 7064 5228
rect 4160 5108 4212 5160
rect 5080 5108 5132 5160
rect 6000 5108 6052 5160
rect 6184 5108 6236 5160
rect 3608 5040 3660 5092
rect 6644 5151 6696 5160
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 6644 5108 6696 5117
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 7472 5108 7524 5160
rect 9680 5176 9732 5228
rect 11152 5176 11204 5228
rect 12532 5176 12584 5228
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 13176 5176 13228 5228
rect 14924 5287 14976 5296
rect 14924 5253 14933 5287
rect 14933 5253 14967 5287
rect 14967 5253 14976 5287
rect 14924 5244 14976 5253
rect 15936 5287 15988 5296
rect 15936 5253 15945 5287
rect 15945 5253 15979 5287
rect 15979 5253 15988 5287
rect 15936 5244 15988 5253
rect 17500 5312 17552 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 21548 5312 21600 5364
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 20352 5244 20404 5296
rect 21088 5244 21140 5296
rect 23756 5244 23808 5296
rect 25320 5312 25372 5364
rect 25780 5312 25832 5364
rect 25872 5312 25924 5364
rect 24124 5287 24176 5296
rect 24124 5253 24133 5287
rect 24133 5253 24167 5287
rect 24167 5253 24176 5287
rect 24124 5244 24176 5253
rect 24400 5244 24452 5296
rect 24768 5244 24820 5296
rect 26332 5244 26384 5296
rect 26608 5355 26660 5364
rect 26608 5321 26617 5355
rect 26617 5321 26651 5355
rect 26651 5321 26660 5355
rect 26608 5312 26660 5321
rect 29828 5312 29880 5364
rect 15108 5176 15160 5228
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 9588 5108 9640 5160
rect 11336 5108 11388 5160
rect 11704 5108 11756 5160
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 4252 4972 4304 5024
rect 6276 4972 6328 5024
rect 6460 4972 6512 5024
rect 6552 4972 6604 5024
rect 9404 5040 9456 5092
rect 13636 5151 13688 5160
rect 13636 5117 13678 5151
rect 13678 5117 13688 5151
rect 13636 5108 13688 5117
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 14832 5151 14884 5160
rect 14832 5117 14841 5151
rect 14841 5117 14875 5151
rect 14875 5117 14884 5151
rect 14832 5108 14884 5117
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 16028 5151 16080 5160
rect 16028 5117 16037 5151
rect 16037 5117 16071 5151
rect 16071 5117 16080 5151
rect 16028 5108 16080 5117
rect 16120 5108 16172 5160
rect 18420 5108 18472 5160
rect 18696 5151 18748 5160
rect 18696 5117 18705 5151
rect 18705 5117 18739 5151
rect 18739 5117 18748 5151
rect 18696 5108 18748 5117
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 18880 5108 18932 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 20260 5108 20312 5160
rect 20352 5108 20404 5160
rect 23112 5176 23164 5228
rect 24676 5176 24728 5228
rect 25964 5176 26016 5228
rect 20904 5151 20956 5160
rect 20904 5117 20913 5151
rect 20913 5117 20947 5151
rect 20947 5117 20956 5151
rect 20904 5108 20956 5117
rect 21456 5151 21508 5160
rect 21456 5117 21465 5151
rect 21465 5117 21499 5151
rect 21499 5117 21508 5151
rect 21456 5108 21508 5117
rect 22652 5108 22704 5160
rect 24216 5108 24268 5160
rect 24400 5151 24452 5160
rect 24400 5117 24409 5151
rect 24409 5117 24443 5151
rect 24443 5117 24452 5151
rect 24400 5108 24452 5117
rect 24492 5108 24544 5160
rect 11152 4972 11204 5024
rect 11336 4972 11388 5024
rect 11704 4972 11756 5024
rect 11888 4972 11940 5024
rect 12900 4972 12952 5024
rect 14280 4972 14332 5024
rect 15660 5083 15712 5092
rect 15660 5049 15669 5083
rect 15669 5049 15703 5083
rect 15703 5049 15712 5083
rect 15660 5040 15712 5049
rect 17960 5040 18012 5092
rect 15752 4972 15804 5024
rect 16396 4972 16448 5024
rect 21272 5015 21324 5024
rect 21272 4981 21281 5015
rect 21281 4981 21315 5015
rect 21315 4981 21324 5015
rect 21272 4972 21324 4981
rect 24584 5015 24636 5024
rect 24584 4981 24593 5015
rect 24593 4981 24627 5015
rect 24627 4981 24636 5015
rect 24584 4972 24636 4981
rect 25044 4972 25096 5024
rect 25412 5151 25464 5160
rect 25412 5117 25421 5151
rect 25421 5117 25455 5151
rect 25455 5117 25464 5151
rect 25412 5108 25464 5117
rect 26608 5108 26660 5160
rect 28080 5244 28132 5296
rect 29552 5176 29604 5228
rect 27712 5151 27764 5160
rect 27712 5117 27721 5151
rect 27721 5117 27755 5151
rect 27755 5117 27764 5151
rect 27712 5108 27764 5117
rect 29276 5151 29328 5160
rect 29276 5117 29285 5151
rect 29285 5117 29319 5151
rect 29319 5117 29328 5151
rect 29276 5108 29328 5117
rect 29460 5108 29512 5160
rect 30840 5151 30892 5160
rect 30840 5117 30849 5151
rect 30849 5117 30883 5151
rect 30883 5117 30892 5151
rect 30840 5108 30892 5117
rect 30288 5040 30340 5092
rect 28540 5015 28592 5024
rect 28540 4981 28549 5015
rect 28549 4981 28583 5015
rect 28583 4981 28592 5015
rect 28540 4972 28592 4981
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 12096 4870 12148 4922
rect 12160 4870 12212 4922
rect 12224 4870 12276 4922
rect 12288 4870 12340 4922
rect 12352 4870 12404 4922
rect 19870 4870 19922 4922
rect 19934 4870 19986 4922
rect 19998 4870 20050 4922
rect 20062 4870 20114 4922
rect 20126 4870 20178 4922
rect 27644 4870 27696 4922
rect 27708 4870 27760 4922
rect 27772 4870 27824 4922
rect 27836 4870 27888 4922
rect 27900 4870 27952 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 3148 4768 3200 4820
rect 4252 4768 4304 4820
rect 4988 4811 5040 4820
rect 4988 4777 4997 4811
rect 4997 4777 5031 4811
rect 5031 4777 5040 4811
rect 4988 4768 5040 4777
rect 5816 4811 5868 4820
rect 5816 4777 5825 4811
rect 5825 4777 5859 4811
rect 5859 4777 5868 4811
rect 5816 4768 5868 4777
rect 6920 4768 6972 4820
rect 2044 4743 2096 4752
rect 2044 4709 2053 4743
rect 2053 4709 2087 4743
rect 2087 4709 2096 4743
rect 2044 4700 2096 4709
rect 7564 4700 7616 4752
rect 9680 4700 9732 4752
rect 10416 4700 10468 4752
rect 12532 4768 12584 4820
rect 13084 4768 13136 4820
rect 15384 4768 15436 4820
rect 16396 4768 16448 4820
rect 17224 4811 17276 4820
rect 17224 4777 17233 4811
rect 17233 4777 17267 4811
rect 17267 4777 17276 4811
rect 17224 4768 17276 4777
rect 17408 4768 17460 4820
rect 18604 4768 18656 4820
rect 18788 4768 18840 4820
rect 21732 4768 21784 4820
rect 22192 4768 22244 4820
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 29368 4811 29420 4820
rect 29368 4777 29377 4811
rect 29377 4777 29411 4811
rect 29411 4777 29420 4811
rect 29368 4768 29420 4777
rect 1308 4632 1360 4684
rect 2780 4632 2832 4684
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 4160 4632 4212 4684
rect 3608 4564 3660 4616
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6092 4632 6144 4684
rect 6460 4632 6512 4684
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 7840 4632 7892 4684
rect 9404 4632 9456 4684
rect 9496 4675 9548 4684
rect 9496 4641 9505 4675
rect 9505 4641 9539 4675
rect 9539 4641 9548 4675
rect 9496 4632 9548 4641
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 8392 4564 8444 4616
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 10968 4632 11020 4684
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 5172 4428 5224 4480
rect 8024 4471 8076 4480
rect 8024 4437 8033 4471
rect 8033 4437 8067 4471
rect 8067 4437 8076 4471
rect 8024 4428 8076 4437
rect 9772 4428 9824 4480
rect 10968 4496 11020 4548
rect 11152 4564 11204 4616
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12532 4632 12584 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 17316 4700 17368 4752
rect 18420 4700 18472 4752
rect 12808 4496 12860 4548
rect 13360 4564 13412 4616
rect 17132 4632 17184 4684
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 18328 4675 18380 4684
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 18604 4632 18656 4684
rect 19708 4700 19760 4752
rect 19984 4700 20036 4752
rect 20352 4743 20404 4752
rect 20352 4709 20361 4743
rect 20361 4709 20395 4743
rect 20395 4709 20404 4743
rect 20352 4700 20404 4709
rect 21088 4700 21140 4752
rect 16212 4564 16264 4616
rect 17408 4564 17460 4616
rect 20536 4675 20588 4684
rect 20536 4641 20575 4675
rect 20575 4641 20588 4675
rect 20536 4632 20588 4641
rect 20812 4632 20864 4684
rect 21548 4564 21600 4616
rect 10324 4428 10376 4480
rect 10416 4428 10468 4480
rect 11796 4428 11848 4480
rect 15384 4428 15436 4480
rect 16856 4428 16908 4480
rect 16948 4471 17000 4480
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 18880 4428 18932 4480
rect 20720 4496 20772 4548
rect 22744 4675 22796 4684
rect 22744 4641 22753 4675
rect 22753 4641 22787 4675
rect 22787 4641 22796 4675
rect 22744 4632 22796 4641
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 23940 4632 23992 4684
rect 25780 4700 25832 4752
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 25136 4632 25188 4684
rect 25320 4632 25372 4684
rect 26700 4607 26752 4616
rect 26700 4573 26709 4607
rect 26709 4573 26743 4607
rect 26743 4573 26752 4607
rect 26700 4564 26752 4573
rect 27436 4675 27488 4684
rect 27436 4641 27445 4675
rect 27445 4641 27479 4675
rect 27479 4641 27488 4675
rect 27436 4632 27488 4641
rect 30012 4632 30064 4684
rect 28908 4496 28960 4548
rect 19524 4428 19576 4480
rect 19616 4428 19668 4480
rect 28540 4428 28592 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 11436 4326 11488 4378
rect 11500 4326 11552 4378
rect 11564 4326 11616 4378
rect 11628 4326 11680 4378
rect 11692 4326 11744 4378
rect 19210 4326 19262 4378
rect 19274 4326 19326 4378
rect 19338 4326 19390 4378
rect 19402 4326 19454 4378
rect 19466 4326 19518 4378
rect 26984 4326 27036 4378
rect 27048 4326 27100 4378
rect 27112 4326 27164 4378
rect 27176 4326 27228 4378
rect 27240 4326 27292 4378
rect 3700 4224 3752 4276
rect 4252 4224 4304 4276
rect 7656 4224 7708 4276
rect 7840 4224 7892 4276
rect 8024 4224 8076 4276
rect 10140 4224 10192 4276
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 12624 4267 12676 4276
rect 12624 4233 12633 4267
rect 12633 4233 12667 4267
rect 12667 4233 12676 4267
rect 12624 4224 12676 4233
rect 16212 4224 16264 4276
rect 16856 4224 16908 4276
rect 19984 4224 20036 4276
rect 20628 4224 20680 4276
rect 6000 4156 6052 4208
rect 12900 4156 12952 4208
rect 6184 4088 6236 4140
rect 6368 4088 6420 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 3516 4020 3568 4072
rect 4160 4063 4212 4072
rect 4160 4029 4169 4063
rect 4169 4029 4203 4063
rect 4203 4029 4212 4063
rect 4160 4020 4212 4029
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 6828 4020 6880 4072
rect 8208 4088 8260 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 7656 4020 7708 4072
rect 8116 4020 8168 4072
rect 3424 3952 3476 4004
rect 5080 3952 5132 4004
rect 7380 3952 7432 4004
rect 9680 4088 9732 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 9496 4020 9548 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 13452 4088 13504 4140
rect 17132 4156 17184 4208
rect 18236 4156 18288 4208
rect 20812 4156 20864 4208
rect 14188 4088 14240 4140
rect 19616 4088 19668 4140
rect 19800 4131 19852 4140
rect 19800 4097 19809 4131
rect 19809 4097 19843 4131
rect 19843 4097 19852 4131
rect 19800 4088 19852 4097
rect 20628 4131 20680 4140
rect 10416 4063 10468 4072
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 11060 4020 11112 4072
rect 12440 4020 12492 4072
rect 13176 4020 13228 4072
rect 13912 4020 13964 4072
rect 14832 4020 14884 4072
rect 3608 3884 3660 3936
rect 6276 3884 6328 3936
rect 10048 3884 10100 3936
rect 10232 3884 10284 3936
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 14464 3952 14516 4004
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 15476 4063 15528 4072
rect 15476 4029 15485 4063
rect 15485 4029 15519 4063
rect 15519 4029 15528 4063
rect 15476 4020 15528 4029
rect 15936 4063 15988 4072
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16120 3952 16172 4004
rect 17960 4020 18012 4072
rect 18972 4020 19024 4072
rect 17684 3884 17736 3936
rect 18420 3952 18472 4004
rect 19340 3995 19392 4004
rect 19340 3961 19349 3995
rect 19349 3961 19383 3995
rect 19383 3961 19392 3995
rect 19340 3952 19392 3961
rect 19708 4063 19760 4072
rect 19708 4029 19717 4063
rect 19717 4029 19751 4063
rect 19751 4029 19760 4063
rect 19708 4020 19760 4029
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 20720 4020 20772 4072
rect 21548 4020 21600 4072
rect 21824 4063 21876 4072
rect 21824 4029 21833 4063
rect 21833 4029 21867 4063
rect 21867 4029 21876 4063
rect 21824 4020 21876 4029
rect 22744 4224 22796 4276
rect 24676 4224 24728 4276
rect 22836 4156 22888 4208
rect 22928 4156 22980 4208
rect 25136 4156 25188 4208
rect 22468 4020 22520 4072
rect 21364 3995 21416 4004
rect 21364 3961 21373 3995
rect 21373 3961 21407 3995
rect 21407 3961 21416 3995
rect 21364 3952 21416 3961
rect 22284 3952 22336 4004
rect 22836 3952 22888 4004
rect 20536 3884 20588 3936
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 21824 3884 21876 3936
rect 22468 3927 22520 3936
rect 22468 3893 22477 3927
rect 22477 3893 22511 3927
rect 22511 3893 22520 3927
rect 23204 4063 23256 4072
rect 23204 4029 23213 4063
rect 23213 4029 23247 4063
rect 23247 4029 23256 4063
rect 23204 4020 23256 4029
rect 24216 4088 24268 4140
rect 25964 4131 26016 4140
rect 25964 4097 25973 4131
rect 25973 4097 26007 4131
rect 26007 4097 26016 4131
rect 25964 4088 26016 4097
rect 25044 3952 25096 4004
rect 25504 4020 25556 4072
rect 25872 4063 25924 4072
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 22468 3884 22520 3893
rect 24032 3884 24084 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 12096 3782 12148 3834
rect 12160 3782 12212 3834
rect 12224 3782 12276 3834
rect 12288 3782 12340 3834
rect 12352 3782 12404 3834
rect 19870 3782 19922 3834
rect 19934 3782 19986 3834
rect 19998 3782 20050 3834
rect 20062 3782 20114 3834
rect 20126 3782 20178 3834
rect 27644 3782 27696 3834
rect 27708 3782 27760 3834
rect 27772 3782 27824 3834
rect 27836 3782 27888 3834
rect 27900 3782 27952 3834
rect 3424 3680 3476 3732
rect 4896 3680 4948 3732
rect 3056 3612 3108 3664
rect 5724 3612 5776 3664
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 3332 3544 3384 3596
rect 4068 3544 4120 3596
rect 8392 3612 8444 3664
rect 6828 3544 6880 3596
rect 6552 3476 6604 3528
rect 12900 3587 12952 3596
rect 12900 3553 12909 3587
rect 12909 3553 12943 3587
rect 12943 3553 12952 3587
rect 12900 3544 12952 3553
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 2412 3408 2464 3460
rect 12348 3408 12400 3460
rect 12900 3408 12952 3460
rect 3700 3340 3752 3392
rect 10508 3383 10560 3392
rect 10508 3349 10517 3383
rect 10517 3349 10551 3383
rect 10551 3349 10560 3383
rect 10508 3340 10560 3349
rect 14004 3476 14056 3528
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 19340 3680 19392 3732
rect 20720 3680 20772 3732
rect 21272 3680 21324 3732
rect 31392 3680 31444 3732
rect 14464 3612 14516 3664
rect 22468 3612 22520 3664
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 14372 3587 14424 3596
rect 14372 3553 14382 3587
rect 14382 3553 14416 3587
rect 14416 3553 14424 3587
rect 14372 3544 14424 3553
rect 16488 3544 16540 3596
rect 21364 3544 21416 3596
rect 24860 3476 24912 3528
rect 14464 3408 14516 3460
rect 14740 3340 14792 3392
rect 15476 3340 15528 3392
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 11436 3238 11488 3290
rect 11500 3238 11552 3290
rect 11564 3238 11616 3290
rect 11628 3238 11680 3290
rect 11692 3238 11744 3290
rect 19210 3238 19262 3290
rect 19274 3238 19326 3290
rect 19338 3238 19390 3290
rect 19402 3238 19454 3290
rect 19466 3238 19518 3290
rect 26984 3238 27036 3290
rect 27048 3238 27100 3290
rect 27112 3238 27164 3290
rect 27176 3238 27228 3290
rect 27240 3238 27292 3290
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 12096 2694 12148 2746
rect 12160 2694 12212 2746
rect 12224 2694 12276 2746
rect 12288 2694 12340 2746
rect 12352 2694 12404 2746
rect 19870 2694 19922 2746
rect 19934 2694 19986 2746
rect 19998 2694 20050 2746
rect 20062 2694 20114 2746
rect 20126 2694 20178 2746
rect 27644 2694 27696 2746
rect 27708 2694 27760 2746
rect 27772 2694 27824 2746
rect 27836 2694 27888 2746
rect 27900 2694 27952 2746
rect 1032 2592 1084 2644
rect 24584 2592 24636 2644
rect 2228 2524 2280 2576
rect 24860 2524 24912 2576
rect 8300 2456 8352 2508
rect 23388 2456 23440 2508
rect 572 2388 624 2440
rect 11888 2388 11940 2440
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 11436 2150 11488 2202
rect 11500 2150 11552 2202
rect 11564 2150 11616 2202
rect 11628 2150 11680 2202
rect 11692 2150 11744 2202
rect 19210 2150 19262 2202
rect 19274 2150 19326 2202
rect 19338 2150 19390 2202
rect 19402 2150 19454 2202
rect 19466 2150 19518 2202
rect 26984 2150 27036 2202
rect 27048 2150 27100 2202
rect 27112 2150 27164 2202
rect 27176 2150 27228 2202
rect 27240 2150 27292 2202
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 12096 1606 12148 1658
rect 12160 1606 12212 1658
rect 12224 1606 12276 1658
rect 12288 1606 12340 1658
rect 12352 1606 12404 1658
rect 19870 1606 19922 1658
rect 19934 1606 19986 1658
rect 19998 1606 20050 1658
rect 20062 1606 20114 1658
rect 20126 1606 20178 1658
rect 27644 1606 27696 1658
rect 27708 1606 27760 1658
rect 27772 1606 27824 1658
rect 27836 1606 27888 1658
rect 27900 1606 27952 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 11436 1062 11488 1114
rect 11500 1062 11552 1114
rect 11564 1062 11616 1114
rect 11628 1062 11680 1114
rect 11692 1062 11744 1114
rect 19210 1062 19262 1114
rect 19274 1062 19326 1114
rect 19338 1062 19390 1114
rect 19402 1062 19454 1114
rect 19466 1062 19518 1114
rect 26984 1062 27036 1114
rect 27048 1062 27100 1114
rect 27112 1062 27164 1114
rect 27176 1062 27228 1114
rect 27240 1062 27292 1114
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 12096 518 12148 570
rect 12160 518 12212 570
rect 12224 518 12276 570
rect 12288 518 12340 570
rect 12352 518 12404 570
rect 19870 518 19922 570
rect 19934 518 19986 570
rect 19998 518 20050 570
rect 20062 518 20114 570
rect 20126 518 20178 570
rect 27644 518 27696 570
rect 27708 518 27760 570
rect 27772 518 27824 570
rect 27836 518 27888 570
rect 27900 518 27952 570
<< metal2 >>
rect 6550 22128 6606 22137
rect 6550 22063 6606 22072
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 6182 21720 6238 21729
rect 6182 21655 6184 21664
rect 6236 21655 6238 21664
rect 6184 21626 6236 21632
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 754 20360 810 20369
rect 754 20295 810 20304
rect 664 16720 716 16726
rect 664 16662 716 16668
rect 572 16176 624 16182
rect 572 16118 624 16124
rect 584 2446 612 16118
rect 676 6905 704 16662
rect 768 7993 796 20295
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 2318 19952 2374 19961
rect 2318 19887 2374 19896
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 1768 18148 1820 18154
rect 1768 18090 1820 18096
rect 1780 17746 1808 18090
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1308 17672 1360 17678
rect 1308 17614 1360 17620
rect 1216 16992 1268 16998
rect 1216 16934 1268 16940
rect 1228 15570 1256 16934
rect 1320 16046 1348 17614
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1308 16040 1360 16046
rect 1492 16040 1544 16046
rect 1308 15982 1360 15988
rect 1412 16000 1492 16028
rect 1216 15564 1268 15570
rect 1136 15524 1216 15552
rect 1032 14340 1084 14346
rect 1032 14282 1084 14288
rect 1044 13394 1072 14282
rect 1032 13388 1084 13394
rect 1032 13330 1084 13336
rect 940 13320 992 13326
rect 846 13288 902 13297
rect 940 13262 992 13268
rect 846 13223 902 13232
rect 754 7984 810 7993
rect 754 7919 810 7928
rect 662 6896 718 6905
rect 662 6831 718 6840
rect 860 6225 888 13223
rect 846 6216 902 6225
rect 846 6151 902 6160
rect 952 5914 980 13262
rect 1044 11898 1072 13330
rect 1136 12374 1164 15524
rect 1216 15506 1268 15512
rect 1216 15020 1268 15026
rect 1216 14962 1268 14968
rect 1124 12368 1176 12374
rect 1124 12310 1176 12316
rect 1032 11892 1084 11898
rect 1032 11834 1084 11840
rect 1122 11112 1178 11121
rect 1122 11047 1178 11056
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 1044 9178 1072 9454
rect 1032 9172 1084 9178
rect 1032 9114 1084 9120
rect 1030 8392 1086 8401
rect 1030 8327 1086 8336
rect 940 5908 992 5914
rect 940 5850 992 5856
rect 1044 2650 1072 8327
rect 1032 2644 1084 2650
rect 1032 2586 1084 2592
rect 572 2440 624 2446
rect 572 2382 624 2388
rect 1136 1465 1164 11047
rect 1228 9586 1256 14962
rect 1320 11218 1348 15982
rect 1412 11354 1440 16000
rect 1596 16017 1624 17070
rect 1688 16794 1716 17478
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1492 15982 1544 15988
rect 1582 16008 1638 16017
rect 1780 15994 1808 17682
rect 1872 16046 1900 17682
rect 1964 17649 1992 18158
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1950 17640 2006 17649
rect 1950 17575 2006 17584
rect 1964 16182 1992 17575
rect 2056 17134 2084 18022
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1952 16176 2004 16182
rect 1952 16118 2004 16124
rect 1582 15943 1638 15952
rect 1688 15966 1808 15994
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15552 1532 15846
rect 1596 15706 1624 15943
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1584 15564 1636 15570
rect 1504 15524 1584 15552
rect 1504 14958 1532 15524
rect 1584 15506 1636 15512
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 13462 1532 14894
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 1688 13274 1716 15966
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 13394 1808 15846
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 14482 1900 14758
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1952 14476 2004 14482
rect 2056 14464 2084 17070
rect 2148 17066 2176 18158
rect 2228 17808 2280 17814
rect 2226 17776 2228 17785
rect 2280 17776 2282 17785
rect 2226 17711 2282 17720
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2240 17542 2268 17614
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2136 17060 2188 17066
rect 2240 17048 2268 17478
rect 2332 17202 2360 19887
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3436 18834 3464 19110
rect 3896 18834 3924 19178
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 5460 18970 5488 19246
rect 6288 19230 6500 19258
rect 6288 19174 6316 19230
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6368 19168 6420 19174
rect 6368 19110 6420 19116
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3238 18728 3294 18737
rect 3238 18663 3240 18672
rect 3292 18663 3294 18672
rect 3240 18634 3292 18640
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2424 18154 2452 18226
rect 2412 18148 2464 18154
rect 2412 18090 2464 18096
rect 2516 17338 2544 18362
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2424 17134 2452 17274
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2240 17020 2360 17048
rect 2136 17002 2188 17008
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2004 14436 2084 14464
rect 1952 14418 2004 14424
rect 1872 13977 1900 14418
rect 1858 13968 1914 13977
rect 1858 13903 1914 13912
rect 1964 13394 1992 14418
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1952 13388 2004 13394
rect 2004 13348 2084 13376
rect 1952 13330 2004 13336
rect 1688 13246 1808 13274
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 12434 1532 13126
rect 1504 12406 1624 12434
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1308 11212 1360 11218
rect 1308 11154 1360 11160
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1320 9654 1348 10202
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1216 9580 1268 9586
rect 1216 9522 1268 9528
rect 1504 9382 1532 12242
rect 1596 11937 1624 12406
rect 1674 12200 1730 12209
rect 1674 12135 1730 12144
rect 1582 11928 1638 11937
rect 1582 11863 1638 11872
rect 1688 11694 1716 12135
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1674 11520 1730 11529
rect 1674 11455 1730 11464
rect 1688 10962 1716 11455
rect 1780 11286 1808 13246
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1688 10934 1808 10962
rect 1780 10742 1808 10934
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 9722 1624 10406
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1780 9178 1808 10678
rect 1872 10062 1900 12378
rect 1964 12374 1992 12786
rect 1952 12368 2004 12374
rect 1952 12310 2004 12316
rect 1964 11694 1992 12310
rect 2056 12306 2084 13348
rect 2148 12782 2176 16186
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2240 15910 2268 16118
rect 2332 16046 2360 17020
rect 2424 16250 2452 17070
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2240 13841 2268 14418
rect 2226 13832 2282 13841
rect 2226 13767 2282 13776
rect 2332 13716 2360 15982
rect 2240 13688 2360 13716
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2134 12608 2190 12617
rect 2134 12543 2190 12552
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2148 11694 2176 12543
rect 2240 12356 2268 13688
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12434 2360 13126
rect 2516 12986 2544 17274
rect 2608 16046 2636 17682
rect 2976 17610 3004 17818
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16658 2912 16934
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2608 13734 2636 15846
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13394 2636 13670
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2332 12406 2452 12434
rect 2240 12328 2360 12356
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11762 2268 12038
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2226 11656 2282 11665
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1228 6866 1256 8978
rect 1596 8430 1624 8978
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1308 8016 1360 8022
rect 1412 8004 1440 8230
rect 1360 7976 1440 8004
rect 1308 7958 1360 7964
rect 1412 7274 1440 7976
rect 1504 7954 1532 8298
rect 1492 7948 1544 7954
rect 1492 7890 1544 7896
rect 1504 7324 1532 7890
rect 1596 7546 1624 8366
rect 1688 7954 1716 8502
rect 1872 8090 1900 9318
rect 1964 8956 1992 11494
rect 2056 9518 2084 11630
rect 2148 11558 2176 11630
rect 2226 11591 2282 11600
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2044 8968 2096 8974
rect 1964 8928 2044 8956
rect 2044 8910 2096 8916
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 7478 1716 7890
rect 1872 7698 1900 8026
rect 1964 8022 1992 8774
rect 2056 8430 2084 8910
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 2056 7750 2084 8366
rect 1780 7670 1900 7698
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1584 7336 1636 7342
rect 1504 7296 1584 7324
rect 1584 7278 1636 7284
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 1596 7002 1624 7278
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1596 6254 1624 6938
rect 1688 6322 1716 7414
rect 1780 6458 1808 7670
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 1964 7342 1992 7482
rect 2148 7342 2176 11154
rect 2240 8362 2268 11591
rect 2332 11529 2360 12328
rect 2424 11778 2452 12406
rect 2504 11892 2556 11898
rect 2608 11880 2636 12718
rect 2700 11898 2728 15438
rect 2884 14482 2912 16458
rect 2976 14906 3004 17546
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 3068 16590 3096 17206
rect 3252 17134 3280 18634
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3330 17096 3386 17105
rect 3330 17031 3386 17040
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3160 16522 3188 16934
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3160 15337 3188 15506
rect 3146 15328 3202 15337
rect 3146 15263 3202 15272
rect 2976 14878 3096 14906
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 12918 2820 13330
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12986 2912 13126
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2884 12594 2912 12922
rect 2792 12566 2912 12594
rect 2556 11852 2636 11880
rect 2688 11892 2740 11898
rect 2504 11834 2556 11840
rect 2688 11834 2740 11840
rect 2424 11750 2544 11778
rect 2410 11656 2466 11665
rect 2410 11591 2466 11600
rect 2424 11558 2452 11591
rect 2412 11552 2464 11558
rect 2318 11520 2374 11529
rect 2412 11494 2464 11500
rect 2318 11455 2374 11464
rect 2332 11286 2360 11455
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2240 7886 2268 8298
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7478 2268 7822
rect 2228 7472 2280 7478
rect 2226 7440 2228 7449
rect 2280 7440 2282 7449
rect 2226 7375 2282 7384
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 2136 7336 2188 7342
rect 2136 7278 2188 7284
rect 1872 7002 1900 7278
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1320 5166 1348 5714
rect 1596 5710 1624 6190
rect 1688 5778 1716 6258
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1872 5273 1900 6734
rect 1964 6390 1992 7278
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1964 5846 1992 6326
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 1858 5264 1914 5273
rect 1858 5199 1914 5208
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4690 1348 5102
rect 2056 4758 2084 6802
rect 2148 5846 2176 7278
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 2240 5710 2268 6938
rect 2332 6798 2360 9998
rect 2424 8566 2452 11086
rect 2516 10033 2544 11750
rect 2792 11642 2820 12566
rect 2976 11880 3004 13874
rect 3068 13394 3096 14878
rect 3160 14550 3188 15263
rect 3252 14618 3280 15506
rect 3344 15450 3372 17031
rect 3436 15570 3464 18770
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 17105 3556 18566
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 4080 18290 4108 18838
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3804 17814 3832 18090
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3988 17746 4016 18158
rect 4080 17814 4108 18226
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 4264 17678 4292 18022
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4724 17882 4752 18158
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 4080 17202 4108 17614
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 3528 16114 3556 16186
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3344 15422 3464 15450
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3344 14958 3372 15302
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 3240 14476 3292 14482
rect 3292 14436 3372 14464
rect 3240 14418 3292 14424
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 3160 11898 3188 12854
rect 3148 11892 3200 11898
rect 2976 11852 3096 11880
rect 2962 11792 3018 11801
rect 2962 11727 2964 11736
rect 3016 11727 3018 11736
rect 2964 11698 3016 11704
rect 2700 11614 2820 11642
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 11354 2636 11494
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2502 10024 2558 10033
rect 2502 9959 2558 9968
rect 2608 9178 2636 10610
rect 2700 9625 2728 11614
rect 2778 11384 2834 11393
rect 2778 11319 2834 11328
rect 2792 10606 2820 11319
rect 2884 11082 2912 11630
rect 2964 11280 3016 11286
rect 2962 11248 2964 11257
rect 3016 11248 3018 11257
rect 2962 11183 3018 11192
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2686 9616 2742 9625
rect 2686 9551 2742 9560
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2516 9058 2544 9114
rect 2516 9030 2636 9058
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2424 8294 2452 8502
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2424 4826 2452 7890
rect 2502 5672 2558 5681
rect 2502 5607 2504 5616
rect 2556 5607 2558 5616
rect 2504 5578 2556 5584
rect 2608 5522 2636 9030
rect 2700 7002 2728 9454
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2792 6882 2820 10406
rect 2884 9110 2912 10746
rect 2976 9450 3004 11086
rect 3068 10810 3096 11852
rect 3148 11834 3200 11840
rect 3160 11626 3188 11834
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3252 11286 3280 14282
rect 3344 13870 3372 14436
rect 3436 14346 3464 15422
rect 3528 15094 3556 16050
rect 4080 15706 4108 17138
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 16726 4200 17070
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4264 16046 4292 17614
rect 4816 17377 4844 17682
rect 4342 17368 4398 17377
rect 4342 17303 4398 17312
rect 4802 17368 4858 17377
rect 4802 17303 4858 17312
rect 4356 17134 4384 17303
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4712 17060 4764 17066
rect 4712 17002 4764 17008
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4724 15638 4752 17002
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4816 16561 4844 16934
rect 4908 16590 4936 18770
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16794 5028 16934
rect 5092 16794 5120 17070
rect 5184 17066 5212 18226
rect 5276 18154 5304 18770
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5276 17338 5304 18090
rect 5368 18086 5396 18770
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5460 17898 5488 18906
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6274 18864 6330 18873
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 5920 18601 5948 18634
rect 5906 18592 5962 18601
rect 5906 18527 5962 18536
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5368 17870 5488 17898
rect 5632 17876 5684 17882
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5172 16720 5224 16726
rect 4986 16688 5042 16697
rect 5172 16662 5224 16668
rect 4986 16623 4988 16632
rect 5040 16623 5042 16632
rect 4988 16594 5040 16600
rect 4896 16584 4948 16590
rect 4802 16552 4858 16561
rect 4896 16526 4948 16532
rect 4802 16487 4858 16496
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 3516 15088 3568 15094
rect 4080 15042 4108 15506
rect 3516 15030 3568 15036
rect 3988 15014 4108 15042
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3424 14340 3476 14346
rect 3620 14328 3648 14894
rect 3988 14822 4016 15014
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3424 14282 3476 14288
rect 3528 14300 3648 14328
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3344 13297 3372 13806
rect 3330 13288 3386 13297
rect 3330 13223 3386 13232
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2884 8838 2912 9046
rect 2976 9042 3004 9386
rect 3068 9353 3096 9454
rect 3054 9344 3110 9353
rect 3054 9279 3110 9288
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 3068 8634 3096 8978
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2700 6854 2820 6882
rect 2700 6066 2728 6854
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6254 2820 6734
rect 2884 6458 2912 8298
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 6730 3004 8230
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3068 6322 3096 6598
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2700 6038 2820 6066
rect 2516 5494 2636 5522
rect 2516 5302 2544 5494
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2516 5137 2544 5238
rect 2792 5166 2820 6038
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2780 5160 2832 5166
rect 2502 5128 2558 5137
rect 2780 5102 2832 5108
rect 2502 5063 2558 5072
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2044 4752 2096 4758
rect 2044 4694 2096 4700
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 2056 2774 2084 4694
rect 2424 3466 2452 4762
rect 2792 4690 2820 5102
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3068 3670 3096 5714
rect 3160 4826 3188 11154
rect 3238 10704 3294 10713
rect 3238 10639 3294 10648
rect 3252 10606 3280 10639
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3252 9722 3280 10066
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3238 9616 3294 9625
rect 3238 9551 3294 9560
rect 3252 8294 3280 9551
rect 3344 8430 3372 13126
rect 3436 12442 3464 13806
rect 3528 13530 3556 14300
rect 3988 14278 4016 14758
rect 4080 14414 4108 14894
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3712 13462 3740 13806
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3988 13258 4016 13670
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3528 12306 3556 12582
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3436 11830 3464 12242
rect 3620 12186 3648 12242
rect 3528 12158 3648 12186
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3436 11132 3464 11562
rect 3528 11393 3556 12158
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3514 11384 3570 11393
rect 3514 11319 3570 11328
rect 3516 11144 3568 11150
rect 3436 11104 3516 11132
rect 3516 11086 3568 11092
rect 3620 10996 3648 11698
rect 3712 11694 3740 11834
rect 4080 11762 4108 14350
rect 4172 13190 4200 14418
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4160 12844 4212 12850
rect 4264 12832 4292 13738
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4212 12804 4292 12832
rect 4160 12786 4212 12792
rect 4172 12170 4200 12786
rect 4356 12628 4384 13194
rect 4448 12889 4476 13194
rect 4434 12880 4490 12889
rect 4434 12815 4490 12824
rect 4540 12782 4568 13466
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12782 4660 13330
rect 4724 12889 4752 13806
rect 4816 13569 4844 16390
rect 5000 16046 5028 16390
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4802 13560 4858 13569
rect 4802 13495 4858 13504
rect 4908 13240 4936 14894
rect 5000 13394 5028 15982
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5184 15450 5212 16662
rect 5276 16250 5304 16934
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5092 15314 5120 15438
rect 5184 15422 5304 15450
rect 5092 15286 5212 15314
rect 5078 15192 5134 15201
rect 5078 15127 5134 15136
rect 5092 15026 5120 15127
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5184 14822 5212 15286
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5078 14104 5134 14113
rect 5078 14039 5134 14048
rect 5092 13841 5120 14039
rect 5172 13864 5224 13870
rect 5078 13832 5134 13841
rect 5172 13806 5224 13812
rect 5078 13767 5134 13776
rect 5184 13530 5212 13806
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 4908 13212 5028 13240
rect 4710 12880 4766 12889
rect 4710 12815 4766 12824
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4264 12600 4384 12628
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3712 11218 3740 11494
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3712 11014 3740 11154
rect 3804 11014 3832 11698
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3528 10968 3648 10996
rect 3700 11008 3752 11014
rect 3528 10656 3556 10968
rect 3700 10950 3752 10956
rect 3792 11008 3844 11014
rect 3896 10996 3924 11630
rect 4068 11620 4120 11626
rect 4120 11580 4200 11608
rect 4068 11562 4120 11568
rect 3976 11552 4028 11558
rect 4172 11529 4200 11580
rect 3976 11494 4028 11500
rect 4158 11520 4214 11529
rect 3988 11354 4016 11494
rect 4158 11455 4214 11464
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3896 10968 4108 10996
rect 3792 10950 3844 10956
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 4080 10810 4108 10968
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3436 10628 3648 10656
rect 3436 10538 3464 10628
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3344 6866 3372 8366
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3436 6662 3464 9930
rect 3528 9081 3556 10474
rect 3620 9926 3648 10628
rect 3700 10600 3752 10606
rect 3698 10568 3700 10577
rect 3752 10568 3754 10577
rect 3698 10503 3754 10512
rect 3804 10418 3832 10746
rect 4172 10690 4200 11455
rect 4264 11218 4292 12600
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 4816 12458 4844 12718
rect 4816 12430 4936 12458
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4802 12336 4858 12345
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11626 4476 12038
rect 4540 11694 4568 12106
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4540 11540 4568 11630
rect 4724 11608 4752 12310
rect 4802 12271 4858 12280
rect 4816 12170 4844 12271
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4908 12102 4936 12430
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4724 11580 4844 11608
rect 4540 11512 4752 11540
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4540 11014 4568 11222
rect 4632 11121 4660 11290
rect 4724 11218 4752 11512
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4618 11112 4674 11121
rect 4618 11047 4674 11056
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4710 10976 4766 10985
rect 4342 10840 4398 10849
rect 4252 10804 4304 10810
rect 4342 10775 4398 10784
rect 4252 10746 4304 10752
rect 4080 10662 4200 10690
rect 3804 10390 3924 10418
rect 3790 10296 3846 10305
rect 3790 10231 3792 10240
rect 3844 10231 3846 10240
rect 3792 10202 3844 10208
rect 3896 10130 3924 10390
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3712 9382 3740 9454
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3514 9072 3570 9081
rect 3514 9007 3570 9016
rect 3712 8974 3740 9318
rect 3804 9178 3832 9454
rect 4080 9178 4108 10662
rect 4264 10520 4292 10746
rect 4356 10606 4384 10775
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4172 10492 4292 10520
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 4080 8809 4108 8978
rect 4066 8800 4122 8809
rect 3662 8732 3970 8741
rect 4066 8735 4122 8744
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 3976 8628 4028 8634
rect 4172 8616 4200 10492
rect 4448 10452 4476 10950
rect 4710 10911 4766 10920
rect 4264 10424 4476 10452
rect 4264 10248 4292 10424
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 4264 10220 4476 10248
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4252 10056 4304 10062
rect 4250 10024 4252 10033
rect 4304 10024 4306 10033
rect 4250 9959 4306 9968
rect 4264 9722 4292 9959
rect 4356 9897 4384 10066
rect 4342 9888 4398 9897
rect 4342 9823 4398 9832
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4448 9382 4476 10220
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4540 9654 4568 10066
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4724 9382 4752 10911
rect 4816 10810 4844 11580
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4816 10606 4844 10746
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4816 9654 4844 10134
rect 4908 9994 4936 10406
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4712 9376 4764 9382
rect 4816 9353 4844 9454
rect 4712 9318 4764 9324
rect 4802 9344 4858 9353
rect 4322 9276 4630 9285
rect 4802 9279 4858 9288
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 8968 4488 8974
rect 4540 8945 4568 8978
rect 4436 8910 4488 8916
rect 4526 8936 4582 8945
rect 4342 8664 4398 8673
rect 4172 8588 4292 8616
rect 4342 8599 4344 8608
rect 3976 8570 4028 8576
rect 3516 8424 3568 8430
rect 3608 8424 3660 8430
rect 3516 8366 3568 8372
rect 3606 8392 3608 8401
rect 3700 8424 3752 8430
rect 3660 8392 3662 8401
rect 3528 7342 3556 8366
rect 3700 8366 3752 8372
rect 3606 8327 3662 8336
rect 3712 8294 3740 8366
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3988 7750 4016 8570
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3620 6866 3648 7210
rect 3712 6866 3740 7482
rect 3976 7336 4028 7342
rect 3974 7304 3976 7313
rect 4028 7304 4030 7313
rect 3974 7239 4030 7248
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3988 6769 4016 7142
rect 4080 6866 4108 7890
rect 4172 7818 4200 8434
rect 4264 8430 4292 8588
rect 4396 8599 4398 8608
rect 4344 8570 4396 8576
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4448 8294 4476 8910
rect 4526 8871 4582 8880
rect 4526 8800 4582 8809
rect 4526 8735 4582 8744
rect 4540 8294 4568 8735
rect 4618 8528 4674 8537
rect 4724 8514 4752 9114
rect 4908 9042 4936 9658
rect 4896 9036 4948 9042
rect 4816 8996 4896 9024
rect 4816 8634 4844 8996
rect 4896 8978 4948 8984
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4724 8486 4844 8514
rect 4618 8463 4674 8472
rect 4632 8430 4660 8463
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4436 8288 4488 8294
rect 4540 8266 4752 8294
rect 4436 8230 4488 8236
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4172 6866 4200 7754
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7546 4292 7686
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3974 6760 4030 6769
rect 3620 6730 3974 6746
rect 3608 6724 3974 6730
rect 3660 6718 3974 6724
rect 4264 6746 4292 7346
rect 4356 7342 4384 7958
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4632 7750 4660 7890
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4724 7426 4752 8266
rect 4816 7546 4844 8486
rect 4908 8430 4936 8774
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4894 7848 4950 7857
rect 4894 7783 4896 7792
rect 4948 7783 4950 7792
rect 4896 7754 4948 7760
rect 4894 7576 4950 7585
rect 4804 7540 4856 7546
rect 5000 7546 5028 13212
rect 5078 13016 5134 13025
rect 5184 12986 5212 13330
rect 5078 12951 5134 12960
rect 5172 12980 5224 12986
rect 5092 12782 5120 12951
rect 5172 12922 5224 12928
rect 5276 12782 5304 15422
rect 5368 14550 5396 17870
rect 5632 17818 5684 17824
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5460 15706 5488 17206
rect 5644 17134 5672 17818
rect 5828 17746 5856 18362
rect 6012 17746 6040 18702
rect 6104 18057 6132 18838
rect 6184 18828 6236 18834
rect 6274 18799 6330 18808
rect 6184 18770 6236 18776
rect 6196 18465 6224 18770
rect 6182 18456 6238 18465
rect 6182 18391 6238 18400
rect 6288 18290 6316 18799
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6090 18048 6146 18057
rect 6090 17983 6146 17992
rect 5816 17740 5868 17746
rect 5736 17700 5816 17728
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5552 16590 5580 17002
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5552 15502 5580 15846
rect 5644 15570 5672 15914
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5540 15496 5592 15502
rect 5538 15464 5540 15473
rect 5592 15464 5594 15473
rect 5538 15399 5594 15408
rect 5736 15314 5764 17700
rect 5816 17682 5868 17688
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 5920 17270 5948 17478
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5814 17096 5870 17105
rect 5814 17031 5870 17040
rect 5644 15286 5764 15314
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5460 14482 5488 15098
rect 5540 14816 5592 14822
rect 5644 14804 5672 15286
rect 5828 15026 5856 17031
rect 6012 16980 6040 17478
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6104 17134 6132 17274
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 5920 16952 6040 16980
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5814 14920 5870 14929
rect 5592 14776 5672 14804
rect 5540 14758 5592 14764
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5368 14074 5396 14350
rect 5552 14346 5580 14758
rect 5736 14482 5764 14894
rect 5814 14855 5870 14864
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5724 14272 5776 14278
rect 5538 14240 5594 14249
rect 5724 14214 5776 14220
rect 5538 14175 5594 14184
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5460 13870 5488 14010
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13734 5488 13806
rect 5552 13802 5580 14175
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5354 13152 5410 13161
rect 5354 13087 5410 13096
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5184 12442 5212 12582
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5276 12306 5304 12582
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5092 9042 5120 12106
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 11898 5212 12038
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5184 11529 5212 11562
rect 5170 11520 5226 11529
rect 5170 11455 5226 11464
rect 5184 11354 5212 11455
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5276 10742 5304 11562
rect 5368 11336 5396 13087
rect 5552 12889 5580 13398
rect 5538 12880 5594 12889
rect 5538 12815 5594 12824
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 12442 5488 12718
rect 5448 12436 5500 12442
rect 5644 12434 5672 13874
rect 5448 12378 5500 12384
rect 5552 12406 5672 12434
rect 5368 11308 5488 11336
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5078 8936 5134 8945
rect 5078 8871 5134 8880
rect 5092 8838 5120 8871
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5092 8430 5120 8570
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5184 8362 5212 10610
rect 5276 10130 5304 10678
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5276 9042 5304 9386
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5078 8256 5134 8265
rect 5078 8191 5134 8200
rect 5092 7721 5120 8191
rect 5184 7954 5212 8298
rect 5276 7954 5304 8570
rect 5368 8022 5396 11154
rect 5460 10674 5488 11308
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5552 10554 5580 12406
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5644 12209 5672 12310
rect 5630 12200 5686 12209
rect 5630 12135 5686 12144
rect 5736 10985 5764 14214
rect 5828 13734 5856 14855
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5828 11830 5856 13670
rect 5920 13462 5948 16952
rect 6196 16794 6224 18158
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6288 17542 6316 18022
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6380 17105 6408 19110
rect 6472 18766 6500 19230
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6564 17678 6592 22063
rect 11980 22024 12032 22030
rect 11886 21992 11942 22001
rect 26884 22024 26936 22030
rect 11980 21966 12032 21972
rect 12254 21992 12310 22001
rect 11886 21927 11942 21936
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 9586 21856 9642 21865
rect 6734 21720 6790 21729
rect 6734 21655 6736 21664
rect 6788 21655 6790 21664
rect 7286 21720 7342 21729
rect 7286 21655 7288 21664
rect 6736 21626 6788 21632
rect 7340 21655 7342 21664
rect 7838 21720 7894 21729
rect 7838 21655 7840 21664
rect 7288 21626 7340 21632
rect 7892 21655 7894 21664
rect 8390 21720 8446 21729
rect 8390 21655 8392 21664
rect 7840 21626 7892 21632
rect 8444 21655 8446 21664
rect 8392 21626 8444 21632
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 7852 21010 7880 21286
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7208 20058 7236 20878
rect 7668 20466 7696 20946
rect 8484 20528 8536 20534
rect 8484 20470 8536 20476
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7562 20360 7618 20369
rect 7562 20295 7618 20304
rect 7286 20088 7342 20097
rect 7196 20052 7248 20058
rect 7286 20023 7342 20032
rect 7196 19994 7248 20000
rect 7208 19922 7236 19994
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18698 6868 19110
rect 7010 18864 7066 18873
rect 7010 18799 7012 18808
rect 7064 18799 7066 18808
rect 7012 18770 7064 18776
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6644 18624 6696 18630
rect 6642 18592 6644 18601
rect 6696 18592 6698 18601
rect 6642 18527 6698 18536
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6656 17882 6684 18158
rect 6734 18048 6790 18057
rect 6734 17983 6790 17992
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6366 17096 6422 17105
rect 6472 17066 6500 17478
rect 6366 17031 6422 17040
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6012 16046 6040 16594
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6012 15910 6040 15982
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6012 14550 6040 15438
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6104 14958 6132 15098
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6012 14074 6040 14486
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6012 13870 6040 14010
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 6012 13462 6040 13806
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5920 13190 5948 13262
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 5816 11008 5868 11014
rect 5722 10976 5778 10985
rect 5816 10950 5868 10956
rect 5722 10911 5778 10920
rect 5460 10526 5580 10554
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5460 9722 5488 10526
rect 5540 10464 5592 10470
rect 5538 10432 5540 10441
rect 5592 10432 5594 10441
rect 5538 10367 5594 10376
rect 5644 10062 5672 10542
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5538 9752 5594 9761
rect 5448 9716 5500 9722
rect 5736 9722 5764 10542
rect 5538 9687 5594 9696
rect 5724 9716 5776 9722
rect 5448 9658 5500 9664
rect 5446 9616 5502 9625
rect 5446 9551 5448 9560
rect 5500 9551 5502 9560
rect 5448 9522 5500 9528
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5460 8634 5488 9386
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5460 7954 5488 8570
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5078 7712 5134 7721
rect 5078 7647 5134 7656
rect 4894 7511 4896 7520
rect 4804 7482 4856 7488
rect 4948 7511 4950 7520
rect 4988 7540 5040 7546
rect 4896 7482 4948 7488
rect 4988 7482 5040 7488
rect 4724 7398 5028 7426
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4172 6730 4292 6746
rect 3974 6695 4030 6704
rect 4160 6724 4292 6730
rect 3608 6666 3660 6672
rect 4212 6718 4292 6724
rect 4160 6666 4212 6672
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 3332 6248 3384 6254
rect 3608 6248 3660 6254
rect 3332 6190 3384 6196
rect 3528 6196 3608 6202
rect 3528 6190 3660 6196
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3252 3602 3280 5714
rect 3344 5658 3372 6190
rect 3528 6174 3648 6190
rect 3976 6180 4028 6186
rect 3528 5846 3556 6174
rect 4080 6168 4108 6598
rect 4632 6254 4660 6938
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4028 6140 4108 6168
rect 3976 6122 4028 6128
rect 4080 5846 4108 6140
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4724 5914 4752 7278
rect 4816 6866 4844 7278
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4802 6352 4858 6361
rect 4802 6287 4858 6296
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3424 5704 3476 5710
rect 3344 5652 3424 5658
rect 3344 5646 3476 5652
rect 3344 5630 3464 5646
rect 3344 3602 3372 5630
rect 3528 5352 3556 5782
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 3528 5324 3648 5352
rect 3620 5098 3648 5324
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3436 4010 3464 4626
rect 3528 4078 3556 4626
rect 3620 4622 3648 5034
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3436 3738 3464 3946
rect 3620 3942 3648 4111
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 3712 3398 3740 4218
rect 4080 3602 4108 5782
rect 4816 5778 4844 6287
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4250 5536 4306 5545
rect 4250 5471 4306 5480
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4172 4690 4200 5102
rect 4264 5030 4292 5471
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 4826 4292 4966
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4078 4200 4626
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4282 4292 4558
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4908 3738 4936 7278
rect 5000 6186 5028 7398
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 5000 4826 5028 5238
rect 5092 5166 5120 7647
rect 5184 6934 5212 7890
rect 5276 7002 5304 7890
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5368 7177 5396 7278
rect 5552 7206 5580 9687
rect 5724 9658 5776 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9110 5672 9454
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5644 8362 5672 9046
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5540 7200 5592 7206
rect 5354 7168 5410 7177
rect 5540 7142 5592 7148
rect 5354 7103 5410 7112
rect 5264 6996 5316 7002
rect 5644 6984 5672 8298
rect 5264 6938 5316 6944
rect 5368 6956 5672 6984
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5368 6866 5396 6956
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6322 5396 6802
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5262 6080 5318 6089
rect 5184 5778 5212 6054
rect 5262 6015 5318 6024
rect 5276 5778 5304 6015
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5092 4010 5120 4626
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4078 5212 4422
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5736 3670 5764 9522
rect 5828 9450 5856 10950
rect 5920 10656 5948 12786
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6012 12345 6040 12718
rect 5998 12336 6054 12345
rect 5998 12271 6054 12280
rect 6012 12238 6040 12271
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6012 10810 6040 11766
rect 6104 11354 6132 14350
rect 6196 13841 6224 14350
rect 6288 14074 6316 16594
rect 6380 16250 6408 16594
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6182 13832 6238 13841
rect 6182 13767 6238 13776
rect 6182 13560 6238 13569
rect 6182 13495 6238 13504
rect 6196 12714 6224 13495
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12850 6316 13126
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6288 12753 6316 12786
rect 6274 12744 6330 12753
rect 6184 12708 6236 12714
rect 6274 12679 6330 12688
rect 6184 12650 6236 12656
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6196 12073 6224 12378
rect 6182 12064 6238 12073
rect 6182 11999 6238 12008
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6104 10810 6132 10950
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5920 10628 6040 10656
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5920 10266 5948 10474
rect 6012 10441 6040 10628
rect 5998 10432 6054 10441
rect 5998 10367 6054 10376
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5828 9042 5856 9386
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5828 6798 5856 8502
rect 5920 8265 5948 10202
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6012 9178 6040 9454
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5998 8936 6054 8945
rect 5998 8871 6054 8880
rect 5906 8256 5962 8265
rect 5906 8191 5962 8200
rect 6012 7936 6040 8871
rect 6104 8498 6132 10746
rect 6196 10470 6224 11999
rect 6288 11642 6316 12679
rect 6380 12617 6408 15098
rect 6472 14362 6500 17002
rect 6564 16658 6592 17614
rect 6656 17338 6684 17818
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 14618 6592 15302
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6472 14334 6592 14362
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6472 13870 6500 14214
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6366 12608 6422 12617
rect 6366 12543 6422 12552
rect 6472 12102 6500 13806
rect 6564 13190 6592 14334
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6564 12782 6592 12922
rect 6552 12776 6604 12782
rect 6550 12744 6552 12753
rect 6604 12744 6606 12753
rect 6550 12679 6606 12688
rect 6550 12608 6606 12617
rect 6550 12543 6606 12552
rect 6564 12170 6592 12543
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6288 11614 6408 11642
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 10606 6316 11494
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6274 10432 6330 10441
rect 6274 10367 6330 10376
rect 6182 10296 6238 10305
rect 6182 10231 6238 10240
rect 6196 10130 6224 10231
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6012 7908 6132 7936
rect 5998 7848 6054 7857
rect 5998 7783 6054 7792
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5814 6352 5870 6361
rect 5814 6287 5870 6296
rect 5828 6118 5856 6287
rect 6012 6186 6040 7783
rect 6104 6866 6132 7908
rect 6196 7177 6224 10066
rect 6288 8945 6316 10367
rect 6380 10044 6408 11614
rect 6472 10198 6500 12038
rect 6656 11898 6684 16730
rect 6748 13138 6776 17983
rect 6840 17746 6868 18294
rect 7024 18154 7052 18770
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7116 18086 7144 18702
rect 7300 18272 7328 20023
rect 7576 19961 7604 20295
rect 7562 19952 7618 19961
rect 7562 19887 7618 19896
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7484 19514 7512 19790
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 8496 19310 8524 20470
rect 9048 20398 9076 21286
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 8864 19700 8892 20334
rect 8956 19854 8984 20334
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8944 19712 8996 19718
rect 8864 19672 8944 19700
rect 8944 19654 8996 19660
rect 8956 19514 8984 19654
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 8390 18864 8446 18873
rect 8390 18799 8392 18808
rect 8444 18799 8446 18808
rect 8576 18828 8628 18834
rect 8392 18770 8444 18776
rect 8576 18770 8628 18776
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7208 18244 7328 18272
rect 7392 18272 7420 18702
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 8298 18592 8354 18601
rect 7484 18426 7512 18566
rect 8298 18527 8354 18536
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7392 18244 7512 18272
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 6920 17672 6972 17678
rect 6918 17640 6920 17649
rect 7012 17672 7064 17678
rect 6972 17640 6974 17649
rect 7012 17614 7064 17620
rect 6918 17575 6974 17584
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6840 16454 6868 17274
rect 6932 17241 6960 17575
rect 7024 17338 7052 17614
rect 7116 17377 7144 17682
rect 7102 17368 7158 17377
rect 7012 17332 7064 17338
rect 7102 17303 7158 17312
rect 7012 17274 7064 17280
rect 6918 17232 6974 17241
rect 6918 17167 6974 17176
rect 7208 17134 7236 18244
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7300 17338 7328 18090
rect 7392 17746 7420 18090
rect 7484 17882 7512 18244
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7576 17921 7604 18090
rect 7562 17912 7618 17921
rect 7472 17876 7524 17882
rect 7562 17847 7618 17856
rect 7930 17912 7986 17921
rect 7930 17847 7986 17856
rect 7472 17818 7524 17824
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7208 16726 7236 17070
rect 7300 16998 7328 17070
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6932 16114 6960 16526
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6840 14958 6868 15506
rect 6932 15026 6960 16050
rect 7024 15638 7052 16050
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14952 6880 14958
rect 7012 14952 7064 14958
rect 6828 14894 6880 14900
rect 6918 14920 6974 14929
rect 7012 14894 7064 14900
rect 6918 14855 6974 14864
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14657 6868 14758
rect 6826 14648 6882 14657
rect 6826 14583 6882 14592
rect 6932 14482 6960 14855
rect 7024 14793 7052 14894
rect 7010 14784 7066 14793
rect 7010 14719 7066 14728
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6840 13852 6868 14282
rect 6932 14006 6960 14282
rect 7024 14074 7052 14554
rect 7116 14482 7144 16186
rect 7300 16153 7328 16934
rect 7286 16144 7342 16153
rect 7286 16079 7342 16088
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6920 14000 6972 14006
rect 7116 13954 7144 14418
rect 6920 13942 6972 13948
rect 7024 13926 7144 13954
rect 6840 13824 6960 13852
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13394 6868 13670
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6748 13110 6868 13138
rect 6840 12986 6868 13110
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6748 12753 6776 12922
rect 6828 12776 6880 12782
rect 6734 12744 6790 12753
rect 6828 12718 6880 12724
rect 6734 12679 6790 12688
rect 6840 12442 6868 12718
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6748 11218 6776 11834
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6642 11112 6698 11121
rect 6642 11047 6698 11056
rect 6736 11076 6788 11082
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10470 6592 10950
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6380 10016 6592 10044
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6380 9110 6408 9386
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6472 9042 6500 9658
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6368 8968 6420 8974
rect 6274 8936 6330 8945
rect 6368 8910 6420 8916
rect 6274 8871 6330 8880
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6182 7168 6238 7177
rect 6182 7103 6238 7112
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5828 4826 5856 5782
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6012 4690 6040 5102
rect 6104 4690 6132 6802
rect 6288 6662 6316 8774
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6288 5914 6316 6122
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5370 6316 5714
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6012 4214 6040 4626
rect 6196 4622 6224 5102
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4622 6316 4966
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 6196 4146 6224 4558
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6288 3942 6316 4558
rect 6380 4146 6408 8910
rect 6472 8634 6500 8978
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6564 8430 6592 10016
rect 6656 9217 6684 11047
rect 6736 11018 6788 11024
rect 6748 10606 6776 11018
rect 6840 11014 6868 11494
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6932 10470 6960 13824
rect 7024 13462 7052 13926
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12918 7052 13262
rect 7116 13190 7144 13806
rect 7208 13546 7236 15982
rect 7286 15056 7342 15065
rect 7286 14991 7288 15000
rect 7340 14991 7342 15000
rect 7288 14962 7340 14968
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7300 14618 7328 14826
rect 7392 14618 7420 17478
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16998 7512 17070
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7484 16522 7512 16934
rect 7668 16833 7696 17614
rect 7654 16824 7710 16833
rect 7654 16759 7710 16768
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15706 7512 15846
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7484 15570 7512 15642
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7576 15502 7604 16526
rect 7668 16289 7696 16759
rect 7654 16280 7710 16289
rect 7654 16215 7710 16224
rect 7852 15960 7880 17682
rect 7944 17610 7972 17847
rect 8036 17678 8064 18362
rect 8312 18154 8340 18527
rect 8484 18216 8536 18222
rect 8588 18193 8616 18770
rect 8956 18630 8984 18770
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8484 18158 8536 18164
rect 8574 18184 8630 18193
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8392 18080 8444 18086
rect 8390 18048 8392 18057
rect 8444 18048 8446 18057
rect 8390 17983 8446 17992
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 8128 17542 8156 17750
rect 8220 17649 8248 17818
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8206 17640 8262 17649
rect 8206 17575 8262 17584
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8404 17338 8432 17682
rect 8496 17377 8524 18158
rect 8574 18119 8630 18128
rect 8482 17368 8538 17377
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8392 17332 8444 17338
rect 8482 17303 8538 17312
rect 8392 17274 8444 17280
rect 8208 16720 8260 16726
rect 8206 16688 8208 16697
rect 8260 16688 8262 16697
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8116 16652 8168 16658
rect 8206 16623 8262 16632
rect 8116 16594 8168 16600
rect 8036 16046 8064 16594
rect 8128 16114 8156 16594
rect 8312 16522 8340 17274
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 7932 15972 7984 15978
rect 7852 15932 7932 15960
rect 7932 15914 7984 15920
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15570 7696 15846
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7564 15496 7616 15502
rect 7748 15496 7800 15502
rect 7564 15438 7616 15444
rect 7668 15444 7748 15450
rect 7668 15438 7800 15444
rect 7470 15328 7526 15337
rect 7470 15263 7526 15272
rect 7484 14929 7512 15263
rect 7576 15042 7604 15438
rect 7668 15422 7788 15438
rect 7668 15162 7696 15422
rect 7944 15348 7972 15914
rect 8220 15620 8248 15982
rect 8312 15745 8340 15982
rect 8298 15736 8354 15745
rect 8298 15671 8354 15680
rect 8220 15592 8340 15620
rect 8404 15609 8432 17070
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8496 16658 8524 17002
rect 8680 16794 8708 18362
rect 8852 18216 8904 18222
rect 8758 18184 8814 18193
rect 8852 18158 8904 18164
rect 8758 18119 8814 18128
rect 8772 17338 8800 18119
rect 8864 18057 8892 18158
rect 8850 18048 8906 18057
rect 8850 17983 8906 17992
rect 8850 17912 8906 17921
rect 8850 17847 8906 17856
rect 8864 17746 8892 17847
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8772 17134 8800 17274
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8956 16833 8984 17614
rect 8942 16824 8998 16833
rect 8668 16788 8720 16794
rect 8942 16759 8998 16768
rect 8668 16730 8720 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16289 8524 16594
rect 8482 16280 8538 16289
rect 8482 16215 8538 16224
rect 8496 15638 8524 16215
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8484 15632 8536 15638
rect 7760 15320 7972 15348
rect 8024 15360 8076 15366
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7760 15042 7788 15320
rect 8024 15302 8076 15308
rect 8036 15201 8064 15302
rect 8022 15192 8078 15201
rect 8022 15127 8078 15136
rect 8036 15094 8064 15127
rect 8024 15088 8076 15094
rect 7576 15014 7696 15042
rect 7760 15014 7880 15042
rect 8024 15030 8076 15036
rect 7564 14952 7616 14958
rect 7470 14920 7526 14929
rect 7668 14940 7696 15014
rect 7668 14912 7788 14940
rect 7564 14894 7616 14900
rect 7470 14855 7526 14864
rect 7470 14784 7526 14793
rect 7470 14719 7526 14728
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7484 14482 7512 14719
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7300 13716 7328 14418
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7392 13870 7420 14282
rect 7472 14272 7524 14278
rect 7470 14240 7472 14249
rect 7524 14240 7526 14249
rect 7470 14175 7526 14184
rect 7380 13864 7432 13870
rect 7576 13841 7604 14894
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7380 13806 7432 13812
rect 7562 13832 7618 13841
rect 7562 13767 7618 13776
rect 7472 13728 7524 13734
rect 7300 13688 7420 13716
rect 7208 13518 7328 13546
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 7024 11898 7052 12854
rect 7116 12374 7144 13126
rect 7208 12986 7236 13398
rect 7300 13326 7328 13518
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 7208 12306 7236 12922
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7194 12200 7250 12209
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11558 7144 12174
rect 7194 12135 7250 12144
rect 7208 11694 7236 12135
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7010 11248 7066 11257
rect 7010 11183 7066 11192
rect 7196 11212 7248 11218
rect 7024 10606 7052 11183
rect 7196 11154 7248 11160
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 7024 10266 7052 10542
rect 7116 10266 7144 11086
rect 7208 10810 7236 11154
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6642 9208 6698 9217
rect 6642 9143 6698 9152
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6472 5930 6500 8366
rect 6656 7750 6684 9143
rect 6748 9110 6776 10066
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 9586 6868 9862
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6932 9518 6960 10134
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7208 9926 7236 10066
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 6920 9512 6972 9518
rect 7104 9512 7156 9518
rect 6920 9454 6972 9460
rect 7024 9472 7104 9500
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 9178 6868 9318
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6748 8566 6776 9046
rect 7024 8906 7052 9472
rect 7104 9454 7156 9460
rect 7208 9382 7236 9862
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6918 8392 6974 8401
rect 6918 8327 6974 8336
rect 6932 7993 6960 8327
rect 6918 7984 6974 7993
rect 6918 7919 6974 7928
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6826 7440 6882 7449
rect 6826 7375 6882 7384
rect 6840 7342 6868 7375
rect 7024 7342 7052 8842
rect 7208 7410 7236 9318
rect 7300 7546 7328 13262
rect 7392 13258 7420 13688
rect 7472 13670 7524 13676
rect 7562 13696 7618 13705
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7484 12986 7512 13670
rect 7562 13631 7618 13640
rect 7576 13530 7604 13631
rect 7668 13530 7696 14758
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7576 12442 7604 13330
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 7668 12288 7696 13194
rect 7760 12986 7788 14912
rect 7852 13802 7880 15014
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 7930 14648 7986 14657
rect 7930 14583 7986 14592
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7944 13512 7972 14583
rect 8128 14550 8156 14758
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8116 14408 8168 14414
rect 8022 14376 8078 14385
rect 8116 14350 8168 14356
rect 8022 14311 8078 14320
rect 7852 13484 7972 13512
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7852 12866 7880 13484
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 13190 7972 13330
rect 8036 13190 8064 14311
rect 8128 13870 8156 14350
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8220 13569 8248 14894
rect 8312 14249 8340 15592
rect 8390 15600 8446 15609
rect 8484 15574 8536 15580
rect 8390 15535 8446 15544
rect 8588 15094 8616 15914
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8680 14906 8708 16730
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8956 15881 8984 15982
rect 9048 15910 9076 19178
rect 9140 17814 9168 21830
rect 9586 21791 9642 21800
rect 9494 21720 9550 21729
rect 9600 21690 9628 21791
rect 11436 21788 11744 21797
rect 11436 21786 11442 21788
rect 11498 21786 11522 21788
rect 11578 21786 11602 21788
rect 11658 21786 11682 21788
rect 11738 21786 11744 21788
rect 11498 21734 11500 21786
rect 11680 21734 11682 21786
rect 11436 21732 11442 21734
rect 11498 21732 11522 21734
rect 11578 21732 11602 21734
rect 11658 21732 11682 21734
rect 11738 21732 11744 21734
rect 10046 21720 10102 21729
rect 9494 21655 9496 21664
rect 9548 21655 9550 21664
rect 9588 21684 9640 21690
rect 9496 21626 9548 21632
rect 10046 21655 10048 21664
rect 9588 21626 9640 21632
rect 10100 21655 10102 21664
rect 10598 21720 10654 21729
rect 10598 21655 10600 21664
rect 10048 21626 10100 21632
rect 10652 21655 10654 21664
rect 11150 21720 11206 21729
rect 11436 21723 11744 21732
rect 11900 21690 11928 21927
rect 11150 21655 11152 21664
rect 10600 21626 10652 21632
rect 11204 21655 11206 21664
rect 11428 21684 11480 21690
rect 11152 21626 11204 21632
rect 11428 21626 11480 21632
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9588 21072 9640 21078
rect 9588 21014 9640 21020
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 9232 19990 9260 20470
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9220 19984 9272 19990
rect 9220 19926 9272 19932
rect 9324 19378 9352 20198
rect 9600 19990 9628 21014
rect 9968 20942 9996 21422
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10612 21146 10640 21286
rect 10600 21140 10652 21146
rect 10520 21100 10600 21128
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 10414 20904 10470 20913
rect 9968 20398 9996 20878
rect 10414 20839 10470 20848
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9588 19984 9640 19990
rect 9588 19926 9640 19932
rect 9496 19712 9548 19718
rect 9600 19700 9628 19926
rect 10138 19816 10194 19825
rect 10138 19751 10194 19760
rect 9548 19672 9628 19700
rect 9496 19654 9548 19660
rect 9678 19408 9734 19417
rect 9312 19372 9364 19378
rect 9678 19343 9734 19352
rect 9312 19314 9364 19320
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18834 9260 19110
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9218 18592 9274 18601
rect 9218 18527 9274 18536
rect 9232 18086 9260 18527
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9220 17876 9272 17882
rect 9324 17864 9352 18770
rect 9494 18456 9550 18465
rect 9494 18391 9550 18400
rect 9272 17836 9352 17864
rect 9220 17818 9272 17824
rect 9128 17808 9180 17814
rect 9128 17750 9180 17756
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9218 17640 9274 17649
rect 9218 17575 9220 17584
rect 9272 17575 9274 17584
rect 9312 17604 9364 17610
rect 9220 17546 9272 17552
rect 9312 17546 9364 17552
rect 9324 17377 9352 17546
rect 9416 17542 9444 17750
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9310 17368 9366 17377
rect 9310 17303 9366 17312
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9036 15904 9088 15910
rect 8942 15872 8998 15881
rect 9036 15846 9088 15852
rect 8942 15807 8998 15816
rect 9048 15638 9076 15846
rect 9036 15632 9088 15638
rect 9036 15574 9088 15580
rect 8944 15496 8996 15502
rect 9220 15496 9272 15502
rect 8996 15456 9168 15484
rect 8944 15438 8996 15444
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 15026 8892 15302
rect 8942 15056 8998 15065
rect 8852 15020 8904 15026
rect 8942 14991 8998 15000
rect 8852 14962 8904 14968
rect 8496 14634 8524 14894
rect 8588 14804 8616 14894
rect 8680 14878 8800 14906
rect 8588 14776 8708 14804
rect 8496 14606 8616 14634
rect 8390 14512 8446 14521
rect 8588 14482 8616 14606
rect 8390 14447 8446 14456
rect 8576 14476 8628 14482
rect 8404 14278 8432 14447
rect 8576 14418 8628 14424
rect 8574 14376 8630 14385
rect 8574 14311 8630 14320
rect 8392 14272 8444 14278
rect 8298 14240 8354 14249
rect 8392 14214 8444 14220
rect 8298 14175 8354 14184
rect 8404 14074 8432 14214
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8588 13870 8616 14311
rect 8680 14278 8708 14776
rect 8772 14657 8800 14878
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8758 14648 8814 14657
rect 8758 14583 8760 14592
rect 8812 14583 8814 14592
rect 8760 14554 8812 14560
rect 8758 14512 8814 14521
rect 8758 14447 8760 14456
rect 8812 14447 8814 14456
rect 8760 14418 8812 14424
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8206 13560 8262 13569
rect 8206 13495 8262 13504
rect 7932 13184 7984 13190
rect 8024 13184 8076 13190
rect 7932 13126 7984 13132
rect 8022 13152 8024 13161
rect 8076 13152 8078 13161
rect 8022 13087 8078 13096
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 7576 12260 7696 12288
rect 7760 12838 7880 12866
rect 7576 12220 7604 12260
rect 7760 12220 7788 12838
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7944 12617 7972 12718
rect 7930 12608 7986 12617
rect 7930 12543 7986 12552
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7484 12192 7604 12220
rect 7668 12192 7788 12220
rect 7484 10606 7512 12192
rect 7668 12050 7696 12192
rect 7576 12022 7696 12050
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7840 12096 7892 12102
rect 7944 12073 7972 12378
rect 7840 12038 7892 12044
rect 7930 12064 7986 12073
rect 7576 11694 7604 12022
rect 7656 11892 7708 11898
rect 7760 11880 7788 12038
rect 7708 11852 7788 11880
rect 7656 11834 7708 11840
rect 7852 11830 7880 12038
rect 7930 11999 7986 12008
rect 7840 11824 7892 11830
rect 7668 11772 7840 11778
rect 7668 11766 7892 11772
rect 7668 11750 7880 11766
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7668 11354 7696 11750
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7748 11552 7800 11558
rect 7852 11529 7880 11630
rect 7748 11494 7800 11500
rect 7838 11520 7894 11529
rect 7760 11370 7788 11494
rect 7838 11455 7894 11464
rect 7656 11348 7708 11354
rect 7760 11342 7880 11370
rect 7656 11290 7708 11296
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7576 10198 7604 10542
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7392 8974 7420 9998
rect 7484 9518 7512 9998
rect 7562 9752 7618 9761
rect 7562 9687 7618 9696
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8566 7420 8774
rect 7484 8634 7512 8871
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6934 6684 7142
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6564 6254 6592 6802
rect 6656 6730 6684 6870
rect 6748 6798 6776 7278
rect 7102 7032 7158 7041
rect 7102 6967 7158 6976
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6550 5944 6606 5953
rect 6472 5902 6550 5930
rect 6656 5914 6684 6258
rect 6550 5879 6606 5888
rect 6644 5908 6696 5914
rect 6564 5846 6592 5879
rect 6644 5850 6696 5856
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5166 6684 5646
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6472 4690 6500 4966
rect 6564 4690 6592 4966
rect 6932 4826 6960 6734
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7024 5234 7052 5782
rect 7116 5710 7144 6967
rect 7288 6248 7340 6254
rect 7392 6236 7420 7958
rect 7340 6208 7420 6236
rect 7288 6190 7340 6196
rect 7300 5914 7328 6190
rect 7576 5914 7604 9687
rect 7668 8430 7696 11290
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10538 7788 10950
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7760 10441 7788 10474
rect 7746 10432 7802 10441
rect 7746 10367 7802 10376
rect 7852 10305 7880 11342
rect 7838 10296 7894 10305
rect 7838 10231 7894 10240
rect 7944 9761 7972 11999
rect 8036 11393 8064 12718
rect 8022 11384 8078 11393
rect 8022 11319 8078 11328
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 10985 8064 11154
rect 8022 10976 8078 10985
rect 8022 10911 8078 10920
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 9353 7788 9522
rect 7840 9512 7892 9518
rect 7892 9472 7972 9500
rect 7840 9454 7892 9460
rect 7746 9344 7802 9353
rect 7746 9279 7802 9288
rect 7746 9072 7802 9081
rect 7746 9007 7802 9016
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7760 8412 7788 9007
rect 7838 8664 7894 8673
rect 7838 8599 7840 8608
rect 7892 8599 7894 8608
rect 7840 8570 7892 8576
rect 7838 8528 7894 8537
rect 7838 8463 7894 8472
rect 7852 8430 7880 8463
rect 7840 8424 7892 8430
rect 7760 8384 7840 8412
rect 7654 7304 7710 7313
rect 7654 7239 7710 7248
rect 7668 7002 7696 7239
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7392 5166 7420 5850
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7470 5536 7526 5545
rect 7470 5471 7526 5480
rect 7484 5166 7512 5471
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6932 4146 6960 4762
rect 7392 4690 7420 5102
rect 7576 4758 7604 5714
rect 7668 5681 7696 6190
rect 7760 5846 7788 8384
rect 7840 8366 7892 8372
rect 7944 8294 7972 9472
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7930 7168 7986 7177
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7748 5704 7800 5710
rect 7654 5672 7710 5681
rect 7748 5646 7800 5652
rect 7654 5607 7710 5616
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7760 4690 7788 5646
rect 7852 5302 7880 7142
rect 7930 7103 7986 7112
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7944 5166 7972 7103
rect 8036 6458 8064 10746
rect 8128 9722 8156 12922
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8220 10962 8248 12854
rect 8312 11830 8340 13806
rect 8390 13696 8446 13705
rect 8390 13631 8446 13640
rect 8404 12306 8432 13631
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8496 13258 8524 13330
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8482 13152 8538 13161
rect 8482 13087 8538 13096
rect 8496 12918 8524 13087
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8588 12753 8616 13330
rect 8680 12900 8708 13942
rect 8772 13841 8800 14418
rect 8864 14006 8892 14826
rect 8956 14550 8984 14991
rect 9140 14940 9168 15456
rect 9220 15438 9272 15444
rect 9232 15094 9260 15438
rect 9220 15088 9272 15094
rect 9220 15030 9272 15036
rect 9140 14912 9260 14940
rect 9036 14884 9088 14890
rect 9088 14844 9168 14872
rect 9036 14826 9088 14832
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9048 14346 9076 14418
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13870 8984 13942
rect 8944 13864 8996 13870
rect 8758 13832 8814 13841
rect 8944 13806 8996 13812
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8758 13767 8814 13776
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8864 13530 8892 13738
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8944 13456 8996 13462
rect 8850 13424 8906 13433
rect 8944 13398 8996 13404
rect 8850 13359 8852 13368
rect 8904 13359 8906 13368
rect 8852 13330 8904 13336
rect 8760 12912 8812 12918
rect 8680 12872 8760 12900
rect 8760 12854 8812 12860
rect 8760 12776 8812 12782
rect 8574 12744 8630 12753
rect 8760 12718 8812 12724
rect 8574 12679 8630 12688
rect 8576 12436 8628 12442
rect 8772 12424 8800 12718
rect 8864 12594 8892 13330
rect 8956 12986 8984 13398
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8864 12566 8984 12594
rect 8576 12378 8628 12384
rect 8680 12396 8800 12424
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8312 11286 8340 11562
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8220 10934 8340 10962
rect 8206 10840 8262 10849
rect 8312 10810 8340 10934
rect 8206 10775 8208 10784
rect 8260 10775 8262 10784
rect 8300 10804 8352 10810
rect 8208 10746 8260 10752
rect 8300 10746 8352 10752
rect 8298 10704 8354 10713
rect 8208 10668 8260 10674
rect 8298 10639 8354 10648
rect 8208 10610 8260 10616
rect 8220 10062 8248 10610
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8128 6730 8156 9386
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9110 8248 9318
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8498 8248 8774
rect 8312 8634 8340 10639
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 8838 8432 9318
rect 8496 8974 8524 12310
rect 8588 12170 8616 12378
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8680 11914 8708 12396
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8588 11886 8708 11914
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8390 8528 8446 8537
rect 8208 8492 8260 8498
rect 8390 8463 8446 8472
rect 8208 8434 8260 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 8265 8340 8366
rect 8298 8256 8354 8265
rect 8298 8191 8354 8200
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 6089 8064 6190
rect 8022 6080 8078 6089
rect 8022 6015 8078 6024
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5724 3664 5776 3670
rect 5724 3606 5776 3612
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 6564 3534 6592 4014
rect 6840 3602 6868 4014
rect 7392 4010 7420 4626
rect 7852 4282 7880 4626
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8036 4282 8064 4422
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7668 4078 7696 4218
rect 8128 4078 8156 6666
rect 8220 4146 8248 7346
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6769 8340 7210
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8404 4622 8432 8463
rect 8496 6866 8524 8774
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 8404 3670 8432 4558
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 8496 2774 8524 6802
rect 8588 5914 8616 11886
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8680 9042 8708 11766
rect 8772 11014 8800 12242
rect 8956 12152 8984 12566
rect 9048 12442 9076 13806
rect 9140 13530 9168 14844
rect 9232 14618 9260 14912
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9140 12714 9168 13466
rect 9218 13288 9274 13297
rect 9218 13223 9274 13232
rect 9232 12730 9260 13223
rect 9324 12850 9352 16050
rect 9508 15978 9536 18391
rect 9692 17954 9720 19343
rect 9862 19272 9918 19281
rect 9862 19207 9918 19216
rect 10048 19236 10100 19242
rect 9876 18834 9904 19207
rect 10048 19178 10100 19184
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9600 17926 9720 17954
rect 9600 17746 9628 17926
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9600 17066 9628 17682
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15881 9536 15914
rect 9494 15872 9550 15881
rect 9494 15807 9550 15816
rect 9600 15706 9628 16594
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9494 15600 9550 15609
rect 9494 15535 9550 15544
rect 9508 15144 9536 15535
rect 9600 15366 9628 15642
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9588 15156 9640 15162
rect 9508 15116 9588 15144
rect 9588 15098 9640 15104
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9600 14550 9628 14894
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9416 13841 9444 14010
rect 9508 14006 9536 14282
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9402 13832 9458 13841
rect 9402 13767 9458 13776
rect 9494 13424 9550 13433
rect 9494 13359 9550 13368
rect 9508 12889 9536 13359
rect 9600 13161 9628 14350
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 9494 12880 9550 12889
rect 9312 12844 9364 12850
rect 9494 12815 9550 12824
rect 9312 12786 9364 12792
rect 9128 12708 9180 12714
rect 9232 12702 9352 12730
rect 9128 12650 9180 12656
rect 9220 12640 9272 12646
rect 9140 12588 9220 12594
rect 9140 12582 9272 12588
rect 9140 12566 9260 12582
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9140 12209 9168 12566
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9126 12200 9182 12209
rect 8956 12124 9076 12152
rect 9232 12170 9260 12242
rect 9324 12209 9352 12702
rect 9496 12232 9548 12238
rect 9310 12200 9366 12209
rect 9126 12135 9182 12144
rect 9220 12164 9272 12170
rect 8942 12064 8998 12073
rect 8942 11999 8998 12008
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11529 8892 11562
rect 8956 11558 8984 11999
rect 9048 11778 9076 12124
rect 9496 12174 9548 12180
rect 9310 12135 9366 12144
rect 9404 12164 9456 12170
rect 9220 12106 9272 12112
rect 9404 12106 9456 12112
rect 9416 12073 9444 12106
rect 9508 12102 9536 12174
rect 9496 12096 9548 12102
rect 9126 12064 9182 12073
rect 9126 11999 9182 12008
rect 9402 12064 9458 12073
rect 9496 12038 9548 12044
rect 9402 11999 9458 12008
rect 9140 11898 9168 11999
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9508 11830 9536 12038
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9496 11824 9548 11830
rect 9048 11750 9260 11778
rect 9496 11766 9548 11772
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8944 11552 8996 11558
rect 8850 11520 8906 11529
rect 8944 11494 8996 11500
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8850 11455 8906 11464
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8850 10976 8906 10985
rect 8850 10911 8906 10920
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8772 10062 8800 10474
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8864 9926 8892 10911
rect 8956 9926 8984 11154
rect 9048 11150 9076 11494
rect 9036 11144 9088 11150
rect 9140 11121 9168 11630
rect 9232 11218 9260 11750
rect 9600 11354 9628 11834
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9220 11212 9272 11218
rect 9496 11212 9548 11218
rect 9220 11154 9272 11160
rect 9324 11172 9496 11200
rect 9036 11086 9088 11092
rect 9126 11112 9182 11121
rect 9126 11047 9182 11056
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10674 9076 10950
rect 9324 10742 9352 11172
rect 9496 11154 9548 11160
rect 9600 11098 9628 11290
rect 9416 11070 9628 11098
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9048 10130 9076 10610
rect 9220 10600 9272 10606
rect 9312 10600 9364 10606
rect 9220 10542 9272 10548
rect 9310 10568 9312 10577
rect 9364 10568 9366 10577
rect 9126 10296 9182 10305
rect 9232 10266 9260 10542
rect 9310 10503 9366 10512
rect 9126 10231 9182 10240
rect 9220 10260 9272 10266
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 9140 9874 9168 10231
rect 9220 10202 9272 10208
rect 9220 9988 9272 9994
rect 9324 9976 9352 10503
rect 9416 10418 9444 11070
rect 9588 11008 9640 11014
rect 9494 10976 9550 10985
rect 9588 10950 9640 10956
rect 9692 10962 9720 17478
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9784 12442 9812 13806
rect 9876 13569 9904 17750
rect 9968 15706 9996 18770
rect 10060 17134 10088 19178
rect 10152 18222 10180 19751
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10244 18057 10272 18770
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10230 18048 10286 18057
rect 10230 17983 10286 17992
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10152 17610 10180 17682
rect 10244 17678 10272 17818
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10244 17134 10272 17614
rect 10336 17542 10364 18158
rect 10428 17882 10456 20839
rect 10520 20398 10548 21100
rect 10600 21082 10652 21088
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10612 20806 10640 20946
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10612 19514 10640 20742
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10508 18148 10560 18154
rect 10508 18090 10560 18096
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10428 17377 10456 17682
rect 10414 17368 10470 17377
rect 10414 17303 10470 17312
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 16250 10088 16526
rect 10152 16250 10180 16662
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 16153 10272 16390
rect 10230 16144 10286 16153
rect 10230 16079 10286 16088
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9954 15328 10010 15337
rect 9954 15263 10010 15272
rect 9968 15026 9996 15263
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9862 13560 9918 13569
rect 9862 13495 9918 13504
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9876 12356 9904 13398
rect 9968 13326 9996 14826
rect 10060 14113 10088 15982
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10060 13161 10088 13330
rect 10046 13152 10102 13161
rect 10046 13087 10102 13096
rect 10152 12696 10180 15846
rect 10244 15570 10272 16079
rect 10336 15570 10364 16458
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10244 15337 10272 15506
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10230 15328 10286 15337
rect 10230 15263 10286 15272
rect 10232 15088 10284 15094
rect 10230 15056 10232 15065
rect 10284 15056 10286 15065
rect 10230 14991 10286 15000
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10244 14385 10272 14554
rect 10230 14376 10286 14385
rect 10230 14311 10286 14320
rect 10336 14328 10364 15370
rect 10428 14482 10456 17070
rect 10520 14958 10548 18090
rect 10612 18057 10640 18090
rect 10598 18048 10654 18057
rect 10598 17983 10654 17992
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10612 17542 10640 17818
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10612 14793 10640 17478
rect 10704 15201 10732 17478
rect 10796 15502 10824 21558
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10980 20806 11008 20946
rect 11152 20868 11204 20874
rect 11256 20856 11284 21082
rect 11348 20942 11376 21490
rect 11440 21146 11468 21626
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11808 21078 11836 21286
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11204 20828 11284 20856
rect 11152 20810 11204 20816
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10980 19990 11008 20334
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 20058 11100 20266
rect 11150 20224 11206 20233
rect 11150 20159 11206 20168
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11072 19514 11100 19858
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11164 18834 11192 20159
rect 11256 19854 11284 20828
rect 11348 20330 11376 20878
rect 11436 20700 11744 20709
rect 11436 20698 11442 20700
rect 11498 20698 11522 20700
rect 11578 20698 11602 20700
rect 11658 20698 11682 20700
rect 11738 20698 11744 20700
rect 11498 20646 11500 20698
rect 11680 20646 11682 20698
rect 11436 20644 11442 20646
rect 11498 20644 11522 20646
rect 11578 20644 11602 20646
rect 11658 20644 11682 20646
rect 11738 20644 11744 20646
rect 11436 20635 11744 20644
rect 11992 20346 12020 21966
rect 26884 21966 26936 21972
rect 12254 21927 12310 21936
rect 13820 21956 13872 21962
rect 12268 21690 12296 21927
rect 13820 21898 13872 21904
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 12806 21720 12862 21729
rect 12256 21684 12308 21690
rect 12806 21655 12808 21664
rect 12256 21626 12308 21632
rect 12860 21655 12862 21664
rect 13358 21720 13414 21729
rect 13358 21655 13360 21664
rect 12808 21626 12860 21632
rect 13412 21655 13414 21664
rect 13360 21626 13412 21632
rect 13832 21622 13860 21898
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 13910 21720 13966 21729
rect 13910 21655 13912 21664
rect 13964 21655 13966 21664
rect 16670 21720 16726 21729
rect 16670 21655 16672 21664
rect 13912 21626 13964 21632
rect 16724 21655 16726 21664
rect 16672 21626 16724 21632
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 18418 21584 18474 21593
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 17224 21548 17276 21554
rect 18418 21519 18420 21528
rect 17224 21490 17276 21496
rect 18472 21519 18474 21528
rect 18420 21490 18472 21496
rect 14370 21448 14426 21457
rect 14280 21412 14332 21418
rect 14370 21383 14426 21392
rect 14280 21354 14332 21360
rect 12096 21244 12404 21253
rect 12096 21242 12102 21244
rect 12158 21242 12182 21244
rect 12238 21242 12262 21244
rect 12318 21242 12342 21244
rect 12398 21242 12404 21244
rect 12158 21190 12160 21242
rect 12340 21190 12342 21242
rect 12096 21188 12102 21190
rect 12158 21188 12182 21190
rect 12238 21188 12262 21190
rect 12318 21188 12342 21190
rect 12398 21188 12404 21190
rect 12096 21179 12404 21188
rect 14292 21146 14320 21354
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 11336 20324 11388 20330
rect 11336 20266 11388 20272
rect 11808 20318 12020 20346
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11348 19378 11376 19722
rect 11436 19612 11744 19621
rect 11436 19610 11442 19612
rect 11498 19610 11522 19612
rect 11578 19610 11602 19612
rect 11658 19610 11682 19612
rect 11738 19610 11744 19612
rect 11498 19558 11500 19610
rect 11680 19558 11682 19610
rect 11436 19556 11442 19558
rect 11498 19556 11522 19558
rect 11578 19556 11602 19558
rect 11658 19556 11682 19558
rect 11738 19556 11744 19558
rect 11436 19547 11744 19556
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11072 18698 11100 18770
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18154 11192 18566
rect 11256 18426 11284 18838
rect 11808 18766 11836 20318
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11900 20097 11928 20198
rect 12096 20156 12404 20165
rect 12096 20154 12102 20156
rect 12158 20154 12182 20156
rect 12238 20154 12262 20156
rect 12318 20154 12342 20156
rect 12398 20154 12404 20156
rect 12158 20102 12160 20154
rect 12340 20102 12342 20154
rect 12096 20100 12102 20102
rect 12158 20100 12182 20102
rect 12238 20100 12262 20102
rect 12318 20100 12342 20102
rect 12398 20100 12404 20102
rect 11886 20088 11942 20097
rect 12096 20091 12404 20100
rect 12452 20058 12480 20878
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12714 20496 12770 20505
rect 12714 20431 12770 20440
rect 11886 20023 11942 20032
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12256 19984 12308 19990
rect 12256 19926 12308 19932
rect 12360 19938 12388 19994
rect 12544 19938 12572 19994
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11992 18952 12020 19858
rect 12084 19514 12112 19858
rect 12268 19802 12296 19926
rect 12360 19910 12572 19938
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12636 19802 12664 19858
rect 12268 19774 12664 19802
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12070 19408 12126 19417
rect 12070 19343 12126 19352
rect 12084 19242 12112 19343
rect 12728 19334 12756 20431
rect 12806 20360 12862 20369
rect 12806 20295 12862 20304
rect 12820 20262 12848 20295
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12820 19446 12848 19858
rect 12912 19718 12940 20742
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 13096 19514 13124 20946
rect 14108 20602 14136 20946
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12440 19304 12492 19310
rect 12728 19306 12940 19334
rect 12440 19246 12492 19252
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12096 19068 12404 19077
rect 12096 19066 12102 19068
rect 12158 19066 12182 19068
rect 12238 19066 12262 19068
rect 12318 19066 12342 19068
rect 12398 19066 12404 19068
rect 12158 19014 12160 19066
rect 12340 19014 12342 19066
rect 12096 19012 12102 19014
rect 12158 19012 12182 19014
rect 12238 19012 12262 19014
rect 12318 19012 12342 19014
rect 12398 19012 12404 19014
rect 12096 19003 12404 19012
rect 12452 18970 12480 19246
rect 12440 18964 12492 18970
rect 11992 18924 12296 18952
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11242 18320 11298 18329
rect 11242 18255 11298 18264
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16833 10916 17070
rect 11072 16998 11100 18090
rect 11256 18086 11284 18255
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11256 17513 11284 17682
rect 11242 17504 11298 17513
rect 11242 17439 11298 17448
rect 11348 17338 11376 18634
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11436 18524 11744 18533
rect 11436 18522 11442 18524
rect 11498 18522 11522 18524
rect 11578 18522 11602 18524
rect 11658 18522 11682 18524
rect 11738 18522 11744 18524
rect 11498 18470 11500 18522
rect 11680 18470 11682 18522
rect 11436 18468 11442 18470
rect 11498 18468 11522 18470
rect 11578 18468 11602 18470
rect 11658 18468 11682 18470
rect 11738 18468 11744 18470
rect 11436 18459 11744 18468
rect 11808 18222 11836 18566
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11436 17436 11744 17445
rect 11436 17434 11442 17436
rect 11498 17434 11522 17436
rect 11578 17434 11602 17436
rect 11658 17434 11682 17436
rect 11738 17434 11744 17436
rect 11498 17382 11500 17434
rect 11680 17382 11682 17434
rect 11436 17380 11442 17382
rect 11498 17380 11522 17382
rect 11578 17380 11602 17382
rect 11658 17380 11682 17382
rect 11738 17380 11744 17382
rect 11436 17371 11744 17380
rect 11808 17338 11836 17682
rect 11992 17542 12020 18702
rect 12084 18290 12112 18702
rect 12176 18630 12204 18770
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12268 18086 12296 18924
rect 12440 18906 12492 18912
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12636 18154 12664 18294
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12096 17980 12404 17989
rect 12096 17978 12102 17980
rect 12158 17978 12182 17980
rect 12238 17978 12262 17980
rect 12318 17978 12342 17980
rect 12398 17978 12404 17980
rect 12158 17926 12160 17978
rect 12340 17926 12342 17978
rect 12096 17924 12102 17926
rect 12158 17924 12182 17926
rect 12238 17924 12262 17926
rect 12318 17924 12342 17926
rect 12398 17924 12404 17926
rect 12096 17915 12404 17924
rect 12530 17912 12586 17921
rect 12452 17870 12530 17898
rect 12452 17728 12480 17870
rect 12530 17847 12586 17856
rect 12360 17700 12480 17728
rect 12622 17776 12678 17785
rect 12820 17746 12848 18090
rect 12622 17711 12678 17720
rect 12716 17740 12768 17746
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 12164 17536 12216 17542
rect 12360 17513 12388 17700
rect 12636 17678 12664 17711
rect 12716 17682 12768 17688
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12164 17478 12216 17484
rect 12346 17504 12402 17513
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12176 17202 12204 17478
rect 12346 17439 12402 17448
rect 12452 17377 12480 17546
rect 12532 17536 12584 17542
rect 12530 17504 12532 17513
rect 12584 17504 12586 17513
rect 12530 17439 12586 17448
rect 12438 17368 12494 17377
rect 12438 17303 12494 17312
rect 12728 17270 12756 17682
rect 12716 17264 12768 17270
rect 12820 17241 12848 17682
rect 12716 17206 12768 17212
rect 12806 17232 12862 17241
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12452 17156 12664 17184
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10874 16824 10930 16833
rect 10874 16759 10930 16768
rect 11150 16824 11206 16833
rect 11150 16759 11206 16768
rect 11164 16658 11192 16759
rect 11348 16674 11376 17070
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11532 16776 11560 16934
rect 11612 16788 11664 16794
rect 11532 16748 11612 16776
rect 11612 16730 11664 16736
rect 11152 16652 11204 16658
rect 11348 16646 11468 16674
rect 11152 16594 11204 16600
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11336 16584 11388 16590
rect 11440 16574 11468 16646
rect 11624 16612 11744 16640
rect 11624 16574 11652 16612
rect 11440 16546 11652 16574
rect 11336 16526 11388 16532
rect 11072 16454 11100 16526
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10966 16280 11022 16289
rect 11348 16250 11376 16526
rect 11716 16522 11744 16612
rect 11808 16572 11836 17070
rect 11992 16794 12020 17138
rect 12452 17066 12480 17156
rect 12530 17096 12586 17105
rect 12440 17060 12492 17066
rect 12530 17031 12586 17040
rect 12440 17002 12492 17008
rect 12096 16892 12404 16901
rect 12096 16890 12102 16892
rect 12158 16890 12182 16892
rect 12238 16890 12262 16892
rect 12318 16890 12342 16892
rect 12398 16890 12404 16892
rect 12158 16838 12160 16890
rect 12340 16838 12342 16890
rect 12096 16836 12102 16838
rect 12158 16836 12182 16838
rect 12238 16836 12262 16838
rect 12318 16836 12342 16838
rect 12398 16836 12404 16838
rect 12096 16827 12404 16836
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12072 16584 12124 16590
rect 11808 16544 12072 16572
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11436 16348 11744 16357
rect 11436 16346 11442 16348
rect 11498 16346 11522 16348
rect 11578 16346 11602 16348
rect 11658 16346 11682 16348
rect 11738 16346 11744 16348
rect 11498 16294 11500 16346
rect 11680 16294 11682 16346
rect 11436 16292 11442 16294
rect 11498 16292 11522 16294
rect 11578 16292 11602 16294
rect 11658 16292 11682 16294
rect 11738 16292 11744 16294
rect 11436 16283 11744 16292
rect 10966 16215 11022 16224
rect 11336 16244 11388 16250
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10888 15638 10916 15914
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10690 15192 10746 15201
rect 10690 15127 10746 15136
rect 10782 15056 10838 15065
rect 10782 14991 10838 15000
rect 10598 14784 10654 14793
rect 10598 14719 10654 14728
rect 10796 14618 10824 14991
rect 10888 14890 10916 15438
rect 10980 15434 11008 16215
rect 11336 16186 11388 16192
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11336 16040 11388 16046
rect 11150 16008 11206 16017
rect 11624 16028 11652 16186
rect 11704 16040 11756 16046
rect 11624 16000 11704 16028
rect 11336 15982 11388 15988
rect 11704 15982 11756 15988
rect 11150 15943 11206 15952
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11072 15201 11100 15370
rect 11058 15192 11114 15201
rect 11058 15127 11114 15136
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10966 14920 11022 14929
rect 10876 14884 10928 14890
rect 10966 14855 11022 14864
rect 10876 14826 10928 14832
rect 10874 14784 10930 14793
rect 10874 14719 10930 14728
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10508 14544 10560 14550
rect 10506 14512 10508 14521
rect 10560 14512 10562 14521
rect 10416 14476 10468 14482
rect 10690 14512 10746 14521
rect 10506 14447 10562 14456
rect 10600 14476 10652 14482
rect 10416 14418 10468 14424
rect 10690 14447 10746 14456
rect 10784 14476 10836 14482
rect 10600 14418 10652 14424
rect 10336 14300 10548 14328
rect 10520 14074 10548 14300
rect 10612 14249 10640 14418
rect 10598 14240 10654 14249
rect 10598 14175 10654 14184
rect 10598 14104 10654 14113
rect 10508 14068 10560 14074
rect 10598 14039 10654 14048
rect 10508 14010 10560 14016
rect 10612 13938 10640 14039
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10336 13394 10364 13806
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10414 13560 10470 13569
rect 10414 13495 10470 13504
rect 10428 13394 10456 13495
rect 10520 13462 10548 13738
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10232 12912 10284 12918
rect 10230 12880 10232 12889
rect 10284 12880 10286 12889
rect 10230 12815 10286 12824
rect 10060 12668 10180 12696
rect 9876 12328 9996 12356
rect 9770 11656 9826 11665
rect 9770 11591 9826 11600
rect 9784 11218 9812 11591
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9494 10911 9550 10920
rect 9508 10674 9536 10911
rect 9600 10742 9628 10950
rect 9692 10934 9904 10962
rect 9770 10840 9826 10849
rect 9692 10798 9770 10826
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9416 10390 9536 10418
rect 9402 10296 9458 10305
rect 9402 10231 9458 10240
rect 9416 10198 9444 10231
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9508 10112 9536 10390
rect 9600 10305 9628 10678
rect 9692 10470 9720 10798
rect 9770 10775 9826 10784
rect 9876 10690 9904 10934
rect 9784 10662 9904 10690
rect 9784 10606 9812 10662
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9784 10470 9812 10542
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9586 10296 9642 10305
rect 9692 10266 9720 10406
rect 9586 10231 9642 10240
rect 9680 10260 9732 10266
rect 9876 10248 9904 10542
rect 9680 10202 9732 10208
rect 9784 10220 9904 10248
rect 9588 10124 9640 10130
rect 9508 10084 9588 10112
rect 9588 10066 9640 10072
rect 9404 10056 9456 10062
rect 9456 10016 9536 10044
rect 9404 9998 9456 10004
rect 9272 9948 9352 9976
rect 9220 9930 9272 9936
rect 9508 9926 9536 10016
rect 9496 9920 9548 9926
rect 8864 9654 8892 9862
rect 9140 9846 9260 9874
rect 9496 9862 9548 9868
rect 9678 9888 9734 9897
rect 8852 9648 8904 9654
rect 9128 9648 9180 9654
rect 8852 9590 8904 9596
rect 9126 9616 9128 9625
rect 9180 9616 9182 9625
rect 9126 9551 9182 9560
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8772 9382 8800 9454
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8758 8528 8814 8537
rect 8758 8463 8760 8472
rect 8812 8463 8814 8472
rect 8760 8434 8812 8440
rect 8852 8424 8904 8430
rect 8772 8372 8852 8378
rect 8772 8366 8904 8372
rect 8772 8350 8892 8366
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 7177 8708 8230
rect 8772 8022 8800 8350
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8864 7886 8892 8230
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8772 7449 8800 7822
rect 8850 7576 8906 7585
rect 8850 7511 8906 7520
rect 8758 7440 8814 7449
rect 8758 7375 8814 7384
rect 8666 7168 8722 7177
rect 8666 7103 8722 7112
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8680 6322 8708 6802
rect 8772 6746 8800 7375
rect 8864 7342 8892 7511
rect 8956 7410 8984 8978
rect 9048 8838 9076 9454
rect 9232 9042 9260 9846
rect 9508 9602 9536 9862
rect 9678 9823 9734 9832
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9324 9574 9536 9602
rect 9324 9518 9352 9574
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9140 8537 9168 8774
rect 9126 8528 9182 8537
rect 9126 8463 9182 8472
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9048 8022 9076 8366
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9324 7886 9352 9318
rect 9416 9178 9444 9454
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9416 8634 9444 8978
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9402 8256 9458 8265
rect 9402 8191 9458 8200
rect 9416 8090 9444 8191
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 7954 9444 8026
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9508 7818 9536 9574
rect 9600 9110 9628 9658
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9128 7744 9180 7750
rect 9034 7712 9090 7721
rect 9128 7686 9180 7692
rect 9034 7647 9090 7656
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8864 6866 8892 7278
rect 8956 7002 8984 7346
rect 9048 7342 9076 7647
rect 9140 7546 9168 7686
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9034 7168 9090 7177
rect 9034 7103 9090 7112
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8772 6718 8892 6746
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 5574 8616 5714
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8772 4146 8800 6598
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 2056 2746 2268 2774
rect 2240 2582 2268 2746
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 8312 2746 8524 2774
rect 2228 2576 2280 2582
rect 2228 2518 2280 2524
rect 8312 2514 8340 2746
rect 8864 2553 8892 6718
rect 9048 5574 9076 7103
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9232 6780 9260 6870
rect 9312 6792 9364 6798
rect 9232 6752 9312 6780
rect 9312 6734 9364 6740
rect 9416 6474 9444 7482
rect 9508 7002 9536 7754
rect 9600 7546 9628 8055
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9600 6866 9628 7375
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9416 6446 9536 6474
rect 9402 6216 9458 6225
rect 9402 6151 9458 6160
rect 9416 5914 9444 6151
rect 9508 6089 9536 6446
rect 9494 6080 9550 6089
rect 9494 6015 9550 6024
rect 9404 5908 9456 5914
rect 9324 5868 9404 5896
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9232 5642 9260 5782
rect 9324 5778 9352 5868
rect 9404 5850 9456 5856
rect 9508 5778 9536 6015
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9416 5098 9444 5714
rect 9692 5710 9720 9823
rect 9784 9722 9812 10220
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9876 9926 9904 10066
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9784 8906 9812 9658
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9770 8800 9826 8809
rect 9770 8735 9826 8744
rect 9784 7868 9812 8735
rect 9876 8294 9904 9862
rect 9968 8430 9996 12328
rect 10060 11914 10088 12668
rect 10244 12628 10272 12815
rect 10428 12782 10456 13330
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10520 12850 10548 13262
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10152 12600 10272 12628
rect 10152 12306 10180 12600
rect 10140 12300 10192 12306
rect 10520 12288 10548 12786
rect 10140 12242 10192 12248
rect 10428 12260 10548 12288
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 12073 10180 12106
rect 10244 12102 10272 12174
rect 10232 12096 10284 12102
rect 10138 12064 10194 12073
rect 10232 12038 10284 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10138 11999 10194 12008
rect 10060 11886 10272 11914
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10060 9160 10088 11766
rect 10152 10985 10180 11766
rect 10244 11257 10272 11886
rect 10336 11830 10364 12038
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10428 11694 10456 12260
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10230 11248 10286 11257
rect 10286 11206 10364 11234
rect 10230 11183 10286 11192
rect 10232 11008 10284 11014
rect 10138 10976 10194 10985
rect 10232 10950 10284 10956
rect 10138 10911 10194 10920
rect 10138 10704 10194 10713
rect 10138 10639 10194 10648
rect 10152 10606 10180 10639
rect 10244 10606 10272 10950
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10266 10272 10406
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10152 9897 10180 10202
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10138 9888 10194 9897
rect 10138 9823 10194 9832
rect 10244 9738 10272 10066
rect 10336 10062 10364 11206
rect 10428 11014 10456 11494
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10152 9710 10272 9738
rect 10152 9382 10180 9710
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10140 9376 10192 9382
rect 10244 9353 10272 9522
rect 10140 9318 10192 9324
rect 10230 9344 10286 9353
rect 10230 9279 10286 9288
rect 10232 9172 10284 9178
rect 10060 9132 10180 9160
rect 10046 9072 10102 9081
rect 10046 9007 10048 9016
rect 10100 9007 10102 9016
rect 10048 8978 10100 8984
rect 10152 8906 10180 9132
rect 10232 9114 10284 9120
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10138 8800 10194 8809
rect 10138 8735 10194 8744
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9968 7954 9996 8366
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9864 7880 9916 7886
rect 9784 7840 9864 7868
rect 9864 7822 9916 7828
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 6934 9812 7142
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9784 5778 9812 6870
rect 9876 5953 9904 7822
rect 9954 7576 10010 7585
rect 9954 7511 10010 7520
rect 9968 7478 9996 7511
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9862 5944 9918 5953
rect 9862 5879 9918 5888
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 5234 9720 5646
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9600 4690 9628 5102
rect 9680 4752 9732 4758
rect 9784 4740 9812 5714
rect 9732 4712 9812 4740
rect 9680 4694 9732 4700
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9416 4185 9444 4626
rect 9402 4176 9458 4185
rect 9402 4111 9458 4120
rect 9508 4078 9536 4626
rect 9678 4584 9734 4593
rect 9678 4519 9734 4528
rect 9692 4146 9720 4519
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9784 4078 9812 4422
rect 9876 4146 9904 5879
rect 9968 4185 9996 7414
rect 10060 6662 10088 7890
rect 10152 7274 10180 8735
rect 10244 8022 10272 9114
rect 10336 9081 10364 9522
rect 10428 9178 10456 10610
rect 10520 10577 10548 12106
rect 10612 11914 10640 13330
rect 10704 12714 10732 14447
rect 10784 14418 10836 14424
rect 10796 13705 10824 14418
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10704 12374 10732 12650
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10704 12073 10732 12310
rect 10796 12102 10824 13398
rect 10888 13161 10916 14719
rect 10980 13258 11008 14855
rect 11072 14113 11100 15030
rect 11164 14940 11192 15943
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11256 15094 11284 15506
rect 11348 15094 11376 15982
rect 11702 15736 11758 15745
rect 11702 15671 11758 15680
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11624 15366 11652 15574
rect 11612 15360 11664 15366
rect 11716 15348 11744 15671
rect 11808 15484 11836 16544
rect 12072 16526 12124 16532
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 11888 16448 11940 16454
rect 11886 16416 11888 16425
rect 11980 16448 12032 16454
rect 11940 16416 11942 16425
rect 11980 16390 12032 16396
rect 11886 16351 11942 16360
rect 11888 16244 11940 16250
rect 11992 16232 12020 16390
rect 12360 16289 12388 16458
rect 11940 16204 12020 16232
rect 12346 16280 12402 16289
rect 12346 16215 12402 16224
rect 11888 16186 11940 16192
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12162 16144 12218 16153
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11900 15706 11928 15982
rect 12084 15978 12112 16118
rect 12452 16114 12480 16730
rect 12544 16658 12572 17031
rect 12636 16810 12664 17156
rect 12728 16998 12756 17206
rect 12806 17167 12862 17176
rect 12716 16992 12768 16998
rect 12714 16960 12716 16969
rect 12768 16960 12770 16969
rect 12714 16895 12770 16904
rect 12714 16824 12770 16833
rect 12636 16782 12714 16810
rect 12912 16794 12940 19306
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 13004 19122 13032 19178
rect 13082 19136 13138 19145
rect 13004 19094 13082 19122
rect 13082 19071 13138 19080
rect 13096 18834 13124 19071
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12990 17912 13046 17921
rect 12990 17847 13046 17856
rect 12714 16759 12770 16768
rect 12900 16788 12952 16794
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12530 16280 12586 16289
rect 12530 16215 12586 16224
rect 12162 16079 12218 16088
rect 12440 16108 12492 16114
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 12176 15910 12204 16079
rect 12440 16050 12492 16056
rect 12544 16046 12572 16215
rect 12728 16114 12756 16759
rect 12900 16730 12952 16736
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12440 15904 12492 15910
rect 12544 15881 12572 15982
rect 12440 15846 12492 15852
rect 12530 15872 12586 15881
rect 12096 15804 12404 15813
rect 12096 15802 12102 15804
rect 12158 15802 12182 15804
rect 12238 15802 12262 15804
rect 12318 15802 12342 15804
rect 12398 15802 12404 15804
rect 12158 15750 12160 15802
rect 12340 15750 12342 15802
rect 12096 15748 12102 15750
rect 12158 15748 12182 15750
rect 12238 15748 12262 15750
rect 12318 15748 12342 15750
rect 12398 15748 12404 15750
rect 12096 15739 12404 15748
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12452 15638 12480 15846
rect 12530 15807 12586 15816
rect 12636 15745 12664 15982
rect 12622 15736 12678 15745
rect 12622 15671 12678 15680
rect 11980 15632 12032 15638
rect 12440 15632 12492 15638
rect 12032 15592 12204 15620
rect 11980 15574 12032 15580
rect 11808 15456 12020 15484
rect 11716 15320 11836 15348
rect 11612 15302 11664 15308
rect 11436 15260 11744 15269
rect 11436 15258 11442 15260
rect 11498 15258 11522 15260
rect 11578 15258 11602 15260
rect 11658 15258 11682 15260
rect 11738 15258 11744 15260
rect 11498 15206 11500 15258
rect 11680 15206 11682 15258
rect 11436 15204 11442 15206
rect 11498 15204 11522 15206
rect 11578 15204 11602 15206
rect 11658 15204 11682 15206
rect 11738 15204 11744 15206
rect 11436 15195 11744 15204
rect 11808 15178 11836 15320
rect 11886 15192 11942 15201
rect 11808 15150 11886 15178
rect 11886 15127 11942 15136
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11518 15056 11574 15065
rect 11164 14912 11284 14940
rect 11256 14414 11284 14912
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11244 14408 11296 14414
rect 11348 14396 11376 15030
rect 11518 14991 11574 15000
rect 11532 14958 11560 14991
rect 11428 14952 11480 14958
rect 11426 14920 11428 14929
rect 11520 14952 11572 14958
rect 11480 14920 11482 14929
rect 11520 14894 11572 14900
rect 11426 14855 11482 14864
rect 11992 14600 12020 15456
rect 12070 15328 12126 15337
rect 12070 15263 12126 15272
rect 12084 14958 12112 15263
rect 12176 14958 12204 15592
rect 12440 15574 12492 15580
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12438 15192 12494 15201
rect 12438 15127 12494 15136
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12096 14716 12404 14725
rect 12096 14714 12102 14716
rect 12158 14714 12182 14716
rect 12238 14714 12262 14716
rect 12318 14714 12342 14716
rect 12398 14714 12404 14716
rect 12158 14662 12160 14714
rect 12340 14662 12342 14714
rect 12096 14660 12102 14662
rect 12158 14660 12182 14662
rect 12238 14660 12262 14662
rect 12318 14660 12342 14662
rect 12398 14660 12404 14662
rect 12096 14651 12404 14660
rect 11992 14572 12204 14600
rect 11612 14476 11664 14482
rect 12072 14476 12124 14482
rect 11664 14436 12020 14464
rect 11612 14418 11664 14424
rect 11520 14408 11572 14414
rect 11348 14368 11520 14396
rect 11244 14350 11296 14356
rect 11520 14350 11572 14356
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10874 13152 10930 13161
rect 10874 13087 10930 13096
rect 10966 13016 11022 13025
rect 10966 12951 11022 12960
rect 10980 12918 11008 12951
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 11072 12617 11100 13942
rect 11164 13734 11192 14350
rect 11992 14249 12020 14436
rect 12072 14418 12124 14424
rect 11978 14240 12034 14249
rect 11436 14172 11744 14181
rect 11978 14175 12034 14184
rect 11436 14170 11442 14172
rect 11498 14170 11522 14172
rect 11578 14170 11602 14172
rect 11658 14170 11682 14172
rect 11738 14170 11744 14172
rect 11498 14118 11500 14170
rect 11680 14118 11682 14170
rect 11436 14116 11442 14118
rect 11498 14116 11522 14118
rect 11578 14116 11602 14118
rect 11658 14116 11682 14118
rect 11738 14116 11744 14118
rect 11242 14104 11298 14113
rect 11436 14107 11744 14116
rect 11242 14039 11298 14048
rect 11612 14068 11664 14074
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11256 13530 11284 14039
rect 11612 14010 11664 14016
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11624 13394 11652 14010
rect 11702 13560 11758 13569
rect 11808 13530 11836 14010
rect 12084 13716 12112 14418
rect 12176 13852 12204 14572
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12268 14006 12296 14350
rect 12452 14346 12480 15127
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12544 14074 12572 15506
rect 12636 15337 12664 15671
rect 12622 15328 12678 15337
rect 12622 15263 12678 15272
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 14249 12664 14418
rect 12622 14240 12678 14249
rect 12622 14175 12678 14184
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12176 13824 12480 13852
rect 11900 13688 12112 13716
rect 11702 13495 11758 13504
rect 11796 13524 11848 13530
rect 11716 13462 11744 13495
rect 11796 13466 11848 13472
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11336 13388 11388 13394
rect 11256 13348 11336 13376
rect 11150 13288 11206 13297
rect 11150 13223 11206 13232
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 11164 12481 11192 13223
rect 11150 12472 11206 12481
rect 11150 12407 11206 12416
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10784 12096 10836 12102
rect 10690 12064 10746 12073
rect 10888 12073 10916 12174
rect 10784 12038 10836 12044
rect 10874 12064 10930 12073
rect 10690 11999 10746 12008
rect 10612 11886 10732 11914
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10506 10568 10562 10577
rect 10506 10503 10562 10512
rect 10612 10452 10640 11766
rect 10704 11150 10732 11886
rect 10796 11676 10824 12038
rect 10874 11999 10930 12008
rect 10980 11937 11008 12310
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10966 11928 11022 11937
rect 10966 11863 11022 11872
rect 11072 11830 11100 12174
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 11164 11694 11192 12106
rect 10876 11688 10928 11694
rect 10796 11648 10876 11676
rect 10876 11630 10928 11636
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11354 10916 11494
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10782 11248 10838 11257
rect 10782 11183 10838 11192
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10704 10742 10732 11086
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10692 10578 10744 10584
rect 10692 10520 10744 10526
rect 10520 10424 10640 10452
rect 10520 10130 10548 10424
rect 10598 10296 10654 10305
rect 10704 10266 10732 10520
rect 10598 10231 10654 10240
rect 10692 10260 10744 10266
rect 10612 10198 10640 10231
rect 10692 10202 10744 10208
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10506 9752 10562 9761
rect 10704 9738 10732 10066
rect 10562 9710 10732 9738
rect 10506 9687 10562 9696
rect 10520 9586 10548 9687
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10322 9072 10378 9081
rect 10322 9007 10378 9016
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10152 6866 10180 7210
rect 10244 7206 10272 7958
rect 10336 7562 10364 8774
rect 10520 8430 10548 9318
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10428 7750 10456 8230
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10336 7534 10456 7562
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10152 6458 10180 6802
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 6633 10272 6666
rect 10230 6624 10286 6633
rect 10230 6559 10286 6568
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10244 6254 10272 6559
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5846 10364 6054
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10046 4856 10102 4865
rect 10046 4791 10102 4800
rect 10060 4622 10088 4791
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10152 4282 10180 5782
rect 10428 5370 10456 7534
rect 10520 7342 10548 8366
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10612 6934 10640 9318
rect 10704 8634 10732 9318
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 8129 10732 8434
rect 10690 8120 10746 8129
rect 10690 8055 10746 8064
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10520 6254 10548 6802
rect 10690 6488 10746 6497
rect 10690 6423 10746 6432
rect 10704 6254 10732 6423
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10416 4752 10468 4758
rect 10336 4712 10416 4740
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4282 10272 4558
rect 10336 4486 10364 4712
rect 10416 4694 10468 4700
rect 10416 4616 10468 4622
rect 10414 4584 10416 4593
rect 10468 4584 10470 4593
rect 10414 4519 10470 4528
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9954 4176 10010 4185
rect 9864 4140 9916 4146
rect 9954 4111 10010 4120
rect 9864 4082 9916 4088
rect 10428 4078 10456 4422
rect 10520 4078 10548 6190
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5778 10640 6054
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 4078 10640 5714
rect 10796 5710 10824 11183
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10606 10916 11086
rect 11256 11064 11284 13348
rect 11336 13330 11388 13336
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 13190 11836 13330
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11436 13084 11744 13093
rect 11436 13082 11442 13084
rect 11498 13082 11522 13084
rect 11578 13082 11602 13084
rect 11658 13082 11682 13084
rect 11738 13082 11744 13084
rect 11498 13030 11500 13082
rect 11680 13030 11682 13082
rect 11436 13028 11442 13030
rect 11498 13028 11522 13030
rect 11578 13028 11602 13030
rect 11658 13028 11682 13030
rect 11738 13028 11744 13030
rect 11436 13019 11744 13028
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11348 12617 11376 12650
rect 11520 12640 11572 12646
rect 11334 12608 11390 12617
rect 11520 12582 11572 12588
rect 11334 12543 11390 12552
rect 11532 12306 11560 12582
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11624 12152 11652 12922
rect 11900 12764 11928 13688
rect 12096 13628 12404 13637
rect 12096 13626 12102 13628
rect 12158 13626 12182 13628
rect 12238 13626 12262 13628
rect 12318 13626 12342 13628
rect 12398 13626 12404 13628
rect 12158 13574 12160 13626
rect 12340 13574 12342 13626
rect 12096 13572 12102 13574
rect 12158 13572 12182 13574
rect 12238 13572 12262 13574
rect 12318 13572 12342 13574
rect 12398 13572 12404 13574
rect 12096 13563 12404 13572
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12256 13524 12308 13530
rect 12452 13512 12480 13824
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12308 13484 12480 13512
rect 12530 13560 12586 13569
rect 12530 13495 12532 13504
rect 12256 13466 12308 13472
rect 12584 13495 12586 13504
rect 12532 13466 12584 13472
rect 11896 12736 11928 12764
rect 11896 12696 11924 12736
rect 11896 12668 11928 12696
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12164 11756 12170
rect 11624 12124 11704 12152
rect 11704 12106 11756 12112
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11808 12050 11836 12582
rect 11900 12238 11928 12668
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11348 11880 11376 12038
rect 11808 12022 11928 12050
rect 11436 11996 11744 12005
rect 11436 11994 11442 11996
rect 11498 11994 11522 11996
rect 11578 11994 11602 11996
rect 11658 11994 11682 11996
rect 11738 11994 11744 11996
rect 11498 11942 11500 11994
rect 11680 11942 11682 11994
rect 11436 11940 11442 11942
rect 11498 11940 11522 11942
rect 11578 11940 11602 11942
rect 11658 11940 11682 11942
rect 11738 11940 11744 11942
rect 11436 11931 11744 11940
rect 11796 11892 11848 11898
rect 11348 11852 11468 11880
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 11558 11376 11698
rect 11440 11694 11468 11852
rect 11796 11834 11848 11840
rect 11702 11792 11758 11801
rect 11702 11727 11758 11736
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11532 11370 11560 11630
rect 11716 11558 11744 11727
rect 11808 11694 11836 11834
rect 11900 11762 11928 12022
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11992 11694 12020 13466
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12084 12628 12112 13262
rect 12268 13025 12296 13262
rect 12254 13016 12310 13025
rect 12164 12980 12216 12986
rect 12254 12951 12310 12960
rect 12348 12980 12400 12986
rect 12164 12922 12216 12928
rect 12348 12922 12400 12928
rect 12176 12889 12204 12922
rect 12162 12880 12218 12889
rect 12360 12866 12388 12922
rect 12452 12866 12480 13262
rect 12360 12838 12480 12866
rect 12162 12815 12218 12824
rect 12440 12776 12492 12782
rect 12544 12764 12572 13262
rect 12636 12918 12664 13670
rect 12728 13326 12756 14894
rect 12820 14346 12848 16594
rect 13004 16096 13032 17847
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13096 17542 13124 17682
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 13096 16658 13124 17206
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12912 16068 13032 16096
rect 12912 15570 12940 16068
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 13004 15881 13032 15914
rect 12990 15872 13046 15881
rect 12990 15807 13046 15816
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 13004 15144 13032 15506
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12912 15116 13032 15144
rect 12912 14890 12940 15116
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 13004 14657 13032 14962
rect 12990 14648 13046 14657
rect 12990 14583 13046 14592
rect 13096 14521 13124 15438
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12806 13696 12862 13705
rect 12806 13631 12862 13640
rect 12820 13410 12848 13631
rect 12912 13530 12940 14350
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 13938 13124 14282
rect 13188 14074 13216 19790
rect 13464 19786 13492 20402
rect 13740 20398 13768 20538
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 14016 20058 14044 20334
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13266 19544 13322 19553
rect 13266 19479 13322 19488
rect 13280 19378 13308 19479
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13372 18952 13400 19654
rect 13464 19242 13492 19722
rect 13556 19428 13584 19858
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13726 19544 13782 19553
rect 13726 19479 13782 19488
rect 13636 19440 13688 19446
rect 13556 19400 13636 19428
rect 13556 19310 13584 19400
rect 13636 19382 13688 19388
rect 13740 19378 13768 19479
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13648 18970 13676 19246
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13740 19145 13768 19178
rect 13726 19136 13782 19145
rect 13782 19094 13860 19122
rect 13726 19071 13782 19080
rect 13280 18924 13400 18952
rect 13636 18964 13688 18970
rect 13280 15094 13308 18924
rect 13636 18906 13688 18912
rect 13452 18896 13504 18902
rect 13372 18856 13452 18884
rect 13372 16794 13400 18856
rect 13452 18838 13504 18844
rect 13542 18864 13598 18873
rect 13542 18799 13598 18808
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13358 15872 13414 15881
rect 13358 15807 13414 15816
rect 13372 15609 13400 15807
rect 13358 15600 13414 15609
rect 13358 15535 13414 15544
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13280 14482 13308 14894
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13266 14376 13322 14385
rect 13266 14311 13322 14320
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13280 13705 13308 14311
rect 13372 13734 13400 15302
rect 13464 15026 13492 18022
rect 13556 17184 13584 18799
rect 13726 18728 13782 18737
rect 13726 18663 13782 18672
rect 13636 18216 13688 18222
rect 13634 18184 13636 18193
rect 13688 18184 13690 18193
rect 13634 18119 13690 18128
rect 13740 17746 13768 18663
rect 13832 18222 13860 19094
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13740 17241 13768 17478
rect 13818 17368 13874 17377
rect 13818 17303 13874 17312
rect 13726 17232 13782 17241
rect 13556 17156 13676 17184
rect 13726 17167 13782 17176
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13556 16833 13584 17002
rect 13542 16824 13598 16833
rect 13542 16759 13598 16768
rect 13648 16674 13676 17156
rect 13726 17096 13782 17105
rect 13726 17031 13782 17040
rect 13740 16998 13768 17031
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13832 16833 13860 17303
rect 13818 16824 13874 16833
rect 13818 16759 13874 16768
rect 13556 16646 13676 16674
rect 13820 16652 13872 16658
rect 13556 16017 13584 16646
rect 13820 16594 13872 16600
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13728 16584 13780 16590
rect 13832 16561 13860 16594
rect 13728 16526 13780 16532
rect 13818 16552 13874 16561
rect 13542 16008 13598 16017
rect 13648 15978 13676 16526
rect 13740 16028 13768 16526
rect 13818 16487 13874 16496
rect 13820 16040 13872 16046
rect 13740 16000 13820 16028
rect 13820 15982 13872 15988
rect 13542 15943 13598 15952
rect 13636 15972 13688 15978
rect 13556 15706 13584 15943
rect 13636 15914 13688 15920
rect 13544 15700 13596 15706
rect 13648 15688 13676 15914
rect 13832 15910 13860 15982
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13820 15700 13872 15706
rect 13648 15660 13820 15688
rect 13544 15642 13596 15648
rect 13820 15642 13872 15648
rect 13636 15564 13688 15570
rect 13556 15524 13636 15552
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13556 14906 13584 15524
rect 13636 15506 13688 15512
rect 13648 15450 13676 15506
rect 13648 15422 13768 15450
rect 13636 15360 13688 15366
rect 13740 15348 13768 15422
rect 13820 15360 13872 15366
rect 13740 15320 13820 15348
rect 13636 15302 13688 15308
rect 13820 15302 13872 15308
rect 13464 14878 13584 14906
rect 13360 13728 13412 13734
rect 13266 13696 13322 13705
rect 13360 13670 13412 13676
rect 13266 13631 13322 13640
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12820 13382 12940 13410
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12716 12776 12768 12782
rect 12492 12736 12572 12764
rect 12636 12736 12716 12764
rect 12440 12718 12492 12724
rect 12084 12600 12572 12628
rect 12096 12540 12404 12549
rect 12096 12538 12102 12540
rect 12158 12538 12182 12540
rect 12238 12538 12262 12540
rect 12318 12538 12342 12540
rect 12398 12538 12404 12540
rect 12158 12486 12160 12538
rect 12340 12486 12342 12538
rect 12096 12484 12102 12486
rect 12158 12484 12182 12486
rect 12238 12484 12262 12486
rect 12318 12484 12342 12486
rect 12398 12484 12404 12486
rect 12096 12475 12404 12484
rect 12072 12368 12124 12374
rect 12124 12316 12204 12322
rect 12072 12310 12204 12316
rect 12084 12294 12204 12310
rect 12070 12200 12126 12209
rect 12070 12135 12126 12144
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11532 11342 11652 11370
rect 11624 11268 11652 11342
rect 11704 11280 11756 11286
rect 11624 11240 11704 11268
rect 11428 11212 11480 11218
rect 11072 11036 11284 11064
rect 11348 11172 11428 11200
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10888 10062 10916 10406
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10888 9761 10916 9998
rect 10874 9752 10930 9761
rect 10874 9687 10930 9696
rect 10874 9344 10930 9353
rect 10874 9279 10930 9288
rect 10888 5817 10916 9279
rect 10980 8809 11008 10678
rect 10966 8800 11022 8809
rect 10966 8735 11022 8744
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 8401 11008 8434
rect 10966 8392 11022 8401
rect 10966 8327 11022 8336
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 7546 11008 7890
rect 11072 7546 11100 11036
rect 11348 10962 11376 11172
rect 11428 11154 11480 11160
rect 11624 11121 11652 11240
rect 11704 11222 11756 11228
rect 11610 11112 11666 11121
rect 11610 11047 11666 11056
rect 11164 10934 11376 10962
rect 11164 10656 11192 10934
rect 11436 10908 11744 10917
rect 11436 10906 11442 10908
rect 11498 10906 11522 10908
rect 11578 10906 11602 10908
rect 11658 10906 11682 10908
rect 11738 10906 11744 10908
rect 11498 10854 11500 10906
rect 11680 10854 11682 10906
rect 11436 10852 11442 10854
rect 11498 10852 11522 10854
rect 11578 10852 11602 10854
rect 11658 10852 11682 10854
rect 11738 10852 11744 10854
rect 11242 10840 11298 10849
rect 11436 10843 11744 10852
rect 11298 10810 11376 10826
rect 11298 10804 11388 10810
rect 11298 10798 11336 10804
rect 11242 10775 11298 10784
rect 11336 10746 11388 10752
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11520 10668 11572 10674
rect 11164 10628 11284 10656
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 8634 11192 9862
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 7342 11192 7822
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6866 11192 7142
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11256 6730 11284 10628
rect 11348 10628 11520 10656
rect 11348 9722 11376 10628
rect 11520 10610 11572 10616
rect 11716 10606 11744 10678
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11808 10520 11836 11630
rect 12084 11540 12112 12135
rect 12176 11801 12204 12294
rect 12348 12232 12400 12238
rect 12268 12192 12348 12220
rect 12162 11792 12218 11801
rect 12162 11727 12218 11736
rect 12268 11608 12296 12192
rect 12348 12174 12400 12180
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12348 11620 12400 11626
rect 12268 11580 12348 11608
rect 12348 11562 12400 11568
rect 11900 11512 12112 11540
rect 11900 11393 11928 11512
rect 12096 11452 12404 11461
rect 12096 11450 12102 11452
rect 12158 11450 12182 11452
rect 12238 11450 12262 11452
rect 12318 11450 12342 11452
rect 12398 11450 12404 11452
rect 12158 11398 12160 11450
rect 12340 11398 12342 11450
rect 12096 11396 12102 11398
rect 12158 11396 12182 11398
rect 12238 11396 12262 11398
rect 12318 11396 12342 11398
rect 12398 11396 12404 11398
rect 11886 11384 11942 11393
rect 12096 11387 12404 11396
rect 11886 11319 11942 11328
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 10532 11940 10538
rect 11808 10492 11888 10520
rect 11888 10474 11940 10480
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11612 10464 11664 10470
rect 11704 10464 11756 10470
rect 11612 10406 11664 10412
rect 11702 10432 11704 10441
rect 11756 10432 11758 10441
rect 11532 9926 11560 10406
rect 11624 10305 11652 10406
rect 11702 10367 11758 10376
rect 11610 10296 11666 10305
rect 11610 10231 11666 10240
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11436 9820 11744 9829
rect 11436 9818 11442 9820
rect 11498 9818 11522 9820
rect 11578 9818 11602 9820
rect 11658 9818 11682 9820
rect 11738 9818 11744 9820
rect 11498 9766 11500 9818
rect 11680 9766 11682 9818
rect 11436 9764 11442 9766
rect 11498 9764 11522 9766
rect 11578 9764 11602 9766
rect 11658 9764 11682 9766
rect 11738 9764 11744 9766
rect 11436 9755 11744 9764
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11440 9602 11468 9658
rect 11348 9574 11468 9602
rect 11348 8294 11376 9574
rect 11520 9512 11572 9518
rect 11518 9480 11520 9489
rect 11796 9512 11848 9518
rect 11572 9480 11574 9489
rect 11796 9454 11848 9460
rect 11518 9415 11574 9424
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11518 9208 11574 9217
rect 11716 9178 11744 9318
rect 11518 9143 11574 9152
rect 11704 9172 11756 9178
rect 11532 9110 11560 9143
rect 11704 9114 11756 9120
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11610 9072 11666 9081
rect 11610 9007 11612 9016
rect 11664 9007 11666 9016
rect 11612 8978 11664 8984
rect 11436 8732 11744 8741
rect 11436 8730 11442 8732
rect 11498 8730 11522 8732
rect 11578 8730 11602 8732
rect 11658 8730 11682 8732
rect 11738 8730 11744 8732
rect 11498 8678 11500 8730
rect 11680 8678 11682 8730
rect 11436 8676 11442 8678
rect 11498 8676 11522 8678
rect 11578 8676 11602 8678
rect 11658 8676 11682 8678
rect 11738 8676 11744 8678
rect 11436 8667 11744 8676
rect 11808 8634 11836 9454
rect 11900 9178 11928 9930
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11992 9058 12020 11154
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10713 12388 11086
rect 12346 10704 12402 10713
rect 12346 10639 12402 10648
rect 12162 10568 12218 10577
rect 12162 10503 12218 10512
rect 12176 10470 12204 10503
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12096 10364 12404 10373
rect 12096 10362 12102 10364
rect 12158 10362 12182 10364
rect 12238 10362 12262 10364
rect 12318 10362 12342 10364
rect 12398 10362 12404 10364
rect 12158 10310 12160 10362
rect 12340 10310 12342 10362
rect 12096 10308 12102 10310
rect 12158 10308 12182 10310
rect 12238 10308 12262 10310
rect 12318 10308 12342 10310
rect 12398 10308 12404 10310
rect 12096 10299 12404 10308
rect 12452 10266 12480 12038
rect 12544 11937 12572 12600
rect 12530 11928 12586 11937
rect 12530 11863 12586 11872
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12544 10674 12572 11766
rect 12636 11762 12664 12736
rect 12716 12718 12768 12724
rect 12820 12050 12848 13194
rect 12912 12714 12940 13382
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12912 12306 12940 12543
rect 13004 12442 13032 13330
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12728 12022 12848 12050
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12636 11218 12664 11698
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12636 10742 12664 11018
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12636 10198 12664 10406
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12360 9722 12388 9930
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 12084 9450 12112 9590
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12096 9276 12404 9285
rect 12096 9274 12102 9276
rect 12158 9274 12182 9276
rect 12238 9274 12262 9276
rect 12318 9274 12342 9276
rect 12398 9274 12404 9276
rect 12158 9222 12160 9274
rect 12340 9222 12342 9274
rect 12096 9220 12102 9222
rect 12158 9220 12182 9222
rect 12238 9220 12262 9222
rect 12318 9220 12342 9222
rect 12398 9220 12404 9222
rect 12096 9211 12404 9220
rect 11900 9030 12020 9058
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7954 11376 8230
rect 11440 8090 11468 8366
rect 11532 8294 11560 8570
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11436 7644 11744 7653
rect 11436 7642 11442 7644
rect 11498 7642 11522 7644
rect 11578 7642 11602 7644
rect 11658 7642 11682 7644
rect 11738 7642 11744 7644
rect 11498 7590 11500 7642
rect 11680 7590 11682 7642
rect 11436 7588 11442 7590
rect 11498 7588 11522 7590
rect 11578 7588 11602 7590
rect 11658 7588 11682 7590
rect 11738 7588 11744 7590
rect 11436 7579 11744 7588
rect 11808 7546 11836 8366
rect 11900 8129 11928 9030
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8809 12020 8910
rect 12452 8906 12480 9658
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12636 9353 12664 9454
rect 12622 9344 12678 9353
rect 12622 9279 12678 9288
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12348 8832 12400 8838
rect 11978 8800 12034 8809
rect 12348 8774 12400 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 11978 8735 12034 8744
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12268 8430 12296 8570
rect 12360 8537 12388 8774
rect 12346 8528 12402 8537
rect 12544 8498 12572 8774
rect 12346 8463 12402 8472
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12636 8430 12664 8910
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12624 8424 12676 8430
rect 12728 8412 12756 12022
rect 12806 11928 12862 11937
rect 12806 11863 12862 11872
rect 12820 8634 12848 11863
rect 12912 11121 12940 12106
rect 13004 11558 13032 12174
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11393 13032 11494
rect 12990 11384 13046 11393
rect 12990 11319 13046 11328
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12898 11112 12954 11121
rect 12898 11047 12954 11056
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10130 12940 10950
rect 13004 10470 13032 11154
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12990 10296 13046 10305
rect 12990 10231 13046 10240
rect 13004 10130 13032 10231
rect 13096 10198 13124 13262
rect 13280 12782 13308 13631
rect 13372 13530 13400 13670
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13464 13462 13492 14878
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14482 13584 14758
rect 13648 14521 13676 15302
rect 13728 14952 13780 14958
rect 13820 14952 13872 14958
rect 13728 14894 13780 14900
rect 13818 14920 13820 14929
rect 13872 14920 13874 14929
rect 13740 14618 13768 14894
rect 13818 14855 13874 14864
rect 13924 14618 13952 19654
rect 14108 19514 14136 20402
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14384 19394 14412 21383
rect 14462 20632 14518 20641
rect 14462 20567 14464 20576
rect 14516 20567 14518 20576
rect 14464 20538 14516 20544
rect 14200 19366 14412 19394
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14108 18834 14136 19246
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14016 17678 14044 18158
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14004 17536 14056 17542
rect 14002 17504 14004 17513
rect 14056 17504 14058 17513
rect 14002 17439 14058 17448
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13634 14512 13690 14521
rect 13544 14476 13596 14482
rect 13634 14447 13690 14456
rect 13544 14418 13596 14424
rect 13648 13977 13676 14447
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13634 13968 13690 13977
rect 13634 13903 13690 13912
rect 13832 13870 13860 14010
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13268 12776 13320 12782
rect 13174 12744 13230 12753
rect 13268 12718 13320 12724
rect 13174 12679 13230 12688
rect 13188 12306 13216 12679
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 11665 13216 12242
rect 13174 11656 13230 11665
rect 13174 11591 13230 11600
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 10742 13216 11494
rect 13280 11286 13308 12718
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13372 12442 13400 12650
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13372 10538 13400 11154
rect 13464 10606 13492 13398
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13556 12753 13584 13262
rect 13740 12986 13768 13262
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13832 12986 13860 13126
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13634 12880 13690 12889
rect 13634 12815 13636 12824
rect 13688 12815 13690 12824
rect 13636 12786 13688 12792
rect 13728 12776 13780 12782
rect 13542 12744 13598 12753
rect 13728 12718 13780 12724
rect 13542 12679 13598 12688
rect 13740 12306 13768 12718
rect 13924 12322 13952 13806
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13832 12294 13952 12322
rect 13544 12232 13596 12238
rect 13648 12209 13676 12242
rect 13544 12174 13596 12180
rect 13634 12200 13690 12209
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13266 10432 13322 10441
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12912 9042 12940 10066
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13004 9518 13032 9590
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 13004 8974 13032 9454
rect 13096 9217 13124 10134
rect 13188 10130 13216 10406
rect 13266 10367 13322 10376
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13176 9648 13228 9654
rect 13280 9636 13308 10367
rect 13228 9608 13308 9636
rect 13176 9590 13228 9596
rect 13372 9568 13400 10474
rect 13464 10130 13492 10542
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13280 9540 13400 9568
rect 13174 9344 13230 9353
rect 13174 9279 13230 9288
rect 13082 9208 13138 9217
rect 13082 9143 13138 9152
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12808 8424 12860 8430
rect 12728 8384 12808 8412
rect 12624 8366 12676 8372
rect 13096 8412 13124 9143
rect 13188 9110 13216 9279
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8430 13216 8774
rect 12808 8366 12860 8372
rect 12912 8384 13124 8412
rect 13176 8424 13228 8430
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11886 8120 11942 8129
rect 11886 8055 11942 8064
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11532 6798 11560 7482
rect 11900 7426 11928 8055
rect 11992 7721 12020 8298
rect 12360 8276 12388 8366
rect 12360 8248 12480 8276
rect 12096 8188 12404 8197
rect 12096 8186 12102 8188
rect 12158 8186 12182 8188
rect 12238 8186 12262 8188
rect 12318 8186 12342 8188
rect 12398 8186 12404 8188
rect 12158 8134 12160 8186
rect 12340 8134 12342 8186
rect 12096 8132 12102 8134
rect 12158 8132 12182 8134
rect 12238 8132 12262 8134
rect 12318 8132 12342 8134
rect 12398 8132 12404 8134
rect 12096 8123 12404 8132
rect 12452 8072 12480 8248
rect 12268 8044 12480 8072
rect 12164 7744 12216 7750
rect 11978 7712 12034 7721
rect 12164 7686 12216 7692
rect 11978 7647 12034 7656
rect 12176 7478 12204 7686
rect 12164 7472 12216 7478
rect 11900 7398 12112 7426
rect 12164 7414 12216 7420
rect 12084 7342 12112 7398
rect 12268 7392 12296 8044
rect 12636 8022 12664 8366
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12452 7449 12480 7890
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7750 12664 7822
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12438 7440 12494 7449
rect 12268 7364 12388 7392
rect 12438 7375 12494 7384
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6458 11100 6598
rect 11436 6556 11744 6565
rect 11436 6554 11442 6556
rect 11498 6554 11522 6556
rect 11578 6554 11602 6556
rect 11658 6554 11682 6556
rect 11738 6554 11744 6556
rect 11498 6502 11500 6554
rect 11680 6502 11682 6554
rect 11436 6500 11442 6502
rect 11498 6500 11522 6502
rect 11578 6500 11602 6502
rect 11658 6500 11682 6502
rect 11738 6500 11744 6502
rect 11436 6491 11744 6500
rect 11808 6458 11836 6802
rect 11992 6730 12020 7278
rect 12360 7188 12388 7364
rect 12532 7200 12584 7206
rect 12360 7160 12480 7188
rect 12096 7100 12404 7109
rect 12096 7098 12102 7100
rect 12158 7098 12182 7100
rect 12238 7098 12262 7100
rect 12318 7098 12342 7100
rect 12398 7098 12404 7100
rect 12158 7046 12160 7098
rect 12340 7046 12342 7098
rect 12096 7044 12102 7046
rect 12158 7044 12182 7046
rect 12238 7044 12262 7046
rect 12318 7044 12342 7046
rect 12398 7044 12404 7046
rect 12096 7035 12404 7044
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12452 6882 12480 7160
rect 12530 7168 12532 7177
rect 12584 7168 12586 7177
rect 12530 7103 12586 7112
rect 12636 7041 12664 7686
rect 12728 7274 12756 7686
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12820 7206 12848 8026
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12622 7032 12678 7041
rect 12622 6967 12678 6976
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11978 6624 12034 6633
rect 11978 6559 12034 6568
rect 11886 6488 11942 6497
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11796 6452 11848 6458
rect 11886 6423 11942 6432
rect 11796 6394 11848 6400
rect 11058 6352 11114 6361
rect 11058 6287 11114 6296
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10784 5704 10836 5710
rect 10968 5704 11020 5710
rect 10784 5646 10836 5652
rect 10874 5672 10930 5681
rect 10796 5574 10824 5646
rect 10968 5646 11020 5652
rect 10874 5607 10930 5616
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10048 3936 10100 3942
rect 10232 3936 10284 3942
rect 10100 3896 10232 3924
rect 10048 3878 10100 3884
rect 10232 3878 10284 3884
rect 10520 3398 10548 4014
rect 10612 3641 10640 4014
rect 10598 3632 10654 3641
rect 10598 3567 10654 3576
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 8850 2544 8906 2553
rect 8300 2508 8352 2514
rect 8850 2479 8906 2488
rect 8300 2450 8352 2456
rect 10888 2417 10916 5607
rect 10980 4690 11008 5646
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10968 4548 11020 4554
rect 11072 4536 11100 6287
rect 11164 6174 11468 6202
rect 11164 6118 11192 6174
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11164 5234 11192 5714
rect 11256 5302 11284 6054
rect 11334 5944 11390 5953
rect 11334 5879 11390 5888
rect 11348 5846 11376 5879
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11348 5166 11376 5782
rect 11440 5778 11468 6174
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5778 11560 6054
rect 11716 5778 11744 6394
rect 11796 6112 11848 6118
rect 11794 6080 11796 6089
rect 11848 6080 11850 6089
rect 11794 6015 11850 6024
rect 11900 5914 11928 6423
rect 11992 6254 12020 6559
rect 12268 6361 12296 6870
rect 12348 6860 12400 6866
rect 12452 6854 12572 6882
rect 12348 6802 12400 6808
rect 12254 6352 12310 6361
rect 12254 6287 12310 6296
rect 11980 6248 12032 6254
rect 12360 6236 12388 6802
rect 12440 6792 12492 6798
rect 12438 6760 12440 6769
rect 12492 6760 12494 6769
rect 12438 6695 12494 6704
rect 12360 6208 12480 6236
rect 11980 6190 12032 6196
rect 11992 5914 12020 6190
rect 12096 6012 12404 6021
rect 12096 6010 12102 6012
rect 12158 6010 12182 6012
rect 12238 6010 12262 6012
rect 12318 6010 12342 6012
rect 12398 6010 12404 6012
rect 12158 5958 12160 6010
rect 12340 5958 12342 6010
rect 12096 5956 12102 5958
rect 12158 5956 12182 5958
rect 12238 5956 12262 5958
rect 12318 5956 12342 5958
rect 12398 5956 12404 5958
rect 12096 5947 12404 5956
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12452 5846 12480 6208
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 12084 5710 12112 5782
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11436 5468 11744 5477
rect 11436 5466 11442 5468
rect 11498 5466 11522 5468
rect 11578 5466 11602 5468
rect 11658 5466 11682 5468
rect 11738 5466 11744 5468
rect 11498 5414 11500 5466
rect 11680 5414 11682 5466
rect 11436 5412 11442 5414
rect 11498 5412 11522 5414
rect 11578 5412 11602 5414
rect 11658 5412 11682 5414
rect 11738 5412 11744 5414
rect 11436 5403 11744 5412
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11716 5166 11744 5238
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11716 5030 11744 5102
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11164 4622 11192 4966
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11020 4508 11100 4536
rect 10968 4490 11020 4496
rect 11072 4078 11100 4508
rect 11348 4146 11376 4966
rect 11808 4486 11836 5578
rect 12348 5568 12400 5574
rect 11900 5516 12348 5522
rect 11900 5510 12400 5516
rect 11900 5494 12388 5510
rect 11900 5030 11928 5494
rect 12544 5370 12572 6854
rect 12820 6746 12848 7142
rect 12912 7002 12940 8384
rect 13176 8366 13228 8372
rect 13188 8294 13216 8366
rect 13096 8266 13216 8294
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13004 7002 13032 7278
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 12992 6860 13044 6866
rect 12728 6718 12848 6746
rect 12912 6820 12992 6848
rect 12728 6186 12756 6718
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6322 12848 6598
rect 12912 6322 12940 6820
rect 12992 6802 13044 6808
rect 13096 6798 13124 8266
rect 13280 8090 13308 9540
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 8537 13400 9386
rect 13358 8528 13414 8537
rect 13358 8463 13414 8472
rect 13464 8362 13492 10066
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7206 13216 7754
rect 13280 7342 13308 7890
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13084 6792 13136 6798
rect 12990 6760 13046 6769
rect 13084 6734 13136 6740
rect 12990 6695 13046 6704
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12716 6180 12768 6186
rect 12768 6140 12848 6168
rect 12716 6122 12768 6128
rect 12714 5536 12770 5545
rect 12714 5471 12770 5480
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 12096 4924 12404 4933
rect 12096 4922 12102 4924
rect 12158 4922 12182 4924
rect 12238 4922 12262 4924
rect 12318 4922 12342 4924
rect 12398 4922 12404 4924
rect 12158 4870 12160 4922
rect 12340 4870 12342 4922
rect 12096 4868 12102 4870
rect 12158 4868 12182 4870
rect 12238 4868 12262 4870
rect 12318 4868 12342 4870
rect 12398 4868 12404 4870
rect 12096 4859 12404 4868
rect 11978 4720 12034 4729
rect 11978 4655 12034 4664
rect 11992 4622 12020 4655
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11796 4480 11848 4486
rect 11796 4422 11848 4428
rect 11436 4380 11744 4389
rect 11436 4378 11442 4380
rect 11498 4378 11522 4380
rect 11578 4378 11602 4380
rect 11658 4378 11682 4380
rect 11738 4378 11744 4380
rect 11498 4326 11500 4378
rect 11680 4326 11682 4378
rect 11436 4324 11442 4326
rect 11498 4324 11522 4326
rect 11578 4324 11602 4326
rect 11658 4324 11682 4326
rect 11738 4324 11744 4326
rect 11436 4315 11744 4324
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11610 4040 11666 4049
rect 11610 3975 11666 3984
rect 11624 3942 11652 3975
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11436 3292 11744 3301
rect 11436 3290 11442 3292
rect 11498 3290 11522 3292
rect 11578 3290 11602 3292
rect 11658 3290 11682 3292
rect 11738 3290 11744 3292
rect 11498 3238 11500 3290
rect 11680 3238 11682 3290
rect 11436 3236 11442 3238
rect 11498 3236 11522 3238
rect 11578 3236 11602 3238
rect 11658 3236 11682 3238
rect 11738 3236 11744 3238
rect 11436 3227 11744 3236
rect 11900 2446 11928 4558
rect 11992 4457 12020 4558
rect 11978 4448 12034 4457
rect 11978 4383 12034 4392
rect 12452 4078 12480 5306
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12544 4826 12572 5170
rect 12728 5166 12756 5471
rect 12716 5160 12768 5166
rect 12714 5128 12716 5137
rect 12768 5128 12770 5137
rect 12714 5063 12770 5072
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12096 3836 12404 3845
rect 12096 3834 12102 3836
rect 12158 3834 12182 3836
rect 12238 3834 12262 3836
rect 12318 3834 12342 3836
rect 12398 3834 12404 3836
rect 12158 3782 12160 3834
rect 12340 3782 12342 3834
rect 12096 3780 12102 3782
rect 12158 3780 12182 3782
rect 12238 3780 12262 3782
rect 12318 3780 12342 3782
rect 12398 3780 12404 3782
rect 12096 3771 12404 3780
rect 12348 3460 12400 3466
rect 12544 3448 12572 4626
rect 12622 4584 12678 4593
rect 12820 4554 12848 6140
rect 12912 5370 12940 6258
rect 13004 6254 13032 6695
rect 13096 6254 13124 6734
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13004 5817 13032 6054
rect 12990 5808 13046 5817
rect 12990 5743 13046 5752
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12912 5030 12940 5170
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12622 4519 12678 4528
rect 12808 4548 12860 4554
rect 12636 4282 12664 4519
rect 12808 4490 12860 4496
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12912 4214 12940 4966
rect 13096 4826 13124 6190
rect 13188 5234 13216 7142
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13280 6118 13308 6802
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13280 5846 13308 6054
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 13096 4060 13124 4762
rect 13372 4622 13400 8298
rect 13450 8120 13506 8129
rect 13450 8055 13506 8064
rect 13464 7750 13492 8055
rect 13556 7886 13584 12174
rect 13634 12135 13690 12144
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13648 11150 13676 11562
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 11218 13768 11290
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13636 11144 13688 11150
rect 13832 11098 13860 12294
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 11121 13952 12174
rect 13636 11086 13688 11092
rect 13648 9489 13676 11086
rect 13740 11070 13860 11098
rect 13910 11112 13966 11121
rect 13740 9926 13768 11070
rect 13910 11047 13966 11056
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10606 13952 10950
rect 14016 10674 14044 15846
rect 14108 15337 14136 18226
rect 14200 17746 14228 19366
rect 14370 19272 14426 19281
rect 14370 19207 14426 19216
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14292 18086 14320 18770
rect 14384 18358 14412 19207
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14384 18222 14412 18294
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14292 17649 14320 17682
rect 14278 17640 14334 17649
rect 14188 17604 14240 17610
rect 14278 17575 14334 17584
rect 14188 17546 14240 17552
rect 14200 17270 14228 17546
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14292 16454 14320 17070
rect 14384 16590 14412 17070
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14476 16250 14504 18702
rect 14568 18465 14596 18702
rect 14554 18456 14610 18465
rect 14554 18391 14610 18400
rect 14660 18290 14688 21490
rect 14752 21418 14780 21490
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 14740 21412 14792 21418
rect 14740 21354 14792 21360
rect 14752 21078 14780 21354
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 14740 21072 14792 21078
rect 14740 21014 14792 21020
rect 15474 21040 15530 21049
rect 14752 20398 14780 21014
rect 15384 21004 15436 21010
rect 16132 21010 16160 21286
rect 15474 20975 15530 20984
rect 16028 21004 16080 21010
rect 15384 20946 15436 20952
rect 15396 20874 15424 20946
rect 15488 20942 15516 20975
rect 16028 20946 16080 20952
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20641 15240 20742
rect 15198 20632 15254 20641
rect 15198 20567 15254 20576
rect 14830 20496 14886 20505
rect 14830 20431 14886 20440
rect 15384 20460 15436 20466
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14752 19922 14780 20198
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14752 19378 14780 19858
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18465 14780 18566
rect 14738 18456 14794 18465
rect 14738 18391 14794 18400
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14568 17134 14596 17274
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14554 16824 14610 16833
rect 14554 16759 14610 16768
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14292 16153 14320 16186
rect 14278 16144 14334 16153
rect 14278 16079 14334 16088
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14186 15872 14242 15881
rect 14186 15807 14242 15816
rect 14094 15328 14150 15337
rect 14094 15263 14150 15272
rect 14200 15162 14228 15807
rect 14292 15162 14320 15982
rect 14568 15638 14596 16759
rect 14660 16522 14688 17682
rect 14752 17542 14780 18391
rect 14844 17864 14872 20431
rect 15384 20402 15436 20408
rect 15396 19961 15424 20402
rect 15568 19984 15620 19990
rect 15014 19952 15070 19961
rect 15014 19887 15016 19896
rect 15068 19887 15070 19896
rect 15382 19952 15438 19961
rect 15568 19926 15620 19932
rect 15382 19887 15438 19896
rect 15016 19858 15068 19864
rect 15580 19242 15608 19926
rect 16040 19718 16068 20946
rect 16408 20890 16436 21422
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16486 21176 16542 21185
rect 16776 21146 16804 21354
rect 16486 21111 16542 21120
rect 16764 21140 16816 21146
rect 16500 21078 16528 21111
rect 16764 21082 16816 21088
rect 17236 21078 17264 21490
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 17328 21146 17356 21286
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 16488 21072 16540 21078
rect 16488 21014 16540 21020
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 17040 20936 17092 20942
rect 16408 20874 16528 20890
rect 17040 20878 17092 20884
rect 16408 20868 16540 20874
rect 16408 20862 16488 20868
rect 16488 20810 16540 20816
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 16132 19854 16160 20266
rect 16408 20074 16436 20538
rect 16500 20466 16528 20810
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16776 20466 16804 20742
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16224 20046 16436 20074
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15764 19553 15792 19654
rect 15750 19544 15806 19553
rect 15750 19479 15806 19488
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15120 19009 15148 19110
rect 15106 19000 15162 19009
rect 15106 18935 15162 18944
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14936 18290 14964 18566
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14844 17836 14964 17864
rect 14830 17776 14886 17785
rect 14830 17711 14886 17720
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14660 15201 14688 15574
rect 14646 15192 14702 15201
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14280 15156 14332 15162
rect 14646 15127 14702 15136
rect 14280 15098 14332 15104
rect 14372 15088 14424 15094
rect 14200 15036 14372 15042
rect 14200 15030 14424 15036
rect 14200 15014 14412 15030
rect 14648 15020 14700 15026
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14108 14482 14136 14894
rect 14200 14822 14228 15014
rect 14648 14962 14700 14968
rect 14660 14890 14688 14962
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14108 13938 14136 14010
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14108 13190 14136 13738
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14094 12744 14150 12753
rect 14094 12679 14150 12688
rect 14108 12374 14136 12679
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13832 9722 13860 10066
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13924 9654 13952 9998
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13728 9512 13780 9518
rect 13634 9480 13690 9489
rect 13728 9454 13780 9460
rect 13634 9415 13690 9424
rect 13740 9081 13768 9454
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13726 9072 13782 9081
rect 13924 9042 13952 9114
rect 14016 9081 14044 10202
rect 14002 9072 14058 9081
rect 13726 9007 13782 9016
rect 13912 9036 13964 9042
rect 14002 9007 14058 9016
rect 13912 8978 13964 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13910 8936 13966 8945
rect 13648 8090 13676 8910
rect 13728 8900 13780 8906
rect 13910 8871 13966 8880
rect 13728 8842 13780 8848
rect 13740 8566 13768 8842
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13740 8430 13768 8502
rect 13924 8430 13952 8871
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13556 7449 13584 7822
rect 13542 7440 13598 7449
rect 13542 7375 13598 7384
rect 13740 6934 13768 8230
rect 13832 7721 13860 8230
rect 14016 7954 14044 9007
rect 14108 7954 14136 12310
rect 14200 12238 14228 14758
rect 14292 14550 14320 14758
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14292 13258 14320 13398
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 12782 14320 13194
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14188 12232 14240 12238
rect 14186 12200 14188 12209
rect 14280 12232 14332 12238
rect 14240 12200 14242 12209
rect 14280 12174 14332 12180
rect 14186 12135 14242 12144
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11778 14228 12038
rect 14292 11898 14320 12174
rect 14384 11898 14412 12242
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14200 11750 14320 11778
rect 14188 11552 14240 11558
rect 14292 11529 14320 11750
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14188 11494 14240 11500
rect 14278 11520 14334 11529
rect 14200 11218 14228 11494
rect 14278 11455 14334 11464
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14200 10713 14228 11018
rect 14186 10704 14242 10713
rect 14186 10639 14242 10648
rect 14200 10606 14228 10639
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14292 9976 14320 11455
rect 14476 11354 14504 11630
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14370 11248 14426 11257
rect 14370 11183 14372 11192
rect 14424 11183 14426 11192
rect 14372 11154 14424 11160
rect 14200 9948 14320 9976
rect 14200 9654 14228 9948
rect 14278 9888 14334 9897
rect 14278 9823 14334 9832
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14200 8945 14228 9386
rect 14292 9042 14320 9823
rect 14384 9738 14412 11154
rect 14462 10704 14518 10713
rect 14462 10639 14518 10648
rect 14476 10606 14504 10639
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14476 10044 14504 10367
rect 14568 10146 14596 13806
rect 14660 13394 14688 14486
rect 14752 13870 14780 17478
rect 14844 17202 14872 17711
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14936 16726 14964 17836
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14924 16720 14976 16726
rect 15028 16697 15056 17070
rect 15396 17066 15424 18362
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 14924 16662 14976 16668
rect 15014 16688 15070 16697
rect 15014 16623 15070 16632
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 14830 16008 14886 16017
rect 14830 15943 14886 15952
rect 14844 15570 14872 15943
rect 15028 15638 15056 16186
rect 15016 15632 15068 15638
rect 14936 15592 15016 15620
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14936 14890 14964 15592
rect 15016 15574 15068 15580
rect 15120 15337 15148 17002
rect 15396 15910 15424 17002
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15106 15328 15162 15337
rect 15106 15263 15162 15272
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14844 14385 14872 14554
rect 15028 14482 15056 15098
rect 15212 15094 15240 15642
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15108 14884 15160 14890
rect 15212 14872 15240 15030
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15160 14844 15240 14872
rect 15108 14826 15160 14832
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14830 14376 14886 14385
rect 14830 14311 14886 14320
rect 14830 14104 14886 14113
rect 14936 14074 14964 14418
rect 15120 14385 15148 14826
rect 15304 14618 15332 14962
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15106 14376 15162 14385
rect 15106 14311 15162 14320
rect 15290 14376 15346 14385
rect 15290 14311 15346 14320
rect 15014 14104 15070 14113
rect 14830 14039 14886 14048
rect 14924 14068 14976 14074
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14738 13560 14794 13569
rect 14738 13495 14794 13504
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14752 13326 14780 13495
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14844 12696 14872 14039
rect 15014 14039 15070 14048
rect 14924 14010 14976 14016
rect 14844 12668 14964 12696
rect 14830 12608 14886 12617
rect 14830 12543 14886 12552
rect 14738 12336 14794 12345
rect 14738 12271 14740 12280
rect 14792 12271 14794 12280
rect 14740 12242 14792 12248
rect 14844 11694 14872 12543
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 11354 14688 11562
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14738 11248 14794 11257
rect 14738 11183 14794 11192
rect 14752 10606 14780 11183
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14844 10266 14872 11630
rect 14936 11286 14964 12668
rect 15028 12442 15056 14039
rect 15108 14000 15160 14006
rect 15106 13968 15108 13977
rect 15160 13968 15162 13977
rect 15106 13903 15162 13912
rect 15120 13870 15148 13903
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 12782 15148 13330
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 11801 15148 12038
rect 15212 11898 15240 13738
rect 15304 13705 15332 14311
rect 15396 13870 15424 15302
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15290 13696 15346 13705
rect 15290 13631 15346 13640
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15304 13258 15332 13330
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15304 12345 15332 12718
rect 15290 12336 15346 12345
rect 15290 12271 15346 12280
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14924 11280 14976 11286
rect 14922 11248 14924 11257
rect 15120 11257 15148 11630
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14976 11248 14978 11257
rect 14922 11183 14978 11192
rect 15106 11248 15162 11257
rect 15106 11183 15162 11192
rect 14936 10266 14964 11183
rect 15212 10985 15240 11494
rect 15396 11218 15424 13806
rect 15488 13530 15516 17614
rect 15580 17338 15608 17614
rect 15764 17542 15792 18702
rect 16224 18630 16252 20046
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16316 18902 16344 19926
rect 16408 19854 16436 20046
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16408 19310 16436 19654
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16316 18290 16344 18838
rect 16500 18766 16528 20402
rect 17052 20058 17080 20878
rect 17236 20330 17264 21014
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17958 20632 18014 20641
rect 17958 20567 17960 20576
rect 18012 20567 18014 20576
rect 17960 20538 18012 20544
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17958 20224 18014 20233
rect 17958 20159 18014 20168
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16592 19514 16620 19790
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16684 19394 16712 19790
rect 17144 19700 17172 19994
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 16868 19672 17172 19700
rect 16868 19553 16896 19672
rect 16854 19544 16910 19553
rect 17512 19514 17540 19858
rect 16854 19479 16910 19488
rect 17132 19508 17184 19514
rect 16592 19366 16712 19394
rect 16592 18834 16620 19366
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16684 18970 16712 19246
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16408 18222 16436 18634
rect 16592 18630 16620 18770
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16776 18426 16804 18770
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 15856 17678 15884 18022
rect 15844 17672 15896 17678
rect 15842 17640 15844 17649
rect 15896 17640 15898 17649
rect 15842 17575 15898 17584
rect 16212 17604 16264 17610
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 16114 15700 16458
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15570 15608 15846
rect 15658 15736 15714 15745
rect 15764 15706 15792 17070
rect 15658 15671 15714 15680
rect 15752 15700 15804 15706
rect 15672 15570 15700 15671
rect 15752 15642 15804 15648
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15752 15564 15804 15570
rect 15856 15552 15884 17575
rect 16212 17546 16264 17552
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16132 16794 16160 17070
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16028 16720 16080 16726
rect 16026 16688 16028 16697
rect 16080 16688 16082 16697
rect 15936 16652 15988 16658
rect 16026 16623 16082 16632
rect 15936 16594 15988 16600
rect 15948 16561 15976 16594
rect 16028 16584 16080 16590
rect 15934 16552 15990 16561
rect 16028 16526 16080 16532
rect 15934 16487 15990 16496
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 16114 15976 16390
rect 16040 16182 16068 16526
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 15620 15976 16050
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 15948 15592 16068 15620
rect 15856 15524 15976 15552
rect 15752 15506 15804 15512
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12782 15516 13262
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 12170 15516 12718
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15198 10976 15254 10985
rect 15198 10911 15254 10920
rect 15396 10742 15424 11018
rect 15292 10736 15344 10742
rect 15014 10704 15070 10713
rect 15198 10704 15254 10713
rect 15292 10678 15344 10684
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15014 10639 15070 10648
rect 15120 10648 15198 10656
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14740 10192 14792 10198
rect 14738 10160 14740 10169
rect 14792 10160 14794 10169
rect 14568 10118 14688 10146
rect 14556 10056 14608 10062
rect 14476 10016 14556 10044
rect 14556 9998 14608 10004
rect 14384 9710 14504 9738
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14186 8936 14242 8945
rect 14186 8871 14242 8880
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14200 8498 14228 8570
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14186 8392 14242 8401
rect 14384 8378 14412 9590
rect 14476 9382 14504 9710
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14568 9450 14596 9590
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 8514 14504 9318
rect 14660 9092 14688 10118
rect 14738 10095 14794 10104
rect 15028 10062 15056 10639
rect 15120 10628 15200 10648
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14740 9920 14792 9926
rect 15120 9874 15148 10628
rect 15252 10639 15254 10648
rect 15200 10610 15252 10616
rect 15304 10538 15332 10678
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 14740 9862 14792 9868
rect 14568 9064 14688 9092
rect 14568 8616 14596 9064
rect 14568 8588 14688 8616
rect 14476 8486 14596 8514
rect 14186 8327 14242 8336
rect 14292 8350 14412 8378
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14200 7954 14228 8327
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14096 7948 14148 7954
rect 14096 7890 14148 7896
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13818 7712 13874 7721
rect 13818 7647 13874 7656
rect 13832 7018 13860 7647
rect 13924 7177 13952 7822
rect 14096 7744 14148 7750
rect 14094 7712 14096 7721
rect 14148 7712 14150 7721
rect 14094 7647 14150 7656
rect 13910 7168 13966 7177
rect 13910 7103 13966 7112
rect 13832 6990 13952 7018
rect 13452 6928 13504 6934
rect 13728 6928 13780 6934
rect 13452 6870 13504 6876
rect 13542 6896 13598 6905
rect 13464 6254 13492 6870
rect 13728 6870 13780 6876
rect 13542 6831 13598 6840
rect 13556 6798 13584 6831
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13556 5914 13584 6734
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13740 6118 13768 6326
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13924 5914 13952 6990
rect 14200 6746 14228 7890
rect 14016 6718 14228 6746
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13464 5534 13492 5850
rect 13740 5556 13768 5850
rect 13464 5506 13676 5534
rect 13740 5528 13860 5556
rect 13648 5166 13676 5506
rect 13832 5522 13860 5528
rect 13832 5494 13952 5522
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13176 4072 13228 4078
rect 13096 4032 13176 4060
rect 13176 4014 13228 4020
rect 13464 3913 13492 4082
rect 13924 4078 13952 5494
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 14016 3924 14044 6718
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6254 14136 6598
rect 14292 6254 14320 8350
rect 14476 8129 14504 8366
rect 14568 8362 14596 8486
rect 14660 8430 14688 8588
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14462 8120 14518 8129
rect 14660 8090 14688 8366
rect 14752 8294 14780 9862
rect 14844 9846 15148 9874
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14462 8055 14518 8064
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14738 7984 14794 7993
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14464 7948 14516 7954
rect 14516 7908 14688 7936
rect 14738 7919 14740 7928
rect 14464 7890 14516 7896
rect 14384 7818 14412 7890
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14568 7342 14596 7482
rect 14660 7342 14688 7908
rect 14792 7919 14794 7928
rect 14740 7890 14792 7896
rect 14752 7410 14780 7890
rect 14844 7886 14872 9846
rect 15304 9738 15332 9930
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15120 9710 15332 9738
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15028 9042 15056 9590
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 8294 14964 8842
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 15028 8566 15056 8599
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 15014 8392 15070 8401
rect 15014 8327 15016 8336
rect 15068 8327 15070 8336
rect 15016 8298 15068 8304
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 15014 8256 15070 8265
rect 15120 8242 15148 9710
rect 15396 9674 15424 9862
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15304 9646 15424 9674
rect 15212 9518 15240 9590
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15070 8214 15148 8242
rect 15014 8191 15070 8200
rect 14924 7948 14976 7954
rect 15028 7936 15056 8191
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 14976 7908 15056 7936
rect 14924 7890 14976 7896
rect 14832 7880 14884 7886
rect 14884 7828 15056 7834
rect 14832 7822 15056 7828
rect 14844 7806 15056 7822
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14922 7712 14978 7721
rect 14844 7546 14872 7686
rect 14922 7647 14978 7656
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14936 7342 14964 7647
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14660 7002 14688 7278
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14476 5953 14504 6938
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14462 5944 14518 5953
rect 14462 5879 14518 5888
rect 14568 5642 14596 6802
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14200 4146 14228 5102
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13450 3904 13506 3913
rect 13450 3839 13506 3848
rect 13924 3896 14044 3924
rect 12898 3768 12954 3777
rect 12898 3703 12954 3712
rect 12912 3602 12940 3703
rect 13818 3632 13874 3641
rect 12900 3596 12952 3602
rect 13924 3618 13952 3896
rect 14292 3777 14320 4966
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14278 3768 14334 3777
rect 14278 3703 14334 3712
rect 13874 3602 13952 3618
rect 14002 3632 14058 3641
rect 13874 3596 13964 3602
rect 13874 3590 13912 3596
rect 13818 3567 13874 3576
rect 12900 3538 12952 3544
rect 14292 3602 14320 3703
rect 14476 3670 14504 3946
rect 14660 3738 14688 6190
rect 14752 6089 14780 6190
rect 14738 6080 14794 6089
rect 14738 6015 14794 6024
rect 14844 5522 14872 6258
rect 15028 6254 15056 7806
rect 15120 7721 15148 8026
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15108 6792 15160 6798
rect 15106 6760 15108 6769
rect 15160 6760 15162 6769
rect 15106 6695 15162 6704
rect 15212 6254 15240 9454
rect 15304 9450 15332 9646
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15396 9330 15424 9522
rect 15304 9302 15424 9330
rect 15304 8820 15332 9302
rect 15382 9208 15438 9217
rect 15382 9143 15438 9152
rect 15396 8974 15424 9143
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15384 8832 15436 8838
rect 15304 8792 15384 8820
rect 15384 8774 15436 8780
rect 15382 8664 15438 8673
rect 15382 8599 15384 8608
rect 15436 8599 15438 8608
rect 15384 8570 15436 8576
rect 15292 8084 15344 8090
rect 15384 8084 15436 8090
rect 15344 8044 15384 8072
rect 15292 8026 15344 8032
rect 15384 8026 15436 8032
rect 15304 7546 15332 8026
rect 15384 7982 15436 7988
rect 15384 7924 15436 7930
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15396 7426 15424 7924
rect 15488 7546 15516 11834
rect 15580 11626 15608 15506
rect 15764 15366 15792 15506
rect 15842 15464 15898 15473
rect 15842 15399 15898 15408
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15672 14482 15700 14894
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 14278 15700 14418
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 12918 15700 13670
rect 15764 13394 15792 14962
rect 15856 13569 15884 15399
rect 15948 13938 15976 15524
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15842 13560 15898 13569
rect 15842 13495 15898 13504
rect 15856 13394 15884 13495
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15660 12776 15712 12782
rect 15658 12744 15660 12753
rect 15712 12744 15714 12753
rect 15658 12679 15714 12688
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 11082 15608 11154
rect 15672 11082 15700 12174
rect 15764 11898 15792 13330
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15750 11792 15806 11801
rect 15750 11727 15806 11736
rect 15764 11694 15792 11727
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15566 10840 15622 10849
rect 15566 10775 15622 10784
rect 15580 10742 15608 10775
rect 15568 10736 15620 10742
rect 15620 10696 15700 10724
rect 15568 10678 15620 10684
rect 15566 9344 15622 9353
rect 15566 9279 15622 9288
rect 15580 8673 15608 9279
rect 15566 8664 15622 8673
rect 15566 8599 15622 8608
rect 15672 8480 15700 10696
rect 15856 10690 15884 12786
rect 15948 12646 15976 13398
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11937 15976 12174
rect 15934 11928 15990 11937
rect 15934 11863 15990 11872
rect 16040 11626 16068 15592
rect 16132 13274 16160 15914
rect 16224 15026 16252 17546
rect 16316 17202 16344 18022
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16316 14482 16344 17138
rect 16408 16697 16436 17750
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16592 17134 16620 17682
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16776 17202 16804 17478
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16394 16688 16450 16697
rect 16394 16623 16396 16632
rect 16448 16623 16450 16632
rect 16396 16594 16448 16600
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 16017 16436 16390
rect 16488 16040 16540 16046
rect 16394 16008 16450 16017
rect 16488 15982 16540 15988
rect 16394 15943 16450 15952
rect 16500 15706 16528 15982
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16408 14618 16436 15370
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 14074 16252 14350
rect 16212 14068 16264 14074
rect 16500 14056 16528 15642
rect 16592 14482 16620 17070
rect 16868 17066 16896 19479
rect 17132 19450 17184 19456
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17144 18902 17172 19450
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17236 18222 17264 18362
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17604 18154 17632 19246
rect 17880 18426 17908 19858
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17224 17808 17276 17814
rect 17276 17768 17540 17796
rect 17224 17750 17276 17756
rect 17052 17105 17080 17750
rect 17130 17504 17186 17513
rect 17130 17439 17186 17448
rect 17038 17096 17094 17105
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16856 17060 16908 17066
rect 17038 17031 17094 17040
rect 16856 17002 16908 17008
rect 16776 16794 16804 17002
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 16289 16712 16594
rect 16670 16280 16726 16289
rect 16670 16215 16726 16224
rect 16684 15609 16712 16215
rect 16670 15600 16726 15609
rect 16670 15535 16726 15544
rect 16764 15496 16816 15502
rect 16762 15464 16764 15473
rect 16816 15464 16818 15473
rect 16762 15399 16818 15408
rect 16764 14816 16816 14822
rect 16868 14804 16896 17002
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 15570 16988 16934
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17052 15978 17080 16594
rect 17144 16522 17172 17439
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 17144 15858 17172 16458
rect 17052 15830 17172 15858
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16946 15192 17002 15201
rect 16946 15127 17002 15136
rect 16960 15026 16988 15127
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16960 14929 16988 14962
rect 16946 14920 17002 14929
rect 16946 14855 17002 14864
rect 16816 14776 16896 14804
rect 16764 14758 16816 14764
rect 16580 14476 16632 14482
rect 16764 14476 16816 14482
rect 16632 14436 16712 14464
rect 16580 14418 16632 14424
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16212 14010 16264 14016
rect 16408 14028 16528 14056
rect 16302 13832 16358 13841
rect 16302 13767 16358 13776
rect 16210 13424 16266 13433
rect 16210 13359 16212 13368
rect 16264 13359 16266 13368
rect 16212 13330 16264 13336
rect 16132 13246 16252 13274
rect 16118 12744 16174 12753
rect 16118 12679 16174 12688
rect 16132 12073 16160 12679
rect 16118 12064 16174 12073
rect 16118 11999 16174 12008
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16132 11150 16160 11999
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15764 10662 15884 10690
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15764 10441 15792 10662
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15750 10432 15806 10441
rect 15750 10367 15806 10376
rect 15856 10198 15884 10542
rect 15948 10282 15976 10678
rect 16040 10538 16068 11086
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15948 10254 16068 10282
rect 16040 10198 16068 10254
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16026 9888 16082 9897
rect 16026 9823 16082 9832
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15856 9382 15884 9590
rect 16040 9489 16068 9823
rect 16026 9480 16082 9489
rect 16026 9415 16082 9424
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15934 9344 15990 9353
rect 15934 9279 15990 9288
rect 15948 9024 15976 9279
rect 15856 8996 15976 9024
rect 15672 8452 15792 8480
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15566 8256 15622 8265
rect 15566 8191 15622 8200
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15304 7398 15424 7426
rect 15304 7342 15332 7398
rect 15292 7336 15344 7342
rect 15476 7336 15528 7342
rect 15292 7278 15344 7284
rect 15384 7302 15436 7308
rect 15580 7324 15608 8191
rect 15672 7342 15700 8298
rect 15528 7296 15608 7324
rect 15660 7336 15712 7342
rect 15476 7278 15528 7284
rect 15660 7278 15712 7284
rect 15384 7244 15436 7250
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15304 6458 15332 6734
rect 15396 6458 15424 7244
rect 15474 7032 15530 7041
rect 15474 6967 15476 6976
rect 15528 6967 15530 6976
rect 15476 6938 15528 6944
rect 15672 6662 15700 7278
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15384 6180 15436 6186
rect 15384 6122 15436 6128
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 14752 5494 14872 5522
rect 14752 5166 14780 5494
rect 14922 5400 14978 5409
rect 14832 5364 14884 5370
rect 14922 5335 14978 5344
rect 15106 5400 15162 5409
rect 15106 5335 15162 5344
rect 14832 5306 14884 5312
rect 14844 5166 14872 5306
rect 14936 5302 14964 5335
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14832 5160 14884 5166
rect 14936 5137 14964 5238
rect 15120 5234 15148 5335
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15304 5166 15332 5850
rect 15396 5846 15424 6122
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15672 5642 15700 6598
rect 15764 5710 15792 8452
rect 15856 8090 15884 8996
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15842 7712 15898 7721
rect 15842 7647 15898 7656
rect 15856 7410 15884 7647
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15292 5160 15344 5166
rect 14832 5102 14884 5108
rect 14922 5128 14978 5137
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14464 3664 14516 3670
rect 14370 3632 14426 3641
rect 14002 3567 14058 3576
rect 14280 3596 14332 3602
rect 13912 3538 13964 3544
rect 12912 3466 12940 3538
rect 14016 3534 14044 3567
rect 14464 3606 14516 3612
rect 14370 3567 14372 3576
rect 14280 3538 14332 3544
rect 14424 3567 14426 3576
rect 14372 3538 14424 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14476 3466 14504 3606
rect 12400 3420 12572 3448
rect 12900 3460 12952 3466
rect 12348 3402 12400 3408
rect 12900 3402 12952 3408
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14752 3398 14780 5102
rect 14844 4078 14872 5102
rect 15292 5102 15344 5108
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14922 5063 14978 5072
rect 15304 4078 15332 5102
rect 15396 4826 15424 5102
rect 15660 5092 15712 5098
rect 15488 5052 15660 5080
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15396 4486 15424 4762
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15488 4078 15516 5052
rect 15660 5034 15712 5040
rect 15764 5030 15792 5646
rect 15948 5302 15976 8842
rect 16040 7721 16068 9415
rect 16026 7712 16082 7721
rect 16026 7647 16082 7656
rect 16132 6934 16160 11086
rect 16120 6928 16172 6934
rect 16118 6896 16120 6905
rect 16172 6896 16174 6905
rect 16118 6831 16174 6840
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16132 6458 16160 6734
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 16026 5264 16082 5273
rect 16026 5199 16082 5208
rect 16040 5166 16068 5199
rect 16132 5166 16160 6190
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15750 4856 15806 4865
rect 15750 4791 15806 4800
rect 15764 4690 15792 4791
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15764 4154 15792 4626
rect 15764 4126 15976 4154
rect 15948 4078 15976 4126
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15488 3398 15516 4014
rect 16132 4010 16160 5102
rect 16224 4622 16252 13246
rect 16316 13190 16344 13767
rect 16408 13274 16436 14028
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16500 13705 16528 13874
rect 16486 13696 16542 13705
rect 16486 13631 16542 13640
rect 16408 13246 16528 13274
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12986 16436 13126
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16500 12434 16528 13246
rect 16592 12628 16620 14282
rect 16684 13938 16712 14436
rect 16764 14418 16816 14424
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16776 12986 16804 14418
rect 16868 14346 16896 14776
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16856 14340 16908 14346
rect 16856 14282 16908 14288
rect 16960 14113 16988 14418
rect 16946 14104 17002 14113
rect 16946 14039 17002 14048
rect 17052 13988 17080 15830
rect 17236 14958 17264 17274
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17224 14952 17276 14958
rect 17144 14912 17224 14940
rect 17144 14550 17172 14912
rect 17224 14894 17276 14900
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17236 14006 17264 14758
rect 17328 14006 17356 15438
rect 17420 15026 17448 17070
rect 17512 17066 17540 17768
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17498 16688 17554 16697
rect 17498 16623 17500 16632
rect 17552 16623 17554 16632
rect 17500 16594 17552 16600
rect 17498 16416 17554 16425
rect 17498 16351 17554 16360
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17512 14414 17540 16351
rect 17604 14958 17632 18090
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17696 17746 17724 17818
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17696 17610 17724 17682
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17788 16574 17816 18022
rect 17696 16546 17816 16574
rect 17696 15502 17724 16546
rect 17972 16522 18000 20159
rect 18064 19922 18092 20878
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18052 19236 18104 19242
rect 18052 19178 18104 19184
rect 18064 18970 18092 19178
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18156 18902 18184 21014
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18248 19990 18276 20266
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18340 19786 18368 21286
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18616 20262 18644 20946
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18156 18358 18184 18838
rect 18340 18601 18368 19382
rect 18432 19378 18460 19926
rect 18616 19514 18644 20198
rect 18708 19718 18736 20266
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18432 18970 18460 19314
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18524 18630 18552 19178
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18512 18624 18564 18630
rect 18326 18592 18382 18601
rect 18512 18566 18564 18572
rect 18326 18527 18382 18536
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18064 17610 18092 17682
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 18064 16998 18092 17138
rect 18052 16992 18104 16998
rect 18050 16960 18052 16969
rect 18104 16960 18106 16969
rect 18050 16895 18106 16904
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17958 15872 18014 15881
rect 17958 15807 18014 15816
rect 17776 15632 17828 15638
rect 17776 15574 17828 15580
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17696 14498 17724 15438
rect 17788 15366 17816 15574
rect 17972 15570 18000 15807
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 15042 17908 15302
rect 17880 15026 18000 15042
rect 17880 15020 18012 15026
rect 17880 15014 17960 15020
rect 17960 14962 18012 14968
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14618 17908 14894
rect 18064 14793 18092 16526
rect 18156 15638 18184 17206
rect 18248 16794 18276 17478
rect 18340 16833 18368 17682
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17338 18460 17478
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18326 16824 18382 16833
rect 18236 16788 18288 16794
rect 18326 16759 18382 16768
rect 18420 16788 18472 16794
rect 18236 16730 18288 16736
rect 18420 16730 18472 16736
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 18050 14784 18106 14793
rect 18050 14719 18106 14728
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17604 14470 17724 14498
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17500 14272 17552 14278
rect 17406 14240 17462 14249
rect 17500 14214 17552 14220
rect 17406 14175 17462 14184
rect 16960 13960 17080 13988
rect 17224 14000 17276 14006
rect 16854 13832 16910 13841
rect 16854 13767 16910 13776
rect 16868 13433 16896 13767
rect 16854 13424 16910 13433
rect 16854 13359 16910 13368
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16960 12696 16988 13960
rect 17224 13942 17276 13948
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17052 13394 17080 13806
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17038 13288 17094 13297
rect 17038 13223 17040 13232
rect 17092 13223 17094 13232
rect 17040 13194 17092 13200
rect 17040 12708 17092 12714
rect 16960 12668 17040 12696
rect 17040 12650 17092 12656
rect 16592 12600 16896 12628
rect 17052 12617 17080 12650
rect 16408 12406 16528 12434
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16316 10742 16344 11834
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16302 9888 16358 9897
rect 16302 9823 16358 9832
rect 16316 8430 16344 9823
rect 16408 9674 16436 12406
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16578 11384 16634 11393
rect 16578 11319 16634 11328
rect 16592 11218 16620 11319
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16500 10674 16528 11154
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16684 10470 16712 12242
rect 16868 11354 16896 12600
rect 17038 12608 17094 12617
rect 17038 12543 17094 12552
rect 17040 12300 17092 12306
rect 16960 12260 17040 12288
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16776 10849 16804 11086
rect 16762 10840 16818 10849
rect 16762 10775 16818 10784
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16408 9646 16528 9674
rect 16500 9586 16528 9646
rect 16592 9625 16620 10066
rect 16684 9926 16712 10202
rect 16776 10169 16804 10542
rect 16762 10160 16818 10169
rect 16762 10095 16818 10104
rect 16868 10062 16896 10542
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16672 9920 16724 9926
rect 16868 9897 16896 9998
rect 16672 9862 16724 9868
rect 16854 9888 16910 9897
rect 16854 9823 16910 9832
rect 16960 9654 16988 12260
rect 17040 12242 17092 12248
rect 17038 12200 17094 12209
rect 17038 12135 17094 12144
rect 17052 10690 17080 12135
rect 17144 10810 17172 13806
rect 17224 13388 17276 13394
rect 17420 13376 17448 14175
rect 17512 14074 17540 14214
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17604 13394 17632 14470
rect 17788 14113 17816 14554
rect 17774 14104 17830 14113
rect 18064 14090 18092 14719
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18064 14062 18184 14090
rect 17774 14039 17830 14048
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17592 13388 17644 13394
rect 17420 13348 17540 13376
rect 17224 13330 17276 13336
rect 17236 12918 17264 13330
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17328 12782 17356 13194
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12073 17264 12582
rect 17420 12442 17448 13194
rect 17512 13138 17540 13348
rect 17592 13330 17644 13336
rect 17604 13297 17632 13330
rect 17590 13288 17646 13297
rect 17590 13223 17646 13232
rect 17512 13110 17632 13138
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17316 12096 17368 12102
rect 17222 12064 17278 12073
rect 17316 12038 17368 12044
rect 17222 11999 17278 12008
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17052 10662 17172 10690
rect 17040 9988 17092 9994
rect 17040 9930 17092 9936
rect 16948 9648 17000 9654
rect 16578 9616 16634 9625
rect 16488 9580 16540 9586
rect 16948 9590 17000 9596
rect 16578 9551 16634 9560
rect 16672 9580 16724 9586
rect 16488 9522 16540 9528
rect 16396 9512 16448 9518
rect 16394 9480 16396 9489
rect 16448 9480 16450 9489
rect 16394 9415 16450 9424
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 8004 16344 8230
rect 16408 8129 16436 9114
rect 16500 8401 16528 9522
rect 16486 8392 16542 8401
rect 16486 8327 16488 8336
rect 16540 8327 16542 8336
rect 16488 8298 16540 8304
rect 16394 8120 16450 8129
rect 16394 8055 16450 8064
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16396 8016 16448 8022
rect 16316 7976 16396 8004
rect 16396 7958 16448 7964
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7342 16344 7686
rect 16408 7342 16436 7958
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16408 6254 16436 7278
rect 16500 7177 16528 8026
rect 16592 7206 16620 9551
rect 16672 9522 16724 9528
rect 16684 8537 16712 9522
rect 17052 9466 17080 9930
rect 16868 9438 17080 9466
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 9042 16804 9318
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16670 8528 16726 8537
rect 16776 8498 16804 8842
rect 16670 8463 16726 8472
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16670 8120 16726 8129
rect 16670 8055 16726 8064
rect 16684 7886 16712 8055
rect 16776 7886 16804 8298
rect 16868 8022 16896 9438
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7342 16712 7686
rect 16868 7546 16896 7822
rect 16960 7546 16988 9318
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17052 8838 17080 9046
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17052 8090 17080 8230
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16580 7200 16632 7206
rect 16486 7168 16542 7177
rect 16580 7142 16632 7148
rect 16486 7103 16542 7112
rect 16500 6866 16528 7103
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16500 5914 16528 6190
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16486 5808 16542 5817
rect 16592 5794 16620 6190
rect 16776 6186 16804 7278
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16542 5766 16620 5794
rect 16868 5778 16896 7346
rect 16946 7032 17002 7041
rect 16946 6967 17002 6976
rect 16856 5772 16908 5778
rect 16486 5743 16488 5752
rect 16540 5743 16542 5752
rect 16488 5714 16540 5720
rect 16856 5714 16908 5720
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4826 16436 4966
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16224 4282 16252 4558
rect 16960 4486 16988 6967
rect 17052 6730 17080 7890
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 17144 4690 17172 10662
rect 17236 9518 17264 11999
rect 17328 10452 17356 12038
rect 17420 11898 17448 12174
rect 17512 12170 17540 12922
rect 17604 12889 17632 13110
rect 17590 12880 17646 12889
rect 17590 12815 17646 12824
rect 17590 12336 17646 12345
rect 17590 12271 17592 12280
rect 17644 12271 17646 12280
rect 17592 12242 17644 12248
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11218 17448 11494
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17512 11121 17540 11290
rect 17498 11112 17554 11121
rect 17498 11047 17554 11056
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17420 10520 17448 10746
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17420 10492 17540 10520
rect 17328 10424 17448 10452
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17328 8838 17356 9862
rect 17420 9382 17448 10424
rect 17512 9738 17540 10492
rect 17604 10266 17632 10542
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17696 10146 17724 13942
rect 17788 13161 17816 14039
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17774 13152 17830 13161
rect 17774 13087 17830 13096
rect 17788 12782 17816 13087
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12306 17816 12582
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17776 10804 17828 10810
rect 17880 10792 17908 13806
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 17972 13025 18000 13194
rect 17958 13016 18014 13025
rect 17958 12951 18014 12960
rect 17960 12776 18012 12782
rect 18064 12764 18092 13942
rect 18156 13394 18184 14062
rect 18248 13938 18276 14554
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18248 13841 18276 13874
rect 18234 13832 18290 13841
rect 18234 13767 18290 13776
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18248 13002 18276 13767
rect 18012 12736 18092 12764
rect 18156 12974 18276 13002
rect 17960 12718 18012 12724
rect 17828 10764 17908 10792
rect 17776 10746 17828 10752
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17788 10305 17816 10542
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17774 10296 17830 10305
rect 17774 10231 17830 10240
rect 17788 10198 17816 10231
rect 17604 10118 17724 10146
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17604 9874 17632 10118
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17788 9897 17816 9930
rect 17774 9888 17830 9897
rect 17604 9846 17724 9874
rect 17512 9710 17632 9738
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17498 9344 17554 9353
rect 17498 9279 17554 9288
rect 17406 9208 17462 9217
rect 17406 9143 17462 9152
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17236 8498 17264 8774
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17328 8362 17356 8434
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17222 8120 17278 8129
rect 17222 8055 17278 8064
rect 17236 8022 17264 8055
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17420 7410 17448 9143
rect 17512 8974 17540 9279
rect 17604 9024 17632 9710
rect 17696 9160 17724 9846
rect 17774 9823 17830 9832
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17788 9586 17816 9658
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17880 9518 17908 10474
rect 17868 9512 17920 9518
rect 17774 9480 17830 9489
rect 17868 9454 17920 9460
rect 17774 9415 17776 9424
rect 17828 9415 17830 9424
rect 17776 9386 17828 9392
rect 17696 9132 17908 9160
rect 17775 9036 17827 9042
rect 17604 8996 17775 9024
rect 17775 8978 17827 8984
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17236 4826 17264 7142
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17328 4758 17356 7142
rect 17512 6866 17540 7482
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17420 6458 17448 6802
rect 17500 6724 17552 6730
rect 17604 6712 17632 8434
rect 17696 7274 17724 8774
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17788 6934 17816 8978
rect 17880 8838 17908 9132
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17880 8129 17908 8366
rect 17972 8294 18000 12718
rect 18156 12696 18184 12974
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18064 12668 18184 12696
rect 18064 12306 18092 12668
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18156 12170 18184 12378
rect 18144 12164 18196 12170
rect 18144 12106 18196 12112
rect 18248 12050 18276 12854
rect 18064 12022 18276 12050
rect 18064 9217 18092 12022
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 10606 18184 11494
rect 18248 10985 18276 11766
rect 18340 11762 18368 16662
rect 18432 14657 18460 16730
rect 18418 14648 18474 14657
rect 18418 14583 18474 14592
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18432 14074 18460 14418
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13530 18460 13874
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18432 12646 18460 13262
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18234 10976 18290 10985
rect 18234 10911 18290 10920
rect 18432 10656 18460 12582
rect 18524 12102 18552 18566
rect 18616 18329 18644 18702
rect 18708 18358 18736 19654
rect 18800 19242 18828 21830
rect 19210 21788 19518 21797
rect 19210 21786 19216 21788
rect 19272 21786 19296 21788
rect 19352 21786 19376 21788
rect 19432 21786 19456 21788
rect 19512 21786 19518 21788
rect 19272 21734 19274 21786
rect 19454 21734 19456 21786
rect 19210 21732 19216 21734
rect 19272 21732 19296 21734
rect 19352 21732 19376 21734
rect 19432 21732 19456 21734
rect 19512 21732 19518 21734
rect 19210 21723 19518 21732
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 22296 21570 22324 21626
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 18972 21412 19024 21418
rect 18972 21354 19024 21360
rect 18984 20602 19012 21354
rect 19064 21072 19116 21078
rect 19062 21040 19064 21049
rect 19116 21040 19118 21049
rect 19062 20975 19118 20984
rect 19444 20874 19472 21490
rect 20260 21412 20312 21418
rect 20628 21412 20680 21418
rect 20312 21372 20392 21400
rect 20260 21354 20312 21360
rect 19870 21244 20178 21253
rect 19870 21242 19876 21244
rect 19932 21242 19956 21244
rect 20012 21242 20036 21244
rect 20092 21242 20116 21244
rect 20172 21242 20178 21244
rect 19932 21190 19934 21242
rect 20114 21190 20116 21242
rect 19870 21188 19876 21190
rect 19932 21188 19956 21190
rect 20012 21188 20036 21190
rect 20092 21188 20116 21190
rect 20172 21188 20178 21190
rect 19870 21179 20178 21188
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19432 20868 19484 20874
rect 19432 20810 19484 20816
rect 19210 20700 19518 20709
rect 19210 20698 19216 20700
rect 19272 20698 19296 20700
rect 19352 20698 19376 20700
rect 19432 20698 19456 20700
rect 19512 20698 19518 20700
rect 19272 20646 19274 20698
rect 19454 20646 19456 20698
rect 19210 20644 19216 20646
rect 19272 20644 19296 20646
rect 19352 20644 19376 20646
rect 19432 20644 19456 20646
rect 19512 20644 19518 20646
rect 19210 20635 19518 20644
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18880 20528 18932 20534
rect 19628 20482 19656 20878
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 20088 20862 20300 20890
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 18880 20470 18932 20476
rect 18892 19990 18920 20470
rect 19536 20454 19656 20482
rect 19720 20466 19748 20742
rect 19708 20460 19760 20466
rect 19536 20398 19564 20454
rect 19708 20402 19760 20408
rect 19156 20392 19208 20398
rect 19524 20392 19576 20398
rect 19156 20334 19208 20340
rect 19444 20352 19524 20380
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18972 19984 19024 19990
rect 19168 19961 19196 20334
rect 19444 20058 19472 20352
rect 19524 20334 19576 20340
rect 19812 20312 19840 20810
rect 20088 20602 20116 20862
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19720 20284 19840 20312
rect 19720 20244 19748 20284
rect 19996 20262 20024 20334
rect 20076 20324 20128 20330
rect 20180 20312 20208 20742
rect 20128 20284 20208 20312
rect 20076 20266 20128 20272
rect 19628 20216 19748 20244
rect 19984 20256 20036 20262
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19524 19984 19576 19990
rect 18972 19926 19024 19932
rect 19154 19952 19210 19961
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18800 18465 18828 18838
rect 18892 18698 18920 19926
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18786 18456 18842 18465
rect 18786 18391 18842 18400
rect 18696 18352 18748 18358
rect 18602 18320 18658 18329
rect 18696 18294 18748 18300
rect 18602 18255 18658 18264
rect 18984 18222 19012 19926
rect 19628 19972 19656 20216
rect 19984 20198 20036 20204
rect 19870 20156 20178 20165
rect 19870 20154 19876 20156
rect 19932 20154 19956 20156
rect 20012 20154 20036 20156
rect 20092 20154 20116 20156
rect 20172 20154 20178 20156
rect 19932 20102 19934 20154
rect 20114 20102 20116 20154
rect 19870 20100 19876 20102
rect 19932 20100 19956 20102
rect 20012 20100 20036 20102
rect 20092 20100 20116 20102
rect 20172 20100 20178 20102
rect 19870 20091 20178 20100
rect 20272 20058 20300 20862
rect 20364 20602 20392 21372
rect 20628 21354 20680 21360
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 20640 21010 20668 21354
rect 20904 21344 20956 21350
rect 20902 21312 20904 21321
rect 20956 21312 20958 21321
rect 20902 21247 20958 21256
rect 21100 21128 21128 21354
rect 20916 21100 21128 21128
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20916 20890 20944 21100
rect 20996 21004 21048 21010
rect 20996 20946 21048 20952
rect 20640 20862 20944 20890
rect 21008 20890 21036 20946
rect 21008 20862 21128 20890
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20442 20224 20498 20233
rect 20442 20159 20498 20168
rect 20350 20088 20406 20097
rect 20260 20052 20312 20058
rect 20350 20023 20406 20032
rect 20260 19994 20312 20000
rect 19576 19944 19656 19972
rect 19524 19926 19576 19932
rect 19154 19887 19210 19896
rect 19340 19780 19392 19786
rect 19392 19740 19656 19768
rect 19340 19722 19392 19728
rect 19064 19712 19116 19718
rect 19628 19689 19656 19740
rect 19064 19654 19116 19660
rect 19614 19680 19670 19689
rect 19076 18902 19104 19654
rect 19210 19612 19518 19621
rect 19614 19615 19670 19624
rect 19210 19610 19216 19612
rect 19272 19610 19296 19612
rect 19352 19610 19376 19612
rect 19432 19610 19456 19612
rect 19512 19610 19518 19612
rect 19272 19558 19274 19610
rect 19454 19558 19456 19610
rect 19210 19556 19216 19558
rect 19272 19556 19296 19558
rect 19352 19556 19376 19558
rect 19432 19556 19456 19558
rect 19512 19556 19518 19558
rect 19210 19547 19518 19556
rect 20364 19446 20392 20023
rect 20456 19514 20484 20159
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20352 19440 20404 19446
rect 19890 19408 19946 19417
rect 19720 19366 19890 19394
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19628 18970 19656 19110
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 19248 18760 19300 18766
rect 19524 18760 19576 18766
rect 19300 18720 19524 18748
rect 19248 18702 19300 18708
rect 19524 18702 19576 18708
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19210 18524 19518 18533
rect 19210 18522 19216 18524
rect 19272 18522 19296 18524
rect 19352 18522 19376 18524
rect 19432 18522 19456 18524
rect 19512 18522 19518 18524
rect 19272 18470 19274 18522
rect 19454 18470 19456 18522
rect 19210 18468 19216 18470
rect 19272 18468 19296 18470
rect 19352 18468 19376 18470
rect 19432 18468 19456 18470
rect 19512 18468 19518 18470
rect 19210 18459 19518 18468
rect 19628 18426 19656 18634
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 18972 18216 19024 18222
rect 19156 18216 19208 18222
rect 18972 18158 19024 18164
rect 19076 18176 19156 18204
rect 18602 17776 18658 17785
rect 18602 17711 18604 17720
rect 18656 17711 18658 17720
rect 18604 17682 18656 17688
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18616 17066 18644 17478
rect 18984 17134 19012 17478
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18616 16794 18644 17002
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18602 16008 18658 16017
rect 18602 15943 18604 15952
rect 18656 15943 18658 15952
rect 18604 15914 18656 15920
rect 18602 14376 18658 14385
rect 18602 14311 18658 14320
rect 18616 12442 18644 14311
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18708 12306 18736 16050
rect 18800 13394 18828 16934
rect 18878 15464 18934 15473
rect 18878 15399 18934 15408
rect 18892 14074 18920 15399
rect 18984 14657 19012 17070
rect 18970 14648 19026 14657
rect 18970 14583 19026 14592
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 19076 14006 19104 18176
rect 19156 18158 19208 18164
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19536 17882 19564 18090
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19628 17814 19656 18022
rect 19720 17921 19748 19366
rect 20352 19382 20404 19388
rect 19890 19343 19946 19352
rect 20352 19304 20404 19310
rect 20536 19304 20588 19310
rect 20404 19264 20484 19292
rect 20352 19246 20404 19252
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19812 18442 19840 19178
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 19870 19068 20178 19077
rect 19870 19066 19876 19068
rect 19932 19066 19956 19068
rect 20012 19066 20036 19068
rect 20092 19066 20116 19068
rect 20172 19066 20178 19068
rect 19932 19014 19934 19066
rect 20114 19014 20116 19066
rect 19870 19012 19876 19014
rect 19932 19012 19956 19014
rect 20012 19012 20036 19014
rect 20092 19012 20116 19014
rect 20172 19012 20178 19014
rect 19870 19003 20178 19012
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19904 18601 19932 18906
rect 20272 18834 20300 19110
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19890 18592 19946 18601
rect 19890 18527 19946 18536
rect 19812 18414 19932 18442
rect 19800 18080 19852 18086
rect 19904 18068 19932 18414
rect 19996 18222 20024 18634
rect 20088 18329 20116 18702
rect 20272 18358 20300 18770
rect 20364 18698 20392 18770
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20260 18352 20312 18358
rect 20074 18320 20130 18329
rect 20260 18294 20312 18300
rect 20074 18255 20130 18264
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19984 18080 20036 18086
rect 19904 18040 19984 18068
rect 19800 18022 19852 18028
rect 20036 18040 20300 18068
rect 19984 18022 20036 18028
rect 19706 17912 19762 17921
rect 19706 17847 19762 17856
rect 19616 17808 19668 17814
rect 19616 17750 19668 17756
rect 19720 17626 19748 17847
rect 19628 17598 19748 17626
rect 19210 17436 19518 17445
rect 19210 17434 19216 17436
rect 19272 17434 19296 17436
rect 19352 17434 19376 17436
rect 19432 17434 19456 17436
rect 19512 17434 19518 17436
rect 19272 17382 19274 17434
rect 19454 17382 19456 17434
rect 19210 17380 19216 17382
rect 19272 17380 19296 17382
rect 19352 17380 19376 17382
rect 19432 17380 19456 17382
rect 19512 17380 19518 17382
rect 19210 17371 19518 17380
rect 19628 17218 19656 17598
rect 19812 17542 19840 18022
rect 19870 17980 20178 17989
rect 19870 17978 19876 17980
rect 19932 17978 19956 17980
rect 20012 17978 20036 17980
rect 20092 17978 20116 17980
rect 20172 17978 20178 17980
rect 19932 17926 19934 17978
rect 20114 17926 20116 17978
rect 19870 17924 19876 17926
rect 19932 17924 19956 17926
rect 20012 17924 20036 17926
rect 20092 17924 20116 17926
rect 20172 17924 20178 17926
rect 19870 17915 20178 17924
rect 20272 17921 20300 18040
rect 20258 17912 20314 17921
rect 19892 17876 19944 17882
rect 20258 17847 20314 17856
rect 19892 17818 19944 17824
rect 19904 17678 19932 17818
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19536 17190 19656 17218
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19352 16658 19380 17070
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19536 16436 19564 17190
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19628 16998 19656 17070
rect 19720 16998 19748 17478
rect 19812 17338 19840 17478
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 20088 17134 20116 17682
rect 20364 17678 20392 18634
rect 20456 18358 20484 19264
rect 20536 19246 20588 19252
rect 20548 18970 20576 19246
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20548 18222 20576 18906
rect 20640 18442 20668 20862
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 19310 20760 20742
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20824 19310 20852 19722
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20810 19000 20866 19009
rect 20916 18970 20944 19246
rect 20810 18935 20866 18944
rect 20904 18964 20956 18970
rect 20824 18834 20852 18935
rect 20904 18906 20956 18912
rect 20902 18864 20958 18873
rect 20812 18828 20864 18834
rect 20902 18799 20958 18808
rect 20812 18770 20864 18776
rect 20916 18630 20944 18799
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20640 18414 20760 18442
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20444 18148 20496 18154
rect 20444 18090 20496 18096
rect 20456 17746 20484 18090
rect 20640 17864 20668 18294
rect 20732 18086 20760 18414
rect 21008 18306 21036 19654
rect 21100 19174 21128 20862
rect 21192 20058 21220 21558
rect 22296 21542 22416 21570
rect 21270 21448 21326 21457
rect 21270 21383 21326 21392
rect 21284 21010 21312 21383
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21548 21004 21600 21010
rect 21600 20964 21680 20992
rect 21548 20946 21600 20952
rect 21456 20936 21508 20942
rect 21508 20884 21588 20890
rect 21456 20878 21588 20884
rect 21468 20862 21588 20878
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21284 20330 21312 20538
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18834 21128 19110
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21192 18766 21220 19994
rect 21284 19990 21312 20266
rect 21272 19984 21324 19990
rect 21272 19926 21324 19932
rect 21376 19836 21404 20402
rect 21284 19808 21404 19836
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 20824 18278 21036 18306
rect 21180 18352 21232 18358
rect 21284 18340 21312 19808
rect 21560 19718 21588 20862
rect 21652 20466 21680 20964
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21640 19984 21692 19990
rect 21640 19926 21692 19932
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21456 19304 21508 19310
rect 21362 19272 21418 19281
rect 21456 19246 21508 19252
rect 21362 19207 21364 19216
rect 21416 19207 21418 19216
rect 21364 19178 21416 19184
rect 21468 19145 21496 19246
rect 21454 19136 21510 19145
rect 21454 19071 21510 19080
rect 21468 18630 21496 19071
rect 21560 18873 21588 19654
rect 21652 19446 21680 19926
rect 21744 19514 21772 20266
rect 21836 19786 21864 20266
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21640 19440 21692 19446
rect 21692 19388 21864 19394
rect 21640 19382 21864 19388
rect 21652 19366 21864 19382
rect 21928 19378 21956 21082
rect 22282 20360 22338 20369
rect 22282 20295 22338 20304
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 21640 19236 21692 19242
rect 21640 19178 21692 19184
rect 21652 19009 21680 19178
rect 21638 19000 21694 19009
rect 21638 18935 21694 18944
rect 21546 18864 21602 18873
rect 21602 18822 21772 18850
rect 21546 18799 21602 18808
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21548 18624 21600 18630
rect 21548 18566 21600 18572
rect 21232 18312 21312 18340
rect 21180 18294 21232 18300
rect 21088 18284 21140 18290
rect 20824 18222 20852 18278
rect 21088 18226 21140 18232
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20548 17836 20668 17864
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20272 17134 20300 17546
rect 19800 17128 19852 17134
rect 19984 17128 20036 17134
rect 19800 17070 19852 17076
rect 19982 17096 19984 17105
rect 20076 17128 20128 17134
rect 20036 17096 20038 17105
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19536 16408 19656 16436
rect 19720 16425 19748 16730
rect 19812 16658 19840 17070
rect 20076 17070 20128 17076
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 19982 17031 20038 17040
rect 19870 16892 20178 16901
rect 19870 16890 19876 16892
rect 19932 16890 19956 16892
rect 20012 16890 20036 16892
rect 20092 16890 20116 16892
rect 20172 16890 20178 16892
rect 19932 16838 19934 16890
rect 20114 16838 20116 16890
rect 19870 16836 19876 16838
rect 19932 16836 19956 16838
rect 20012 16836 20036 16838
rect 20092 16836 20116 16838
rect 20172 16836 20178 16838
rect 19870 16827 20178 16836
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19210 16348 19518 16357
rect 19210 16346 19216 16348
rect 19272 16346 19296 16348
rect 19352 16346 19376 16348
rect 19432 16346 19456 16348
rect 19512 16346 19518 16348
rect 19272 16294 19274 16346
rect 19454 16294 19456 16346
rect 19210 16292 19216 16294
rect 19272 16292 19296 16294
rect 19352 16292 19376 16294
rect 19432 16292 19456 16294
rect 19512 16292 19518 16294
rect 19210 16283 19518 16292
rect 19628 16164 19656 16408
rect 19706 16416 19762 16425
rect 19706 16351 19762 16360
rect 19706 16280 19762 16289
rect 19812 16250 19840 16458
rect 19982 16280 20038 16289
rect 19706 16215 19762 16224
rect 19800 16244 19852 16250
rect 19444 16136 19656 16164
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15978 19288 16050
rect 19444 15978 19472 16136
rect 19720 16096 19748 16215
rect 20272 16250 20300 17070
rect 20548 16776 20576 17836
rect 20732 17746 20760 17847
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20720 17740 20772 17746
rect 20772 17700 20852 17728
rect 20720 17682 20772 17688
rect 20640 17338 20668 17682
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20626 17096 20682 17105
rect 20626 17031 20682 17040
rect 20364 16748 20576 16776
rect 19982 16215 19984 16224
rect 19800 16186 19852 16192
rect 20036 16215 20038 16224
rect 20260 16244 20312 16250
rect 19984 16186 20036 16192
rect 20260 16186 20312 16192
rect 19536 16068 19748 16096
rect 19800 16108 19852 16114
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19352 15366 19380 15846
rect 19536 15570 19564 16068
rect 19800 16050 19852 16056
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19708 15496 19760 15502
rect 19706 15464 19708 15473
rect 19760 15464 19762 15473
rect 19706 15399 19762 15408
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19614 15328 19670 15337
rect 19210 15260 19518 15269
rect 19614 15263 19670 15272
rect 19210 15258 19216 15260
rect 19272 15258 19296 15260
rect 19352 15258 19376 15260
rect 19432 15258 19456 15260
rect 19512 15258 19518 15260
rect 19272 15206 19274 15258
rect 19454 15206 19456 15258
rect 19210 15204 19216 15206
rect 19272 15204 19296 15206
rect 19352 15204 19376 15206
rect 19432 15204 19456 15206
rect 19512 15204 19518 15206
rect 19210 15195 19518 15204
rect 19628 15144 19656 15263
rect 19444 15116 19656 15144
rect 19338 15056 19394 15065
rect 19338 14991 19340 15000
rect 19392 14991 19394 15000
rect 19340 14962 19392 14968
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 14657 19380 14758
rect 19338 14648 19394 14657
rect 19444 14618 19472 15116
rect 19720 15008 19748 15399
rect 19536 14980 19748 15008
rect 19338 14583 19394 14592
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19536 14482 19564 14980
rect 19812 14940 19840 16050
rect 19870 15804 20178 15813
rect 19870 15802 19876 15804
rect 19932 15802 19956 15804
rect 20012 15802 20036 15804
rect 20092 15802 20116 15804
rect 20172 15802 20178 15804
rect 19932 15750 19934 15802
rect 20114 15750 20116 15802
rect 19870 15748 19876 15750
rect 19932 15748 19956 15750
rect 20012 15748 20036 15750
rect 20092 15748 20116 15750
rect 20172 15748 20178 15750
rect 19870 15739 20178 15748
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 15026 20116 15506
rect 20180 15502 20208 15642
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20272 15042 20300 15642
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20180 15014 20300 15042
rect 19628 14912 19840 14940
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19340 14408 19392 14414
rect 19154 14376 19210 14385
rect 19154 14311 19156 14320
rect 19208 14311 19210 14320
rect 19338 14376 19340 14385
rect 19432 14408 19484 14414
rect 19392 14376 19394 14385
rect 19432 14350 19484 14356
rect 19338 14311 19394 14320
rect 19156 14282 19208 14288
rect 19444 14260 19472 14350
rect 19628 14328 19656 14912
rect 20180 14890 20208 15014
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 19892 14884 19944 14890
rect 19812 14844 19892 14872
rect 19706 14648 19762 14657
rect 19706 14583 19708 14592
rect 19760 14583 19762 14592
rect 19708 14554 19760 14560
rect 19628 14300 19748 14328
rect 19444 14232 19656 14260
rect 19210 14172 19518 14181
rect 19210 14170 19216 14172
rect 19272 14170 19296 14172
rect 19352 14170 19376 14172
rect 19432 14170 19456 14172
rect 19512 14170 19518 14172
rect 19272 14118 19274 14170
rect 19454 14118 19456 14170
rect 19210 14116 19216 14118
rect 19272 14116 19296 14118
rect 19352 14116 19376 14118
rect 19432 14116 19456 14118
rect 19512 14116 19518 14118
rect 19210 14107 19518 14116
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19432 14068 19484 14074
rect 19628 14056 19656 14232
rect 19432 14010 19484 14016
rect 19536 14028 19656 14056
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19156 13864 19208 13870
rect 18892 13824 19156 13852
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18892 13297 18920 13824
rect 19156 13806 19208 13812
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19156 13728 19208 13734
rect 18970 13696 19026 13705
rect 18970 13631 19026 13640
rect 19154 13696 19156 13705
rect 19208 13696 19210 13705
rect 19154 13631 19210 13640
rect 18984 13530 19012 13631
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19260 13394 19288 13806
rect 19064 13388 19116 13394
rect 18984 13348 19064 13376
rect 18878 13288 18934 13297
rect 18878 13223 18934 13232
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18616 11914 18644 12174
rect 18708 11937 18736 12242
rect 18800 12073 18828 12922
rect 18984 12594 19012 13348
rect 19064 13330 19116 13336
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19168 13297 19196 13330
rect 19154 13288 19210 13297
rect 19154 13223 19210 13232
rect 19260 13172 19288 13330
rect 19352 13326 19380 14010
rect 19444 13870 19472 14010
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19536 13190 19564 14028
rect 19616 13728 19668 13734
rect 19614 13696 19616 13705
rect 19668 13696 19670 13705
rect 19614 13631 19670 13640
rect 19076 13144 19288 13172
rect 19524 13184 19576 13190
rect 19076 12968 19104 13144
rect 19524 13126 19576 13132
rect 19210 13084 19518 13093
rect 19210 13082 19216 13084
rect 19272 13082 19296 13084
rect 19352 13082 19376 13084
rect 19432 13082 19456 13084
rect 19512 13082 19518 13084
rect 19272 13030 19274 13082
rect 19454 13030 19456 13082
rect 19210 13028 19216 13030
rect 19272 13028 19296 13030
rect 19352 13028 19376 13030
rect 19432 13028 19456 13030
rect 19512 13028 19518 13030
rect 19210 13019 19518 13028
rect 19720 12968 19748 14300
rect 19812 14074 19840 14844
rect 19892 14826 19944 14832
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 19870 14716 20178 14725
rect 19870 14714 19876 14716
rect 19932 14714 19956 14716
rect 20012 14714 20036 14716
rect 20092 14714 20116 14716
rect 20172 14714 20178 14716
rect 19932 14662 19934 14714
rect 20114 14662 20116 14714
rect 19870 14660 19876 14662
rect 19932 14660 19956 14662
rect 20012 14660 20036 14662
rect 20092 14660 20116 14662
rect 20172 14660 20178 14662
rect 19870 14651 20178 14660
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19996 14482 20024 14554
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19904 14074 19932 14282
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19890 13832 19946 13841
rect 19076 12940 19196 12968
rect 19168 12782 19196 12940
rect 19628 12940 19748 12968
rect 19812 13790 19890 13818
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19156 12776 19208 12782
rect 19444 12753 19472 12786
rect 19156 12718 19208 12724
rect 19430 12744 19486 12753
rect 19340 12708 19392 12714
rect 19430 12679 19486 12688
rect 19524 12708 19576 12714
rect 19340 12650 19392 12656
rect 19524 12650 19576 12656
rect 18984 12566 19104 12594
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18786 12064 18842 12073
rect 18786 11999 18842 12008
rect 18248 10628 18460 10656
rect 18524 11886 18644 11914
rect 18694 11928 18750 11937
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18050 9208 18106 9217
rect 18050 9143 18106 9152
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18064 8430 18092 8910
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17866 8120 17922 8129
rect 17866 8055 17922 8064
rect 17880 7041 17908 8055
rect 18064 7410 18092 8366
rect 18156 7546 18184 10542
rect 18248 10130 18276 10628
rect 18524 10606 18552 11886
rect 18694 11863 18750 11872
rect 18694 11792 18750 11801
rect 18694 11727 18696 11736
rect 18748 11727 18750 11736
rect 18696 11698 18748 11704
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18512 10600 18564 10606
rect 18432 10560 18512 10588
rect 18326 10296 18382 10305
rect 18326 10231 18382 10240
rect 18340 10198 18368 10231
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18234 9888 18290 9897
rect 18234 9823 18290 9832
rect 18248 9722 18276 9823
rect 18340 9761 18368 9998
rect 18326 9752 18382 9761
rect 18236 9716 18288 9722
rect 18326 9687 18382 9696
rect 18236 9658 18288 9664
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18248 8634 18276 9454
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18248 8129 18276 8366
rect 18234 8120 18290 8129
rect 18234 8055 18290 8064
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17866 7032 17922 7041
rect 17866 6967 17922 6976
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17552 6684 17632 6712
rect 17500 6666 17552 6672
rect 17696 6610 17724 6802
rect 17512 6582 17724 6610
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17512 5370 17540 6582
rect 17682 6352 17738 6361
rect 17682 6287 17738 6296
rect 17696 5778 17724 6287
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16868 4282 16896 4422
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 17144 4214 17172 4626
rect 17420 4622 17448 4762
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 4457 17448 4558
rect 17406 4448 17462 4457
rect 17406 4383 17462 4392
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 17696 3942 17724 5714
rect 17788 5710 17816 6870
rect 17972 6866 18000 7210
rect 18248 6984 18276 7822
rect 18156 6956 18276 6984
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17880 6225 17908 6802
rect 18156 6497 18184 6956
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18142 6488 18198 6497
rect 17960 6452 18012 6458
rect 18142 6423 18198 6432
rect 17960 6394 18012 6400
rect 17866 6216 17922 6225
rect 17866 6151 17922 6160
rect 17972 5778 18000 6394
rect 18248 6390 18276 6802
rect 18340 6458 18368 9454
rect 18432 6662 18460 10560
rect 18512 10542 18564 10548
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18524 9024 18552 10066
rect 18616 9722 18644 11630
rect 18892 11626 18920 12174
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18786 11112 18842 11121
rect 18786 11047 18842 11056
rect 18696 10464 18748 10470
rect 18694 10432 18696 10441
rect 18748 10432 18750 10441
rect 18694 10367 18750 10376
rect 18800 9874 18828 11047
rect 18892 11014 18920 11562
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18880 10600 18932 10606
rect 18984 10588 19012 12378
rect 19076 12306 19104 12566
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19076 11121 19104 12242
rect 19260 12170 19288 12378
rect 19352 12170 19380 12650
rect 19536 12481 19564 12650
rect 19522 12472 19578 12481
rect 19522 12407 19578 12416
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19210 11996 19518 12005
rect 19210 11994 19216 11996
rect 19272 11994 19296 11996
rect 19352 11994 19376 11996
rect 19432 11994 19456 11996
rect 19512 11994 19518 11996
rect 19272 11942 19274 11994
rect 19454 11942 19456 11994
rect 19210 11940 19216 11942
rect 19272 11940 19296 11942
rect 19352 11940 19376 11942
rect 19432 11940 19456 11942
rect 19512 11940 19518 11942
rect 19210 11931 19518 11940
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19444 11694 19472 11834
rect 19522 11792 19578 11801
rect 19522 11727 19524 11736
rect 19576 11727 19578 11736
rect 19524 11698 19576 11704
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19524 11552 19576 11558
rect 19522 11520 19524 11529
rect 19576 11520 19578 11529
rect 19522 11455 19578 11464
rect 19628 11218 19656 12940
rect 19812 12866 19840 13790
rect 20180 13802 20208 14214
rect 19890 13767 19946 13776
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 20272 13705 20300 14894
rect 20364 14414 20392 16748
rect 20640 16658 20668 17031
rect 20824 16726 20852 17700
rect 21008 17270 21036 18022
rect 21100 17882 21128 18226
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21192 17746 21220 18294
rect 21468 18170 21496 18566
rect 21560 18358 21588 18566
rect 21652 18465 21680 18634
rect 21638 18456 21694 18465
rect 21638 18391 21694 18400
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21284 18142 21496 18170
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21086 17640 21142 17649
rect 21086 17575 21142 17584
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20902 16688 20958 16697
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20442 15736 20498 15745
rect 20442 15671 20498 15680
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20456 14074 20484 15671
rect 20548 14793 20576 16594
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20534 14784 20590 14793
rect 20640 14770 20668 16458
rect 20824 15910 20852 16662
rect 20902 16623 20904 16632
rect 20956 16623 20958 16632
rect 20904 16594 20956 16600
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20916 16289 20944 16390
rect 20902 16280 20958 16289
rect 20902 16215 20958 16224
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20824 15706 20852 15846
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20732 14890 20760 15574
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20640 14742 20760 14770
rect 20534 14719 20590 14728
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20548 13954 20576 14350
rect 20548 13926 20668 13954
rect 20536 13864 20588 13870
rect 20534 13832 20536 13841
rect 20588 13832 20590 13841
rect 20352 13796 20404 13802
rect 20534 13767 20590 13776
rect 20352 13738 20404 13744
rect 20258 13696 20314 13705
rect 19870 13628 20178 13637
rect 20258 13631 20314 13640
rect 19870 13626 19876 13628
rect 19932 13626 19956 13628
rect 20012 13626 20036 13628
rect 20092 13626 20116 13628
rect 20172 13626 20178 13628
rect 19932 13574 19934 13626
rect 20114 13574 20116 13626
rect 19870 13572 19876 13574
rect 19932 13572 19956 13574
rect 20012 13572 20036 13574
rect 20092 13572 20116 13574
rect 20172 13572 20178 13574
rect 19870 13563 20178 13572
rect 20076 13456 20128 13462
rect 20272 13410 20300 13631
rect 20076 13398 20128 13404
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19720 12838 19840 12866
rect 19720 12617 19748 12838
rect 19800 12776 19852 12782
rect 19798 12744 19800 12753
rect 19852 12744 19854 12753
rect 19798 12679 19854 12688
rect 19904 12628 19932 13330
rect 20088 13190 20116 13398
rect 20180 13382 20300 13410
rect 20364 13394 20392 13738
rect 20352 13388 20404 13394
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 19996 12646 20024 13126
rect 20180 12986 20208 13382
rect 20352 13330 20404 13336
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 13025 20300 13262
rect 20640 13190 20668 13926
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20258 13016 20314 13025
rect 20168 12980 20220 12986
rect 20258 12951 20314 12960
rect 20168 12922 20220 12928
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 19706 12608 19762 12617
rect 19706 12543 19762 12552
rect 19812 12600 19932 12628
rect 19984 12640 20036 12646
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19720 11354 19748 12242
rect 19812 11642 19840 12600
rect 19984 12582 20036 12588
rect 19870 12540 20178 12549
rect 19870 12538 19876 12540
rect 19932 12538 19956 12540
rect 20012 12538 20036 12540
rect 20092 12538 20116 12540
rect 20172 12538 20178 12540
rect 19932 12486 19934 12538
rect 20114 12486 20116 12538
rect 19870 12484 19876 12486
rect 19932 12484 19956 12486
rect 20012 12484 20036 12486
rect 20092 12484 20116 12486
rect 20172 12484 20178 12486
rect 19870 12475 20178 12484
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20076 11824 20128 11830
rect 20180 11812 20208 12174
rect 20128 11784 20208 11812
rect 20076 11766 20128 11772
rect 19812 11626 20116 11642
rect 19812 11620 20128 11626
rect 19812 11614 20076 11620
rect 20076 11562 20128 11568
rect 19870 11452 20178 11461
rect 19870 11450 19876 11452
rect 19932 11450 19956 11452
rect 20012 11450 20036 11452
rect 20092 11450 20116 11452
rect 20172 11450 20178 11452
rect 19932 11398 19934 11450
rect 20114 11398 20116 11450
rect 19870 11396 19876 11398
rect 19932 11396 19956 11398
rect 20012 11396 20036 11398
rect 20092 11396 20116 11398
rect 20172 11396 20178 11398
rect 19870 11387 20178 11396
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19062 11112 19118 11121
rect 19062 11047 19118 11056
rect 19168 10996 19196 11154
rect 19720 11064 19748 11154
rect 19904 11082 19932 11290
rect 20272 11234 20300 12718
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 12442 20392 12582
rect 20456 12481 20484 13126
rect 20732 12850 20760 14742
rect 20824 14618 20852 15370
rect 20916 15337 20944 15642
rect 21008 15366 21036 17206
rect 21100 17105 21128 17575
rect 21086 17096 21142 17105
rect 21086 17031 21142 17040
rect 21088 16992 21140 16998
rect 21086 16960 21088 16969
rect 21140 16960 21142 16969
rect 21086 16895 21142 16904
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 20996 15360 21048 15366
rect 20902 15328 20958 15337
rect 20996 15302 21048 15308
rect 20902 15263 20958 15272
rect 21100 15178 21128 16730
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21192 15745 21220 15982
rect 21178 15736 21234 15745
rect 21178 15671 21234 15680
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 15473 21220 15506
rect 21178 15464 21234 15473
rect 21178 15399 21234 15408
rect 20916 15150 21128 15178
rect 21180 15156 21232 15162
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20824 13841 20852 14010
rect 20916 13938 20944 15150
rect 21180 15098 21232 15104
rect 20994 15056 21050 15065
rect 20994 14991 21050 15000
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20810 13832 20866 13841
rect 20810 13767 20866 13776
rect 20916 13394 20944 13874
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20534 12608 20590 12617
rect 20534 12543 20590 12552
rect 20442 12472 20498 12481
rect 20352 12436 20404 12442
rect 20442 12407 20498 12416
rect 20352 12378 20404 12384
rect 20364 12322 20392 12378
rect 20548 12374 20576 12543
rect 20536 12368 20588 12374
rect 20364 12294 20484 12322
rect 20536 12310 20588 12316
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 19996 11218 20300 11234
rect 19984 11212 20300 11218
rect 20036 11206 20300 11212
rect 19984 11154 20036 11160
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19076 10968 19196 10996
rect 19628 11036 19748 11064
rect 19892 11076 19944 11082
rect 19076 10792 19104 10968
rect 19210 10908 19518 10917
rect 19210 10906 19216 10908
rect 19272 10906 19296 10908
rect 19352 10906 19376 10908
rect 19432 10906 19456 10908
rect 19512 10906 19518 10908
rect 19272 10854 19274 10906
rect 19454 10854 19456 10906
rect 19210 10852 19216 10854
rect 19272 10852 19296 10854
rect 19352 10852 19376 10854
rect 19432 10852 19456 10854
rect 19512 10852 19518 10854
rect 19210 10843 19518 10852
rect 19076 10764 19380 10792
rect 19246 10704 19302 10713
rect 19246 10639 19302 10648
rect 19156 10600 19208 10606
rect 18984 10560 19156 10588
rect 18880 10542 18932 10548
rect 19156 10542 19208 10548
rect 18708 9846 18828 9874
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18604 9376 18656 9382
rect 18602 9344 18604 9353
rect 18656 9344 18658 9353
rect 18602 9279 18658 9288
rect 18524 8996 18644 9024
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18524 8809 18552 8842
rect 18510 8800 18566 8809
rect 18510 8735 18566 8744
rect 18510 8392 18566 8401
rect 18510 8327 18566 8336
rect 18524 8294 18552 8327
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18616 8106 18644 8996
rect 18708 8809 18736 9846
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18800 9042 18828 9658
rect 18892 9568 18920 10542
rect 19154 10432 19210 10441
rect 19154 10367 19210 10376
rect 19168 9994 19196 10367
rect 19260 10062 19288 10639
rect 19352 10470 19380 10764
rect 19628 10656 19656 11036
rect 19892 11018 19944 11024
rect 19984 11008 20036 11014
rect 19720 10956 19984 10962
rect 19720 10950 20036 10956
rect 20088 10962 20116 11086
rect 19720 10934 20024 10950
rect 20088 10934 20300 10962
rect 19720 10674 19748 10934
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 19536 10628 19656 10656
rect 19708 10668 19760 10674
rect 19430 10568 19486 10577
rect 19430 10503 19486 10512
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19338 10296 19394 10305
rect 19338 10231 19394 10240
rect 19352 10062 19380 10231
rect 19444 10062 19472 10503
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19536 9908 19564 10628
rect 19708 10610 19760 10616
rect 19614 10568 19670 10577
rect 20180 10538 20208 10678
rect 19614 10503 19616 10512
rect 19668 10503 19670 10512
rect 20168 10532 20220 10538
rect 19616 10474 19668 10480
rect 20168 10474 20220 10480
rect 19708 10464 19760 10470
rect 19614 10432 19670 10441
rect 19892 10464 19944 10470
rect 19708 10406 19760 10412
rect 19812 10424 19892 10452
rect 19614 10367 19670 10376
rect 19628 10010 19656 10367
rect 19720 10112 19748 10406
rect 19812 10180 19840 10424
rect 19892 10406 19944 10412
rect 19870 10364 20178 10373
rect 19870 10362 19876 10364
rect 19932 10362 19956 10364
rect 20012 10362 20036 10364
rect 20092 10362 20116 10364
rect 20172 10362 20178 10364
rect 19932 10310 19934 10362
rect 20114 10310 20116 10362
rect 19870 10308 19876 10310
rect 19932 10308 19956 10310
rect 20012 10308 20036 10310
rect 20092 10308 20116 10310
rect 20172 10308 20178 10310
rect 19870 10299 20178 10308
rect 19812 10152 20116 10180
rect 19720 10084 20024 10112
rect 19890 10024 19946 10033
rect 19628 9982 19890 10010
rect 19890 9959 19946 9968
rect 19536 9880 19656 9908
rect 19210 9820 19518 9829
rect 19210 9818 19216 9820
rect 19272 9818 19296 9820
rect 19352 9818 19376 9820
rect 19432 9818 19456 9820
rect 19512 9818 19518 9820
rect 19272 9766 19274 9818
rect 19454 9766 19456 9818
rect 19210 9764 19216 9766
rect 19272 9764 19296 9766
rect 19352 9764 19376 9766
rect 19432 9764 19456 9766
rect 19512 9764 19518 9766
rect 19210 9755 19518 9764
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19156 9648 19208 9654
rect 19208 9608 19288 9636
rect 19156 9590 19208 9596
rect 18972 9580 19024 9586
rect 18892 9540 18972 9568
rect 18892 9489 18920 9540
rect 18972 9522 19024 9528
rect 19156 9512 19208 9518
rect 18878 9480 18934 9489
rect 19156 9454 19208 9460
rect 18878 9415 18934 9424
rect 18972 9444 19024 9450
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18694 8800 18750 8809
rect 18694 8735 18750 8744
rect 18694 8528 18750 8537
rect 18694 8463 18696 8472
rect 18748 8463 18750 8472
rect 18696 8434 18748 8440
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18524 8078 18644 8106
rect 18708 8090 18736 8298
rect 18800 8129 18828 8298
rect 18786 8120 18842 8129
rect 18696 8084 18748 8090
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18248 5914 18276 6326
rect 18524 6304 18552 8078
rect 18786 8055 18842 8064
rect 18696 8026 18748 8032
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18786 7984 18842 7993
rect 18432 6276 18552 6304
rect 18432 6089 18460 6276
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18418 6080 18474 6089
rect 18418 6015 18474 6024
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 18432 5166 18460 6015
rect 18524 5778 18552 6122
rect 18616 5846 18644 7958
rect 18786 7919 18788 7928
rect 18840 7919 18842 7928
rect 18788 7890 18840 7896
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18708 6934 18736 7686
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18708 5624 18736 6598
rect 18800 6186 18828 7346
rect 18892 6866 18920 9415
rect 18972 9386 19024 9392
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 18984 9353 19012 9386
rect 18970 9344 19026 9353
rect 18970 9279 19026 9288
rect 18984 9178 19012 9279
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18984 8362 19012 8570
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18970 8120 19026 8129
rect 18970 8055 18972 8064
rect 19024 8055 19026 8064
rect 18972 8026 19024 8032
rect 18984 7954 19012 8026
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18970 7304 19026 7313
rect 18970 7239 19026 7248
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18878 6488 18934 6497
rect 18878 6423 18934 6432
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18892 6118 18920 6423
rect 18880 6112 18932 6118
rect 18984 6089 19012 7239
rect 18880 6054 18932 6060
rect 18970 6080 19026 6089
rect 18616 5596 18736 5624
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4078 18000 5034
rect 18432 4758 18460 5102
rect 18616 4826 18644 5596
rect 18694 5536 18750 5545
rect 18694 5471 18750 5480
rect 18708 5166 18736 5471
rect 18892 5409 18920 6054
rect 18970 6015 19026 6024
rect 19076 5914 19104 9386
rect 19168 9042 19196 9454
rect 19260 9382 19288 9608
rect 19340 9580 19392 9586
rect 19444 9568 19472 9658
rect 19392 9540 19472 9568
rect 19340 9522 19392 9528
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19352 8838 19380 9386
rect 19536 8906 19564 9454
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19210 8732 19518 8741
rect 19210 8730 19216 8732
rect 19272 8730 19296 8732
rect 19352 8730 19376 8732
rect 19432 8730 19456 8732
rect 19512 8730 19518 8732
rect 19272 8678 19274 8730
rect 19454 8678 19456 8730
rect 19210 8676 19216 8678
rect 19272 8676 19296 8678
rect 19352 8676 19376 8678
rect 19432 8676 19456 8678
rect 19512 8676 19518 8678
rect 19210 8667 19518 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19168 7954 19196 8230
rect 19260 7954 19288 8502
rect 19444 7954 19472 8570
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19260 7750 19288 7890
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 7750 19380 7822
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19210 7644 19518 7653
rect 19210 7642 19216 7644
rect 19272 7642 19296 7644
rect 19352 7642 19376 7644
rect 19432 7642 19456 7644
rect 19512 7642 19518 7644
rect 19272 7590 19274 7642
rect 19454 7590 19456 7642
rect 19210 7588 19216 7590
rect 19272 7588 19296 7590
rect 19352 7588 19376 7590
rect 19432 7588 19456 7590
rect 19512 7588 19518 7590
rect 19210 7579 19518 7588
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 6934 19564 7346
rect 19524 6928 19576 6934
rect 19524 6870 19576 6876
rect 19628 6866 19656 9880
rect 19890 9888 19946 9897
rect 19812 9846 19890 9874
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19720 9353 19748 9454
rect 19706 9344 19762 9353
rect 19706 9279 19762 9288
rect 19706 9208 19762 9217
rect 19706 9143 19708 9152
rect 19760 9143 19762 9152
rect 19708 9114 19760 9120
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19720 8809 19748 8978
rect 19812 8838 19840 9846
rect 19890 9823 19946 9832
rect 19996 9722 20024 10084
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20088 9586 20116 10152
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19870 9276 20178 9285
rect 19870 9274 19876 9276
rect 19932 9274 19956 9276
rect 20012 9274 20036 9276
rect 20092 9274 20116 9276
rect 20172 9274 20178 9276
rect 19932 9222 19934 9274
rect 20114 9222 20116 9274
rect 19870 9220 19876 9222
rect 19932 9220 19956 9222
rect 20012 9220 20036 9222
rect 20092 9220 20116 9222
rect 20172 9220 20178 9222
rect 19870 9211 20178 9220
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19800 8832 19852 8838
rect 19706 8800 19762 8809
rect 19800 8774 19852 8780
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19706 8735 19762 8744
rect 19812 8650 19840 8774
rect 19720 8622 19840 8650
rect 19720 8265 19748 8622
rect 19904 8548 19932 8774
rect 19996 8566 20024 8842
rect 19812 8520 19932 8548
rect 19984 8560 20036 8566
rect 19706 8256 19762 8265
rect 19706 8191 19762 8200
rect 19812 8106 19840 8520
rect 19984 8502 20036 8508
rect 20074 8392 20130 8401
rect 20074 8327 20076 8336
rect 20128 8327 20130 8336
rect 20180 8344 20208 8978
rect 20272 8838 20300 10934
rect 20364 10674 20392 12174
rect 20456 12073 20484 12294
rect 20442 12064 20498 12073
rect 20442 11999 20498 12008
rect 20534 11928 20590 11937
rect 20534 11863 20536 11872
rect 20588 11863 20590 11872
rect 20536 11834 20588 11840
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20456 11218 20484 11290
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20442 10976 20498 10985
rect 20442 10911 20498 10920
rect 20456 10674 20484 10911
rect 20548 10792 20576 11834
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20548 10764 20606 10792
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20444 10566 20496 10572
rect 20364 10526 20444 10554
rect 20364 9674 20392 10526
rect 20444 10508 20496 10514
rect 20578 10452 20606 10764
rect 20640 10588 20668 11562
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10742 20760 10950
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20640 10560 20760 10588
rect 20456 10424 20606 10452
rect 20732 10441 20760 10560
rect 20718 10432 20774 10441
rect 20456 9897 20484 10424
rect 20718 10367 20774 10376
rect 20718 10296 20774 10305
rect 20718 10231 20774 10240
rect 20732 10198 20760 10231
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20640 9897 20668 10066
rect 20824 10044 20852 12922
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20916 11257 20944 12582
rect 21008 12345 21036 14991
rect 21088 14884 21140 14890
rect 21192 14872 21220 15098
rect 21140 14844 21220 14872
rect 21088 14826 21140 14832
rect 21100 12986 21128 14826
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21192 13802 21220 14282
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21284 13410 21312 18142
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21376 17134 21404 18022
rect 21560 17954 21588 18022
rect 21468 17926 21588 17954
rect 21468 17814 21496 17926
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21560 17649 21588 17926
rect 21546 17640 21602 17649
rect 21546 17575 21602 17584
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 16454 21404 16934
rect 21560 16658 21588 17575
rect 21640 17536 21692 17542
rect 21640 17478 21692 17484
rect 21652 17202 21680 17478
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21744 17134 21772 18822
rect 21836 18290 21864 19366
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 22112 19174 22140 19654
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22190 18864 22246 18873
rect 22190 18799 22246 18808
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21822 18184 21878 18193
rect 21822 18119 21878 18128
rect 21916 18148 21968 18154
rect 21836 17377 21864 18119
rect 21916 18090 21968 18096
rect 21928 17882 21956 18090
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22006 17912 22062 17921
rect 21916 17876 21968 17882
rect 22006 17847 22062 17856
rect 21916 17818 21968 17824
rect 21822 17368 21878 17377
rect 21822 17303 21878 17312
rect 21836 17134 21864 17303
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 22020 16998 22048 17847
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22112 16833 22140 18022
rect 22204 17270 22232 18799
rect 22192 17264 22244 17270
rect 22192 17206 22244 17212
rect 22296 17066 22324 20295
rect 22388 18601 22416 21542
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 23020 21480 23072 21486
rect 23020 21422 23072 21428
rect 22940 21010 22968 21422
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22834 20768 22890 20777
rect 22834 20703 22890 20712
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22756 18834 22784 20198
rect 22848 19242 22876 20703
rect 22940 20602 22968 20946
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22940 19990 22968 20538
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 23032 19689 23060 21422
rect 23124 21350 23152 21626
rect 24124 21412 24176 21418
rect 24124 21354 24176 21360
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 23112 21344 23164 21350
rect 24032 21344 24084 21350
rect 23112 21286 23164 21292
rect 23938 21312 23994 21321
rect 23124 21146 23152 21286
rect 24032 21286 24084 21292
rect 23938 21247 23994 21256
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23492 20466 23520 20946
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23492 20058 23520 20402
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23296 19984 23348 19990
rect 23348 19944 23428 19972
rect 23296 19926 23348 19932
rect 23018 19680 23074 19689
rect 23018 19615 23074 19624
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 23112 19236 23164 19242
rect 23112 19178 23164 19184
rect 22926 19000 22982 19009
rect 23124 18970 23152 19178
rect 22926 18935 22982 18944
rect 23112 18964 23164 18970
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22374 18592 22430 18601
rect 22374 18527 22430 18536
rect 22388 18426 22416 18527
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22466 18184 22522 18193
rect 22466 18119 22522 18128
rect 22480 17134 22508 18119
rect 22468 17128 22520 17134
rect 22374 17096 22430 17105
rect 22284 17060 22336 17066
rect 22468 17070 22520 17076
rect 22374 17031 22430 17040
rect 22284 17002 22336 17008
rect 22098 16824 22154 16833
rect 22098 16759 22154 16768
rect 22190 16688 22246 16697
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 22100 16652 22152 16658
rect 22296 16658 22324 17002
rect 22388 16658 22416 17031
rect 22480 16658 22508 17070
rect 22190 16623 22246 16632
rect 22284 16652 22336 16658
rect 22100 16594 22152 16600
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21822 16552 21878 16561
rect 21364 16448 21416 16454
rect 21744 16425 21772 16526
rect 21822 16487 21878 16496
rect 21364 16390 21416 16396
rect 21730 16416 21786 16425
rect 21376 13716 21404 16390
rect 21730 16351 21786 16360
rect 21456 16040 21508 16046
rect 21454 16008 21456 16017
rect 21548 16040 21600 16046
rect 21508 16008 21510 16017
rect 21732 16040 21784 16046
rect 21548 15982 21600 15988
rect 21638 16008 21694 16017
rect 21454 15943 21510 15952
rect 21468 15337 21496 15943
rect 21454 15328 21510 15337
rect 21454 15263 21510 15272
rect 21454 15192 21510 15201
rect 21454 15127 21510 15136
rect 21468 15026 21496 15127
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21468 13977 21496 14826
rect 21560 14249 21588 15982
rect 21732 15982 21784 15988
rect 21638 15943 21694 15952
rect 21652 15910 21680 15943
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21652 14958 21680 15098
rect 21744 15042 21772 15982
rect 21836 15473 21864 16487
rect 21822 15464 21878 15473
rect 21822 15399 21878 15408
rect 21744 15026 21864 15042
rect 21744 15020 21876 15026
rect 21744 15014 21824 15020
rect 21824 14962 21876 14968
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21652 14822 21680 14894
rect 21640 14816 21692 14822
rect 21744 14793 21772 14894
rect 21824 14816 21876 14822
rect 21640 14758 21692 14764
rect 21730 14784 21786 14793
rect 21546 14240 21602 14249
rect 21546 14175 21602 14184
rect 21560 14074 21588 14175
rect 21652 14074 21680 14758
rect 21824 14758 21876 14764
rect 21730 14719 21786 14728
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21836 13977 21864 14758
rect 21454 13968 21510 13977
rect 21822 13968 21878 13977
rect 21454 13903 21510 13912
rect 21732 13932 21784 13938
rect 21468 13870 21496 13903
rect 21822 13903 21878 13912
rect 21732 13874 21784 13880
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21376 13688 21588 13716
rect 21454 13424 21510 13433
rect 21192 13326 21220 13398
rect 21284 13382 21404 13410
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21086 12880 21142 12889
rect 21086 12815 21142 12824
rect 20994 12336 21050 12345
rect 20994 12271 21050 12280
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20902 11248 20958 11257
rect 20902 11183 20958 11192
rect 20904 11008 20956 11014
rect 21008 10985 21036 11834
rect 20904 10950 20956 10956
rect 20994 10976 21050 10985
rect 20916 10305 20944 10950
rect 20994 10911 21050 10920
rect 21008 10674 21036 10911
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 20902 10296 20958 10305
rect 21008 10266 21036 10610
rect 21100 10266 21128 12815
rect 21192 12306 21220 13262
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 20902 10231 20958 10240
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20732 10016 20852 10044
rect 20442 9888 20498 9897
rect 20442 9823 20498 9832
rect 20626 9888 20682 9897
rect 20626 9823 20682 9832
rect 20364 9646 20484 9674
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20364 8634 20392 9454
rect 20456 9178 20484 9646
rect 20536 9512 20588 9518
rect 20640 9500 20668 9823
rect 20588 9472 20668 9500
rect 20536 9454 20588 9460
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20548 9024 20576 9114
rect 20456 8996 20576 9024
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20352 8356 20404 8362
rect 20180 8316 20300 8344
rect 20076 8298 20128 8304
rect 19870 8188 20178 8197
rect 19870 8186 19876 8188
rect 19932 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20178 8188
rect 19932 8134 19934 8186
rect 20114 8134 20116 8186
rect 19870 8132 19876 8134
rect 19932 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20178 8134
rect 19870 8123 20178 8132
rect 19720 8078 19840 8106
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19720 6798 19748 8078
rect 20272 8072 20300 8316
rect 20352 8298 20404 8304
rect 20180 8044 20300 8072
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19812 7721 19840 7890
rect 19798 7712 19854 7721
rect 19798 7647 19854 7656
rect 19812 7342 19840 7647
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19904 7188 19932 7890
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 20088 7342 20116 7754
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 19812 7160 19932 7188
rect 20180 7188 20208 8044
rect 20364 7954 20392 8298
rect 20456 8022 20484 8996
rect 20640 8922 20668 9472
rect 20548 8906 20668 8922
rect 20536 8900 20668 8906
rect 20588 8894 20668 8900
rect 20536 8842 20588 8848
rect 20628 8832 20680 8838
rect 20626 8800 20628 8809
rect 20680 8800 20682 8809
rect 20626 8735 20682 8744
rect 20732 8430 20760 10016
rect 20916 9722 20944 10066
rect 20996 10056 21048 10062
rect 21048 10016 21128 10044
rect 20996 9998 21048 10004
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20996 9580 21048 9586
rect 20824 9217 20852 9551
rect 20996 9522 21048 9528
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20916 9353 20944 9386
rect 20902 9344 20958 9353
rect 20902 9279 20958 9288
rect 20810 9208 20866 9217
rect 20916 9178 20944 9279
rect 20810 9143 20866 9152
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20810 9072 20866 9081
rect 21008 9042 21036 9522
rect 20810 9007 20866 9016
rect 20996 9036 21048 9042
rect 20824 8634 20852 9007
rect 20996 8978 21048 8984
rect 21100 8906 21128 10016
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20904 8418 20956 8424
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 20352 7948 20404 7954
rect 20628 7948 20680 7954
rect 20352 7890 20404 7896
rect 20548 7908 20628 7936
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 7478 20300 7686
rect 20350 7576 20406 7585
rect 20456 7546 20484 7822
rect 20548 7818 20576 7908
rect 20628 7890 20680 7896
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20350 7511 20406 7520
rect 20444 7540 20496 7546
rect 20260 7472 20312 7478
rect 20260 7414 20312 7420
rect 20260 7336 20312 7342
rect 20364 7324 20392 7511
rect 20444 7482 20496 7488
rect 20312 7296 20392 7324
rect 20260 7278 20312 7284
rect 20180 7160 20300 7188
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19260 6662 19288 6734
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19210 6556 19518 6565
rect 19210 6554 19216 6556
rect 19272 6554 19296 6556
rect 19352 6554 19376 6556
rect 19432 6554 19456 6556
rect 19512 6554 19518 6556
rect 19272 6502 19274 6554
rect 19454 6502 19456 6554
rect 19210 6500 19216 6502
rect 19272 6500 19296 6502
rect 19352 6500 19376 6502
rect 19432 6500 19456 6502
rect 19512 6500 19518 6502
rect 19210 6491 19518 6500
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19168 6118 19196 6190
rect 19156 6112 19208 6118
rect 19444 6089 19472 6190
rect 19156 6054 19208 6060
rect 19430 6080 19486 6089
rect 19430 6015 19486 6024
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18878 5400 18934 5409
rect 18878 5335 18934 5344
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18800 4826 18828 5102
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18248 4214 18276 4626
rect 18236 4208 18288 4214
rect 18340 4185 18368 4626
rect 18236 4150 18288 4156
rect 18326 4176 18382 4185
rect 18326 4111 18382 4120
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18432 4010 18460 4694
rect 18616 4690 18644 4762
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18892 4486 18920 5102
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18984 4078 19012 5714
rect 19444 5710 19472 6015
rect 19340 5704 19392 5710
rect 19338 5672 19340 5681
rect 19432 5704 19484 5710
rect 19392 5672 19394 5681
rect 19064 5636 19116 5642
rect 19432 5646 19484 5652
rect 19338 5607 19394 5616
rect 19064 5578 19116 5584
rect 19076 5370 19104 5578
rect 19210 5468 19518 5477
rect 19210 5466 19216 5468
rect 19272 5466 19296 5468
rect 19352 5466 19376 5468
rect 19432 5466 19456 5468
rect 19512 5466 19518 5468
rect 19272 5414 19274 5466
rect 19454 5414 19456 5466
rect 19210 5412 19216 5414
rect 19272 5412 19296 5414
rect 19352 5412 19376 5414
rect 19432 5412 19456 5414
rect 19512 5412 19518 5414
rect 19210 5403 19518 5412
rect 19064 5364 19116 5370
rect 19628 5352 19656 6666
rect 19812 6644 19840 7160
rect 19870 7100 20178 7109
rect 19870 7098 19876 7100
rect 19932 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20178 7100
rect 19932 7046 19934 7098
rect 20114 7046 20116 7098
rect 19870 7044 19876 7046
rect 19932 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20178 7046
rect 19870 7035 20178 7044
rect 19890 6896 19946 6905
rect 19890 6831 19946 6840
rect 20166 6896 20222 6905
rect 20166 6831 20222 6840
rect 19064 5306 19116 5312
rect 19536 5324 19656 5352
rect 19720 6616 19840 6644
rect 19904 6633 19932 6831
rect 20180 6798 20208 6831
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 19890 6624 19946 6633
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4865 19104 5102
rect 19062 4856 19118 4865
rect 19062 4791 19118 4800
rect 19536 4570 19564 5324
rect 19720 4758 19748 6616
rect 19890 6559 19946 6568
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 19536 4542 19748 4570
rect 19536 4486 19564 4542
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19210 4380 19518 4389
rect 19210 4378 19216 4380
rect 19272 4378 19296 4380
rect 19352 4378 19376 4380
rect 19432 4378 19456 4380
rect 19512 4378 19518 4380
rect 19272 4326 19274 4378
rect 19454 4326 19456 4378
rect 19210 4324 19216 4326
rect 19272 4324 19296 4326
rect 19352 4324 19376 4326
rect 19432 4324 19456 4326
rect 19512 4324 19518 4326
rect 19210 4315 19518 4324
rect 19628 4146 19656 4422
rect 19720 4162 19748 4542
rect 19812 4264 19840 6394
rect 20088 6186 20116 6734
rect 20076 6180 20128 6186
rect 20076 6122 20128 6128
rect 20180 6118 20208 6734
rect 20272 6118 20300 7160
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20456 6458 20484 6802
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 19870 6012 20178 6021
rect 19870 6010 19876 6012
rect 19932 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20178 6012
rect 19932 5958 19934 6010
rect 20114 5958 20116 6010
rect 19870 5956 19876 5958
rect 19932 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20178 5958
rect 19870 5947 20178 5956
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 20088 5574 20116 5714
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20272 5166 20300 6054
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20364 5302 20392 5714
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 19870 4924 20178 4933
rect 19870 4922 19876 4924
rect 19932 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20178 4924
rect 19932 4870 19934 4922
rect 20114 4870 20116 4922
rect 19870 4868 19876 4870
rect 19932 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20178 4870
rect 19870 4859 20178 4868
rect 20364 4758 20392 5102
rect 19984 4752 20036 4758
rect 19984 4694 20036 4700
rect 20352 4752 20404 4758
rect 20352 4694 20404 4700
rect 19996 4282 20024 4694
rect 20548 4690 20576 7754
rect 20732 7750 20760 8230
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20640 7313 20668 7414
rect 20626 7304 20682 7313
rect 20626 7239 20682 7248
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 6866 20668 7142
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20732 6662 20760 7686
rect 20824 7546 20852 8366
rect 20904 8360 20956 8366
rect 20916 8090 20944 8360
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20812 7336 20864 7342
rect 20810 7304 20812 7313
rect 20864 7304 20866 7313
rect 20810 7239 20866 7248
rect 20916 6905 20944 7346
rect 21008 7342 21036 7890
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 20902 6896 20958 6905
rect 20902 6831 20958 6840
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20902 6624 20958 6633
rect 20640 6458 20668 6598
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 19984 4276 20036 4282
rect 19812 4236 19932 4264
rect 19720 4146 19840 4162
rect 19616 4140 19668 4146
rect 19720 4140 19852 4146
rect 19720 4134 19800 4140
rect 19616 4082 19668 4088
rect 19800 4082 19852 4088
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 19708 4072 19760 4078
rect 19904 4026 19932 4236
rect 19984 4218 20036 4224
rect 19760 4020 19932 4026
rect 19708 4014 19932 4020
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 19340 4004 19392 4010
rect 19720 3998 19932 4014
rect 19340 3946 19392 3952
rect 17684 3936 17736 3942
rect 16486 3904 16542 3913
rect 17684 3878 17736 3884
rect 16486 3839 16542 3848
rect 16500 3602 16528 3839
rect 19352 3738 19380 3946
rect 20548 3942 20576 4626
rect 20732 4554 20760 6598
rect 20902 6559 20958 6568
rect 20916 5817 20944 6559
rect 20902 5808 20958 5817
rect 20902 5743 20958 5752
rect 20902 5400 20958 5409
rect 20902 5335 20958 5344
rect 20916 5166 20944 5335
rect 20904 5160 20956 5166
rect 21008 5137 21036 7278
rect 21100 6186 21128 7686
rect 21192 7478 21220 11222
rect 21284 10742 21312 13262
rect 21376 11898 21404 13382
rect 21454 13359 21510 13368
rect 21468 12170 21496 13359
rect 21560 12889 21588 13688
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21546 12880 21602 12889
rect 21546 12815 21602 12824
rect 21652 12442 21680 13330
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21560 11744 21588 12378
rect 21744 11898 21772 13874
rect 21928 13394 21956 16594
rect 22112 16561 22140 16594
rect 22098 16552 22154 16561
rect 22020 16510 22098 16538
rect 22020 15978 22048 16510
rect 22098 16487 22154 16496
rect 22204 16250 22232 16623
rect 22284 16594 22336 16600
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22480 16538 22508 16594
rect 22388 16510 22508 16538
rect 22572 16522 22600 16594
rect 22560 16516 22612 16522
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22192 16244 22244 16250
rect 22192 16186 22244 16192
rect 22112 15978 22140 16186
rect 22284 16040 22336 16046
rect 22282 16008 22284 16017
rect 22336 16008 22338 16017
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 22100 15972 22152 15978
rect 22282 15943 22338 15952
rect 22100 15914 22152 15920
rect 22112 14872 22140 15914
rect 22388 15638 22416 16510
rect 22560 16458 22612 16464
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22480 16114 22508 16390
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22572 15994 22600 16186
rect 22480 15966 22600 15994
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22282 15192 22338 15201
rect 22282 15127 22338 15136
rect 22192 14884 22244 14890
rect 22112 14844 22192 14872
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12782 21956 13330
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 22020 12714 22048 13670
rect 22112 13530 22140 14844
rect 22192 14826 22244 14832
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22204 13954 22232 14554
rect 22296 14346 22324 15127
rect 22388 14958 22416 15574
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22296 14074 22324 14282
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22204 13926 22324 13954
rect 22190 13696 22246 13705
rect 22190 13631 22246 13640
rect 22204 13530 22232 13631
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22112 12850 22140 13330
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 22204 12889 22232 13126
rect 22190 12880 22246 12889
rect 22100 12844 22152 12850
rect 22190 12815 22246 12824
rect 22100 12786 22152 12792
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21640 11756 21692 11762
rect 21560 11716 21640 11744
rect 21640 11698 21692 11704
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21270 8528 21326 8537
rect 21270 8463 21326 8472
rect 21284 8430 21312 8463
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21192 7002 21220 7278
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21088 6180 21140 6186
rect 21088 6122 21140 6128
rect 21100 5302 21128 6122
rect 21192 5914 21220 6734
rect 21284 6361 21312 7958
rect 21270 6352 21326 6361
rect 21270 6287 21326 6296
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21284 5710 21312 6190
rect 21376 5914 21404 11630
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21468 10606 21496 11494
rect 21652 11286 21680 11698
rect 21836 11694 21864 12582
rect 22190 12336 22246 12345
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22008 12300 22060 12306
rect 22190 12271 22246 12280
rect 22008 12242 22060 12248
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21928 11540 21956 12242
rect 22020 11898 22048 12242
rect 22204 12238 22232 12271
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22112 11694 22140 12038
rect 22296 11898 22324 13926
rect 22388 13394 22416 14894
rect 22480 14822 22508 15966
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22466 14648 22522 14657
rect 22466 14583 22468 14592
rect 22520 14583 22522 14592
rect 22468 14554 22520 14560
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22480 13870 22508 14214
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22374 12608 22430 12617
rect 22374 12543 22430 12552
rect 22388 12374 22416 12543
rect 22376 12368 22428 12374
rect 22376 12310 22428 12316
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 21744 11512 21956 11540
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21454 10432 21510 10441
rect 21454 10367 21510 10376
rect 21468 9654 21496 10367
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21560 9194 21588 11086
rect 21640 10600 21692 10606
rect 21640 10542 21692 10548
rect 21652 10266 21680 10542
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21652 9926 21680 10066
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21468 9166 21588 9194
rect 21468 8344 21496 9166
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21560 8566 21588 8978
rect 21652 8956 21680 9522
rect 21744 9110 21772 11512
rect 22006 11112 22062 11121
rect 21916 11076 21968 11082
rect 22006 11047 22062 11056
rect 21916 11018 21968 11024
rect 21928 10674 21956 11018
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21836 9722 21864 10542
rect 21914 10024 21970 10033
rect 21914 9959 21970 9968
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21928 9518 21956 9959
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21824 9376 21876 9382
rect 21876 9336 21956 9364
rect 21824 9318 21876 9324
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21652 8928 21772 8956
rect 21836 8945 21864 8978
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21548 8560 21600 8566
rect 21652 8537 21680 8570
rect 21744 8566 21772 8928
rect 21822 8936 21878 8945
rect 21822 8871 21878 8880
rect 21732 8560 21784 8566
rect 21548 8502 21600 8508
rect 21638 8528 21694 8537
rect 21732 8502 21784 8508
rect 21638 8463 21694 8472
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21640 8356 21692 8362
rect 21468 8316 21640 8344
rect 21640 8298 21692 8304
rect 21744 8129 21772 8366
rect 21730 8120 21786 8129
rect 21640 8084 21692 8090
rect 21730 8055 21786 8064
rect 21640 8026 21692 8032
rect 21652 7818 21680 8026
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21836 7698 21864 8366
rect 21560 7670 21864 7698
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21468 6934 21496 7511
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 21560 6066 21588 7670
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21836 7342 21864 7482
rect 21732 7336 21784 7342
rect 21652 7296 21732 7324
rect 21652 6934 21680 7296
rect 21732 7278 21784 7284
rect 21824 7336 21876 7342
rect 21824 7278 21876 7284
rect 21730 7032 21786 7041
rect 21730 6967 21786 6976
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21744 6866 21772 6967
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21744 6662 21772 6802
rect 21928 6798 21956 9336
rect 22020 9042 22048 11047
rect 22112 10130 22140 11630
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22204 11121 22232 11154
rect 22190 11112 22246 11121
rect 22190 11047 22246 11056
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22204 10606 22232 10950
rect 22282 10840 22338 10849
rect 22282 10775 22284 10784
rect 22336 10775 22338 10784
rect 22284 10746 22336 10752
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22204 10198 22232 10542
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22282 9616 22338 9625
rect 22282 9551 22338 9560
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22020 8430 22048 8774
rect 22008 8424 22060 8430
rect 22112 8401 22140 9046
rect 22008 8366 22060 8372
rect 22098 8392 22154 8401
rect 22098 8327 22154 8336
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22098 8256 22154 8265
rect 22020 7954 22048 8230
rect 22098 8191 22154 8200
rect 22112 8090 22140 8191
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22112 6662 22140 7890
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 21928 6254 21956 6598
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 21916 6248 21968 6254
rect 21822 6216 21878 6225
rect 21916 6190 21968 6196
rect 21822 6151 21878 6160
rect 21468 6038 21588 6066
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21088 5296 21140 5302
rect 21088 5238 21140 5244
rect 20904 5102 20956 5108
rect 20994 5128 21050 5137
rect 20994 5063 21050 5072
rect 20810 4856 20866 4865
rect 20810 4791 20866 4800
rect 20824 4690 20852 4791
rect 21100 4758 21128 5238
rect 21468 5166 21496 6038
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21560 5370 21588 5714
rect 21652 5574 21680 5850
rect 21836 5778 21864 6151
rect 22020 5778 22048 6394
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20720 4548 20772 4554
rect 20720 4490 20772 4496
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20640 4146 20668 4218
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20732 4078 20760 4490
rect 20824 4214 20852 4626
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 19870 3836 20178 3845
rect 19870 3834 19876 3836
rect 19932 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20178 3836
rect 19932 3782 19934 3834
rect 20114 3782 20116 3834
rect 19870 3780 19876 3782
rect 19932 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20178 3782
rect 19870 3771 20178 3780
rect 20732 3738 20760 3878
rect 21284 3738 21312 4966
rect 21468 4729 21496 5102
rect 21744 4826 21772 5578
rect 22204 4826 22232 9454
rect 22296 8294 22324 9551
rect 22388 8634 22416 11630
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22388 8022 22416 8366
rect 22376 8016 22428 8022
rect 22376 7958 22428 7964
rect 22480 7392 22508 13670
rect 22572 12374 22600 15846
rect 22664 15706 22692 18702
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22756 17270 22784 18294
rect 22836 18080 22888 18086
rect 22836 18022 22888 18028
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22744 17128 22796 17134
rect 22742 17096 22744 17105
rect 22796 17096 22798 17105
rect 22742 17031 22798 17040
rect 22848 16697 22876 18022
rect 22940 16998 22968 18935
rect 23112 18906 23164 18912
rect 23296 18896 23348 18902
rect 23296 18838 23348 18844
rect 23112 18624 23164 18630
rect 23018 18592 23074 18601
rect 23112 18566 23164 18572
rect 23018 18527 23074 18536
rect 23032 17134 23060 18527
rect 23124 17241 23152 18566
rect 23204 18420 23256 18426
rect 23308 18408 23336 18838
rect 23400 18766 23428 19944
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23388 18420 23440 18426
rect 23308 18380 23388 18408
rect 23204 18362 23256 18368
rect 23388 18362 23440 18368
rect 23216 17785 23244 18362
rect 23584 18358 23612 19722
rect 23572 18352 23624 18358
rect 23386 18320 23442 18329
rect 23572 18294 23624 18300
rect 23386 18255 23442 18264
rect 23676 18272 23704 20810
rect 23952 20602 23980 21247
rect 24044 21010 24072 21286
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24136 20806 24164 21354
rect 24228 21146 24256 21354
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24216 20936 24268 20942
rect 24216 20878 24268 20884
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 24136 20466 24164 20742
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23756 19984 23808 19990
rect 23756 19926 23808 19932
rect 23768 19310 23796 19926
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23860 19514 23888 19790
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23768 18970 23796 19246
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23860 18873 23888 19246
rect 23846 18864 23902 18873
rect 23846 18799 23902 18808
rect 23952 18465 23980 19994
rect 24044 19514 24072 20334
rect 24136 19990 24164 20402
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 24228 19718 24256 20878
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 24228 19310 24256 19654
rect 24216 19304 24268 19310
rect 24216 19246 24268 19252
rect 24124 19236 24176 19242
rect 24124 19178 24176 19184
rect 24032 18896 24084 18902
rect 24136 18884 24164 19178
rect 24084 18856 24164 18884
rect 24032 18838 24084 18844
rect 24044 18766 24072 18838
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 23938 18456 23994 18465
rect 23938 18391 23994 18400
rect 23846 18320 23902 18329
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23202 17776 23258 17785
rect 23202 17711 23258 17720
rect 23110 17232 23166 17241
rect 23110 17167 23166 17176
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 22928 16992 22980 16998
rect 23124 16969 23152 17167
rect 22928 16934 22980 16940
rect 23110 16960 23166 16969
rect 23110 16895 23166 16904
rect 22834 16688 22890 16697
rect 22834 16623 22836 16632
rect 22888 16623 22890 16632
rect 22836 16594 22888 16600
rect 22928 16584 22980 16590
rect 22926 16552 22928 16561
rect 23020 16584 23072 16590
rect 22980 16552 22982 16561
rect 22836 16516 22888 16522
rect 23216 16561 23244 17711
rect 23020 16526 23072 16532
rect 23202 16552 23258 16561
rect 22926 16487 22982 16496
rect 22836 16458 22888 16464
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22664 15026 22692 15642
rect 22848 15434 22876 16458
rect 23032 16250 23060 16526
rect 23202 16487 23258 16496
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 22940 15706 22968 15914
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 23032 15609 23060 16050
rect 23018 15600 23074 15609
rect 23018 15535 23074 15544
rect 22836 15428 22888 15434
rect 22836 15370 22888 15376
rect 23124 15178 23152 16390
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23216 15910 23244 16186
rect 23204 15904 23256 15910
rect 23308 15892 23336 18158
rect 23400 17785 23428 18255
rect 23676 18244 23796 18272
rect 23846 18255 23902 18264
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23492 18057 23520 18090
rect 23478 18048 23534 18057
rect 23478 17983 23534 17992
rect 23480 17808 23532 17814
rect 23386 17776 23442 17785
rect 23480 17750 23532 17756
rect 23386 17711 23442 17720
rect 23388 17332 23440 17338
rect 23492 17320 23520 17750
rect 23440 17292 23520 17320
rect 23388 17274 23440 17280
rect 23386 17232 23442 17241
rect 23386 17167 23442 17176
rect 23480 17196 23532 17202
rect 23400 17066 23428 17167
rect 23480 17138 23532 17144
rect 23388 17060 23440 17066
rect 23388 17002 23440 17008
rect 23492 16454 23520 17138
rect 23572 17060 23624 17066
rect 23572 17002 23624 17008
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23400 16250 23428 16390
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23492 15994 23520 16390
rect 23584 16114 23612 17002
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23676 16046 23704 16759
rect 23768 16726 23796 18244
rect 23860 18222 23888 18255
rect 23952 18222 23980 18391
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23940 18216 23992 18222
rect 23940 18158 23992 18164
rect 24044 17882 24072 18702
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 23940 17672 23992 17678
rect 24136 17660 24164 18090
rect 24216 17876 24268 17882
rect 24216 17818 24268 17824
rect 23992 17632 24164 17660
rect 23940 17614 23992 17620
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23860 17270 23888 17478
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23952 17202 23980 17614
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 24044 17134 24072 17274
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 23756 16720 23808 16726
rect 23756 16662 23808 16668
rect 23860 16522 23888 17070
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23952 16402 23980 16594
rect 23860 16374 23980 16402
rect 23664 16040 23716 16046
rect 23492 15966 23612 15994
rect 23664 15982 23716 15988
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23584 15910 23612 15966
rect 23480 15904 23532 15910
rect 23308 15864 23428 15892
rect 23204 15846 23256 15852
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22940 15150 23152 15178
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22756 14958 22784 15098
rect 22744 14952 22796 14958
rect 22650 14920 22706 14929
rect 22744 14894 22796 14900
rect 22650 14855 22706 14864
rect 22664 13410 22692 14855
rect 22756 13977 22784 14894
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22848 14074 22876 14214
rect 22836 14068 22888 14074
rect 22836 14010 22888 14016
rect 22742 13968 22798 13977
rect 22742 13903 22798 13912
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22756 13530 22784 13670
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22664 13382 22784 13410
rect 22650 13288 22706 13297
rect 22650 13223 22706 13232
rect 22664 12986 22692 13223
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22650 12880 22706 12889
rect 22650 12815 22652 12824
rect 22704 12815 22706 12824
rect 22652 12786 22704 12792
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22756 12306 22784 13382
rect 22848 13326 22876 13670
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22572 11354 22600 11630
rect 22652 11552 22704 11558
rect 22756 11529 22784 11630
rect 22652 11494 22704 11500
rect 22742 11520 22798 11529
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 10198 22600 10406
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22560 10056 22612 10062
rect 22664 10033 22692 11494
rect 22742 11455 22798 11464
rect 22742 11248 22798 11257
rect 22848 11218 22876 12786
rect 22940 12442 22968 15150
rect 23112 14952 23164 14958
rect 23112 14894 23164 14900
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 23032 14482 23060 14826
rect 23020 14476 23072 14482
rect 23020 14418 23072 14424
rect 23032 14385 23060 14418
rect 23124 14396 23152 14894
rect 23216 14793 23244 15506
rect 23400 14958 23428 15864
rect 23480 15846 23532 15852
rect 23572 15904 23624 15910
rect 23624 15864 23704 15892
rect 23572 15846 23624 15852
rect 23492 15638 23520 15846
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23492 15502 23520 15574
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 23202 14784 23258 14793
rect 23202 14719 23258 14728
rect 23204 14408 23256 14414
rect 23018 14376 23074 14385
rect 23124 14368 23204 14396
rect 23204 14350 23256 14356
rect 23018 14311 23074 14320
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22742 11183 22798 11192
rect 22836 11212 22888 11218
rect 22756 10577 22784 11183
rect 22836 11154 22888 11160
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22848 10606 22876 10950
rect 22836 10600 22888 10606
rect 22742 10568 22798 10577
rect 22836 10542 22888 10548
rect 22742 10503 22798 10512
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22560 9998 22612 10004
rect 22650 10024 22706 10033
rect 22572 7585 22600 9998
rect 22650 9959 22706 9968
rect 22756 9722 22784 10406
rect 22848 9994 22876 10542
rect 22836 9988 22888 9994
rect 22836 9930 22888 9936
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22940 9518 22968 12242
rect 23032 11694 23060 14311
rect 23400 13977 23428 14894
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23202 13968 23258 13977
rect 23202 13903 23258 13912
rect 23386 13968 23442 13977
rect 23386 13903 23442 13912
rect 23110 13832 23166 13841
rect 23110 13767 23166 13776
rect 23124 13530 23152 13767
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23124 12306 23152 12922
rect 23216 12850 23244 13903
rect 23400 13802 23428 13903
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23296 12300 23348 12306
rect 23296 12242 23348 12248
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 23124 11529 23152 12038
rect 23110 11520 23166 11529
rect 23110 11455 23166 11464
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23032 10810 23060 11290
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23018 10296 23074 10305
rect 23018 10231 23074 10240
rect 23032 10130 23060 10231
rect 23112 10192 23164 10198
rect 23112 10134 23164 10140
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23124 10033 23152 10134
rect 23110 10024 23166 10033
rect 23110 9959 23166 9968
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 22836 9444 22888 9450
rect 22836 9386 22888 9392
rect 22650 9344 22706 9353
rect 22650 9279 22706 9288
rect 22664 8430 22692 9279
rect 22848 9178 22876 9386
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22940 9081 22968 9318
rect 23032 9178 23060 9454
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 22926 9072 22982 9081
rect 23124 9058 23152 9590
rect 23032 9042 23152 9058
rect 22926 9007 22982 9016
rect 23020 9036 23152 9042
rect 23072 9030 23152 9036
rect 23020 8978 23072 8984
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22650 8256 22706 8265
rect 22650 8191 22706 8200
rect 22664 7954 22692 8191
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22756 7698 22784 8502
rect 22836 8424 22888 8430
rect 22836 8366 22888 8372
rect 22848 7818 22876 8366
rect 22940 8129 22968 8910
rect 23032 8566 23060 8978
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23124 8634 23152 8910
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23112 8356 23164 8362
rect 23112 8298 23164 8304
rect 22926 8120 22982 8129
rect 22926 8055 22982 8064
rect 22836 7812 22888 7818
rect 22836 7754 22888 7760
rect 22558 7576 22614 7585
rect 22558 7511 22614 7520
rect 22388 7364 22508 7392
rect 22284 7336 22336 7342
rect 22388 7324 22416 7364
rect 22336 7296 22416 7324
rect 22284 7278 22336 7284
rect 22468 7268 22520 7274
rect 22572 7256 22600 7511
rect 22520 7228 22600 7256
rect 22468 7210 22520 7216
rect 22558 7032 22614 7041
rect 22558 6967 22614 6976
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22376 6860 22428 6866
rect 22376 6802 22428 6808
rect 22296 6458 22324 6802
rect 22388 6497 22416 6802
rect 22374 6488 22430 6497
rect 22284 6452 22336 6458
rect 22374 6423 22430 6432
rect 22284 6394 22336 6400
rect 22572 6390 22600 6967
rect 22664 6934 22692 7686
rect 22756 7670 22968 7698
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22744 7268 22796 7274
rect 22744 7210 22796 7216
rect 22652 6928 22704 6934
rect 22756 6905 22784 7210
rect 22652 6870 22704 6876
rect 22742 6896 22798 6905
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 21454 4720 21510 4729
rect 21454 4655 21510 4664
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21560 4078 21588 4558
rect 21822 4176 21878 4185
rect 21822 4111 21878 4120
rect 21836 4078 21864 4111
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 19210 3292 19518 3301
rect 19210 3290 19216 3292
rect 19272 3290 19296 3292
rect 19352 3290 19376 3292
rect 19432 3290 19456 3292
rect 19512 3290 19518 3292
rect 19272 3238 19274 3290
rect 19454 3238 19456 3290
rect 19210 3236 19216 3238
rect 19272 3236 19296 3238
rect 19352 3236 19376 3238
rect 19432 3236 19456 3238
rect 19512 3236 19518 3238
rect 19210 3227 19518 3236
rect 21284 2961 21312 3674
rect 21376 3602 21404 3946
rect 21836 3942 21864 4014
rect 22296 4010 22324 5714
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 22480 4078 22508 5510
rect 22664 5166 22692 6870
rect 22742 6831 22798 6840
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22756 6118 22784 6734
rect 22848 6730 22876 7278
rect 22836 6724 22888 6730
rect 22836 6666 22888 6672
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22652 5160 22704 5166
rect 22652 5102 22704 5108
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22756 4282 22784 4626
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22848 4214 22876 4626
rect 22940 4214 22968 7670
rect 23018 7576 23074 7585
rect 23018 7511 23074 7520
rect 23032 7002 23060 7511
rect 23020 6996 23072 7002
rect 23020 6938 23072 6944
rect 23032 6730 23060 6938
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 23124 5234 23152 8298
rect 23216 8090 23244 12242
rect 23308 11762 23336 12242
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23308 10538 23336 10746
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23294 10432 23350 10441
rect 23294 10367 23350 10376
rect 23308 10130 23336 10367
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23294 9208 23350 9217
rect 23294 9143 23350 9152
rect 23308 9042 23336 9143
rect 23296 9036 23348 9042
rect 23296 8978 23348 8984
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23308 8265 23336 8434
rect 23400 8412 23428 12378
rect 23492 11354 23520 14214
rect 23584 14113 23612 15030
rect 23676 14482 23704 15864
rect 23768 15638 23796 15982
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23860 15484 23888 16374
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 23952 15570 23980 15914
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23768 15456 23888 15484
rect 23768 15162 23796 15456
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23768 14929 23796 15098
rect 23754 14920 23810 14929
rect 23754 14855 23810 14864
rect 23860 14793 23888 15302
rect 24044 15201 24072 17070
rect 24136 16046 24164 17478
rect 24228 16522 24256 17818
rect 24320 16726 24348 21286
rect 24780 20942 24808 21830
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24582 20360 24638 20369
rect 24582 20295 24638 20304
rect 24676 20324 24728 20330
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24412 19310 24440 19790
rect 24596 19689 24624 20295
rect 24676 20266 24728 20272
rect 24582 19680 24638 19689
rect 24582 19615 24638 19624
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24504 18358 24532 18702
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24596 18222 24624 19615
rect 24688 18290 24716 20266
rect 24872 19990 24900 21490
rect 24860 19984 24912 19990
rect 24780 19944 24860 19972
rect 24780 19242 24808 19944
rect 24860 19926 24912 19932
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25056 19310 25084 19722
rect 25240 19310 25268 21558
rect 26056 21480 26108 21486
rect 26252 21457 26280 21898
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 26056 21422 26108 21428
rect 26238 21448 26294 21457
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25412 20460 25464 20466
rect 25412 20402 25464 20408
rect 25318 19952 25374 19961
rect 25318 19887 25374 19896
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 24768 19236 24820 19242
rect 24768 19178 24820 19184
rect 24872 18698 24900 19246
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24964 18698 24992 19110
rect 25056 18834 25084 19246
rect 25332 19174 25360 19887
rect 25424 19514 25452 20402
rect 25688 19712 25740 19718
rect 25688 19654 25740 19660
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25700 19310 25728 19654
rect 25792 19310 25820 20878
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25976 20602 26004 20810
rect 25964 20596 26016 20602
rect 25964 20538 26016 20544
rect 26068 20330 26096 21422
rect 26148 21412 26200 21418
rect 26238 21383 26294 21392
rect 26148 21354 26200 21360
rect 26160 20777 26188 21354
rect 26344 20806 26372 21490
rect 26436 21162 26464 21626
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 26436 21134 26556 21162
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26332 20800 26384 20806
rect 26146 20768 26202 20777
rect 26332 20742 26384 20748
rect 26146 20703 26202 20712
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26056 20324 26108 20330
rect 26056 20266 26108 20272
rect 25962 19816 26018 19825
rect 25962 19751 26018 19760
rect 25870 19408 25926 19417
rect 25870 19343 25926 19352
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25228 18896 25280 18902
rect 25226 18864 25228 18873
rect 25424 18873 25452 19246
rect 25884 18970 25912 19343
rect 25976 19310 26004 19751
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25872 18964 25924 18970
rect 25872 18906 25924 18912
rect 25280 18864 25282 18873
rect 25044 18828 25096 18834
rect 25226 18799 25282 18808
rect 25410 18864 25466 18873
rect 25410 18799 25466 18808
rect 25044 18770 25096 18776
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25962 18728 26018 18737
rect 24860 18692 24912 18698
rect 24860 18634 24912 18640
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24412 17882 24440 18158
rect 24964 18086 24992 18634
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25148 18154 25176 18566
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24398 17776 24454 17785
rect 25148 17746 25176 18090
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 24398 17711 24454 17720
rect 25136 17740 25188 17746
rect 24412 17678 24440 17711
rect 25136 17682 25188 17688
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24308 16720 24360 16726
rect 24308 16662 24360 16668
rect 24412 16590 24440 17614
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24768 17332 24820 17338
rect 24820 17292 24900 17320
rect 24768 17274 24820 17280
rect 24766 17232 24822 17241
rect 24766 17167 24822 17176
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24490 16824 24546 16833
rect 24490 16759 24546 16768
rect 24504 16658 24532 16759
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 24306 16144 24362 16153
rect 24306 16079 24308 16088
rect 24360 16079 24362 16088
rect 24308 16050 24360 16056
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24030 15192 24086 15201
rect 24030 15127 24032 15136
rect 24084 15127 24086 15136
rect 24032 15098 24084 15104
rect 23940 14816 23992 14822
rect 23846 14784 23902 14793
rect 23940 14758 23992 14764
rect 23846 14719 23902 14728
rect 23754 14648 23810 14657
rect 23754 14583 23810 14592
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23570 14104 23626 14113
rect 23570 14039 23626 14048
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23584 12306 23612 13806
rect 23676 13802 23704 14418
rect 23664 13796 23716 13802
rect 23664 13738 23716 13744
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23676 12617 23704 13330
rect 23662 12608 23718 12617
rect 23662 12543 23718 12552
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23478 10568 23534 10577
rect 23478 10503 23534 10512
rect 23492 9761 23520 10503
rect 23584 9926 23612 12038
rect 23676 10577 23704 12543
rect 23662 10568 23718 10577
rect 23662 10503 23718 10512
rect 23768 10130 23796 14583
rect 23860 11286 23888 14719
rect 23952 14074 23980 14758
rect 24030 14512 24086 14521
rect 24030 14447 24032 14456
rect 24084 14447 24086 14456
rect 24032 14418 24084 14424
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 24044 13394 24072 14418
rect 24136 14006 24164 15506
rect 24228 14550 24256 15982
rect 24412 15688 24440 16526
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24596 15881 24624 15982
rect 24582 15872 24638 15881
rect 24582 15807 24638 15816
rect 24320 15660 24440 15688
rect 24584 15700 24636 15706
rect 24320 15609 24348 15660
rect 24584 15642 24636 15648
rect 24306 15600 24362 15609
rect 24596 15570 24624 15642
rect 24306 15535 24362 15544
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24320 14958 24348 15302
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24216 14544 24268 14550
rect 24216 14486 24268 14492
rect 24306 14512 24362 14521
rect 24306 14447 24308 14456
rect 24360 14447 24362 14456
rect 24308 14418 24360 14424
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24122 13696 24178 13705
rect 24122 13631 24178 13640
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24044 12866 24072 13194
rect 23952 12838 24072 12866
rect 23952 11694 23980 12838
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 24044 12442 24072 12718
rect 24136 12696 24164 13631
rect 24228 13569 24256 14214
rect 24214 13560 24270 13569
rect 24214 13495 24270 13504
rect 24228 13326 24256 13495
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24216 13184 24268 13190
rect 24214 13152 24216 13161
rect 24308 13184 24360 13190
rect 24268 13152 24270 13161
rect 24308 13126 24360 13132
rect 24214 13087 24270 13096
rect 24320 12714 24348 13126
rect 24216 12708 24268 12714
rect 24136 12668 24216 12696
rect 24216 12650 24268 12656
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24216 12368 24268 12374
rect 24216 12310 24268 12316
rect 24030 12200 24086 12209
rect 24030 12135 24086 12144
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23938 11520 23994 11529
rect 23938 11455 23994 11464
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 23848 11144 23900 11150
rect 23952 11132 23980 11455
rect 24044 11354 24072 12135
rect 24228 11830 24256 12310
rect 24412 11898 24440 15506
rect 24688 15502 24716 16934
rect 24780 16153 24808 17167
rect 24872 16946 24900 17292
rect 24964 17202 24992 17478
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24872 16918 24992 16946
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24872 16697 24900 16730
rect 24858 16688 24914 16697
rect 24964 16658 24992 16918
rect 24858 16623 24914 16632
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 25056 16250 25084 17614
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 16590 25176 17546
rect 25240 17513 25268 18022
rect 25424 17785 25452 18702
rect 25516 17921 25544 18702
rect 25962 18663 26018 18672
rect 26068 18714 26096 20266
rect 26146 20088 26202 20097
rect 26146 20023 26202 20032
rect 26160 19145 26188 20023
rect 26252 19718 26280 20334
rect 26344 19922 26372 20742
rect 26436 20233 26464 20946
rect 26528 20602 26556 21134
rect 26620 20806 26648 21286
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26528 20398 26556 20538
rect 26896 20482 26924 21966
rect 27988 21956 28040 21962
rect 27988 21898 28040 21904
rect 30932 21956 30984 21962
rect 30932 21898 30984 21904
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 26984 21788 27292 21797
rect 26984 21786 26990 21788
rect 27046 21786 27070 21788
rect 27126 21786 27150 21788
rect 27206 21786 27230 21788
rect 27286 21786 27292 21788
rect 27046 21734 27048 21786
rect 27228 21734 27230 21786
rect 26984 21732 26990 21734
rect 27046 21732 27070 21734
rect 27126 21732 27150 21734
rect 27206 21732 27230 21734
rect 27286 21732 27292 21734
rect 26984 21723 27292 21732
rect 27540 21010 27568 21830
rect 28000 21418 28028 21898
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 28356 21616 28408 21622
rect 28356 21558 28408 21564
rect 27988 21412 28040 21418
rect 27988 21354 28040 21360
rect 28264 21412 28316 21418
rect 28264 21354 28316 21360
rect 27644 21244 27952 21253
rect 27644 21242 27650 21244
rect 27706 21242 27730 21244
rect 27786 21242 27810 21244
rect 27866 21242 27890 21244
rect 27946 21242 27952 21244
rect 27706 21190 27708 21242
rect 27888 21190 27890 21242
rect 27644 21188 27650 21190
rect 27706 21188 27730 21190
rect 27786 21188 27810 21190
rect 27866 21188 27890 21190
rect 27946 21188 27952 21190
rect 27644 21179 27952 21188
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27356 20806 27384 20946
rect 27344 20800 27396 20806
rect 27344 20742 27396 20748
rect 26984 20700 27292 20709
rect 26984 20698 26990 20700
rect 27046 20698 27070 20700
rect 27126 20698 27150 20700
rect 27206 20698 27230 20700
rect 27286 20698 27292 20700
rect 27046 20646 27048 20698
rect 27228 20646 27230 20698
rect 26984 20644 26990 20646
rect 27046 20644 27070 20646
rect 27126 20644 27150 20646
rect 27206 20644 27230 20646
rect 27286 20644 27292 20646
rect 26984 20635 27292 20644
rect 27632 20505 27660 20946
rect 28000 20890 28028 21354
rect 28080 21344 28132 21350
rect 28080 21286 28132 21292
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 28092 21146 28120 21286
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 28078 20904 28134 20913
rect 28000 20862 28078 20890
rect 28078 20839 28134 20848
rect 27618 20496 27674 20505
rect 26896 20454 27108 20482
rect 26516 20392 26568 20398
rect 26884 20392 26936 20398
rect 26516 20334 26568 20340
rect 26606 20360 26662 20369
rect 26884 20334 26936 20340
rect 26606 20295 26662 20304
rect 26422 20224 26478 20233
rect 26422 20159 26478 20168
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26240 19712 26292 19718
rect 26240 19654 26292 19660
rect 26330 19680 26386 19689
rect 26330 19615 26386 19624
rect 26344 19310 26372 19615
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 26146 19136 26202 19145
rect 26146 19071 26202 19080
rect 26252 19009 26280 19178
rect 26238 19000 26294 19009
rect 26238 18935 26294 18944
rect 26436 18902 26464 20159
rect 26620 19689 26648 20295
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26804 19854 26832 20198
rect 26896 20058 26924 20334
rect 26976 20324 27028 20330
rect 26976 20266 27028 20272
rect 26988 20058 27016 20266
rect 26884 20052 26936 20058
rect 26884 19994 26936 20000
rect 26976 20052 27028 20058
rect 26976 19994 27028 20000
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26606 19680 26662 19689
rect 26606 19615 26662 19624
rect 26712 19514 26740 19790
rect 26700 19508 26752 19514
rect 26700 19450 26752 19456
rect 26804 19242 26832 19790
rect 27080 19768 27108 20454
rect 27160 20460 27212 20466
rect 27618 20431 27674 20440
rect 27160 20402 27212 20408
rect 27172 20097 27200 20402
rect 27632 20398 27660 20431
rect 27344 20392 27396 20398
rect 27620 20392 27672 20398
rect 27396 20352 27476 20380
rect 27344 20334 27396 20340
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27158 20088 27214 20097
rect 27158 20023 27214 20032
rect 26896 19740 27108 19768
rect 26792 19236 26844 19242
rect 26792 19178 26844 19184
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26424 18760 26476 18766
rect 26068 18686 26372 18714
rect 26424 18702 26476 18708
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25502 17912 25558 17921
rect 25558 17870 25636 17898
rect 25502 17847 25558 17856
rect 25410 17776 25466 17785
rect 25410 17711 25466 17720
rect 25318 17640 25374 17649
rect 25318 17575 25374 17584
rect 25504 17604 25556 17610
rect 25226 17504 25282 17513
rect 25226 17439 25282 17448
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24766 16144 24822 16153
rect 24766 16079 24822 16088
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 25044 16108 25096 16114
rect 25148 16096 25176 16526
rect 25096 16068 25176 16096
rect 25044 16050 25096 16056
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24780 15706 24808 15982
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24766 15600 24822 15609
rect 24766 15535 24822 15544
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 24596 14958 24624 15370
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24504 13841 24532 14894
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24596 14278 24624 14418
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24490 13832 24546 13841
rect 24490 13767 24546 13776
rect 24492 13388 24544 13394
rect 24492 13330 24544 13336
rect 24504 13297 24532 13330
rect 24490 13288 24546 13297
rect 24490 13223 24546 13232
rect 24490 13016 24546 13025
rect 24490 12951 24546 12960
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24136 11558 24164 11698
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24124 11280 24176 11286
rect 24030 11248 24086 11257
rect 24124 11222 24176 11228
rect 24030 11183 24086 11192
rect 23900 11104 23980 11132
rect 23848 11086 23900 11092
rect 24044 11082 24072 11183
rect 24032 11076 24084 11082
rect 24032 11018 24084 11024
rect 24136 10962 24164 11222
rect 23952 10934 24164 10962
rect 23848 10260 23900 10266
rect 23952 10248 23980 10934
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24044 10266 24072 10746
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 23900 10220 23980 10248
rect 24032 10260 24084 10266
rect 23848 10202 23900 10208
rect 24032 10202 24084 10208
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23478 9752 23534 9761
rect 23478 9687 23534 9696
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23572 9512 23624 9518
rect 23572 9454 23624 9460
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23492 8838 23520 9114
rect 23584 9042 23612 9454
rect 23664 9444 23716 9450
rect 23664 9386 23716 9392
rect 23676 9110 23704 9386
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23480 8424 23532 8430
rect 23400 8384 23480 8412
rect 23532 8384 23612 8412
rect 23480 8366 23532 8372
rect 23294 8256 23350 8265
rect 23294 8191 23350 8200
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23216 7410 23244 7482
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22836 4004 22888 4010
rect 22940 3992 22968 4150
rect 23216 4078 23244 6598
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 22888 3964 22968 3992
rect 22836 3946 22888 3952
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3670 22508 3878
rect 22468 3664 22520 3670
rect 22468 3606 22520 3612
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21270 2952 21326 2961
rect 21270 2887 21326 2896
rect 23308 2774 23336 8191
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23400 7954 23428 8026
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23400 7002 23428 7890
rect 23492 7002 23520 7890
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23400 6882 23428 6938
rect 23400 6854 23520 6882
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23400 6662 23428 6734
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23492 6390 23520 6854
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 23584 5642 23612 8384
rect 23676 7954 23704 8910
rect 23768 8809 23796 9658
rect 23952 9489 23980 9862
rect 23938 9480 23994 9489
rect 23938 9415 23994 9424
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 9110 23888 9318
rect 23848 9104 23900 9110
rect 23848 9046 23900 9052
rect 23754 8800 23810 8809
rect 23754 8735 23810 8744
rect 23754 8528 23810 8537
rect 23754 8463 23810 8472
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23768 7834 23796 8463
rect 23846 8392 23902 8401
rect 23846 8327 23848 8336
rect 23900 8327 23902 8336
rect 23848 8298 23900 8304
rect 23676 7806 23796 7834
rect 23848 7812 23900 7818
rect 23676 6866 23704 7806
rect 23848 7754 23900 7760
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23768 6769 23796 7686
rect 23860 7546 23888 7754
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23754 6760 23810 6769
rect 23664 6724 23716 6730
rect 23754 6695 23810 6704
rect 23664 6666 23716 6672
rect 23676 6633 23704 6666
rect 23662 6624 23718 6633
rect 23662 6559 23718 6568
rect 23662 6352 23718 6361
rect 23662 6287 23718 6296
rect 23676 5953 23704 6287
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23662 5944 23718 5953
rect 23662 5879 23718 5888
rect 23572 5636 23624 5642
rect 23572 5578 23624 5584
rect 23768 5574 23796 6190
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23768 5302 23796 5510
rect 23756 5296 23808 5302
rect 23756 5238 23808 5244
rect 23860 3505 23888 6054
rect 23952 5370 23980 9415
rect 24030 9344 24086 9353
rect 24030 9279 24086 9288
rect 24044 9042 24072 9279
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 24030 8256 24086 8265
rect 24030 8191 24086 8200
rect 24044 8090 24072 8191
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24136 7993 24164 10542
rect 24228 10198 24256 11766
rect 24504 11694 24532 12951
rect 24596 12782 24624 13942
rect 24688 13818 24716 15438
rect 24780 15337 24808 15535
rect 24872 15502 24900 16050
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24766 15328 24822 15337
rect 24766 15263 24822 15272
rect 24872 15178 24900 15438
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24780 15150 24900 15178
rect 24780 14793 24808 15150
rect 24964 15026 24992 15302
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 24860 14884 24912 14890
rect 24912 14844 24992 14872
rect 24860 14826 24912 14832
rect 24766 14784 24822 14793
rect 24766 14719 24822 14728
rect 24964 14346 24992 14844
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24780 13938 24808 14214
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24688 13790 24808 13818
rect 24674 13560 24730 13569
rect 24674 13495 24730 13504
rect 24688 13258 24716 13495
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24674 13152 24730 13161
rect 24674 13087 24730 13096
rect 24688 12850 24716 13087
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 24584 12776 24636 12782
rect 24584 12718 24636 12724
rect 24596 12345 24624 12718
rect 24582 12336 24638 12345
rect 24582 12271 24638 12280
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 24320 11354 24348 11562
rect 24492 11552 24544 11558
rect 24398 11520 24454 11529
rect 24454 11500 24492 11506
rect 24454 11494 24544 11500
rect 24454 11478 24532 11494
rect 24398 11455 24454 11464
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24320 10538 24348 10950
rect 24412 10606 24440 11086
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 24320 10198 24348 10474
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24308 10192 24360 10198
rect 24308 10134 24360 10140
rect 24216 9512 24268 9518
rect 24214 9480 24216 9489
rect 24268 9480 24270 9489
rect 24214 9415 24270 9424
rect 24214 9208 24270 9217
rect 24214 9143 24270 9152
rect 24228 9042 24256 9143
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24320 8242 24348 10134
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24412 8906 24440 9998
rect 24504 9625 24532 11478
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24596 10606 24624 11290
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24490 9616 24546 9625
rect 24490 9551 24546 9560
rect 24504 9518 24532 9551
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24504 8809 24532 8978
rect 24490 8800 24546 8809
rect 24490 8735 24546 8744
rect 24398 8664 24454 8673
rect 24398 8599 24454 8608
rect 24412 8430 24440 8599
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24504 8242 24532 8735
rect 24596 8634 24624 10542
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24228 8214 24348 8242
rect 24412 8214 24532 8242
rect 24122 7984 24178 7993
rect 24032 7948 24084 7954
rect 24122 7919 24178 7928
rect 24032 7890 24084 7896
rect 24044 7342 24072 7890
rect 24124 7472 24176 7478
rect 24124 7414 24176 7420
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24044 6780 24072 7278
rect 24136 6934 24164 7414
rect 24228 7177 24256 8214
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24214 7168 24270 7177
rect 24214 7103 24270 7112
rect 24124 6928 24176 6934
rect 24124 6870 24176 6876
rect 24044 6752 24164 6780
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24044 6361 24072 6394
rect 24030 6352 24086 6361
rect 24030 6287 24086 6296
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24044 5817 24072 6054
rect 24030 5808 24086 5817
rect 24030 5743 24086 5752
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23952 4690 23980 5306
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 24044 3942 24072 5646
rect 24136 5302 24164 6752
rect 24228 6186 24256 7103
rect 24320 6730 24348 8026
rect 24412 7478 24440 8214
rect 24490 8120 24546 8129
rect 24596 8090 24624 8366
rect 24490 8055 24546 8064
rect 24584 8084 24636 8090
rect 24504 7954 24532 8055
rect 24584 8026 24636 8032
rect 24582 7984 24638 7993
rect 24492 7948 24544 7954
rect 24688 7954 24716 12786
rect 24780 11286 24808 13790
rect 24872 12102 24900 14214
rect 24964 13705 24992 14282
rect 24950 13696 25006 13705
rect 24950 13631 25006 13640
rect 25056 13546 25084 15914
rect 25148 15026 25176 16068
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 25240 14929 25268 17439
rect 25332 16658 25360 17575
rect 25504 17546 25556 17552
rect 25410 16824 25466 16833
rect 25410 16759 25466 16768
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25332 15502 25360 16594
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25332 15162 25360 15302
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 25226 14920 25282 14929
rect 25136 14884 25188 14890
rect 25226 14855 25282 14864
rect 25136 14826 25188 14832
rect 25148 14226 25176 14826
rect 25424 14822 25452 16759
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25332 14550 25360 14758
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25148 14198 25268 14226
rect 25134 14104 25190 14113
rect 25134 14039 25190 14048
rect 25148 13802 25176 14039
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 24964 13518 25084 13546
rect 24964 13394 24992 13518
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24964 13025 24992 13330
rect 24950 13016 25006 13025
rect 24950 12951 25006 12960
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24950 12064 25006 12073
rect 24950 11999 25006 12008
rect 24964 11762 24992 11999
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24952 11212 25004 11218
rect 24952 11154 25004 11160
rect 24964 10849 24992 11154
rect 24950 10840 25006 10849
rect 24950 10775 25006 10784
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24768 10056 24820 10062
rect 24820 10004 24900 10010
rect 24768 9998 24900 10004
rect 24780 9982 24900 9998
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9518 24808 9862
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24872 9450 24900 9982
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24872 9092 24900 9386
rect 24964 9382 24992 10542
rect 25056 10266 25084 13398
rect 25148 13326 25176 13738
rect 25240 13569 25268 14198
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25332 13841 25360 14010
rect 25412 13864 25464 13870
rect 25318 13832 25374 13841
rect 25412 13806 25464 13812
rect 25318 13767 25374 13776
rect 25226 13560 25282 13569
rect 25226 13495 25282 13504
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25332 13433 25360 13466
rect 25318 13424 25374 13433
rect 25424 13394 25452 13806
rect 25516 13734 25544 17546
rect 25608 17105 25636 17870
rect 25884 17814 25912 18022
rect 25872 17808 25924 17814
rect 25872 17750 25924 17756
rect 25872 17672 25924 17678
rect 25976 17649 26004 18663
rect 25872 17614 25924 17620
rect 25962 17640 26018 17649
rect 25884 17184 25912 17614
rect 25962 17575 26018 17584
rect 25962 17504 26018 17513
rect 25962 17439 26018 17448
rect 25976 17338 26004 17439
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25884 17156 26004 17184
rect 25594 17096 25650 17105
rect 25594 17031 25650 17040
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 16522 25636 16934
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25596 16516 25648 16522
rect 25596 16458 25648 16464
rect 25686 16416 25742 16425
rect 25686 16351 25742 16360
rect 25700 16182 25728 16351
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25688 15972 25740 15978
rect 25688 15914 25740 15920
rect 25596 15564 25648 15570
rect 25596 15506 25648 15512
rect 25608 14890 25636 15506
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25608 14657 25636 14826
rect 25594 14648 25650 14657
rect 25594 14583 25650 14592
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25608 14074 25636 14350
rect 25700 14278 25728 15914
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25700 14006 25728 14214
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25504 13728 25556 13734
rect 25504 13670 25556 13676
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25516 13530 25544 13670
rect 25608 13530 25636 13670
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25318 13359 25374 13368
rect 25412 13388 25464 13394
rect 25412 13330 25464 13336
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25134 13016 25190 13025
rect 25134 12951 25190 12960
rect 25148 12714 25176 12951
rect 25136 12708 25188 12714
rect 25136 12650 25188 12656
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 25148 11393 25176 12242
rect 25318 11792 25374 11801
rect 25318 11727 25374 11736
rect 25332 11694 25360 11727
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25424 11529 25452 13330
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25516 12073 25544 12242
rect 25596 12096 25648 12102
rect 25502 12064 25558 12073
rect 25596 12038 25648 12044
rect 25502 11999 25558 12008
rect 25504 11824 25556 11830
rect 25504 11766 25556 11772
rect 25516 11694 25544 11766
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25504 11552 25556 11558
rect 25410 11520 25466 11529
rect 25504 11494 25556 11500
rect 25410 11455 25466 11464
rect 25134 11384 25190 11393
rect 25134 11319 25190 11328
rect 25412 11280 25464 11286
rect 25412 11222 25464 11228
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24780 9064 24900 9092
rect 24780 8430 24808 9064
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24582 7919 24638 7928
rect 24676 7948 24728 7954
rect 24492 7890 24544 7896
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24412 7177 24440 7278
rect 24398 7168 24454 7177
rect 24398 7103 24454 7112
rect 24308 6724 24360 6730
rect 24308 6666 24360 6672
rect 24400 6724 24452 6730
rect 24400 6666 24452 6672
rect 24412 6322 24440 6666
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24504 5914 24532 7890
rect 24596 7478 24624 7919
rect 24676 7890 24728 7896
rect 24780 7546 24808 8230
rect 24964 8090 24992 9318
rect 25056 8838 25084 10066
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25056 8294 25084 8774
rect 25148 8430 25176 10950
rect 25226 10432 25282 10441
rect 25226 10367 25282 10376
rect 25240 9654 25268 10367
rect 25424 10305 25452 11222
rect 25516 11218 25544 11494
rect 25608 11354 25636 12038
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25700 10810 25728 13806
rect 25792 13326 25820 16730
rect 25884 16425 25912 16730
rect 25870 16416 25926 16425
rect 25870 16351 25926 16360
rect 25872 16176 25924 16182
rect 25872 16118 25924 16124
rect 25884 15366 25912 16118
rect 25976 16114 26004 17156
rect 26068 17134 26096 18686
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 26160 17678 26188 18566
rect 26344 18154 26372 18686
rect 26332 18148 26384 18154
rect 26332 18090 26384 18096
rect 26238 17912 26294 17921
rect 26238 17847 26294 17856
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 26252 17270 26280 17847
rect 26344 17814 26372 18090
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26436 17746 26464 18702
rect 26896 18272 26924 19740
rect 26984 19612 27292 19621
rect 26984 19610 26990 19612
rect 27046 19610 27070 19612
rect 27126 19610 27150 19612
rect 27206 19610 27230 19612
rect 27286 19610 27292 19612
rect 27046 19558 27048 19610
rect 27228 19558 27230 19610
rect 26984 19556 26990 19558
rect 27046 19556 27070 19558
rect 27126 19556 27150 19558
rect 27206 19556 27230 19558
rect 27286 19556 27292 19558
rect 26984 19547 27292 19556
rect 27356 19242 27384 20198
rect 27344 19236 27396 19242
rect 27344 19178 27396 19184
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 26984 18524 27292 18533
rect 26984 18522 26990 18524
rect 27046 18522 27070 18524
rect 27126 18522 27150 18524
rect 27206 18522 27230 18524
rect 27286 18522 27292 18524
rect 27046 18470 27048 18522
rect 27228 18470 27230 18522
rect 26984 18468 26990 18470
rect 27046 18468 27070 18470
rect 27126 18468 27150 18470
rect 27206 18468 27230 18470
rect 27286 18468 27292 18470
rect 26984 18459 27292 18468
rect 26804 18244 26924 18272
rect 26606 18184 26662 18193
rect 26516 18148 26568 18154
rect 26606 18119 26662 18128
rect 26516 18090 26568 18096
rect 26528 17882 26556 18090
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26424 17740 26476 17746
rect 26424 17682 26476 17688
rect 26620 17542 26648 18119
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26436 17377 26464 17478
rect 26422 17368 26478 17377
rect 26422 17303 26478 17312
rect 26240 17264 26292 17270
rect 26146 17232 26202 17241
rect 26240 17206 26292 17212
rect 26330 17232 26386 17241
rect 26146 17167 26202 17176
rect 26804 17218 26832 18244
rect 26884 18148 26936 18154
rect 26884 18090 26936 18096
rect 26896 17610 26924 18090
rect 26884 17604 26936 17610
rect 26884 17546 26936 17552
rect 26984 17436 27292 17445
rect 26984 17434 26990 17436
rect 27046 17434 27070 17436
rect 27126 17434 27150 17436
rect 27206 17434 27230 17436
rect 27286 17434 27292 17436
rect 27046 17382 27048 17434
rect 27228 17382 27230 17434
rect 26984 17380 26990 17382
rect 27046 17380 27070 17382
rect 27126 17380 27150 17382
rect 27206 17380 27230 17382
rect 27286 17380 27292 17382
rect 26984 17371 27292 17380
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 26804 17190 27108 17218
rect 26330 17167 26386 17176
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 26056 16992 26108 16998
rect 26056 16934 26108 16940
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25884 15201 25912 15302
rect 25870 15192 25926 15201
rect 25870 15127 25926 15136
rect 25872 14816 25924 14822
rect 25976 14804 26004 16050
rect 26068 16046 26096 16934
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 26068 15162 26096 15982
rect 26160 15638 26188 17167
rect 26344 16833 26372 17167
rect 26976 17128 27028 17134
rect 26896 17088 26976 17116
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26330 16824 26386 16833
rect 26330 16759 26386 16768
rect 26330 16688 26386 16697
rect 26330 16623 26386 16632
rect 26424 16652 26476 16658
rect 26344 16590 26372 16623
rect 26424 16594 26476 16600
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26332 16584 26384 16590
rect 26238 16552 26294 16561
rect 26436 16561 26464 16594
rect 26332 16526 26384 16532
rect 26422 16552 26478 16561
rect 26238 16487 26294 16496
rect 26422 16487 26478 16496
rect 26252 16250 26280 16487
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26344 16046 26372 16390
rect 26422 16280 26478 16289
rect 26528 16250 26556 16594
rect 26422 16215 26478 16224
rect 26516 16244 26568 16250
rect 26436 16114 26464 16215
rect 26516 16186 26568 16192
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26148 15632 26200 15638
rect 26148 15574 26200 15580
rect 26344 15570 26372 15982
rect 26528 15706 26556 16186
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 25924 14776 26004 14804
rect 26148 14816 26200 14822
rect 25872 14758 25924 14764
rect 26148 14758 26200 14764
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 25884 13394 25912 14758
rect 25962 14648 26018 14657
rect 25962 14583 25964 14592
rect 26016 14583 26018 14592
rect 25964 14554 26016 14560
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25976 14249 26004 14418
rect 26056 14408 26108 14414
rect 26056 14350 26108 14356
rect 25962 14240 26018 14249
rect 25962 14175 26018 14184
rect 25964 14000 26016 14006
rect 25962 13968 25964 13977
rect 26016 13968 26018 13977
rect 25962 13903 26018 13912
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 25872 13388 25924 13394
rect 25872 13330 25924 13336
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25884 13161 25912 13330
rect 25870 13152 25926 13161
rect 25870 13087 25926 13096
rect 25976 12442 26004 13806
rect 25964 12436 26016 12442
rect 25964 12378 26016 12384
rect 25778 12336 25834 12345
rect 25778 12271 25780 12280
rect 25832 12271 25834 12280
rect 25780 12242 25832 12248
rect 25792 11665 25820 12242
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 25884 11694 25912 11834
rect 25872 11688 25924 11694
rect 25778 11656 25834 11665
rect 25872 11630 25924 11636
rect 25962 11656 26018 11665
rect 25778 11591 25834 11600
rect 25778 11520 25834 11529
rect 25778 11455 25834 11464
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25410 10296 25466 10305
rect 25410 10231 25466 10240
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25240 9382 25268 9454
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25134 8120 25190 8129
rect 24952 8084 25004 8090
rect 25134 8055 25190 8064
rect 24952 8026 25004 8032
rect 25044 8016 25096 8022
rect 25044 7958 25096 7964
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24674 7440 24730 7449
rect 24872 7426 24900 7890
rect 25056 7721 25084 7958
rect 25148 7954 25176 8055
rect 25136 7948 25188 7954
rect 25136 7890 25188 7896
rect 25042 7712 25098 7721
rect 25042 7647 25098 7656
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24674 7375 24730 7384
rect 24780 7398 24900 7426
rect 24584 7336 24636 7342
rect 24688 7324 24716 7375
rect 24636 7296 24716 7324
rect 24584 7278 24636 7284
rect 24780 7206 24808 7398
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24768 7200 24820 7206
rect 24872 7177 24900 7210
rect 24964 7206 24992 7482
rect 25044 7472 25096 7478
rect 25240 7426 25268 8910
rect 25332 8888 25360 9862
rect 25516 9722 25544 10406
rect 25608 10198 25636 10406
rect 25596 10192 25648 10198
rect 25596 10134 25648 10140
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25424 9042 25452 9658
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 25332 8860 25452 8888
rect 25320 7948 25372 7954
rect 25320 7890 25372 7896
rect 25332 7449 25360 7890
rect 25424 7562 25452 8860
rect 25516 8294 25544 9318
rect 25608 8634 25636 9930
rect 25792 9926 25820 11455
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 25686 9616 25742 9625
rect 25686 9551 25742 9560
rect 25700 9450 25728 9551
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25792 9217 25820 9386
rect 25778 9208 25834 9217
rect 25778 9143 25834 9152
rect 25686 9072 25742 9081
rect 25686 9007 25742 9016
rect 25700 8838 25728 9007
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25516 7818 25544 8230
rect 25504 7812 25556 7818
rect 25504 7754 25556 7760
rect 25502 7576 25558 7585
rect 25424 7534 25502 7562
rect 25502 7511 25558 7520
rect 25044 7414 25096 7420
rect 25056 7342 25084 7414
rect 25148 7398 25268 7426
rect 25318 7440 25374 7449
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 24952 7200 25004 7206
rect 24768 7142 24820 7148
rect 24858 7168 24914 7177
rect 24952 7142 25004 7148
rect 24858 7103 24914 7112
rect 24582 7032 24638 7041
rect 24582 6967 24584 6976
rect 24636 6967 24638 6976
rect 24584 6938 24636 6944
rect 24768 6928 24820 6934
rect 24768 6870 24820 6876
rect 24858 6896 24914 6905
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24596 6458 24624 6598
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 24688 6186 24716 6802
rect 24780 6390 24808 6870
rect 24858 6831 24914 6840
rect 24872 6662 24900 6831
rect 24964 6798 24992 7142
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24768 6384 24820 6390
rect 24768 6326 24820 6332
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24412 5166 24440 5238
rect 24504 5166 24532 5850
rect 24780 5778 24808 6326
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24780 5302 24808 5714
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 24228 4146 24256 5102
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23846 3496 23902 3505
rect 23846 3431 23902 3440
rect 12096 2748 12404 2757
rect 12096 2746 12102 2748
rect 12158 2746 12182 2748
rect 12238 2746 12262 2748
rect 12318 2746 12342 2748
rect 12398 2746 12404 2748
rect 12158 2694 12160 2746
rect 12340 2694 12342 2746
rect 12096 2692 12102 2694
rect 12158 2692 12182 2694
rect 12238 2692 12262 2694
rect 12318 2692 12342 2694
rect 12398 2692 12404 2694
rect 12096 2683 12404 2692
rect 19870 2748 20178 2757
rect 19870 2746 19876 2748
rect 19932 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20178 2748
rect 23308 2746 23428 2774
rect 19932 2694 19934 2746
rect 20114 2694 20116 2746
rect 19870 2692 19876 2694
rect 19932 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20178 2694
rect 19706 2680 19762 2689
rect 19870 2683 20178 2692
rect 19706 2615 19762 2624
rect 11888 2440 11940 2446
rect 10874 2408 10930 2417
rect 11888 2382 11940 2388
rect 10874 2343 10930 2352
rect 19720 2281 19748 2615
rect 23400 2514 23428 2746
rect 24596 2650 24624 4966
rect 24688 4282 24716 5170
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24872 3534 24900 6394
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 25056 4826 25084 4966
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25148 4690 25176 7398
rect 25318 7375 25374 7384
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25228 7268 25280 7274
rect 25228 7210 25280 7216
rect 25240 6662 25268 7210
rect 25424 7002 25452 7346
rect 25516 7342 25544 7511
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25412 6996 25464 7002
rect 25412 6938 25464 6944
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25332 6610 25360 6802
rect 25608 6798 25636 8434
rect 25700 7970 25728 8774
rect 25792 8634 25820 9143
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25792 8090 25820 8366
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25700 7942 25820 7970
rect 25792 7818 25820 7942
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25780 7812 25832 7818
rect 25780 7754 25832 7760
rect 25596 6792 25648 6798
rect 25516 6752 25596 6780
rect 25240 6236 25268 6598
rect 25332 6582 25452 6610
rect 25320 6248 25372 6254
rect 25240 6208 25320 6236
rect 25320 6190 25372 6196
rect 25332 5914 25360 6190
rect 25424 6186 25452 6582
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25332 5710 25360 5850
rect 25424 5710 25452 6122
rect 25516 5760 25544 6752
rect 25700 6769 25728 7754
rect 25778 7168 25834 7177
rect 25778 7103 25834 7112
rect 25792 7002 25820 7103
rect 25780 6996 25832 7002
rect 25780 6938 25832 6944
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25596 6734 25648 6740
rect 25686 6760 25742 6769
rect 25686 6695 25742 6704
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25608 6497 25636 6598
rect 25594 6488 25650 6497
rect 25594 6423 25650 6432
rect 25792 6390 25820 6802
rect 25884 6458 25912 11630
rect 25962 11591 26018 11600
rect 25976 11121 26004 11591
rect 25962 11112 26018 11121
rect 26068 11082 26096 14350
rect 26160 13462 26188 14758
rect 26252 14482 26280 14758
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26238 13696 26294 13705
rect 26238 13631 26294 13640
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 26252 13258 26280 13631
rect 26344 13462 26372 14962
rect 26436 14618 26464 15574
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26620 14006 26648 16934
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26804 16658 26832 16730
rect 26896 16697 26924 17088
rect 26976 17070 27028 17076
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 26882 16688 26938 16697
rect 26792 16652 26844 16658
rect 26712 16612 26792 16640
rect 26712 16114 26740 16612
rect 26882 16623 26938 16632
rect 26792 16594 26844 16600
rect 26792 16448 26844 16454
rect 26792 16390 26844 16396
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26712 15745 26740 16050
rect 26698 15736 26754 15745
rect 26698 15671 26754 15680
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26712 14657 26740 15302
rect 26698 14648 26754 14657
rect 26698 14583 26754 14592
rect 26698 14104 26754 14113
rect 26698 14039 26700 14048
rect 26752 14039 26754 14048
rect 26700 14010 26752 14016
rect 26608 14000 26660 14006
rect 26608 13942 26660 13948
rect 26698 13968 26754 13977
rect 26698 13903 26754 13912
rect 26332 13456 26384 13462
rect 26332 13398 26384 13404
rect 26516 13456 26568 13462
rect 26516 13398 26568 13404
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26148 13184 26200 13190
rect 26148 13126 26200 13132
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26422 13152 26478 13161
rect 26160 12850 26188 13126
rect 26344 13025 26372 13126
rect 26422 13087 26478 13096
rect 26330 13016 26386 13025
rect 26330 12951 26386 12960
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26148 12708 26200 12714
rect 26148 12650 26200 12656
rect 26160 12345 26188 12650
rect 26436 12424 26464 13087
rect 26528 12850 26556 13398
rect 26608 13388 26660 13394
rect 26712 13376 26740 13903
rect 26804 13705 26832 16390
rect 26896 16182 26924 16623
rect 26988 16522 27016 16730
rect 26976 16516 27028 16522
rect 26976 16458 27028 16464
rect 27080 16454 27108 17190
rect 27172 16590 27200 17274
rect 27356 17202 27384 18702
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27344 17060 27396 17066
rect 27344 17002 27396 17008
rect 27356 16969 27384 17002
rect 27342 16960 27398 16969
rect 27342 16895 27398 16904
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 26984 16348 27292 16357
rect 26984 16346 26990 16348
rect 27046 16346 27070 16348
rect 27126 16346 27150 16348
rect 27206 16346 27230 16348
rect 27286 16346 27292 16348
rect 27046 16294 27048 16346
rect 27228 16294 27230 16346
rect 26984 16292 26990 16294
rect 27046 16292 27070 16294
rect 27126 16292 27150 16294
rect 27206 16292 27230 16294
rect 27286 16292 27292 16294
rect 26984 16283 27292 16292
rect 26884 16176 26936 16182
rect 26884 16118 26936 16124
rect 27068 16176 27120 16182
rect 27068 16118 27120 16124
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 26896 15910 26924 15982
rect 26884 15904 26936 15910
rect 26884 15846 26936 15852
rect 26896 15065 26924 15846
rect 27080 15473 27108 16118
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27172 15910 27200 16050
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27160 15564 27212 15570
rect 27160 15506 27212 15512
rect 27066 15464 27122 15473
rect 27066 15399 27122 15408
rect 27172 15366 27200 15506
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 26984 15260 27292 15269
rect 26984 15258 26990 15260
rect 27046 15258 27070 15260
rect 27126 15258 27150 15260
rect 27206 15258 27230 15260
rect 27286 15258 27292 15260
rect 27046 15206 27048 15258
rect 27228 15206 27230 15258
rect 26984 15204 26990 15206
rect 27046 15204 27070 15206
rect 27126 15204 27150 15206
rect 27206 15204 27230 15206
rect 27286 15204 27292 15206
rect 26984 15195 27292 15204
rect 26882 15056 26938 15065
rect 26882 14991 26938 15000
rect 27356 14958 27384 16895
rect 27448 15094 27476 20352
rect 27620 20334 27672 20340
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27540 19258 27568 20198
rect 27644 20156 27952 20165
rect 27644 20154 27650 20156
rect 27706 20154 27730 20156
rect 27786 20154 27810 20156
rect 27866 20154 27890 20156
rect 27946 20154 27952 20156
rect 27706 20102 27708 20154
rect 27888 20102 27890 20154
rect 27644 20100 27650 20102
rect 27706 20100 27730 20102
rect 27786 20100 27810 20102
rect 27866 20100 27890 20102
rect 27946 20100 27952 20102
rect 27644 20091 27952 20100
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27816 19378 27844 19654
rect 28000 19378 28028 19858
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 28092 19334 28120 20839
rect 28184 20210 28212 21286
rect 28276 20398 28304 21354
rect 28264 20392 28316 20398
rect 28264 20334 28316 20340
rect 28184 20182 28304 20210
rect 28170 20088 28226 20097
rect 28170 20023 28226 20032
rect 28184 19854 28212 20023
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 28276 19718 28304 20182
rect 28368 19854 28396 21558
rect 28814 21448 28870 21457
rect 28814 21383 28870 21392
rect 29368 21412 29420 21418
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28632 21344 28684 21350
rect 28828 21332 28856 21383
rect 29368 21354 29420 21360
rect 29000 21344 29052 21350
rect 28828 21304 28948 21332
rect 28632 21286 28684 21292
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28460 20602 28488 20878
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28460 19786 28488 20334
rect 28552 20058 28580 21286
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28552 19922 28580 19994
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 28448 19780 28500 19786
rect 28448 19722 28500 19728
rect 28540 19780 28592 19786
rect 28540 19722 28592 19728
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28276 19446 28304 19654
rect 28264 19440 28316 19446
rect 28264 19382 28316 19388
rect 27540 19230 27660 19258
rect 27632 19174 27660 19230
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27540 18630 27568 19110
rect 27644 19068 27952 19077
rect 27644 19066 27650 19068
rect 27706 19066 27730 19068
rect 27786 19066 27810 19068
rect 27866 19066 27890 19068
rect 27946 19066 27952 19068
rect 27706 19014 27708 19066
rect 27888 19014 27890 19066
rect 27644 19012 27650 19014
rect 27706 19012 27730 19014
rect 27786 19012 27810 19014
rect 27866 19012 27890 19014
rect 27946 19012 27952 19014
rect 27644 19003 27952 19012
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27540 18290 27568 18566
rect 27724 18465 27752 18906
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 27710 18456 27766 18465
rect 27710 18391 27766 18400
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27540 17796 27568 18226
rect 27908 18222 27936 18770
rect 27712 18216 27764 18222
rect 27710 18184 27712 18193
rect 27896 18216 27948 18222
rect 27764 18184 27766 18193
rect 27710 18119 27766 18128
rect 27894 18184 27896 18193
rect 27948 18184 27950 18193
rect 27894 18119 27950 18128
rect 27644 17980 27952 17989
rect 27644 17978 27650 17980
rect 27706 17978 27730 17980
rect 27786 17978 27810 17980
rect 27866 17978 27890 17980
rect 27946 17978 27952 17980
rect 27706 17926 27708 17978
rect 27888 17926 27890 17978
rect 27644 17924 27650 17926
rect 27706 17924 27730 17926
rect 27786 17924 27810 17926
rect 27866 17924 27890 17926
rect 27946 17924 27952 17926
rect 27644 17915 27952 17924
rect 28000 17882 28028 19314
rect 28092 19306 28212 19334
rect 28080 18828 28132 18834
rect 28080 18770 28132 18776
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 27620 17808 27672 17814
rect 27540 17768 27620 17796
rect 27620 17750 27672 17756
rect 28092 17524 28120 18770
rect 28184 18714 28212 19306
rect 28460 18714 28488 19722
rect 28552 19689 28580 19722
rect 28644 19718 28672 21286
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28724 21072 28776 21078
rect 28724 21014 28776 21020
rect 28736 20602 28764 21014
rect 28828 21010 28856 21082
rect 28920 21078 28948 21304
rect 29000 21286 29052 21292
rect 28908 21072 28960 21078
rect 28908 21014 28960 21020
rect 28816 21004 28868 21010
rect 28816 20946 28868 20952
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28816 20596 28868 20602
rect 28816 20538 28868 20544
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28632 19712 28684 19718
rect 28538 19680 28594 19689
rect 28632 19654 28684 19660
rect 28538 19615 28594 19624
rect 28736 19514 28764 20334
rect 28828 20058 28856 20538
rect 29012 20466 29040 21286
rect 29274 21176 29330 21185
rect 29380 21146 29408 21354
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 29274 21111 29276 21120
rect 29328 21111 29330 21120
rect 29368 21140 29420 21146
rect 29276 21082 29328 21088
rect 29368 21082 29420 21088
rect 29472 21100 29776 21128
rect 29472 20874 29500 21100
rect 29748 21010 29776 21100
rect 29828 21072 29880 21078
rect 29828 21014 29880 21020
rect 29552 21004 29604 21010
rect 29552 20946 29604 20952
rect 29644 21004 29696 21010
rect 29644 20946 29696 20952
rect 29736 21004 29788 21010
rect 29736 20946 29788 20952
rect 29460 20868 29512 20874
rect 29460 20810 29512 20816
rect 29092 20800 29144 20806
rect 29144 20760 29224 20788
rect 29092 20742 29144 20748
rect 28908 20460 28960 20466
rect 28908 20402 28960 20408
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28920 20346 28948 20402
rect 28920 20318 29132 20346
rect 29000 20256 29052 20262
rect 28906 20224 28962 20233
rect 29000 20198 29052 20204
rect 28906 20159 28962 20168
rect 28920 20058 28948 20159
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28908 20052 28960 20058
rect 28908 19994 28960 20000
rect 29012 19825 29040 20198
rect 28998 19816 29054 19825
rect 28998 19751 29054 19760
rect 28816 19712 28868 19718
rect 28816 19654 28868 19660
rect 28828 19514 28856 19654
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28736 19145 28764 19450
rect 28908 19440 28960 19446
rect 28908 19382 28960 19388
rect 28816 19168 28868 19174
rect 28722 19136 28778 19145
rect 28816 19110 28868 19116
rect 28722 19071 28778 19080
rect 28828 18714 28856 19110
rect 28184 18686 28396 18714
rect 28460 18686 28856 18714
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 27894 17504 27950 17513
rect 27894 17439 27950 17448
rect 28000 17496 28120 17524
rect 28184 17513 28212 18566
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 28276 18222 28304 18294
rect 28264 18216 28316 18222
rect 28264 18158 28316 18164
rect 28368 18057 28396 18686
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28460 18222 28488 18362
rect 28448 18216 28500 18222
rect 28448 18158 28500 18164
rect 28354 18048 28410 18057
rect 28354 17983 28410 17992
rect 28368 17814 28396 17983
rect 28356 17808 28408 17814
rect 28356 17750 28408 17756
rect 28356 17604 28408 17610
rect 28356 17546 28408 17552
rect 28264 17536 28316 17542
rect 28170 17504 28226 17513
rect 27526 17368 27582 17377
rect 27526 17303 27528 17312
rect 27580 17303 27582 17312
rect 27528 17274 27580 17280
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27540 16182 27568 17138
rect 27908 17134 27936 17439
rect 28000 17202 28028 17496
rect 28264 17478 28316 17484
rect 28170 17439 28226 17448
rect 28078 17232 28134 17241
rect 27988 17196 28040 17202
rect 28078 17167 28134 17176
rect 27988 17138 28040 17144
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 28092 17082 28120 17167
rect 28092 17054 28212 17082
rect 27804 16992 27856 16998
rect 27856 16952 28028 16980
rect 27804 16934 27856 16940
rect 28000 16946 28028 16952
rect 28078 16960 28134 16969
rect 28000 16918 28078 16946
rect 27644 16892 27952 16901
rect 27644 16890 27650 16892
rect 27706 16890 27730 16892
rect 27786 16890 27810 16892
rect 27866 16890 27890 16892
rect 27946 16890 27952 16892
rect 27706 16838 27708 16890
rect 27888 16838 27890 16890
rect 27644 16836 27650 16838
rect 27706 16836 27730 16838
rect 27786 16836 27810 16838
rect 27866 16836 27890 16838
rect 27946 16836 27952 16838
rect 27644 16827 27952 16836
rect 27804 16788 27856 16794
rect 28000 16776 28028 16918
rect 28078 16895 28134 16904
rect 27856 16748 28028 16776
rect 27804 16730 27856 16736
rect 28080 16720 28132 16726
rect 28078 16688 28080 16697
rect 28132 16688 28134 16697
rect 28184 16658 28212 17054
rect 28078 16623 28134 16632
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27988 16584 28040 16590
rect 27988 16526 28040 16532
rect 27528 16176 27580 16182
rect 27620 16176 27672 16182
rect 27528 16118 27580 16124
rect 27618 16144 27620 16153
rect 27672 16144 27674 16153
rect 27540 15688 27568 16118
rect 27618 16079 27674 16088
rect 27816 16046 27844 16526
rect 27896 16448 27948 16454
rect 27896 16390 27948 16396
rect 28000 16402 28028 16526
rect 28080 16516 28132 16522
rect 28132 16476 28212 16504
rect 28080 16458 28132 16464
rect 27804 16040 27856 16046
rect 27908 16028 27936 16390
rect 28000 16374 28120 16402
rect 27988 16176 28040 16182
rect 27986 16144 27988 16153
rect 28040 16144 28042 16153
rect 27986 16079 28042 16088
rect 27908 16000 28028 16028
rect 27804 15982 27856 15988
rect 27644 15804 27952 15813
rect 27644 15802 27650 15804
rect 27706 15802 27730 15804
rect 27786 15802 27810 15804
rect 27866 15802 27890 15804
rect 27946 15802 27952 15804
rect 27706 15750 27708 15802
rect 27888 15750 27890 15802
rect 27644 15748 27650 15750
rect 27706 15748 27730 15750
rect 27786 15748 27810 15750
rect 27866 15748 27890 15750
rect 27946 15748 27952 15750
rect 27644 15739 27952 15748
rect 27620 15700 27672 15706
rect 27540 15660 27620 15688
rect 27896 15700 27948 15706
rect 27672 15660 27752 15688
rect 27620 15642 27672 15648
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27632 15162 27660 15506
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27724 14822 27752 15660
rect 27896 15642 27948 15648
rect 27908 14929 27936 15642
rect 27894 14920 27950 14929
rect 27894 14855 27950 14864
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27356 14482 27384 14758
rect 27644 14716 27952 14725
rect 27644 14714 27650 14716
rect 27706 14714 27730 14716
rect 27786 14714 27810 14716
rect 27866 14714 27890 14716
rect 27946 14714 27952 14716
rect 27706 14662 27708 14714
rect 27888 14662 27890 14714
rect 27644 14660 27650 14662
rect 27706 14660 27730 14662
rect 27786 14660 27810 14662
rect 27866 14660 27890 14662
rect 27946 14660 27952 14662
rect 27644 14651 27952 14660
rect 28000 14600 28028 16000
rect 28092 15706 28120 16374
rect 28184 15994 28212 16476
rect 28276 16114 28304 17478
rect 28368 17184 28396 17546
rect 28460 17377 28488 18158
rect 28552 18086 28580 18686
rect 28920 18358 28948 19382
rect 29000 19304 29052 19310
rect 29000 19246 29052 19252
rect 28908 18352 28960 18358
rect 28908 18294 28960 18300
rect 29012 18290 29040 19246
rect 29104 18902 29132 20318
rect 29196 18970 29224 20760
rect 29276 20324 29328 20330
rect 29276 20266 29328 20272
rect 29288 20058 29316 20266
rect 29472 20097 29500 20810
rect 29458 20088 29514 20097
rect 29276 20052 29328 20058
rect 29458 20023 29514 20032
rect 29276 19994 29328 20000
rect 29472 19990 29500 20023
rect 29460 19984 29512 19990
rect 29564 19961 29592 20946
rect 29460 19926 29512 19932
rect 29550 19952 29606 19961
rect 29368 19916 29420 19922
rect 29656 19938 29684 20946
rect 29840 20505 29868 21014
rect 30208 20942 30236 21286
rect 30196 20936 30248 20942
rect 30196 20878 30248 20884
rect 29826 20496 29882 20505
rect 29826 20431 29882 20440
rect 29840 20233 29868 20431
rect 29826 20224 29882 20233
rect 29826 20159 29882 20168
rect 29840 20058 29868 20159
rect 29828 20052 29880 20058
rect 29828 19994 29880 20000
rect 29656 19910 29868 19938
rect 29550 19887 29606 19896
rect 29368 19858 29420 19864
rect 29276 19712 29328 19718
rect 29276 19654 29328 19660
rect 29288 19242 29316 19654
rect 29276 19236 29328 19242
rect 29276 19178 29328 19184
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 29092 18896 29144 18902
rect 29092 18838 29144 18844
rect 29276 18828 29328 18834
rect 29276 18770 29328 18776
rect 29288 18426 29316 18770
rect 29092 18420 29144 18426
rect 29092 18362 29144 18368
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 28632 18216 28684 18222
rect 28630 18184 28632 18193
rect 28684 18184 28686 18193
rect 28630 18119 28686 18128
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 28446 17368 28502 17377
rect 28446 17303 28502 17312
rect 28448 17196 28500 17202
rect 28368 17156 28448 17184
rect 28368 16658 28396 17156
rect 28448 17138 28500 17144
rect 28448 17060 28500 17066
rect 28448 17002 28500 17008
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28354 16552 28410 16561
rect 28354 16487 28410 16496
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28184 15966 28304 15994
rect 28276 15892 28304 15966
rect 28184 15864 28304 15892
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 28184 15502 28212 15864
rect 28368 15570 28396 16487
rect 28460 16454 28488 17002
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28446 16144 28502 16153
rect 28446 16079 28502 16088
rect 28460 15706 28488 16079
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28446 15600 28502 15609
rect 28356 15564 28408 15570
rect 28446 15535 28448 15544
rect 28356 15506 28408 15512
rect 28500 15535 28502 15544
rect 28448 15506 28500 15512
rect 28172 15496 28224 15502
rect 27908 14572 28028 14600
rect 28092 15456 28172 15484
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 27344 14476 27396 14482
rect 27344 14418 27396 14424
rect 26988 14385 27016 14418
rect 26974 14376 27030 14385
rect 26974 14311 27030 14320
rect 26984 14172 27292 14181
rect 26984 14170 26990 14172
rect 27046 14170 27070 14172
rect 27126 14170 27150 14172
rect 27206 14170 27230 14172
rect 27286 14170 27292 14172
rect 27046 14118 27048 14170
rect 27228 14118 27230 14170
rect 26984 14116 26990 14118
rect 27046 14116 27070 14118
rect 27126 14116 27150 14118
rect 27206 14116 27230 14118
rect 27286 14116 27292 14118
rect 26984 14107 27292 14116
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26790 13696 26846 13705
rect 26790 13631 26846 13640
rect 26660 13348 26740 13376
rect 26608 13330 26660 13336
rect 26516 12844 26568 12850
rect 26568 12804 26648 12832
rect 26516 12786 26568 12792
rect 26516 12436 26568 12442
rect 26436 12396 26516 12424
rect 26516 12378 26568 12384
rect 26146 12336 26202 12345
rect 26146 12271 26202 12280
rect 26240 12300 26292 12306
rect 26160 11694 26188 12271
rect 26240 12242 26292 12248
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 26252 11898 26280 12242
rect 26436 12209 26464 12242
rect 26422 12200 26478 12209
rect 26422 12135 26478 12144
rect 26516 12164 26568 12170
rect 26516 12106 26568 12112
rect 26424 12096 26476 12102
rect 26424 12038 26476 12044
rect 26330 11928 26386 11937
rect 26240 11892 26292 11898
rect 26436 11898 26464 12038
rect 26330 11863 26386 11872
rect 26424 11892 26476 11898
rect 26240 11834 26292 11840
rect 26344 11830 26372 11863
rect 26424 11834 26476 11840
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26330 11520 26386 11529
rect 26330 11455 26386 11464
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 25962 11047 26018 11056
rect 26056 11076 26108 11082
rect 26056 11018 26108 11024
rect 25962 10976 26018 10985
rect 25962 10911 26018 10920
rect 25976 10606 26004 10911
rect 26056 10736 26108 10742
rect 26056 10678 26108 10684
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 25976 10198 26004 10542
rect 25964 10192 26016 10198
rect 25964 10134 26016 10140
rect 26068 10130 26096 10678
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 26056 10124 26108 10130
rect 26056 10066 26108 10072
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 25976 9178 26004 9998
rect 26160 9897 26188 10474
rect 26146 9888 26202 9897
rect 26146 9823 26202 9832
rect 26148 9580 26200 9586
rect 26252 9568 26280 11154
rect 26344 10606 26372 11455
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26436 10606 26464 10746
rect 26332 10600 26384 10606
rect 26332 10542 26384 10548
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26330 10296 26386 10305
rect 26436 10266 26464 10542
rect 26330 10231 26386 10240
rect 26424 10260 26476 10266
rect 26344 10044 26372 10231
rect 26424 10202 26476 10208
rect 26344 10016 26464 10044
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26200 9540 26280 9568
rect 26148 9522 26200 9528
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26068 9178 26096 9454
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25976 8430 26004 8774
rect 26054 8528 26110 8537
rect 26160 8514 26188 9318
rect 26110 8486 26188 8514
rect 26252 8498 26280 9540
rect 26344 9382 26372 9862
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26436 8838 26464 10016
rect 26528 9994 26556 12106
rect 26620 11762 26648 12804
rect 26712 12714 26740 13348
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26700 12708 26752 12714
rect 26700 12650 26752 12656
rect 26698 12608 26754 12617
rect 26804 12594 26832 13262
rect 26754 12566 26832 12594
rect 26698 12543 26754 12552
rect 26712 12374 26740 12543
rect 26700 12368 26752 12374
rect 26700 12310 26752 12316
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 26804 12209 26832 12242
rect 26790 12200 26846 12209
rect 26790 12135 26846 12144
rect 26896 12102 26924 13942
rect 26974 13560 27030 13569
rect 26974 13495 27030 13504
rect 26988 13394 27016 13495
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26984 13084 27292 13093
rect 26984 13082 26990 13084
rect 27046 13082 27070 13084
rect 27126 13082 27150 13084
rect 27206 13082 27230 13084
rect 27286 13082 27292 13084
rect 27046 13030 27048 13082
rect 27228 13030 27230 13082
rect 26984 13028 26990 13030
rect 27046 13028 27070 13030
rect 27126 13028 27150 13030
rect 27206 13028 27230 13030
rect 27286 13028 27292 13030
rect 26984 13019 27292 13028
rect 27356 12968 27384 14418
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27264 12940 27384 12968
rect 27160 12912 27212 12918
rect 26974 12880 27030 12889
rect 26974 12815 26976 12824
rect 27028 12815 27030 12824
rect 27080 12872 27160 12900
rect 26976 12786 27028 12792
rect 27080 12306 27108 12872
rect 27160 12854 27212 12860
rect 27160 12436 27212 12442
rect 27160 12378 27212 12384
rect 27172 12345 27200 12378
rect 27158 12336 27214 12345
rect 27068 12300 27120 12306
rect 27264 12306 27292 12940
rect 27448 12832 27476 13126
rect 27356 12804 27476 12832
rect 27158 12271 27214 12280
rect 27252 12300 27304 12306
rect 27068 12242 27120 12248
rect 27252 12242 27304 12248
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26712 10742 26740 12038
rect 26984 11996 27292 12005
rect 26984 11994 26990 11996
rect 27046 11994 27070 11996
rect 27126 11994 27150 11996
rect 27206 11994 27230 11996
rect 27286 11994 27292 11996
rect 27046 11942 27048 11994
rect 27228 11942 27230 11994
rect 26984 11940 26990 11942
rect 27046 11940 27070 11942
rect 27126 11940 27150 11942
rect 27206 11940 27230 11942
rect 27286 11940 27292 11942
rect 26984 11931 27292 11940
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27068 11688 27120 11694
rect 27068 11630 27120 11636
rect 26882 11384 26938 11393
rect 26882 11319 26938 11328
rect 26896 11014 26924 11319
rect 27080 11257 27108 11630
rect 27066 11248 27122 11257
rect 27264 11218 27292 11698
rect 27066 11183 27122 11192
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 26884 11008 26936 11014
rect 26884 10950 26936 10956
rect 26896 10792 26924 10950
rect 26984 10908 27292 10917
rect 26984 10906 26990 10908
rect 27046 10906 27070 10908
rect 27126 10906 27150 10908
rect 27206 10906 27230 10908
rect 27286 10906 27292 10908
rect 27046 10854 27048 10906
rect 27228 10854 27230 10906
rect 26984 10852 26990 10854
rect 27046 10852 27070 10854
rect 27126 10852 27150 10854
rect 27206 10852 27230 10854
rect 27286 10852 27292 10854
rect 26984 10843 27292 10852
rect 26896 10764 27292 10792
rect 26700 10736 26752 10742
rect 26700 10678 26752 10684
rect 26792 10736 26844 10742
rect 26792 10678 26844 10684
rect 26608 10056 26660 10062
rect 26606 10024 26608 10033
rect 26660 10024 26662 10033
rect 26516 9988 26568 9994
rect 26606 9959 26662 9968
rect 26516 9930 26568 9936
rect 26698 9752 26754 9761
rect 26804 9722 26832 10678
rect 26884 10600 26936 10606
rect 26884 10542 26936 10548
rect 26698 9687 26754 9696
rect 26792 9716 26844 9722
rect 26516 9648 26568 9654
rect 26516 9590 26568 9596
rect 26528 9217 26556 9590
rect 26712 9586 26740 9687
rect 26792 9658 26844 9664
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26514 9208 26570 9217
rect 26514 9143 26570 9152
rect 26514 9072 26570 9081
rect 26514 9007 26570 9016
rect 26528 8838 26556 9007
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26422 8664 26478 8673
rect 26332 8628 26384 8634
rect 26422 8599 26478 8608
rect 26332 8570 26384 8576
rect 26240 8492 26292 8498
rect 26054 8463 26110 8472
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 25976 8265 26004 8366
rect 25962 8256 26018 8265
rect 25962 8191 26018 8200
rect 25964 8016 26016 8022
rect 26068 8004 26096 8463
rect 26240 8434 26292 8440
rect 26148 8424 26200 8430
rect 26148 8366 26200 8372
rect 26016 7976 26096 8004
rect 25964 7958 26016 7964
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25872 6452 25924 6458
rect 25872 6394 25924 6400
rect 25780 6384 25832 6390
rect 25780 6326 25832 6332
rect 25792 6254 25820 6326
rect 25780 6248 25832 6254
rect 25780 6190 25832 6196
rect 25596 5772 25648 5778
rect 25516 5732 25596 5760
rect 25596 5714 25648 5720
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 25332 4690 25360 5306
rect 25424 5273 25452 5646
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 25410 5264 25466 5273
rect 25410 5199 25466 5208
rect 25424 5166 25452 5199
rect 25412 5160 25464 5166
rect 25412 5102 25464 5108
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25056 4010 25084 4626
rect 25148 4214 25176 4626
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25516 4078 25544 5578
rect 25792 5370 25820 6190
rect 25976 5778 26004 7822
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 26068 7410 26096 7686
rect 26160 7546 26188 8366
rect 26252 8265 26280 8434
rect 26238 8256 26294 8265
rect 26238 8191 26294 8200
rect 26344 7954 26372 8570
rect 26436 8566 26464 8599
rect 26424 8560 26476 8566
rect 26424 8502 26476 8508
rect 26528 8412 26556 8774
rect 26436 8384 26556 8412
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 26238 7848 26294 7857
rect 26238 7783 26294 7792
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26252 7342 26280 7783
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 25872 5772 25924 5778
rect 25872 5714 25924 5720
rect 25964 5772 26016 5778
rect 25964 5714 26016 5720
rect 25884 5370 25912 5714
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25792 4758 25820 5306
rect 25780 4752 25832 4758
rect 25780 4694 25832 4700
rect 25884 4078 25912 5306
rect 25976 5234 26004 5714
rect 26068 5574 26096 7142
rect 26344 6866 26372 7890
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 26160 6390 26188 6734
rect 26148 6384 26200 6390
rect 26148 6326 26200 6332
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26344 5302 26372 5714
rect 26332 5296 26384 5302
rect 26332 5238 26384 5244
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25976 4146 26004 5170
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25044 4004 25096 4010
rect 25044 3946 25096 3952
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24858 2680 24914 2689
rect 24584 2644 24636 2650
rect 24858 2615 24914 2624
rect 24584 2586 24636 2592
rect 24872 2582 24900 2615
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 19706 2272 19762 2281
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 11436 2204 11744 2213
rect 11436 2202 11442 2204
rect 11498 2202 11522 2204
rect 11578 2202 11602 2204
rect 11658 2202 11682 2204
rect 11738 2202 11744 2204
rect 11498 2150 11500 2202
rect 11680 2150 11682 2202
rect 11436 2148 11442 2150
rect 11498 2148 11522 2150
rect 11578 2148 11602 2150
rect 11658 2148 11682 2150
rect 11738 2148 11744 2150
rect 11436 2139 11744 2148
rect 19210 2204 19518 2213
rect 19706 2207 19762 2216
rect 19210 2202 19216 2204
rect 19272 2202 19296 2204
rect 19352 2202 19376 2204
rect 19432 2202 19456 2204
rect 19512 2202 19518 2204
rect 19272 2150 19274 2202
rect 19454 2150 19456 2202
rect 19210 2148 19216 2150
rect 19272 2148 19296 2150
rect 19352 2148 19376 2150
rect 19432 2148 19456 2150
rect 19512 2148 19518 2150
rect 19210 2139 19518 2148
rect 26436 2009 26464 8384
rect 26516 7744 26568 7750
rect 26514 7712 26516 7721
rect 26568 7712 26570 7721
rect 26514 7647 26570 7656
rect 26528 7410 26556 7647
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26620 6322 26648 9454
rect 26804 8974 26832 9658
rect 26896 9042 26924 10542
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 26976 10464 27028 10470
rect 27080 10441 27108 10474
rect 27160 10464 27212 10470
rect 26976 10406 27028 10412
rect 27066 10432 27122 10441
rect 26988 10305 27016 10406
rect 27160 10406 27212 10412
rect 27066 10367 27122 10376
rect 26974 10296 27030 10305
rect 26974 10231 27030 10240
rect 26988 9994 27016 10231
rect 27172 9994 27200 10406
rect 27264 10130 27292 10764
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 26976 9988 27028 9994
rect 26976 9930 27028 9936
rect 27160 9988 27212 9994
rect 27160 9930 27212 9936
rect 26984 9820 27292 9829
rect 26984 9818 26990 9820
rect 27046 9818 27070 9820
rect 27126 9818 27150 9820
rect 27206 9818 27230 9820
rect 27286 9818 27292 9820
rect 27046 9766 27048 9818
rect 27228 9766 27230 9818
rect 26984 9764 26990 9766
rect 27046 9764 27070 9766
rect 27126 9764 27150 9766
rect 27206 9764 27230 9766
rect 27286 9764 27292 9766
rect 26984 9755 27292 9764
rect 27160 9648 27212 9654
rect 27160 9590 27212 9596
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26988 9353 27016 9522
rect 27172 9518 27200 9590
rect 27356 9518 27384 12804
rect 27540 12764 27568 14282
rect 27908 13734 27936 14572
rect 28092 14278 28120 15456
rect 28172 15438 28224 15444
rect 28264 15496 28316 15502
rect 28368 15473 28396 15506
rect 28264 15438 28316 15444
rect 28354 15464 28410 15473
rect 28172 14952 28224 14958
rect 28172 14894 28224 14900
rect 28184 14414 28212 14894
rect 28276 14521 28304 15438
rect 28354 15399 28410 15408
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28368 14890 28396 15302
rect 28448 15088 28500 15094
rect 28448 15030 28500 15036
rect 28460 14929 28488 15030
rect 28552 15026 28580 18022
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28644 16969 28672 17478
rect 28630 16960 28686 16969
rect 28630 16895 28686 16904
rect 28644 16046 28672 16895
rect 28736 16794 28764 18226
rect 29012 17882 29040 18226
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 28998 17096 29054 17105
rect 28908 17060 28960 17066
rect 28998 17031 29054 17040
rect 28908 17002 28960 17008
rect 28816 16992 28868 16998
rect 28816 16934 28868 16940
rect 28828 16794 28856 16934
rect 28920 16833 28948 17002
rect 28906 16824 28962 16833
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 28816 16788 28868 16794
rect 28906 16759 28908 16768
rect 28816 16730 28868 16736
rect 28960 16759 28962 16768
rect 28908 16730 28960 16736
rect 28736 16674 28764 16730
rect 28906 16688 28962 16697
rect 28736 16646 28856 16674
rect 28724 16244 28776 16250
rect 28724 16186 28776 16192
rect 28632 16040 28684 16046
rect 28632 15982 28684 15988
rect 28632 15904 28684 15910
rect 28632 15846 28684 15852
rect 28644 15502 28672 15846
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28446 14920 28502 14929
rect 28356 14884 28408 14890
rect 28446 14855 28502 14864
rect 28356 14826 28408 14832
rect 28262 14512 28318 14521
rect 28262 14447 28318 14456
rect 28356 14476 28408 14482
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 28080 14272 28132 14278
rect 28080 14214 28132 14220
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27644 13628 27952 13637
rect 27644 13626 27650 13628
rect 27706 13626 27730 13628
rect 27786 13626 27810 13628
rect 27866 13626 27890 13628
rect 27946 13626 27952 13628
rect 27706 13574 27708 13626
rect 27888 13574 27890 13626
rect 27644 13572 27650 13574
rect 27706 13572 27730 13574
rect 27786 13572 27810 13574
rect 27866 13572 27890 13574
rect 27946 13572 27952 13574
rect 27644 13563 27952 13572
rect 27804 13456 27856 13462
rect 27804 13398 27856 13404
rect 27896 13456 27948 13462
rect 27896 13398 27948 13404
rect 27620 13388 27672 13394
rect 27620 13330 27672 13336
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27632 13161 27660 13330
rect 27618 13152 27674 13161
rect 27618 13087 27674 13096
rect 27448 12736 27568 12764
rect 27448 12288 27476 12736
rect 27632 12696 27660 13087
rect 27724 12918 27752 13330
rect 27712 12912 27764 12918
rect 27712 12854 27764 12860
rect 27816 12782 27844 13398
rect 27908 13258 27936 13398
rect 28000 13297 28028 14214
rect 28172 14000 28224 14006
rect 28172 13942 28224 13948
rect 28080 13524 28132 13530
rect 28080 13466 28132 13472
rect 27986 13288 28042 13297
rect 27896 13252 27948 13258
rect 27986 13223 28042 13232
rect 27896 13194 27948 13200
rect 27988 13184 28040 13190
rect 27988 13126 28040 13132
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27540 12668 27660 12696
rect 27540 12356 27568 12668
rect 27644 12540 27952 12549
rect 27644 12538 27650 12540
rect 27706 12538 27730 12540
rect 27786 12538 27810 12540
rect 27866 12538 27890 12540
rect 27946 12538 27952 12540
rect 27706 12486 27708 12538
rect 27888 12486 27890 12538
rect 27644 12484 27650 12486
rect 27706 12484 27730 12486
rect 27786 12484 27810 12486
rect 27866 12484 27890 12486
rect 27946 12484 27952 12486
rect 27644 12475 27952 12484
rect 28000 12434 28028 13126
rect 28092 12832 28120 13466
rect 28184 13394 28212 13942
rect 28276 13870 28304 14447
rect 28356 14418 28408 14424
rect 28632 14476 28684 14482
rect 28736 14464 28764 16186
rect 28684 14436 28764 14464
rect 28632 14418 28684 14424
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28172 13388 28224 13394
rect 28224 13348 28304 13376
rect 28172 13330 28224 13336
rect 28092 12804 28212 12832
rect 28078 12744 28134 12753
rect 28078 12679 28134 12688
rect 27908 12406 28028 12434
rect 27620 12368 27672 12374
rect 27540 12328 27620 12356
rect 27620 12310 27672 12316
rect 27448 12260 27568 12288
rect 27436 12164 27488 12170
rect 27436 12106 27488 12112
rect 27448 11558 27476 12106
rect 27540 11626 27568 12260
rect 27632 12209 27660 12310
rect 27618 12200 27674 12209
rect 27618 12135 27674 12144
rect 27804 12096 27856 12102
rect 27804 12038 27856 12044
rect 27710 11928 27766 11937
rect 27710 11863 27766 11872
rect 27724 11762 27752 11863
rect 27712 11756 27764 11762
rect 27712 11698 27764 11704
rect 27816 11665 27844 12038
rect 27908 11694 27936 12406
rect 27986 12336 28042 12345
rect 28092 12306 28120 12679
rect 27986 12271 28042 12280
rect 28080 12300 28132 12306
rect 27896 11688 27948 11694
rect 27618 11656 27674 11665
rect 27528 11620 27580 11626
rect 27618 11591 27674 11600
rect 27802 11656 27858 11665
rect 27896 11630 27948 11636
rect 27802 11591 27858 11600
rect 27528 11562 27580 11568
rect 27436 11552 27488 11558
rect 27436 11494 27488 11500
rect 27436 11348 27488 11354
rect 27540 11336 27568 11562
rect 27632 11558 27660 11591
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27644 11452 27952 11461
rect 27644 11450 27650 11452
rect 27706 11450 27730 11452
rect 27786 11450 27810 11452
rect 27866 11450 27890 11452
rect 27946 11450 27952 11452
rect 27706 11398 27708 11450
rect 27888 11398 27890 11450
rect 27644 11396 27650 11398
rect 27706 11396 27730 11398
rect 27786 11396 27810 11398
rect 27866 11396 27890 11398
rect 27946 11396 27952 11398
rect 27644 11387 27952 11396
rect 28000 11354 28028 12271
rect 28080 12242 28132 12248
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 27488 11308 27568 11336
rect 27988 11348 28040 11354
rect 27436 11290 27488 11296
rect 27988 11290 28040 11296
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 26974 9344 27030 9353
rect 26974 9279 27030 9288
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26792 8968 26844 8974
rect 26792 8910 26844 8916
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 26712 8401 26740 8842
rect 26804 8548 26832 8910
rect 26988 8820 27016 9279
rect 27344 9036 27396 9042
rect 27448 9024 27476 11290
rect 27804 11280 27856 11286
rect 27526 11248 27582 11257
rect 27856 11240 27936 11268
rect 27804 11222 27856 11228
rect 27526 11183 27528 11192
rect 27580 11183 27582 11192
rect 27712 11212 27764 11218
rect 27528 11154 27580 11160
rect 27712 11154 27764 11160
rect 27618 11112 27674 11121
rect 27724 11082 27752 11154
rect 27618 11047 27674 11056
rect 27712 11076 27764 11082
rect 27528 11008 27580 11014
rect 27528 10950 27580 10956
rect 27540 10538 27568 10950
rect 27632 10724 27660 11047
rect 27712 11018 27764 11024
rect 27712 10736 27764 10742
rect 27632 10696 27712 10724
rect 27712 10678 27764 10684
rect 27908 10606 27936 11240
rect 28092 10810 28120 11834
rect 28184 11744 28212 12804
rect 28276 11898 28304 13348
rect 28368 12374 28396 14418
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28460 14006 28488 14214
rect 28644 14074 28672 14418
rect 28828 14074 28856 16646
rect 28906 16623 28962 16632
rect 28920 16153 28948 16623
rect 29012 16522 29040 17031
rect 29000 16516 29052 16522
rect 29000 16458 29052 16464
rect 28906 16144 28962 16153
rect 28906 16079 28962 16088
rect 28908 16040 28960 16046
rect 28908 15982 28960 15988
rect 28920 15434 28948 15982
rect 28908 15428 28960 15434
rect 28908 15370 28960 15376
rect 28920 14482 28948 15370
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 29012 15201 29040 15302
rect 28998 15192 29054 15201
rect 28998 15127 29054 15136
rect 29104 14618 29132 18362
rect 29184 18148 29236 18154
rect 29184 18090 29236 18096
rect 29276 18148 29328 18154
rect 29276 18090 29328 18096
rect 29196 17066 29224 18090
rect 29288 17338 29316 18090
rect 29276 17332 29328 17338
rect 29276 17274 29328 17280
rect 29276 17128 29328 17134
rect 29274 17096 29276 17105
rect 29328 17096 29330 17105
rect 29184 17060 29236 17066
rect 29274 17031 29330 17040
rect 29184 17002 29236 17008
rect 29274 16552 29330 16561
rect 29274 16487 29330 16496
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29196 16182 29224 16390
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29196 15570 29224 16118
rect 29288 15706 29316 16487
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29274 15600 29330 15609
rect 29184 15564 29236 15570
rect 29274 15535 29330 15544
rect 29184 15506 29236 15512
rect 29196 14822 29224 15506
rect 29288 15366 29316 15535
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29380 15162 29408 19858
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29460 19780 29512 19786
rect 29460 19722 29512 19728
rect 29472 19281 29500 19722
rect 29458 19272 29514 19281
rect 29458 19207 29514 19216
rect 29472 18873 29500 19207
rect 29656 18902 29684 19790
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29748 19417 29776 19654
rect 29734 19408 29790 19417
rect 29734 19343 29790 19352
rect 29734 19136 29790 19145
rect 29734 19071 29790 19080
rect 29644 18896 29696 18902
rect 29458 18864 29514 18873
rect 29644 18838 29696 18844
rect 29748 18834 29776 19071
rect 29458 18799 29514 18808
rect 29736 18828 29788 18834
rect 29736 18770 29788 18776
rect 29644 18692 29696 18698
rect 29644 18634 29696 18640
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29472 17338 29500 18362
rect 29656 17814 29684 18634
rect 29748 18426 29776 18770
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29736 18148 29788 18154
rect 29736 18090 29788 18096
rect 29748 18057 29776 18090
rect 29734 18048 29790 18057
rect 29734 17983 29790 17992
rect 29644 17808 29696 17814
rect 29644 17750 29696 17756
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29550 17368 29606 17377
rect 29460 17332 29512 17338
rect 29550 17303 29606 17312
rect 29460 17274 29512 17280
rect 29458 17232 29514 17241
rect 29458 17167 29514 17176
rect 29472 16590 29500 17167
rect 29564 16726 29592 17303
rect 29552 16720 29604 16726
rect 29552 16662 29604 16668
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29552 16448 29604 16454
rect 29552 16390 29604 16396
rect 29564 16289 29592 16390
rect 29550 16280 29606 16289
rect 29550 16215 29606 16224
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29458 16008 29514 16017
rect 29458 15943 29460 15952
rect 29512 15943 29514 15952
rect 29460 15914 29512 15920
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29276 14952 29328 14958
rect 29274 14920 29276 14929
rect 29328 14920 29330 14929
rect 29274 14855 29330 14864
rect 29184 14816 29236 14822
rect 29184 14758 29236 14764
rect 29092 14612 29144 14618
rect 29092 14554 29144 14560
rect 28908 14476 28960 14482
rect 28908 14418 28960 14424
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28816 14068 28868 14074
rect 28816 14010 28868 14016
rect 28448 14000 28500 14006
rect 28828 13977 28856 14010
rect 28448 13942 28500 13948
rect 28814 13968 28870 13977
rect 28814 13903 28870 13912
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 28448 13728 28500 13734
rect 28448 13670 28500 13676
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28460 13394 28488 13670
rect 28448 13388 28500 13394
rect 28448 13330 28500 13336
rect 28920 13326 28948 13670
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28736 12782 28764 13262
rect 29012 12986 29040 13398
rect 29104 13190 29132 13806
rect 29092 13184 29144 13190
rect 29196 13161 29224 14758
rect 29368 13796 29420 13802
rect 29368 13738 29420 13744
rect 29380 13462 29408 13738
rect 29368 13456 29420 13462
rect 29368 13398 29420 13404
rect 29092 13126 29144 13132
rect 29182 13152 29238 13161
rect 29182 13087 29238 13096
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 28632 12776 28684 12782
rect 28632 12718 28684 12724
rect 28724 12776 28776 12782
rect 29184 12776 29236 12782
rect 28724 12718 28776 12724
rect 28906 12744 28962 12753
rect 28356 12368 28408 12374
rect 28408 12328 28580 12356
rect 28356 12310 28408 12316
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28368 11830 28396 12174
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 28184 11716 28304 11744
rect 28170 11656 28226 11665
rect 28276 11626 28304 11716
rect 28356 11688 28408 11694
rect 28356 11630 28408 11636
rect 28170 11591 28226 11600
rect 28264 11620 28316 11626
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 27896 10600 27948 10606
rect 27896 10542 27948 10548
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 27644 10364 27952 10373
rect 27644 10362 27650 10364
rect 27706 10362 27730 10364
rect 27786 10362 27810 10364
rect 27866 10362 27890 10364
rect 27946 10362 27952 10364
rect 27706 10310 27708 10362
rect 27888 10310 27890 10362
rect 27644 10308 27650 10310
rect 27706 10308 27730 10310
rect 27786 10308 27810 10310
rect 27866 10308 27890 10310
rect 27946 10308 27952 10310
rect 27644 10299 27952 10308
rect 27986 10160 28042 10169
rect 27528 10124 27580 10130
rect 27986 10095 28042 10104
rect 27528 10066 27580 10072
rect 27540 9586 27568 10066
rect 28000 10062 28028 10095
rect 27988 10056 28040 10062
rect 27618 10024 27674 10033
rect 27988 9998 28040 10004
rect 28092 10010 28120 10406
rect 28184 10130 28212 11591
rect 28264 11562 28316 11568
rect 28368 11354 28396 11630
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 28262 11248 28318 11257
rect 28262 11183 28264 11192
rect 28316 11183 28318 11192
rect 28264 11154 28316 11160
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 28276 10062 28304 11154
rect 28460 10538 28488 11834
rect 28552 11762 28580 12328
rect 28644 12170 28672 12718
rect 28736 12306 28764 12718
rect 29184 12718 29236 12724
rect 28906 12679 28962 12688
rect 28724 12300 28776 12306
rect 28920 12288 28948 12679
rect 29196 12481 29224 12718
rect 29182 12472 29238 12481
rect 29182 12407 29238 12416
rect 29092 12368 29144 12374
rect 29090 12336 29092 12345
rect 29144 12336 29146 12345
rect 29380 12322 29408 12922
rect 28920 12260 29040 12288
rect 29090 12271 29146 12280
rect 29196 12294 29408 12322
rect 28724 12242 28776 12248
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28540 11756 28592 11762
rect 28540 11698 28592 11704
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28448 10532 28500 10538
rect 28448 10474 28500 10480
rect 28264 10056 28316 10062
rect 28092 9982 28212 10010
rect 28264 9998 28316 10004
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 27618 9959 27674 9968
rect 27632 9722 27660 9959
rect 28080 9920 28132 9926
rect 28080 9862 28132 9868
rect 27620 9716 27672 9722
rect 27620 9658 27672 9664
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27724 9586 27752 9658
rect 27986 9616 28042 9625
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 27712 9580 27764 9586
rect 27986 9551 27988 9560
rect 27712 9522 27764 9528
rect 28040 9551 28042 9560
rect 27988 9522 28040 9528
rect 27644 9276 27952 9285
rect 27644 9274 27650 9276
rect 27706 9274 27730 9276
rect 27786 9274 27810 9276
rect 27866 9274 27890 9276
rect 27946 9274 27952 9276
rect 27706 9222 27708 9274
rect 27888 9222 27890 9274
rect 27644 9220 27650 9222
rect 27706 9220 27730 9222
rect 27786 9220 27810 9222
rect 27866 9220 27890 9222
rect 27946 9220 27952 9222
rect 27644 9211 27952 9220
rect 27528 9172 27580 9178
rect 27580 9132 27752 9160
rect 27528 9114 27580 9120
rect 27620 9036 27672 9042
rect 27396 8996 27476 9024
rect 27540 8996 27620 9024
rect 27344 8978 27396 8984
rect 27540 8945 27568 8996
rect 27620 8978 27672 8984
rect 27724 8974 27752 9132
rect 27712 8968 27764 8974
rect 27526 8936 27582 8945
rect 27436 8900 27488 8906
rect 27712 8910 27764 8916
rect 28092 8922 28120 9862
rect 28184 9024 28212 9982
rect 28276 9178 28304 9998
rect 28368 9178 28396 9998
rect 28460 9382 28488 10474
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 28446 9208 28502 9217
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28356 9172 28408 9178
rect 28446 9143 28502 9152
rect 28356 9114 28408 9120
rect 28356 9036 28408 9042
rect 28184 8996 28304 9024
rect 28092 8894 28212 8922
rect 27526 8871 27582 8880
rect 27436 8842 27488 8848
rect 26896 8792 27016 8820
rect 26896 8616 26924 8792
rect 26984 8732 27292 8741
rect 26984 8730 26990 8732
rect 27046 8730 27070 8732
rect 27126 8730 27150 8732
rect 27206 8730 27230 8732
rect 27286 8730 27292 8732
rect 27046 8678 27048 8730
rect 27228 8678 27230 8730
rect 26984 8676 26990 8678
rect 27046 8676 27070 8678
rect 27126 8676 27150 8678
rect 27206 8676 27230 8678
rect 27286 8676 27292 8678
rect 26984 8667 27292 8676
rect 27344 8628 27396 8634
rect 26896 8588 27292 8616
rect 26804 8520 26924 8548
rect 26698 8392 26754 8401
rect 26698 8327 26754 8336
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26698 8120 26754 8129
rect 26698 8055 26754 8064
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26620 5370 26648 6258
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26620 5166 26648 5306
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26712 4622 26740 8055
rect 26804 7274 26832 8230
rect 26896 7954 26924 8520
rect 26974 8528 27030 8537
rect 26974 8463 27030 8472
rect 26988 7954 27016 8463
rect 27264 8362 27292 8588
rect 27344 8570 27396 8576
rect 27068 8356 27120 8362
rect 27068 8298 27120 8304
rect 27252 8356 27304 8362
rect 27252 8298 27304 8304
rect 27080 8265 27108 8298
rect 27066 8256 27122 8265
rect 27066 8191 27122 8200
rect 26884 7948 26936 7954
rect 26884 7890 26936 7896
rect 26976 7948 27028 7954
rect 26976 7890 27028 7896
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26804 5710 26832 7210
rect 26896 6934 26924 7890
rect 26984 7644 27292 7653
rect 26984 7642 26990 7644
rect 27046 7642 27070 7644
rect 27126 7642 27150 7644
rect 27206 7642 27230 7644
rect 27286 7642 27292 7644
rect 27046 7590 27048 7642
rect 27228 7590 27230 7642
rect 26984 7588 26990 7590
rect 27046 7588 27070 7590
rect 27126 7588 27150 7590
rect 27206 7588 27230 7590
rect 27286 7588 27292 7590
rect 26984 7579 27292 7588
rect 27356 7342 27384 8570
rect 27448 8362 27476 8842
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 28080 8832 28132 8838
rect 28080 8774 28132 8780
rect 27540 8566 27568 8774
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 27528 8560 27580 8566
rect 27908 8537 27936 8570
rect 27528 8502 27580 8508
rect 27894 8528 27950 8537
rect 27894 8463 27950 8472
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27802 8392 27858 8401
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27344 7336 27396 7342
rect 27436 7336 27488 7342
rect 27344 7278 27396 7284
rect 27434 7304 27436 7313
rect 27488 7304 27490 7313
rect 26884 6928 26936 6934
rect 26884 6870 26936 6876
rect 26896 6254 26924 6870
rect 27080 6730 27108 7278
rect 27434 7239 27490 7248
rect 27344 6792 27396 6798
rect 27344 6734 27396 6740
rect 27068 6724 27120 6730
rect 27068 6666 27120 6672
rect 26984 6556 27292 6565
rect 26984 6554 26990 6556
rect 27046 6554 27070 6556
rect 27126 6554 27150 6556
rect 27206 6554 27230 6556
rect 27286 6554 27292 6556
rect 27046 6502 27048 6554
rect 27228 6502 27230 6554
rect 26984 6500 26990 6502
rect 27046 6500 27070 6502
rect 27126 6500 27150 6502
rect 27206 6500 27230 6502
rect 27286 6500 27292 6502
rect 26984 6491 27292 6500
rect 27356 6458 27384 6734
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 26884 6248 26936 6254
rect 26884 6190 26936 6196
rect 26976 6180 27028 6186
rect 26976 6122 27028 6128
rect 26988 5846 27016 6122
rect 27356 5846 27384 6394
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 27344 5840 27396 5846
rect 27344 5782 27396 5788
rect 26884 5772 26936 5778
rect 26884 5714 26936 5720
rect 26792 5704 26844 5710
rect 26896 5681 26924 5714
rect 26792 5646 26844 5652
rect 26882 5672 26938 5681
rect 26882 5607 26884 5616
rect 26936 5607 26938 5616
rect 26884 5578 26936 5584
rect 26984 5468 27292 5477
rect 26984 5466 26990 5468
rect 27046 5466 27070 5468
rect 27126 5466 27150 5468
rect 27206 5466 27230 5468
rect 27286 5466 27292 5468
rect 27046 5414 27048 5466
rect 27228 5414 27230 5466
rect 26984 5412 26990 5414
rect 27046 5412 27070 5414
rect 27126 5412 27150 5414
rect 27206 5412 27230 5414
rect 27286 5412 27292 5414
rect 26984 5403 27292 5412
rect 27448 4690 27476 5850
rect 27540 5710 27568 8366
rect 27802 8327 27858 8336
rect 27816 8294 27844 8327
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27644 8188 27952 8197
rect 27644 8186 27650 8188
rect 27706 8186 27730 8188
rect 27786 8186 27810 8188
rect 27866 8186 27890 8188
rect 27946 8186 27952 8188
rect 27706 8134 27708 8186
rect 27888 8134 27890 8186
rect 27644 8132 27650 8134
rect 27706 8132 27730 8134
rect 27786 8132 27810 8134
rect 27866 8132 27890 8134
rect 27946 8132 27952 8134
rect 27644 8123 27952 8132
rect 28000 8072 28028 8434
rect 27908 8044 28028 8072
rect 27908 7954 27936 8044
rect 27896 7948 27948 7954
rect 27896 7890 27948 7896
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 27908 7256 27936 7890
rect 28000 7857 28028 7890
rect 28092 7886 28120 8774
rect 28080 7880 28132 7886
rect 27986 7848 28042 7857
rect 28080 7822 28132 7828
rect 27986 7783 28042 7792
rect 27988 7268 28040 7274
rect 27908 7228 27988 7256
rect 27988 7210 28040 7216
rect 27644 7100 27952 7109
rect 27644 7098 27650 7100
rect 27706 7098 27730 7100
rect 27786 7098 27810 7100
rect 27866 7098 27890 7100
rect 27946 7098 27952 7100
rect 27706 7046 27708 7098
rect 27888 7046 27890 7098
rect 27644 7044 27650 7046
rect 27706 7044 27730 7046
rect 27786 7044 27810 7046
rect 27866 7044 27890 7046
rect 27946 7044 27952 7046
rect 27644 7035 27952 7044
rect 27644 6012 27952 6021
rect 27644 6010 27650 6012
rect 27706 6010 27730 6012
rect 27786 6010 27810 6012
rect 27866 6010 27890 6012
rect 27946 6010 27952 6012
rect 27706 5958 27708 6010
rect 27888 5958 27890 6010
rect 27644 5956 27650 5958
rect 27706 5956 27730 5958
rect 27786 5956 27810 5958
rect 27866 5956 27890 5958
rect 27946 5956 27952 5958
rect 27644 5947 27952 5956
rect 28000 5778 28028 7210
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 27724 5166 27752 5714
rect 28092 5302 28120 7822
rect 28184 7818 28212 8894
rect 28276 8362 28304 8996
rect 28356 8978 28408 8984
rect 28264 8356 28316 8362
rect 28264 8298 28316 8304
rect 28172 7812 28224 7818
rect 28172 7754 28224 7760
rect 28170 7712 28226 7721
rect 28170 7647 28226 7656
rect 28184 7274 28212 7647
rect 28172 7268 28224 7274
rect 28172 7210 28224 7216
rect 28184 6730 28212 7210
rect 28172 6724 28224 6730
rect 28172 6666 28224 6672
rect 28276 6458 28304 8298
rect 28368 7954 28396 8978
rect 28356 7948 28408 7954
rect 28356 7890 28408 7896
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28368 7546 28396 7754
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28368 6934 28396 7482
rect 28356 6928 28408 6934
rect 28356 6870 28408 6876
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28460 6254 28488 9143
rect 28552 7546 28580 11562
rect 28644 10470 28672 12106
rect 28736 12084 28764 12242
rect 28736 12056 28856 12084
rect 28724 11892 28776 11898
rect 28724 11834 28776 11840
rect 28736 11218 28764 11834
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 28630 9616 28686 9625
rect 28630 9551 28686 9560
rect 28644 8294 28672 9551
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28736 8090 28764 11154
rect 28828 11014 28856 12056
rect 29012 11694 29040 12260
rect 29000 11688 29052 11694
rect 29196 11642 29224 12294
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29274 11928 29330 11937
rect 29274 11863 29330 11872
rect 29000 11630 29052 11636
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 29104 11614 29224 11642
rect 28816 11008 28868 11014
rect 28816 10950 28868 10956
rect 28816 10464 28868 10470
rect 28816 10406 28868 10412
rect 28828 9994 28856 10406
rect 28816 9988 28868 9994
rect 28816 9930 28868 9936
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 28630 7984 28686 7993
rect 28630 7919 28632 7928
rect 28684 7919 28686 7928
rect 28632 7890 28684 7896
rect 28540 7540 28592 7546
rect 28540 7482 28592 7488
rect 28552 6866 28580 7482
rect 28828 7410 28856 9930
rect 28920 9042 28948 11562
rect 29104 11558 29132 11614
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29184 11552 29236 11558
rect 29184 11494 29236 11500
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 29012 9722 29040 10542
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 29104 9330 29132 11494
rect 29196 10674 29224 11494
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29288 10606 29316 11863
rect 29380 11132 29408 12174
rect 29472 11694 29500 15914
rect 29564 15706 29592 16050
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29552 15564 29604 15570
rect 29552 15506 29604 15512
rect 29564 15434 29592 15506
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29550 15056 29606 15065
rect 29550 14991 29552 15000
rect 29604 14991 29606 15000
rect 29552 14962 29604 14968
rect 29656 14890 29684 17614
rect 29748 17066 29776 17983
rect 29736 17060 29788 17066
rect 29736 17002 29788 17008
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 29748 15552 29776 16594
rect 29840 16250 29868 19910
rect 29920 19916 29972 19922
rect 29920 19858 29972 19864
rect 29932 18970 29960 19858
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 30024 18970 30052 19450
rect 30208 19281 30236 20878
rect 30300 20754 30328 21830
rect 30564 21412 30616 21418
rect 30564 21354 30616 21360
rect 30576 21146 30604 21354
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30852 21185 30880 21286
rect 30838 21176 30894 21185
rect 30564 21140 30616 21146
rect 30838 21111 30894 21120
rect 30564 21082 30616 21088
rect 30300 20726 30420 20754
rect 30288 20596 30340 20602
rect 30288 20538 30340 20544
rect 30300 19990 30328 20538
rect 30392 20534 30420 20726
rect 30380 20528 30432 20534
rect 30380 20470 30432 20476
rect 30576 20398 30604 21082
rect 30944 21078 30972 21898
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 30932 21072 30984 21078
rect 30932 21014 30984 21020
rect 31220 20942 31248 21422
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 30564 20392 30616 20398
rect 30840 20392 30892 20398
rect 30564 20334 30616 20340
rect 30838 20360 30840 20369
rect 30892 20360 30894 20369
rect 30288 19984 30340 19990
rect 30288 19926 30340 19932
rect 30194 19272 30250 19281
rect 30194 19207 30250 19216
rect 29920 18964 29972 18970
rect 29920 18906 29972 18912
rect 30012 18964 30064 18970
rect 30012 18906 30064 18912
rect 30024 18850 30052 18906
rect 29932 18822 30052 18850
rect 30300 18834 30328 19926
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30288 18828 30340 18834
rect 29932 18766 29960 18822
rect 30288 18770 30340 18776
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 29828 16244 29880 16250
rect 29828 16186 29880 16192
rect 29828 15564 29880 15570
rect 29748 15524 29828 15552
rect 29828 15506 29880 15512
rect 29736 15360 29788 15366
rect 29736 15302 29788 15308
rect 29644 14884 29696 14890
rect 29644 14826 29696 14832
rect 29748 14550 29776 15302
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29840 14482 29868 15506
rect 29932 14958 29960 18702
rect 30012 18284 30064 18290
rect 30116 18272 30144 18702
rect 30064 18244 30144 18272
rect 30012 18226 30064 18232
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30024 17202 30052 17682
rect 30116 17678 30144 18244
rect 30208 18086 30236 18702
rect 30484 18193 30512 19790
rect 30576 19310 30604 20334
rect 30838 20295 30894 20304
rect 30656 19780 30708 19786
rect 30656 19722 30708 19728
rect 30564 19304 30616 19310
rect 30564 19246 30616 19252
rect 30470 18184 30526 18193
rect 30470 18119 30526 18128
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30012 17196 30064 17202
rect 30012 17138 30064 17144
rect 30104 17060 30156 17066
rect 30104 17002 30156 17008
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 30024 15502 30052 16526
rect 30116 15858 30144 17002
rect 30208 15978 30236 17682
rect 30378 17640 30434 17649
rect 30378 17575 30434 17584
rect 30288 17536 30340 17542
rect 30288 17478 30340 17484
rect 30300 16658 30328 17478
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 30116 15830 30236 15858
rect 30208 15706 30236 15830
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29920 14816 29972 14822
rect 29918 14784 29920 14793
rect 29972 14784 29974 14793
rect 29918 14719 29974 14728
rect 30024 14482 30052 15438
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 30012 14476 30064 14482
rect 30012 14418 30064 14424
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29552 13728 29604 13734
rect 29552 13670 29604 13676
rect 29564 13258 29592 13670
rect 29644 13388 29696 13394
rect 29644 13330 29696 13336
rect 29552 13252 29604 13258
rect 29552 13194 29604 13200
rect 29656 12714 29684 13330
rect 29644 12708 29696 12714
rect 29644 12650 29696 12656
rect 29460 11688 29512 11694
rect 29460 11630 29512 11636
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29564 11354 29592 11630
rect 29644 11552 29696 11558
rect 29644 11494 29696 11500
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29656 11286 29684 11494
rect 29644 11280 29696 11286
rect 29644 11222 29696 11228
rect 29748 11218 29776 14282
rect 29840 12889 29868 14418
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 29932 12918 29960 13126
rect 29920 12912 29972 12918
rect 29826 12880 29882 12889
rect 29920 12854 29972 12860
rect 29826 12815 29882 12824
rect 29840 11762 29868 12815
rect 29932 12374 29960 12854
rect 29920 12368 29972 12374
rect 29920 12310 29972 12316
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 30024 11694 30052 14418
rect 30116 13802 30144 15642
rect 30300 15450 30328 16594
rect 30392 16046 30420 17575
rect 30472 16992 30524 16998
rect 30472 16934 30524 16940
rect 30484 16658 30512 16934
rect 30472 16652 30524 16658
rect 30472 16594 30524 16600
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30380 15564 30432 15570
rect 30380 15506 30432 15512
rect 30392 15473 30420 15506
rect 30208 15422 30328 15450
rect 30378 15464 30434 15473
rect 30208 14482 30236 15422
rect 30484 15434 30512 16594
rect 30562 16416 30618 16425
rect 30562 16351 30618 16360
rect 30378 15399 30434 15408
rect 30472 15428 30524 15434
rect 30288 15360 30340 15366
rect 30286 15328 30288 15337
rect 30340 15328 30342 15337
rect 30286 15263 30342 15272
rect 30286 15192 30342 15201
rect 30286 15127 30342 15136
rect 30300 15094 30328 15127
rect 30288 15088 30340 15094
rect 30288 15030 30340 15036
rect 30392 14958 30420 15399
rect 30472 15370 30524 15376
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30208 13870 30236 14418
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 30104 13796 30156 13802
rect 30104 13738 30156 13744
rect 30104 13456 30156 13462
rect 30104 13398 30156 13404
rect 30012 11688 30064 11694
rect 30012 11630 30064 11636
rect 30116 11540 30144 13398
rect 30208 12434 30236 13806
rect 30300 13734 30328 14214
rect 30392 13841 30420 14758
rect 30484 14482 30512 15370
rect 30576 14958 30604 16351
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30668 14618 30696 19722
rect 31220 19689 31248 20878
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31206 19680 31262 19689
rect 31206 19615 31262 19624
rect 30930 19272 30986 19281
rect 30930 19207 30986 19216
rect 31024 19236 31076 19242
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30760 18970 30788 19110
rect 30748 18964 30800 18970
rect 30748 18906 30800 18912
rect 30840 18964 30892 18970
rect 30840 18906 30892 18912
rect 30852 18698 30880 18906
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30746 18456 30802 18465
rect 30944 18426 30972 19207
rect 31024 19178 31076 19184
rect 31116 19236 31168 19242
rect 31116 19178 31168 19184
rect 31036 18902 31064 19178
rect 31024 18896 31076 18902
rect 31024 18838 31076 18844
rect 31128 18834 31156 19178
rect 31116 18828 31168 18834
rect 31116 18770 31168 18776
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 31036 18630 31064 18702
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 30746 18391 30802 18400
rect 30932 18420 30984 18426
rect 30760 18358 30788 18391
rect 30932 18362 30984 18368
rect 30748 18352 30800 18358
rect 30748 18294 30800 18300
rect 30838 18184 30894 18193
rect 30838 18119 30894 18128
rect 30748 17332 30800 17338
rect 30748 17274 30800 17280
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30760 14074 30788 17274
rect 30852 15570 30880 18119
rect 30944 16046 30972 18362
rect 31128 18290 31156 18770
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 31220 18154 31248 19615
rect 31312 18630 31340 19858
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31312 18329 31340 18566
rect 31298 18320 31354 18329
rect 31298 18255 31354 18264
rect 31208 18148 31260 18154
rect 31208 18090 31260 18096
rect 31404 18086 31432 21422
rect 31574 20360 31630 20369
rect 31574 20295 31630 20304
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31496 18737 31524 18770
rect 31482 18728 31538 18737
rect 31482 18663 31538 18672
rect 31392 18080 31444 18086
rect 31392 18022 31444 18028
rect 31114 17640 31170 17649
rect 31114 17575 31170 17584
rect 31128 17338 31156 17575
rect 31116 17332 31168 17338
rect 31116 17274 31168 17280
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 30932 16040 30984 16046
rect 30932 15982 30984 15988
rect 30840 15564 30892 15570
rect 30840 15506 30892 15512
rect 30852 14346 30880 15506
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 30944 14482 30972 15098
rect 30932 14476 30984 14482
rect 30932 14418 30984 14424
rect 30840 14340 30892 14346
rect 30840 14282 30892 14288
rect 30748 14068 30800 14074
rect 30748 14010 30800 14016
rect 30656 13932 30708 13938
rect 30656 13874 30708 13880
rect 30378 13832 30434 13841
rect 30378 13767 30434 13776
rect 30288 13728 30340 13734
rect 30288 13670 30340 13676
rect 30300 13161 30328 13670
rect 30286 13152 30342 13161
rect 30286 13087 30342 13096
rect 30208 12406 30328 12434
rect 30300 12238 30328 12406
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 30300 11694 30328 12174
rect 30668 11937 30696 13874
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30852 12782 30880 13262
rect 30748 12776 30800 12782
rect 30748 12718 30800 12724
rect 30840 12776 30892 12782
rect 30840 12718 30892 12724
rect 30654 11928 30710 11937
rect 30654 11863 30710 11872
rect 30472 11824 30524 11830
rect 30472 11766 30524 11772
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 30024 11512 30144 11540
rect 29736 11212 29788 11218
rect 29736 11154 29788 11160
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 29460 11144 29512 11150
rect 29380 11104 29460 11132
rect 29460 11086 29512 11092
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29184 10532 29236 10538
rect 29184 10474 29236 10480
rect 29196 10198 29224 10474
rect 29472 10248 29500 11086
rect 29932 11082 29960 11154
rect 29920 11076 29972 11082
rect 29920 11018 29972 11024
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 29380 10220 29592 10248
rect 29184 10192 29236 10198
rect 29184 10134 29236 10140
rect 29276 10056 29328 10062
rect 29276 9998 29328 10004
rect 29184 9580 29236 9586
rect 29184 9522 29236 9528
rect 29012 9302 29132 9330
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 29012 8906 29040 9302
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 29000 8900 29052 8906
rect 28920 8860 29000 8888
rect 28920 8294 28948 8860
rect 29000 8842 29052 8848
rect 28908 8288 28960 8294
rect 28908 8230 28960 8236
rect 29000 8288 29052 8294
rect 29000 8230 29052 8236
rect 29012 7818 29040 8230
rect 29000 7812 29052 7818
rect 29000 7754 29052 7760
rect 29104 7698 29132 9114
rect 29196 7886 29224 9522
rect 29288 9518 29316 9998
rect 29380 9518 29408 10220
rect 29564 10130 29592 10220
rect 29748 10130 29776 10950
rect 29932 10690 29960 11018
rect 29840 10662 29960 10690
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29552 10124 29604 10130
rect 29552 10066 29604 10072
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 29380 9178 29408 9454
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29472 9042 29500 10066
rect 29748 10010 29776 10066
rect 29564 9982 29776 10010
rect 29460 9036 29512 9042
rect 29460 8978 29512 8984
rect 29368 8900 29420 8906
rect 29368 8842 29420 8848
rect 29380 8498 29408 8842
rect 29564 8514 29592 9982
rect 29644 9920 29696 9926
rect 29644 9862 29696 9868
rect 29656 9704 29684 9862
rect 29656 9676 29776 9704
rect 29748 9518 29776 9676
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29656 9178 29684 9454
rect 29734 9344 29790 9353
rect 29734 9279 29790 9288
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 29368 8492 29420 8498
rect 29564 8486 29684 8514
rect 29368 8434 29420 8440
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 29458 8392 29514 8401
rect 29288 8265 29316 8366
rect 29458 8327 29514 8336
rect 29274 8256 29330 8265
rect 29274 8191 29330 8200
rect 29276 8016 29328 8022
rect 29276 7958 29328 7964
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 29012 7670 29132 7698
rect 28816 7404 28868 7410
rect 28816 7346 28868 7352
rect 28724 7336 28776 7342
rect 28724 7278 28776 7284
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28644 6866 28672 7142
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28736 6769 28764 7278
rect 29012 7206 29040 7670
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29092 7268 29144 7274
rect 29092 7210 29144 7216
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 6934 29040 7142
rect 29000 6928 29052 6934
rect 29000 6870 29052 6876
rect 28722 6760 28778 6769
rect 28722 6695 28778 6704
rect 28908 6724 28960 6730
rect 28908 6666 28960 6672
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28460 5914 28488 6190
rect 28448 5908 28500 5914
rect 28448 5850 28500 5856
rect 28460 5574 28488 5850
rect 28448 5568 28500 5574
rect 28448 5510 28500 5516
rect 28080 5296 28132 5302
rect 28080 5238 28132 5244
rect 27712 5160 27764 5166
rect 27712 5102 27764 5108
rect 28538 5128 28594 5137
rect 28538 5063 28594 5072
rect 28552 5030 28580 5063
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 27644 4924 27952 4933
rect 27644 4922 27650 4924
rect 27706 4922 27730 4924
rect 27786 4922 27810 4924
rect 27866 4922 27890 4924
rect 27946 4922 27952 4924
rect 27706 4870 27708 4922
rect 27888 4870 27890 4922
rect 27644 4868 27650 4870
rect 27706 4868 27730 4870
rect 27786 4868 27810 4870
rect 27866 4868 27890 4870
rect 27946 4868 27952 4870
rect 27644 4859 27952 4868
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 26700 4616 26752 4622
rect 26700 4558 26752 4564
rect 28552 4486 28580 4966
rect 28920 4554 28948 6666
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 29012 6322 29040 6598
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 28908 4548 28960 4554
rect 28908 4490 28960 4496
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 26984 4380 27292 4389
rect 26984 4378 26990 4380
rect 27046 4378 27070 4380
rect 27126 4378 27150 4380
rect 27206 4378 27230 4380
rect 27286 4378 27292 4380
rect 27046 4326 27048 4378
rect 27228 4326 27230 4378
rect 26984 4324 26990 4326
rect 27046 4324 27070 4326
rect 27126 4324 27150 4326
rect 27206 4324 27230 4326
rect 27286 4324 27292 4326
rect 26984 4315 27292 4324
rect 27644 3836 27952 3845
rect 27644 3834 27650 3836
rect 27706 3834 27730 3836
rect 27786 3834 27810 3836
rect 27866 3834 27890 3836
rect 27946 3834 27952 3836
rect 27706 3782 27708 3834
rect 27888 3782 27890 3834
rect 27644 3780 27650 3782
rect 27706 3780 27730 3782
rect 27786 3780 27810 3782
rect 27866 3780 27890 3782
rect 27946 3780 27952 3782
rect 27644 3771 27952 3780
rect 26984 3292 27292 3301
rect 26984 3290 26990 3292
rect 27046 3290 27070 3292
rect 27126 3290 27150 3292
rect 27206 3290 27230 3292
rect 27286 3290 27292 3292
rect 27046 3238 27048 3290
rect 27228 3238 27230 3290
rect 26984 3236 26990 3238
rect 27046 3236 27070 3238
rect 27126 3236 27150 3238
rect 27206 3236 27230 3238
rect 27286 3236 27292 3238
rect 26984 3227 27292 3236
rect 29012 3097 29040 6054
rect 29104 5778 29132 7210
rect 29196 7206 29224 7278
rect 29184 7200 29236 7206
rect 29184 7142 29236 7148
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29196 5914 29224 6190
rect 29184 5908 29236 5914
rect 29184 5850 29236 5856
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 29288 5642 29316 7958
rect 29472 7342 29500 8327
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29564 8090 29592 8230
rect 29656 8090 29684 8486
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29460 7336 29512 7342
rect 29460 7278 29512 7284
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29472 6225 29500 6802
rect 29458 6216 29514 6225
rect 29380 6174 29458 6202
rect 29276 5636 29328 5642
rect 29276 5578 29328 5584
rect 29288 5166 29316 5578
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 29380 4826 29408 6174
rect 29458 6151 29514 6160
rect 29564 5778 29592 7890
rect 29644 7744 29696 7750
rect 29748 7732 29776 9279
rect 29696 7704 29776 7732
rect 29644 7686 29696 7692
rect 29656 5817 29684 7686
rect 29840 7002 29868 10662
rect 29920 10192 29972 10198
rect 29920 10134 29972 10140
rect 29932 9042 29960 10134
rect 29920 9036 29972 9042
rect 29920 8978 29972 8984
rect 29932 8498 29960 8978
rect 30024 8514 30052 11512
rect 30380 10736 30432 10742
rect 30378 10704 30380 10713
rect 30432 10704 30434 10713
rect 30378 10639 30434 10648
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 10130 30144 10406
rect 30208 10266 30236 10542
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 30300 10198 30328 10542
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30104 10124 30156 10130
rect 30104 10066 30156 10072
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 30116 9330 30144 10066
rect 30208 9926 30236 10066
rect 30196 9920 30248 9926
rect 30196 9862 30248 9868
rect 30392 9704 30420 10639
rect 30300 9676 30420 9704
rect 30300 9636 30328 9676
rect 30208 9608 30328 9636
rect 30208 9518 30236 9608
rect 30196 9512 30248 9518
rect 30380 9512 30432 9518
rect 30196 9454 30248 9460
rect 30300 9460 30380 9466
rect 30300 9454 30432 9460
rect 30300 9438 30420 9454
rect 30300 9330 30328 9438
rect 30116 9302 30328 9330
rect 30300 9178 30328 9302
rect 30288 9172 30340 9178
rect 30288 9114 30340 9120
rect 30484 9058 30512 11766
rect 30564 11212 30616 11218
rect 30564 11154 30616 11160
rect 30208 9042 30512 9058
rect 30576 9042 30604 11154
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30104 9036 30156 9042
rect 30104 8978 30156 8984
rect 30196 9036 30512 9042
rect 30248 9030 30512 9036
rect 30564 9036 30616 9042
rect 30196 8978 30248 8984
rect 30564 8978 30616 8984
rect 30116 8634 30144 8978
rect 30380 8968 30432 8974
rect 30378 8936 30380 8945
rect 30432 8936 30434 8945
rect 30196 8900 30248 8906
rect 30378 8871 30434 8880
rect 30472 8900 30524 8906
rect 30196 8842 30248 8848
rect 30472 8842 30524 8848
rect 30208 8786 30236 8842
rect 30208 8758 30328 8786
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 29920 8492 29972 8498
rect 30024 8486 30236 8514
rect 29920 8434 29972 8440
rect 30012 8424 30064 8430
rect 29918 8392 29974 8401
rect 29974 8372 30012 8378
rect 29974 8366 30064 8372
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 29974 8350 30052 8366
rect 29918 8327 29974 8336
rect 30024 8090 30052 8350
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 30012 8084 30064 8090
rect 30012 8026 30064 8032
rect 29932 7954 29960 8026
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29828 6996 29880 7002
rect 29828 6938 29880 6944
rect 29840 6322 29868 6938
rect 29932 6644 29960 7890
rect 30012 7812 30064 7818
rect 30012 7754 30064 7760
rect 30024 6746 30052 7754
rect 30116 7546 30144 8366
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30116 7274 30144 7482
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 30116 6866 30144 7210
rect 30208 7206 30236 8486
rect 30300 8430 30328 8758
rect 30288 8424 30340 8430
rect 30340 8384 30420 8412
rect 30288 8366 30340 8372
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 30300 7410 30328 7754
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30104 6860 30156 6866
rect 30104 6802 30156 6808
rect 30024 6718 30144 6746
rect 29932 6616 30052 6644
rect 30024 6322 30052 6616
rect 30116 6322 30144 6718
rect 29828 6316 29880 6322
rect 29828 6258 29880 6264
rect 30012 6316 30064 6322
rect 30012 6258 30064 6264
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 29642 5808 29698 5817
rect 29460 5772 29512 5778
rect 29460 5714 29512 5720
rect 29552 5772 29604 5778
rect 29840 5778 29868 6258
rect 30024 6118 30052 6258
rect 30300 6254 30328 7346
rect 30392 7342 30420 8384
rect 30484 7954 30512 8842
rect 30576 8634 30604 8978
rect 30564 8628 30616 8634
rect 30564 8570 30616 8576
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30576 7449 30604 8570
rect 30668 7478 30696 10542
rect 30760 9625 30788 12718
rect 30944 11286 30972 14418
rect 31036 13870 31064 16730
rect 31114 16688 31170 16697
rect 31114 16623 31116 16632
rect 31168 16623 31170 16632
rect 31116 16594 31168 16600
rect 31300 16516 31352 16522
rect 31300 16458 31352 16464
rect 31208 16448 31260 16454
rect 31208 16390 31260 16396
rect 31116 16040 31168 16046
rect 31116 15982 31168 15988
rect 31128 14550 31156 15982
rect 31220 15638 31248 16390
rect 31208 15632 31260 15638
rect 31208 15574 31260 15580
rect 31312 15570 31340 16458
rect 31404 16046 31432 18022
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31300 15564 31352 15570
rect 31352 15524 31524 15552
rect 31300 15506 31352 15512
rect 31390 14920 31446 14929
rect 31390 14855 31446 14864
rect 31116 14544 31168 14550
rect 31116 14486 31168 14492
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 31036 11762 31064 13806
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30932 11280 30984 11286
rect 30932 11222 30984 11228
rect 31024 10600 31076 10606
rect 31024 10542 31076 10548
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30852 9994 30880 10066
rect 30840 9988 30892 9994
rect 30840 9930 30892 9936
rect 30746 9616 30802 9625
rect 30746 9551 30802 9560
rect 31036 9518 31064 10542
rect 31116 10532 31168 10538
rect 31116 10474 31168 10480
rect 31128 9926 31156 10474
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 31128 9518 31156 9862
rect 30748 9512 30800 9518
rect 31024 9512 31076 9518
rect 30800 9460 30972 9466
rect 30748 9454 30972 9460
rect 31024 9454 31076 9460
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 30760 9438 30972 9454
rect 30840 9376 30892 9382
rect 30840 9318 30892 9324
rect 30852 9110 30880 9318
rect 30840 9104 30892 9110
rect 30840 9046 30892 9052
rect 30944 9042 30972 9438
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30840 8424 30892 8430
rect 30840 8366 30892 8372
rect 30852 7546 30880 8366
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30656 7472 30708 7478
rect 30562 7440 30618 7449
rect 30656 7414 30708 7420
rect 30562 7375 30618 7384
rect 30380 7336 30432 7342
rect 30380 7278 30432 7284
rect 30668 6866 30696 7414
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30840 6860 30892 6866
rect 30840 6802 30892 6808
rect 30668 6390 30696 6802
rect 30656 6384 30708 6390
rect 30656 6326 30708 6332
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 29642 5743 29698 5752
rect 29828 5772 29880 5778
rect 29552 5714 29604 5720
rect 29828 5714 29880 5720
rect 29472 5166 29500 5714
rect 29564 5234 29592 5714
rect 29840 5370 29868 5714
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 30024 4690 30052 6054
rect 30300 5846 30328 6190
rect 30288 5840 30340 5846
rect 30288 5782 30340 5788
rect 30300 5098 30328 5782
rect 30852 5166 30880 6802
rect 30944 6361 30972 8978
rect 31036 8265 31064 9454
rect 31220 9110 31248 14350
rect 31300 9920 31352 9926
rect 31300 9862 31352 9868
rect 31312 9586 31340 9862
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 31300 9444 31352 9450
rect 31300 9386 31352 9392
rect 31208 9104 31260 9110
rect 31208 9046 31260 9052
rect 31312 8906 31340 9386
rect 31300 8900 31352 8906
rect 31300 8842 31352 8848
rect 31022 8256 31078 8265
rect 31022 8191 31078 8200
rect 31036 6866 31064 8191
rect 31024 6860 31076 6866
rect 31024 6802 31076 6808
rect 30930 6352 30986 6361
rect 30930 6287 30986 6296
rect 30840 5160 30892 5166
rect 30840 5102 30892 5108
rect 30288 5092 30340 5098
rect 30288 5034 30340 5040
rect 30012 4684 30064 4690
rect 30012 4626 30064 4632
rect 31404 3738 31432 14855
rect 31496 9042 31524 15524
rect 31588 14958 31616 20295
rect 31760 20052 31812 20058
rect 31760 19994 31812 20000
rect 31666 17504 31722 17513
rect 31666 17439 31722 17448
rect 31680 15502 31708 17439
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31772 15162 31800 19994
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 31576 14952 31628 14958
rect 31576 14894 31628 14900
rect 31576 12640 31628 12646
rect 31576 12582 31628 12588
rect 31484 9036 31536 9042
rect 31484 8978 31536 8984
rect 31588 8090 31616 12582
rect 31668 9988 31720 9994
rect 31668 9930 31720 9936
rect 31680 8362 31708 9930
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 31668 8356 31720 8362
rect 31668 8298 31720 8304
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31772 7954 31800 9454
rect 31760 7948 31812 7954
rect 31760 7890 31812 7896
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 28998 3088 29054 3097
rect 28998 3023 29054 3032
rect 27644 2748 27952 2757
rect 27644 2746 27650 2748
rect 27706 2746 27730 2748
rect 27786 2746 27810 2748
rect 27866 2746 27890 2748
rect 27946 2746 27952 2748
rect 27706 2694 27708 2746
rect 27888 2694 27890 2746
rect 27644 2692 27650 2694
rect 27706 2692 27730 2694
rect 27786 2692 27810 2694
rect 27866 2692 27890 2694
rect 27946 2692 27952 2694
rect 27644 2683 27952 2692
rect 26984 2204 27292 2213
rect 26984 2202 26990 2204
rect 27046 2202 27070 2204
rect 27126 2202 27150 2204
rect 27206 2202 27230 2204
rect 27286 2202 27292 2204
rect 27046 2150 27048 2202
rect 27228 2150 27230 2202
rect 26984 2148 26990 2150
rect 27046 2148 27070 2150
rect 27126 2148 27150 2150
rect 27206 2148 27230 2150
rect 27286 2148 27292 2150
rect 26984 2139 27292 2148
rect 26422 2000 26478 2009
rect 26422 1935 26478 1944
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 12096 1660 12404 1669
rect 12096 1658 12102 1660
rect 12158 1658 12182 1660
rect 12238 1658 12262 1660
rect 12318 1658 12342 1660
rect 12398 1658 12404 1660
rect 12158 1606 12160 1658
rect 12340 1606 12342 1658
rect 12096 1604 12102 1606
rect 12158 1604 12182 1606
rect 12238 1604 12262 1606
rect 12318 1604 12342 1606
rect 12398 1604 12404 1606
rect 12096 1595 12404 1604
rect 19870 1660 20178 1669
rect 19870 1658 19876 1660
rect 19932 1658 19956 1660
rect 20012 1658 20036 1660
rect 20092 1658 20116 1660
rect 20172 1658 20178 1660
rect 19932 1606 19934 1658
rect 20114 1606 20116 1658
rect 19870 1604 19876 1606
rect 19932 1604 19956 1606
rect 20012 1604 20036 1606
rect 20092 1604 20116 1606
rect 20172 1604 20178 1606
rect 19870 1595 20178 1604
rect 27644 1660 27952 1669
rect 27644 1658 27650 1660
rect 27706 1658 27730 1660
rect 27786 1658 27810 1660
rect 27866 1658 27890 1660
rect 27946 1658 27952 1660
rect 27706 1606 27708 1658
rect 27888 1606 27890 1658
rect 27644 1604 27650 1606
rect 27706 1604 27730 1606
rect 27786 1604 27810 1606
rect 27866 1604 27890 1606
rect 27946 1604 27952 1606
rect 27644 1595 27952 1604
rect 1122 1456 1178 1465
rect 1122 1391 1178 1400
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 11436 1116 11744 1125
rect 11436 1114 11442 1116
rect 11498 1114 11522 1116
rect 11578 1114 11602 1116
rect 11658 1114 11682 1116
rect 11738 1114 11744 1116
rect 11498 1062 11500 1114
rect 11680 1062 11682 1114
rect 11436 1060 11442 1062
rect 11498 1060 11522 1062
rect 11578 1060 11602 1062
rect 11658 1060 11682 1062
rect 11738 1060 11744 1062
rect 11436 1051 11744 1060
rect 19210 1116 19518 1125
rect 19210 1114 19216 1116
rect 19272 1114 19296 1116
rect 19352 1114 19376 1116
rect 19432 1114 19456 1116
rect 19512 1114 19518 1116
rect 19272 1062 19274 1114
rect 19454 1062 19456 1114
rect 19210 1060 19216 1062
rect 19272 1060 19296 1062
rect 19352 1060 19376 1062
rect 19432 1060 19456 1062
rect 19512 1060 19518 1062
rect 19210 1051 19518 1060
rect 26984 1116 27292 1125
rect 26984 1114 26990 1116
rect 27046 1114 27070 1116
rect 27126 1114 27150 1116
rect 27206 1114 27230 1116
rect 27286 1114 27292 1116
rect 27046 1062 27048 1114
rect 27228 1062 27230 1114
rect 26984 1060 26990 1062
rect 27046 1060 27070 1062
rect 27126 1060 27150 1062
rect 27206 1060 27230 1062
rect 27286 1060 27292 1062
rect 26984 1051 27292 1060
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 12096 572 12404 581
rect 12096 570 12102 572
rect 12158 570 12182 572
rect 12238 570 12262 572
rect 12318 570 12342 572
rect 12398 570 12404 572
rect 12158 518 12160 570
rect 12340 518 12342 570
rect 12096 516 12102 518
rect 12158 516 12182 518
rect 12238 516 12262 518
rect 12318 516 12342 518
rect 12398 516 12404 518
rect 12096 507 12404 516
rect 19870 572 20178 581
rect 19870 570 19876 572
rect 19932 570 19956 572
rect 20012 570 20036 572
rect 20092 570 20116 572
rect 20172 570 20178 572
rect 19932 518 19934 570
rect 20114 518 20116 570
rect 19870 516 19876 518
rect 19932 516 19956 518
rect 20012 516 20036 518
rect 20092 516 20116 518
rect 20172 516 20178 518
rect 19870 507 20178 516
rect 27644 572 27952 581
rect 27644 570 27650 572
rect 27706 570 27730 572
rect 27786 570 27810 572
rect 27866 570 27890 572
rect 27946 570 27952 572
rect 27706 518 27708 570
rect 27888 518 27890 570
rect 27644 516 27650 518
rect 27706 516 27730 518
rect 27786 516 27810 518
rect 27866 516 27890 518
rect 27946 516 27952 518
rect 27644 507 27952 516
<< via2 >>
rect 6550 22072 6606 22128
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 6182 21684 6238 21720
rect 6182 21664 6184 21684
rect 6184 21664 6236 21684
rect 6236 21664 6238 21684
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 754 20304 810 20360
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 2318 19896 2374 19952
rect 846 13232 902 13288
rect 754 7928 810 7984
rect 662 6840 718 6896
rect 846 6160 902 6216
rect 1122 11056 1178 11112
rect 1030 8336 1086 8392
rect 1582 15952 1638 16008
rect 1950 17584 2006 17640
rect 2226 17756 2228 17776
rect 2228 17756 2280 17776
rect 2280 17756 2282 17776
rect 2226 17720 2282 17756
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 3238 18692 3294 18728
rect 3238 18672 3240 18692
rect 3240 18672 3292 18692
rect 3292 18672 3294 18692
rect 1858 13912 1914 13968
rect 1674 12144 1730 12200
rect 1582 11872 1638 11928
rect 1674 11464 1730 11520
rect 2226 13776 2282 13832
rect 2134 12552 2190 12608
rect 2226 11600 2282 11656
rect 3330 17040 3386 17096
rect 3146 15272 3202 15328
rect 2410 11600 2466 11656
rect 2318 11464 2374 11520
rect 2226 7420 2228 7440
rect 2228 7420 2280 7440
rect 2280 7420 2282 7440
rect 2226 7384 2282 7420
rect 1858 5208 1914 5264
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 3514 17040 3570 17096
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 2962 11756 3018 11792
rect 2962 11736 2964 11756
rect 2964 11736 3016 11756
rect 3016 11736 3018 11756
rect 2502 9968 2558 10024
rect 2778 11328 2834 11384
rect 2962 11228 2964 11248
rect 2964 11228 3016 11248
rect 3016 11228 3018 11248
rect 2962 11192 3018 11228
rect 2686 9560 2742 9616
rect 2502 5636 2558 5672
rect 2502 5616 2504 5636
rect 2504 5616 2556 5636
rect 2556 5616 2558 5636
rect 4342 17312 4398 17368
rect 4802 17312 4858 17368
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 5906 18536 5962 18592
rect 4986 16652 5042 16688
rect 4986 16632 4988 16652
rect 4988 16632 5040 16652
rect 5040 16632 5042 16652
rect 4802 16496 4858 16552
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 3330 13232 3386 13288
rect 3054 9288 3110 9344
rect 2502 5072 2558 5128
rect 3238 10648 3294 10704
rect 3238 9560 3294 9616
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 3514 11328 3570 11384
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 4434 12824 4490 12880
rect 4802 13504 4858 13560
rect 5078 15136 5134 15192
rect 5078 14048 5134 14104
rect 5078 13776 5134 13832
rect 4710 12824 4766 12880
rect 4158 11464 4214 11520
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 3698 10548 3700 10568
rect 3700 10548 3752 10568
rect 3752 10548 3754 10568
rect 3698 10512 3754 10548
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 4802 12280 4858 12336
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 4618 11056 4674 11112
rect 4342 10784 4398 10840
rect 3790 10260 3846 10296
rect 3790 10240 3792 10260
rect 3792 10240 3844 10260
rect 3844 10240 3846 10260
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 3514 9016 3570 9072
rect 4066 8744 4122 8800
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 4710 10920 4766 10976
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 4250 10004 4252 10024
rect 4252 10004 4304 10024
rect 4304 10004 4306 10024
rect 4250 9968 4306 10004
rect 4342 9832 4398 9888
rect 4802 9288 4858 9344
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 4342 8628 4398 8664
rect 4342 8608 4344 8628
rect 4344 8608 4396 8628
rect 4396 8608 4398 8628
rect 3606 8372 3608 8392
rect 3608 8372 3660 8392
rect 3660 8372 3662 8392
rect 3606 8336 3662 8372
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 3974 7284 3976 7304
rect 3976 7284 4028 7304
rect 4028 7284 4030 7304
rect 3974 7248 4030 7284
rect 4526 8880 4582 8936
rect 4526 8744 4582 8800
rect 4618 8472 4674 8528
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 3974 6704 4030 6760
rect 4894 7812 4950 7848
rect 4894 7792 4896 7812
rect 4896 7792 4948 7812
rect 4948 7792 4950 7812
rect 4894 7540 4950 7576
rect 5078 12960 5134 13016
rect 6274 18808 6330 18864
rect 6182 18400 6238 18456
rect 6090 17992 6146 18048
rect 5538 15444 5540 15464
rect 5540 15444 5592 15464
rect 5592 15444 5594 15464
rect 5538 15408 5594 15444
rect 5814 17040 5870 17096
rect 5814 14864 5870 14920
rect 5538 14184 5594 14240
rect 5354 13096 5410 13152
rect 5170 11464 5226 11520
rect 5538 12824 5594 12880
rect 5078 8880 5134 8936
rect 5078 8200 5134 8256
rect 5630 12144 5686 12200
rect 11886 21936 11942 21992
rect 6734 21684 6790 21720
rect 6734 21664 6736 21684
rect 6736 21664 6788 21684
rect 6788 21664 6790 21684
rect 7286 21684 7342 21720
rect 7286 21664 7288 21684
rect 7288 21664 7340 21684
rect 7340 21664 7342 21684
rect 7838 21684 7894 21720
rect 7838 21664 7840 21684
rect 7840 21664 7892 21684
rect 7892 21664 7894 21684
rect 8390 21684 8446 21720
rect 8390 21664 8392 21684
rect 8392 21664 8444 21684
rect 8444 21664 8446 21684
rect 7562 20304 7618 20360
rect 7286 20032 7342 20088
rect 7010 18828 7066 18864
rect 7010 18808 7012 18828
rect 7012 18808 7064 18828
rect 7064 18808 7066 18828
rect 6642 18572 6644 18592
rect 6644 18572 6696 18592
rect 6696 18572 6698 18592
rect 6642 18536 6698 18572
rect 6734 17992 6790 18048
rect 6366 17040 6422 17096
rect 5722 10920 5778 10976
rect 5538 10412 5540 10432
rect 5540 10412 5592 10432
rect 5592 10412 5594 10432
rect 5538 10376 5594 10412
rect 5538 9696 5594 9752
rect 5446 9580 5502 9616
rect 5446 9560 5448 9580
rect 5448 9560 5500 9580
rect 5500 9560 5502 9580
rect 5078 7656 5134 7712
rect 4894 7520 4896 7540
rect 4896 7520 4948 7540
rect 4948 7520 4950 7540
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 4802 6296 4858 6352
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 3606 4120 3662 4176
rect 4250 5480 4306 5536
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 5354 7112 5410 7168
rect 5262 6024 5318 6080
rect 5998 12280 6054 12336
rect 6182 13776 6238 13832
rect 6182 13504 6238 13560
rect 6274 12688 6330 12744
rect 6182 12008 6238 12064
rect 5998 10376 6054 10432
rect 5998 8880 6054 8936
rect 5906 8200 5962 8256
rect 6366 12552 6422 12608
rect 6550 12724 6552 12744
rect 6552 12724 6604 12744
rect 6604 12724 6606 12744
rect 6550 12688 6606 12724
rect 6550 12552 6606 12608
rect 6274 10376 6330 10432
rect 6182 10240 6238 10296
rect 5998 7792 6054 7848
rect 5814 6296 5870 6352
rect 7562 19896 7618 19952
rect 8390 18828 8446 18864
rect 8390 18808 8392 18828
rect 8392 18808 8444 18828
rect 8444 18808 8446 18828
rect 8298 18536 8354 18592
rect 6918 17620 6920 17640
rect 6920 17620 6972 17640
rect 6972 17620 6974 17640
rect 6918 17584 6974 17620
rect 7102 17312 7158 17368
rect 6918 17176 6974 17232
rect 7562 17856 7618 17912
rect 7930 17856 7986 17912
rect 6918 14864 6974 14920
rect 6826 14592 6882 14648
rect 7010 14728 7066 14784
rect 7286 16088 7342 16144
rect 6734 12688 6790 12744
rect 6642 11056 6698 11112
rect 6274 8880 6330 8936
rect 6182 7112 6238 7168
rect 7286 15020 7342 15056
rect 7286 15000 7288 15020
rect 7288 15000 7340 15020
rect 7340 15000 7342 15020
rect 7654 16768 7710 16824
rect 7654 16224 7710 16280
rect 8390 18028 8392 18048
rect 8392 18028 8444 18048
rect 8444 18028 8446 18048
rect 8390 17992 8446 18028
rect 8206 17584 8262 17640
rect 8574 18128 8630 18184
rect 8482 17312 8538 17368
rect 8206 16668 8208 16688
rect 8208 16668 8260 16688
rect 8260 16668 8262 16688
rect 8206 16632 8262 16668
rect 7470 15272 7526 15328
rect 8298 15680 8354 15736
rect 8758 18128 8814 18184
rect 8850 17992 8906 18048
rect 8850 17856 8906 17912
rect 8942 16768 8998 16824
rect 8482 16224 8538 16280
rect 8022 15136 8078 15192
rect 7470 14864 7526 14920
rect 7470 14728 7526 14784
rect 7470 14220 7472 14240
rect 7472 14220 7524 14240
rect 7524 14220 7526 14240
rect 7470 14184 7526 14220
rect 7562 13776 7618 13832
rect 7194 12144 7250 12200
rect 7010 11192 7066 11248
rect 6642 9152 6698 9208
rect 6918 8336 6974 8392
rect 6918 7928 6974 7984
rect 6826 7384 6882 7440
rect 7562 13640 7618 13696
rect 7930 14592 7986 14648
rect 8022 14320 8078 14376
rect 8390 15544 8446 15600
rect 9586 21800 9642 21856
rect 9494 21684 9550 21720
rect 11442 21786 11498 21788
rect 11522 21786 11578 21788
rect 11602 21786 11658 21788
rect 11682 21786 11738 21788
rect 11442 21734 11488 21786
rect 11488 21734 11498 21786
rect 11522 21734 11552 21786
rect 11552 21734 11564 21786
rect 11564 21734 11578 21786
rect 11602 21734 11616 21786
rect 11616 21734 11628 21786
rect 11628 21734 11658 21786
rect 11682 21734 11692 21786
rect 11692 21734 11738 21786
rect 11442 21732 11498 21734
rect 11522 21732 11578 21734
rect 11602 21732 11658 21734
rect 11682 21732 11738 21734
rect 9494 21664 9496 21684
rect 9496 21664 9548 21684
rect 9548 21664 9550 21684
rect 10046 21684 10102 21720
rect 10046 21664 10048 21684
rect 10048 21664 10100 21684
rect 10100 21664 10102 21684
rect 10598 21684 10654 21720
rect 10598 21664 10600 21684
rect 10600 21664 10652 21684
rect 10652 21664 10654 21684
rect 11150 21684 11206 21720
rect 11150 21664 11152 21684
rect 11152 21664 11204 21684
rect 11204 21664 11206 21684
rect 10414 20848 10470 20904
rect 10138 19760 10194 19816
rect 9678 19352 9734 19408
rect 9218 18536 9274 18592
rect 9494 18400 9550 18456
rect 9218 17604 9274 17640
rect 9218 17584 9220 17604
rect 9220 17584 9272 17604
rect 9272 17584 9274 17604
rect 9310 17312 9366 17368
rect 8942 15816 8998 15872
rect 8942 15000 8998 15056
rect 8390 14456 8446 14512
rect 8574 14320 8630 14376
rect 8298 14184 8354 14240
rect 8758 14612 8814 14648
rect 8758 14592 8760 14612
rect 8760 14592 8812 14612
rect 8812 14592 8814 14612
rect 8758 14476 8814 14512
rect 8758 14456 8760 14476
rect 8760 14456 8812 14476
rect 8812 14456 8814 14476
rect 8206 13504 8262 13560
rect 8022 13132 8024 13152
rect 8024 13132 8076 13152
rect 8076 13132 8078 13152
rect 8022 13096 8078 13132
rect 7930 12552 7986 12608
rect 7930 12008 7986 12064
rect 7838 11464 7894 11520
rect 7562 9696 7618 9752
rect 7470 8880 7526 8936
rect 7102 6976 7158 7032
rect 6550 5888 6606 5944
rect 7746 10376 7802 10432
rect 7838 10240 7894 10296
rect 8022 11328 8078 11384
rect 8022 10920 8078 10976
rect 7930 9696 7986 9752
rect 7746 9288 7802 9344
rect 7746 9016 7802 9072
rect 7838 8628 7894 8664
rect 7838 8608 7840 8628
rect 7840 8608 7892 8628
rect 7892 8608 7894 8628
rect 7838 8472 7894 8528
rect 7654 7248 7710 7304
rect 7470 5480 7526 5536
rect 7654 5616 7710 5672
rect 7930 7112 7986 7168
rect 8390 13640 8446 13696
rect 8482 13096 8538 13152
rect 8758 13776 8814 13832
rect 8850 13388 8906 13424
rect 8850 13368 8852 13388
rect 8852 13368 8904 13388
rect 8904 13368 8906 13388
rect 8574 12688 8630 12744
rect 8206 10804 8262 10840
rect 8206 10784 8208 10804
rect 8208 10784 8260 10804
rect 8260 10784 8262 10804
rect 8298 10648 8354 10704
rect 8390 8472 8446 8528
rect 8298 8200 8354 8256
rect 8022 6024 8078 6080
rect 8298 6704 8354 6760
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 9218 13232 9274 13288
rect 9862 19216 9918 19272
rect 9494 15816 9550 15872
rect 9494 15544 9550 15600
rect 9402 13776 9458 13832
rect 9494 13368 9550 13424
rect 9586 13096 9642 13152
rect 9494 12824 9550 12880
rect 9126 12144 9182 12200
rect 8942 12008 8998 12064
rect 9310 12144 9366 12200
rect 9126 12008 9182 12064
rect 9402 12008 9458 12064
rect 8850 11464 8906 11520
rect 8850 10920 8906 10976
rect 9126 11056 9182 11112
rect 9310 10548 9312 10568
rect 9312 10548 9364 10568
rect 9364 10548 9366 10568
rect 9126 10240 9182 10296
rect 9310 10512 9366 10548
rect 9494 10920 9550 10976
rect 10230 17992 10286 18048
rect 10414 17312 10470 17368
rect 10230 16088 10286 16144
rect 9954 15272 10010 15328
rect 9862 13504 9918 13560
rect 10046 14048 10102 14104
rect 10046 13096 10102 13152
rect 10230 15272 10286 15328
rect 10230 15036 10232 15056
rect 10232 15036 10284 15056
rect 10284 15036 10286 15056
rect 10230 15000 10286 15036
rect 10230 14320 10286 14376
rect 10598 17992 10654 18048
rect 11150 20168 11206 20224
rect 11442 20698 11498 20700
rect 11522 20698 11578 20700
rect 11602 20698 11658 20700
rect 11682 20698 11738 20700
rect 11442 20646 11488 20698
rect 11488 20646 11498 20698
rect 11522 20646 11552 20698
rect 11552 20646 11564 20698
rect 11564 20646 11578 20698
rect 11602 20646 11616 20698
rect 11616 20646 11628 20698
rect 11628 20646 11658 20698
rect 11682 20646 11692 20698
rect 11692 20646 11738 20698
rect 11442 20644 11498 20646
rect 11522 20644 11578 20646
rect 11602 20644 11658 20646
rect 11682 20644 11738 20646
rect 12254 21936 12310 21992
rect 12806 21684 12862 21720
rect 12806 21664 12808 21684
rect 12808 21664 12860 21684
rect 12860 21664 12862 21684
rect 13358 21684 13414 21720
rect 13358 21664 13360 21684
rect 13360 21664 13412 21684
rect 13412 21664 13414 21684
rect 13910 21684 13966 21720
rect 13910 21664 13912 21684
rect 13912 21664 13964 21684
rect 13964 21664 13966 21684
rect 16670 21684 16726 21720
rect 16670 21664 16672 21684
rect 16672 21664 16724 21684
rect 16724 21664 16726 21684
rect 18418 21548 18474 21584
rect 18418 21528 18420 21548
rect 18420 21528 18472 21548
rect 18472 21528 18474 21548
rect 14370 21392 14426 21448
rect 12102 21242 12158 21244
rect 12182 21242 12238 21244
rect 12262 21242 12318 21244
rect 12342 21242 12398 21244
rect 12102 21190 12148 21242
rect 12148 21190 12158 21242
rect 12182 21190 12212 21242
rect 12212 21190 12224 21242
rect 12224 21190 12238 21242
rect 12262 21190 12276 21242
rect 12276 21190 12288 21242
rect 12288 21190 12318 21242
rect 12342 21190 12352 21242
rect 12352 21190 12398 21242
rect 12102 21188 12158 21190
rect 12182 21188 12238 21190
rect 12262 21188 12318 21190
rect 12342 21188 12398 21190
rect 11442 19610 11498 19612
rect 11522 19610 11578 19612
rect 11602 19610 11658 19612
rect 11682 19610 11738 19612
rect 11442 19558 11488 19610
rect 11488 19558 11498 19610
rect 11522 19558 11552 19610
rect 11552 19558 11564 19610
rect 11564 19558 11578 19610
rect 11602 19558 11616 19610
rect 11616 19558 11628 19610
rect 11628 19558 11658 19610
rect 11682 19558 11692 19610
rect 11692 19558 11738 19610
rect 11442 19556 11498 19558
rect 11522 19556 11578 19558
rect 11602 19556 11658 19558
rect 11682 19556 11738 19558
rect 12102 20154 12158 20156
rect 12182 20154 12238 20156
rect 12262 20154 12318 20156
rect 12342 20154 12398 20156
rect 12102 20102 12148 20154
rect 12148 20102 12158 20154
rect 12182 20102 12212 20154
rect 12212 20102 12224 20154
rect 12224 20102 12238 20154
rect 12262 20102 12276 20154
rect 12276 20102 12288 20154
rect 12288 20102 12318 20154
rect 12342 20102 12352 20154
rect 12352 20102 12398 20154
rect 12102 20100 12158 20102
rect 12182 20100 12238 20102
rect 12262 20100 12318 20102
rect 12342 20100 12398 20102
rect 11886 20032 11942 20088
rect 12714 20440 12770 20496
rect 12070 19352 12126 19408
rect 12806 20304 12862 20360
rect 12102 19066 12158 19068
rect 12182 19066 12238 19068
rect 12262 19066 12318 19068
rect 12342 19066 12398 19068
rect 12102 19014 12148 19066
rect 12148 19014 12158 19066
rect 12182 19014 12212 19066
rect 12212 19014 12224 19066
rect 12224 19014 12238 19066
rect 12262 19014 12276 19066
rect 12276 19014 12288 19066
rect 12288 19014 12318 19066
rect 12342 19014 12352 19066
rect 12352 19014 12398 19066
rect 12102 19012 12158 19014
rect 12182 19012 12238 19014
rect 12262 19012 12318 19014
rect 12342 19012 12398 19014
rect 11242 18264 11298 18320
rect 11242 17448 11298 17504
rect 11442 18522 11498 18524
rect 11522 18522 11578 18524
rect 11602 18522 11658 18524
rect 11682 18522 11738 18524
rect 11442 18470 11488 18522
rect 11488 18470 11498 18522
rect 11522 18470 11552 18522
rect 11552 18470 11564 18522
rect 11564 18470 11578 18522
rect 11602 18470 11616 18522
rect 11616 18470 11628 18522
rect 11628 18470 11658 18522
rect 11682 18470 11692 18522
rect 11692 18470 11738 18522
rect 11442 18468 11498 18470
rect 11522 18468 11578 18470
rect 11602 18468 11658 18470
rect 11682 18468 11738 18470
rect 11442 17434 11498 17436
rect 11522 17434 11578 17436
rect 11602 17434 11658 17436
rect 11682 17434 11738 17436
rect 11442 17382 11488 17434
rect 11488 17382 11498 17434
rect 11522 17382 11552 17434
rect 11552 17382 11564 17434
rect 11564 17382 11578 17434
rect 11602 17382 11616 17434
rect 11616 17382 11628 17434
rect 11628 17382 11658 17434
rect 11682 17382 11692 17434
rect 11692 17382 11738 17434
rect 11442 17380 11498 17382
rect 11522 17380 11578 17382
rect 11602 17380 11658 17382
rect 11682 17380 11738 17382
rect 12102 17978 12158 17980
rect 12182 17978 12238 17980
rect 12262 17978 12318 17980
rect 12342 17978 12398 17980
rect 12102 17926 12148 17978
rect 12148 17926 12158 17978
rect 12182 17926 12212 17978
rect 12212 17926 12224 17978
rect 12224 17926 12238 17978
rect 12262 17926 12276 17978
rect 12276 17926 12288 17978
rect 12288 17926 12318 17978
rect 12342 17926 12352 17978
rect 12352 17926 12398 17978
rect 12102 17924 12158 17926
rect 12182 17924 12238 17926
rect 12262 17924 12318 17926
rect 12342 17924 12398 17926
rect 12530 17856 12586 17912
rect 12622 17720 12678 17776
rect 12346 17448 12402 17504
rect 12530 17484 12532 17504
rect 12532 17484 12584 17504
rect 12584 17484 12586 17504
rect 12530 17448 12586 17484
rect 12438 17312 12494 17368
rect 10874 16768 10930 16824
rect 11150 16768 11206 16824
rect 10966 16224 11022 16280
rect 12530 17040 12586 17096
rect 12102 16890 12158 16892
rect 12182 16890 12238 16892
rect 12262 16890 12318 16892
rect 12342 16890 12398 16892
rect 12102 16838 12148 16890
rect 12148 16838 12158 16890
rect 12182 16838 12212 16890
rect 12212 16838 12224 16890
rect 12224 16838 12238 16890
rect 12262 16838 12276 16890
rect 12276 16838 12288 16890
rect 12288 16838 12318 16890
rect 12342 16838 12352 16890
rect 12352 16838 12398 16890
rect 12102 16836 12158 16838
rect 12182 16836 12238 16838
rect 12262 16836 12318 16838
rect 12342 16836 12398 16838
rect 11442 16346 11498 16348
rect 11522 16346 11578 16348
rect 11602 16346 11658 16348
rect 11682 16346 11738 16348
rect 11442 16294 11488 16346
rect 11488 16294 11498 16346
rect 11522 16294 11552 16346
rect 11552 16294 11564 16346
rect 11564 16294 11578 16346
rect 11602 16294 11616 16346
rect 11616 16294 11628 16346
rect 11628 16294 11658 16346
rect 11682 16294 11692 16346
rect 11692 16294 11738 16346
rect 11442 16292 11498 16294
rect 11522 16292 11578 16294
rect 11602 16292 11658 16294
rect 11682 16292 11738 16294
rect 10690 15136 10746 15192
rect 10782 15000 10838 15056
rect 10598 14728 10654 14784
rect 11150 15952 11206 16008
rect 11058 15136 11114 15192
rect 10966 14864 11022 14920
rect 10874 14728 10930 14784
rect 10506 14492 10508 14512
rect 10508 14492 10560 14512
rect 10560 14492 10562 14512
rect 10506 14456 10562 14492
rect 10690 14456 10746 14512
rect 10598 14184 10654 14240
rect 10598 14048 10654 14104
rect 10414 13504 10470 13560
rect 10230 12860 10232 12880
rect 10232 12860 10284 12880
rect 10284 12860 10286 12880
rect 10230 12824 10286 12860
rect 9770 11600 9826 11656
rect 9402 10240 9458 10296
rect 9770 10784 9826 10840
rect 9586 10240 9642 10296
rect 9126 9596 9128 9616
rect 9128 9596 9180 9616
rect 9180 9596 9182 9616
rect 9126 9560 9182 9596
rect 8758 8492 8814 8528
rect 8758 8472 8760 8492
rect 8760 8472 8812 8492
rect 8812 8472 8814 8492
rect 8850 7520 8906 7576
rect 8758 7384 8814 7440
rect 8666 7112 8722 7168
rect 9678 9832 9734 9888
rect 9126 8472 9182 8528
rect 9402 8200 9458 8256
rect 9586 8064 9642 8120
rect 9034 7656 9090 7712
rect 9034 7112 9090 7168
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 9586 7384 9642 7440
rect 9402 6160 9458 6216
rect 9494 6024 9550 6080
rect 9770 8744 9826 8800
rect 10138 12008 10194 12064
rect 10230 11192 10286 11248
rect 10138 10920 10194 10976
rect 10138 10648 10194 10704
rect 10138 9832 10194 9888
rect 10230 9288 10286 9344
rect 10046 9036 10102 9072
rect 10046 9016 10048 9036
rect 10048 9016 10100 9036
rect 10100 9016 10102 9036
rect 10138 8744 10194 8800
rect 9954 7520 10010 7576
rect 9862 5888 9918 5944
rect 9402 4120 9458 4176
rect 9678 4528 9734 4584
rect 10782 13640 10838 13696
rect 11702 15680 11758 15736
rect 11886 16396 11888 16416
rect 11888 16396 11940 16416
rect 11940 16396 11942 16416
rect 11886 16360 11942 16396
rect 12346 16224 12402 16280
rect 12162 16088 12218 16144
rect 12806 17176 12862 17232
rect 12714 16940 12716 16960
rect 12716 16940 12768 16960
rect 12768 16940 12770 16960
rect 12714 16904 12770 16940
rect 12714 16768 12770 16824
rect 13082 19080 13138 19136
rect 12990 17856 13046 17912
rect 12530 16224 12586 16280
rect 12102 15802 12158 15804
rect 12182 15802 12238 15804
rect 12262 15802 12318 15804
rect 12342 15802 12398 15804
rect 12102 15750 12148 15802
rect 12148 15750 12158 15802
rect 12182 15750 12212 15802
rect 12212 15750 12224 15802
rect 12224 15750 12238 15802
rect 12262 15750 12276 15802
rect 12276 15750 12288 15802
rect 12288 15750 12318 15802
rect 12342 15750 12352 15802
rect 12352 15750 12398 15802
rect 12102 15748 12158 15750
rect 12182 15748 12238 15750
rect 12262 15748 12318 15750
rect 12342 15748 12398 15750
rect 12530 15816 12586 15872
rect 12622 15680 12678 15736
rect 11442 15258 11498 15260
rect 11522 15258 11578 15260
rect 11602 15258 11658 15260
rect 11682 15258 11738 15260
rect 11442 15206 11488 15258
rect 11488 15206 11498 15258
rect 11522 15206 11552 15258
rect 11552 15206 11564 15258
rect 11564 15206 11578 15258
rect 11602 15206 11616 15258
rect 11616 15206 11628 15258
rect 11628 15206 11658 15258
rect 11682 15206 11692 15258
rect 11692 15206 11738 15258
rect 11442 15204 11498 15206
rect 11522 15204 11578 15206
rect 11602 15204 11658 15206
rect 11682 15204 11738 15206
rect 11886 15136 11942 15192
rect 11518 15000 11574 15056
rect 11426 14900 11428 14920
rect 11428 14900 11480 14920
rect 11480 14900 11482 14920
rect 11426 14864 11482 14900
rect 12070 15272 12126 15328
rect 12438 15136 12494 15192
rect 12102 14714 12158 14716
rect 12182 14714 12238 14716
rect 12262 14714 12318 14716
rect 12342 14714 12398 14716
rect 12102 14662 12148 14714
rect 12148 14662 12158 14714
rect 12182 14662 12212 14714
rect 12212 14662 12224 14714
rect 12224 14662 12238 14714
rect 12262 14662 12276 14714
rect 12276 14662 12288 14714
rect 12288 14662 12318 14714
rect 12342 14662 12352 14714
rect 12352 14662 12398 14714
rect 12102 14660 12158 14662
rect 12182 14660 12238 14662
rect 12262 14660 12318 14662
rect 12342 14660 12398 14662
rect 11058 14048 11114 14104
rect 10874 13096 10930 13152
rect 10966 12960 11022 13016
rect 11978 14184 12034 14240
rect 11442 14170 11498 14172
rect 11522 14170 11578 14172
rect 11602 14170 11658 14172
rect 11682 14170 11738 14172
rect 11442 14118 11488 14170
rect 11488 14118 11498 14170
rect 11522 14118 11552 14170
rect 11552 14118 11564 14170
rect 11564 14118 11578 14170
rect 11602 14118 11616 14170
rect 11616 14118 11628 14170
rect 11628 14118 11658 14170
rect 11682 14118 11692 14170
rect 11692 14118 11738 14170
rect 11442 14116 11498 14118
rect 11522 14116 11578 14118
rect 11602 14116 11658 14118
rect 11682 14116 11738 14118
rect 11242 14048 11298 14104
rect 11702 13504 11758 13560
rect 12622 15272 12678 15328
rect 12622 14184 12678 14240
rect 11150 13232 11206 13288
rect 11058 12552 11114 12608
rect 11150 12416 11206 12472
rect 10690 12008 10746 12064
rect 10506 10512 10562 10568
rect 10874 12008 10930 12064
rect 10966 11872 11022 11928
rect 10782 11192 10838 11248
rect 10598 10240 10654 10296
rect 10506 9696 10562 9752
rect 10322 9016 10378 9072
rect 10230 6568 10286 6624
rect 10046 4800 10102 4856
rect 10690 8064 10746 8120
rect 10690 6432 10746 6488
rect 10414 4564 10416 4584
rect 10416 4564 10468 4584
rect 10468 4564 10470 4584
rect 10414 4528 10470 4564
rect 9954 4120 10010 4176
rect 11442 13082 11498 13084
rect 11522 13082 11578 13084
rect 11602 13082 11658 13084
rect 11682 13082 11738 13084
rect 11442 13030 11488 13082
rect 11488 13030 11498 13082
rect 11522 13030 11552 13082
rect 11552 13030 11564 13082
rect 11564 13030 11578 13082
rect 11602 13030 11616 13082
rect 11616 13030 11628 13082
rect 11628 13030 11658 13082
rect 11682 13030 11692 13082
rect 11692 13030 11738 13082
rect 11442 13028 11498 13030
rect 11522 13028 11578 13030
rect 11602 13028 11658 13030
rect 11682 13028 11738 13030
rect 11334 12552 11390 12608
rect 12102 13626 12158 13628
rect 12182 13626 12238 13628
rect 12262 13626 12318 13628
rect 12342 13626 12398 13628
rect 12102 13574 12148 13626
rect 12148 13574 12158 13626
rect 12182 13574 12212 13626
rect 12212 13574 12224 13626
rect 12224 13574 12238 13626
rect 12262 13574 12276 13626
rect 12276 13574 12288 13626
rect 12288 13574 12318 13626
rect 12342 13574 12352 13626
rect 12352 13574 12398 13626
rect 12102 13572 12158 13574
rect 12182 13572 12238 13574
rect 12262 13572 12318 13574
rect 12342 13572 12398 13574
rect 12530 13524 12586 13560
rect 12530 13504 12532 13524
rect 12532 13504 12584 13524
rect 12584 13504 12586 13524
rect 11442 11994 11498 11996
rect 11522 11994 11578 11996
rect 11602 11994 11658 11996
rect 11682 11994 11738 11996
rect 11442 11942 11488 11994
rect 11488 11942 11498 11994
rect 11522 11942 11552 11994
rect 11552 11942 11564 11994
rect 11564 11942 11578 11994
rect 11602 11942 11616 11994
rect 11616 11942 11628 11994
rect 11628 11942 11658 11994
rect 11682 11942 11692 11994
rect 11692 11942 11738 11994
rect 11442 11940 11498 11942
rect 11522 11940 11578 11942
rect 11602 11940 11658 11942
rect 11682 11940 11738 11942
rect 11702 11736 11758 11792
rect 12254 12960 12310 13016
rect 12162 12824 12218 12880
rect 12990 15816 13046 15872
rect 12990 14592 13046 14648
rect 13082 14456 13138 14512
rect 12806 13640 12862 13696
rect 13266 19488 13322 19544
rect 13726 19488 13782 19544
rect 13726 19080 13782 19136
rect 13542 18808 13598 18864
rect 13358 15816 13414 15872
rect 13358 15544 13414 15600
rect 13266 14320 13322 14376
rect 13726 18672 13782 18728
rect 13634 18164 13636 18184
rect 13636 18164 13688 18184
rect 13688 18164 13690 18184
rect 13634 18128 13690 18164
rect 13818 17312 13874 17368
rect 13726 17176 13782 17232
rect 13542 16768 13598 16824
rect 13726 17040 13782 17096
rect 13818 16768 13874 16824
rect 13542 15952 13598 16008
rect 13818 16496 13874 16552
rect 13266 13640 13322 13696
rect 12102 12538 12158 12540
rect 12182 12538 12238 12540
rect 12262 12538 12318 12540
rect 12342 12538 12398 12540
rect 12102 12486 12148 12538
rect 12148 12486 12158 12538
rect 12182 12486 12212 12538
rect 12212 12486 12224 12538
rect 12224 12486 12238 12538
rect 12262 12486 12276 12538
rect 12276 12486 12288 12538
rect 12288 12486 12318 12538
rect 12342 12486 12352 12538
rect 12352 12486 12398 12538
rect 12102 12484 12158 12486
rect 12182 12484 12238 12486
rect 12262 12484 12318 12486
rect 12342 12484 12398 12486
rect 12070 12144 12126 12200
rect 10874 9696 10930 9752
rect 10874 9288 10930 9344
rect 10966 8744 11022 8800
rect 10966 8336 11022 8392
rect 11610 11056 11666 11112
rect 11442 10906 11498 10908
rect 11522 10906 11578 10908
rect 11602 10906 11658 10908
rect 11682 10906 11738 10908
rect 11442 10854 11488 10906
rect 11488 10854 11498 10906
rect 11522 10854 11552 10906
rect 11552 10854 11564 10906
rect 11564 10854 11578 10906
rect 11602 10854 11616 10906
rect 11616 10854 11628 10906
rect 11628 10854 11658 10906
rect 11682 10854 11692 10906
rect 11692 10854 11738 10906
rect 11442 10852 11498 10854
rect 11522 10852 11578 10854
rect 11602 10852 11658 10854
rect 11682 10852 11738 10854
rect 11242 10784 11298 10840
rect 12162 11736 12218 11792
rect 12102 11450 12158 11452
rect 12182 11450 12238 11452
rect 12262 11450 12318 11452
rect 12342 11450 12398 11452
rect 12102 11398 12148 11450
rect 12148 11398 12158 11450
rect 12182 11398 12212 11450
rect 12212 11398 12224 11450
rect 12224 11398 12238 11450
rect 12262 11398 12276 11450
rect 12276 11398 12288 11450
rect 12288 11398 12318 11450
rect 12342 11398 12352 11450
rect 12352 11398 12398 11450
rect 12102 11396 12158 11398
rect 12182 11396 12238 11398
rect 12262 11396 12318 11398
rect 12342 11396 12398 11398
rect 11886 11328 11942 11384
rect 11702 10412 11704 10432
rect 11704 10412 11756 10432
rect 11756 10412 11758 10432
rect 11702 10376 11758 10412
rect 11610 10240 11666 10296
rect 11442 9818 11498 9820
rect 11522 9818 11578 9820
rect 11602 9818 11658 9820
rect 11682 9818 11738 9820
rect 11442 9766 11488 9818
rect 11488 9766 11498 9818
rect 11522 9766 11552 9818
rect 11552 9766 11564 9818
rect 11564 9766 11578 9818
rect 11602 9766 11616 9818
rect 11616 9766 11628 9818
rect 11628 9766 11658 9818
rect 11682 9766 11692 9818
rect 11692 9766 11738 9818
rect 11442 9764 11498 9766
rect 11522 9764 11578 9766
rect 11602 9764 11658 9766
rect 11682 9764 11738 9766
rect 11518 9460 11520 9480
rect 11520 9460 11572 9480
rect 11572 9460 11574 9480
rect 11518 9424 11574 9460
rect 11518 9152 11574 9208
rect 11610 9036 11666 9072
rect 11610 9016 11612 9036
rect 11612 9016 11664 9036
rect 11664 9016 11666 9036
rect 11442 8730 11498 8732
rect 11522 8730 11578 8732
rect 11602 8730 11658 8732
rect 11682 8730 11738 8732
rect 11442 8678 11488 8730
rect 11488 8678 11498 8730
rect 11522 8678 11552 8730
rect 11552 8678 11564 8730
rect 11564 8678 11578 8730
rect 11602 8678 11616 8730
rect 11616 8678 11628 8730
rect 11628 8678 11658 8730
rect 11682 8678 11692 8730
rect 11692 8678 11738 8730
rect 11442 8676 11498 8678
rect 11522 8676 11578 8678
rect 11602 8676 11658 8678
rect 11682 8676 11738 8678
rect 12346 10648 12402 10704
rect 12162 10512 12218 10568
rect 12102 10362 12158 10364
rect 12182 10362 12238 10364
rect 12262 10362 12318 10364
rect 12342 10362 12398 10364
rect 12102 10310 12148 10362
rect 12148 10310 12158 10362
rect 12182 10310 12212 10362
rect 12212 10310 12224 10362
rect 12224 10310 12238 10362
rect 12262 10310 12276 10362
rect 12276 10310 12288 10362
rect 12288 10310 12318 10362
rect 12342 10310 12352 10362
rect 12352 10310 12398 10362
rect 12102 10308 12158 10310
rect 12182 10308 12238 10310
rect 12262 10308 12318 10310
rect 12342 10308 12398 10310
rect 12530 11872 12586 11928
rect 12898 12552 12954 12608
rect 12102 9274 12158 9276
rect 12182 9274 12238 9276
rect 12262 9274 12318 9276
rect 12342 9274 12398 9276
rect 12102 9222 12148 9274
rect 12148 9222 12158 9274
rect 12182 9222 12212 9274
rect 12212 9222 12224 9274
rect 12224 9222 12238 9274
rect 12262 9222 12276 9274
rect 12276 9222 12288 9274
rect 12288 9222 12318 9274
rect 12342 9222 12352 9274
rect 12352 9222 12398 9274
rect 12102 9220 12158 9222
rect 12182 9220 12238 9222
rect 12262 9220 12318 9222
rect 12342 9220 12398 9222
rect 11442 7642 11498 7644
rect 11522 7642 11578 7644
rect 11602 7642 11658 7644
rect 11682 7642 11738 7644
rect 11442 7590 11488 7642
rect 11488 7590 11498 7642
rect 11522 7590 11552 7642
rect 11552 7590 11564 7642
rect 11564 7590 11578 7642
rect 11602 7590 11616 7642
rect 11616 7590 11628 7642
rect 11628 7590 11658 7642
rect 11682 7590 11692 7642
rect 11692 7590 11738 7642
rect 11442 7588 11498 7590
rect 11522 7588 11578 7590
rect 11602 7588 11658 7590
rect 11682 7588 11738 7590
rect 12622 9288 12678 9344
rect 11978 8744 12034 8800
rect 12346 8472 12402 8528
rect 12806 11872 12862 11928
rect 12990 11328 13046 11384
rect 12898 11056 12954 11112
rect 12990 10240 13046 10296
rect 13818 14900 13820 14920
rect 13820 14900 13872 14920
rect 13872 14900 13874 14920
rect 13818 14864 13874 14900
rect 14462 20596 14518 20632
rect 14462 20576 14464 20596
rect 14464 20576 14516 20596
rect 14516 20576 14518 20596
rect 14002 17484 14004 17504
rect 14004 17484 14056 17504
rect 14056 17484 14058 17504
rect 14002 17448 14058 17484
rect 13634 14456 13690 14512
rect 13634 13912 13690 13968
rect 13174 12688 13230 12744
rect 13174 11600 13230 11656
rect 13634 12844 13690 12880
rect 13634 12824 13636 12844
rect 13636 12824 13688 12844
rect 13688 12824 13690 12844
rect 13542 12688 13598 12744
rect 13266 10376 13322 10432
rect 13174 9288 13230 9344
rect 13082 9152 13138 9208
rect 11886 8064 11942 8120
rect 12102 8186 12158 8188
rect 12182 8186 12238 8188
rect 12262 8186 12318 8188
rect 12342 8186 12398 8188
rect 12102 8134 12148 8186
rect 12148 8134 12158 8186
rect 12182 8134 12212 8186
rect 12212 8134 12224 8186
rect 12224 8134 12238 8186
rect 12262 8134 12276 8186
rect 12276 8134 12288 8186
rect 12288 8134 12318 8186
rect 12342 8134 12352 8186
rect 12352 8134 12398 8186
rect 12102 8132 12158 8134
rect 12182 8132 12238 8134
rect 12262 8132 12318 8134
rect 12342 8132 12398 8134
rect 11978 7656 12034 7712
rect 12438 7384 12494 7440
rect 11442 6554 11498 6556
rect 11522 6554 11578 6556
rect 11602 6554 11658 6556
rect 11682 6554 11738 6556
rect 11442 6502 11488 6554
rect 11488 6502 11498 6554
rect 11522 6502 11552 6554
rect 11552 6502 11564 6554
rect 11564 6502 11578 6554
rect 11602 6502 11616 6554
rect 11616 6502 11628 6554
rect 11628 6502 11658 6554
rect 11682 6502 11692 6554
rect 11692 6502 11738 6554
rect 11442 6500 11498 6502
rect 11522 6500 11578 6502
rect 11602 6500 11658 6502
rect 11682 6500 11738 6502
rect 12102 7098 12158 7100
rect 12182 7098 12238 7100
rect 12262 7098 12318 7100
rect 12342 7098 12398 7100
rect 12102 7046 12148 7098
rect 12148 7046 12158 7098
rect 12182 7046 12212 7098
rect 12212 7046 12224 7098
rect 12224 7046 12238 7098
rect 12262 7046 12276 7098
rect 12276 7046 12288 7098
rect 12288 7046 12318 7098
rect 12342 7046 12352 7098
rect 12352 7046 12398 7098
rect 12102 7044 12158 7046
rect 12182 7044 12238 7046
rect 12262 7044 12318 7046
rect 12342 7044 12398 7046
rect 12530 7148 12532 7168
rect 12532 7148 12584 7168
rect 12584 7148 12586 7168
rect 12530 7112 12586 7148
rect 12622 6976 12678 7032
rect 11978 6568 12034 6624
rect 11886 6432 11942 6488
rect 11058 6296 11114 6352
rect 10874 5752 10930 5808
rect 10874 5616 10930 5672
rect 10598 3576 10654 3632
rect 8850 2488 8906 2544
rect 11334 5888 11390 5944
rect 11794 6060 11796 6080
rect 11796 6060 11848 6080
rect 11848 6060 11850 6080
rect 11794 6024 11850 6060
rect 12254 6296 12310 6352
rect 12438 6740 12440 6760
rect 12440 6740 12492 6760
rect 12492 6740 12494 6760
rect 12438 6704 12494 6740
rect 12102 6010 12158 6012
rect 12182 6010 12238 6012
rect 12262 6010 12318 6012
rect 12342 6010 12398 6012
rect 12102 5958 12148 6010
rect 12148 5958 12158 6010
rect 12182 5958 12212 6010
rect 12212 5958 12224 6010
rect 12224 5958 12238 6010
rect 12262 5958 12276 6010
rect 12276 5958 12288 6010
rect 12288 5958 12318 6010
rect 12342 5958 12352 6010
rect 12352 5958 12398 6010
rect 12102 5956 12158 5958
rect 12182 5956 12238 5958
rect 12262 5956 12318 5958
rect 12342 5956 12398 5958
rect 11442 5466 11498 5468
rect 11522 5466 11578 5468
rect 11602 5466 11658 5468
rect 11682 5466 11738 5468
rect 11442 5414 11488 5466
rect 11488 5414 11498 5466
rect 11522 5414 11552 5466
rect 11552 5414 11564 5466
rect 11564 5414 11578 5466
rect 11602 5414 11616 5466
rect 11616 5414 11628 5466
rect 11628 5414 11658 5466
rect 11682 5414 11692 5466
rect 11692 5414 11738 5466
rect 11442 5412 11498 5414
rect 11522 5412 11578 5414
rect 11602 5412 11658 5414
rect 11682 5412 11738 5414
rect 13358 8472 13414 8528
rect 12990 6704 13046 6760
rect 12714 5480 12770 5536
rect 12102 4922 12158 4924
rect 12182 4922 12238 4924
rect 12262 4922 12318 4924
rect 12342 4922 12398 4924
rect 12102 4870 12148 4922
rect 12148 4870 12158 4922
rect 12182 4870 12212 4922
rect 12212 4870 12224 4922
rect 12224 4870 12238 4922
rect 12262 4870 12276 4922
rect 12276 4870 12288 4922
rect 12288 4870 12318 4922
rect 12342 4870 12352 4922
rect 12352 4870 12398 4922
rect 12102 4868 12158 4870
rect 12182 4868 12238 4870
rect 12262 4868 12318 4870
rect 12342 4868 12398 4870
rect 11978 4664 12034 4720
rect 11442 4378 11498 4380
rect 11522 4378 11578 4380
rect 11602 4378 11658 4380
rect 11682 4378 11738 4380
rect 11442 4326 11488 4378
rect 11488 4326 11498 4378
rect 11522 4326 11552 4378
rect 11552 4326 11564 4378
rect 11564 4326 11578 4378
rect 11602 4326 11616 4378
rect 11616 4326 11628 4378
rect 11628 4326 11658 4378
rect 11682 4326 11692 4378
rect 11692 4326 11738 4378
rect 11442 4324 11498 4326
rect 11522 4324 11578 4326
rect 11602 4324 11658 4326
rect 11682 4324 11738 4326
rect 11610 3984 11666 4040
rect 11442 3290 11498 3292
rect 11522 3290 11578 3292
rect 11602 3290 11658 3292
rect 11682 3290 11738 3292
rect 11442 3238 11488 3290
rect 11488 3238 11498 3290
rect 11522 3238 11552 3290
rect 11552 3238 11564 3290
rect 11564 3238 11578 3290
rect 11602 3238 11616 3290
rect 11616 3238 11628 3290
rect 11628 3238 11658 3290
rect 11682 3238 11692 3290
rect 11692 3238 11738 3290
rect 11442 3236 11498 3238
rect 11522 3236 11578 3238
rect 11602 3236 11658 3238
rect 11682 3236 11738 3238
rect 11978 4392 12034 4448
rect 12714 5108 12716 5128
rect 12716 5108 12768 5128
rect 12768 5108 12770 5128
rect 12714 5072 12770 5108
rect 12102 3834 12158 3836
rect 12182 3834 12238 3836
rect 12262 3834 12318 3836
rect 12342 3834 12398 3836
rect 12102 3782 12148 3834
rect 12148 3782 12158 3834
rect 12182 3782 12212 3834
rect 12212 3782 12224 3834
rect 12224 3782 12238 3834
rect 12262 3782 12276 3834
rect 12276 3782 12288 3834
rect 12288 3782 12318 3834
rect 12342 3782 12352 3834
rect 12352 3782 12398 3834
rect 12102 3780 12158 3782
rect 12182 3780 12238 3782
rect 12262 3780 12318 3782
rect 12342 3780 12398 3782
rect 12622 4528 12678 4584
rect 12990 5752 13046 5808
rect 13450 8064 13506 8120
rect 13634 12144 13690 12200
rect 13910 11056 13966 11112
rect 14370 19216 14426 19272
rect 14278 17584 14334 17640
rect 14554 18400 14610 18456
rect 15474 20984 15530 21040
rect 15198 20576 15254 20632
rect 14830 20440 14886 20496
rect 14738 18400 14794 18456
rect 14554 16768 14610 16824
rect 14278 16088 14334 16144
rect 14186 15816 14242 15872
rect 14094 15272 14150 15328
rect 15014 19916 15070 19952
rect 15014 19896 15016 19916
rect 15016 19896 15068 19916
rect 15068 19896 15070 19916
rect 15382 19896 15438 19952
rect 16486 21120 16542 21176
rect 15750 19488 15806 19544
rect 15106 18944 15162 19000
rect 14830 17720 14886 17776
rect 14646 15136 14702 15192
rect 14094 12688 14150 12744
rect 13634 9424 13690 9480
rect 13726 9016 13782 9072
rect 14002 9016 14058 9072
rect 13910 8880 13966 8936
rect 13542 7384 13598 7440
rect 14186 12180 14188 12200
rect 14188 12180 14240 12200
rect 14240 12180 14242 12200
rect 14186 12144 14242 12180
rect 14278 11464 14334 11520
rect 14186 10648 14242 10704
rect 14370 11212 14426 11248
rect 14370 11192 14372 11212
rect 14372 11192 14424 11212
rect 14424 11192 14426 11212
rect 14278 9832 14334 9888
rect 14462 10648 14518 10704
rect 14462 10376 14518 10432
rect 15014 16632 15070 16688
rect 14830 15952 14886 16008
rect 15106 15272 15162 15328
rect 14830 14320 14886 14376
rect 14830 14048 14886 14104
rect 15106 14320 15162 14376
rect 15290 14320 15346 14376
rect 14738 13504 14794 13560
rect 15014 14048 15070 14104
rect 14830 12552 14886 12608
rect 14738 12300 14794 12336
rect 14738 12280 14740 12300
rect 14740 12280 14792 12300
rect 14792 12280 14794 12300
rect 14738 11192 14794 11248
rect 15106 13948 15108 13968
rect 15108 13948 15160 13968
rect 15160 13948 15162 13968
rect 15106 13912 15162 13948
rect 15290 13640 15346 13696
rect 15290 12280 15346 12336
rect 15106 11736 15162 11792
rect 14922 11228 14924 11248
rect 14924 11228 14976 11248
rect 14976 11228 14978 11248
rect 14922 11192 14978 11228
rect 15106 11192 15162 11248
rect 17958 20596 18014 20632
rect 17958 20576 17960 20596
rect 17960 20576 18012 20596
rect 18012 20576 18014 20596
rect 17958 20168 18014 20224
rect 16854 19488 16910 19544
rect 15842 17620 15844 17640
rect 15844 17620 15896 17640
rect 15896 17620 15898 17640
rect 15842 17584 15898 17620
rect 15658 15680 15714 15736
rect 16026 16668 16028 16688
rect 16028 16668 16080 16688
rect 16080 16668 16082 16688
rect 16026 16632 16082 16668
rect 15934 16496 15990 16552
rect 15198 10920 15254 10976
rect 15014 10648 15070 10704
rect 15198 10668 15254 10704
rect 15198 10648 15200 10668
rect 15200 10648 15252 10668
rect 15252 10648 15254 10668
rect 14186 8880 14242 8936
rect 14186 8336 14242 8392
rect 14738 10140 14740 10160
rect 14740 10140 14792 10160
rect 14792 10140 14794 10160
rect 14738 10104 14794 10140
rect 13818 7656 13874 7712
rect 14094 7692 14096 7712
rect 14096 7692 14148 7712
rect 14148 7692 14150 7712
rect 14094 7656 14150 7692
rect 13910 7112 13966 7168
rect 13542 6840 13598 6896
rect 14462 8064 14518 8120
rect 14738 7948 14794 7984
rect 14738 7928 14740 7948
rect 14740 7928 14792 7948
rect 14792 7928 14794 7948
rect 15014 8608 15070 8664
rect 15014 8356 15070 8392
rect 15014 8336 15016 8356
rect 15016 8336 15068 8356
rect 15068 8336 15070 8356
rect 15014 8200 15070 8256
rect 14922 7656 14978 7712
rect 14462 5888 14518 5944
rect 13450 3848 13506 3904
rect 12898 3712 12954 3768
rect 13818 3576 13874 3632
rect 14278 3712 14334 3768
rect 14002 3576 14058 3632
rect 14738 6024 14794 6080
rect 15106 7656 15162 7712
rect 15106 6740 15108 6760
rect 15108 6740 15160 6760
rect 15160 6740 15162 6760
rect 15106 6704 15162 6740
rect 15382 9152 15438 9208
rect 15382 8628 15438 8664
rect 15382 8608 15384 8628
rect 15384 8608 15436 8628
rect 15436 8608 15438 8628
rect 15842 15408 15898 15464
rect 15842 13504 15898 13560
rect 15658 12724 15660 12744
rect 15660 12724 15712 12744
rect 15712 12724 15714 12744
rect 15658 12688 15714 12724
rect 15750 11736 15806 11792
rect 15566 10784 15622 10840
rect 15566 9288 15622 9344
rect 15566 8608 15622 8664
rect 15934 11872 15990 11928
rect 16394 16652 16450 16688
rect 16394 16632 16396 16652
rect 16396 16632 16448 16652
rect 16448 16632 16450 16652
rect 16394 15952 16450 16008
rect 17130 17448 17186 17504
rect 17038 17040 17094 17096
rect 16670 16224 16726 16280
rect 16670 15544 16726 15600
rect 16762 15444 16764 15464
rect 16764 15444 16816 15464
rect 16816 15444 16818 15464
rect 16762 15408 16818 15444
rect 16946 15136 17002 15192
rect 16946 14864 17002 14920
rect 16302 13776 16358 13832
rect 16210 13388 16266 13424
rect 16210 13368 16212 13388
rect 16212 13368 16264 13388
rect 16264 13368 16266 13388
rect 16118 12688 16174 12744
rect 16118 12008 16174 12064
rect 15750 10376 15806 10432
rect 16026 9832 16082 9888
rect 16026 9424 16082 9480
rect 15934 9288 15990 9344
rect 15566 8200 15622 8256
rect 15474 6996 15530 7032
rect 15474 6976 15476 6996
rect 15476 6976 15528 6996
rect 15528 6976 15530 6996
rect 14922 5344 14978 5400
rect 15106 5344 15162 5400
rect 15842 7656 15898 7712
rect 14370 3596 14426 3632
rect 14370 3576 14372 3596
rect 14372 3576 14424 3596
rect 14424 3576 14426 3596
rect 14922 5072 14978 5128
rect 16026 7656 16082 7712
rect 16118 6876 16120 6896
rect 16120 6876 16172 6896
rect 16172 6876 16174 6896
rect 16118 6840 16174 6876
rect 16026 5208 16082 5264
rect 15750 4800 15806 4856
rect 16486 13640 16542 13696
rect 16946 14048 17002 14104
rect 17498 16652 17554 16688
rect 17498 16632 17500 16652
rect 17500 16632 17552 16652
rect 17552 16632 17554 16652
rect 17498 16360 17554 16416
rect 18326 18536 18382 18592
rect 18050 16940 18052 16960
rect 18052 16940 18104 16960
rect 18104 16940 18106 16960
rect 18050 16904 18106 16940
rect 17958 15816 18014 15872
rect 18326 16768 18382 16824
rect 18050 14728 18106 14784
rect 17406 14184 17462 14240
rect 16854 13776 16910 13832
rect 16854 13368 16910 13424
rect 17038 13252 17094 13288
rect 17038 13232 17040 13252
rect 17040 13232 17092 13252
rect 17092 13232 17094 13252
rect 16302 9832 16358 9888
rect 16578 11328 16634 11384
rect 17038 12552 17094 12608
rect 16762 10784 16818 10840
rect 16762 10104 16818 10160
rect 16854 9832 16910 9888
rect 17038 12144 17094 12200
rect 17774 14048 17830 14104
rect 17590 13232 17646 13288
rect 17222 12008 17278 12064
rect 16578 9560 16634 9616
rect 16394 9460 16396 9480
rect 16396 9460 16448 9480
rect 16448 9460 16450 9480
rect 16394 9424 16450 9460
rect 16486 8356 16542 8392
rect 16486 8336 16488 8356
rect 16488 8336 16540 8356
rect 16540 8336 16542 8356
rect 16394 8064 16450 8120
rect 16670 8472 16726 8528
rect 16670 8064 16726 8120
rect 16486 7112 16542 7168
rect 16486 5772 16542 5808
rect 16486 5752 16488 5772
rect 16488 5752 16540 5772
rect 16540 5752 16542 5772
rect 16946 6976 17002 7032
rect 17590 12824 17646 12880
rect 17590 12300 17646 12336
rect 17590 12280 17592 12300
rect 17592 12280 17644 12300
rect 17644 12280 17646 12300
rect 17498 11056 17554 11112
rect 17774 13096 17830 13152
rect 17958 12960 18014 13016
rect 18234 13776 18290 13832
rect 17774 10240 17830 10296
rect 17498 9288 17554 9344
rect 17406 9152 17462 9208
rect 17222 8064 17278 8120
rect 17774 9832 17830 9888
rect 17774 9444 17830 9480
rect 17774 9424 17776 9444
rect 17776 9424 17828 9444
rect 17828 9424 17830 9444
rect 18418 14592 18474 14648
rect 18234 10920 18290 10976
rect 19216 21786 19272 21788
rect 19296 21786 19352 21788
rect 19376 21786 19432 21788
rect 19456 21786 19512 21788
rect 19216 21734 19262 21786
rect 19262 21734 19272 21786
rect 19296 21734 19326 21786
rect 19326 21734 19338 21786
rect 19338 21734 19352 21786
rect 19376 21734 19390 21786
rect 19390 21734 19402 21786
rect 19402 21734 19432 21786
rect 19456 21734 19466 21786
rect 19466 21734 19512 21786
rect 19216 21732 19272 21734
rect 19296 21732 19352 21734
rect 19376 21732 19432 21734
rect 19456 21732 19512 21734
rect 19062 21020 19064 21040
rect 19064 21020 19116 21040
rect 19116 21020 19118 21040
rect 19062 20984 19118 21020
rect 19876 21242 19932 21244
rect 19956 21242 20012 21244
rect 20036 21242 20092 21244
rect 20116 21242 20172 21244
rect 19876 21190 19922 21242
rect 19922 21190 19932 21242
rect 19956 21190 19986 21242
rect 19986 21190 19998 21242
rect 19998 21190 20012 21242
rect 20036 21190 20050 21242
rect 20050 21190 20062 21242
rect 20062 21190 20092 21242
rect 20116 21190 20126 21242
rect 20126 21190 20172 21242
rect 19876 21188 19932 21190
rect 19956 21188 20012 21190
rect 20036 21188 20092 21190
rect 20116 21188 20172 21190
rect 19216 20698 19272 20700
rect 19296 20698 19352 20700
rect 19376 20698 19432 20700
rect 19456 20698 19512 20700
rect 19216 20646 19262 20698
rect 19262 20646 19272 20698
rect 19296 20646 19326 20698
rect 19326 20646 19338 20698
rect 19338 20646 19352 20698
rect 19376 20646 19390 20698
rect 19390 20646 19402 20698
rect 19402 20646 19432 20698
rect 19456 20646 19466 20698
rect 19466 20646 19512 20698
rect 19216 20644 19272 20646
rect 19296 20644 19352 20646
rect 19376 20644 19432 20646
rect 19456 20644 19512 20646
rect 18786 18400 18842 18456
rect 18602 18264 18658 18320
rect 19154 19896 19210 19952
rect 19876 20154 19932 20156
rect 19956 20154 20012 20156
rect 20036 20154 20092 20156
rect 20116 20154 20172 20156
rect 19876 20102 19922 20154
rect 19922 20102 19932 20154
rect 19956 20102 19986 20154
rect 19986 20102 19998 20154
rect 19998 20102 20012 20154
rect 20036 20102 20050 20154
rect 20050 20102 20062 20154
rect 20062 20102 20092 20154
rect 20116 20102 20126 20154
rect 20126 20102 20172 20154
rect 19876 20100 19932 20102
rect 19956 20100 20012 20102
rect 20036 20100 20092 20102
rect 20116 20100 20172 20102
rect 20902 21292 20904 21312
rect 20904 21292 20956 21312
rect 20956 21292 20958 21312
rect 20902 21256 20958 21292
rect 20442 20168 20498 20224
rect 20350 20032 20406 20088
rect 19614 19624 19670 19680
rect 19216 19610 19272 19612
rect 19296 19610 19352 19612
rect 19376 19610 19432 19612
rect 19456 19610 19512 19612
rect 19216 19558 19262 19610
rect 19262 19558 19272 19610
rect 19296 19558 19326 19610
rect 19326 19558 19338 19610
rect 19338 19558 19352 19610
rect 19376 19558 19390 19610
rect 19390 19558 19402 19610
rect 19402 19558 19432 19610
rect 19456 19558 19466 19610
rect 19466 19558 19512 19610
rect 19216 19556 19272 19558
rect 19296 19556 19352 19558
rect 19376 19556 19432 19558
rect 19456 19556 19512 19558
rect 19216 18522 19272 18524
rect 19296 18522 19352 18524
rect 19376 18522 19432 18524
rect 19456 18522 19512 18524
rect 19216 18470 19262 18522
rect 19262 18470 19272 18522
rect 19296 18470 19326 18522
rect 19326 18470 19338 18522
rect 19338 18470 19352 18522
rect 19376 18470 19390 18522
rect 19390 18470 19402 18522
rect 19402 18470 19432 18522
rect 19456 18470 19466 18522
rect 19466 18470 19512 18522
rect 19216 18468 19272 18470
rect 19296 18468 19352 18470
rect 19376 18468 19432 18470
rect 19456 18468 19512 18470
rect 18602 17740 18658 17776
rect 18602 17720 18604 17740
rect 18604 17720 18656 17740
rect 18656 17720 18658 17740
rect 18602 15972 18658 16008
rect 18602 15952 18604 15972
rect 18604 15952 18656 15972
rect 18656 15952 18658 15972
rect 18602 14320 18658 14376
rect 18878 15408 18934 15464
rect 18970 14592 19026 14648
rect 19890 19352 19946 19408
rect 19876 19066 19932 19068
rect 19956 19066 20012 19068
rect 20036 19066 20092 19068
rect 20116 19066 20172 19068
rect 19876 19014 19922 19066
rect 19922 19014 19932 19066
rect 19956 19014 19986 19066
rect 19986 19014 19998 19066
rect 19998 19014 20012 19066
rect 20036 19014 20050 19066
rect 20050 19014 20062 19066
rect 20062 19014 20092 19066
rect 20116 19014 20126 19066
rect 20126 19014 20172 19066
rect 19876 19012 19932 19014
rect 19956 19012 20012 19014
rect 20036 19012 20092 19014
rect 20116 19012 20172 19014
rect 19890 18536 19946 18592
rect 20074 18264 20130 18320
rect 19706 17856 19762 17912
rect 19216 17434 19272 17436
rect 19296 17434 19352 17436
rect 19376 17434 19432 17436
rect 19456 17434 19512 17436
rect 19216 17382 19262 17434
rect 19262 17382 19272 17434
rect 19296 17382 19326 17434
rect 19326 17382 19338 17434
rect 19338 17382 19352 17434
rect 19376 17382 19390 17434
rect 19390 17382 19402 17434
rect 19402 17382 19432 17434
rect 19456 17382 19466 17434
rect 19466 17382 19512 17434
rect 19216 17380 19272 17382
rect 19296 17380 19352 17382
rect 19376 17380 19432 17382
rect 19456 17380 19512 17382
rect 19876 17978 19932 17980
rect 19956 17978 20012 17980
rect 20036 17978 20092 17980
rect 20116 17978 20172 17980
rect 19876 17926 19922 17978
rect 19922 17926 19932 17978
rect 19956 17926 19986 17978
rect 19986 17926 19998 17978
rect 19998 17926 20012 17978
rect 20036 17926 20050 17978
rect 20050 17926 20062 17978
rect 20062 17926 20092 17978
rect 20116 17926 20126 17978
rect 20126 17926 20172 17978
rect 19876 17924 19932 17926
rect 19956 17924 20012 17926
rect 20036 17924 20092 17926
rect 20116 17924 20172 17926
rect 20258 17856 20314 17912
rect 20810 18944 20866 19000
rect 20902 18808 20958 18864
rect 21270 21392 21326 21448
rect 21362 19236 21418 19272
rect 21362 19216 21364 19236
rect 21364 19216 21416 19236
rect 21416 19216 21418 19236
rect 21454 19080 21510 19136
rect 22282 20304 22338 20360
rect 21638 18944 21694 19000
rect 21546 18808 21602 18864
rect 20718 17856 20774 17912
rect 19982 17076 19984 17096
rect 19984 17076 20036 17096
rect 20036 17076 20038 17096
rect 19982 17040 20038 17076
rect 19876 16890 19932 16892
rect 19956 16890 20012 16892
rect 20036 16890 20092 16892
rect 20116 16890 20172 16892
rect 19876 16838 19922 16890
rect 19922 16838 19932 16890
rect 19956 16838 19986 16890
rect 19986 16838 19998 16890
rect 19998 16838 20012 16890
rect 20036 16838 20050 16890
rect 20050 16838 20062 16890
rect 20062 16838 20092 16890
rect 20116 16838 20126 16890
rect 20126 16838 20172 16890
rect 19876 16836 19932 16838
rect 19956 16836 20012 16838
rect 20036 16836 20092 16838
rect 20116 16836 20172 16838
rect 19216 16346 19272 16348
rect 19296 16346 19352 16348
rect 19376 16346 19432 16348
rect 19456 16346 19512 16348
rect 19216 16294 19262 16346
rect 19262 16294 19272 16346
rect 19296 16294 19326 16346
rect 19326 16294 19338 16346
rect 19338 16294 19352 16346
rect 19376 16294 19390 16346
rect 19390 16294 19402 16346
rect 19402 16294 19432 16346
rect 19456 16294 19466 16346
rect 19466 16294 19512 16346
rect 19216 16292 19272 16294
rect 19296 16292 19352 16294
rect 19376 16292 19432 16294
rect 19456 16292 19512 16294
rect 19706 16360 19762 16416
rect 19706 16224 19762 16280
rect 19982 16244 20038 16280
rect 20626 17040 20682 17096
rect 19982 16224 19984 16244
rect 19984 16224 20036 16244
rect 20036 16224 20038 16244
rect 19706 15444 19708 15464
rect 19708 15444 19760 15464
rect 19760 15444 19762 15464
rect 19706 15408 19762 15444
rect 19614 15272 19670 15328
rect 19216 15258 19272 15260
rect 19296 15258 19352 15260
rect 19376 15258 19432 15260
rect 19456 15258 19512 15260
rect 19216 15206 19262 15258
rect 19262 15206 19272 15258
rect 19296 15206 19326 15258
rect 19326 15206 19338 15258
rect 19338 15206 19352 15258
rect 19376 15206 19390 15258
rect 19390 15206 19402 15258
rect 19402 15206 19432 15258
rect 19456 15206 19466 15258
rect 19466 15206 19512 15258
rect 19216 15204 19272 15206
rect 19296 15204 19352 15206
rect 19376 15204 19432 15206
rect 19456 15204 19512 15206
rect 19338 15020 19394 15056
rect 19338 15000 19340 15020
rect 19340 15000 19392 15020
rect 19392 15000 19394 15020
rect 19338 14592 19394 14648
rect 19876 15802 19932 15804
rect 19956 15802 20012 15804
rect 20036 15802 20092 15804
rect 20116 15802 20172 15804
rect 19876 15750 19922 15802
rect 19922 15750 19932 15802
rect 19956 15750 19986 15802
rect 19986 15750 19998 15802
rect 19998 15750 20012 15802
rect 20036 15750 20050 15802
rect 20050 15750 20062 15802
rect 20062 15750 20092 15802
rect 20116 15750 20126 15802
rect 20126 15750 20172 15802
rect 19876 15748 19932 15750
rect 19956 15748 20012 15750
rect 20036 15748 20092 15750
rect 20116 15748 20172 15750
rect 19154 14340 19210 14376
rect 19154 14320 19156 14340
rect 19156 14320 19208 14340
rect 19208 14320 19210 14340
rect 19338 14356 19340 14376
rect 19340 14356 19392 14376
rect 19392 14356 19394 14376
rect 19338 14320 19394 14356
rect 19706 14612 19762 14648
rect 19706 14592 19708 14612
rect 19708 14592 19760 14612
rect 19760 14592 19762 14612
rect 19216 14170 19272 14172
rect 19296 14170 19352 14172
rect 19376 14170 19432 14172
rect 19456 14170 19512 14172
rect 19216 14118 19262 14170
rect 19262 14118 19272 14170
rect 19296 14118 19326 14170
rect 19326 14118 19338 14170
rect 19338 14118 19352 14170
rect 19376 14118 19390 14170
rect 19390 14118 19402 14170
rect 19402 14118 19432 14170
rect 19456 14118 19466 14170
rect 19466 14118 19512 14170
rect 19216 14116 19272 14118
rect 19296 14116 19352 14118
rect 19376 14116 19432 14118
rect 19456 14116 19512 14118
rect 18970 13640 19026 13696
rect 19154 13676 19156 13696
rect 19156 13676 19208 13696
rect 19208 13676 19210 13696
rect 19154 13640 19210 13676
rect 18878 13232 18934 13288
rect 19154 13232 19210 13288
rect 19614 13676 19616 13696
rect 19616 13676 19668 13696
rect 19668 13676 19670 13696
rect 19614 13640 19670 13676
rect 19216 13082 19272 13084
rect 19296 13082 19352 13084
rect 19376 13082 19432 13084
rect 19456 13082 19512 13084
rect 19216 13030 19262 13082
rect 19262 13030 19272 13082
rect 19296 13030 19326 13082
rect 19326 13030 19338 13082
rect 19338 13030 19352 13082
rect 19376 13030 19390 13082
rect 19390 13030 19402 13082
rect 19402 13030 19432 13082
rect 19456 13030 19466 13082
rect 19466 13030 19512 13082
rect 19216 13028 19272 13030
rect 19296 13028 19352 13030
rect 19376 13028 19432 13030
rect 19456 13028 19512 13030
rect 19876 14714 19932 14716
rect 19956 14714 20012 14716
rect 20036 14714 20092 14716
rect 20116 14714 20172 14716
rect 19876 14662 19922 14714
rect 19922 14662 19932 14714
rect 19956 14662 19986 14714
rect 19986 14662 19998 14714
rect 19998 14662 20012 14714
rect 20036 14662 20050 14714
rect 20050 14662 20062 14714
rect 20062 14662 20092 14714
rect 20116 14662 20126 14714
rect 20126 14662 20172 14714
rect 19876 14660 19932 14662
rect 19956 14660 20012 14662
rect 20036 14660 20092 14662
rect 20116 14660 20172 14662
rect 19430 12688 19486 12744
rect 18786 12008 18842 12064
rect 18050 9152 18106 9208
rect 17866 8064 17922 8120
rect 18694 11872 18750 11928
rect 18694 11756 18750 11792
rect 18694 11736 18696 11756
rect 18696 11736 18748 11756
rect 18748 11736 18750 11756
rect 18326 10240 18382 10296
rect 18234 9832 18290 9888
rect 18326 9696 18382 9752
rect 18234 8064 18290 8120
rect 17866 6976 17922 7032
rect 17682 6296 17738 6352
rect 17406 4392 17462 4448
rect 18142 6432 18198 6488
rect 17866 6160 17922 6216
rect 18786 11056 18842 11112
rect 18694 10412 18696 10432
rect 18696 10412 18748 10432
rect 18748 10412 18750 10432
rect 18694 10376 18750 10412
rect 19522 12416 19578 12472
rect 19216 11994 19272 11996
rect 19296 11994 19352 11996
rect 19376 11994 19432 11996
rect 19456 11994 19512 11996
rect 19216 11942 19262 11994
rect 19262 11942 19272 11994
rect 19296 11942 19326 11994
rect 19326 11942 19338 11994
rect 19338 11942 19352 11994
rect 19376 11942 19390 11994
rect 19390 11942 19402 11994
rect 19402 11942 19432 11994
rect 19456 11942 19466 11994
rect 19466 11942 19512 11994
rect 19216 11940 19272 11942
rect 19296 11940 19352 11942
rect 19376 11940 19432 11942
rect 19456 11940 19512 11942
rect 19522 11756 19578 11792
rect 19522 11736 19524 11756
rect 19524 11736 19576 11756
rect 19576 11736 19578 11756
rect 19522 11500 19524 11520
rect 19524 11500 19576 11520
rect 19576 11500 19578 11520
rect 19522 11464 19578 11500
rect 19890 13776 19946 13832
rect 21638 18400 21694 18456
rect 21086 17584 21142 17640
rect 20442 15680 20498 15736
rect 20534 14728 20590 14784
rect 20902 16652 20958 16688
rect 20902 16632 20904 16652
rect 20904 16632 20956 16652
rect 20956 16632 20958 16652
rect 20902 16224 20958 16280
rect 20534 13812 20536 13832
rect 20536 13812 20588 13832
rect 20588 13812 20590 13832
rect 20534 13776 20590 13812
rect 20258 13640 20314 13696
rect 19876 13626 19932 13628
rect 19956 13626 20012 13628
rect 20036 13626 20092 13628
rect 20116 13626 20172 13628
rect 19876 13574 19922 13626
rect 19922 13574 19932 13626
rect 19956 13574 19986 13626
rect 19986 13574 19998 13626
rect 19998 13574 20012 13626
rect 20036 13574 20050 13626
rect 20050 13574 20062 13626
rect 20062 13574 20092 13626
rect 20116 13574 20126 13626
rect 20126 13574 20172 13626
rect 19876 13572 19932 13574
rect 19956 13572 20012 13574
rect 20036 13572 20092 13574
rect 20116 13572 20172 13574
rect 19798 12724 19800 12744
rect 19800 12724 19852 12744
rect 19852 12724 19854 12744
rect 19798 12688 19854 12724
rect 20258 12960 20314 13016
rect 19706 12552 19762 12608
rect 19876 12538 19932 12540
rect 19956 12538 20012 12540
rect 20036 12538 20092 12540
rect 20116 12538 20172 12540
rect 19876 12486 19922 12538
rect 19922 12486 19932 12538
rect 19956 12486 19986 12538
rect 19986 12486 19998 12538
rect 19998 12486 20012 12538
rect 20036 12486 20050 12538
rect 20050 12486 20062 12538
rect 20062 12486 20092 12538
rect 20116 12486 20126 12538
rect 20126 12486 20172 12538
rect 19876 12484 19932 12486
rect 19956 12484 20012 12486
rect 20036 12484 20092 12486
rect 20116 12484 20172 12486
rect 19876 11450 19932 11452
rect 19956 11450 20012 11452
rect 20036 11450 20092 11452
rect 20116 11450 20172 11452
rect 19876 11398 19922 11450
rect 19922 11398 19932 11450
rect 19956 11398 19986 11450
rect 19986 11398 19998 11450
rect 19998 11398 20012 11450
rect 20036 11398 20050 11450
rect 20050 11398 20062 11450
rect 20062 11398 20092 11450
rect 20116 11398 20126 11450
rect 20126 11398 20172 11450
rect 19876 11396 19932 11398
rect 19956 11396 20012 11398
rect 20036 11396 20092 11398
rect 20116 11396 20172 11398
rect 19062 11056 19118 11112
rect 21086 17040 21142 17096
rect 21086 16940 21088 16960
rect 21088 16940 21140 16960
rect 21140 16940 21142 16960
rect 21086 16904 21142 16940
rect 20902 15272 20958 15328
rect 21178 15680 21234 15736
rect 21178 15408 21234 15464
rect 20994 15000 21050 15056
rect 20810 13776 20866 13832
rect 20534 12552 20590 12608
rect 20442 12416 20498 12472
rect 19216 10906 19272 10908
rect 19296 10906 19352 10908
rect 19376 10906 19432 10908
rect 19456 10906 19512 10908
rect 19216 10854 19262 10906
rect 19262 10854 19272 10906
rect 19296 10854 19326 10906
rect 19326 10854 19338 10906
rect 19338 10854 19352 10906
rect 19376 10854 19390 10906
rect 19390 10854 19402 10906
rect 19402 10854 19432 10906
rect 19456 10854 19466 10906
rect 19466 10854 19512 10906
rect 19216 10852 19272 10854
rect 19296 10852 19352 10854
rect 19376 10852 19432 10854
rect 19456 10852 19512 10854
rect 19246 10648 19302 10704
rect 18602 9324 18604 9344
rect 18604 9324 18656 9344
rect 18656 9324 18658 9344
rect 18602 9288 18658 9324
rect 18510 8744 18566 8800
rect 18510 8336 18566 8392
rect 19154 10376 19210 10432
rect 19430 10512 19486 10568
rect 19338 10240 19394 10296
rect 19614 10532 19670 10568
rect 19614 10512 19616 10532
rect 19616 10512 19668 10532
rect 19668 10512 19670 10532
rect 19614 10376 19670 10432
rect 19876 10362 19932 10364
rect 19956 10362 20012 10364
rect 20036 10362 20092 10364
rect 20116 10362 20172 10364
rect 19876 10310 19922 10362
rect 19922 10310 19932 10362
rect 19956 10310 19986 10362
rect 19986 10310 19998 10362
rect 19998 10310 20012 10362
rect 20036 10310 20050 10362
rect 20050 10310 20062 10362
rect 20062 10310 20092 10362
rect 20116 10310 20126 10362
rect 20126 10310 20172 10362
rect 19876 10308 19932 10310
rect 19956 10308 20012 10310
rect 20036 10308 20092 10310
rect 20116 10308 20172 10310
rect 19890 9968 19946 10024
rect 19216 9818 19272 9820
rect 19296 9818 19352 9820
rect 19376 9818 19432 9820
rect 19456 9818 19512 9820
rect 19216 9766 19262 9818
rect 19262 9766 19272 9818
rect 19296 9766 19326 9818
rect 19326 9766 19338 9818
rect 19338 9766 19352 9818
rect 19376 9766 19390 9818
rect 19390 9766 19402 9818
rect 19402 9766 19432 9818
rect 19456 9766 19466 9818
rect 19466 9766 19512 9818
rect 19216 9764 19272 9766
rect 19296 9764 19352 9766
rect 19376 9764 19432 9766
rect 19456 9764 19512 9766
rect 18878 9424 18934 9480
rect 18694 8744 18750 8800
rect 18694 8492 18750 8528
rect 18694 8472 18696 8492
rect 18696 8472 18748 8492
rect 18748 8472 18750 8492
rect 18786 8064 18842 8120
rect 18418 6024 18474 6080
rect 18786 7948 18842 7984
rect 18786 7928 18788 7948
rect 18788 7928 18840 7948
rect 18840 7928 18842 7948
rect 18970 9288 19026 9344
rect 18970 8084 19026 8120
rect 18970 8064 18972 8084
rect 18972 8064 19024 8084
rect 19024 8064 19026 8084
rect 18970 7248 19026 7304
rect 18878 6432 18934 6488
rect 18694 5480 18750 5536
rect 18970 6024 19026 6080
rect 19216 8730 19272 8732
rect 19296 8730 19352 8732
rect 19376 8730 19432 8732
rect 19456 8730 19512 8732
rect 19216 8678 19262 8730
rect 19262 8678 19272 8730
rect 19296 8678 19326 8730
rect 19326 8678 19338 8730
rect 19338 8678 19352 8730
rect 19376 8678 19390 8730
rect 19390 8678 19402 8730
rect 19402 8678 19432 8730
rect 19456 8678 19466 8730
rect 19466 8678 19512 8730
rect 19216 8676 19272 8678
rect 19296 8676 19352 8678
rect 19376 8676 19432 8678
rect 19456 8676 19512 8678
rect 19216 7642 19272 7644
rect 19296 7642 19352 7644
rect 19376 7642 19432 7644
rect 19456 7642 19512 7644
rect 19216 7590 19262 7642
rect 19262 7590 19272 7642
rect 19296 7590 19326 7642
rect 19326 7590 19338 7642
rect 19338 7590 19352 7642
rect 19376 7590 19390 7642
rect 19390 7590 19402 7642
rect 19402 7590 19432 7642
rect 19456 7590 19466 7642
rect 19466 7590 19512 7642
rect 19216 7588 19272 7590
rect 19296 7588 19352 7590
rect 19376 7588 19432 7590
rect 19456 7588 19512 7590
rect 19706 9288 19762 9344
rect 19706 9172 19762 9208
rect 19706 9152 19708 9172
rect 19708 9152 19760 9172
rect 19760 9152 19762 9172
rect 19890 9832 19946 9888
rect 19876 9274 19932 9276
rect 19956 9274 20012 9276
rect 20036 9274 20092 9276
rect 20116 9274 20172 9276
rect 19876 9222 19922 9274
rect 19922 9222 19932 9274
rect 19956 9222 19986 9274
rect 19986 9222 19998 9274
rect 19998 9222 20012 9274
rect 20036 9222 20050 9274
rect 20050 9222 20062 9274
rect 20062 9222 20092 9274
rect 20116 9222 20126 9274
rect 20126 9222 20172 9274
rect 19876 9220 19932 9222
rect 19956 9220 20012 9222
rect 20036 9220 20092 9222
rect 20116 9220 20172 9222
rect 19706 8744 19762 8800
rect 19706 8200 19762 8256
rect 20074 8356 20130 8392
rect 20074 8336 20076 8356
rect 20076 8336 20128 8356
rect 20128 8336 20130 8356
rect 20442 12008 20498 12064
rect 20534 11892 20590 11928
rect 20534 11872 20536 11892
rect 20536 11872 20588 11892
rect 20588 11872 20590 11892
rect 20442 10920 20498 10976
rect 20718 10376 20774 10432
rect 20718 10240 20774 10296
rect 21546 17584 21602 17640
rect 22190 18808 22246 18864
rect 21822 18128 21878 18184
rect 22006 17856 22062 17912
rect 21822 17312 21878 17368
rect 22834 20712 22890 20768
rect 23938 21256 23994 21312
rect 23018 19624 23074 19680
rect 22926 18944 22982 19000
rect 22374 18536 22430 18592
rect 22466 18128 22522 18184
rect 22374 17040 22430 17096
rect 22098 16768 22154 16824
rect 22190 16632 22246 16688
rect 21822 16496 21878 16552
rect 21730 16360 21786 16416
rect 21454 15988 21456 16008
rect 21456 15988 21508 16008
rect 21508 15988 21510 16008
rect 21454 15952 21510 15988
rect 21454 15272 21510 15328
rect 21454 15136 21510 15192
rect 21638 15952 21694 16008
rect 21822 15408 21878 15464
rect 21546 14184 21602 14240
rect 21730 14728 21786 14784
rect 21454 13912 21510 13968
rect 21822 13912 21878 13968
rect 21086 12824 21142 12880
rect 20994 12280 21050 12336
rect 20902 11192 20958 11248
rect 20994 10920 21050 10976
rect 20902 10240 20958 10296
rect 20442 9832 20498 9888
rect 20626 9832 20682 9888
rect 19876 8186 19932 8188
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 19876 8134 19922 8186
rect 19922 8134 19932 8186
rect 19956 8134 19986 8186
rect 19986 8134 19998 8186
rect 19998 8134 20012 8186
rect 20036 8134 20050 8186
rect 20050 8134 20062 8186
rect 20062 8134 20092 8186
rect 20116 8134 20126 8186
rect 20126 8134 20172 8186
rect 19876 8132 19932 8134
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 19798 7656 19854 7712
rect 20626 8780 20628 8800
rect 20628 8780 20680 8800
rect 20680 8780 20682 8800
rect 20626 8744 20682 8780
rect 20810 9560 20866 9616
rect 20902 9288 20958 9344
rect 20810 9152 20866 9208
rect 20810 9016 20866 9072
rect 20350 7520 20406 7576
rect 19216 6554 19272 6556
rect 19296 6554 19352 6556
rect 19376 6554 19432 6556
rect 19456 6554 19512 6556
rect 19216 6502 19262 6554
rect 19262 6502 19272 6554
rect 19296 6502 19326 6554
rect 19326 6502 19338 6554
rect 19338 6502 19352 6554
rect 19376 6502 19390 6554
rect 19390 6502 19402 6554
rect 19402 6502 19432 6554
rect 19456 6502 19466 6554
rect 19466 6502 19512 6554
rect 19216 6500 19272 6502
rect 19296 6500 19352 6502
rect 19376 6500 19432 6502
rect 19456 6500 19512 6502
rect 19430 6024 19486 6080
rect 18878 5344 18934 5400
rect 18326 4120 18382 4176
rect 19338 5652 19340 5672
rect 19340 5652 19392 5672
rect 19392 5652 19394 5672
rect 19338 5616 19394 5652
rect 19216 5466 19272 5468
rect 19296 5466 19352 5468
rect 19376 5466 19432 5468
rect 19456 5466 19512 5468
rect 19216 5414 19262 5466
rect 19262 5414 19272 5466
rect 19296 5414 19326 5466
rect 19326 5414 19338 5466
rect 19338 5414 19352 5466
rect 19376 5414 19390 5466
rect 19390 5414 19402 5466
rect 19402 5414 19432 5466
rect 19456 5414 19466 5466
rect 19466 5414 19512 5466
rect 19216 5412 19272 5414
rect 19296 5412 19352 5414
rect 19376 5412 19432 5414
rect 19456 5412 19512 5414
rect 19876 7098 19932 7100
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 19876 7046 19922 7098
rect 19922 7046 19932 7098
rect 19956 7046 19986 7098
rect 19986 7046 19998 7098
rect 19998 7046 20012 7098
rect 20036 7046 20050 7098
rect 20050 7046 20062 7098
rect 20062 7046 20092 7098
rect 20116 7046 20126 7098
rect 20126 7046 20172 7098
rect 19876 7044 19932 7046
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 19890 6840 19946 6896
rect 20166 6840 20222 6896
rect 19062 4800 19118 4856
rect 19890 6568 19946 6624
rect 19216 4378 19272 4380
rect 19296 4378 19352 4380
rect 19376 4378 19432 4380
rect 19456 4378 19512 4380
rect 19216 4326 19262 4378
rect 19262 4326 19272 4378
rect 19296 4326 19326 4378
rect 19326 4326 19338 4378
rect 19338 4326 19352 4378
rect 19376 4326 19390 4378
rect 19390 4326 19402 4378
rect 19402 4326 19432 4378
rect 19456 4326 19466 4378
rect 19466 4326 19512 4378
rect 19216 4324 19272 4326
rect 19296 4324 19352 4326
rect 19376 4324 19432 4326
rect 19456 4324 19512 4326
rect 19876 6010 19932 6012
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 19876 5958 19922 6010
rect 19922 5958 19932 6010
rect 19956 5958 19986 6010
rect 19986 5958 19998 6010
rect 19998 5958 20012 6010
rect 20036 5958 20050 6010
rect 20050 5958 20062 6010
rect 20062 5958 20092 6010
rect 20116 5958 20126 6010
rect 20126 5958 20172 6010
rect 19876 5956 19932 5958
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 19876 4922 19932 4924
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 19876 4870 19922 4922
rect 19922 4870 19932 4922
rect 19956 4870 19986 4922
rect 19986 4870 19998 4922
rect 19998 4870 20012 4922
rect 20036 4870 20050 4922
rect 20050 4870 20062 4922
rect 20062 4870 20092 4922
rect 20116 4870 20126 4922
rect 20126 4870 20172 4922
rect 19876 4868 19932 4870
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20626 7248 20682 7304
rect 20810 7284 20812 7304
rect 20812 7284 20864 7304
rect 20864 7284 20866 7304
rect 20810 7248 20866 7284
rect 20902 6840 20958 6896
rect 16486 3848 16542 3904
rect 20902 6568 20958 6624
rect 20902 5752 20958 5808
rect 20902 5344 20958 5400
rect 21454 13368 21510 13424
rect 21546 12824 21602 12880
rect 22098 16496 22154 16552
rect 22282 15988 22284 16008
rect 22284 15988 22336 16008
rect 22336 15988 22338 16008
rect 22282 15952 22338 15988
rect 22282 15136 22338 15192
rect 22190 13640 22246 13696
rect 22190 12824 22246 12880
rect 21270 8472 21326 8528
rect 21270 6296 21326 6352
rect 22190 12280 22246 12336
rect 22466 14612 22522 14648
rect 22466 14592 22468 14612
rect 22468 14592 22520 14612
rect 22520 14592 22522 14612
rect 22374 12552 22430 12608
rect 21454 10376 21510 10432
rect 22006 11056 22062 11112
rect 21914 9968 21970 10024
rect 21822 8880 21878 8936
rect 21638 8472 21694 8528
rect 21730 8064 21786 8120
rect 21454 7520 21510 7576
rect 21730 6976 21786 7032
rect 22190 11056 22246 11112
rect 22282 10804 22338 10840
rect 22282 10784 22284 10804
rect 22284 10784 22336 10804
rect 22336 10784 22338 10804
rect 22282 9560 22338 9616
rect 22098 8336 22154 8392
rect 22098 8200 22154 8256
rect 21822 6160 21878 6216
rect 20994 5072 21050 5128
rect 20810 4800 20866 4856
rect 19876 3834 19932 3836
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 19876 3782 19922 3834
rect 19922 3782 19932 3834
rect 19956 3782 19986 3834
rect 19986 3782 19998 3834
rect 19998 3782 20012 3834
rect 20036 3782 20050 3834
rect 20050 3782 20062 3834
rect 20062 3782 20092 3834
rect 20116 3782 20126 3834
rect 20126 3782 20172 3834
rect 19876 3780 19932 3782
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 22742 17076 22744 17096
rect 22744 17076 22796 17096
rect 22796 17076 22798 17096
rect 22742 17040 22798 17076
rect 23018 18536 23074 18592
rect 23386 18264 23442 18320
rect 23846 18808 23902 18864
rect 23938 18400 23994 18456
rect 23202 17720 23258 17776
rect 23110 17176 23166 17232
rect 23110 16904 23166 16960
rect 22834 16652 22890 16688
rect 22834 16632 22836 16652
rect 22836 16632 22888 16652
rect 22888 16632 22890 16652
rect 22926 16532 22928 16552
rect 22928 16532 22980 16552
rect 22980 16532 22982 16552
rect 22926 16496 22982 16532
rect 23202 16496 23258 16552
rect 23018 15544 23074 15600
rect 23846 18264 23902 18320
rect 23478 17992 23534 18048
rect 23386 17720 23442 17776
rect 23386 17176 23442 17232
rect 23662 16768 23718 16824
rect 22650 14864 22706 14920
rect 22742 13912 22798 13968
rect 22650 13232 22706 13288
rect 22650 12844 22706 12880
rect 22650 12824 22652 12844
rect 22652 12824 22704 12844
rect 22704 12824 22706 12844
rect 22742 11464 22798 11520
rect 22742 11192 22798 11248
rect 23202 14728 23258 14784
rect 23018 14320 23074 14376
rect 22742 10512 22798 10568
rect 22650 9968 22706 10024
rect 23202 13912 23258 13968
rect 23386 13912 23442 13968
rect 23110 13776 23166 13832
rect 23110 11464 23166 11520
rect 23018 10240 23074 10296
rect 23110 9968 23166 10024
rect 22650 9288 22706 9344
rect 22926 9016 22982 9072
rect 22650 8200 22706 8256
rect 22926 8064 22982 8120
rect 22558 7520 22614 7576
rect 22558 6976 22614 7032
rect 22374 6432 22430 6488
rect 21454 4664 21510 4720
rect 21822 4120 21878 4176
rect 19216 3290 19272 3292
rect 19296 3290 19352 3292
rect 19376 3290 19432 3292
rect 19456 3290 19512 3292
rect 19216 3238 19262 3290
rect 19262 3238 19272 3290
rect 19296 3238 19326 3290
rect 19326 3238 19338 3290
rect 19338 3238 19352 3290
rect 19376 3238 19390 3290
rect 19390 3238 19402 3290
rect 19402 3238 19432 3290
rect 19456 3238 19466 3290
rect 19466 3238 19512 3290
rect 19216 3236 19272 3238
rect 19296 3236 19352 3238
rect 19376 3236 19432 3238
rect 19456 3236 19512 3238
rect 22742 6840 22798 6896
rect 23018 7520 23074 7576
rect 23294 10376 23350 10432
rect 23294 9152 23350 9208
rect 23754 14864 23810 14920
rect 24582 20304 24638 20360
rect 24582 19624 24638 19680
rect 25318 19896 25374 19952
rect 26238 21392 26294 21448
rect 26146 20712 26202 20768
rect 25962 19760 26018 19816
rect 25870 19352 25926 19408
rect 25226 18844 25228 18864
rect 25228 18844 25280 18864
rect 25280 18844 25282 18864
rect 25226 18808 25282 18844
rect 25410 18808 25466 18864
rect 24398 17720 24454 17776
rect 24766 17176 24822 17232
rect 24490 16768 24546 16824
rect 24306 16108 24362 16144
rect 24306 16088 24308 16108
rect 24308 16088 24360 16108
rect 24360 16088 24362 16108
rect 24030 15156 24086 15192
rect 24030 15136 24032 15156
rect 24032 15136 24084 15156
rect 24084 15136 24086 15156
rect 23846 14728 23902 14784
rect 23754 14592 23810 14648
rect 23570 14048 23626 14104
rect 23662 12552 23718 12608
rect 23478 10512 23534 10568
rect 23662 10512 23718 10568
rect 24030 14476 24086 14512
rect 24030 14456 24032 14476
rect 24032 14456 24084 14476
rect 24084 14456 24086 14476
rect 24582 15816 24638 15872
rect 24306 15544 24362 15600
rect 24306 14476 24362 14512
rect 24306 14456 24308 14476
rect 24308 14456 24360 14476
rect 24360 14456 24362 14476
rect 24122 13640 24178 13696
rect 24214 13504 24270 13560
rect 24214 13132 24216 13152
rect 24216 13132 24268 13152
rect 24268 13132 24270 13152
rect 24214 13096 24270 13132
rect 24030 12144 24086 12200
rect 23938 11464 23994 11520
rect 24858 16632 24914 16688
rect 25962 18672 26018 18728
rect 26146 20032 26202 20088
rect 26990 21786 27046 21788
rect 27070 21786 27126 21788
rect 27150 21786 27206 21788
rect 27230 21786 27286 21788
rect 26990 21734 27036 21786
rect 27036 21734 27046 21786
rect 27070 21734 27100 21786
rect 27100 21734 27112 21786
rect 27112 21734 27126 21786
rect 27150 21734 27164 21786
rect 27164 21734 27176 21786
rect 27176 21734 27206 21786
rect 27230 21734 27240 21786
rect 27240 21734 27286 21786
rect 26990 21732 27046 21734
rect 27070 21732 27126 21734
rect 27150 21732 27206 21734
rect 27230 21732 27286 21734
rect 27650 21242 27706 21244
rect 27730 21242 27786 21244
rect 27810 21242 27866 21244
rect 27890 21242 27946 21244
rect 27650 21190 27696 21242
rect 27696 21190 27706 21242
rect 27730 21190 27760 21242
rect 27760 21190 27772 21242
rect 27772 21190 27786 21242
rect 27810 21190 27824 21242
rect 27824 21190 27836 21242
rect 27836 21190 27866 21242
rect 27890 21190 27900 21242
rect 27900 21190 27946 21242
rect 27650 21188 27706 21190
rect 27730 21188 27786 21190
rect 27810 21188 27866 21190
rect 27890 21188 27946 21190
rect 26990 20698 27046 20700
rect 27070 20698 27126 20700
rect 27150 20698 27206 20700
rect 27230 20698 27286 20700
rect 26990 20646 27036 20698
rect 27036 20646 27046 20698
rect 27070 20646 27100 20698
rect 27100 20646 27112 20698
rect 27112 20646 27126 20698
rect 27150 20646 27164 20698
rect 27164 20646 27176 20698
rect 27176 20646 27206 20698
rect 27230 20646 27240 20698
rect 27240 20646 27286 20698
rect 26990 20644 27046 20646
rect 27070 20644 27126 20646
rect 27150 20644 27206 20646
rect 27230 20644 27286 20646
rect 28078 20848 28134 20904
rect 26606 20304 26662 20360
rect 26422 20168 26478 20224
rect 26330 19624 26386 19680
rect 26146 19080 26202 19136
rect 26238 18944 26294 19000
rect 26606 19624 26662 19680
rect 27618 20440 27674 20496
rect 27158 20032 27214 20088
rect 25502 17856 25558 17912
rect 25410 17720 25466 17776
rect 25318 17584 25374 17640
rect 25226 17448 25282 17504
rect 24766 16088 24822 16144
rect 24766 15544 24822 15600
rect 24490 13776 24546 13832
rect 24490 13232 24546 13288
rect 24490 12960 24546 13016
rect 24030 11192 24086 11248
rect 23478 9696 23534 9752
rect 23294 8200 23350 8256
rect 21270 2896 21326 2952
rect 23938 9424 23994 9480
rect 23754 8744 23810 8800
rect 23754 8472 23810 8528
rect 23846 8356 23902 8392
rect 23846 8336 23848 8356
rect 23848 8336 23900 8356
rect 23900 8336 23902 8356
rect 23754 6704 23810 6760
rect 23662 6568 23718 6624
rect 23662 6296 23718 6352
rect 23662 5888 23718 5944
rect 24030 9288 24086 9344
rect 24030 8200 24086 8256
rect 24766 15272 24822 15328
rect 24766 14728 24822 14784
rect 24674 13504 24730 13560
rect 24674 13096 24730 13152
rect 24582 12280 24638 12336
rect 24398 11464 24454 11520
rect 24214 9460 24216 9480
rect 24216 9460 24268 9480
rect 24268 9460 24270 9480
rect 24214 9424 24270 9460
rect 24214 9152 24270 9208
rect 24490 9560 24546 9616
rect 24490 8744 24546 8800
rect 24398 8608 24454 8664
rect 24122 7928 24178 7984
rect 24214 7112 24270 7168
rect 24030 6296 24086 6352
rect 24030 5752 24086 5808
rect 24490 8064 24546 8120
rect 24582 7928 24638 7984
rect 24950 13640 25006 13696
rect 25410 16768 25466 16824
rect 25226 14864 25282 14920
rect 25134 14048 25190 14104
rect 24950 12960 25006 13016
rect 24950 12008 25006 12064
rect 24950 10784 25006 10840
rect 25318 13776 25374 13832
rect 25226 13504 25282 13560
rect 25318 13368 25374 13424
rect 25962 17584 26018 17640
rect 25962 17448 26018 17504
rect 25594 17040 25650 17096
rect 25686 16360 25742 16416
rect 25594 14592 25650 14648
rect 25134 12960 25190 13016
rect 25318 11736 25374 11792
rect 25502 12008 25558 12064
rect 25410 11464 25466 11520
rect 25134 11328 25190 11384
rect 24398 7112 24454 7168
rect 25226 10376 25282 10432
rect 25870 16360 25926 16416
rect 26238 17856 26294 17912
rect 26990 19610 27046 19612
rect 27070 19610 27126 19612
rect 27150 19610 27206 19612
rect 27230 19610 27286 19612
rect 26990 19558 27036 19610
rect 27036 19558 27046 19610
rect 27070 19558 27100 19610
rect 27100 19558 27112 19610
rect 27112 19558 27126 19610
rect 27150 19558 27164 19610
rect 27164 19558 27176 19610
rect 27176 19558 27206 19610
rect 27230 19558 27240 19610
rect 27240 19558 27286 19610
rect 26990 19556 27046 19558
rect 27070 19556 27126 19558
rect 27150 19556 27206 19558
rect 27230 19556 27286 19558
rect 26990 18522 27046 18524
rect 27070 18522 27126 18524
rect 27150 18522 27206 18524
rect 27230 18522 27286 18524
rect 26990 18470 27036 18522
rect 27036 18470 27046 18522
rect 27070 18470 27100 18522
rect 27100 18470 27112 18522
rect 27112 18470 27126 18522
rect 27150 18470 27164 18522
rect 27164 18470 27176 18522
rect 27176 18470 27206 18522
rect 27230 18470 27240 18522
rect 27240 18470 27286 18522
rect 26990 18468 27046 18470
rect 27070 18468 27126 18470
rect 27150 18468 27206 18470
rect 27230 18468 27286 18470
rect 26606 18128 26662 18184
rect 26422 17312 26478 17368
rect 26146 17176 26202 17232
rect 26330 17176 26386 17232
rect 26990 17434 27046 17436
rect 27070 17434 27126 17436
rect 27150 17434 27206 17436
rect 27230 17434 27286 17436
rect 26990 17382 27036 17434
rect 27036 17382 27046 17434
rect 27070 17382 27100 17434
rect 27100 17382 27112 17434
rect 27112 17382 27126 17434
rect 27150 17382 27164 17434
rect 27164 17382 27176 17434
rect 27176 17382 27206 17434
rect 27230 17382 27240 17434
rect 27240 17382 27286 17434
rect 26990 17380 27046 17382
rect 27070 17380 27126 17382
rect 27150 17380 27206 17382
rect 27230 17380 27286 17382
rect 25870 15136 25926 15192
rect 26330 16768 26386 16824
rect 26330 16632 26386 16688
rect 26238 16496 26294 16552
rect 26422 16496 26478 16552
rect 26422 16224 26478 16280
rect 25962 14612 26018 14648
rect 25962 14592 25964 14612
rect 25964 14592 26016 14612
rect 26016 14592 26018 14612
rect 25962 14184 26018 14240
rect 25962 13948 25964 13968
rect 25964 13948 26016 13968
rect 26016 13948 26018 13968
rect 25962 13912 26018 13948
rect 25870 13096 25926 13152
rect 25778 12300 25834 12336
rect 25778 12280 25780 12300
rect 25780 12280 25832 12300
rect 25832 12280 25834 12300
rect 25778 11600 25834 11656
rect 25778 11464 25834 11520
rect 25410 10240 25466 10296
rect 25134 8064 25190 8120
rect 24674 7384 24730 7440
rect 25042 7656 25098 7712
rect 25686 9560 25742 9616
rect 25778 9152 25834 9208
rect 25686 9016 25742 9072
rect 25502 7520 25558 7576
rect 24858 7112 24914 7168
rect 24582 6996 24638 7032
rect 24582 6976 24584 6996
rect 24584 6976 24636 6996
rect 24636 6976 24638 6996
rect 24858 6840 24914 6896
rect 23846 3440 23902 3496
rect 12102 2746 12158 2748
rect 12182 2746 12238 2748
rect 12262 2746 12318 2748
rect 12342 2746 12398 2748
rect 12102 2694 12148 2746
rect 12148 2694 12158 2746
rect 12182 2694 12212 2746
rect 12212 2694 12224 2746
rect 12224 2694 12238 2746
rect 12262 2694 12276 2746
rect 12276 2694 12288 2746
rect 12288 2694 12318 2746
rect 12342 2694 12352 2746
rect 12352 2694 12398 2746
rect 12102 2692 12158 2694
rect 12182 2692 12238 2694
rect 12262 2692 12318 2694
rect 12342 2692 12398 2694
rect 19876 2746 19932 2748
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 19876 2694 19922 2746
rect 19922 2694 19932 2746
rect 19956 2694 19986 2746
rect 19986 2694 19998 2746
rect 19998 2694 20012 2746
rect 20036 2694 20050 2746
rect 20050 2694 20062 2746
rect 20062 2694 20092 2746
rect 20116 2694 20126 2746
rect 20126 2694 20172 2746
rect 19876 2692 19932 2694
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 19706 2624 19762 2680
rect 10874 2352 10930 2408
rect 25318 7384 25374 7440
rect 25778 7112 25834 7168
rect 25686 6704 25742 6760
rect 25594 6432 25650 6488
rect 25962 11600 26018 11656
rect 25962 11056 26018 11112
rect 26238 13640 26294 13696
rect 26882 16632 26938 16688
rect 26698 15680 26754 15736
rect 26698 14592 26754 14648
rect 26698 14068 26754 14104
rect 26698 14048 26700 14068
rect 26700 14048 26752 14068
rect 26752 14048 26754 14068
rect 26698 13912 26754 13968
rect 26422 13096 26478 13152
rect 26330 12960 26386 13016
rect 27342 16904 27398 16960
rect 26990 16346 27046 16348
rect 27070 16346 27126 16348
rect 27150 16346 27206 16348
rect 27230 16346 27286 16348
rect 26990 16294 27036 16346
rect 27036 16294 27046 16346
rect 27070 16294 27100 16346
rect 27100 16294 27112 16346
rect 27112 16294 27126 16346
rect 27150 16294 27164 16346
rect 27164 16294 27176 16346
rect 27176 16294 27206 16346
rect 27230 16294 27240 16346
rect 27240 16294 27286 16346
rect 26990 16292 27046 16294
rect 27070 16292 27126 16294
rect 27150 16292 27206 16294
rect 27230 16292 27286 16294
rect 27066 15408 27122 15464
rect 26990 15258 27046 15260
rect 27070 15258 27126 15260
rect 27150 15258 27206 15260
rect 27230 15258 27286 15260
rect 26990 15206 27036 15258
rect 27036 15206 27046 15258
rect 27070 15206 27100 15258
rect 27100 15206 27112 15258
rect 27112 15206 27126 15258
rect 27150 15206 27164 15258
rect 27164 15206 27176 15258
rect 27176 15206 27206 15258
rect 27230 15206 27240 15258
rect 27240 15206 27286 15258
rect 26990 15204 27046 15206
rect 27070 15204 27126 15206
rect 27150 15204 27206 15206
rect 27230 15204 27286 15206
rect 26882 15000 26938 15056
rect 27650 20154 27706 20156
rect 27730 20154 27786 20156
rect 27810 20154 27866 20156
rect 27890 20154 27946 20156
rect 27650 20102 27696 20154
rect 27696 20102 27706 20154
rect 27730 20102 27760 20154
rect 27760 20102 27772 20154
rect 27772 20102 27786 20154
rect 27810 20102 27824 20154
rect 27824 20102 27836 20154
rect 27836 20102 27866 20154
rect 27890 20102 27900 20154
rect 27900 20102 27946 20154
rect 27650 20100 27706 20102
rect 27730 20100 27786 20102
rect 27810 20100 27866 20102
rect 27890 20100 27946 20102
rect 28170 20032 28226 20088
rect 28814 21392 28870 21448
rect 27650 19066 27706 19068
rect 27730 19066 27786 19068
rect 27810 19066 27866 19068
rect 27890 19066 27946 19068
rect 27650 19014 27696 19066
rect 27696 19014 27706 19066
rect 27730 19014 27760 19066
rect 27760 19014 27772 19066
rect 27772 19014 27786 19066
rect 27810 19014 27824 19066
rect 27824 19014 27836 19066
rect 27836 19014 27866 19066
rect 27890 19014 27900 19066
rect 27900 19014 27946 19066
rect 27650 19012 27706 19014
rect 27730 19012 27786 19014
rect 27810 19012 27866 19014
rect 27890 19012 27946 19014
rect 27710 18400 27766 18456
rect 27710 18164 27712 18184
rect 27712 18164 27764 18184
rect 27764 18164 27766 18184
rect 27710 18128 27766 18164
rect 27894 18164 27896 18184
rect 27896 18164 27948 18184
rect 27948 18164 27950 18184
rect 27894 18128 27950 18164
rect 27650 17978 27706 17980
rect 27730 17978 27786 17980
rect 27810 17978 27866 17980
rect 27890 17978 27946 17980
rect 27650 17926 27696 17978
rect 27696 17926 27706 17978
rect 27730 17926 27760 17978
rect 27760 17926 27772 17978
rect 27772 17926 27786 17978
rect 27810 17926 27824 17978
rect 27824 17926 27836 17978
rect 27836 17926 27866 17978
rect 27890 17926 27900 17978
rect 27900 17926 27946 17978
rect 27650 17924 27706 17926
rect 27730 17924 27786 17926
rect 27810 17924 27866 17926
rect 27890 17924 27946 17926
rect 28538 19624 28594 19680
rect 29274 21140 29330 21176
rect 29274 21120 29276 21140
rect 29276 21120 29328 21140
rect 29328 21120 29330 21140
rect 28906 20168 28962 20224
rect 28998 19760 29054 19816
rect 28722 19080 28778 19136
rect 27894 17448 27950 17504
rect 28354 17992 28410 18048
rect 27526 17332 27582 17368
rect 27526 17312 27528 17332
rect 27528 17312 27580 17332
rect 27580 17312 27582 17332
rect 28170 17448 28226 17504
rect 28078 17176 28134 17232
rect 27650 16890 27706 16892
rect 27730 16890 27786 16892
rect 27810 16890 27866 16892
rect 27890 16890 27946 16892
rect 27650 16838 27696 16890
rect 27696 16838 27706 16890
rect 27730 16838 27760 16890
rect 27760 16838 27772 16890
rect 27772 16838 27786 16890
rect 27810 16838 27824 16890
rect 27824 16838 27836 16890
rect 27836 16838 27866 16890
rect 27890 16838 27900 16890
rect 27900 16838 27946 16890
rect 27650 16836 27706 16838
rect 27730 16836 27786 16838
rect 27810 16836 27866 16838
rect 27890 16836 27946 16838
rect 28078 16904 28134 16960
rect 28078 16668 28080 16688
rect 28080 16668 28132 16688
rect 28132 16668 28134 16688
rect 28078 16632 28134 16668
rect 27618 16124 27620 16144
rect 27620 16124 27672 16144
rect 27672 16124 27674 16144
rect 27618 16088 27674 16124
rect 27986 16124 27988 16144
rect 27988 16124 28040 16144
rect 28040 16124 28042 16144
rect 27986 16088 28042 16124
rect 27650 15802 27706 15804
rect 27730 15802 27786 15804
rect 27810 15802 27866 15804
rect 27890 15802 27946 15804
rect 27650 15750 27696 15802
rect 27696 15750 27706 15802
rect 27730 15750 27760 15802
rect 27760 15750 27772 15802
rect 27772 15750 27786 15802
rect 27810 15750 27824 15802
rect 27824 15750 27836 15802
rect 27836 15750 27866 15802
rect 27890 15750 27900 15802
rect 27900 15750 27946 15802
rect 27650 15748 27706 15750
rect 27730 15748 27786 15750
rect 27810 15748 27866 15750
rect 27890 15748 27946 15750
rect 27894 14864 27950 14920
rect 27650 14714 27706 14716
rect 27730 14714 27786 14716
rect 27810 14714 27866 14716
rect 27890 14714 27946 14716
rect 27650 14662 27696 14714
rect 27696 14662 27706 14714
rect 27730 14662 27760 14714
rect 27760 14662 27772 14714
rect 27772 14662 27786 14714
rect 27810 14662 27824 14714
rect 27824 14662 27836 14714
rect 27836 14662 27866 14714
rect 27890 14662 27900 14714
rect 27900 14662 27946 14714
rect 27650 14660 27706 14662
rect 27730 14660 27786 14662
rect 27810 14660 27866 14662
rect 27890 14660 27946 14662
rect 29458 20032 29514 20088
rect 29550 19896 29606 19952
rect 29826 20440 29882 20496
rect 29826 20168 29882 20224
rect 28630 18164 28632 18184
rect 28632 18164 28684 18184
rect 28684 18164 28686 18184
rect 28630 18128 28686 18164
rect 28446 17312 28502 17368
rect 28354 16496 28410 16552
rect 28446 16088 28502 16144
rect 28446 15564 28502 15600
rect 28446 15544 28448 15564
rect 28448 15544 28500 15564
rect 28500 15544 28502 15564
rect 26974 14320 27030 14376
rect 26990 14170 27046 14172
rect 27070 14170 27126 14172
rect 27150 14170 27206 14172
rect 27230 14170 27286 14172
rect 26990 14118 27036 14170
rect 27036 14118 27046 14170
rect 27070 14118 27100 14170
rect 27100 14118 27112 14170
rect 27112 14118 27126 14170
rect 27150 14118 27164 14170
rect 27164 14118 27176 14170
rect 27176 14118 27206 14170
rect 27230 14118 27240 14170
rect 27240 14118 27286 14170
rect 26990 14116 27046 14118
rect 27070 14116 27126 14118
rect 27150 14116 27206 14118
rect 27230 14116 27286 14118
rect 26790 13640 26846 13696
rect 26146 12280 26202 12336
rect 26422 12144 26478 12200
rect 26330 11872 26386 11928
rect 26330 11464 26386 11520
rect 25962 10920 26018 10976
rect 26146 9832 26202 9888
rect 26330 10240 26386 10296
rect 26054 8472 26110 8528
rect 26698 12552 26754 12608
rect 26790 12144 26846 12200
rect 26974 13504 27030 13560
rect 26990 13082 27046 13084
rect 27070 13082 27126 13084
rect 27150 13082 27206 13084
rect 27230 13082 27286 13084
rect 26990 13030 27036 13082
rect 27036 13030 27046 13082
rect 27070 13030 27100 13082
rect 27100 13030 27112 13082
rect 27112 13030 27126 13082
rect 27150 13030 27164 13082
rect 27164 13030 27176 13082
rect 27176 13030 27206 13082
rect 27230 13030 27240 13082
rect 27240 13030 27286 13082
rect 26990 13028 27046 13030
rect 27070 13028 27126 13030
rect 27150 13028 27206 13030
rect 27230 13028 27286 13030
rect 26974 12844 27030 12880
rect 26974 12824 26976 12844
rect 26976 12824 27028 12844
rect 27028 12824 27030 12844
rect 27158 12280 27214 12336
rect 26990 11994 27046 11996
rect 27070 11994 27126 11996
rect 27150 11994 27206 11996
rect 27230 11994 27286 11996
rect 26990 11942 27036 11994
rect 27036 11942 27046 11994
rect 27070 11942 27100 11994
rect 27100 11942 27112 11994
rect 27112 11942 27126 11994
rect 27150 11942 27164 11994
rect 27164 11942 27176 11994
rect 27176 11942 27206 11994
rect 27230 11942 27240 11994
rect 27240 11942 27286 11994
rect 26990 11940 27046 11942
rect 27070 11940 27126 11942
rect 27150 11940 27206 11942
rect 27230 11940 27286 11942
rect 26882 11328 26938 11384
rect 27066 11192 27122 11248
rect 26990 10906 27046 10908
rect 27070 10906 27126 10908
rect 27150 10906 27206 10908
rect 27230 10906 27286 10908
rect 26990 10854 27036 10906
rect 27036 10854 27046 10906
rect 27070 10854 27100 10906
rect 27100 10854 27112 10906
rect 27112 10854 27126 10906
rect 27150 10854 27164 10906
rect 27164 10854 27176 10906
rect 27176 10854 27206 10906
rect 27230 10854 27240 10906
rect 27240 10854 27286 10906
rect 26990 10852 27046 10854
rect 27070 10852 27126 10854
rect 27150 10852 27206 10854
rect 27230 10852 27286 10854
rect 26606 10004 26608 10024
rect 26608 10004 26660 10024
rect 26660 10004 26662 10024
rect 26606 9968 26662 10004
rect 26698 9696 26754 9752
rect 26514 9152 26570 9208
rect 26514 9016 26570 9072
rect 26422 8608 26478 8664
rect 25962 8200 26018 8256
rect 25410 5208 25466 5264
rect 26238 8200 26294 8256
rect 26238 7792 26294 7848
rect 24858 2624 24914 2680
rect 19706 2216 19762 2272
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 11442 2202 11498 2204
rect 11522 2202 11578 2204
rect 11602 2202 11658 2204
rect 11682 2202 11738 2204
rect 11442 2150 11488 2202
rect 11488 2150 11498 2202
rect 11522 2150 11552 2202
rect 11552 2150 11564 2202
rect 11564 2150 11578 2202
rect 11602 2150 11616 2202
rect 11616 2150 11628 2202
rect 11628 2150 11658 2202
rect 11682 2150 11692 2202
rect 11692 2150 11738 2202
rect 11442 2148 11498 2150
rect 11522 2148 11578 2150
rect 11602 2148 11658 2150
rect 11682 2148 11738 2150
rect 19216 2202 19272 2204
rect 19296 2202 19352 2204
rect 19376 2202 19432 2204
rect 19456 2202 19512 2204
rect 19216 2150 19262 2202
rect 19262 2150 19272 2202
rect 19296 2150 19326 2202
rect 19326 2150 19338 2202
rect 19338 2150 19352 2202
rect 19376 2150 19390 2202
rect 19390 2150 19402 2202
rect 19402 2150 19432 2202
rect 19456 2150 19466 2202
rect 19466 2150 19512 2202
rect 19216 2148 19272 2150
rect 19296 2148 19352 2150
rect 19376 2148 19432 2150
rect 19456 2148 19512 2150
rect 26514 7692 26516 7712
rect 26516 7692 26568 7712
rect 26568 7692 26570 7712
rect 26514 7656 26570 7692
rect 27066 10376 27122 10432
rect 26974 10240 27030 10296
rect 26990 9818 27046 9820
rect 27070 9818 27126 9820
rect 27150 9818 27206 9820
rect 27230 9818 27286 9820
rect 26990 9766 27036 9818
rect 27036 9766 27046 9818
rect 27070 9766 27100 9818
rect 27100 9766 27112 9818
rect 27112 9766 27126 9818
rect 27150 9766 27164 9818
rect 27164 9766 27176 9818
rect 27176 9766 27206 9818
rect 27230 9766 27240 9818
rect 27240 9766 27286 9818
rect 26990 9764 27046 9766
rect 27070 9764 27126 9766
rect 27150 9764 27206 9766
rect 27230 9764 27286 9766
rect 28354 15408 28410 15464
rect 28630 16904 28686 16960
rect 28998 17040 29054 17096
rect 28906 16788 28962 16824
rect 28906 16768 28908 16788
rect 28908 16768 28960 16788
rect 28960 16768 28962 16788
rect 28446 14864 28502 14920
rect 28262 14456 28318 14512
rect 27650 13626 27706 13628
rect 27730 13626 27786 13628
rect 27810 13626 27866 13628
rect 27890 13626 27946 13628
rect 27650 13574 27696 13626
rect 27696 13574 27706 13626
rect 27730 13574 27760 13626
rect 27760 13574 27772 13626
rect 27772 13574 27786 13626
rect 27810 13574 27824 13626
rect 27824 13574 27836 13626
rect 27836 13574 27866 13626
rect 27890 13574 27900 13626
rect 27900 13574 27946 13626
rect 27650 13572 27706 13574
rect 27730 13572 27786 13574
rect 27810 13572 27866 13574
rect 27890 13572 27946 13574
rect 27618 13096 27674 13152
rect 27986 13232 28042 13288
rect 27650 12538 27706 12540
rect 27730 12538 27786 12540
rect 27810 12538 27866 12540
rect 27890 12538 27946 12540
rect 27650 12486 27696 12538
rect 27696 12486 27706 12538
rect 27730 12486 27760 12538
rect 27760 12486 27772 12538
rect 27772 12486 27786 12538
rect 27810 12486 27824 12538
rect 27824 12486 27836 12538
rect 27836 12486 27866 12538
rect 27890 12486 27900 12538
rect 27900 12486 27946 12538
rect 27650 12484 27706 12486
rect 27730 12484 27786 12486
rect 27810 12484 27866 12486
rect 27890 12484 27946 12486
rect 28078 12688 28134 12744
rect 27618 12144 27674 12200
rect 27710 11872 27766 11928
rect 27986 12280 28042 12336
rect 27618 11600 27674 11656
rect 27802 11600 27858 11656
rect 27650 11450 27706 11452
rect 27730 11450 27786 11452
rect 27810 11450 27866 11452
rect 27890 11450 27946 11452
rect 27650 11398 27696 11450
rect 27696 11398 27706 11450
rect 27730 11398 27760 11450
rect 27760 11398 27772 11450
rect 27772 11398 27786 11450
rect 27810 11398 27824 11450
rect 27824 11398 27836 11450
rect 27836 11398 27866 11450
rect 27890 11398 27900 11450
rect 27900 11398 27946 11450
rect 27650 11396 27706 11398
rect 27730 11396 27786 11398
rect 27810 11396 27866 11398
rect 27890 11396 27946 11398
rect 26974 9288 27030 9344
rect 27526 11212 27582 11248
rect 27526 11192 27528 11212
rect 27528 11192 27580 11212
rect 27580 11192 27582 11212
rect 27618 11056 27674 11112
rect 28906 16632 28962 16688
rect 28906 16088 28962 16144
rect 28998 15136 29054 15192
rect 29274 17076 29276 17096
rect 29276 17076 29328 17096
rect 29328 17076 29330 17096
rect 29274 17040 29330 17076
rect 29274 16496 29330 16552
rect 29274 15544 29330 15600
rect 29458 19216 29514 19272
rect 29734 19352 29790 19408
rect 29734 19080 29790 19136
rect 29458 18808 29514 18864
rect 29734 17992 29790 18048
rect 29550 17312 29606 17368
rect 29458 17176 29514 17232
rect 29550 16224 29606 16280
rect 29458 15972 29514 16008
rect 29458 15952 29460 15972
rect 29460 15952 29512 15972
rect 29512 15952 29514 15972
rect 29274 14900 29276 14920
rect 29276 14900 29328 14920
rect 29328 14900 29330 14920
rect 29274 14864 29330 14900
rect 28814 13912 28870 13968
rect 29182 13096 29238 13152
rect 28170 11600 28226 11656
rect 27650 10362 27706 10364
rect 27730 10362 27786 10364
rect 27810 10362 27866 10364
rect 27890 10362 27946 10364
rect 27650 10310 27696 10362
rect 27696 10310 27706 10362
rect 27730 10310 27760 10362
rect 27760 10310 27772 10362
rect 27772 10310 27786 10362
rect 27810 10310 27824 10362
rect 27824 10310 27836 10362
rect 27836 10310 27866 10362
rect 27890 10310 27900 10362
rect 27900 10310 27946 10362
rect 27650 10308 27706 10310
rect 27730 10308 27786 10310
rect 27810 10308 27866 10310
rect 27890 10308 27946 10310
rect 27986 10104 28042 10160
rect 27618 9968 27674 10024
rect 28262 11212 28318 11248
rect 28262 11192 28264 11212
rect 28264 11192 28316 11212
rect 28316 11192 28318 11212
rect 28906 12688 28962 12744
rect 29182 12416 29238 12472
rect 29090 12316 29092 12336
rect 29092 12316 29144 12336
rect 29144 12316 29146 12336
rect 29090 12280 29146 12316
rect 27986 9580 28042 9616
rect 27986 9560 27988 9580
rect 27988 9560 28040 9580
rect 28040 9560 28042 9580
rect 27650 9274 27706 9276
rect 27730 9274 27786 9276
rect 27810 9274 27866 9276
rect 27890 9274 27946 9276
rect 27650 9222 27696 9274
rect 27696 9222 27706 9274
rect 27730 9222 27760 9274
rect 27760 9222 27772 9274
rect 27772 9222 27786 9274
rect 27810 9222 27824 9274
rect 27824 9222 27836 9274
rect 27836 9222 27866 9274
rect 27890 9222 27900 9274
rect 27900 9222 27946 9274
rect 27650 9220 27706 9222
rect 27730 9220 27786 9222
rect 27810 9220 27866 9222
rect 27890 9220 27946 9222
rect 27526 8880 27582 8936
rect 28446 9152 28502 9208
rect 26990 8730 27046 8732
rect 27070 8730 27126 8732
rect 27150 8730 27206 8732
rect 27230 8730 27286 8732
rect 26990 8678 27036 8730
rect 27036 8678 27046 8730
rect 27070 8678 27100 8730
rect 27100 8678 27112 8730
rect 27112 8678 27126 8730
rect 27150 8678 27164 8730
rect 27164 8678 27176 8730
rect 27176 8678 27206 8730
rect 27230 8678 27240 8730
rect 27240 8678 27286 8730
rect 26990 8676 27046 8678
rect 27070 8676 27126 8678
rect 27150 8676 27206 8678
rect 27230 8676 27286 8678
rect 26698 8336 26754 8392
rect 26698 8064 26754 8120
rect 26974 8472 27030 8528
rect 27066 8200 27122 8256
rect 26990 7642 27046 7644
rect 27070 7642 27126 7644
rect 27150 7642 27206 7644
rect 27230 7642 27286 7644
rect 26990 7590 27036 7642
rect 27036 7590 27046 7642
rect 27070 7590 27100 7642
rect 27100 7590 27112 7642
rect 27112 7590 27126 7642
rect 27150 7590 27164 7642
rect 27164 7590 27176 7642
rect 27176 7590 27206 7642
rect 27230 7590 27240 7642
rect 27240 7590 27286 7642
rect 26990 7588 27046 7590
rect 27070 7588 27126 7590
rect 27150 7588 27206 7590
rect 27230 7588 27286 7590
rect 27894 8472 27950 8528
rect 27434 7284 27436 7304
rect 27436 7284 27488 7304
rect 27488 7284 27490 7304
rect 27434 7248 27490 7284
rect 26990 6554 27046 6556
rect 27070 6554 27126 6556
rect 27150 6554 27206 6556
rect 27230 6554 27286 6556
rect 26990 6502 27036 6554
rect 27036 6502 27046 6554
rect 27070 6502 27100 6554
rect 27100 6502 27112 6554
rect 27112 6502 27126 6554
rect 27150 6502 27164 6554
rect 27164 6502 27176 6554
rect 27176 6502 27206 6554
rect 27230 6502 27240 6554
rect 27240 6502 27286 6554
rect 26990 6500 27046 6502
rect 27070 6500 27126 6502
rect 27150 6500 27206 6502
rect 27230 6500 27286 6502
rect 26882 5636 26938 5672
rect 26882 5616 26884 5636
rect 26884 5616 26936 5636
rect 26936 5616 26938 5636
rect 26990 5466 27046 5468
rect 27070 5466 27126 5468
rect 27150 5466 27206 5468
rect 27230 5466 27286 5468
rect 26990 5414 27036 5466
rect 27036 5414 27046 5466
rect 27070 5414 27100 5466
rect 27100 5414 27112 5466
rect 27112 5414 27126 5466
rect 27150 5414 27164 5466
rect 27164 5414 27176 5466
rect 27176 5414 27206 5466
rect 27230 5414 27240 5466
rect 27240 5414 27286 5466
rect 26990 5412 27046 5414
rect 27070 5412 27126 5414
rect 27150 5412 27206 5414
rect 27230 5412 27286 5414
rect 27802 8336 27858 8392
rect 27650 8186 27706 8188
rect 27730 8186 27786 8188
rect 27810 8186 27866 8188
rect 27890 8186 27946 8188
rect 27650 8134 27696 8186
rect 27696 8134 27706 8186
rect 27730 8134 27760 8186
rect 27760 8134 27772 8186
rect 27772 8134 27786 8186
rect 27810 8134 27824 8186
rect 27824 8134 27836 8186
rect 27836 8134 27866 8186
rect 27890 8134 27900 8186
rect 27900 8134 27946 8186
rect 27650 8132 27706 8134
rect 27730 8132 27786 8134
rect 27810 8132 27866 8134
rect 27890 8132 27946 8134
rect 27986 7792 28042 7848
rect 27650 7098 27706 7100
rect 27730 7098 27786 7100
rect 27810 7098 27866 7100
rect 27890 7098 27946 7100
rect 27650 7046 27696 7098
rect 27696 7046 27706 7098
rect 27730 7046 27760 7098
rect 27760 7046 27772 7098
rect 27772 7046 27786 7098
rect 27810 7046 27824 7098
rect 27824 7046 27836 7098
rect 27836 7046 27866 7098
rect 27890 7046 27900 7098
rect 27900 7046 27946 7098
rect 27650 7044 27706 7046
rect 27730 7044 27786 7046
rect 27810 7044 27866 7046
rect 27890 7044 27946 7046
rect 27650 6010 27706 6012
rect 27730 6010 27786 6012
rect 27810 6010 27866 6012
rect 27890 6010 27946 6012
rect 27650 5958 27696 6010
rect 27696 5958 27706 6010
rect 27730 5958 27760 6010
rect 27760 5958 27772 6010
rect 27772 5958 27786 6010
rect 27810 5958 27824 6010
rect 27824 5958 27836 6010
rect 27836 5958 27866 6010
rect 27890 5958 27900 6010
rect 27900 5958 27946 6010
rect 27650 5956 27706 5958
rect 27730 5956 27786 5958
rect 27810 5956 27866 5958
rect 27890 5956 27946 5958
rect 28170 7656 28226 7712
rect 28630 9560 28686 9616
rect 29274 11872 29330 11928
rect 28630 7948 28686 7984
rect 28630 7928 28632 7948
rect 28632 7928 28684 7948
rect 28684 7928 28686 7948
rect 29550 15020 29606 15056
rect 29550 15000 29552 15020
rect 29552 15000 29604 15020
rect 29604 15000 29606 15020
rect 30838 21120 30894 21176
rect 30838 20340 30840 20360
rect 30840 20340 30892 20360
rect 30892 20340 30894 20360
rect 30194 19216 30250 19272
rect 30838 20304 30894 20340
rect 30470 18128 30526 18184
rect 30378 17584 30434 17640
rect 29918 14764 29920 14784
rect 29920 14764 29972 14784
rect 29972 14764 29974 14784
rect 29918 14728 29974 14764
rect 29826 12824 29882 12880
rect 30378 15408 30434 15464
rect 30562 16360 30618 16416
rect 30286 15308 30288 15328
rect 30288 15308 30340 15328
rect 30340 15308 30342 15328
rect 30286 15272 30342 15308
rect 30286 15136 30342 15192
rect 31206 19624 31262 19680
rect 30930 19216 30986 19272
rect 30746 18400 30802 18456
rect 30838 18128 30894 18184
rect 31298 18264 31354 18320
rect 31574 20304 31630 20360
rect 31482 18672 31538 18728
rect 31114 17584 31170 17640
rect 30378 13776 30434 13832
rect 30286 13096 30342 13152
rect 30654 11872 30710 11928
rect 29734 9288 29790 9344
rect 29458 8336 29514 8392
rect 29274 8200 29330 8256
rect 28722 6704 28778 6760
rect 28538 5072 28594 5128
rect 27650 4922 27706 4924
rect 27730 4922 27786 4924
rect 27810 4922 27866 4924
rect 27890 4922 27946 4924
rect 27650 4870 27696 4922
rect 27696 4870 27706 4922
rect 27730 4870 27760 4922
rect 27760 4870 27772 4922
rect 27772 4870 27786 4922
rect 27810 4870 27824 4922
rect 27824 4870 27836 4922
rect 27836 4870 27866 4922
rect 27890 4870 27900 4922
rect 27900 4870 27946 4922
rect 27650 4868 27706 4870
rect 27730 4868 27786 4870
rect 27810 4868 27866 4870
rect 27890 4868 27946 4870
rect 26990 4378 27046 4380
rect 27070 4378 27126 4380
rect 27150 4378 27206 4380
rect 27230 4378 27286 4380
rect 26990 4326 27036 4378
rect 27036 4326 27046 4378
rect 27070 4326 27100 4378
rect 27100 4326 27112 4378
rect 27112 4326 27126 4378
rect 27150 4326 27164 4378
rect 27164 4326 27176 4378
rect 27176 4326 27206 4378
rect 27230 4326 27240 4378
rect 27240 4326 27286 4378
rect 26990 4324 27046 4326
rect 27070 4324 27126 4326
rect 27150 4324 27206 4326
rect 27230 4324 27286 4326
rect 27650 3834 27706 3836
rect 27730 3834 27786 3836
rect 27810 3834 27866 3836
rect 27890 3834 27946 3836
rect 27650 3782 27696 3834
rect 27696 3782 27706 3834
rect 27730 3782 27760 3834
rect 27760 3782 27772 3834
rect 27772 3782 27786 3834
rect 27810 3782 27824 3834
rect 27824 3782 27836 3834
rect 27836 3782 27866 3834
rect 27890 3782 27900 3834
rect 27900 3782 27946 3834
rect 27650 3780 27706 3782
rect 27730 3780 27786 3782
rect 27810 3780 27866 3782
rect 27890 3780 27946 3782
rect 26990 3290 27046 3292
rect 27070 3290 27126 3292
rect 27150 3290 27206 3292
rect 27230 3290 27286 3292
rect 26990 3238 27036 3290
rect 27036 3238 27046 3290
rect 27070 3238 27100 3290
rect 27100 3238 27112 3290
rect 27112 3238 27126 3290
rect 27150 3238 27164 3290
rect 27164 3238 27176 3290
rect 27176 3238 27206 3290
rect 27230 3238 27240 3290
rect 27240 3238 27286 3290
rect 26990 3236 27046 3238
rect 27070 3236 27126 3238
rect 27150 3236 27206 3238
rect 27230 3236 27286 3238
rect 29458 6160 29514 6216
rect 30378 10684 30380 10704
rect 30380 10684 30432 10704
rect 30432 10684 30434 10704
rect 30378 10648 30434 10684
rect 30378 8916 30380 8936
rect 30380 8916 30432 8936
rect 30432 8916 30434 8936
rect 30378 8880 30434 8916
rect 29918 8336 29974 8392
rect 29642 5752 29698 5808
rect 31114 16652 31170 16688
rect 31114 16632 31116 16652
rect 31116 16632 31168 16652
rect 31168 16632 31170 16652
rect 31390 14864 31446 14920
rect 30746 9560 30802 9616
rect 30562 7384 30618 7440
rect 31022 8200 31078 8256
rect 30930 6296 30986 6352
rect 31666 17448 31722 17504
rect 28998 3032 29054 3088
rect 27650 2746 27706 2748
rect 27730 2746 27786 2748
rect 27810 2746 27866 2748
rect 27890 2746 27946 2748
rect 27650 2694 27696 2746
rect 27696 2694 27706 2746
rect 27730 2694 27760 2746
rect 27760 2694 27772 2746
rect 27772 2694 27786 2746
rect 27810 2694 27824 2746
rect 27824 2694 27836 2746
rect 27836 2694 27866 2746
rect 27890 2694 27900 2746
rect 27900 2694 27946 2746
rect 27650 2692 27706 2694
rect 27730 2692 27786 2694
rect 27810 2692 27866 2694
rect 27890 2692 27946 2694
rect 26990 2202 27046 2204
rect 27070 2202 27126 2204
rect 27150 2202 27206 2204
rect 27230 2202 27286 2204
rect 26990 2150 27036 2202
rect 27036 2150 27046 2202
rect 27070 2150 27100 2202
rect 27100 2150 27112 2202
rect 27112 2150 27126 2202
rect 27150 2150 27164 2202
rect 27164 2150 27176 2202
rect 27176 2150 27206 2202
rect 27230 2150 27240 2202
rect 27240 2150 27286 2202
rect 26990 2148 27046 2150
rect 27070 2148 27126 2150
rect 27150 2148 27206 2150
rect 27230 2148 27286 2150
rect 26422 1944 26478 2000
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 12102 1658 12158 1660
rect 12182 1658 12238 1660
rect 12262 1658 12318 1660
rect 12342 1658 12398 1660
rect 12102 1606 12148 1658
rect 12148 1606 12158 1658
rect 12182 1606 12212 1658
rect 12212 1606 12224 1658
rect 12224 1606 12238 1658
rect 12262 1606 12276 1658
rect 12276 1606 12288 1658
rect 12288 1606 12318 1658
rect 12342 1606 12352 1658
rect 12352 1606 12398 1658
rect 12102 1604 12158 1606
rect 12182 1604 12238 1606
rect 12262 1604 12318 1606
rect 12342 1604 12398 1606
rect 19876 1658 19932 1660
rect 19956 1658 20012 1660
rect 20036 1658 20092 1660
rect 20116 1658 20172 1660
rect 19876 1606 19922 1658
rect 19922 1606 19932 1658
rect 19956 1606 19986 1658
rect 19986 1606 19998 1658
rect 19998 1606 20012 1658
rect 20036 1606 20050 1658
rect 20050 1606 20062 1658
rect 20062 1606 20092 1658
rect 20116 1606 20126 1658
rect 20126 1606 20172 1658
rect 19876 1604 19932 1606
rect 19956 1604 20012 1606
rect 20036 1604 20092 1606
rect 20116 1604 20172 1606
rect 27650 1658 27706 1660
rect 27730 1658 27786 1660
rect 27810 1658 27866 1660
rect 27890 1658 27946 1660
rect 27650 1606 27696 1658
rect 27696 1606 27706 1658
rect 27730 1606 27760 1658
rect 27760 1606 27772 1658
rect 27772 1606 27786 1658
rect 27810 1606 27824 1658
rect 27824 1606 27836 1658
rect 27836 1606 27866 1658
rect 27890 1606 27900 1658
rect 27900 1606 27946 1658
rect 27650 1604 27706 1606
rect 27730 1604 27786 1606
rect 27810 1604 27866 1606
rect 27890 1604 27946 1606
rect 1122 1400 1178 1456
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 11442 1114 11498 1116
rect 11522 1114 11578 1116
rect 11602 1114 11658 1116
rect 11682 1114 11738 1116
rect 11442 1062 11488 1114
rect 11488 1062 11498 1114
rect 11522 1062 11552 1114
rect 11552 1062 11564 1114
rect 11564 1062 11578 1114
rect 11602 1062 11616 1114
rect 11616 1062 11628 1114
rect 11628 1062 11658 1114
rect 11682 1062 11692 1114
rect 11692 1062 11738 1114
rect 11442 1060 11498 1062
rect 11522 1060 11578 1062
rect 11602 1060 11658 1062
rect 11682 1060 11738 1062
rect 19216 1114 19272 1116
rect 19296 1114 19352 1116
rect 19376 1114 19432 1116
rect 19456 1114 19512 1116
rect 19216 1062 19262 1114
rect 19262 1062 19272 1114
rect 19296 1062 19326 1114
rect 19326 1062 19338 1114
rect 19338 1062 19352 1114
rect 19376 1062 19390 1114
rect 19390 1062 19402 1114
rect 19402 1062 19432 1114
rect 19456 1062 19466 1114
rect 19466 1062 19512 1114
rect 19216 1060 19272 1062
rect 19296 1060 19352 1062
rect 19376 1060 19432 1062
rect 19456 1060 19512 1062
rect 26990 1114 27046 1116
rect 27070 1114 27126 1116
rect 27150 1114 27206 1116
rect 27230 1114 27286 1116
rect 26990 1062 27036 1114
rect 27036 1062 27046 1114
rect 27070 1062 27100 1114
rect 27100 1062 27112 1114
rect 27112 1062 27126 1114
rect 27150 1062 27164 1114
rect 27164 1062 27176 1114
rect 27176 1062 27206 1114
rect 27230 1062 27240 1114
rect 27240 1062 27286 1114
rect 26990 1060 27046 1062
rect 27070 1060 27126 1062
rect 27150 1060 27206 1062
rect 27230 1060 27286 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 12102 570 12158 572
rect 12182 570 12238 572
rect 12262 570 12318 572
rect 12342 570 12398 572
rect 12102 518 12148 570
rect 12148 518 12158 570
rect 12182 518 12212 570
rect 12212 518 12224 570
rect 12224 518 12238 570
rect 12262 518 12276 570
rect 12276 518 12288 570
rect 12288 518 12318 570
rect 12342 518 12352 570
rect 12352 518 12398 570
rect 12102 516 12158 518
rect 12182 516 12238 518
rect 12262 516 12318 518
rect 12342 516 12398 518
rect 19876 570 19932 572
rect 19956 570 20012 572
rect 20036 570 20092 572
rect 20116 570 20172 572
rect 19876 518 19922 570
rect 19922 518 19932 570
rect 19956 518 19986 570
rect 19986 518 19998 570
rect 19998 518 20012 570
rect 20036 518 20050 570
rect 20050 518 20062 570
rect 20062 518 20092 570
rect 20116 518 20126 570
rect 20126 518 20172 570
rect 19876 516 19932 518
rect 19956 516 20012 518
rect 20036 516 20092 518
rect 20116 516 20172 518
rect 27650 570 27706 572
rect 27730 570 27786 572
rect 27810 570 27866 572
rect 27890 570 27946 572
rect 27650 518 27696 570
rect 27696 518 27706 570
rect 27730 518 27760 570
rect 27760 518 27772 570
rect 27772 518 27786 570
rect 27810 518 27824 570
rect 27824 518 27836 570
rect 27836 518 27866 570
rect 27890 518 27900 570
rect 27900 518 27946 570
rect 27650 516 27706 518
rect 27730 516 27786 518
rect 27810 516 27866 518
rect 27890 516 27946 518
<< metal3 >>
rect 6545 22130 6611 22133
rect 20294 22130 20300 22132
rect 6545 22128 20300 22130
rect 6545 22072 6550 22128
rect 6606 22072 20300 22128
rect 6545 22070 20300 22072
rect 6545 22067 6611 22070
rect 20294 22068 20300 22070
rect 20364 22068 20370 22132
rect 11646 21932 11652 21996
rect 11716 21994 11722 21996
rect 11881 21994 11947 21997
rect 12249 21996 12315 21997
rect 11716 21992 11947 21994
rect 11716 21936 11886 21992
rect 11942 21936 11947 21992
rect 11716 21934 11947 21936
rect 11716 21932 11722 21934
rect 11881 21931 11947 21934
rect 12198 21932 12204 21996
rect 12268 21994 12315 21996
rect 24342 21994 24348 21996
rect 12268 21992 12360 21994
rect 12310 21936 12360 21992
rect 12268 21934 12360 21936
rect 17174 21934 24348 21994
rect 12268 21932 12315 21934
rect 12249 21931 12315 21932
rect 8886 21796 8892 21860
rect 8956 21858 8962 21860
rect 9581 21858 9647 21861
rect 8956 21856 9647 21858
rect 8956 21800 9586 21856
rect 9642 21800 9647 21856
rect 8956 21798 9647 21800
rect 8956 21796 8962 21798
rect 9581 21795 9647 21798
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 11432 21792 11748 21793
rect 11432 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11748 21792
rect 11432 21727 11748 21728
rect 6177 21724 6243 21725
rect 6729 21724 6795 21725
rect 7281 21724 7347 21725
rect 7833 21724 7899 21725
rect 8385 21724 8451 21725
rect 9489 21724 9555 21725
rect 10041 21724 10107 21725
rect 10593 21724 10659 21725
rect 11145 21724 11211 21725
rect 12801 21724 12867 21725
rect 13353 21724 13419 21725
rect 13905 21724 13971 21725
rect 16665 21724 16731 21725
rect 6126 21660 6132 21724
rect 6196 21722 6243 21724
rect 6196 21720 6288 21722
rect 6238 21664 6288 21720
rect 6196 21662 6288 21664
rect 6196 21660 6243 21662
rect 6678 21660 6684 21724
rect 6748 21722 6795 21724
rect 6748 21720 6840 21722
rect 6790 21664 6840 21720
rect 6748 21662 6840 21664
rect 6748 21660 6795 21662
rect 7230 21660 7236 21724
rect 7300 21722 7347 21724
rect 7300 21720 7392 21722
rect 7342 21664 7392 21720
rect 7300 21662 7392 21664
rect 7300 21660 7347 21662
rect 7782 21660 7788 21724
rect 7852 21722 7899 21724
rect 7852 21720 7944 21722
rect 7894 21664 7944 21720
rect 7852 21662 7944 21664
rect 7852 21660 7899 21662
rect 8334 21660 8340 21724
rect 8404 21722 8451 21724
rect 8404 21720 8496 21722
rect 8446 21664 8496 21720
rect 8404 21662 8496 21664
rect 8404 21660 8451 21662
rect 9438 21660 9444 21724
rect 9508 21722 9555 21724
rect 9508 21720 9600 21722
rect 9550 21664 9600 21720
rect 9508 21662 9600 21664
rect 9508 21660 9555 21662
rect 9990 21660 9996 21724
rect 10060 21722 10107 21724
rect 10060 21720 10152 21722
rect 10102 21664 10152 21720
rect 10060 21662 10152 21664
rect 10060 21660 10107 21662
rect 10542 21660 10548 21724
rect 10612 21722 10659 21724
rect 10612 21720 10704 21722
rect 10654 21664 10704 21720
rect 10612 21662 10704 21664
rect 10612 21660 10659 21662
rect 11094 21660 11100 21724
rect 11164 21722 11211 21724
rect 11164 21720 11256 21722
rect 11206 21664 11256 21720
rect 11164 21662 11256 21664
rect 11164 21660 11211 21662
rect 12750 21660 12756 21724
rect 12820 21722 12867 21724
rect 12820 21720 12912 21722
rect 12862 21664 12912 21720
rect 12820 21662 12912 21664
rect 12820 21660 12867 21662
rect 13302 21660 13308 21724
rect 13372 21722 13419 21724
rect 13372 21720 13464 21722
rect 13414 21664 13464 21720
rect 13372 21662 13464 21664
rect 13372 21660 13419 21662
rect 13854 21660 13860 21724
rect 13924 21722 13971 21724
rect 13924 21720 14016 21722
rect 13966 21664 14016 21720
rect 13924 21662 14016 21664
rect 13924 21660 13971 21662
rect 16614 21660 16620 21724
rect 16684 21722 16731 21724
rect 16684 21720 16776 21722
rect 16726 21664 16776 21720
rect 16684 21662 16776 21664
rect 16684 21660 16731 21662
rect 6177 21659 6243 21660
rect 6729 21659 6795 21660
rect 7281 21659 7347 21660
rect 7833 21659 7899 21660
rect 8385 21659 8451 21660
rect 9489 21659 9555 21660
rect 10041 21659 10107 21660
rect 10593 21659 10659 21660
rect 11145 21659 11211 21660
rect 12801 21659 12867 21660
rect 13353 21659 13419 21660
rect 13905 21659 13971 21660
rect 16665 21659 16731 21660
rect 8150 21524 8156 21588
rect 8220 21586 8226 21588
rect 17174 21586 17234 21934
rect 24342 21932 24348 21934
rect 24412 21932 24418 21996
rect 19206 21792 19522 21793
rect 19206 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19522 21792
rect 19206 21727 19522 21728
rect 26980 21792 27296 21793
rect 26980 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27296 21792
rect 26980 21727 27296 21728
rect 8220 21526 17234 21586
rect 18094 21662 19074 21722
rect 8220 21524 8226 21526
rect 14365 21450 14431 21453
rect 18094 21450 18154 21662
rect 18413 21586 18479 21589
rect 18822 21586 18828 21588
rect 18413 21584 18828 21586
rect 18413 21528 18418 21584
rect 18474 21528 18828 21584
rect 18413 21526 18828 21528
rect 18413 21523 18479 21526
rect 18822 21524 18828 21526
rect 18892 21524 18898 21588
rect 19014 21586 19074 21662
rect 25814 21586 25820 21588
rect 19014 21526 25820 21586
rect 25814 21524 25820 21526
rect 25884 21524 25890 21588
rect 14365 21448 18154 21450
rect 14365 21392 14370 21448
rect 14426 21392 18154 21448
rect 14365 21390 18154 21392
rect 14365 21387 14431 21390
rect 18270 21388 18276 21452
rect 18340 21450 18346 21452
rect 21265 21450 21331 21453
rect 18340 21448 21331 21450
rect 18340 21392 21270 21448
rect 21326 21392 21331 21448
rect 18340 21390 21331 21392
rect 18340 21388 18346 21390
rect 21265 21387 21331 21390
rect 26233 21450 26299 21453
rect 26550 21450 26556 21452
rect 26233 21448 26556 21450
rect 26233 21392 26238 21448
rect 26294 21392 26556 21448
rect 26233 21390 26556 21392
rect 26233 21387 26299 21390
rect 26550 21388 26556 21390
rect 26620 21388 26626 21452
rect 28809 21450 28875 21453
rect 26742 21448 28875 21450
rect 26742 21392 28814 21448
rect 28870 21392 28875 21448
rect 26742 21390 28875 21392
rect 20897 21314 20963 21317
rect 21030 21314 21036 21316
rect 20897 21312 21036 21314
rect 20897 21256 20902 21312
rect 20958 21256 21036 21312
rect 20897 21254 21036 21256
rect 20897 21251 20963 21254
rect 21030 21252 21036 21254
rect 21100 21252 21106 21316
rect 23933 21314 23999 21317
rect 26742 21314 26802 21390
rect 28809 21387 28875 21390
rect 23933 21312 26802 21314
rect 23933 21256 23938 21312
rect 23994 21256 26802 21312
rect 23933 21254 26802 21256
rect 23933 21251 23999 21254
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 12092 21248 12408 21249
rect 12092 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12408 21248
rect 12092 21183 12408 21184
rect 19866 21248 20182 21249
rect 19866 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20182 21248
rect 19866 21183 20182 21184
rect 27640 21248 27956 21249
rect 27640 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27956 21248
rect 27640 21183 27956 21184
rect 16481 21178 16547 21181
rect 17166 21178 17172 21180
rect 16481 21176 17172 21178
rect 16481 21120 16486 21176
rect 16542 21120 17172 21176
rect 16481 21118 17172 21120
rect 16481 21115 16547 21118
rect 17166 21116 17172 21118
rect 17236 21116 17242 21180
rect 29269 21178 29335 21181
rect 30833 21178 30899 21181
rect 29269 21176 30899 21178
rect 29269 21120 29274 21176
rect 29330 21120 30838 21176
rect 30894 21120 30899 21176
rect 29269 21118 30899 21120
rect 29269 21115 29335 21118
rect 30833 21115 30899 21118
rect 15469 21044 15535 21045
rect 15469 21042 15516 21044
rect 15424 21040 15516 21042
rect 15424 20984 15474 21040
rect 15424 20982 15516 20984
rect 15469 20980 15516 20982
rect 15580 20980 15586 21044
rect 19057 21042 19123 21045
rect 27470 21042 27476 21044
rect 19057 21040 27476 21042
rect 19057 20984 19062 21040
rect 19118 20984 27476 21040
rect 19057 20982 27476 20984
rect 15469 20979 15535 20980
rect 19057 20979 19123 20982
rect 27470 20980 27476 20982
rect 27540 20980 27546 21044
rect 10409 20906 10475 20909
rect 24158 20906 24164 20908
rect 10409 20904 24164 20906
rect 10409 20848 10414 20904
rect 10470 20848 24164 20904
rect 10409 20846 24164 20848
rect 10409 20843 10475 20846
rect 24158 20844 24164 20846
rect 24228 20844 24234 20908
rect 28073 20906 28139 20909
rect 26742 20904 28139 20906
rect 26742 20848 28078 20904
rect 28134 20848 28139 20904
rect 26742 20846 28139 20848
rect 22829 20770 22895 20773
rect 26141 20770 26207 20773
rect 26742 20770 26802 20846
rect 28073 20843 28139 20846
rect 22829 20768 26802 20770
rect 22829 20712 22834 20768
rect 22890 20712 26146 20768
rect 26202 20712 26802 20768
rect 22829 20710 26802 20712
rect 22829 20707 22895 20710
rect 26141 20707 26207 20710
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 11432 20704 11748 20705
rect 11432 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11748 20704
rect 11432 20639 11748 20640
rect 19206 20704 19522 20705
rect 19206 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19522 20704
rect 19206 20639 19522 20640
rect 26980 20704 27296 20705
rect 26980 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27296 20704
rect 26980 20639 27296 20640
rect 14457 20636 14523 20637
rect 14406 20572 14412 20636
rect 14476 20634 14523 20636
rect 15193 20634 15259 20637
rect 16062 20634 16068 20636
rect 14476 20632 14568 20634
rect 14518 20576 14568 20632
rect 14476 20574 14568 20576
rect 15193 20632 16068 20634
rect 15193 20576 15198 20632
rect 15254 20576 16068 20632
rect 15193 20574 16068 20576
rect 14476 20572 14523 20574
rect 14457 20571 14523 20572
rect 15193 20571 15259 20574
rect 16062 20572 16068 20574
rect 16132 20572 16138 20636
rect 17718 20572 17724 20636
rect 17788 20634 17794 20636
rect 17953 20634 18019 20637
rect 17788 20632 18019 20634
rect 17788 20576 17958 20632
rect 18014 20576 18019 20632
rect 17788 20574 18019 20576
rect 17788 20572 17794 20574
rect 17953 20571 18019 20574
rect 974 20436 980 20500
rect 1044 20498 1050 20500
rect 12709 20498 12775 20501
rect 1044 20496 12775 20498
rect 1044 20440 12714 20496
rect 12770 20440 12775 20496
rect 1044 20438 12775 20440
rect 1044 20436 1050 20438
rect 12709 20435 12775 20438
rect 14825 20498 14891 20501
rect 26182 20498 26188 20500
rect 14825 20496 26188 20498
rect 14825 20440 14830 20496
rect 14886 20440 26188 20496
rect 14825 20438 26188 20440
rect 14825 20435 14891 20438
rect 26182 20436 26188 20438
rect 26252 20436 26258 20500
rect 27613 20498 27679 20501
rect 29821 20498 29887 20501
rect 26374 20496 29887 20498
rect 26374 20440 27618 20496
rect 27674 20440 29826 20496
rect 29882 20440 29887 20496
rect 26374 20438 29887 20440
rect 749 20362 815 20365
rect 7557 20362 7623 20365
rect 12801 20362 12867 20365
rect 22277 20362 22343 20365
rect 749 20360 7114 20362
rect 749 20304 754 20360
rect 810 20304 7114 20360
rect 749 20302 7114 20304
rect 749 20299 815 20302
rect 7054 20226 7114 20302
rect 7557 20360 12634 20362
rect 7557 20304 7562 20360
rect 7618 20304 12634 20360
rect 7557 20302 12634 20304
rect 7557 20299 7623 20302
rect 11145 20226 11211 20229
rect 7054 20224 11211 20226
rect 7054 20168 11150 20224
rect 11206 20168 11211 20224
rect 7054 20166 11211 20168
rect 12574 20226 12634 20302
rect 12801 20360 22343 20362
rect 12801 20304 12806 20360
rect 12862 20304 22282 20360
rect 22338 20304 22343 20360
rect 12801 20302 22343 20304
rect 12801 20299 12867 20302
rect 22277 20299 22343 20302
rect 24577 20362 24643 20365
rect 26374 20362 26434 20438
rect 27613 20435 27679 20438
rect 29821 20435 29887 20438
rect 24577 20360 26434 20362
rect 24577 20304 24582 20360
rect 24638 20304 26434 20360
rect 24577 20302 26434 20304
rect 26601 20362 26667 20365
rect 30833 20362 30899 20365
rect 31569 20362 31635 20365
rect 26601 20360 31635 20362
rect 26601 20304 26606 20360
rect 26662 20304 30838 20360
rect 30894 20304 31574 20360
rect 31630 20304 31635 20360
rect 26601 20302 31635 20304
rect 24577 20299 24643 20302
rect 26601 20299 26667 20302
rect 30833 20299 30899 20302
rect 31569 20299 31635 20302
rect 17953 20226 18019 20229
rect 12574 20224 18019 20226
rect 12574 20168 17958 20224
rect 18014 20168 18019 20224
rect 12574 20166 18019 20168
rect 11145 20163 11211 20166
rect 17953 20163 18019 20166
rect 20437 20226 20503 20229
rect 26417 20226 26483 20229
rect 20437 20224 26483 20226
rect 20437 20168 20442 20224
rect 20498 20168 26422 20224
rect 26478 20168 26483 20224
rect 20437 20166 26483 20168
rect 20437 20163 20503 20166
rect 26417 20163 26483 20166
rect 28901 20226 28967 20229
rect 29821 20226 29887 20229
rect 28901 20224 29887 20226
rect 28901 20168 28906 20224
rect 28962 20168 29826 20224
rect 29882 20168 29887 20224
rect 28901 20166 29887 20168
rect 28901 20163 28967 20166
rect 29821 20163 29887 20166
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 12092 20160 12408 20161
rect 12092 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12408 20160
rect 12092 20095 12408 20096
rect 19866 20160 20182 20161
rect 19866 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20182 20160
rect 19866 20095 20182 20096
rect 27640 20160 27956 20161
rect 27640 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27956 20160
rect 27640 20095 27956 20096
rect 7281 20090 7347 20093
rect 11881 20090 11947 20093
rect 7281 20088 11947 20090
rect 7281 20032 7286 20088
rect 7342 20032 11886 20088
rect 11942 20032 11947 20088
rect 7281 20030 11947 20032
rect 7281 20027 7347 20030
rect 11881 20027 11947 20030
rect 20345 20090 20411 20093
rect 21030 20090 21036 20092
rect 20345 20088 21036 20090
rect 20345 20032 20350 20088
rect 20406 20032 21036 20088
rect 20345 20030 21036 20032
rect 20345 20027 20411 20030
rect 21030 20028 21036 20030
rect 21100 20028 21106 20092
rect 26141 20090 26207 20093
rect 27153 20090 27219 20093
rect 26141 20088 27219 20090
rect 26141 20032 26146 20088
rect 26202 20032 27158 20088
rect 27214 20032 27219 20088
rect 26141 20030 27219 20032
rect 26141 20027 26207 20030
rect 27153 20027 27219 20030
rect 28165 20090 28231 20093
rect 29453 20090 29519 20093
rect 28165 20088 29519 20090
rect 28165 20032 28170 20088
rect 28226 20032 29458 20088
rect 29514 20032 29519 20088
rect 28165 20030 29519 20032
rect 28165 20027 28231 20030
rect 29453 20027 29519 20030
rect 2313 19954 2379 19957
rect 7557 19954 7623 19957
rect 15009 19956 15075 19957
rect 2313 19952 7623 19954
rect 2313 19896 2318 19952
rect 2374 19896 7562 19952
rect 7618 19896 7623 19952
rect 2313 19894 7623 19896
rect 2313 19891 2379 19894
rect 7557 19891 7623 19894
rect 14958 19892 14964 19956
rect 15028 19954 15075 19956
rect 15377 19954 15443 19957
rect 19149 19954 19215 19957
rect 25313 19954 25379 19957
rect 29545 19954 29611 19957
rect 15028 19952 15120 19954
rect 15070 19896 15120 19952
rect 15028 19894 15120 19896
rect 15377 19952 25146 19954
rect 15377 19896 15382 19952
rect 15438 19896 19154 19952
rect 19210 19896 25146 19952
rect 15377 19894 25146 19896
rect 15028 19892 15075 19894
rect 15009 19891 15075 19892
rect 15377 19891 15443 19894
rect 19149 19891 19215 19894
rect 10133 19818 10199 19821
rect 24710 19818 24716 19820
rect 10133 19816 24716 19818
rect 10133 19760 10138 19816
rect 10194 19760 24716 19816
rect 10133 19758 24716 19760
rect 10133 19755 10199 19758
rect 24710 19756 24716 19758
rect 24780 19756 24786 19820
rect 19609 19682 19675 19685
rect 23013 19682 23079 19685
rect 24577 19682 24643 19685
rect 11838 19622 17234 19682
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 11432 19616 11748 19617
rect 11432 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11748 19616
rect 11432 19551 11748 19552
rect 9673 19410 9739 19413
rect 11838 19410 11898 19622
rect 13261 19546 13327 19549
rect 13721 19546 13787 19549
rect 13261 19544 13787 19546
rect 13261 19488 13266 19544
rect 13322 19488 13726 19544
rect 13782 19488 13787 19544
rect 13261 19486 13787 19488
rect 13261 19483 13327 19486
rect 13721 19483 13787 19486
rect 15745 19546 15811 19549
rect 16849 19546 16915 19549
rect 15745 19544 16915 19546
rect 15745 19488 15750 19544
rect 15806 19488 16854 19544
rect 16910 19488 16915 19544
rect 15745 19486 16915 19488
rect 15745 19483 15811 19486
rect 16849 19483 16915 19486
rect 9673 19408 11898 19410
rect 9673 19352 9678 19408
rect 9734 19352 11898 19408
rect 9673 19350 11898 19352
rect 12065 19410 12131 19413
rect 16430 19410 16436 19412
rect 12065 19408 16436 19410
rect 12065 19352 12070 19408
rect 12126 19352 16436 19408
rect 12065 19350 16436 19352
rect 9673 19347 9739 19350
rect 12065 19347 12131 19350
rect 16430 19348 16436 19350
rect 16500 19348 16506 19412
rect 17174 19410 17234 19622
rect 19609 19680 24643 19682
rect 19609 19624 19614 19680
rect 19670 19624 23018 19680
rect 23074 19624 24582 19680
rect 24638 19624 24643 19680
rect 19609 19622 24643 19624
rect 25086 19682 25146 19894
rect 25313 19952 29611 19954
rect 25313 19896 25318 19952
rect 25374 19896 29550 19952
rect 29606 19896 29611 19952
rect 25313 19894 29611 19896
rect 25313 19891 25379 19894
rect 29545 19891 29611 19894
rect 25957 19818 26023 19821
rect 28993 19818 29059 19821
rect 25957 19816 29059 19818
rect 25957 19760 25962 19816
rect 26018 19760 28998 19816
rect 29054 19760 29059 19816
rect 25957 19758 29059 19760
rect 25957 19755 26023 19758
rect 28993 19755 29059 19758
rect 26325 19682 26391 19685
rect 26601 19682 26667 19685
rect 25086 19680 26667 19682
rect 25086 19624 26330 19680
rect 26386 19624 26606 19680
rect 26662 19624 26667 19680
rect 25086 19622 26667 19624
rect 19609 19619 19675 19622
rect 23013 19619 23079 19622
rect 24577 19619 24643 19622
rect 26325 19619 26391 19622
rect 26601 19619 26667 19622
rect 28533 19682 28599 19685
rect 31201 19682 31267 19685
rect 28533 19680 31267 19682
rect 28533 19624 28538 19680
rect 28594 19624 31206 19680
rect 31262 19624 31267 19680
rect 28533 19622 31267 19624
rect 28533 19619 28599 19622
rect 31201 19619 31267 19622
rect 19206 19616 19522 19617
rect 19206 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19522 19616
rect 19206 19551 19522 19552
rect 26980 19616 27296 19617
rect 26980 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27296 19616
rect 26980 19551 27296 19552
rect 22502 19546 22508 19548
rect 19750 19486 22508 19546
rect 19750 19410 19810 19486
rect 22502 19484 22508 19486
rect 22572 19484 22578 19548
rect 25998 19546 26004 19548
rect 25638 19486 26004 19546
rect 17174 19350 19810 19410
rect 19885 19410 19951 19413
rect 25638 19410 25698 19486
rect 25998 19484 26004 19486
rect 26068 19484 26074 19548
rect 19885 19408 25698 19410
rect 19885 19352 19890 19408
rect 19946 19352 25698 19408
rect 19885 19350 25698 19352
rect 25865 19410 25931 19413
rect 29729 19410 29795 19413
rect 25865 19408 29795 19410
rect 25865 19352 25870 19408
rect 25926 19352 29734 19408
rect 29790 19352 29795 19408
rect 25865 19350 29795 19352
rect 19885 19347 19951 19350
rect 25865 19347 25931 19350
rect 29729 19347 29795 19350
rect 9857 19274 9923 19277
rect 14038 19274 14044 19276
rect 9857 19272 14044 19274
rect 9857 19216 9862 19272
rect 9918 19216 14044 19272
rect 9857 19214 14044 19216
rect 9857 19211 9923 19214
rect 14038 19212 14044 19214
rect 14108 19212 14114 19276
rect 14365 19274 14431 19277
rect 20662 19274 20668 19276
rect 14365 19272 20668 19274
rect 14365 19216 14370 19272
rect 14426 19216 20668 19272
rect 14365 19214 20668 19216
rect 14365 19211 14431 19214
rect 20662 19212 20668 19214
rect 20732 19212 20738 19276
rect 21357 19274 21423 19277
rect 28758 19274 28764 19276
rect 21357 19272 28764 19274
rect 21357 19216 21362 19272
rect 21418 19216 28764 19272
rect 21357 19214 28764 19216
rect 21357 19211 21423 19214
rect 28758 19212 28764 19214
rect 28828 19212 28834 19276
rect 29453 19274 29519 19277
rect 30189 19274 30255 19277
rect 30925 19274 30991 19277
rect 29453 19272 30991 19274
rect 29453 19216 29458 19272
rect 29514 19216 30194 19272
rect 30250 19216 30930 19272
rect 30986 19216 30991 19272
rect 29453 19214 30991 19216
rect 29453 19211 29519 19214
rect 30189 19211 30255 19214
rect 30925 19211 30991 19214
rect 13077 19138 13143 19141
rect 13721 19138 13787 19141
rect 13077 19136 13787 19138
rect 13077 19080 13082 19136
rect 13138 19080 13726 19136
rect 13782 19080 13787 19136
rect 13077 19078 13787 19080
rect 13077 19075 13143 19078
rect 13721 19075 13787 19078
rect 21449 19138 21515 19141
rect 26141 19138 26207 19141
rect 21449 19136 26207 19138
rect 21449 19080 21454 19136
rect 21510 19080 26146 19136
rect 26202 19080 26207 19136
rect 21449 19078 26207 19080
rect 21449 19075 21515 19078
rect 26141 19075 26207 19078
rect 28717 19138 28783 19141
rect 29729 19138 29795 19141
rect 28717 19136 29795 19138
rect 28717 19080 28722 19136
rect 28778 19080 29734 19136
rect 29790 19080 29795 19136
rect 28717 19078 29795 19080
rect 28717 19075 28783 19078
rect 29729 19075 29795 19078
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12092 19072 12408 19073
rect 12092 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12408 19072
rect 12092 19007 12408 19008
rect 19866 19072 20182 19073
rect 19866 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20182 19072
rect 19866 19007 20182 19008
rect 27640 19072 27956 19073
rect 27640 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27956 19072
rect 27640 19007 27956 19008
rect 15101 19002 15167 19005
rect 20805 19002 20871 19005
rect 21633 19002 21699 19005
rect 13356 19000 15167 19002
rect 13356 18944 15106 19000
rect 15162 18944 15167 19000
rect 13356 18942 15167 18944
rect 6269 18866 6335 18869
rect 7005 18866 7071 18869
rect 6269 18864 7071 18866
rect 6269 18808 6274 18864
rect 6330 18808 7010 18864
rect 7066 18808 7071 18864
rect 6269 18806 7071 18808
rect 6269 18803 6335 18806
rect 7005 18803 7071 18806
rect 8385 18866 8451 18869
rect 13356 18866 13416 18942
rect 15101 18939 15167 18942
rect 20670 19000 21699 19002
rect 20670 18944 20810 19000
rect 20866 18944 21638 19000
rect 21694 18944 21699 19000
rect 20670 18942 21699 18944
rect 8385 18864 13416 18866
rect 8385 18808 8390 18864
rect 8446 18808 13416 18864
rect 8385 18806 13416 18808
rect 13537 18866 13603 18869
rect 20670 18866 20730 18942
rect 20805 18939 20871 18942
rect 21633 18939 21699 18942
rect 22921 19002 22987 19005
rect 26233 19002 26299 19005
rect 22921 19000 26299 19002
rect 22921 18944 22926 19000
rect 22982 18944 26238 19000
rect 26294 18944 26299 19000
rect 22921 18942 26299 18944
rect 22921 18939 22987 18942
rect 26233 18939 26299 18942
rect 13537 18864 20730 18866
rect 13537 18808 13542 18864
rect 13598 18808 20730 18864
rect 13537 18806 20730 18808
rect 20897 18866 20963 18869
rect 21541 18866 21607 18869
rect 20897 18864 21607 18866
rect 20897 18808 20902 18864
rect 20958 18808 21546 18864
rect 21602 18808 21607 18864
rect 20897 18806 21607 18808
rect 8385 18803 8451 18806
rect 13537 18803 13603 18806
rect 20897 18803 20963 18806
rect 21541 18803 21607 18806
rect 22185 18866 22251 18869
rect 23841 18866 23907 18869
rect 22185 18864 23907 18866
rect 22185 18808 22190 18864
rect 22246 18808 23846 18864
rect 23902 18808 23907 18864
rect 22185 18806 23907 18808
rect 22185 18803 22251 18806
rect 23841 18803 23907 18806
rect 24710 18804 24716 18868
rect 24780 18866 24786 18868
rect 25221 18866 25287 18869
rect 24780 18864 25287 18866
rect 24780 18808 25226 18864
rect 25282 18808 25287 18864
rect 24780 18806 25287 18808
rect 24780 18804 24786 18806
rect 25221 18803 25287 18806
rect 25405 18866 25471 18869
rect 29453 18866 29519 18869
rect 25405 18864 29519 18866
rect 25405 18808 25410 18864
rect 25466 18808 29458 18864
rect 29514 18808 29519 18864
rect 25405 18806 29519 18808
rect 25405 18803 25471 18806
rect 29453 18803 29519 18806
rect 3233 18730 3299 18733
rect 13721 18730 13787 18733
rect 25957 18730 26023 18733
rect 31477 18730 31543 18733
rect 3233 18728 13600 18730
rect 3233 18672 3238 18728
rect 3294 18672 13600 18728
rect 3233 18670 13600 18672
rect 3233 18667 3299 18670
rect 5758 18532 5764 18596
rect 5828 18594 5834 18596
rect 5901 18594 5967 18597
rect 6637 18596 6703 18597
rect 6637 18594 6684 18596
rect 5828 18592 5967 18594
rect 5828 18536 5906 18592
rect 5962 18536 5967 18592
rect 5828 18534 5967 18536
rect 6592 18592 6684 18594
rect 6592 18536 6642 18592
rect 6592 18534 6684 18536
rect 5828 18532 5834 18534
rect 5901 18531 5967 18534
rect 6637 18532 6684 18534
rect 6748 18532 6754 18596
rect 8293 18594 8359 18597
rect 9213 18594 9279 18597
rect 8293 18592 9279 18594
rect 8293 18536 8298 18592
rect 8354 18536 9218 18592
rect 9274 18536 9279 18592
rect 8293 18534 9279 18536
rect 13540 18594 13600 18670
rect 13721 18728 26023 18730
rect 13721 18672 13726 18728
rect 13782 18672 25962 18728
rect 26018 18672 26023 18728
rect 13721 18670 26023 18672
rect 13721 18667 13787 18670
rect 25957 18667 26023 18670
rect 26190 18728 31543 18730
rect 26190 18672 31482 18728
rect 31538 18672 31543 18728
rect 26190 18670 31543 18672
rect 18321 18594 18387 18597
rect 13540 18592 18387 18594
rect 13540 18536 18326 18592
rect 18382 18536 18387 18592
rect 13540 18534 18387 18536
rect 6637 18531 6703 18532
rect 8293 18531 8359 18534
rect 9213 18531 9279 18534
rect 18321 18531 18387 18534
rect 19885 18594 19951 18597
rect 20294 18594 20300 18596
rect 19885 18592 20300 18594
rect 19885 18536 19890 18592
rect 19946 18536 20300 18592
rect 19885 18534 20300 18536
rect 19885 18531 19951 18534
rect 20294 18532 20300 18534
rect 20364 18532 20370 18596
rect 22369 18594 22435 18597
rect 23013 18594 23079 18597
rect 26190 18594 26250 18670
rect 31477 18667 31543 18670
rect 22369 18592 26250 18594
rect 22369 18536 22374 18592
rect 22430 18536 23018 18592
rect 23074 18536 26250 18592
rect 22369 18534 26250 18536
rect 22369 18531 22435 18534
rect 23013 18531 23079 18534
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 11432 18528 11748 18529
rect 11432 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11748 18528
rect 11432 18463 11748 18464
rect 19206 18528 19522 18529
rect 19206 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19522 18528
rect 19206 18463 19522 18464
rect 26980 18528 27296 18529
rect 26980 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27296 18528
rect 26980 18463 27296 18464
rect 6177 18458 6243 18461
rect 9489 18458 9555 18461
rect 6177 18456 9555 18458
rect 6177 18400 6182 18456
rect 6238 18400 9494 18456
rect 9550 18400 9555 18456
rect 6177 18398 9555 18400
rect 6177 18395 6243 18398
rect 9489 18395 9555 18398
rect 11830 18396 11836 18460
rect 11900 18458 11906 18460
rect 14549 18458 14615 18461
rect 11900 18456 14615 18458
rect 11900 18400 14554 18456
rect 14610 18400 14615 18456
rect 11900 18398 14615 18400
rect 11900 18396 11906 18398
rect 14549 18395 14615 18398
rect 14733 18458 14799 18461
rect 18781 18458 18847 18461
rect 14733 18456 18847 18458
rect 14733 18400 14738 18456
rect 14794 18400 18786 18456
rect 18842 18400 18847 18456
rect 14733 18398 18847 18400
rect 14733 18395 14799 18398
rect 18781 18395 18847 18398
rect 21633 18458 21699 18461
rect 23933 18458 23999 18461
rect 21633 18456 23999 18458
rect 21633 18400 21638 18456
rect 21694 18400 23938 18456
rect 23994 18400 23999 18456
rect 21633 18398 23999 18400
rect 21633 18395 21699 18398
rect 23933 18395 23999 18398
rect 27705 18458 27771 18461
rect 29862 18458 29868 18460
rect 27705 18456 29868 18458
rect 27705 18400 27710 18456
rect 27766 18400 29868 18456
rect 27705 18398 29868 18400
rect 27705 18395 27771 18398
rect 29862 18396 29868 18398
rect 29932 18458 29938 18460
rect 30741 18458 30807 18461
rect 29932 18456 30807 18458
rect 29932 18400 30746 18456
rect 30802 18400 30807 18456
rect 29932 18398 30807 18400
rect 29932 18396 29938 18398
rect 30741 18395 30807 18398
rect 2630 18260 2636 18324
rect 2700 18322 2706 18324
rect 11237 18322 11303 18325
rect 18597 18322 18663 18325
rect 2700 18320 11303 18322
rect 2700 18264 11242 18320
rect 11298 18264 11303 18320
rect 2700 18262 11303 18264
rect 2700 18260 2706 18262
rect 11237 18259 11303 18262
rect 11516 18320 18663 18322
rect 11516 18264 18602 18320
rect 18658 18264 18663 18320
rect 11516 18262 18663 18264
rect 4102 18124 4108 18188
rect 4172 18186 4178 18188
rect 8569 18186 8635 18189
rect 4172 18184 8635 18186
rect 4172 18128 8574 18184
rect 8630 18128 8635 18184
rect 4172 18126 8635 18128
rect 4172 18124 4178 18126
rect 8569 18123 8635 18126
rect 8753 18186 8819 18189
rect 11516 18186 11576 18262
rect 18597 18259 18663 18262
rect 20069 18322 20135 18325
rect 23381 18322 23447 18325
rect 20069 18320 23447 18322
rect 20069 18264 20074 18320
rect 20130 18264 23386 18320
rect 23442 18264 23447 18320
rect 20069 18262 23447 18264
rect 20069 18259 20135 18262
rect 23381 18259 23447 18262
rect 23841 18322 23907 18325
rect 31293 18322 31359 18325
rect 23841 18320 31359 18322
rect 23841 18264 23846 18320
rect 23902 18264 31298 18320
rect 31354 18264 31359 18320
rect 23841 18262 31359 18264
rect 23841 18259 23907 18262
rect 31293 18259 31359 18262
rect 13629 18186 13695 18189
rect 21817 18186 21883 18189
rect 8753 18184 11576 18186
rect 8753 18128 8758 18184
rect 8814 18128 11576 18184
rect 8753 18126 11576 18128
rect 11654 18126 12588 18186
rect 8753 18123 8819 18126
rect 6085 18050 6151 18053
rect 6729 18050 6795 18053
rect 6085 18048 6795 18050
rect 6085 17992 6090 18048
rect 6146 17992 6734 18048
rect 6790 17992 6795 18048
rect 6085 17990 6795 17992
rect 6085 17987 6151 17990
rect 6729 17987 6795 17990
rect 8385 18050 8451 18053
rect 8845 18050 8911 18053
rect 10225 18052 10291 18053
rect 10174 18050 10180 18052
rect 8385 18048 8911 18050
rect 8385 17992 8390 18048
rect 8446 17992 8850 18048
rect 8906 17992 8911 18048
rect 8385 17990 8911 17992
rect 10134 17990 10180 18050
rect 10244 18048 10291 18052
rect 10286 17992 10291 18048
rect 8385 17987 8451 17990
rect 8845 17987 8911 17990
rect 10174 17988 10180 17990
rect 10244 17988 10291 17992
rect 10225 17987 10291 17988
rect 10593 18050 10659 18053
rect 11654 18050 11714 18126
rect 10593 18048 11714 18050
rect 10593 17992 10598 18048
rect 10654 17992 11714 18048
rect 10593 17990 11714 17992
rect 12528 18050 12588 18126
rect 13629 18184 17970 18186
rect 13629 18128 13634 18184
rect 13690 18128 17970 18184
rect 13629 18126 17970 18128
rect 13629 18123 13695 18126
rect 15510 18050 15516 18052
rect 12528 17990 15516 18050
rect 10593 17987 10659 17990
rect 15510 17988 15516 17990
rect 15580 17988 15586 18052
rect 17910 18050 17970 18126
rect 19382 18184 21883 18186
rect 19382 18128 21822 18184
rect 21878 18128 21883 18184
rect 19382 18126 21883 18128
rect 19382 18050 19442 18126
rect 21817 18123 21883 18126
rect 22461 18186 22527 18189
rect 26601 18186 26667 18189
rect 22461 18184 26667 18186
rect 22461 18128 22466 18184
rect 22522 18128 26606 18184
rect 26662 18128 26667 18184
rect 22461 18126 26667 18128
rect 22461 18123 22527 18126
rect 26601 18123 26667 18126
rect 26734 18124 26740 18188
rect 26804 18186 26810 18188
rect 27705 18186 27771 18189
rect 26804 18184 27771 18186
rect 26804 18128 27710 18184
rect 27766 18128 27771 18184
rect 26804 18126 27771 18128
rect 26804 18124 26810 18126
rect 27705 18123 27771 18126
rect 27889 18186 27955 18189
rect 28625 18186 28691 18189
rect 30465 18186 30531 18189
rect 30833 18186 30899 18189
rect 27889 18184 30899 18186
rect 27889 18128 27894 18184
rect 27950 18128 28630 18184
rect 28686 18128 30470 18184
rect 30526 18128 30838 18184
rect 30894 18128 30899 18184
rect 27889 18126 30899 18128
rect 27889 18123 27955 18126
rect 28625 18123 28691 18126
rect 30465 18123 30531 18126
rect 30833 18123 30899 18126
rect 17910 17990 19442 18050
rect 21950 17988 21956 18052
rect 22020 18050 22026 18052
rect 23473 18050 23539 18053
rect 22020 18048 23539 18050
rect 22020 17992 23478 18048
rect 23534 17992 23539 18048
rect 22020 17990 23539 17992
rect 22020 17988 22026 17990
rect 23473 17987 23539 17990
rect 28349 18050 28415 18053
rect 29729 18050 29795 18053
rect 28349 18048 29795 18050
rect 28349 17992 28354 18048
rect 28410 17992 29734 18048
rect 29790 17992 29795 18048
rect 28349 17990 29795 17992
rect 28349 17987 28415 17990
rect 29729 17987 29795 17990
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 12092 17984 12408 17985
rect 12092 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12408 17984
rect 12092 17919 12408 17920
rect 19866 17984 20182 17985
rect 19866 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20182 17984
rect 19866 17919 20182 17920
rect 27640 17984 27956 17985
rect 27640 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27956 17984
rect 27640 17919 27956 17920
rect 6310 17852 6316 17916
rect 6380 17914 6386 17916
rect 7557 17914 7623 17917
rect 6380 17912 7623 17914
rect 6380 17856 7562 17912
rect 7618 17856 7623 17912
rect 6380 17854 7623 17856
rect 6380 17852 6386 17854
rect 7557 17851 7623 17854
rect 7925 17914 7991 17917
rect 8845 17914 8911 17917
rect 7925 17912 8911 17914
rect 7925 17856 7930 17912
rect 7986 17856 8850 17912
rect 8906 17856 8911 17912
rect 7925 17854 8911 17856
rect 7925 17851 7991 17854
rect 8845 17851 8911 17854
rect 11094 17852 11100 17916
rect 11164 17914 11170 17916
rect 11830 17914 11836 17916
rect 11164 17854 11836 17914
rect 11164 17852 11170 17854
rect 11830 17852 11836 17854
rect 11900 17852 11906 17916
rect 12525 17914 12591 17917
rect 12985 17914 13051 17917
rect 19701 17914 19767 17917
rect 12525 17912 12818 17914
rect 12525 17856 12530 17912
rect 12586 17856 12818 17912
rect 12525 17854 12818 17856
rect 12525 17851 12591 17854
rect 2221 17778 2287 17781
rect 12617 17778 12683 17781
rect 2221 17776 12683 17778
rect 2221 17720 2226 17776
rect 2282 17720 12622 17776
rect 12678 17720 12683 17776
rect 2221 17718 12683 17720
rect 12758 17778 12818 17854
rect 12985 17912 19767 17914
rect 12985 17856 12990 17912
rect 13046 17856 19706 17912
rect 19762 17856 19767 17912
rect 12985 17854 19767 17856
rect 12985 17851 13051 17854
rect 19701 17851 19767 17854
rect 20253 17914 20319 17917
rect 20713 17914 20779 17917
rect 20253 17912 20779 17914
rect 20253 17856 20258 17912
rect 20314 17856 20718 17912
rect 20774 17856 20779 17912
rect 20253 17854 20779 17856
rect 20253 17851 20319 17854
rect 20713 17851 20779 17854
rect 22001 17914 22067 17917
rect 25497 17914 25563 17917
rect 22001 17912 25563 17914
rect 22001 17856 22006 17912
rect 22062 17856 25502 17912
rect 25558 17856 25563 17912
rect 22001 17854 25563 17856
rect 22001 17851 22067 17854
rect 25497 17851 25563 17854
rect 25998 17852 26004 17916
rect 26068 17914 26074 17916
rect 26233 17914 26299 17917
rect 26068 17912 26299 17914
rect 26068 17856 26238 17912
rect 26294 17856 26299 17912
rect 26068 17854 26299 17856
rect 26068 17852 26074 17854
rect 26233 17851 26299 17854
rect 14825 17778 14891 17781
rect 12758 17776 14891 17778
rect 12758 17720 14830 17776
rect 14886 17720 14891 17776
rect 12758 17718 14891 17720
rect 2221 17715 2287 17718
rect 12617 17715 12683 17718
rect 14825 17715 14891 17718
rect 18597 17778 18663 17781
rect 23197 17778 23263 17781
rect 18597 17776 23263 17778
rect 18597 17720 18602 17776
rect 18658 17720 23202 17776
rect 23258 17720 23263 17776
rect 18597 17718 23263 17720
rect 18597 17715 18663 17718
rect 23197 17715 23263 17718
rect 23381 17778 23447 17781
rect 24393 17778 24459 17781
rect 23381 17776 24459 17778
rect 23381 17720 23386 17776
rect 23442 17720 24398 17776
rect 24454 17720 24459 17776
rect 23381 17718 24459 17720
rect 23381 17715 23447 17718
rect 24393 17715 24459 17718
rect 25405 17778 25471 17781
rect 28390 17778 28396 17780
rect 25405 17776 28396 17778
rect 25405 17720 25410 17776
rect 25466 17720 28396 17776
rect 25405 17718 28396 17720
rect 25405 17715 25471 17718
rect 28390 17716 28396 17718
rect 28460 17716 28466 17780
rect 1945 17642 2011 17645
rect 6913 17642 6979 17645
rect 1945 17640 6979 17642
rect 1945 17584 1950 17640
rect 2006 17584 6918 17640
rect 6974 17584 6979 17640
rect 1945 17582 6979 17584
rect 1945 17579 2011 17582
rect 6913 17579 6979 17582
rect 8201 17642 8267 17645
rect 8886 17642 8892 17644
rect 8201 17640 8892 17642
rect 8201 17584 8206 17640
rect 8262 17584 8892 17640
rect 8201 17582 8892 17584
rect 8201 17579 8267 17582
rect 8886 17580 8892 17582
rect 8956 17580 8962 17644
rect 9213 17642 9279 17645
rect 13854 17642 13860 17644
rect 9213 17640 13860 17642
rect 9213 17584 9218 17640
rect 9274 17584 13860 17640
rect 9213 17582 13860 17584
rect 8894 17506 8954 17580
rect 9213 17579 9279 17582
rect 13854 17580 13860 17582
rect 13924 17580 13930 17644
rect 14038 17580 14044 17644
rect 14108 17642 14114 17644
rect 14273 17642 14339 17645
rect 15837 17642 15903 17645
rect 21081 17642 21147 17645
rect 14108 17640 15903 17642
rect 14108 17584 14278 17640
rect 14334 17584 15842 17640
rect 15898 17584 15903 17640
rect 14108 17582 15903 17584
rect 14108 17580 14114 17582
rect 14273 17579 14339 17582
rect 15837 17579 15903 17582
rect 18600 17640 21147 17642
rect 18600 17584 21086 17640
rect 21142 17584 21147 17640
rect 18600 17582 21147 17584
rect 11237 17506 11303 17509
rect 8894 17504 11303 17506
rect 8894 17448 11242 17504
rect 11298 17448 11303 17504
rect 8894 17446 11303 17448
rect 11237 17443 11303 17446
rect 11830 17444 11836 17508
rect 11900 17506 11906 17508
rect 12341 17506 12407 17509
rect 11900 17504 12407 17506
rect 11900 17448 12346 17504
rect 12402 17448 12407 17504
rect 11900 17446 12407 17448
rect 11900 17444 11906 17446
rect 12341 17443 12407 17446
rect 12525 17506 12591 17509
rect 12934 17506 12940 17508
rect 12525 17504 12940 17506
rect 12525 17448 12530 17504
rect 12586 17448 12940 17504
rect 12525 17446 12940 17448
rect 12525 17443 12591 17446
rect 12934 17444 12940 17446
rect 13004 17444 13010 17508
rect 13997 17506 14063 17509
rect 14406 17506 14412 17508
rect 13997 17504 14412 17506
rect 13997 17448 14002 17504
rect 14058 17448 14412 17504
rect 13997 17446 14412 17448
rect 13997 17443 14063 17446
rect 14406 17444 14412 17446
rect 14476 17444 14482 17508
rect 17125 17506 17191 17509
rect 18600 17506 18660 17582
rect 21081 17579 21147 17582
rect 21541 17642 21607 17645
rect 25313 17642 25379 17645
rect 21541 17640 25379 17642
rect 21541 17584 21546 17640
rect 21602 17584 25318 17640
rect 25374 17584 25379 17640
rect 21541 17582 25379 17584
rect 21541 17579 21607 17582
rect 25313 17579 25379 17582
rect 25957 17642 26023 17645
rect 30373 17642 30439 17645
rect 31109 17642 31175 17645
rect 25957 17640 31175 17642
rect 25957 17584 25962 17640
rect 26018 17584 30378 17640
rect 30434 17584 31114 17640
rect 31170 17584 31175 17640
rect 25957 17582 31175 17584
rect 25957 17579 26023 17582
rect 30373 17579 30439 17582
rect 31109 17579 31175 17582
rect 25221 17506 25287 17509
rect 17125 17504 18660 17506
rect 17125 17448 17130 17504
rect 17186 17448 18660 17504
rect 17125 17446 18660 17448
rect 20716 17504 25287 17506
rect 20716 17448 25226 17504
rect 25282 17448 25287 17504
rect 20716 17446 25287 17448
rect 17125 17443 17191 17446
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 11432 17440 11748 17441
rect 11432 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11748 17440
rect 11432 17375 11748 17376
rect 19206 17440 19522 17441
rect 19206 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19522 17440
rect 19206 17375 19522 17376
rect 4337 17370 4403 17373
rect 4797 17370 4863 17373
rect 7097 17370 7163 17373
rect 4337 17368 7163 17370
rect 4337 17312 4342 17368
rect 4398 17312 4802 17368
rect 4858 17312 7102 17368
rect 7158 17312 7163 17368
rect 4337 17310 7163 17312
rect 4337 17307 4403 17310
rect 4797 17307 4863 17310
rect 7097 17307 7163 17310
rect 8477 17370 8543 17373
rect 9305 17370 9371 17373
rect 8477 17368 9371 17370
rect 8477 17312 8482 17368
rect 8538 17312 9310 17368
rect 9366 17312 9371 17368
rect 8477 17310 9371 17312
rect 8477 17307 8543 17310
rect 9305 17307 9371 17310
rect 10409 17370 10475 17373
rect 10542 17370 10548 17372
rect 10409 17368 10548 17370
rect 10409 17312 10414 17368
rect 10470 17312 10548 17368
rect 10409 17310 10548 17312
rect 10409 17307 10475 17310
rect 10542 17308 10548 17310
rect 10612 17308 10618 17372
rect 12433 17370 12499 17373
rect 13813 17370 13879 17373
rect 12433 17368 13879 17370
rect 12433 17312 12438 17368
rect 12494 17312 13818 17368
rect 13874 17312 13879 17368
rect 12433 17310 13879 17312
rect 12433 17307 12499 17310
rect 13813 17307 13879 17310
rect 6913 17234 6979 17237
rect 12801 17234 12867 17237
rect 6913 17232 12867 17234
rect 6913 17176 6918 17232
rect 6974 17176 12806 17232
rect 12862 17176 12867 17232
rect 6913 17174 12867 17176
rect 6913 17171 6979 17174
rect 12801 17171 12867 17174
rect 13721 17234 13787 17237
rect 14038 17234 14044 17236
rect 13721 17232 14044 17234
rect 13721 17176 13726 17232
rect 13782 17176 14044 17232
rect 13721 17174 14044 17176
rect 13721 17171 13787 17174
rect 14038 17172 14044 17174
rect 14108 17172 14114 17236
rect 20716 17234 20776 17446
rect 25221 17443 25287 17446
rect 25814 17444 25820 17508
rect 25884 17506 25890 17508
rect 25957 17506 26023 17509
rect 25884 17504 26023 17506
rect 25884 17448 25962 17504
rect 26018 17448 26023 17504
rect 25884 17446 26023 17448
rect 25884 17444 25890 17446
rect 25957 17443 26023 17446
rect 27889 17506 27955 17509
rect 28165 17506 28231 17509
rect 31661 17506 31727 17509
rect 27889 17504 31727 17506
rect 27889 17448 27894 17504
rect 27950 17448 28170 17504
rect 28226 17448 31666 17504
rect 31722 17448 31727 17504
rect 27889 17446 31727 17448
rect 27889 17443 27955 17446
rect 28165 17443 28231 17446
rect 31661 17443 31727 17446
rect 26980 17440 27296 17441
rect 26980 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27296 17440
rect 26980 17375 27296 17376
rect 21817 17370 21883 17373
rect 26417 17370 26483 17373
rect 21817 17368 26483 17370
rect 21817 17312 21822 17368
rect 21878 17312 26422 17368
rect 26478 17312 26483 17368
rect 21817 17310 26483 17312
rect 21817 17307 21883 17310
rect 26417 17307 26483 17310
rect 27521 17370 27587 17373
rect 28022 17370 28028 17372
rect 27521 17368 28028 17370
rect 27521 17312 27526 17368
rect 27582 17312 28028 17368
rect 27521 17310 28028 17312
rect 27521 17307 27587 17310
rect 28022 17308 28028 17310
rect 28092 17308 28098 17372
rect 28441 17370 28507 17373
rect 29545 17370 29611 17373
rect 28441 17368 29611 17370
rect 28441 17312 28446 17368
rect 28502 17312 29550 17368
rect 29606 17312 29611 17368
rect 28441 17310 29611 17312
rect 28441 17307 28507 17310
rect 29545 17307 29611 17310
rect 23105 17234 23171 17237
rect 14184 17174 20776 17234
rect 20854 17232 23171 17234
rect 20854 17176 23110 17232
rect 23166 17176 23171 17232
rect 20854 17174 23171 17176
rect 3325 17098 3391 17101
rect 3509 17098 3575 17101
rect 5809 17098 5875 17101
rect 6361 17098 6427 17101
rect 11094 17098 11100 17100
rect 3325 17096 4860 17098
rect 3325 17040 3330 17096
rect 3386 17040 3514 17096
rect 3570 17040 4860 17096
rect 3325 17038 4860 17040
rect 3325 17035 3391 17038
rect 3509 17035 3575 17038
rect 4800 16962 4860 17038
rect 5809 17096 11100 17098
rect 5809 17040 5814 17096
rect 5870 17040 6366 17096
rect 6422 17040 11100 17096
rect 5809 17038 11100 17040
rect 5809 17035 5875 17038
rect 6361 17035 6427 17038
rect 11094 17036 11100 17038
rect 11164 17036 11170 17100
rect 12525 17098 12591 17101
rect 11240 17096 12591 17098
rect 11240 17040 12530 17096
rect 12586 17040 12591 17096
rect 11240 17038 12591 17040
rect 11240 16962 11300 17038
rect 12525 17035 12591 17038
rect 13721 17098 13787 17101
rect 14184 17098 14244 17174
rect 13721 17096 14244 17098
rect 13721 17040 13726 17096
rect 13782 17040 14244 17096
rect 13721 17038 14244 17040
rect 17033 17098 17099 17101
rect 19977 17098 20043 17101
rect 20621 17098 20687 17101
rect 17033 17096 20687 17098
rect 17033 17040 17038 17096
rect 17094 17040 19982 17096
rect 20038 17040 20626 17096
rect 20682 17040 20687 17096
rect 17033 17038 20687 17040
rect 13721 17035 13787 17038
rect 17033 17035 17099 17038
rect 19977 17035 20043 17038
rect 20621 17035 20687 17038
rect 12709 16964 12775 16965
rect 12709 16962 12756 16964
rect 4800 16902 11300 16962
rect 12664 16960 12756 16962
rect 12664 16904 12714 16960
rect 12664 16902 12756 16904
rect 12709 16900 12756 16902
rect 12820 16900 12826 16964
rect 15142 16962 15148 16964
rect 13678 16902 15148 16962
rect 12709 16899 12775 16900
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 12092 16896 12408 16897
rect 12092 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12408 16896
rect 12092 16831 12408 16832
rect 7649 16826 7715 16829
rect 8937 16826 9003 16829
rect 10869 16828 10935 16829
rect 10869 16826 10916 16828
rect 7649 16824 9003 16826
rect 7649 16768 7654 16824
rect 7710 16768 8942 16824
rect 8998 16768 9003 16824
rect 7649 16766 9003 16768
rect 10824 16824 10916 16826
rect 10824 16768 10874 16824
rect 10824 16766 10916 16768
rect 7649 16763 7715 16766
rect 8937 16763 9003 16766
rect 10869 16764 10916 16766
rect 10980 16764 10986 16828
rect 11145 16826 11211 16829
rect 11830 16826 11836 16828
rect 11145 16824 11836 16826
rect 11145 16768 11150 16824
rect 11206 16768 11836 16824
rect 11145 16766 11836 16768
rect 10869 16763 10935 16764
rect 11145 16763 11211 16766
rect 11830 16764 11836 16766
rect 11900 16764 11906 16828
rect 12709 16826 12775 16829
rect 13537 16826 13603 16829
rect 12709 16824 13603 16826
rect 12709 16768 12714 16824
rect 12770 16768 13542 16824
rect 13598 16768 13603 16824
rect 12709 16766 13603 16768
rect 12709 16763 12775 16766
rect 13537 16763 13603 16766
rect 4981 16690 5047 16693
rect 5206 16690 5212 16692
rect 4981 16688 5212 16690
rect 4981 16632 4986 16688
rect 5042 16632 5212 16688
rect 4981 16630 5212 16632
rect 4981 16627 5047 16630
rect 5206 16628 5212 16630
rect 5276 16628 5282 16692
rect 8201 16690 8267 16693
rect 13678 16690 13738 16902
rect 15142 16900 15148 16902
rect 15212 16962 15218 16964
rect 18045 16962 18111 16965
rect 15212 16960 18111 16962
rect 15212 16904 18050 16960
rect 18106 16904 18111 16960
rect 15212 16902 18111 16904
rect 15212 16900 15218 16902
rect 18045 16899 18111 16902
rect 19866 16896 20182 16897
rect 19866 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20182 16896
rect 19866 16831 20182 16832
rect 13813 16826 13879 16829
rect 14549 16826 14615 16829
rect 18321 16826 18387 16829
rect 18638 16826 18644 16828
rect 13813 16824 17786 16826
rect 13813 16768 13818 16824
rect 13874 16768 14554 16824
rect 14610 16768 17786 16824
rect 13813 16766 17786 16768
rect 13813 16763 13879 16766
rect 14549 16763 14615 16766
rect 8201 16688 13738 16690
rect 8201 16632 8206 16688
rect 8262 16632 13738 16688
rect 8201 16630 13738 16632
rect 15009 16690 15075 16693
rect 15326 16690 15332 16692
rect 15009 16688 15332 16690
rect 15009 16632 15014 16688
rect 15070 16632 15332 16688
rect 15009 16630 15332 16632
rect 8201 16627 8267 16630
rect 15009 16627 15075 16630
rect 15326 16628 15332 16630
rect 15396 16628 15402 16692
rect 15878 16628 15884 16692
rect 15948 16690 15954 16692
rect 16021 16690 16087 16693
rect 15948 16688 16087 16690
rect 15948 16632 16026 16688
rect 16082 16632 16087 16688
rect 15948 16630 16087 16632
rect 15948 16628 15954 16630
rect 16021 16627 16087 16630
rect 16246 16628 16252 16692
rect 16316 16690 16322 16692
rect 16389 16690 16455 16693
rect 16316 16688 16455 16690
rect 16316 16632 16394 16688
rect 16450 16632 16455 16688
rect 16316 16630 16455 16632
rect 16316 16628 16322 16630
rect 16389 16627 16455 16630
rect 16798 16628 16804 16692
rect 16868 16690 16874 16692
rect 17493 16690 17559 16693
rect 16868 16688 17559 16690
rect 16868 16632 17498 16688
rect 17554 16632 17559 16688
rect 16868 16630 17559 16632
rect 17726 16690 17786 16766
rect 18321 16824 18644 16826
rect 18321 16768 18326 16824
rect 18382 16768 18644 16824
rect 18321 16766 18644 16768
rect 18321 16763 18387 16766
rect 18638 16764 18644 16766
rect 18708 16764 18714 16828
rect 20854 16826 20914 17174
rect 23105 17171 23171 17174
rect 23381 17234 23447 17237
rect 24761 17234 24827 17237
rect 26141 17234 26207 17237
rect 23381 17232 24827 17234
rect 23381 17176 23386 17232
rect 23442 17176 24766 17232
rect 24822 17176 24827 17232
rect 23381 17174 24827 17176
rect 23381 17171 23447 17174
rect 24761 17171 24827 17174
rect 24902 17232 26207 17234
rect 24902 17176 26146 17232
rect 26202 17176 26207 17232
rect 24902 17174 26207 17176
rect 21081 17098 21147 17101
rect 22369 17098 22435 17101
rect 22737 17100 22803 17101
rect 22686 17098 22692 17100
rect 21081 17096 22435 17098
rect 21081 17040 21086 17096
rect 21142 17040 22374 17096
rect 22430 17040 22435 17096
rect 21081 17038 22435 17040
rect 22610 17038 22692 17098
rect 22756 17098 22803 17100
rect 24902 17098 24962 17174
rect 26141 17171 26207 17174
rect 26325 17234 26391 17237
rect 28073 17234 28139 17237
rect 29453 17234 29519 17237
rect 26325 17232 29519 17234
rect 26325 17176 26330 17232
rect 26386 17176 28078 17232
rect 28134 17176 29458 17232
rect 29514 17176 29519 17232
rect 26325 17174 29519 17176
rect 26325 17171 26391 17174
rect 28073 17171 28139 17174
rect 29453 17171 29519 17174
rect 22756 17096 24962 17098
rect 22798 17040 24962 17096
rect 21081 17035 21147 17038
rect 22369 17035 22435 17038
rect 22686 17036 22692 17038
rect 22756 17038 24962 17040
rect 25589 17098 25655 17101
rect 28993 17098 29059 17101
rect 25589 17096 29059 17098
rect 25589 17040 25594 17096
rect 25650 17040 28998 17096
rect 29054 17040 29059 17096
rect 25589 17038 29059 17040
rect 22756 17036 22803 17038
rect 22737 17035 22803 17036
rect 25589 17035 25655 17038
rect 28993 17035 29059 17038
rect 29269 17098 29335 17101
rect 29494 17098 29500 17100
rect 29269 17096 29500 17098
rect 29269 17040 29274 17096
rect 29330 17040 29500 17096
rect 29269 17038 29500 17040
rect 29269 17035 29335 17038
rect 29494 17036 29500 17038
rect 29564 17036 29570 17100
rect 21081 16962 21147 16965
rect 23105 16962 23171 16965
rect 27337 16962 27403 16965
rect 21081 16960 22524 16962
rect 21081 16904 21086 16960
rect 21142 16904 22524 16960
rect 21081 16902 22524 16904
rect 21081 16899 21147 16902
rect 20302 16766 20914 16826
rect 22093 16826 22159 16829
rect 22318 16826 22324 16828
rect 22093 16824 22324 16826
rect 22093 16768 22098 16824
rect 22154 16768 22324 16824
rect 22093 16766 22324 16768
rect 20302 16690 20362 16766
rect 22093 16763 22159 16766
rect 22318 16764 22324 16766
rect 22388 16764 22394 16828
rect 22464 16826 22524 16902
rect 23105 16960 27403 16962
rect 23105 16904 23110 16960
rect 23166 16904 27342 16960
rect 27398 16904 27403 16960
rect 23105 16902 27403 16904
rect 23105 16899 23171 16902
rect 27337 16899 27403 16902
rect 28073 16962 28139 16965
rect 28625 16962 28691 16965
rect 28073 16960 28691 16962
rect 28073 16904 28078 16960
rect 28134 16904 28630 16960
rect 28686 16904 28691 16960
rect 28073 16902 28691 16904
rect 28073 16899 28139 16902
rect 28625 16899 28691 16902
rect 27640 16896 27956 16897
rect 27640 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27956 16896
rect 27640 16831 27956 16832
rect 23657 16826 23723 16829
rect 22464 16824 23723 16826
rect 22464 16768 23662 16824
rect 23718 16768 23723 16824
rect 22464 16766 23723 16768
rect 23657 16763 23723 16766
rect 24485 16826 24551 16829
rect 25405 16826 25471 16829
rect 26325 16826 26391 16829
rect 28901 16826 28967 16829
rect 24485 16824 26391 16826
rect 24485 16768 24490 16824
rect 24546 16768 25410 16824
rect 25466 16768 26330 16824
rect 26386 16768 26391 16824
rect 24485 16766 26391 16768
rect 24485 16763 24551 16766
rect 25405 16763 25471 16766
rect 26325 16763 26391 16766
rect 28076 16824 28967 16826
rect 28076 16768 28906 16824
rect 28962 16768 28967 16824
rect 28076 16766 28967 16768
rect 28076 16693 28136 16766
rect 28901 16763 28967 16766
rect 17726 16630 20362 16690
rect 20897 16690 20963 16693
rect 22185 16690 22251 16693
rect 20897 16688 22251 16690
rect 20897 16632 20902 16688
rect 20958 16632 22190 16688
rect 22246 16632 22251 16688
rect 20897 16630 22251 16632
rect 16868 16628 16874 16630
rect 17493 16627 17559 16630
rect 20897 16627 20963 16630
rect 22185 16627 22251 16630
rect 22829 16690 22895 16693
rect 24853 16690 24919 16693
rect 26325 16690 26391 16693
rect 22829 16688 24919 16690
rect 22829 16632 22834 16688
rect 22890 16632 24858 16688
rect 24914 16632 24919 16688
rect 22829 16630 24919 16632
rect 22829 16627 22895 16630
rect 24853 16627 24919 16630
rect 25132 16688 26391 16690
rect 25132 16632 26330 16688
rect 26386 16632 26391 16688
rect 25132 16630 26391 16632
rect 4797 16554 4863 16557
rect 13813 16554 13879 16557
rect 4797 16552 13879 16554
rect 4797 16496 4802 16552
rect 4858 16496 13818 16552
rect 13874 16496 13879 16552
rect 4797 16494 13879 16496
rect 4797 16491 4863 16494
rect 13813 16491 13879 16494
rect 14590 16492 14596 16556
rect 14660 16554 14666 16556
rect 15929 16554 15995 16557
rect 21817 16554 21883 16557
rect 22093 16556 22159 16557
rect 22093 16554 22140 16556
rect 14660 16552 21883 16554
rect 14660 16496 15934 16552
rect 15990 16496 21822 16552
rect 21878 16496 21883 16552
rect 14660 16494 21883 16496
rect 22048 16552 22140 16554
rect 22048 16496 22098 16552
rect 22048 16494 22140 16496
rect 14660 16492 14666 16494
rect 15929 16491 15995 16494
rect 21817 16491 21883 16494
rect 22093 16492 22140 16494
rect 22204 16492 22210 16556
rect 22502 16492 22508 16556
rect 22572 16554 22578 16556
rect 22921 16554 22987 16557
rect 22572 16552 22987 16554
rect 22572 16496 22926 16552
rect 22982 16496 22987 16552
rect 22572 16494 22987 16496
rect 22572 16492 22578 16494
rect 22093 16491 22159 16492
rect 22921 16491 22987 16494
rect 23197 16554 23263 16557
rect 25132 16554 25192 16630
rect 26325 16627 26391 16630
rect 26877 16690 26943 16693
rect 28073 16690 28139 16693
rect 26877 16688 28139 16690
rect 26877 16632 26882 16688
rect 26938 16632 28078 16688
rect 28134 16632 28139 16688
rect 26877 16630 28139 16632
rect 26877 16627 26943 16630
rect 28073 16627 28139 16630
rect 28390 16628 28396 16692
rect 28460 16690 28466 16692
rect 28901 16690 28967 16693
rect 31109 16690 31175 16693
rect 28460 16688 31175 16690
rect 28460 16632 28906 16688
rect 28962 16632 31114 16688
rect 31170 16632 31175 16688
rect 28460 16630 31175 16632
rect 28460 16628 28466 16630
rect 28901 16627 28967 16630
rect 31109 16627 31175 16630
rect 26233 16556 26299 16557
rect 26182 16554 26188 16556
rect 23197 16552 25192 16554
rect 23197 16496 23202 16552
rect 23258 16496 25192 16552
rect 23197 16494 25192 16496
rect 26142 16494 26188 16554
rect 26252 16552 26299 16556
rect 26294 16496 26299 16552
rect 23197 16491 23263 16494
rect 26182 16492 26188 16494
rect 26252 16492 26299 16496
rect 26233 16491 26299 16492
rect 26417 16554 26483 16557
rect 28349 16554 28415 16557
rect 26417 16552 28415 16554
rect 26417 16496 26422 16552
rect 26478 16496 28354 16552
rect 28410 16496 28415 16552
rect 26417 16494 28415 16496
rect 26417 16491 26483 16494
rect 28349 16491 28415 16494
rect 29269 16556 29335 16557
rect 29269 16552 29316 16556
rect 29380 16554 29386 16556
rect 29269 16496 29274 16552
rect 29269 16492 29316 16496
rect 29380 16494 29426 16554
rect 29380 16492 29386 16494
rect 29269 16491 29335 16492
rect 11881 16418 11947 16421
rect 17493 16418 17559 16421
rect 11881 16416 17559 16418
rect 11881 16360 11886 16416
rect 11942 16360 17498 16416
rect 17554 16360 17559 16416
rect 11881 16358 17559 16360
rect 11881 16355 11947 16358
rect 17493 16355 17559 16358
rect 19701 16418 19767 16421
rect 21725 16418 21791 16421
rect 25681 16418 25747 16421
rect 19701 16416 21791 16418
rect 19701 16360 19706 16416
rect 19762 16360 21730 16416
rect 21786 16360 21791 16416
rect 19701 16358 21791 16360
rect 19701 16355 19767 16358
rect 21725 16355 21791 16358
rect 22188 16416 25747 16418
rect 22188 16360 25686 16416
rect 25742 16360 25747 16416
rect 22188 16358 25747 16360
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 11432 16352 11748 16353
rect 11432 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11748 16352
rect 11432 16287 11748 16288
rect 19206 16352 19522 16353
rect 19206 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19522 16352
rect 19206 16287 19522 16288
rect 7230 16220 7236 16284
rect 7300 16282 7306 16284
rect 7649 16282 7715 16285
rect 7300 16280 7715 16282
rect 7300 16224 7654 16280
rect 7710 16224 7715 16280
rect 7300 16222 7715 16224
rect 7300 16220 7306 16222
rect 7649 16219 7715 16222
rect 8477 16282 8543 16285
rect 10542 16282 10548 16284
rect 8477 16280 10548 16282
rect 8477 16224 8482 16280
rect 8538 16224 10548 16280
rect 8477 16222 10548 16224
rect 8477 16219 8543 16222
rect 10542 16220 10548 16222
rect 10612 16282 10618 16284
rect 10961 16282 11027 16285
rect 12341 16282 12407 16285
rect 10612 16280 11027 16282
rect 10612 16224 10966 16280
rect 11022 16224 11027 16280
rect 10612 16222 11027 16224
rect 10612 16220 10618 16222
rect 10961 16219 11027 16222
rect 12022 16280 12407 16282
rect 12022 16224 12346 16280
rect 12402 16224 12407 16280
rect 12022 16222 12407 16224
rect 7281 16146 7347 16149
rect 7414 16146 7420 16148
rect 7281 16144 7420 16146
rect 7281 16088 7286 16144
rect 7342 16088 7420 16144
rect 7281 16086 7420 16088
rect 7281 16083 7347 16086
rect 7414 16084 7420 16086
rect 7484 16084 7490 16148
rect 10225 16146 10291 16149
rect 12022 16146 12082 16222
rect 12341 16219 12407 16222
rect 12525 16282 12591 16285
rect 16665 16282 16731 16285
rect 12525 16280 16731 16282
rect 12525 16224 12530 16280
rect 12586 16224 16670 16280
rect 16726 16224 16731 16280
rect 12525 16222 16731 16224
rect 12525 16219 12591 16222
rect 16665 16219 16731 16222
rect 19701 16282 19767 16285
rect 19977 16282 20043 16285
rect 19701 16280 20043 16282
rect 19701 16224 19706 16280
rect 19762 16224 19982 16280
rect 20038 16224 20043 16280
rect 19701 16222 20043 16224
rect 19701 16219 19767 16222
rect 19977 16219 20043 16222
rect 20897 16282 20963 16285
rect 21214 16282 21220 16284
rect 20897 16280 21220 16282
rect 20897 16224 20902 16280
rect 20958 16224 21220 16280
rect 20897 16222 21220 16224
rect 20897 16219 20963 16222
rect 21214 16220 21220 16222
rect 21284 16282 21290 16284
rect 22188 16282 22248 16358
rect 25681 16355 25747 16358
rect 25865 16418 25931 16421
rect 26182 16418 26188 16420
rect 25865 16416 26188 16418
rect 25865 16360 25870 16416
rect 25926 16360 26188 16416
rect 25865 16358 26188 16360
rect 25865 16355 25931 16358
rect 26182 16356 26188 16358
rect 26252 16356 26258 16420
rect 28206 16356 28212 16420
rect 28276 16418 28282 16420
rect 30557 16418 30623 16421
rect 28276 16416 30623 16418
rect 28276 16360 30562 16416
rect 30618 16360 30623 16416
rect 28276 16358 30623 16360
rect 28276 16356 28282 16358
rect 30557 16355 30623 16358
rect 26980 16352 27296 16353
rect 26980 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27296 16352
rect 26980 16287 27296 16288
rect 21284 16222 22248 16282
rect 21284 16220 21290 16222
rect 22318 16220 22324 16284
rect 22388 16282 22394 16284
rect 26417 16282 26483 16285
rect 29545 16282 29611 16285
rect 22388 16280 26483 16282
rect 22388 16224 26422 16280
rect 26478 16224 26483 16280
rect 22388 16222 26483 16224
rect 22388 16220 22394 16222
rect 26417 16219 26483 16222
rect 27478 16280 29611 16282
rect 27478 16224 29550 16280
rect 29606 16224 29611 16280
rect 27478 16222 29611 16224
rect 10225 16144 12082 16146
rect 10225 16088 10230 16144
rect 10286 16088 12082 16144
rect 10225 16086 12082 16088
rect 12157 16146 12223 16149
rect 14273 16146 14339 16149
rect 24301 16146 24367 16149
rect 12157 16144 13876 16146
rect 12157 16088 12162 16144
rect 12218 16088 13876 16144
rect 12157 16086 13876 16088
rect 10225 16083 10291 16086
rect 12157 16083 12223 16086
rect 1577 16010 1643 16013
rect 11145 16010 11211 16013
rect 13537 16010 13603 16013
rect 1577 16008 11211 16010
rect 1577 15952 1582 16008
rect 1638 15952 11150 16008
rect 11206 15952 11211 16008
rect 1577 15950 11211 15952
rect 1577 15947 1643 15950
rect 11145 15947 11211 15950
rect 11884 16008 13603 16010
rect 11884 15952 13542 16008
rect 13598 15952 13603 16008
rect 11884 15950 13603 15952
rect 13816 16010 13876 16086
rect 14273 16144 24367 16146
rect 14273 16088 14278 16144
rect 14334 16088 24306 16144
rect 24362 16088 24367 16144
rect 14273 16086 24367 16088
rect 14273 16083 14339 16086
rect 24301 16083 24367 16086
rect 24761 16146 24827 16149
rect 27478 16146 27538 16222
rect 29545 16219 29611 16222
rect 24761 16144 27538 16146
rect 24761 16088 24766 16144
rect 24822 16088 27538 16144
rect 24761 16086 27538 16088
rect 27613 16146 27679 16149
rect 27981 16146 28047 16149
rect 27613 16144 28047 16146
rect 27613 16088 27618 16144
rect 27674 16088 27986 16144
rect 28042 16088 28047 16144
rect 27613 16086 28047 16088
rect 24761 16083 24827 16086
rect 27613 16083 27679 16086
rect 27981 16083 28047 16086
rect 28441 16146 28507 16149
rect 28901 16146 28967 16149
rect 28441 16144 28967 16146
rect 28441 16088 28446 16144
rect 28502 16088 28906 16144
rect 28962 16088 28967 16144
rect 28441 16086 28967 16088
rect 28441 16083 28507 16086
rect 28901 16083 28967 16086
rect 14825 16010 14891 16013
rect 16389 16010 16455 16013
rect 13816 16008 16455 16010
rect 13816 15952 14830 16008
rect 14886 15952 16394 16008
rect 16450 15952 16455 16008
rect 13816 15950 16455 15952
rect 8518 15812 8524 15876
rect 8588 15874 8594 15876
rect 8937 15874 9003 15877
rect 8588 15872 9003 15874
rect 8588 15816 8942 15872
rect 8998 15816 9003 15872
rect 8588 15814 9003 15816
rect 8588 15812 8594 15814
rect 8937 15811 9003 15814
rect 9489 15874 9555 15877
rect 11884 15874 11944 15950
rect 13537 15947 13603 15950
rect 14825 15947 14891 15950
rect 16389 15947 16455 15950
rect 18597 16010 18663 16013
rect 21449 16010 21515 16013
rect 18597 16008 21515 16010
rect 18597 15952 18602 16008
rect 18658 15952 21454 16008
rect 21510 15952 21515 16008
rect 18597 15950 21515 15952
rect 18597 15947 18663 15950
rect 21449 15947 21515 15950
rect 21633 16010 21699 16013
rect 21766 16010 21772 16012
rect 21633 16008 21772 16010
rect 21633 15952 21638 16008
rect 21694 15952 21772 16008
rect 21633 15950 21772 15952
rect 21633 15947 21699 15950
rect 21766 15948 21772 15950
rect 21836 15948 21842 16012
rect 22277 16010 22343 16013
rect 22502 16010 22508 16012
rect 22277 16008 22508 16010
rect 22277 15952 22282 16008
rect 22338 15952 22508 16008
rect 22277 15950 22508 15952
rect 22277 15947 22343 15950
rect 22502 15948 22508 15950
rect 22572 16010 22578 16012
rect 29453 16010 29519 16013
rect 22572 16008 29519 16010
rect 22572 15952 29458 16008
rect 29514 15952 29519 16008
rect 22572 15950 29519 15952
rect 22572 15948 22578 15950
rect 29453 15947 29519 15950
rect 9489 15872 11944 15874
rect 9489 15816 9494 15872
rect 9550 15816 11944 15872
rect 9489 15814 11944 15816
rect 12525 15876 12591 15877
rect 12525 15872 12572 15876
rect 12636 15874 12642 15876
rect 12985 15874 13051 15877
rect 13118 15874 13124 15876
rect 12525 15816 12530 15872
rect 9489 15811 9555 15814
rect 12525 15812 12572 15816
rect 12636 15814 12682 15874
rect 12985 15872 13124 15874
rect 12985 15816 12990 15872
rect 13046 15816 13124 15872
rect 12985 15814 13124 15816
rect 12636 15812 12642 15814
rect 12525 15811 12591 15812
rect 12985 15811 13051 15814
rect 13118 15812 13124 15814
rect 13188 15812 13194 15876
rect 13353 15874 13419 15877
rect 14181 15874 14247 15877
rect 17953 15874 18019 15877
rect 24577 15874 24643 15877
rect 13353 15872 14106 15874
rect 13353 15816 13358 15872
rect 13414 15816 14106 15872
rect 13353 15814 14106 15816
rect 13353 15811 13419 15814
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 12092 15808 12408 15809
rect 12092 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12408 15808
rect 12092 15743 12408 15744
rect 8293 15738 8359 15741
rect 9254 15738 9260 15740
rect 8293 15736 9260 15738
rect 8293 15680 8298 15736
rect 8354 15680 9260 15736
rect 8293 15678 9260 15680
rect 8293 15675 8359 15678
rect 9254 15676 9260 15678
rect 9324 15738 9330 15740
rect 11697 15738 11763 15741
rect 9324 15736 11763 15738
rect 9324 15680 11702 15736
rect 11758 15680 11763 15736
rect 9324 15678 11763 15680
rect 9324 15676 9330 15678
rect 11697 15675 11763 15678
rect 12617 15738 12683 15741
rect 14046 15738 14106 15814
rect 14181 15872 18019 15874
rect 14181 15816 14186 15872
rect 14242 15816 17958 15872
rect 18014 15816 18019 15872
rect 14181 15814 18019 15816
rect 14181 15811 14247 15814
rect 17953 15811 18019 15814
rect 20302 15872 24643 15874
rect 20302 15816 24582 15872
rect 24638 15816 24643 15872
rect 20302 15814 24643 15816
rect 19866 15808 20182 15809
rect 19866 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20182 15808
rect 19866 15743 20182 15744
rect 15653 15738 15719 15741
rect 12617 15736 13554 15738
rect 12617 15680 12622 15736
rect 12678 15680 13554 15736
rect 12617 15678 13554 15680
rect 14046 15736 15719 15738
rect 14046 15680 15658 15736
rect 15714 15680 15719 15736
rect 14046 15678 15719 15680
rect 12617 15675 12683 15678
rect 8385 15604 8451 15605
rect 8334 15602 8340 15604
rect 8294 15542 8340 15602
rect 8404 15600 8451 15604
rect 8446 15544 8451 15600
rect 8334 15540 8340 15542
rect 8404 15540 8451 15544
rect 8702 15540 8708 15604
rect 8772 15602 8778 15604
rect 9489 15602 9555 15605
rect 13353 15602 13419 15605
rect 8772 15600 13419 15602
rect 8772 15544 9494 15600
rect 9550 15544 13358 15600
rect 13414 15544 13419 15600
rect 8772 15542 13419 15544
rect 13494 15602 13554 15678
rect 15653 15675 15719 15678
rect 16665 15602 16731 15605
rect 20302 15602 20362 15814
rect 24577 15811 24643 15814
rect 28022 15812 28028 15876
rect 28092 15874 28098 15876
rect 28092 15814 29194 15874
rect 28092 15812 28098 15814
rect 27640 15808 27956 15809
rect 27640 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27956 15808
rect 27640 15743 27956 15744
rect 20437 15738 20503 15741
rect 21173 15738 21239 15741
rect 26182 15738 26188 15740
rect 20437 15736 26188 15738
rect 20437 15680 20442 15736
rect 20498 15680 21178 15736
rect 21234 15680 26188 15736
rect 20437 15678 26188 15680
rect 20437 15675 20503 15678
rect 21173 15675 21239 15678
rect 26182 15676 26188 15678
rect 26252 15676 26258 15740
rect 26366 15676 26372 15740
rect 26436 15738 26442 15740
rect 26693 15738 26759 15741
rect 26436 15736 26759 15738
rect 26436 15680 26698 15736
rect 26754 15680 26759 15736
rect 26436 15678 26759 15680
rect 26436 15676 26442 15678
rect 26693 15675 26759 15678
rect 23013 15604 23079 15605
rect 21950 15602 21956 15604
rect 13494 15542 16130 15602
rect 8772 15540 8778 15542
rect 8385 15539 8451 15540
rect 9489 15539 9555 15542
rect 13353 15539 13419 15542
rect 5533 15466 5599 15469
rect 15837 15466 15903 15469
rect 5533 15464 15903 15466
rect 5533 15408 5538 15464
rect 5594 15408 15842 15464
rect 15898 15408 15903 15464
rect 5533 15406 15903 15408
rect 16070 15466 16130 15542
rect 16665 15600 20362 15602
rect 16665 15544 16670 15600
rect 16726 15544 20362 15600
rect 16665 15542 20362 15544
rect 21406 15542 21956 15602
rect 16665 15539 16731 15542
rect 16757 15466 16823 15469
rect 18873 15466 18939 15469
rect 16070 15464 18939 15466
rect 16070 15408 16762 15464
rect 16818 15408 18878 15464
rect 18934 15408 18939 15464
rect 16070 15406 18939 15408
rect 5533 15403 5599 15406
rect 15837 15403 15903 15406
rect 16757 15403 16823 15406
rect 18873 15403 18939 15406
rect 19701 15466 19767 15469
rect 21173 15466 21239 15469
rect 21406 15468 21466 15542
rect 21950 15540 21956 15542
rect 22020 15540 22026 15604
rect 23013 15602 23060 15604
rect 22968 15600 23060 15602
rect 22968 15544 23018 15600
rect 22968 15542 23060 15544
rect 23013 15540 23060 15542
rect 23124 15540 23130 15604
rect 23238 15540 23244 15604
rect 23308 15602 23314 15604
rect 24301 15602 24367 15605
rect 23308 15600 24367 15602
rect 23308 15544 24306 15600
rect 24362 15544 24367 15600
rect 23308 15542 24367 15544
rect 23308 15540 23314 15542
rect 23013 15539 23079 15540
rect 24301 15539 24367 15542
rect 24761 15602 24827 15605
rect 28441 15602 28507 15605
rect 29134 15604 29194 15814
rect 28574 15602 28580 15604
rect 24761 15600 28580 15602
rect 24761 15544 24766 15600
rect 24822 15544 28446 15600
rect 28502 15544 28580 15600
rect 24761 15542 28580 15544
rect 24761 15539 24827 15542
rect 28441 15539 28507 15542
rect 28574 15540 28580 15542
rect 28644 15540 28650 15604
rect 29126 15602 29132 15604
rect 29044 15542 29132 15602
rect 29126 15540 29132 15542
rect 29196 15602 29202 15604
rect 29269 15602 29335 15605
rect 29196 15600 29335 15602
rect 29196 15544 29274 15600
rect 29330 15544 29335 15600
rect 29196 15542 29335 15544
rect 29196 15540 29202 15542
rect 29269 15539 29335 15542
rect 21398 15466 21404 15468
rect 19701 15464 21404 15466
rect 19701 15408 19706 15464
rect 19762 15408 21178 15464
rect 21234 15408 21404 15464
rect 19701 15406 21404 15408
rect 19701 15403 19767 15406
rect 21173 15403 21239 15406
rect 21398 15404 21404 15406
rect 21468 15404 21474 15468
rect 21817 15466 21883 15469
rect 27061 15466 27127 15469
rect 28022 15466 28028 15468
rect 21817 15464 28028 15466
rect 21817 15408 21822 15464
rect 21878 15408 27066 15464
rect 27122 15408 28028 15464
rect 21817 15406 28028 15408
rect 21817 15403 21883 15406
rect 27061 15403 27127 15406
rect 28022 15404 28028 15406
rect 28092 15404 28098 15468
rect 28206 15404 28212 15468
rect 28276 15466 28282 15468
rect 28349 15466 28415 15469
rect 30373 15466 30439 15469
rect 28276 15464 28415 15466
rect 28276 15408 28354 15464
rect 28410 15408 28415 15464
rect 28276 15406 28415 15408
rect 28276 15404 28282 15406
rect 28349 15403 28415 15406
rect 30100 15464 30439 15466
rect 30100 15408 30378 15464
rect 30434 15408 30439 15464
rect 30100 15406 30439 15408
rect 1158 15268 1164 15332
rect 1228 15330 1234 15332
rect 3141 15330 3207 15333
rect 1228 15328 3207 15330
rect 1228 15272 3146 15328
rect 3202 15272 3207 15328
rect 1228 15270 3207 15272
rect 1228 15268 1234 15270
rect 3141 15267 3207 15270
rect 7465 15330 7531 15333
rect 9949 15330 10015 15333
rect 7465 15328 10015 15330
rect 7465 15272 7470 15328
rect 7526 15272 9954 15328
rect 10010 15272 10015 15328
rect 7465 15270 10015 15272
rect 7465 15267 7531 15270
rect 9949 15267 10015 15270
rect 10225 15330 10291 15333
rect 11094 15330 11100 15332
rect 10225 15328 11100 15330
rect 10225 15272 10230 15328
rect 10286 15272 11100 15328
rect 10225 15270 11100 15272
rect 10225 15267 10291 15270
rect 11094 15268 11100 15270
rect 11164 15268 11170 15332
rect 11830 15268 11836 15332
rect 11900 15330 11906 15332
rect 12065 15330 12131 15333
rect 12617 15330 12683 15333
rect 11900 15328 12131 15330
rect 11900 15272 12070 15328
rect 12126 15272 12131 15328
rect 11900 15270 12131 15272
rect 11900 15268 11906 15270
rect 12065 15267 12131 15270
rect 12206 15328 12683 15330
rect 12206 15272 12622 15328
rect 12678 15272 12683 15328
rect 12206 15270 12683 15272
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 11432 15264 11748 15265
rect 11432 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11748 15264
rect 11432 15199 11748 15200
rect 5073 15194 5139 15197
rect 5758 15194 5764 15196
rect 5073 15192 5764 15194
rect 5073 15136 5078 15192
rect 5134 15136 5764 15192
rect 5073 15134 5764 15136
rect 5073 15131 5139 15134
rect 5758 15132 5764 15134
rect 5828 15132 5834 15196
rect 8017 15194 8083 15197
rect 10685 15194 10751 15197
rect 6870 15192 8083 15194
rect 6870 15136 8022 15192
rect 8078 15136 8083 15192
rect 6870 15134 8083 15136
rect 6870 15058 6930 15134
rect 8017 15131 8083 15134
rect 8158 15192 10751 15194
rect 8158 15136 10690 15192
rect 10746 15136 10751 15192
rect 8158 15134 10751 15136
rect 5812 14998 6930 15058
rect 7281 15058 7347 15061
rect 7966 15058 7972 15060
rect 7281 15056 7972 15058
rect 7281 15000 7286 15056
rect 7342 15000 7972 15056
rect 7281 14998 7972 15000
rect 5812 14925 5872 14998
rect 7281 14995 7347 14998
rect 7966 14996 7972 14998
rect 8036 15058 8042 15060
rect 8158 15058 8218 15134
rect 10685 15131 10751 15134
rect 11053 15194 11119 15197
rect 11278 15194 11284 15196
rect 11053 15192 11284 15194
rect 11053 15136 11058 15192
rect 11114 15136 11284 15192
rect 11053 15134 11284 15136
rect 11053 15131 11119 15134
rect 11278 15132 11284 15134
rect 11348 15132 11354 15196
rect 11881 15194 11947 15197
rect 12206 15194 12266 15270
rect 12617 15267 12683 15270
rect 13670 15268 13676 15332
rect 13740 15330 13746 15332
rect 14089 15330 14155 15333
rect 13740 15328 14155 15330
rect 13740 15272 14094 15328
rect 14150 15272 14155 15328
rect 13740 15270 14155 15272
rect 13740 15268 13746 15270
rect 14089 15267 14155 15270
rect 15101 15330 15167 15333
rect 15694 15330 15700 15332
rect 15101 15328 15700 15330
rect 15101 15272 15106 15328
rect 15162 15272 15700 15328
rect 15101 15270 15700 15272
rect 15101 15267 15167 15270
rect 15694 15268 15700 15270
rect 15764 15268 15770 15332
rect 19609 15330 19675 15333
rect 20897 15330 20963 15333
rect 19609 15328 20963 15330
rect 19609 15272 19614 15328
rect 19670 15272 20902 15328
rect 20958 15272 20963 15328
rect 19609 15270 20963 15272
rect 19609 15267 19675 15270
rect 20897 15267 20963 15270
rect 21449 15330 21515 15333
rect 24761 15330 24827 15333
rect 21449 15328 24827 15330
rect 21449 15272 21454 15328
rect 21510 15272 24766 15328
rect 24822 15272 24827 15328
rect 21449 15270 24827 15272
rect 21449 15267 21515 15270
rect 24761 15267 24827 15270
rect 27470 15268 27476 15332
rect 27540 15330 27546 15332
rect 30100 15330 30160 15406
rect 30373 15403 30439 15406
rect 30281 15332 30347 15333
rect 27540 15270 30160 15330
rect 27540 15268 27546 15270
rect 30230 15268 30236 15332
rect 30300 15330 30347 15332
rect 30300 15328 30392 15330
rect 30342 15272 30392 15328
rect 30300 15270 30392 15272
rect 30300 15268 30347 15270
rect 30281 15267 30347 15268
rect 19206 15264 19522 15265
rect 19206 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19522 15264
rect 19206 15199 19522 15200
rect 26980 15264 27296 15265
rect 26980 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27296 15264
rect 26980 15199 27296 15200
rect 11881 15192 12266 15194
rect 11881 15136 11886 15192
rect 11942 15136 12266 15192
rect 11881 15134 12266 15136
rect 12433 15194 12499 15197
rect 14641 15194 14707 15197
rect 12433 15192 14707 15194
rect 12433 15136 12438 15192
rect 12494 15136 14646 15192
rect 14702 15136 14707 15192
rect 12433 15134 14707 15136
rect 11881 15131 11947 15134
rect 12433 15131 12499 15134
rect 14641 15131 14707 15134
rect 16430 15132 16436 15196
rect 16500 15194 16506 15196
rect 16941 15194 17007 15197
rect 16500 15192 17007 15194
rect 16500 15136 16946 15192
rect 17002 15136 17007 15192
rect 16500 15134 17007 15136
rect 16500 15132 16506 15134
rect 16941 15131 17007 15134
rect 21449 15194 21515 15197
rect 22277 15194 22343 15197
rect 24025 15194 24091 15197
rect 25865 15196 25931 15197
rect 25814 15194 25820 15196
rect 21449 15192 24091 15194
rect 21449 15136 21454 15192
rect 21510 15136 22282 15192
rect 22338 15136 24030 15192
rect 24086 15136 24091 15192
rect 21449 15134 24091 15136
rect 25774 15134 25820 15194
rect 25884 15192 25931 15196
rect 25926 15136 25931 15192
rect 21449 15131 21515 15134
rect 22277 15131 22343 15134
rect 24025 15131 24091 15134
rect 25814 15132 25820 15134
rect 25884 15132 25931 15136
rect 25865 15131 25931 15132
rect 28993 15194 29059 15197
rect 30281 15194 30347 15197
rect 28993 15192 30347 15194
rect 28993 15136 28998 15192
rect 29054 15136 30286 15192
rect 30342 15136 30347 15192
rect 28993 15134 30347 15136
rect 28993 15131 29059 15134
rect 30281 15131 30347 15134
rect 8036 14998 8218 15058
rect 8937 15058 9003 15061
rect 10225 15058 10291 15061
rect 8937 15056 10291 15058
rect 8937 15000 8942 15056
rect 8998 15000 10230 15056
rect 10286 15000 10291 15056
rect 8937 14998 10291 15000
rect 8036 14996 8042 14998
rect 8937 14995 9003 14998
rect 10225 14995 10291 14998
rect 10777 15058 10843 15061
rect 11513 15058 11579 15061
rect 19333 15058 19399 15061
rect 10777 15056 11579 15058
rect 10777 15000 10782 15056
rect 10838 15000 11518 15056
rect 11574 15000 11579 15056
rect 10777 14998 11579 15000
rect 10777 14995 10843 14998
rect 11513 14995 11579 14998
rect 11654 15056 19399 15058
rect 11654 15000 19338 15056
rect 19394 15000 19399 15056
rect 11654 14998 19399 15000
rect 5809 14920 5875 14925
rect 5809 14864 5814 14920
rect 5870 14864 5875 14920
rect 5809 14859 5875 14864
rect 6913 14922 6979 14925
rect 7465 14922 7531 14925
rect 6913 14920 7531 14922
rect 6913 14864 6918 14920
rect 6974 14864 7470 14920
rect 7526 14864 7531 14920
rect 6913 14862 7531 14864
rect 6913 14859 6979 14862
rect 7465 14859 7531 14862
rect 7598 14860 7604 14924
rect 7668 14922 7674 14924
rect 10961 14922 11027 14925
rect 11421 14922 11487 14925
rect 7668 14862 10794 14922
rect 7668 14860 7674 14862
rect 7005 14786 7071 14789
rect 7465 14786 7531 14789
rect 9806 14786 9812 14788
rect 7005 14784 9812 14786
rect 7005 14728 7010 14784
rect 7066 14728 7470 14784
rect 7526 14728 9812 14784
rect 7005 14726 9812 14728
rect 7005 14723 7071 14726
rect 7465 14723 7531 14726
rect 9806 14724 9812 14726
rect 9876 14786 9882 14788
rect 10593 14786 10659 14789
rect 9876 14784 10659 14786
rect 9876 14728 10598 14784
rect 10654 14728 10659 14784
rect 9876 14726 10659 14728
rect 9876 14724 9882 14726
rect 10593 14723 10659 14726
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 6821 14650 6887 14653
rect 7598 14650 7604 14652
rect 6821 14648 7604 14650
rect 6821 14592 6826 14648
rect 6882 14592 7604 14648
rect 6821 14590 7604 14592
rect 6821 14587 6887 14590
rect 7598 14588 7604 14590
rect 7668 14588 7674 14652
rect 7925 14650 7991 14653
rect 8753 14650 8819 14653
rect 7925 14648 8819 14650
rect 7925 14592 7930 14648
rect 7986 14592 8758 14648
rect 8814 14592 8819 14648
rect 7925 14590 8819 14592
rect 10734 14650 10794 14862
rect 10961 14920 11487 14922
rect 10961 14864 10966 14920
rect 11022 14864 11426 14920
rect 11482 14864 11487 14920
rect 10961 14862 11487 14864
rect 10961 14859 11027 14862
rect 11421 14859 11487 14862
rect 10869 14786 10935 14789
rect 11654 14786 11714 14998
rect 19333 14995 19399 14998
rect 20989 15058 21055 15061
rect 26877 15058 26943 15061
rect 29545 15058 29611 15061
rect 20989 15056 26943 15058
rect 20989 15000 20994 15056
rect 21050 15000 26882 15056
rect 26938 15000 26943 15056
rect 20989 14998 26943 15000
rect 20989 14995 21055 14998
rect 26877 14995 26943 14998
rect 27064 15056 29611 15058
rect 27064 15000 29550 15056
rect 29606 15000 29611 15056
rect 27064 14998 29611 15000
rect 13813 14922 13879 14925
rect 10869 14784 11714 14786
rect 10869 14728 10874 14784
rect 10930 14728 11714 14784
rect 10869 14726 11714 14728
rect 11838 14920 13879 14922
rect 11838 14864 13818 14920
rect 13874 14864 13879 14920
rect 11838 14862 13879 14864
rect 10869 14723 10935 14726
rect 11838 14650 11898 14862
rect 13813 14859 13879 14862
rect 16941 14922 17007 14925
rect 22645 14922 22711 14925
rect 16941 14920 22711 14922
rect 16941 14864 16946 14920
rect 17002 14864 22650 14920
rect 22706 14864 22711 14920
rect 16941 14862 22711 14864
rect 16941 14859 17007 14862
rect 22645 14859 22711 14862
rect 23749 14922 23815 14925
rect 25221 14922 25287 14925
rect 27064 14922 27124 14998
rect 29545 14995 29611 14998
rect 27889 14922 27955 14925
rect 28441 14922 28507 14925
rect 23749 14920 25146 14922
rect 23749 14864 23754 14920
rect 23810 14864 25146 14920
rect 23749 14862 25146 14864
rect 23749 14859 23815 14862
rect 18045 14786 18111 14789
rect 12528 14784 18111 14786
rect 12528 14728 18050 14784
rect 18106 14728 18111 14784
rect 12528 14726 18111 14728
rect 12092 14720 12408 14721
rect 12092 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12408 14720
rect 12092 14655 12408 14656
rect 10734 14590 11898 14650
rect 7925 14587 7991 14590
rect 8753 14587 8819 14590
rect 8385 14516 8451 14517
rect 8334 14452 8340 14516
rect 8404 14514 8451 14516
rect 8753 14514 8819 14517
rect 10501 14514 10567 14517
rect 8404 14512 8496 14514
rect 8446 14456 8496 14512
rect 8404 14454 8496 14456
rect 8753 14512 10567 14514
rect 8753 14456 8758 14512
rect 8814 14456 10506 14512
rect 10562 14456 10567 14512
rect 8753 14454 10567 14456
rect 8404 14452 8451 14454
rect 8385 14451 8451 14452
rect 8753 14451 8819 14454
rect 10501 14451 10567 14454
rect 10685 14514 10751 14517
rect 12528 14514 12588 14726
rect 18045 14723 18111 14726
rect 20529 14786 20595 14789
rect 20846 14786 20852 14788
rect 20529 14784 20852 14786
rect 20529 14728 20534 14784
rect 20590 14728 20852 14784
rect 20529 14726 20852 14728
rect 20529 14723 20595 14726
rect 20846 14724 20852 14726
rect 20916 14786 20922 14788
rect 21725 14786 21791 14789
rect 23197 14786 23263 14789
rect 20916 14784 23263 14786
rect 20916 14728 21730 14784
rect 21786 14728 23202 14784
rect 23258 14728 23263 14784
rect 20916 14726 23263 14728
rect 20916 14724 20922 14726
rect 21725 14723 21791 14726
rect 23197 14723 23263 14726
rect 23841 14786 23907 14789
rect 24761 14786 24827 14789
rect 23841 14784 24827 14786
rect 23841 14728 23846 14784
rect 23902 14728 24766 14784
rect 24822 14728 24827 14784
rect 23841 14726 24827 14728
rect 25086 14786 25146 14862
rect 25221 14920 27124 14922
rect 25221 14864 25226 14920
rect 25282 14864 27124 14920
rect 25221 14862 27124 14864
rect 27478 14920 28507 14922
rect 27478 14864 27894 14920
rect 27950 14864 28446 14920
rect 28502 14864 28507 14920
rect 27478 14862 28507 14864
rect 25221 14859 25287 14862
rect 27478 14786 27538 14862
rect 27889 14859 27955 14862
rect 28441 14859 28507 14862
rect 29269 14922 29335 14925
rect 31385 14922 31451 14925
rect 29269 14920 31451 14922
rect 29269 14864 29274 14920
rect 29330 14864 31390 14920
rect 31446 14864 31451 14920
rect 29269 14862 31451 14864
rect 29269 14859 29335 14862
rect 31385 14859 31451 14862
rect 29913 14788 29979 14789
rect 25086 14726 27538 14786
rect 23841 14723 23907 14726
rect 24761 14723 24827 14726
rect 29862 14724 29868 14788
rect 29932 14786 29979 14788
rect 29932 14784 30024 14786
rect 29974 14728 30024 14784
rect 29932 14726 30024 14728
rect 29932 14724 29979 14726
rect 29913 14723 29979 14724
rect 19866 14720 20182 14721
rect 19866 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20182 14720
rect 19866 14655 20182 14656
rect 27640 14720 27956 14721
rect 27640 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27956 14720
rect 27640 14655 27956 14656
rect 12985 14650 13051 14653
rect 14038 14650 14044 14652
rect 12985 14648 14044 14650
rect 12985 14592 12990 14648
rect 13046 14592 14044 14648
rect 12985 14590 14044 14592
rect 12985 14587 13051 14590
rect 14038 14588 14044 14590
rect 14108 14588 14114 14652
rect 18086 14588 18092 14652
rect 18156 14650 18162 14652
rect 18413 14650 18479 14653
rect 18156 14648 18479 14650
rect 18156 14592 18418 14648
rect 18474 14592 18479 14648
rect 18156 14590 18479 14592
rect 18156 14588 18162 14590
rect 18413 14587 18479 14590
rect 18822 14588 18828 14652
rect 18892 14650 18898 14652
rect 18965 14650 19031 14653
rect 18892 14648 19031 14650
rect 18892 14592 18970 14648
rect 19026 14592 19031 14648
rect 18892 14590 19031 14592
rect 18892 14588 18898 14590
rect 18965 14587 19031 14590
rect 19333 14650 19399 14653
rect 19701 14650 19767 14653
rect 19333 14648 19767 14650
rect 19333 14592 19338 14648
rect 19394 14592 19706 14648
rect 19762 14592 19767 14648
rect 19333 14590 19767 14592
rect 19333 14587 19399 14590
rect 19701 14587 19767 14590
rect 20662 14588 20668 14652
rect 20732 14650 20738 14652
rect 22461 14650 22527 14653
rect 20732 14648 22527 14650
rect 20732 14592 22466 14648
rect 22522 14592 22527 14648
rect 20732 14590 22527 14592
rect 20732 14588 20738 14590
rect 22461 14587 22527 14590
rect 23749 14650 23815 14653
rect 25589 14650 25655 14653
rect 23749 14648 25655 14650
rect 23749 14592 23754 14648
rect 23810 14592 25594 14648
rect 25650 14592 25655 14648
rect 23749 14590 25655 14592
rect 23749 14587 23815 14590
rect 25589 14587 25655 14590
rect 25957 14650 26023 14653
rect 26693 14650 26759 14653
rect 25957 14648 26759 14650
rect 25957 14592 25962 14648
rect 26018 14592 26698 14648
rect 26754 14592 26759 14648
rect 25957 14590 26759 14592
rect 25957 14587 26023 14590
rect 26693 14587 26759 14590
rect 10685 14512 12588 14514
rect 10685 14456 10690 14512
rect 10746 14456 12588 14512
rect 10685 14454 12588 14456
rect 13077 14514 13143 14517
rect 13629 14514 13695 14517
rect 24025 14514 24091 14517
rect 13077 14512 13554 14514
rect 13077 14456 13082 14512
rect 13138 14456 13554 14512
rect 13077 14454 13554 14456
rect 10685 14451 10751 14454
rect 13077 14451 13143 14454
rect 7230 14316 7236 14380
rect 7300 14378 7306 14380
rect 8017 14378 8083 14381
rect 8569 14380 8635 14381
rect 8518 14378 8524 14380
rect 7300 14376 8083 14378
rect 7300 14320 8022 14376
rect 8078 14320 8083 14376
rect 7300 14318 8083 14320
rect 8478 14318 8524 14378
rect 8588 14376 8635 14380
rect 8630 14320 8635 14376
rect 7300 14316 7306 14318
rect 8017 14315 8083 14318
rect 8518 14316 8524 14318
rect 8588 14316 8635 14320
rect 8569 14315 8635 14316
rect 10225 14378 10291 14381
rect 13261 14378 13327 14381
rect 10225 14376 13327 14378
rect 10225 14320 10230 14376
rect 10286 14320 13266 14376
rect 13322 14320 13327 14376
rect 10225 14318 13327 14320
rect 13494 14378 13554 14454
rect 13629 14512 24091 14514
rect 13629 14456 13634 14512
rect 13690 14456 24030 14512
rect 24086 14456 24091 14512
rect 13629 14454 24091 14456
rect 13629 14451 13695 14454
rect 24025 14451 24091 14454
rect 24158 14452 24164 14516
rect 24228 14514 24234 14516
rect 24301 14514 24367 14517
rect 28257 14514 28323 14517
rect 24228 14512 28323 14514
rect 24228 14456 24306 14512
rect 24362 14456 28262 14512
rect 28318 14456 28323 14512
rect 24228 14454 28323 14456
rect 24228 14452 24234 14454
rect 24301 14451 24367 14454
rect 28257 14451 28323 14454
rect 14825 14378 14891 14381
rect 13494 14376 14891 14378
rect 13494 14320 14830 14376
rect 14886 14320 14891 14376
rect 13494 14318 14891 14320
rect 10225 14315 10291 14318
rect 13261 14315 13327 14318
rect 14825 14315 14891 14318
rect 14958 14316 14964 14380
rect 15028 14378 15034 14380
rect 15101 14378 15167 14381
rect 15028 14376 15167 14378
rect 15028 14320 15106 14376
rect 15162 14320 15167 14376
rect 15028 14318 15167 14320
rect 15028 14316 15034 14318
rect 15101 14315 15167 14318
rect 15285 14378 15351 14381
rect 18597 14378 18663 14381
rect 19149 14378 19215 14381
rect 15285 14376 19215 14378
rect 15285 14320 15290 14376
rect 15346 14320 18602 14376
rect 18658 14320 19154 14376
rect 19210 14320 19215 14376
rect 15285 14318 19215 14320
rect 15285 14315 15351 14318
rect 18597 14315 18663 14318
rect 19149 14315 19215 14318
rect 19333 14378 19399 14381
rect 23013 14378 23079 14381
rect 19333 14376 23079 14378
rect 19333 14320 19338 14376
rect 19394 14320 23018 14376
rect 23074 14320 23079 14376
rect 19333 14318 23079 14320
rect 19333 14315 19399 14318
rect 23013 14315 23079 14318
rect 25998 14316 26004 14380
rect 26068 14378 26074 14380
rect 26969 14378 27035 14381
rect 26068 14376 27035 14378
rect 26068 14320 26974 14376
rect 27030 14320 27035 14376
rect 26068 14318 27035 14320
rect 26068 14316 26074 14318
rect 26969 14315 27035 14318
rect 5533 14242 5599 14245
rect 7465 14242 7531 14245
rect 5533 14240 7531 14242
rect 5533 14184 5538 14240
rect 5594 14184 7470 14240
rect 7526 14184 7531 14240
rect 5533 14182 7531 14184
rect 5533 14179 5599 14182
rect 7465 14179 7531 14182
rect 8293 14242 8359 14245
rect 10593 14242 10659 14245
rect 10726 14242 10732 14244
rect 8293 14240 10732 14242
rect 8293 14184 8298 14240
rect 8354 14184 10598 14240
rect 10654 14184 10732 14240
rect 8293 14182 10732 14184
rect 8293 14179 8359 14182
rect 10593 14179 10659 14182
rect 10726 14180 10732 14182
rect 10796 14180 10802 14244
rect 11973 14240 12039 14245
rect 11973 14184 11978 14240
rect 12034 14184 12039 14240
rect 11973 14179 12039 14184
rect 12617 14242 12683 14245
rect 17401 14242 17467 14245
rect 12617 14240 17467 14242
rect 12617 14184 12622 14240
rect 12678 14184 17406 14240
rect 17462 14184 17467 14240
rect 12617 14182 17467 14184
rect 12617 14179 12683 14182
rect 17401 14179 17467 14182
rect 21541 14242 21607 14245
rect 25957 14242 26023 14245
rect 21541 14240 26023 14242
rect 21541 14184 21546 14240
rect 21602 14184 25962 14240
rect 26018 14184 26023 14240
rect 21541 14182 26023 14184
rect 21541 14179 21607 14182
rect 25957 14179 26023 14182
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 11432 14176 11748 14177
rect 11432 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11748 14176
rect 11432 14111 11748 14112
rect 5073 14106 5139 14109
rect 10041 14106 10107 14109
rect 10593 14106 10659 14109
rect 5073 14104 10659 14106
rect 5073 14048 5078 14104
rect 5134 14048 10046 14104
rect 10102 14048 10598 14104
rect 10654 14048 10659 14104
rect 5073 14046 10659 14048
rect 5073 14043 5139 14046
rect 10041 14043 10107 14046
rect 10593 14043 10659 14046
rect 11053 14106 11119 14109
rect 11237 14106 11303 14109
rect 11053 14104 11303 14106
rect 11053 14048 11058 14104
rect 11114 14048 11242 14104
rect 11298 14048 11303 14104
rect 11053 14046 11303 14048
rect 11976 14106 12036 14179
rect 19206 14176 19522 14177
rect 19206 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19522 14176
rect 19206 14111 19522 14112
rect 26980 14176 27296 14177
rect 26980 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27296 14176
rect 26980 14111 27296 14112
rect 14825 14106 14891 14109
rect 11976 14104 14891 14106
rect 11976 14048 14830 14104
rect 14886 14048 14891 14104
rect 11976 14046 14891 14048
rect 11053 14043 11119 14046
rect 11237 14043 11303 14046
rect 14825 14043 14891 14046
rect 15009 14106 15075 14109
rect 16941 14106 17007 14109
rect 15009 14104 17007 14106
rect 15009 14048 15014 14104
rect 15070 14048 16946 14104
rect 17002 14048 17007 14104
rect 15009 14046 17007 14048
rect 15009 14043 15075 14046
rect 16941 14043 17007 14046
rect 17769 14106 17835 14109
rect 23565 14106 23631 14109
rect 17769 14104 19120 14106
rect 17769 14048 17774 14104
rect 17830 14048 19120 14104
rect 17769 14046 19120 14048
rect 17769 14043 17835 14046
rect 19060 14004 19120 14046
rect 19612 14104 23631 14106
rect 19612 14048 23570 14104
rect 23626 14048 23631 14104
rect 19612 14046 23631 14048
rect 19612 14004 19672 14046
rect 23565 14043 23631 14046
rect 25129 14106 25195 14109
rect 26693 14106 26759 14109
rect 25129 14104 26759 14106
rect 25129 14048 25134 14104
rect 25190 14048 26698 14104
rect 26754 14048 26759 14104
rect 25129 14046 26759 14048
rect 25129 14043 25195 14046
rect 26693 14043 26759 14046
rect 1853 13970 1919 13973
rect 13629 13970 13695 13973
rect 1853 13968 13695 13970
rect 1853 13912 1858 13968
rect 1914 13912 13634 13968
rect 13690 13912 13695 13968
rect 1853 13910 13695 13912
rect 1853 13907 1919 13910
rect 13629 13907 13695 13910
rect 15101 13970 15167 13973
rect 15101 13968 18522 13970
rect 15101 13912 15106 13968
rect 15162 13912 18522 13968
rect 19060 13944 19672 14004
rect 21449 13970 21515 13973
rect 21817 13972 21883 13973
rect 19750 13968 21515 13970
rect 15101 13910 18522 13912
rect 15101 13907 15167 13910
rect 2221 13834 2287 13837
rect 5073 13834 5139 13837
rect 2221 13832 5139 13834
rect 2221 13776 2226 13832
rect 2282 13776 5078 13832
rect 5134 13776 5139 13832
rect 2221 13774 5139 13776
rect 2221 13771 2287 13774
rect 5073 13771 5139 13774
rect 5758 13772 5764 13836
rect 5828 13834 5834 13836
rect 6177 13834 6243 13837
rect 7557 13834 7623 13837
rect 8753 13836 8819 13837
rect 5828 13832 6243 13834
rect 5828 13776 6182 13832
rect 6238 13776 6243 13832
rect 5828 13774 6243 13776
rect 5828 13772 5834 13774
rect 6177 13771 6243 13774
rect 6318 13832 7623 13834
rect 6318 13776 7562 13832
rect 7618 13776 7623 13832
rect 6318 13774 7623 13776
rect 6126 13636 6132 13700
rect 6196 13698 6202 13700
rect 6318 13698 6378 13774
rect 7557 13771 7623 13774
rect 8702 13772 8708 13836
rect 8772 13834 8819 13836
rect 9397 13834 9463 13837
rect 16297 13834 16363 13837
rect 8772 13832 8864 13834
rect 8814 13776 8864 13832
rect 8772 13774 8864 13776
rect 9397 13832 16363 13834
rect 9397 13776 9402 13832
rect 9458 13776 16302 13832
rect 16358 13776 16363 13832
rect 9397 13774 16363 13776
rect 8772 13772 8819 13774
rect 8753 13771 8819 13772
rect 9397 13771 9463 13774
rect 16297 13771 16363 13774
rect 16849 13834 16915 13837
rect 18229 13834 18295 13837
rect 16849 13832 18295 13834
rect 16849 13776 16854 13832
rect 16910 13776 18234 13832
rect 18290 13776 18295 13832
rect 16849 13774 18295 13776
rect 18462 13834 18522 13910
rect 19750 13912 21454 13968
rect 21510 13912 21515 13968
rect 19750 13910 21515 13912
rect 19290 13834 19488 13868
rect 19750 13834 19810 13910
rect 21449 13907 21515 13910
rect 21766 13908 21772 13972
rect 21836 13970 21883 13972
rect 22737 13970 22803 13973
rect 23197 13970 23263 13973
rect 21836 13968 21928 13970
rect 21878 13912 21928 13968
rect 21836 13910 21928 13912
rect 22737 13968 23263 13970
rect 22737 13912 22742 13968
rect 22798 13912 23202 13968
rect 23258 13912 23263 13968
rect 22737 13910 23263 13912
rect 21836 13908 21883 13910
rect 21817 13907 21883 13908
rect 22737 13907 22803 13910
rect 23197 13907 23263 13910
rect 23381 13970 23447 13973
rect 25957 13970 26023 13973
rect 26693 13972 26759 13973
rect 28809 13972 28875 13973
rect 26693 13970 26740 13972
rect 23381 13968 26023 13970
rect 23381 13912 23386 13968
rect 23442 13912 25962 13968
rect 26018 13912 26023 13968
rect 23381 13910 26023 13912
rect 26648 13968 26740 13970
rect 26648 13912 26698 13968
rect 26648 13910 26740 13912
rect 23381 13907 23447 13910
rect 25957 13907 26023 13910
rect 26693 13908 26740 13910
rect 26804 13908 26810 13972
rect 28758 13908 28764 13972
rect 28828 13970 28875 13972
rect 28828 13968 28920 13970
rect 28870 13912 28920 13968
rect 28828 13910 28920 13912
rect 28828 13908 28875 13910
rect 26693 13907 26759 13908
rect 28809 13907 28875 13908
rect 18462 13808 19810 13834
rect 18462 13774 19350 13808
rect 19428 13774 19810 13808
rect 19885 13834 19951 13837
rect 20529 13834 20595 13837
rect 19885 13832 20595 13834
rect 19885 13776 19890 13832
rect 19946 13776 20534 13832
rect 20590 13776 20595 13832
rect 19885 13774 20595 13776
rect 16849 13771 16915 13774
rect 18229 13771 18295 13774
rect 19885 13771 19951 13774
rect 20529 13771 20595 13774
rect 20805 13834 20871 13837
rect 22134 13834 22140 13836
rect 20805 13832 22140 13834
rect 20805 13776 20810 13832
rect 20866 13776 22140 13832
rect 20805 13774 22140 13776
rect 20805 13771 20871 13774
rect 22134 13772 22140 13774
rect 22204 13834 22210 13836
rect 23105 13834 23171 13837
rect 22204 13832 23171 13834
rect 22204 13776 23110 13832
rect 23166 13776 23171 13832
rect 22204 13774 23171 13776
rect 22204 13772 22210 13774
rect 23105 13771 23171 13774
rect 24485 13836 24551 13837
rect 24485 13832 24532 13836
rect 24596 13834 24602 13836
rect 25313 13834 25379 13837
rect 29494 13834 29500 13836
rect 24485 13776 24490 13832
rect 24485 13772 24532 13776
rect 24596 13774 24642 13834
rect 25313 13832 29500 13834
rect 25313 13776 25318 13832
rect 25374 13776 29500 13832
rect 25313 13774 29500 13776
rect 24596 13772 24602 13774
rect 24485 13771 24551 13772
rect 25313 13771 25379 13774
rect 29494 13772 29500 13774
rect 29564 13834 29570 13836
rect 30373 13834 30439 13837
rect 29564 13832 30439 13834
rect 29564 13776 30378 13832
rect 30434 13776 30439 13832
rect 29564 13774 30439 13776
rect 29564 13772 29570 13774
rect 30373 13771 30439 13774
rect 6196 13638 6378 13698
rect 7557 13698 7623 13701
rect 7966 13698 7972 13700
rect 7557 13696 7972 13698
rect 7557 13640 7562 13696
rect 7618 13640 7972 13696
rect 7557 13638 7972 13640
rect 6196 13636 6202 13638
rect 7557 13635 7623 13638
rect 7966 13636 7972 13638
rect 8036 13636 8042 13700
rect 8385 13698 8451 13701
rect 10777 13698 10843 13701
rect 8385 13696 10843 13698
rect 8385 13640 8390 13696
rect 8446 13640 10782 13696
rect 10838 13640 10843 13696
rect 8385 13638 10843 13640
rect 8385 13635 8451 13638
rect 10777 13635 10843 13638
rect 10910 13636 10916 13700
rect 10980 13698 10986 13700
rect 11830 13698 11836 13700
rect 10980 13638 11836 13698
rect 10980 13636 10986 13638
rect 11830 13636 11836 13638
rect 11900 13636 11906 13700
rect 12801 13698 12867 13701
rect 12934 13698 12940 13700
rect 12801 13696 12940 13698
rect 12801 13640 12806 13696
rect 12862 13640 12940 13696
rect 12801 13638 12940 13640
rect 12801 13635 12867 13638
rect 12934 13636 12940 13638
rect 13004 13636 13010 13700
rect 13261 13698 13327 13701
rect 15285 13698 15351 13701
rect 13261 13696 15351 13698
rect 13261 13640 13266 13696
rect 13322 13640 15290 13696
rect 15346 13640 15351 13696
rect 13261 13638 15351 13640
rect 13261 13635 13327 13638
rect 15285 13635 15351 13638
rect 16481 13698 16547 13701
rect 18965 13698 19031 13701
rect 16481 13696 19031 13698
rect 16481 13640 16486 13696
rect 16542 13640 18970 13696
rect 19026 13640 19031 13696
rect 16481 13638 19031 13640
rect 16481 13635 16547 13638
rect 18965 13635 19031 13638
rect 19149 13698 19215 13701
rect 19609 13698 19675 13701
rect 19149 13696 19675 13698
rect 19149 13640 19154 13696
rect 19210 13640 19614 13696
rect 19670 13640 19675 13696
rect 19149 13638 19675 13640
rect 19149 13635 19215 13638
rect 19609 13635 19675 13638
rect 20253 13698 20319 13701
rect 22185 13698 22251 13701
rect 20253 13696 22251 13698
rect 20253 13640 20258 13696
rect 20314 13640 22190 13696
rect 22246 13640 22251 13696
rect 20253 13638 22251 13640
rect 20253 13635 20319 13638
rect 22185 13635 22251 13638
rect 24117 13698 24183 13701
rect 24945 13698 25011 13701
rect 26233 13698 26299 13701
rect 26785 13700 26851 13701
rect 26734 13698 26740 13700
rect 24117 13696 25011 13698
rect 24117 13640 24122 13696
rect 24178 13640 24950 13696
rect 25006 13640 25011 13696
rect 24117 13638 25011 13640
rect 24117 13635 24183 13638
rect 24945 13635 25011 13638
rect 25086 13696 26299 13698
rect 25086 13640 26238 13696
rect 26294 13640 26299 13696
rect 25086 13638 26299 13640
rect 26694 13638 26740 13698
rect 26804 13696 26851 13700
rect 26846 13640 26851 13696
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 12092 13632 12408 13633
rect 12092 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12408 13632
rect 12092 13567 12408 13568
rect 19866 13632 20182 13633
rect 19866 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20182 13632
rect 19866 13567 20182 13568
rect 4797 13562 4863 13565
rect 6177 13562 6243 13565
rect 4797 13560 6243 13562
rect 4797 13504 4802 13560
rect 4858 13504 6182 13560
rect 6238 13504 6243 13560
rect 4797 13502 6243 13504
rect 4797 13499 4863 13502
rect 6177 13499 6243 13502
rect 8201 13562 8267 13565
rect 9438 13562 9444 13564
rect 8201 13560 9444 13562
rect 8201 13504 8206 13560
rect 8262 13504 9444 13560
rect 8201 13502 9444 13504
rect 8201 13499 8267 13502
rect 9438 13500 9444 13502
rect 9508 13500 9514 13564
rect 9857 13562 9923 13565
rect 10409 13562 10475 13565
rect 9857 13560 10475 13562
rect 9857 13504 9862 13560
rect 9918 13504 10414 13560
rect 10470 13504 10475 13560
rect 9857 13502 10475 13504
rect 9857 13499 9923 13502
rect 10409 13499 10475 13502
rect 10726 13500 10732 13564
rect 10796 13562 10802 13564
rect 11697 13562 11763 13565
rect 10796 13560 11763 13562
rect 10796 13504 11702 13560
rect 11758 13504 11763 13560
rect 10796 13502 11763 13504
rect 10796 13500 10802 13502
rect 11697 13499 11763 13502
rect 12525 13562 12591 13565
rect 12934 13562 12940 13564
rect 12525 13560 12940 13562
rect 12525 13504 12530 13560
rect 12586 13504 12940 13560
rect 12525 13502 12940 13504
rect 12525 13499 12591 13502
rect 12934 13500 12940 13502
rect 13004 13500 13010 13564
rect 13854 13500 13860 13564
rect 13924 13562 13930 13564
rect 14733 13562 14799 13565
rect 13924 13560 14799 13562
rect 13924 13504 14738 13560
rect 14794 13504 14799 13560
rect 13924 13502 14799 13504
rect 13924 13500 13930 13502
rect 14733 13499 14799 13502
rect 15837 13562 15903 13565
rect 22318 13562 22324 13564
rect 15837 13560 19764 13562
rect 15837 13504 15842 13560
rect 15898 13504 19764 13560
rect 15837 13502 19764 13504
rect 15837 13499 15903 13502
rect 8845 13426 8911 13429
rect 2730 13424 8911 13426
rect 2730 13368 8850 13424
rect 8906 13368 8911 13424
rect 2730 13366 8911 13368
rect 841 13290 907 13293
rect 2730 13290 2790 13366
rect 8845 13363 8911 13366
rect 9489 13426 9555 13429
rect 16205 13426 16271 13429
rect 16849 13426 16915 13429
rect 19704 13426 19764 13502
rect 20348 13502 22324 13562
rect 20348 13426 20408 13502
rect 22318 13500 22324 13502
rect 22388 13562 22394 13564
rect 24209 13562 24275 13565
rect 22388 13560 24275 13562
rect 22388 13504 24214 13560
rect 24270 13504 24275 13560
rect 22388 13502 24275 13504
rect 22388 13500 22394 13502
rect 24209 13499 24275 13502
rect 24342 13500 24348 13564
rect 24412 13562 24418 13564
rect 24669 13562 24735 13565
rect 24412 13560 24735 13562
rect 24412 13504 24674 13560
rect 24730 13504 24735 13560
rect 24412 13502 24735 13504
rect 24412 13500 24418 13502
rect 24669 13499 24735 13502
rect 9489 13424 16915 13426
rect 9489 13368 9494 13424
rect 9550 13368 16210 13424
rect 16266 13368 16854 13424
rect 16910 13368 16915 13424
rect 9489 13366 16915 13368
rect 9489 13363 9555 13366
rect 16205 13363 16271 13366
rect 16849 13363 16915 13366
rect 17174 13366 19442 13426
rect 19704 13366 20408 13426
rect 21449 13426 21515 13429
rect 25086 13426 25146 13638
rect 26233 13635 26299 13638
rect 26734 13636 26740 13638
rect 26804 13636 26851 13640
rect 26785 13635 26851 13636
rect 27640 13632 27956 13633
rect 27640 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27956 13632
rect 27640 13567 27956 13568
rect 25221 13562 25287 13565
rect 26969 13562 27035 13565
rect 25221 13560 27035 13562
rect 25221 13504 25226 13560
rect 25282 13504 26974 13560
rect 27030 13504 27035 13560
rect 25221 13502 27035 13504
rect 25221 13499 25287 13502
rect 26969 13499 27035 13502
rect 21449 13424 25146 13426
rect 21449 13368 21454 13424
rect 21510 13368 25146 13424
rect 21449 13366 25146 13368
rect 25313 13426 25379 13429
rect 28206 13426 28212 13428
rect 25313 13424 28212 13426
rect 25313 13368 25318 13424
rect 25374 13368 28212 13424
rect 25313 13366 28212 13368
rect 841 13288 2790 13290
rect 841 13232 846 13288
rect 902 13232 2790 13288
rect 841 13230 2790 13232
rect 3325 13290 3391 13293
rect 9213 13290 9279 13293
rect 3325 13288 9279 13290
rect 3325 13232 3330 13288
rect 3386 13232 9218 13288
rect 9274 13232 9279 13288
rect 3325 13230 9279 13232
rect 841 13227 907 13230
rect 3325 13227 3391 13230
rect 9213 13227 9279 13230
rect 11145 13290 11211 13293
rect 17033 13290 17099 13293
rect 11145 13288 17099 13290
rect 11145 13232 11150 13288
rect 11206 13232 17038 13288
rect 17094 13232 17099 13288
rect 11145 13230 17099 13232
rect 11145 13227 11211 13230
rect 17033 13227 17099 13230
rect 5349 13154 5415 13157
rect 8017 13154 8083 13157
rect 5349 13152 8083 13154
rect 5349 13096 5354 13152
rect 5410 13096 8022 13152
rect 8078 13096 8083 13152
rect 5349 13094 8083 13096
rect 5349 13091 5415 13094
rect 8017 13091 8083 13094
rect 8150 13092 8156 13156
rect 8220 13154 8226 13156
rect 8477 13154 8543 13157
rect 8220 13152 8543 13154
rect 8220 13096 8482 13152
rect 8538 13096 8543 13152
rect 8220 13094 8543 13096
rect 8220 13092 8226 13094
rect 8477 13091 8543 13094
rect 9581 13156 9647 13157
rect 9581 13152 9628 13156
rect 9692 13154 9698 13156
rect 10041 13154 10107 13157
rect 10869 13154 10935 13157
rect 17174 13154 17234 13366
rect 17585 13290 17651 13293
rect 18873 13290 18939 13293
rect 17585 13288 18939 13290
rect 17585 13232 17590 13288
rect 17646 13232 18878 13288
rect 18934 13232 18939 13288
rect 17585 13230 18939 13232
rect 17585 13227 17651 13230
rect 18873 13227 18939 13230
rect 19006 13228 19012 13292
rect 19076 13290 19082 13292
rect 19149 13290 19215 13293
rect 19076 13288 19215 13290
rect 19076 13232 19154 13288
rect 19210 13232 19215 13288
rect 19076 13230 19215 13232
rect 19382 13290 19442 13366
rect 21449 13363 21515 13366
rect 25313 13363 25379 13366
rect 28206 13364 28212 13366
rect 28276 13364 28282 13428
rect 22645 13290 22711 13293
rect 24485 13290 24551 13293
rect 27981 13290 28047 13293
rect 19382 13288 22711 13290
rect 19382 13232 22650 13288
rect 22706 13232 22711 13288
rect 19382 13230 22711 13232
rect 19076 13228 19082 13230
rect 19149 13227 19215 13230
rect 22645 13227 22711 13230
rect 22832 13288 28047 13290
rect 22832 13232 24490 13288
rect 24546 13232 27986 13288
rect 28042 13232 28047 13288
rect 22832 13230 28047 13232
rect 9581 13096 9586 13152
rect 9581 13092 9628 13096
rect 9692 13094 9738 13154
rect 10041 13152 10935 13154
rect 10041 13096 10046 13152
rect 10102 13096 10874 13152
rect 10930 13096 10935 13152
rect 10041 13094 10935 13096
rect 9692 13092 9698 13094
rect 9581 13091 9647 13092
rect 10041 13091 10107 13094
rect 10869 13091 10935 13094
rect 11838 13094 17234 13154
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 11432 13088 11748 13089
rect 11432 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11748 13088
rect 11432 13023 11748 13024
rect 5073 13020 5139 13021
rect 5022 13018 5028 13020
rect 4982 12958 5028 13018
rect 5092 13018 5139 13020
rect 10961 13018 11027 13021
rect 5092 13016 11027 13018
rect 5134 12960 10966 13016
rect 11022 12960 11027 13016
rect 5022 12956 5028 12958
rect 5092 12958 11027 12960
rect 5092 12956 5139 12958
rect 5073 12955 5139 12956
rect 10961 12955 11027 12958
rect 2998 12820 3004 12884
rect 3068 12882 3074 12884
rect 4429 12882 4495 12885
rect 3068 12880 4495 12882
rect 3068 12824 4434 12880
rect 4490 12824 4495 12880
rect 3068 12822 4495 12824
rect 3068 12820 3074 12822
rect 4429 12819 4495 12822
rect 4705 12882 4771 12885
rect 4838 12882 4844 12884
rect 4705 12880 4844 12882
rect 4705 12824 4710 12880
rect 4766 12824 4844 12880
rect 4705 12822 4844 12824
rect 4705 12819 4771 12822
rect 4838 12820 4844 12822
rect 4908 12820 4914 12884
rect 5533 12882 5599 12885
rect 9489 12882 9555 12885
rect 5533 12880 9555 12882
rect 5533 12824 5538 12880
rect 5594 12824 9494 12880
rect 9550 12824 9555 12880
rect 5533 12822 9555 12824
rect 5533 12819 5599 12822
rect 9489 12819 9555 12822
rect 10225 12882 10291 12885
rect 11838 12882 11898 13094
rect 17350 13092 17356 13156
rect 17420 13154 17426 13156
rect 17769 13154 17835 13157
rect 22832 13154 22892 13230
rect 24485 13227 24551 13230
rect 27981 13227 28047 13230
rect 17420 13152 17835 13154
rect 17420 13096 17774 13152
rect 17830 13096 17835 13152
rect 17420 13094 17835 13096
rect 17420 13092 17426 13094
rect 17769 13091 17835 13094
rect 19612 13094 22892 13154
rect 24209 13154 24275 13157
rect 24669 13154 24735 13157
rect 24209 13152 24735 13154
rect 24209 13096 24214 13152
rect 24270 13096 24674 13152
rect 24730 13096 24735 13152
rect 24209 13094 24735 13096
rect 19206 13088 19522 13089
rect 19206 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19522 13088
rect 19206 13023 19522 13024
rect 12249 13018 12315 13021
rect 17953 13018 18019 13021
rect 12249 13016 18019 13018
rect 12249 12960 12254 13016
rect 12310 12960 17958 13016
rect 18014 12960 18019 13016
rect 12249 12958 18019 12960
rect 12249 12955 12315 12958
rect 17953 12955 18019 12958
rect 10225 12880 11898 12882
rect 10225 12824 10230 12880
rect 10286 12824 11898 12880
rect 10225 12822 11898 12824
rect 12157 12882 12223 12885
rect 13629 12882 13695 12885
rect 16614 12882 16620 12884
rect 12157 12880 16620 12882
rect 12157 12824 12162 12880
rect 12218 12824 13634 12880
rect 13690 12824 16620 12880
rect 12157 12822 16620 12824
rect 10225 12819 10291 12822
rect 12157 12819 12223 12822
rect 13629 12819 13695 12822
rect 16614 12820 16620 12822
rect 16684 12820 16690 12884
rect 17585 12882 17651 12885
rect 18270 12882 18276 12884
rect 17585 12880 18276 12882
rect 17585 12824 17590 12880
rect 17646 12824 18276 12880
rect 17585 12822 18276 12824
rect 17585 12819 17651 12822
rect 18270 12820 18276 12822
rect 18340 12882 18346 12884
rect 19612 12882 19672 13094
rect 24209 13091 24275 13094
rect 24669 13091 24735 13094
rect 25865 13154 25931 13157
rect 26417 13154 26483 13157
rect 25865 13152 26483 13154
rect 25865 13096 25870 13152
rect 25926 13096 26422 13152
rect 26478 13096 26483 13152
rect 25865 13094 26483 13096
rect 25865 13091 25931 13094
rect 26417 13091 26483 13094
rect 27613 13154 27679 13157
rect 29177 13154 29243 13157
rect 30281 13154 30347 13157
rect 27613 13152 30347 13154
rect 27613 13096 27618 13152
rect 27674 13096 29182 13152
rect 29238 13096 30286 13152
rect 30342 13096 30347 13152
rect 27613 13094 30347 13096
rect 27613 13091 27679 13094
rect 29177 13091 29243 13094
rect 30281 13091 30347 13094
rect 26980 13088 27296 13089
rect 26980 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27296 13088
rect 26980 13023 27296 13024
rect 20253 13018 20319 13021
rect 20662 13018 20668 13020
rect 20253 13016 20668 13018
rect 20253 12960 20258 13016
rect 20314 12960 20668 13016
rect 20253 12958 20668 12960
rect 20253 12955 20319 12958
rect 20662 12956 20668 12958
rect 20732 13018 20738 13020
rect 24485 13018 24551 13021
rect 20732 13016 24551 13018
rect 20732 12960 24490 13016
rect 24546 12960 24551 13016
rect 20732 12958 24551 12960
rect 20732 12956 20738 12958
rect 24485 12955 24551 12958
rect 24945 13018 25011 13021
rect 25129 13018 25195 13021
rect 24945 13016 25195 13018
rect 24945 12960 24950 13016
rect 25006 12960 25134 13016
rect 25190 12960 25195 13016
rect 24945 12958 25195 12960
rect 24945 12955 25011 12958
rect 25129 12955 25195 12958
rect 25262 12956 25268 13020
rect 25332 13018 25338 13020
rect 26325 13018 26391 13021
rect 25332 13016 26391 13018
rect 25332 12960 26330 13016
rect 26386 12960 26391 13016
rect 25332 12958 26391 12960
rect 25332 12956 25338 12958
rect 26325 12955 26391 12958
rect 21081 12884 21147 12885
rect 21030 12882 21036 12884
rect 18340 12822 19672 12882
rect 20990 12822 21036 12882
rect 21100 12880 21147 12884
rect 21142 12824 21147 12880
rect 18340 12820 18346 12822
rect 21030 12820 21036 12822
rect 21100 12820 21147 12824
rect 21081 12819 21147 12820
rect 21541 12882 21607 12885
rect 22185 12884 22251 12885
rect 21950 12882 21956 12884
rect 21541 12880 21956 12882
rect 21541 12824 21546 12880
rect 21602 12824 21956 12880
rect 21541 12822 21956 12824
rect 21541 12819 21607 12822
rect 21950 12820 21956 12822
rect 22020 12820 22026 12884
rect 22134 12820 22140 12884
rect 22204 12882 22251 12884
rect 22645 12882 22711 12885
rect 26734 12882 26740 12884
rect 22204 12880 22296 12882
rect 22246 12824 22296 12880
rect 22204 12822 22296 12824
rect 22645 12880 26740 12882
rect 22645 12824 22650 12880
rect 22706 12824 26740 12880
rect 22645 12822 26740 12824
rect 22204 12820 22251 12822
rect 22185 12819 22251 12820
rect 22645 12819 22711 12822
rect 26734 12820 26740 12822
rect 26804 12820 26810 12884
rect 26969 12882 27035 12885
rect 29821 12882 29887 12885
rect 26969 12880 29887 12882
rect 26969 12824 26974 12880
rect 27030 12824 29826 12880
rect 29882 12824 29887 12880
rect 26969 12822 29887 12824
rect 26969 12819 27035 12822
rect 29821 12819 29887 12822
rect 6269 12746 6335 12749
rect 6545 12748 6611 12749
rect 2270 12744 6335 12746
rect 2270 12688 6274 12744
rect 6330 12688 6335 12744
rect 2270 12686 6335 12688
rect 2129 12610 2195 12613
rect 2270 12610 2330 12686
rect 6269 12683 6335 12686
rect 6494 12684 6500 12748
rect 6564 12746 6611 12748
rect 6729 12746 6795 12749
rect 8569 12746 8635 12749
rect 13169 12746 13235 12749
rect 13537 12748 13603 12749
rect 6564 12744 6656 12746
rect 6606 12688 6656 12744
rect 6564 12686 6656 12688
rect 6729 12744 8402 12746
rect 6729 12688 6734 12744
rect 6790 12688 8402 12744
rect 6729 12686 8402 12688
rect 6564 12684 6611 12686
rect 6545 12683 6611 12684
rect 6729 12683 6795 12686
rect 2129 12608 2330 12610
rect 2129 12552 2134 12608
rect 2190 12552 2330 12608
rect 2129 12550 2330 12552
rect 6361 12610 6427 12613
rect 6545 12610 6611 12613
rect 6361 12608 6611 12610
rect 6361 12552 6366 12608
rect 6422 12552 6550 12608
rect 6606 12552 6611 12608
rect 6361 12550 6611 12552
rect 2129 12547 2195 12550
rect 6361 12547 6427 12550
rect 6545 12547 6611 12550
rect 7782 12548 7788 12612
rect 7852 12610 7858 12612
rect 7925 12610 7991 12613
rect 7852 12608 7991 12610
rect 7852 12552 7930 12608
rect 7986 12552 7991 12608
rect 7852 12550 7991 12552
rect 8342 12610 8402 12686
rect 8569 12744 13235 12746
rect 8569 12688 8574 12744
rect 8630 12688 13174 12744
rect 13230 12688 13235 12744
rect 8569 12686 13235 12688
rect 8569 12683 8635 12686
rect 13169 12683 13235 12686
rect 13486 12684 13492 12748
rect 13556 12746 13603 12748
rect 14089 12746 14155 12749
rect 14958 12746 14964 12748
rect 13556 12744 13648 12746
rect 13598 12688 13648 12744
rect 13556 12686 13648 12688
rect 14089 12744 14964 12746
rect 14089 12688 14094 12744
rect 14150 12688 14964 12744
rect 14089 12686 14964 12688
rect 13556 12684 13603 12686
rect 13537 12683 13603 12684
rect 14089 12683 14155 12686
rect 14958 12684 14964 12686
rect 15028 12684 15034 12748
rect 15653 12746 15719 12749
rect 15878 12746 15884 12748
rect 15653 12744 15884 12746
rect 15653 12688 15658 12744
rect 15714 12688 15884 12744
rect 15653 12686 15884 12688
rect 15653 12683 15719 12686
rect 15878 12684 15884 12686
rect 15948 12684 15954 12748
rect 16113 12746 16179 12749
rect 16113 12744 17970 12746
rect 16113 12688 16118 12744
rect 16174 12688 17970 12744
rect 16113 12686 17970 12688
rect 16113 12683 16179 12686
rect 11053 12610 11119 12613
rect 11329 12612 11395 12613
rect 11278 12610 11284 12612
rect 8342 12608 11119 12610
rect 8342 12552 11058 12608
rect 11114 12552 11119 12608
rect 8342 12550 11119 12552
rect 11238 12550 11284 12610
rect 11348 12608 11395 12612
rect 11390 12552 11395 12608
rect 7852 12548 7858 12550
rect 7925 12547 7991 12550
rect 11053 12547 11119 12550
rect 11278 12548 11284 12550
rect 11348 12548 11395 12552
rect 11329 12547 11395 12548
rect 12893 12610 12959 12613
rect 14825 12610 14891 12613
rect 12893 12608 14891 12610
rect 12893 12552 12898 12608
rect 12954 12552 14830 12608
rect 14886 12552 14891 12608
rect 12893 12550 14891 12552
rect 12893 12547 12959 12550
rect 14825 12547 14891 12550
rect 16062 12548 16068 12612
rect 16132 12610 16138 12612
rect 17033 12610 17099 12613
rect 16132 12608 17099 12610
rect 16132 12552 17038 12608
rect 17094 12552 17099 12608
rect 16132 12550 17099 12552
rect 17910 12610 17970 12686
rect 18454 12684 18460 12748
rect 18524 12746 18530 12748
rect 19425 12746 19491 12749
rect 18524 12744 19491 12746
rect 18524 12688 19430 12744
rect 19486 12688 19491 12744
rect 18524 12686 19491 12688
rect 18524 12684 18530 12686
rect 19425 12683 19491 12686
rect 19793 12746 19859 12749
rect 28073 12746 28139 12749
rect 28901 12746 28967 12749
rect 19793 12744 28967 12746
rect 19793 12688 19798 12744
rect 19854 12688 28078 12744
rect 28134 12688 28906 12744
rect 28962 12688 28967 12744
rect 19793 12686 28967 12688
rect 19793 12683 19859 12686
rect 28073 12683 28139 12686
rect 28901 12683 28967 12686
rect 19701 12610 19767 12613
rect 17910 12608 19767 12610
rect 17910 12552 19706 12608
rect 19762 12552 19767 12608
rect 17910 12550 19767 12552
rect 16132 12548 16138 12550
rect 17033 12547 17099 12550
rect 19701 12547 19767 12550
rect 20529 12610 20595 12613
rect 22369 12610 22435 12613
rect 20529 12608 22435 12610
rect 20529 12552 20534 12608
rect 20590 12552 22374 12608
rect 22430 12552 22435 12608
rect 20529 12550 22435 12552
rect 20529 12547 20595 12550
rect 22369 12547 22435 12550
rect 23657 12610 23723 12613
rect 26693 12610 26759 12613
rect 23657 12608 26759 12610
rect 23657 12552 23662 12608
rect 23718 12552 26698 12608
rect 26754 12552 26759 12608
rect 23657 12550 26759 12552
rect 23657 12547 23723 12550
rect 26693 12547 26759 12550
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 12092 12544 12408 12545
rect 12092 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12408 12544
rect 12092 12479 12408 12480
rect 19866 12544 20182 12545
rect 19866 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20182 12544
rect 19866 12479 20182 12480
rect 27640 12544 27956 12545
rect 27640 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27956 12544
rect 27640 12479 27956 12480
rect 11145 12474 11211 12477
rect 4846 12472 11211 12474
rect 4846 12416 11150 12472
rect 11206 12416 11211 12472
rect 4846 12414 11211 12416
rect 4846 12341 4906 12414
rect 11145 12411 11211 12414
rect 12934 12412 12940 12476
rect 13004 12474 13010 12476
rect 19517 12474 19583 12477
rect 13004 12472 19583 12474
rect 13004 12416 19522 12472
rect 19578 12416 19583 12472
rect 13004 12414 19583 12416
rect 13004 12412 13010 12414
rect 19517 12411 19583 12414
rect 20437 12474 20503 12477
rect 29177 12474 29243 12477
rect 29494 12474 29500 12476
rect 20437 12472 27538 12474
rect 20437 12416 20442 12472
rect 20498 12416 27538 12472
rect 20437 12414 27538 12416
rect 20437 12411 20503 12414
rect 4797 12336 4906 12341
rect 4797 12280 4802 12336
rect 4858 12280 4906 12336
rect 4797 12278 4906 12280
rect 5993 12338 6059 12341
rect 14733 12338 14799 12341
rect 5993 12336 14799 12338
rect 5993 12280 5998 12336
rect 6054 12280 14738 12336
rect 14794 12280 14799 12336
rect 5993 12278 14799 12280
rect 4797 12275 4863 12278
rect 5993 12275 6059 12278
rect 14733 12275 14799 12278
rect 14958 12276 14964 12340
rect 15028 12338 15034 12340
rect 15285 12338 15351 12341
rect 17585 12338 17651 12341
rect 20989 12338 21055 12341
rect 15028 12278 15210 12338
rect 15028 12276 15034 12278
rect 1669 12202 1735 12205
rect 5625 12202 5691 12205
rect 7189 12202 7255 12205
rect 1669 12200 4952 12202
rect 1669 12144 1674 12200
rect 1730 12144 4952 12200
rect 1669 12142 4952 12144
rect 1669 12139 1735 12142
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 1577 11930 1643 11933
rect 1534 11928 1643 11930
rect 1534 11872 1582 11928
rect 1638 11872 1643 11928
rect 1534 11867 1643 11872
rect 4892 11930 4952 12142
rect 5625 12200 7255 12202
rect 5625 12144 5630 12200
rect 5686 12144 7194 12200
rect 7250 12144 7255 12200
rect 5625 12142 7255 12144
rect 5625 12139 5691 12142
rect 7189 12139 7255 12142
rect 7414 12140 7420 12204
rect 7484 12202 7490 12204
rect 7484 12142 8218 12202
rect 7484 12140 7490 12142
rect 6177 12066 6243 12069
rect 7925 12066 7991 12069
rect 8158 12068 8218 12142
rect 8886 12140 8892 12204
rect 8956 12202 8962 12204
rect 9121 12202 9187 12205
rect 8956 12200 9187 12202
rect 8956 12144 9126 12200
rect 9182 12144 9187 12200
rect 8956 12142 9187 12144
rect 8956 12140 8962 12142
rect 9121 12139 9187 12142
rect 9305 12202 9371 12205
rect 9990 12202 9996 12204
rect 9305 12200 9996 12202
rect 9305 12144 9310 12200
rect 9366 12144 9996 12200
rect 9305 12142 9996 12144
rect 9305 12139 9371 12142
rect 9990 12140 9996 12142
rect 10060 12202 10066 12204
rect 12065 12202 12131 12205
rect 13629 12202 13695 12205
rect 10060 12142 11898 12202
rect 10060 12140 10066 12142
rect 6177 12064 7991 12066
rect 6177 12008 6182 12064
rect 6238 12008 7930 12064
rect 7986 12008 7991 12064
rect 6177 12006 7991 12008
rect 6177 12003 6243 12006
rect 7925 12003 7991 12006
rect 8150 12004 8156 12068
rect 8220 12066 8226 12068
rect 8937 12066 9003 12069
rect 9121 12068 9187 12069
rect 8220 12064 9003 12066
rect 8220 12008 8942 12064
rect 8998 12008 9003 12064
rect 8220 12006 9003 12008
rect 8220 12004 8226 12006
rect 8937 12003 9003 12006
rect 9070 12004 9076 12068
rect 9140 12066 9187 12068
rect 9397 12066 9463 12069
rect 10133 12066 10199 12069
rect 9140 12064 9232 12066
rect 9182 12008 9232 12064
rect 9140 12006 9232 12008
rect 9397 12064 10199 12066
rect 9397 12008 9402 12064
rect 9458 12008 10138 12064
rect 10194 12008 10199 12064
rect 9397 12006 10199 12008
rect 9140 12004 9187 12006
rect 9121 12003 9187 12004
rect 9397 12003 9463 12006
rect 10133 12003 10199 12006
rect 10542 12004 10548 12068
rect 10612 12066 10618 12068
rect 10685 12066 10751 12069
rect 10612 12064 10751 12066
rect 10612 12008 10690 12064
rect 10746 12008 10751 12064
rect 10612 12006 10751 12008
rect 10612 12004 10618 12006
rect 10685 12003 10751 12006
rect 10869 12068 10935 12069
rect 10869 12064 10916 12068
rect 10980 12066 10986 12068
rect 11838 12066 11898 12142
rect 12065 12200 13695 12202
rect 12065 12144 12070 12200
rect 12126 12144 13634 12200
rect 13690 12144 13695 12200
rect 12065 12142 13695 12144
rect 12065 12139 12131 12142
rect 13629 12139 13695 12142
rect 14181 12202 14247 12205
rect 14958 12202 14964 12204
rect 14181 12200 14964 12202
rect 14181 12144 14186 12200
rect 14242 12144 14964 12200
rect 14181 12142 14964 12144
rect 14181 12139 14247 12142
rect 14958 12140 14964 12142
rect 15028 12140 15034 12204
rect 15150 12202 15210 12278
rect 15285 12336 17096 12338
rect 15285 12280 15290 12336
rect 15346 12280 17096 12336
rect 15285 12278 17096 12280
rect 15285 12275 15351 12278
rect 17036 12205 17096 12278
rect 17585 12336 21055 12338
rect 17585 12280 17590 12336
rect 17646 12280 20994 12336
rect 21050 12280 21055 12336
rect 17585 12278 21055 12280
rect 17585 12275 17651 12278
rect 20989 12275 21055 12278
rect 22185 12338 22251 12341
rect 24577 12338 24643 12341
rect 22185 12336 24643 12338
rect 22185 12280 22190 12336
rect 22246 12280 24582 12336
rect 24638 12280 24643 12336
rect 22185 12278 24643 12280
rect 22185 12275 22251 12278
rect 24577 12275 24643 12278
rect 25773 12338 25839 12341
rect 25998 12338 26004 12340
rect 25773 12336 26004 12338
rect 25773 12280 25778 12336
rect 25834 12280 26004 12336
rect 25773 12278 26004 12280
rect 25773 12275 25839 12278
rect 25998 12276 26004 12278
rect 26068 12276 26074 12340
rect 26141 12338 26207 12341
rect 27153 12338 27219 12341
rect 26141 12336 27219 12338
rect 26141 12280 26146 12336
rect 26202 12280 27158 12336
rect 27214 12280 27219 12336
rect 26141 12278 27219 12280
rect 27478 12338 27538 12414
rect 29177 12472 29500 12474
rect 29177 12416 29182 12472
rect 29238 12416 29500 12472
rect 29177 12414 29500 12416
rect 29177 12411 29243 12414
rect 29494 12412 29500 12414
rect 29564 12412 29570 12476
rect 27981 12338 28047 12341
rect 29085 12340 29151 12341
rect 29085 12338 29132 12340
rect 27478 12336 28047 12338
rect 27478 12280 27986 12336
rect 28042 12280 28047 12336
rect 27478 12278 28047 12280
rect 29040 12336 29132 12338
rect 29040 12280 29090 12336
rect 29040 12278 29132 12280
rect 26141 12275 26207 12278
rect 27153 12275 27219 12278
rect 27981 12275 28047 12278
rect 29085 12276 29132 12278
rect 29196 12276 29202 12340
rect 29085 12275 29151 12276
rect 15150 12142 16590 12202
rect 16113 12066 16179 12069
rect 10869 12008 10874 12064
rect 10869 12004 10916 12008
rect 10980 12006 11026 12066
rect 11838 12064 16179 12066
rect 11838 12008 16118 12064
rect 16174 12008 16179 12064
rect 11838 12006 16179 12008
rect 10980 12004 10986 12006
rect 10869 12003 10935 12004
rect 16113 12003 16179 12006
rect 11432 12000 11748 12001
rect 11432 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11748 12000
rect 11432 11935 11748 11936
rect 7414 11930 7420 11932
rect 4892 11870 7420 11930
rect 7414 11868 7420 11870
rect 7484 11868 7490 11932
rect 7782 11868 7788 11932
rect 7852 11930 7858 11932
rect 10961 11930 11027 11933
rect 7852 11928 11027 11930
rect 7852 11872 10966 11928
rect 11022 11872 11027 11928
rect 7852 11870 11027 11872
rect 7852 11868 7858 11870
rect 10961 11867 11027 11870
rect 12525 11930 12591 11933
rect 12801 11930 12867 11933
rect 15929 11930 15995 11933
rect 12525 11928 15995 11930
rect 12525 11872 12530 11928
rect 12586 11872 12806 11928
rect 12862 11872 15934 11928
rect 15990 11872 15995 11928
rect 12525 11870 15995 11872
rect 16530 11930 16590 12142
rect 17033 12200 17099 12205
rect 17033 12144 17038 12200
rect 17094 12144 17099 12200
rect 17033 12139 17099 12144
rect 17902 12140 17908 12204
rect 17972 12202 17978 12204
rect 24025 12202 24091 12205
rect 26417 12202 26483 12205
rect 26785 12202 26851 12205
rect 27613 12202 27679 12205
rect 17972 12200 26664 12202
rect 17972 12144 24030 12200
rect 24086 12144 26422 12200
rect 26478 12144 26664 12200
rect 17972 12142 26664 12144
rect 17972 12140 17978 12142
rect 24025 12139 24091 12142
rect 26417 12139 26483 12142
rect 17217 12066 17283 12069
rect 18781 12066 18847 12069
rect 17217 12064 18847 12066
rect 17217 12008 17222 12064
rect 17278 12008 18786 12064
rect 18842 12008 18847 12064
rect 17217 12006 18847 12008
rect 17217 12003 17283 12006
rect 18781 12003 18847 12006
rect 20437 12066 20503 12069
rect 24945 12066 25011 12069
rect 20437 12064 25011 12066
rect 20437 12008 20442 12064
rect 20498 12008 24950 12064
rect 25006 12008 25011 12064
rect 20437 12006 25011 12008
rect 20437 12003 20503 12006
rect 24945 12003 25011 12006
rect 25497 12066 25563 12069
rect 25630 12066 25636 12068
rect 25497 12064 25636 12066
rect 25497 12008 25502 12064
rect 25558 12008 25636 12064
rect 25497 12006 25636 12008
rect 25497 12003 25563 12006
rect 25630 12004 25636 12006
rect 25700 12004 25706 12068
rect 19206 12000 19522 12001
rect 19206 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19522 12000
rect 19206 11935 19522 11936
rect 18689 11930 18755 11933
rect 20529 11932 20595 11933
rect 20478 11930 20484 11932
rect 16530 11928 18755 11930
rect 16530 11872 18694 11928
rect 18750 11872 18755 11928
rect 16530 11870 18755 11872
rect 20438 11870 20484 11930
rect 20548 11928 20595 11932
rect 20590 11872 20595 11928
rect 12525 11867 12591 11870
rect 12801 11867 12867 11870
rect 15929 11867 15995 11870
rect 18689 11867 18755 11870
rect 20478 11868 20484 11870
rect 20548 11868 20595 11872
rect 21950 11868 21956 11932
rect 22020 11930 22026 11932
rect 26325 11930 26391 11933
rect 22020 11928 26391 11930
rect 22020 11872 26330 11928
rect 26386 11872 26391 11928
rect 22020 11870 26391 11872
rect 22020 11868 22026 11870
rect 20529 11867 20595 11868
rect 26325 11867 26391 11870
rect 1534 11522 1594 11867
rect 2957 11794 3023 11797
rect 11697 11794 11763 11797
rect 2270 11792 11763 11794
rect 2270 11736 2962 11792
rect 3018 11736 11702 11792
rect 11758 11736 11763 11792
rect 2270 11734 11763 11736
rect 2270 11661 2330 11734
rect 2957 11731 3023 11734
rect 11697 11731 11763 11734
rect 12157 11794 12223 11797
rect 15101 11794 15167 11797
rect 12157 11792 15167 11794
rect 12157 11736 12162 11792
rect 12218 11736 15106 11792
rect 15162 11736 15167 11792
rect 12157 11734 15167 11736
rect 12157 11731 12223 11734
rect 15101 11731 15167 11734
rect 15510 11732 15516 11796
rect 15580 11794 15586 11796
rect 15745 11794 15811 11797
rect 15580 11792 15811 11794
rect 15580 11736 15750 11792
rect 15806 11736 15811 11792
rect 15580 11734 15811 11736
rect 15580 11732 15586 11734
rect 15745 11731 15811 11734
rect 18689 11794 18755 11797
rect 18822 11794 18828 11796
rect 18689 11792 18828 11794
rect 18689 11736 18694 11792
rect 18750 11736 18828 11792
rect 18689 11734 18828 11736
rect 18689 11731 18755 11734
rect 18822 11732 18828 11734
rect 18892 11732 18898 11796
rect 19517 11794 19583 11797
rect 21214 11794 21220 11796
rect 19517 11792 21220 11794
rect 19517 11736 19522 11792
rect 19578 11736 21220 11792
rect 19517 11734 21220 11736
rect 19517 11731 19583 11734
rect 21214 11732 21220 11734
rect 21284 11794 21290 11796
rect 25313 11794 25379 11797
rect 21284 11792 25379 11794
rect 21284 11736 25318 11792
rect 25374 11736 25379 11792
rect 21284 11734 25379 11736
rect 26604 11794 26664 12142
rect 26785 12200 27679 12202
rect 26785 12144 26790 12200
rect 26846 12144 27618 12200
rect 27674 12144 27679 12200
rect 26785 12142 27679 12144
rect 26785 12139 26851 12142
rect 27613 12139 27679 12142
rect 26980 12000 27296 12001
rect 26980 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27296 12000
rect 26980 11935 27296 11936
rect 27705 11930 27771 11933
rect 28022 11930 28028 11932
rect 27705 11928 28028 11930
rect 27705 11872 27710 11928
rect 27766 11872 28028 11928
rect 27705 11870 28028 11872
rect 27705 11867 27771 11870
rect 28022 11868 28028 11870
rect 28092 11930 28098 11932
rect 29269 11930 29335 11933
rect 30649 11930 30715 11933
rect 28092 11928 30715 11930
rect 28092 11872 29274 11928
rect 29330 11872 30654 11928
rect 30710 11872 30715 11928
rect 28092 11870 30715 11872
rect 28092 11868 28098 11870
rect 29269 11867 29335 11870
rect 30649 11867 30715 11870
rect 28390 11794 28396 11796
rect 26604 11734 28396 11794
rect 21284 11732 21290 11734
rect 25313 11731 25379 11734
rect 28390 11732 28396 11734
rect 28460 11732 28466 11796
rect 2221 11656 2330 11661
rect 2221 11600 2226 11656
rect 2282 11600 2330 11656
rect 2221 11598 2330 11600
rect 2405 11658 2471 11661
rect 9765 11658 9831 11661
rect 13169 11658 13235 11661
rect 25773 11658 25839 11661
rect 2405 11656 9831 11658
rect 2405 11600 2410 11656
rect 2466 11600 9770 11656
rect 9826 11600 9831 11656
rect 2405 11598 9831 11600
rect 2221 11595 2287 11598
rect 2405 11595 2471 11598
rect 9765 11595 9831 11598
rect 11884 11598 12864 11658
rect 1669 11522 1735 11525
rect 1534 11520 1735 11522
rect 1534 11464 1674 11520
rect 1730 11464 1735 11520
rect 1534 11462 1735 11464
rect 1669 11459 1735 11462
rect 2313 11522 2379 11525
rect 4153 11522 4219 11525
rect 2313 11520 4219 11522
rect 2313 11464 2318 11520
rect 2374 11464 4158 11520
rect 4214 11464 4219 11520
rect 2313 11462 4219 11464
rect 2313 11459 2379 11462
rect 4153 11459 4219 11462
rect 5165 11522 5231 11525
rect 7833 11522 7899 11525
rect 5165 11520 7899 11522
rect 5165 11464 5170 11520
rect 5226 11464 7838 11520
rect 7894 11464 7899 11520
rect 5165 11462 7899 11464
rect 5165 11459 5231 11462
rect 7833 11459 7899 11462
rect 8518 11460 8524 11524
rect 8588 11522 8594 11524
rect 8845 11522 8911 11525
rect 11884 11522 11944 11598
rect 8588 11520 11944 11522
rect 8588 11464 8850 11520
rect 8906 11464 11944 11520
rect 8588 11462 11944 11464
rect 8588 11460 8594 11462
rect 8845 11459 8911 11462
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 12092 11456 12408 11457
rect 12092 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12408 11456
rect 12092 11391 12408 11392
rect 2773 11386 2839 11389
rect 3509 11386 3575 11389
rect 8017 11386 8083 11389
rect 11881 11386 11947 11389
rect 2773 11384 3575 11386
rect 2773 11328 2778 11384
rect 2834 11328 3514 11384
rect 3570 11328 3575 11384
rect 2773 11326 3575 11328
rect 2773 11323 2839 11326
rect 3509 11323 3575 11326
rect 5766 11384 11947 11386
rect 5766 11328 8022 11384
rect 8078 11328 11886 11384
rect 11942 11328 11947 11384
rect 5766 11326 11947 11328
rect 2957 11252 3023 11253
rect 2957 11250 3004 11252
rect 2912 11248 3004 11250
rect 2912 11192 2962 11248
rect 2912 11190 3004 11192
rect 2957 11188 3004 11190
rect 3068 11188 3074 11252
rect 3366 11188 3372 11252
rect 3436 11250 3442 11252
rect 5766 11250 5826 11326
rect 8017 11323 8083 11326
rect 11881 11323 11947 11326
rect 3436 11190 5826 11250
rect 7005 11250 7071 11253
rect 10225 11250 10291 11253
rect 7005 11248 10291 11250
rect 7005 11192 7010 11248
rect 7066 11192 10230 11248
rect 10286 11192 10291 11248
rect 7005 11190 10291 11192
rect 3436 11188 3442 11190
rect 2957 11187 3023 11188
rect 7005 11187 7071 11190
rect 10225 11187 10291 11190
rect 10542 11188 10548 11252
rect 10612 11250 10618 11252
rect 10777 11250 10843 11253
rect 10612 11248 10843 11250
rect 10612 11192 10782 11248
rect 10838 11192 10843 11248
rect 10612 11190 10843 11192
rect 10612 11188 10618 11190
rect 10777 11187 10843 11190
rect 11094 11188 11100 11252
rect 11164 11250 11170 11252
rect 12566 11250 12572 11252
rect 11164 11190 12572 11250
rect 11164 11188 11170 11190
rect 12566 11188 12572 11190
rect 12636 11188 12642 11252
rect 12804 11250 12864 11598
rect 13169 11656 25839 11658
rect 13169 11600 13174 11656
rect 13230 11600 25778 11656
rect 25834 11600 25839 11656
rect 13169 11598 25839 11600
rect 13169 11595 13235 11598
rect 25773 11595 25839 11598
rect 25957 11658 26023 11661
rect 27613 11658 27679 11661
rect 25957 11656 27679 11658
rect 25957 11600 25962 11656
rect 26018 11600 27618 11656
rect 27674 11600 27679 11656
rect 25957 11598 27679 11600
rect 25957 11595 26023 11598
rect 27613 11595 27679 11598
rect 27797 11658 27863 11661
rect 28165 11658 28231 11661
rect 27797 11656 28231 11658
rect 27797 11600 27802 11656
rect 27858 11600 28170 11656
rect 28226 11600 28231 11656
rect 27797 11598 28231 11600
rect 27797 11595 27863 11598
rect 28165 11595 28231 11598
rect 14038 11460 14044 11524
rect 14108 11522 14114 11524
rect 14273 11522 14339 11525
rect 14108 11520 14339 11522
rect 14108 11464 14278 11520
rect 14334 11464 14339 11520
rect 14108 11462 14339 11464
rect 14108 11460 14114 11462
rect 14273 11459 14339 11462
rect 19517 11522 19583 11525
rect 19696 11522 19702 11524
rect 19517 11520 19702 11522
rect 19517 11464 19522 11520
rect 19578 11464 19702 11520
rect 19517 11462 19702 11464
rect 19517 11459 19583 11462
rect 19696 11460 19702 11462
rect 19766 11460 19772 11524
rect 20662 11460 20668 11524
rect 20732 11522 20738 11524
rect 22737 11522 22803 11525
rect 20732 11520 22803 11522
rect 20732 11464 22742 11520
rect 22798 11464 22803 11520
rect 20732 11462 22803 11464
rect 20732 11460 20738 11462
rect 22737 11459 22803 11462
rect 22870 11460 22876 11524
rect 22940 11522 22946 11524
rect 23105 11522 23171 11525
rect 22940 11520 23171 11522
rect 22940 11464 23110 11520
rect 23166 11464 23171 11520
rect 22940 11462 23171 11464
rect 22940 11460 22946 11462
rect 23105 11459 23171 11462
rect 23933 11522 23999 11525
rect 24393 11522 24459 11525
rect 23933 11520 24459 11522
rect 23933 11464 23938 11520
rect 23994 11464 24398 11520
rect 24454 11464 24459 11520
rect 23933 11462 24459 11464
rect 23933 11459 23999 11462
rect 24393 11459 24459 11462
rect 25405 11522 25471 11525
rect 25773 11522 25839 11525
rect 25405 11520 25839 11522
rect 25405 11464 25410 11520
rect 25466 11464 25778 11520
rect 25834 11464 25839 11520
rect 25405 11462 25839 11464
rect 25405 11459 25471 11462
rect 25773 11459 25839 11462
rect 26182 11460 26188 11524
rect 26252 11522 26258 11524
rect 26325 11522 26391 11525
rect 26252 11520 26391 11522
rect 26252 11464 26330 11520
rect 26386 11464 26391 11520
rect 26252 11462 26391 11464
rect 26252 11460 26258 11462
rect 26325 11459 26391 11462
rect 19866 11456 20182 11457
rect 19866 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20182 11456
rect 19866 11391 20182 11392
rect 27640 11456 27956 11457
rect 27640 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27956 11456
rect 27640 11391 27956 11392
rect 12985 11386 13051 11389
rect 15510 11386 15516 11388
rect 12985 11384 15516 11386
rect 12985 11328 12990 11384
rect 13046 11328 15516 11384
rect 12985 11326 15516 11328
rect 12985 11323 13051 11326
rect 15510 11324 15516 11326
rect 15580 11324 15586 11388
rect 16430 11324 16436 11388
rect 16500 11386 16506 11388
rect 16573 11386 16639 11389
rect 25129 11386 25195 11389
rect 16500 11384 19764 11386
rect 16500 11328 16578 11384
rect 16634 11352 19764 11384
rect 20256 11384 25195 11386
rect 16634 11328 19810 11352
rect 16500 11326 19810 11328
rect 16500 11324 16506 11326
rect 16573 11323 16639 11326
rect 19704 11292 19810 11326
rect 19750 11284 19810 11292
rect 20256 11328 25134 11384
rect 25190 11328 25195 11384
rect 20256 11326 25195 11328
rect 14365 11250 14431 11253
rect 14590 11250 14596 11252
rect 12804 11190 13186 11250
rect 1117 11114 1183 11117
rect 4613 11114 4679 11117
rect 1117 11112 4679 11114
rect 1117 11056 1122 11112
rect 1178 11056 4618 11112
rect 4674 11056 4679 11112
rect 1117 11054 4679 11056
rect 1117 11051 1183 11054
rect 4613 11051 4679 11054
rect 6637 11116 6703 11117
rect 9121 11116 9187 11117
rect 6637 11112 6684 11116
rect 6748 11114 6754 11116
rect 9070 11114 9076 11116
rect 6637 11056 6642 11112
rect 6637 11052 6684 11056
rect 6748 11054 6794 11114
rect 9030 11054 9076 11114
rect 9140 11112 9187 11116
rect 11605 11114 11671 11117
rect 9182 11056 9187 11112
rect 6748 11052 6754 11054
rect 9070 11052 9076 11054
rect 9140 11052 9187 11056
rect 6637 11051 6703 11052
rect 9121 11051 9187 11052
rect 9308 11112 11671 11114
rect 9308 11056 11610 11112
rect 11666 11056 11671 11112
rect 9308 11054 11671 11056
rect 4705 10978 4771 10981
rect 4838 10978 4844 10980
rect 4705 10976 4844 10978
rect 4705 10920 4710 10976
rect 4766 10920 4844 10976
rect 4705 10918 4844 10920
rect 4705 10915 4771 10918
rect 4838 10916 4844 10918
rect 4908 10916 4914 10980
rect 5717 10978 5783 10981
rect 8017 10978 8083 10981
rect 5717 10976 8083 10978
rect 5717 10920 5722 10976
rect 5778 10920 8022 10976
rect 8078 10920 8083 10976
rect 5717 10918 8083 10920
rect 5717 10915 5783 10918
rect 8017 10915 8083 10918
rect 8845 10978 8911 10981
rect 9308 10978 9368 11054
rect 11605 11051 11671 11054
rect 12893 11116 12959 11117
rect 12893 11112 12940 11116
rect 13004 11114 13010 11116
rect 13126 11114 13186 11190
rect 14365 11248 14596 11250
rect 14365 11192 14370 11248
rect 14426 11192 14596 11248
rect 14365 11190 14596 11192
rect 14365 11187 14431 11190
rect 14590 11188 14596 11190
rect 14660 11188 14666 11252
rect 14733 11250 14799 11253
rect 14917 11250 14983 11253
rect 14733 11248 14983 11250
rect 14733 11192 14738 11248
rect 14794 11192 14922 11248
rect 14978 11192 14983 11248
rect 14733 11190 14983 11192
rect 14733 11187 14799 11190
rect 14917 11187 14983 11190
rect 15101 11250 15167 11253
rect 19750 11250 19948 11284
rect 20256 11250 20316 11326
rect 25129 11323 25195 11326
rect 26366 11324 26372 11388
rect 26436 11386 26442 11388
rect 26877 11386 26943 11389
rect 26436 11384 26943 11386
rect 26436 11328 26882 11384
rect 26938 11328 26943 11384
rect 26436 11326 26943 11328
rect 26436 11324 26442 11326
rect 26877 11323 26943 11326
rect 15101 11248 19580 11250
rect 15101 11192 15106 11248
rect 15162 11192 19580 11248
rect 19750 11224 20316 11250
rect 15101 11190 19580 11192
rect 19888 11190 20316 11224
rect 20897 11250 20963 11253
rect 22737 11250 22803 11253
rect 20897 11248 22803 11250
rect 20897 11192 20902 11248
rect 20958 11192 22742 11248
rect 22798 11192 22803 11248
rect 20897 11190 22803 11192
rect 15101 11187 15167 11190
rect 19520 11148 19580 11190
rect 20897 11187 20963 11190
rect 22737 11187 22803 11190
rect 24025 11250 24091 11253
rect 27061 11250 27127 11253
rect 24025 11248 27127 11250
rect 24025 11192 24030 11248
rect 24086 11192 27066 11248
rect 27122 11192 27127 11248
rect 24025 11190 27127 11192
rect 24025 11187 24091 11190
rect 27061 11187 27127 11190
rect 27521 11250 27587 11253
rect 28257 11250 28323 11253
rect 27521 11248 28323 11250
rect 27521 11192 27526 11248
rect 27582 11192 28262 11248
rect 28318 11192 28323 11248
rect 27521 11190 28323 11192
rect 27521 11187 27587 11190
rect 28257 11187 28323 11190
rect 13905 11114 13971 11117
rect 17493 11114 17559 11117
rect 12893 11056 12898 11112
rect 12893 11052 12940 11056
rect 13004 11054 13050 11114
rect 13126 11112 17559 11114
rect 13126 11056 13910 11112
rect 13966 11056 17498 11112
rect 17554 11056 17559 11112
rect 13126 11054 17559 11056
rect 13004 11052 13010 11054
rect 12893 11051 12959 11052
rect 13905 11051 13971 11054
rect 17493 11051 17559 11054
rect 18781 11114 18847 11117
rect 19057 11114 19123 11117
rect 18781 11112 19123 11114
rect 18781 11056 18786 11112
rect 18842 11056 19062 11112
rect 19118 11056 19123 11112
rect 19520 11114 19764 11148
rect 22001 11114 22067 11117
rect 19520 11112 22067 11114
rect 19520 11088 22006 11112
rect 18781 11054 19123 11056
rect 19704 11056 22006 11088
rect 22062 11056 22067 11112
rect 19704 11054 22067 11056
rect 18781 11051 18847 11054
rect 19057 11051 19123 11054
rect 22001 11051 22067 11054
rect 22185 11114 22251 11117
rect 25957 11114 26023 11117
rect 22185 11112 26023 11114
rect 22185 11056 22190 11112
rect 22246 11056 25962 11112
rect 26018 11056 26023 11112
rect 22185 11054 26023 11056
rect 22185 11051 22251 11054
rect 25957 11051 26023 11054
rect 26550 11052 26556 11116
rect 26620 11114 26626 11116
rect 27613 11114 27679 11117
rect 26620 11112 27679 11114
rect 26620 11056 27618 11112
rect 27674 11056 27679 11112
rect 26620 11054 27679 11056
rect 26620 11052 26626 11054
rect 27613 11051 27679 11054
rect 8845 10976 9368 10978
rect 8845 10920 8850 10976
rect 8906 10920 9368 10976
rect 8845 10918 9368 10920
rect 9489 10978 9555 10981
rect 10133 10978 10199 10981
rect 10542 10978 10548 10980
rect 9489 10976 10548 10978
rect 9489 10920 9494 10976
rect 9550 10920 10138 10976
rect 10194 10920 10548 10976
rect 9489 10918 10548 10920
rect 8845 10915 8911 10918
rect 9489 10915 9555 10918
rect 10133 10915 10199 10918
rect 10542 10916 10548 10918
rect 10612 10916 10618 10980
rect 13118 10978 13124 10980
rect 11838 10918 13124 10978
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 11432 10912 11748 10913
rect 11432 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11748 10912
rect 11432 10847 11748 10848
rect 4337 10842 4403 10845
rect 4838 10842 4844 10844
rect 4337 10840 4844 10842
rect 4337 10784 4342 10840
rect 4398 10784 4844 10840
rect 4337 10782 4844 10784
rect 4337 10779 4403 10782
rect 4838 10780 4844 10782
rect 4908 10780 4914 10844
rect 8201 10842 8267 10845
rect 9622 10842 9628 10844
rect 8201 10840 9628 10842
rect 8201 10784 8206 10840
rect 8262 10784 9628 10840
rect 8201 10782 9628 10784
rect 8201 10779 8267 10782
rect 9622 10780 9628 10782
rect 9692 10780 9698 10844
rect 9765 10842 9831 10845
rect 11237 10842 11303 10845
rect 9765 10840 11303 10842
rect 9765 10784 9770 10840
rect 9826 10784 11242 10840
rect 11298 10784 11303 10840
rect 9765 10782 11303 10784
rect 9765 10779 9831 10782
rect 11237 10779 11303 10782
rect 3233 10706 3299 10709
rect 8293 10706 8359 10709
rect 3233 10704 8359 10706
rect 3233 10648 3238 10704
rect 3294 10648 8298 10704
rect 8354 10648 8359 10704
rect 3233 10646 8359 10648
rect 3233 10643 3299 10646
rect 8293 10643 8359 10646
rect 9438 10644 9444 10708
rect 9508 10706 9514 10708
rect 10133 10706 10199 10709
rect 11838 10706 11898 10918
rect 13118 10916 13124 10918
rect 13188 10978 13194 10980
rect 14038 10978 14044 10980
rect 13188 10918 14044 10978
rect 13188 10916 13194 10918
rect 14038 10916 14044 10918
rect 14108 10916 14114 10980
rect 14222 10916 14228 10980
rect 14292 10978 14298 10980
rect 15193 10978 15259 10981
rect 18229 10978 18295 10981
rect 14292 10976 15259 10978
rect 14292 10920 15198 10976
rect 15254 10920 15259 10976
rect 14292 10918 15259 10920
rect 14292 10916 14298 10918
rect 15193 10915 15259 10918
rect 15334 10976 18295 10978
rect 15334 10920 18234 10976
rect 18290 10920 18295 10976
rect 15334 10918 18295 10920
rect 15334 10842 15394 10918
rect 18229 10915 18295 10918
rect 19696 10916 19702 10980
rect 19766 10978 19772 10980
rect 20437 10978 20503 10981
rect 19766 10976 20503 10978
rect 19766 10920 20442 10976
rect 20498 10920 20503 10976
rect 19766 10918 20503 10920
rect 19766 10916 19772 10918
rect 20437 10915 20503 10918
rect 20989 10978 21055 10981
rect 25957 10978 26023 10981
rect 20989 10976 26023 10978
rect 20989 10920 20994 10976
rect 21050 10920 25962 10976
rect 26018 10920 26023 10976
rect 20989 10918 26023 10920
rect 20989 10915 21055 10918
rect 25957 10915 26023 10918
rect 19206 10912 19522 10913
rect 19206 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19522 10912
rect 19206 10847 19522 10848
rect 26980 10912 27296 10913
rect 26980 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27296 10912
rect 26980 10847 27296 10848
rect 9508 10704 11898 10706
rect 9508 10648 10138 10704
rect 10194 10648 11898 10704
rect 9508 10646 11898 10648
rect 11976 10782 15394 10842
rect 15561 10842 15627 10845
rect 16757 10842 16823 10845
rect 15561 10840 16823 10842
rect 15561 10784 15566 10840
rect 15622 10784 16762 10840
rect 16818 10784 16823 10840
rect 15561 10782 16823 10784
rect 9508 10644 9514 10646
rect 10133 10643 10199 10646
rect 2446 10508 2452 10572
rect 2516 10570 2522 10572
rect 3693 10570 3759 10573
rect 6126 10570 6132 10572
rect 2516 10568 6132 10570
rect 2516 10512 3698 10568
rect 3754 10512 6132 10568
rect 2516 10510 6132 10512
rect 2516 10508 2522 10510
rect 3693 10507 3759 10510
rect 6126 10508 6132 10510
rect 6196 10508 6202 10572
rect 9305 10570 9371 10573
rect 9990 10570 9996 10572
rect 6272 10510 7988 10570
rect 6272 10437 6332 10510
rect 5390 10372 5396 10436
rect 5460 10434 5466 10436
rect 5533 10434 5599 10437
rect 5460 10432 5599 10434
rect 5460 10376 5538 10432
rect 5594 10376 5599 10432
rect 5460 10374 5599 10376
rect 5460 10372 5466 10374
rect 5533 10371 5599 10374
rect 5993 10434 6059 10437
rect 6269 10434 6335 10437
rect 7741 10436 7807 10437
rect 7741 10434 7788 10436
rect 5993 10432 6335 10434
rect 5993 10376 5998 10432
rect 6054 10376 6274 10432
rect 6330 10376 6335 10432
rect 5993 10374 6335 10376
rect 7696 10432 7788 10434
rect 7696 10376 7746 10432
rect 7696 10374 7788 10376
rect 5993 10371 6059 10374
rect 6269 10371 6335 10374
rect 7741 10372 7788 10374
rect 7852 10372 7858 10436
rect 7928 10434 7988 10510
rect 9305 10568 9996 10570
rect 9305 10512 9310 10568
rect 9366 10512 9996 10568
rect 9305 10510 9996 10512
rect 9305 10507 9371 10510
rect 9990 10508 9996 10510
rect 10060 10508 10066 10572
rect 10501 10570 10567 10573
rect 11976 10570 12036 10782
rect 15561 10779 15627 10782
rect 16757 10779 16823 10782
rect 20294 10780 20300 10844
rect 20364 10842 20370 10844
rect 22277 10842 22343 10845
rect 20364 10840 22343 10842
rect 20364 10784 22282 10840
rect 22338 10784 22343 10840
rect 20364 10782 22343 10784
rect 20364 10780 20370 10782
rect 22277 10779 22343 10782
rect 24945 10842 25011 10845
rect 25078 10842 25084 10844
rect 24945 10840 25084 10842
rect 24945 10784 24950 10840
rect 25006 10784 25084 10840
rect 24945 10782 25084 10784
rect 24945 10779 25011 10782
rect 25078 10780 25084 10782
rect 25148 10780 25154 10844
rect 12341 10706 12407 10709
rect 14181 10706 14247 10709
rect 12341 10704 14247 10706
rect 12341 10648 12346 10704
rect 12402 10648 14186 10704
rect 14242 10648 14247 10704
rect 12341 10646 14247 10648
rect 12341 10643 12407 10646
rect 14181 10643 14247 10646
rect 14457 10706 14523 10709
rect 15009 10706 15075 10709
rect 14457 10704 15075 10706
rect 14457 10648 14462 10704
rect 14518 10648 15014 10704
rect 15070 10648 15075 10704
rect 14457 10646 15075 10648
rect 14457 10643 14523 10646
rect 15009 10643 15075 10646
rect 15193 10706 15259 10709
rect 18454 10706 18460 10708
rect 15193 10704 18460 10706
rect 15193 10648 15198 10704
rect 15254 10648 18460 10704
rect 15193 10646 18460 10648
rect 15193 10643 15259 10646
rect 18454 10644 18460 10646
rect 18524 10644 18530 10708
rect 19241 10706 19307 10709
rect 30373 10706 30439 10709
rect 19241 10704 30439 10706
rect 19241 10648 19246 10704
rect 19302 10648 30378 10704
rect 30434 10648 30439 10704
rect 19241 10646 30439 10648
rect 19241 10643 19307 10646
rect 30373 10643 30439 10646
rect 10501 10568 12036 10570
rect 10501 10512 10506 10568
rect 10562 10512 12036 10568
rect 10501 10510 12036 10512
rect 12157 10570 12223 10573
rect 19425 10570 19491 10573
rect 12157 10568 19491 10570
rect 12157 10512 12162 10568
rect 12218 10512 19430 10568
rect 19486 10512 19491 10568
rect 12157 10510 19491 10512
rect 10501 10507 10567 10510
rect 12157 10507 12223 10510
rect 19425 10507 19491 10510
rect 19609 10570 19675 10573
rect 21582 10570 21588 10572
rect 19609 10568 21588 10570
rect 19609 10512 19614 10568
rect 19670 10512 21588 10568
rect 19609 10510 21588 10512
rect 19609 10507 19675 10510
rect 21582 10508 21588 10510
rect 21652 10508 21658 10572
rect 22737 10568 22803 10573
rect 22737 10512 22742 10568
rect 22798 10512 22803 10568
rect 22737 10507 22803 10512
rect 23473 10570 23539 10573
rect 23657 10570 23723 10573
rect 30230 10570 30236 10572
rect 23473 10568 23723 10570
rect 23473 10512 23478 10568
rect 23534 10512 23662 10568
rect 23718 10512 23723 10568
rect 23473 10510 23723 10512
rect 23473 10507 23539 10510
rect 23657 10507 23723 10510
rect 23798 10510 30236 10570
rect 11697 10434 11763 10437
rect 7928 10432 11763 10434
rect 7928 10376 11702 10432
rect 11758 10376 11763 10432
rect 7928 10374 11763 10376
rect 7741 10371 7807 10372
rect 11697 10371 11763 10374
rect 13261 10434 13327 10437
rect 14457 10434 14523 10437
rect 13261 10432 14523 10434
rect 13261 10376 13266 10432
rect 13322 10376 14462 10432
rect 14518 10376 14523 10432
rect 13261 10374 14523 10376
rect 13261 10371 13327 10374
rect 14457 10371 14523 10374
rect 14774 10372 14780 10436
rect 14844 10434 14850 10436
rect 15745 10434 15811 10437
rect 14844 10432 15811 10434
rect 14844 10376 15750 10432
rect 15806 10376 15811 10432
rect 14844 10374 15811 10376
rect 14844 10372 14850 10374
rect 15745 10371 15811 10374
rect 15878 10372 15884 10436
rect 15948 10434 15954 10436
rect 18689 10434 18755 10437
rect 15948 10432 18755 10434
rect 15948 10376 18694 10432
rect 18750 10376 18755 10432
rect 15948 10374 18755 10376
rect 15948 10372 15954 10374
rect 18689 10371 18755 10374
rect 19149 10434 19215 10437
rect 19609 10434 19675 10437
rect 19149 10432 19675 10434
rect 19149 10376 19154 10432
rect 19210 10376 19614 10432
rect 19670 10376 19675 10432
rect 19149 10374 19675 10376
rect 19149 10371 19215 10374
rect 19609 10371 19675 10374
rect 20294 10372 20300 10436
rect 20364 10434 20370 10436
rect 20713 10434 20779 10437
rect 20364 10432 20779 10434
rect 20364 10376 20718 10432
rect 20774 10376 20779 10432
rect 20364 10374 20779 10376
rect 20364 10372 20370 10374
rect 20713 10371 20779 10374
rect 21030 10372 21036 10436
rect 21100 10434 21106 10436
rect 21449 10434 21515 10437
rect 21100 10432 21515 10434
rect 21100 10376 21454 10432
rect 21510 10376 21515 10432
rect 21100 10374 21515 10376
rect 22740 10434 22800 10507
rect 23289 10434 23355 10437
rect 23798 10434 23858 10510
rect 30230 10508 30236 10510
rect 30300 10508 30306 10572
rect 22740 10432 23858 10434
rect 22740 10376 23294 10432
rect 23350 10376 23858 10432
rect 22740 10374 23858 10376
rect 25221 10434 25287 10437
rect 27061 10434 27127 10437
rect 25221 10432 27127 10434
rect 25221 10376 25226 10432
rect 25282 10376 27066 10432
rect 27122 10376 27127 10432
rect 25221 10374 27127 10376
rect 21100 10372 21106 10374
rect 21449 10371 21515 10374
rect 23289 10371 23355 10374
rect 25221 10371 25287 10374
rect 27061 10371 27127 10374
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 12092 10368 12408 10369
rect 12092 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12408 10368
rect 12092 10303 12408 10304
rect 19866 10368 20182 10369
rect 19866 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20182 10368
rect 19866 10303 20182 10304
rect 27640 10368 27956 10369
rect 27640 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27956 10368
rect 27640 10303 27956 10304
rect 3785 10298 3851 10301
rect 4102 10298 4108 10300
rect 3785 10296 4108 10298
rect 3785 10240 3790 10296
rect 3846 10240 4108 10296
rect 3785 10238 4108 10240
rect 3785 10235 3851 10238
rect 4102 10236 4108 10238
rect 4172 10236 4178 10300
rect 6177 10298 6243 10301
rect 6310 10298 6316 10300
rect 6177 10296 6316 10298
rect 6177 10240 6182 10296
rect 6238 10240 6316 10296
rect 6177 10238 6316 10240
rect 6177 10235 6243 10238
rect 6310 10236 6316 10238
rect 6380 10236 6386 10300
rect 7833 10298 7899 10301
rect 9121 10298 9187 10301
rect 7833 10296 9187 10298
rect 7833 10240 7838 10296
rect 7894 10240 9126 10296
rect 9182 10240 9187 10296
rect 7833 10238 9187 10240
rect 7833 10235 7899 10238
rect 9121 10235 9187 10238
rect 9397 10298 9463 10301
rect 9581 10298 9647 10301
rect 9397 10296 9647 10298
rect 9397 10240 9402 10296
rect 9458 10240 9586 10296
rect 9642 10240 9647 10296
rect 9397 10238 9647 10240
rect 9397 10235 9463 10238
rect 9581 10235 9647 10238
rect 9990 10236 9996 10300
rect 10060 10298 10066 10300
rect 10593 10298 10659 10301
rect 10060 10296 10659 10298
rect 10060 10240 10598 10296
rect 10654 10240 10659 10296
rect 10060 10238 10659 10240
rect 10060 10236 10066 10238
rect 10593 10235 10659 10238
rect 11278 10236 11284 10300
rect 11348 10298 11354 10300
rect 11605 10298 11671 10301
rect 11348 10296 11671 10298
rect 11348 10240 11610 10296
rect 11666 10240 11671 10296
rect 11348 10238 11671 10240
rect 11348 10236 11354 10238
rect 11605 10235 11671 10238
rect 12985 10298 13051 10301
rect 17534 10298 17540 10300
rect 12985 10296 17540 10298
rect 12985 10240 12990 10296
rect 13046 10240 17540 10296
rect 12985 10238 17540 10240
rect 12985 10235 13051 10238
rect 17534 10236 17540 10238
rect 17604 10236 17610 10300
rect 17769 10298 17835 10301
rect 18321 10298 18387 10301
rect 17769 10296 18387 10298
rect 17769 10240 17774 10296
rect 17830 10240 18326 10296
rect 18382 10240 18387 10296
rect 17769 10238 18387 10240
rect 17769 10235 17835 10238
rect 18321 10235 18387 10238
rect 18822 10236 18828 10300
rect 18892 10298 18898 10300
rect 19333 10298 19399 10301
rect 18892 10296 19399 10298
rect 18892 10240 19338 10296
rect 19394 10240 19399 10296
rect 18892 10238 19399 10240
rect 18892 10236 18898 10238
rect 19333 10235 19399 10238
rect 20713 10298 20779 10301
rect 20897 10298 20963 10301
rect 20713 10296 20963 10298
rect 20713 10240 20718 10296
rect 20774 10240 20902 10296
rect 20958 10240 20963 10296
rect 20713 10238 20963 10240
rect 20713 10235 20779 10238
rect 20897 10235 20963 10238
rect 21398 10236 21404 10300
rect 21468 10298 21474 10300
rect 23013 10298 23079 10301
rect 21468 10296 23079 10298
rect 21468 10240 23018 10296
rect 23074 10240 23079 10296
rect 21468 10238 23079 10240
rect 21468 10236 21474 10238
rect 23013 10235 23079 10238
rect 24894 10236 24900 10300
rect 24964 10298 24970 10300
rect 25405 10298 25471 10301
rect 24964 10296 25471 10298
rect 24964 10240 25410 10296
rect 25466 10240 25471 10296
rect 24964 10238 25471 10240
rect 24964 10236 24970 10238
rect 25405 10235 25471 10238
rect 26325 10298 26391 10301
rect 26969 10298 27035 10301
rect 26325 10296 27035 10298
rect 26325 10240 26330 10296
rect 26386 10240 26974 10296
rect 27030 10240 27035 10296
rect 26325 10238 27035 10240
rect 26325 10235 26391 10238
rect 26969 10235 27035 10238
rect 14222 10162 14228 10164
rect 2730 10102 14228 10162
rect 2497 10026 2563 10029
rect 2730 10026 2790 10102
rect 14222 10100 14228 10102
rect 14292 10100 14298 10164
rect 14733 10162 14799 10165
rect 15142 10162 15148 10164
rect 14733 10160 15148 10162
rect 14733 10104 14738 10160
rect 14794 10104 15148 10160
rect 14733 10102 15148 10104
rect 14733 10099 14799 10102
rect 15142 10100 15148 10102
rect 15212 10100 15218 10164
rect 16757 10162 16823 10165
rect 27981 10162 28047 10165
rect 16757 10160 28047 10162
rect 16757 10104 16762 10160
rect 16818 10104 27986 10160
rect 28042 10104 28047 10160
rect 16757 10102 28047 10104
rect 16757 10099 16823 10102
rect 27981 10099 28047 10102
rect 2497 10024 2790 10026
rect 2497 9968 2502 10024
rect 2558 9968 2790 10024
rect 2497 9966 2790 9968
rect 4245 10026 4311 10029
rect 19885 10026 19951 10029
rect 21909 10026 21975 10029
rect 22645 10026 22711 10029
rect 23105 10026 23171 10029
rect 26601 10026 26667 10029
rect 27613 10026 27679 10029
rect 4245 10024 15210 10026
rect 4245 9968 4250 10024
rect 4306 9968 15210 10024
rect 4245 9966 15210 9968
rect 2497 9963 2563 9966
rect 4245 9963 4311 9966
rect 4337 9890 4403 9893
rect 9254 9890 9260 9892
rect 4337 9888 9260 9890
rect 4337 9832 4342 9888
rect 4398 9832 9260 9888
rect 4337 9830 9260 9832
rect 4337 9827 4403 9830
rect 9254 9828 9260 9830
rect 9324 9828 9330 9892
rect 9673 9890 9739 9893
rect 9806 9890 9812 9892
rect 9673 9888 9812 9890
rect 9673 9832 9678 9888
rect 9734 9832 9812 9888
rect 9673 9830 9812 9832
rect 9673 9827 9739 9830
rect 9806 9828 9812 9830
rect 9876 9828 9882 9892
rect 10133 9890 10199 9893
rect 10358 9890 10364 9892
rect 10133 9888 10364 9890
rect 10133 9832 10138 9888
rect 10194 9832 10364 9888
rect 10133 9830 10364 9832
rect 10133 9827 10199 9830
rect 10358 9828 10364 9830
rect 10428 9890 10434 9892
rect 11094 9890 11100 9892
rect 10428 9830 11100 9890
rect 10428 9828 10434 9830
rect 11094 9828 11100 9830
rect 11164 9828 11170 9892
rect 12566 9828 12572 9892
rect 12636 9890 12642 9892
rect 13854 9890 13860 9892
rect 12636 9830 13860 9890
rect 12636 9828 12642 9830
rect 13854 9828 13860 9830
rect 13924 9828 13930 9892
rect 14273 9890 14339 9893
rect 14590 9890 14596 9892
rect 14273 9888 14596 9890
rect 14273 9832 14278 9888
rect 14334 9832 14596 9888
rect 14273 9830 14596 9832
rect 14273 9827 14339 9830
rect 14590 9828 14596 9830
rect 14660 9828 14666 9892
rect 15150 9890 15210 9966
rect 15288 9966 19764 10026
rect 15288 9890 15348 9966
rect 15150 9830 15348 9890
rect 15510 9828 15516 9892
rect 15580 9890 15586 9892
rect 16021 9890 16087 9893
rect 15580 9888 16087 9890
rect 15580 9832 16026 9888
rect 16082 9832 16087 9888
rect 15580 9830 16087 9832
rect 15580 9828 15586 9830
rect 16021 9827 16087 9830
rect 16297 9890 16363 9893
rect 16614 9890 16620 9892
rect 16297 9888 16620 9890
rect 16297 9832 16302 9888
rect 16358 9832 16620 9888
rect 16297 9830 16620 9832
rect 16297 9827 16363 9830
rect 16614 9828 16620 9830
rect 16684 9828 16690 9892
rect 16849 9890 16915 9893
rect 16982 9890 16988 9892
rect 16849 9888 16988 9890
rect 16849 9832 16854 9888
rect 16910 9832 16988 9888
rect 16849 9830 16988 9832
rect 16849 9827 16915 9830
rect 16982 9828 16988 9830
rect 17052 9890 17058 9892
rect 17769 9890 17835 9893
rect 18229 9892 18295 9893
rect 18229 9890 18276 9892
rect 17052 9888 17835 9890
rect 17052 9832 17774 9888
rect 17830 9832 17835 9888
rect 17052 9830 17835 9832
rect 18184 9888 18276 9890
rect 18184 9832 18234 9888
rect 18184 9830 18276 9832
rect 17052 9828 17058 9830
rect 17769 9827 17835 9830
rect 18229 9828 18276 9830
rect 18340 9828 18346 9892
rect 18229 9827 18295 9828
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 11432 9824 11748 9825
rect 11432 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11748 9824
rect 11432 9759 11748 9760
rect 19206 9824 19522 9825
rect 19206 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19522 9824
rect 19206 9759 19522 9760
rect 5533 9754 5599 9757
rect 5758 9754 5764 9756
rect 5533 9752 5764 9754
rect 5533 9696 5538 9752
rect 5594 9696 5764 9752
rect 5533 9694 5764 9696
rect 5533 9691 5599 9694
rect 5758 9692 5764 9694
rect 5828 9692 5834 9756
rect 7557 9754 7623 9757
rect 7925 9754 7991 9757
rect 10501 9754 10567 9757
rect 7557 9752 10567 9754
rect 7557 9696 7562 9752
rect 7618 9696 7930 9752
rect 7986 9696 10506 9752
rect 10562 9696 10567 9752
rect 7557 9694 10567 9696
rect 7557 9691 7623 9694
rect 7925 9691 7991 9694
rect 10501 9691 10567 9694
rect 10869 9754 10935 9757
rect 11094 9754 11100 9756
rect 10869 9752 11100 9754
rect 10869 9696 10874 9752
rect 10930 9696 11100 9752
rect 10869 9694 11100 9696
rect 10869 9691 10935 9694
rect 11094 9692 11100 9694
rect 11164 9692 11170 9756
rect 18321 9754 18387 9757
rect 11838 9752 18387 9754
rect 11838 9696 18326 9752
rect 18382 9696 18387 9752
rect 11838 9694 18387 9696
rect 19704 9754 19764 9966
rect 19885 10024 22892 10026
rect 19885 9968 19890 10024
rect 19946 9968 21914 10024
rect 21970 9968 22650 10024
rect 22706 9968 22892 10024
rect 19885 9966 22892 9968
rect 19885 9963 19951 9966
rect 21909 9963 21975 9966
rect 22645 9963 22711 9966
rect 19885 9890 19951 9893
rect 20437 9890 20503 9893
rect 19885 9888 20503 9890
rect 19885 9832 19890 9888
rect 19946 9832 20442 9888
rect 20498 9832 20503 9888
rect 19885 9830 20503 9832
rect 19885 9827 19951 9830
rect 20437 9827 20503 9830
rect 20621 9890 20687 9893
rect 22686 9890 22692 9892
rect 20621 9888 22692 9890
rect 20621 9832 20626 9888
rect 20682 9832 22692 9888
rect 20621 9830 22692 9832
rect 20621 9827 20687 9830
rect 22686 9828 22692 9830
rect 22756 9828 22762 9892
rect 22832 9890 22892 9966
rect 23105 10024 26667 10026
rect 23105 9968 23110 10024
rect 23166 9968 26606 10024
rect 26662 9968 26667 10024
rect 23105 9966 26667 9968
rect 23105 9963 23171 9966
rect 26601 9963 26667 9966
rect 26788 10024 27679 10026
rect 26788 9968 27618 10024
rect 27674 9968 27679 10024
rect 26788 9966 27679 9968
rect 24710 9890 24716 9892
rect 22832 9830 24716 9890
rect 24710 9828 24716 9830
rect 24780 9828 24786 9892
rect 26141 9890 26207 9893
rect 26788 9890 26848 9966
rect 27613 9963 27679 9966
rect 26141 9888 26848 9890
rect 26141 9832 26146 9888
rect 26202 9832 26848 9888
rect 26141 9830 26848 9832
rect 26141 9827 26207 9830
rect 26980 9824 27296 9825
rect 26980 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27296 9824
rect 26980 9759 27296 9760
rect 23473 9754 23539 9757
rect 26550 9754 26556 9756
rect 19704 9752 23539 9754
rect 19704 9696 23478 9752
rect 23534 9696 23539 9752
rect 19704 9694 23539 9696
rect 2681 9618 2747 9621
rect 2681 9616 2790 9618
rect 2681 9560 2686 9616
rect 2742 9560 2790 9616
rect 2681 9555 2790 9560
rect 2998 9556 3004 9620
rect 3068 9618 3074 9620
rect 3233 9618 3299 9621
rect 3068 9616 3299 9618
rect 3068 9560 3238 9616
rect 3294 9560 3299 9616
rect 3068 9558 3299 9560
rect 3068 9556 3074 9558
rect 3233 9555 3299 9558
rect 5441 9618 5507 9621
rect 6494 9618 6500 9620
rect 5441 9616 6500 9618
rect 5441 9560 5446 9616
rect 5502 9560 6500 9616
rect 5441 9558 6500 9560
rect 5441 9555 5507 9558
rect 6494 9556 6500 9558
rect 6564 9618 6570 9620
rect 9121 9618 9187 9621
rect 11838 9618 11898 9694
rect 18321 9691 18387 9694
rect 23473 9691 23539 9694
rect 24350 9694 26556 9754
rect 13486 9618 13492 9620
rect 6564 9616 11898 9618
rect 6564 9560 9126 9616
rect 9182 9560 11898 9616
rect 6564 9558 11898 9560
rect 13404 9558 13492 9618
rect 6564 9556 6570 9558
rect 9121 9555 9187 9558
rect 13486 9556 13492 9558
rect 13556 9618 13562 9620
rect 16573 9618 16639 9621
rect 13556 9616 16639 9618
rect 13556 9560 16578 9616
rect 16634 9560 16639 9616
rect 13556 9558 16639 9560
rect 13556 9556 13562 9558
rect 2730 9482 2790 9555
rect 11513 9482 11579 9485
rect 13118 9482 13124 9484
rect 2730 9422 9690 9482
rect 3049 9346 3115 9349
rect 3182 9346 3188 9348
rect 3049 9344 3188 9346
rect 3049 9288 3054 9344
rect 3110 9288 3188 9344
rect 3049 9286 3188 9288
rect 3049 9283 3115 9286
rect 3182 9284 3188 9286
rect 3252 9284 3258 9348
rect 4797 9346 4863 9349
rect 7741 9346 7807 9349
rect 4797 9344 7807 9346
rect 4797 9288 4802 9344
rect 4858 9288 7746 9344
rect 7802 9288 7807 9344
rect 4797 9286 7807 9288
rect 9630 9346 9690 9422
rect 11513 9480 13124 9482
rect 11513 9424 11518 9480
rect 11574 9424 13124 9480
rect 11513 9422 13124 9424
rect 11513 9419 11579 9422
rect 13118 9420 13124 9422
rect 13188 9420 13194 9484
rect 10225 9346 10291 9349
rect 10869 9346 10935 9349
rect 12617 9348 12683 9349
rect 9630 9344 10935 9346
rect 9630 9288 10230 9344
rect 10286 9288 10874 9344
rect 10930 9288 10935 9344
rect 9630 9286 10935 9288
rect 4797 9283 4863 9286
rect 7741 9283 7807 9286
rect 10225 9283 10291 9286
rect 10869 9283 10935 9286
rect 12566 9284 12572 9348
rect 12636 9346 12683 9348
rect 13169 9346 13235 9349
rect 13494 9346 13554 9556
rect 16573 9555 16639 9558
rect 18638 9556 18644 9620
rect 18708 9618 18714 9620
rect 20805 9618 20871 9621
rect 18708 9616 20871 9618
rect 18708 9560 20810 9616
rect 20866 9560 20871 9616
rect 18708 9558 20871 9560
rect 18708 9556 18714 9558
rect 20805 9555 20871 9558
rect 22277 9618 22343 9621
rect 22870 9618 22876 9620
rect 22277 9616 22876 9618
rect 22277 9560 22282 9616
rect 22338 9560 22876 9616
rect 22277 9558 22876 9560
rect 22277 9555 22343 9558
rect 22870 9556 22876 9558
rect 22940 9618 22946 9620
rect 24350 9618 24410 9694
rect 26550 9692 26556 9694
rect 26620 9754 26626 9756
rect 26693 9754 26759 9757
rect 26620 9752 26759 9754
rect 26620 9696 26698 9752
rect 26754 9696 26759 9752
rect 26620 9694 26759 9696
rect 26620 9692 26626 9694
rect 26693 9691 26759 9694
rect 22940 9558 24410 9618
rect 24485 9618 24551 9621
rect 25446 9618 25452 9620
rect 24485 9616 25452 9618
rect 24485 9560 24490 9616
rect 24546 9560 25452 9616
rect 24485 9558 25452 9560
rect 22940 9556 22946 9558
rect 24485 9555 24551 9558
rect 25446 9556 25452 9558
rect 25516 9556 25522 9620
rect 25681 9618 25747 9621
rect 27981 9618 28047 9621
rect 25681 9616 28047 9618
rect 25681 9560 25686 9616
rect 25742 9560 27986 9616
rect 28042 9560 28047 9616
rect 25681 9558 28047 9560
rect 25681 9555 25747 9558
rect 27981 9555 28047 9558
rect 28625 9618 28691 9621
rect 30741 9618 30807 9621
rect 28625 9616 30807 9618
rect 28625 9560 28630 9616
rect 28686 9560 30746 9616
rect 30802 9560 30807 9616
rect 28625 9558 30807 9560
rect 28625 9555 28691 9558
rect 30741 9555 30807 9558
rect 13629 9482 13695 9485
rect 16021 9482 16087 9485
rect 16389 9482 16455 9485
rect 13629 9480 15946 9482
rect 13629 9424 13634 9480
rect 13690 9424 15946 9480
rect 13629 9422 15946 9424
rect 13629 9419 13695 9422
rect 15886 9349 15946 9422
rect 16021 9480 16455 9482
rect 16021 9424 16026 9480
rect 16082 9424 16394 9480
rect 16450 9424 16455 9480
rect 16021 9422 16455 9424
rect 16021 9419 16087 9422
rect 16389 9419 16455 9422
rect 16798 9420 16804 9484
rect 16868 9482 16874 9484
rect 17769 9482 17835 9485
rect 16868 9480 17835 9482
rect 16868 9424 17774 9480
rect 17830 9424 17835 9480
rect 16868 9422 17835 9424
rect 16868 9420 16874 9422
rect 17769 9419 17835 9422
rect 18873 9482 18939 9485
rect 23933 9482 23999 9485
rect 18873 9480 23999 9482
rect 18873 9424 18878 9480
rect 18934 9424 23938 9480
rect 23994 9424 23999 9480
rect 18873 9422 23999 9424
rect 18873 9419 18939 9422
rect 23933 9419 23999 9422
rect 24209 9482 24275 9485
rect 29126 9482 29132 9484
rect 24209 9480 29132 9482
rect 24209 9424 24214 9480
rect 24270 9424 29132 9480
rect 24209 9422 29132 9424
rect 24209 9419 24275 9422
rect 29126 9420 29132 9422
rect 29196 9420 29202 9484
rect 12636 9344 12728 9346
rect 12678 9288 12728 9344
rect 12636 9286 12728 9288
rect 13169 9344 13554 9346
rect 13169 9288 13174 9344
rect 13230 9288 13554 9344
rect 13169 9286 13554 9288
rect 12636 9284 12683 9286
rect 12617 9283 12683 9284
rect 13169 9283 13235 9286
rect 13854 9284 13860 9348
rect 13924 9346 13930 9348
rect 15561 9346 15627 9349
rect 13924 9344 15627 9346
rect 13924 9288 15566 9344
rect 15622 9288 15627 9344
rect 13924 9286 15627 9288
rect 15886 9344 15995 9349
rect 15886 9288 15934 9344
rect 15990 9288 15995 9344
rect 15886 9286 15995 9288
rect 13924 9284 13930 9286
rect 15561 9283 15627 9286
rect 15929 9283 15995 9286
rect 16614 9284 16620 9348
rect 16684 9346 16690 9348
rect 17493 9346 17559 9349
rect 17902 9346 17908 9348
rect 16684 9344 17908 9346
rect 16684 9288 17498 9344
rect 17554 9288 17908 9344
rect 16684 9286 17908 9288
rect 16684 9284 16690 9286
rect 17493 9283 17559 9286
rect 17902 9284 17908 9286
rect 17972 9284 17978 9348
rect 18454 9284 18460 9348
rect 18524 9346 18530 9348
rect 18597 9346 18663 9349
rect 18524 9344 18663 9346
rect 18524 9288 18602 9344
rect 18658 9288 18663 9344
rect 18524 9286 18663 9288
rect 18524 9284 18530 9286
rect 18597 9283 18663 9286
rect 18965 9346 19031 9349
rect 19701 9346 19767 9349
rect 18965 9344 19767 9346
rect 18965 9288 18970 9344
rect 19026 9288 19706 9344
rect 19762 9288 19767 9344
rect 18965 9286 19767 9288
rect 18965 9283 19031 9286
rect 19701 9283 19767 9286
rect 20897 9346 20963 9349
rect 22645 9346 22711 9349
rect 20897 9344 22711 9346
rect 20897 9288 20902 9344
rect 20958 9288 22650 9344
rect 22706 9288 22711 9344
rect 20897 9286 22711 9288
rect 20897 9283 20963 9286
rect 22645 9283 22711 9286
rect 24025 9346 24091 9349
rect 26969 9346 27035 9349
rect 24025 9344 27035 9346
rect 24025 9288 24030 9344
rect 24086 9288 26974 9344
rect 27030 9288 27035 9344
rect 24025 9286 27035 9288
rect 24025 9283 24091 9286
rect 26969 9283 27035 9286
rect 29494 9284 29500 9348
rect 29564 9346 29570 9348
rect 29729 9346 29795 9349
rect 29564 9344 29795 9346
rect 29564 9288 29734 9344
rect 29790 9288 29795 9344
rect 29564 9286 29795 9288
rect 29564 9284 29570 9286
rect 29729 9283 29795 9286
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 12092 9280 12408 9281
rect 12092 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12408 9280
rect 12092 9215 12408 9216
rect 19866 9280 20182 9281
rect 19866 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20182 9280
rect 19866 9215 20182 9216
rect 27640 9280 27956 9281
rect 27640 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27956 9280
rect 27640 9215 27956 9216
rect 6637 9210 6703 9213
rect 11513 9210 11579 9213
rect 6637 9208 11579 9210
rect 6637 9152 6642 9208
rect 6698 9152 11518 9208
rect 11574 9152 11579 9208
rect 6637 9150 11579 9152
rect 6637 9147 6703 9150
rect 11513 9147 11579 9150
rect 13077 9210 13143 9213
rect 15377 9210 15443 9213
rect 13077 9208 15443 9210
rect 13077 9152 13082 9208
rect 13138 9152 15382 9208
rect 15438 9152 15443 9208
rect 13077 9150 15443 9152
rect 13077 9147 13143 9150
rect 15377 9147 15443 9150
rect 17401 9210 17467 9213
rect 18045 9210 18111 9213
rect 19701 9210 19767 9213
rect 17401 9208 19767 9210
rect 17401 9152 17406 9208
rect 17462 9152 18050 9208
rect 18106 9152 19706 9208
rect 19762 9152 19767 9208
rect 17401 9150 19767 9152
rect 17401 9147 17467 9150
rect 18045 9147 18111 9150
rect 19701 9147 19767 9150
rect 20805 9210 20871 9213
rect 23289 9210 23355 9213
rect 20805 9208 23355 9210
rect 20805 9152 20810 9208
rect 20866 9152 23294 9208
rect 23350 9152 23355 9208
rect 20805 9150 23355 9152
rect 20805 9147 20871 9150
rect 23289 9147 23355 9150
rect 24209 9210 24275 9213
rect 25773 9210 25839 9213
rect 24209 9208 25839 9210
rect 24209 9152 24214 9208
rect 24270 9152 25778 9208
rect 25834 9152 25839 9208
rect 24209 9150 25839 9152
rect 24209 9147 24275 9150
rect 25773 9147 25839 9150
rect 26182 9148 26188 9212
rect 26252 9210 26258 9212
rect 26509 9210 26575 9213
rect 28441 9212 28507 9213
rect 26252 9208 26575 9210
rect 26252 9152 26514 9208
rect 26570 9152 26575 9208
rect 26252 9150 26575 9152
rect 26252 9148 26258 9150
rect 26509 9147 26575 9150
rect 28390 9148 28396 9212
rect 28460 9210 28507 9212
rect 28460 9208 28552 9210
rect 28502 9152 28552 9208
rect 28460 9150 28552 9152
rect 28460 9148 28507 9150
rect 28441 9147 28507 9148
rect 3509 9074 3575 9077
rect 7741 9074 7807 9077
rect 3509 9072 7807 9074
rect 3509 9016 3514 9072
rect 3570 9016 7746 9072
rect 7802 9016 7807 9072
rect 3509 9014 7807 9016
rect 3509 9011 3575 9014
rect 7741 9011 7807 9014
rect 9254 9012 9260 9076
rect 9324 9074 9330 9076
rect 10041 9074 10107 9077
rect 9324 9072 10107 9074
rect 9324 9016 10046 9072
rect 10102 9016 10107 9072
rect 9324 9014 10107 9016
rect 9324 9012 9330 9014
rect 10041 9011 10107 9014
rect 10317 9074 10383 9077
rect 11278 9074 11284 9076
rect 10317 9072 11284 9074
rect 10317 9016 10322 9072
rect 10378 9016 11284 9072
rect 10317 9014 11284 9016
rect 10317 9011 10383 9014
rect 11278 9012 11284 9014
rect 11348 9012 11354 9076
rect 11605 9074 11671 9077
rect 11830 9074 11836 9076
rect 11605 9072 11836 9074
rect 11605 9016 11610 9072
rect 11666 9016 11836 9072
rect 11605 9014 11836 9016
rect 11605 9011 11671 9014
rect 11830 9012 11836 9014
rect 11900 9074 11906 9076
rect 13302 9074 13308 9076
rect 11900 9014 13308 9074
rect 11900 9012 11906 9014
rect 13302 9012 13308 9014
rect 13372 9012 13378 9076
rect 13721 9074 13787 9077
rect 13854 9074 13860 9076
rect 13721 9072 13860 9074
rect 13721 9016 13726 9072
rect 13782 9016 13860 9072
rect 13721 9014 13860 9016
rect 13721 9011 13787 9014
rect 13854 9012 13860 9014
rect 13924 9012 13930 9076
rect 13997 9074 14063 9077
rect 16246 9074 16252 9076
rect 13997 9072 16252 9074
rect 13997 9016 14002 9072
rect 14058 9016 16252 9072
rect 13997 9014 16252 9016
rect 13997 9011 14063 9014
rect 16246 9012 16252 9014
rect 16316 9074 16322 9076
rect 20805 9074 20871 9077
rect 22921 9074 22987 9077
rect 23054 9074 23060 9076
rect 16316 9072 20871 9074
rect 16316 9016 20810 9072
rect 20866 9016 20871 9072
rect 16316 9014 20871 9016
rect 16316 9012 16322 9014
rect 20805 9011 20871 9014
rect 21636 9072 23060 9074
rect 21636 9016 22926 9072
rect 22982 9016 23060 9072
rect 21636 9014 23060 9016
rect 4102 8876 4108 8940
rect 4172 8938 4178 8940
rect 4521 8938 4587 8941
rect 4838 8938 4844 8940
rect 4172 8936 4844 8938
rect 4172 8880 4526 8936
rect 4582 8880 4844 8936
rect 4172 8878 4844 8880
rect 4172 8876 4178 8878
rect 4521 8875 4587 8878
rect 4838 8876 4844 8878
rect 4908 8876 4914 8940
rect 5073 8938 5139 8941
rect 5206 8938 5212 8940
rect 5073 8936 5212 8938
rect 5073 8880 5078 8936
rect 5134 8880 5212 8936
rect 5073 8878 5212 8880
rect 5073 8875 5139 8878
rect 5206 8876 5212 8878
rect 5276 8876 5282 8940
rect 5993 8938 6059 8941
rect 6269 8938 6335 8941
rect 5993 8936 6335 8938
rect 5993 8880 5998 8936
rect 6054 8880 6274 8936
rect 6330 8880 6335 8936
rect 5993 8878 6335 8880
rect 5993 8875 6059 8878
rect 6269 8875 6335 8878
rect 7465 8938 7531 8941
rect 13905 8938 13971 8941
rect 7465 8936 13971 8938
rect 7465 8880 7470 8936
rect 7526 8880 13910 8936
rect 13966 8880 13971 8936
rect 7465 8878 13971 8880
rect 7465 8875 7531 8878
rect 13905 8875 13971 8878
rect 14038 8876 14044 8940
rect 14108 8938 14114 8940
rect 14181 8938 14247 8941
rect 21636 8938 21696 9014
rect 22921 9011 22987 9014
rect 23054 9012 23060 9014
rect 23124 9012 23130 9076
rect 25446 9012 25452 9076
rect 25516 9074 25522 9076
rect 25681 9074 25747 9077
rect 25516 9072 25747 9074
rect 25516 9016 25686 9072
rect 25742 9016 25747 9072
rect 25516 9014 25747 9016
rect 25516 9012 25522 9014
rect 25681 9011 25747 9014
rect 26509 9074 26575 9077
rect 26734 9074 26740 9076
rect 26509 9072 26740 9074
rect 26509 9016 26514 9072
rect 26570 9016 26740 9072
rect 26509 9014 26740 9016
rect 26509 9011 26575 9014
rect 26734 9012 26740 9014
rect 26804 9012 26810 9076
rect 14108 8936 21696 8938
rect 14108 8880 14186 8936
rect 14242 8880 21696 8936
rect 14108 8878 21696 8880
rect 21817 8938 21883 8941
rect 27521 8938 27587 8941
rect 21817 8936 27587 8938
rect 21817 8880 21822 8936
rect 21878 8880 27526 8936
rect 27582 8880 27587 8936
rect 21817 8878 27587 8880
rect 14108 8876 14114 8878
rect 14181 8875 14247 8878
rect 21817 8875 21883 8878
rect 27521 8875 27587 8878
rect 30230 8876 30236 8940
rect 30300 8938 30306 8940
rect 30373 8938 30439 8941
rect 30300 8936 30439 8938
rect 30300 8880 30378 8936
rect 30434 8880 30439 8936
rect 30300 8878 30439 8880
rect 30300 8876 30306 8878
rect 30373 8875 30439 8878
rect 4061 8802 4127 8805
rect 4521 8802 4587 8805
rect 7598 8802 7604 8804
rect 4061 8800 7604 8802
rect 4061 8744 4066 8800
rect 4122 8744 4526 8800
rect 4582 8744 7604 8800
rect 4061 8742 7604 8744
rect 4061 8739 4127 8742
rect 4521 8739 4587 8742
rect 7598 8740 7604 8742
rect 7668 8740 7674 8804
rect 8886 8740 8892 8804
rect 8956 8802 8962 8804
rect 9765 8802 9831 8805
rect 8956 8800 9831 8802
rect 8956 8744 9770 8800
rect 9826 8744 9831 8800
rect 8956 8742 9831 8744
rect 8956 8740 8962 8742
rect 9765 8739 9831 8742
rect 10133 8802 10199 8805
rect 10961 8802 11027 8805
rect 10133 8800 11027 8802
rect 10133 8744 10138 8800
rect 10194 8744 10966 8800
rect 11022 8744 11027 8800
rect 10133 8742 11027 8744
rect 10133 8739 10199 8742
rect 10961 8739 11027 8742
rect 11973 8802 12039 8805
rect 18505 8802 18571 8805
rect 18689 8804 18755 8805
rect 11973 8800 18571 8802
rect 11973 8744 11978 8800
rect 12034 8744 18510 8800
rect 18566 8744 18571 8800
rect 11973 8742 18571 8744
rect 11973 8739 12039 8742
rect 18505 8739 18571 8742
rect 18638 8740 18644 8804
rect 18708 8802 18755 8804
rect 19701 8802 19767 8805
rect 20621 8802 20687 8805
rect 18708 8800 18800 8802
rect 18750 8744 18800 8800
rect 18708 8742 18800 8744
rect 19701 8800 20687 8802
rect 19701 8744 19706 8800
rect 19762 8744 20626 8800
rect 20682 8744 20687 8800
rect 19701 8742 20687 8744
rect 18708 8740 18755 8742
rect 18689 8739 18755 8740
rect 19701 8739 19767 8742
rect 20621 8739 20687 8742
rect 21030 8740 21036 8804
rect 21100 8802 21106 8804
rect 22134 8802 22140 8804
rect 21100 8742 22140 8802
rect 21100 8740 21106 8742
rect 22134 8740 22140 8742
rect 22204 8802 22210 8804
rect 23749 8802 23815 8805
rect 22204 8800 23815 8802
rect 22204 8744 23754 8800
rect 23810 8744 23815 8800
rect 22204 8742 23815 8744
rect 22204 8740 22210 8742
rect 23749 8739 23815 8742
rect 24485 8802 24551 8805
rect 24485 8800 26618 8802
rect 24485 8744 24490 8800
rect 24546 8744 26618 8800
rect 24485 8742 26618 8744
rect 24485 8739 24551 8742
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 11432 8736 11748 8737
rect 11432 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11748 8736
rect 11432 8671 11748 8672
rect 19206 8736 19522 8737
rect 19206 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19522 8736
rect 19206 8671 19522 8672
rect 4337 8666 4403 8669
rect 7833 8666 7899 8669
rect 4337 8664 7899 8666
rect 4337 8608 4342 8664
rect 4398 8608 7838 8664
rect 7894 8608 7899 8664
rect 4337 8606 7899 8608
rect 4337 8603 4403 8606
rect 7833 8603 7899 8606
rect 8158 8606 10058 8666
rect 4613 8530 4679 8533
rect 5390 8530 5396 8532
rect 4613 8528 5396 8530
rect 4613 8472 4618 8528
rect 4674 8472 5396 8528
rect 4613 8470 5396 8472
rect 4613 8467 4679 8470
rect 5390 8468 5396 8470
rect 5460 8468 5466 8532
rect 7833 8530 7899 8533
rect 8158 8530 8218 8606
rect 7833 8528 8218 8530
rect 7833 8472 7838 8528
rect 7894 8472 8218 8528
rect 7833 8470 8218 8472
rect 8385 8530 8451 8533
rect 8518 8530 8524 8532
rect 8385 8528 8524 8530
rect 8385 8472 8390 8528
rect 8446 8472 8524 8528
rect 8385 8470 8524 8472
rect 7833 8467 7899 8470
rect 8385 8467 8451 8470
rect 8518 8468 8524 8470
rect 8588 8468 8594 8532
rect 8753 8530 8819 8533
rect 9121 8530 9187 8533
rect 8753 8528 9187 8530
rect 8753 8472 8758 8528
rect 8814 8472 9126 8528
rect 9182 8472 9187 8528
rect 8753 8470 9187 8472
rect 9998 8530 10058 8606
rect 12068 8606 13600 8666
rect 12068 8530 12128 8606
rect 9998 8470 12128 8530
rect 12341 8530 12407 8533
rect 13353 8530 13419 8533
rect 12341 8528 13419 8530
rect 12341 8472 12346 8528
rect 12402 8472 13358 8528
rect 13414 8472 13419 8528
rect 12341 8470 13419 8472
rect 13540 8530 13600 8606
rect 13670 8604 13676 8668
rect 13740 8666 13746 8668
rect 15009 8666 15075 8669
rect 15377 8668 15443 8669
rect 15326 8666 15332 8668
rect 13740 8664 15075 8666
rect 13740 8608 15014 8664
rect 15070 8608 15075 8664
rect 13740 8606 15075 8608
rect 15286 8606 15332 8666
rect 15396 8664 15443 8668
rect 15438 8608 15443 8664
rect 13740 8604 13746 8606
rect 15009 8603 15075 8606
rect 15326 8604 15332 8606
rect 15396 8604 15443 8608
rect 15377 8603 15443 8604
rect 15561 8666 15627 8669
rect 24393 8666 24459 8669
rect 15561 8664 19120 8666
rect 15561 8608 15566 8664
rect 15622 8608 19120 8664
rect 15561 8606 19120 8608
rect 15561 8603 15627 8606
rect 16665 8530 16731 8533
rect 13540 8528 16731 8530
rect 13540 8472 16670 8528
rect 16726 8472 16731 8528
rect 13540 8470 16731 8472
rect 8753 8467 8819 8470
rect 9121 8467 9187 8470
rect 12341 8467 12407 8470
rect 13353 8467 13419 8470
rect 16665 8467 16731 8470
rect 17534 8468 17540 8532
rect 17604 8530 17610 8532
rect 18689 8530 18755 8533
rect 17604 8528 18755 8530
rect 17604 8472 18694 8528
rect 18750 8472 18755 8528
rect 17604 8470 18755 8472
rect 19060 8530 19120 8606
rect 19612 8664 24459 8666
rect 19612 8608 24398 8664
rect 24454 8608 24459 8664
rect 19612 8606 24459 8608
rect 19612 8530 19672 8606
rect 24393 8603 24459 8606
rect 25814 8604 25820 8668
rect 25884 8666 25890 8668
rect 26417 8666 26483 8669
rect 25884 8664 26483 8666
rect 25884 8608 26422 8664
rect 26478 8608 26483 8664
rect 25884 8606 26483 8608
rect 25884 8604 25890 8606
rect 26417 8603 26483 8606
rect 21265 8530 21331 8533
rect 19060 8470 19672 8530
rect 19750 8528 21331 8530
rect 19750 8472 21270 8528
rect 21326 8472 21331 8528
rect 19750 8470 21331 8472
rect 17604 8468 17610 8470
rect 18689 8467 18755 8470
rect 1025 8396 1091 8397
rect 974 8394 980 8396
rect 934 8334 980 8394
rect 1044 8392 1091 8396
rect 1086 8336 1091 8392
rect 974 8332 980 8334
rect 1044 8332 1091 8336
rect 1025 8331 1091 8332
rect 3601 8394 3667 8397
rect 5206 8394 5212 8396
rect 3601 8392 5212 8394
rect 3601 8336 3606 8392
rect 3662 8336 5212 8392
rect 3601 8334 5212 8336
rect 3601 8331 3667 8334
rect 5206 8332 5212 8334
rect 5276 8394 5282 8396
rect 6913 8394 6979 8397
rect 10961 8394 11027 8397
rect 14181 8394 14247 8397
rect 15009 8394 15075 8397
rect 5276 8334 6792 8394
rect 5276 8332 5282 8334
rect 5073 8258 5139 8261
rect 5901 8258 5967 8261
rect 5073 8256 5967 8258
rect 5073 8200 5078 8256
rect 5134 8200 5906 8256
rect 5962 8200 5967 8256
rect 5073 8198 5967 8200
rect 6732 8258 6792 8334
rect 6913 8392 11027 8394
rect 6913 8336 6918 8392
rect 6974 8336 10966 8392
rect 11022 8336 11027 8392
rect 6913 8334 11027 8336
rect 6913 8331 6979 8334
rect 10961 8331 11027 8334
rect 11286 8334 12588 8394
rect 8293 8260 8359 8261
rect 8293 8258 8340 8260
rect 6732 8198 7114 8258
rect 8248 8256 8340 8258
rect 8248 8200 8298 8256
rect 8248 8198 8340 8200
rect 5073 8195 5139 8198
rect 5901 8195 5967 8198
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 749 7986 815 7989
rect 6913 7986 6979 7989
rect 749 7984 6979 7986
rect 749 7928 754 7984
rect 810 7928 6918 7984
rect 6974 7928 6979 7984
rect 749 7926 6979 7928
rect 7054 7986 7114 8198
rect 8293 8196 8340 8198
rect 8404 8196 8410 8260
rect 9397 8258 9463 8261
rect 11286 8258 11346 8334
rect 9397 8256 11346 8258
rect 9397 8200 9402 8256
rect 9458 8200 11346 8256
rect 9397 8198 11346 8200
rect 12528 8258 12588 8334
rect 14181 8392 15075 8394
rect 14181 8336 14186 8392
rect 14242 8336 15014 8392
rect 15070 8336 15075 8392
rect 14181 8334 15075 8336
rect 14181 8331 14247 8334
rect 15009 8331 15075 8334
rect 16481 8394 16547 8397
rect 18505 8394 18571 8397
rect 16481 8392 18571 8394
rect 16481 8336 16486 8392
rect 16542 8336 18510 8392
rect 18566 8336 18571 8392
rect 16481 8334 18571 8336
rect 18692 8394 18752 8467
rect 19750 8394 19810 8470
rect 21265 8467 21331 8470
rect 21633 8530 21699 8533
rect 23749 8530 23815 8533
rect 26049 8530 26115 8533
rect 21633 8528 26115 8530
rect 21633 8472 21638 8528
rect 21694 8472 23754 8528
rect 23810 8472 26054 8528
rect 26110 8472 26115 8528
rect 21633 8470 26115 8472
rect 26558 8530 26618 8742
rect 26980 8736 27296 8737
rect 26980 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27296 8736
rect 26980 8671 27296 8672
rect 26969 8530 27035 8533
rect 26558 8528 27035 8530
rect 26558 8472 26974 8528
rect 27030 8472 27035 8528
rect 26558 8470 27035 8472
rect 21633 8467 21699 8470
rect 23749 8467 23815 8470
rect 26049 8467 26115 8470
rect 26969 8467 27035 8470
rect 27889 8530 27955 8533
rect 27889 8528 29976 8530
rect 27889 8472 27894 8528
rect 27950 8472 29976 8528
rect 27889 8470 29976 8472
rect 27889 8467 27955 8470
rect 29916 8397 29976 8470
rect 18692 8334 19810 8394
rect 20069 8394 20135 8397
rect 22093 8394 22159 8397
rect 20069 8392 22159 8394
rect 20069 8336 20074 8392
rect 20130 8336 22098 8392
rect 22154 8336 22159 8392
rect 20069 8334 22159 8336
rect 16481 8331 16547 8334
rect 18505 8331 18571 8334
rect 20069 8331 20135 8334
rect 22093 8331 22159 8334
rect 23606 8332 23612 8396
rect 23676 8394 23682 8396
rect 23841 8394 23907 8397
rect 26693 8394 26759 8397
rect 23676 8392 26759 8394
rect 23676 8336 23846 8392
rect 23902 8336 26698 8392
rect 26754 8336 26759 8392
rect 23676 8334 26759 8336
rect 23676 8332 23682 8334
rect 23841 8331 23907 8334
rect 26693 8331 26759 8334
rect 27470 8332 27476 8396
rect 27540 8394 27546 8396
rect 27797 8394 27863 8397
rect 27540 8392 27863 8394
rect 27540 8336 27802 8392
rect 27858 8336 27863 8392
rect 27540 8334 27863 8336
rect 27540 8332 27546 8334
rect 27797 8331 27863 8334
rect 29126 8332 29132 8396
rect 29196 8394 29202 8396
rect 29453 8394 29519 8397
rect 29196 8392 29519 8394
rect 29196 8336 29458 8392
rect 29514 8336 29519 8392
rect 29196 8334 29519 8336
rect 29196 8332 29202 8334
rect 29453 8331 29519 8334
rect 29913 8392 29979 8397
rect 29913 8336 29918 8392
rect 29974 8336 29979 8392
rect 29913 8331 29979 8336
rect 15009 8260 15075 8261
rect 14590 8258 14596 8260
rect 12528 8198 14596 8258
rect 8293 8195 8402 8196
rect 9397 8195 9463 8198
rect 14590 8196 14596 8198
rect 14660 8196 14666 8260
rect 14958 8196 14964 8260
rect 15028 8258 15075 8260
rect 15561 8258 15627 8261
rect 19701 8258 19767 8261
rect 15028 8256 15120 8258
rect 15070 8200 15120 8256
rect 15028 8198 15120 8200
rect 15561 8256 19767 8258
rect 15561 8200 15566 8256
rect 15622 8200 19706 8256
rect 19762 8200 19767 8256
rect 15561 8198 19767 8200
rect 15028 8196 15075 8198
rect 15009 8195 15075 8196
rect 15561 8195 15627 8198
rect 19701 8195 19767 8198
rect 21950 8196 21956 8260
rect 22020 8258 22026 8260
rect 22093 8258 22159 8261
rect 22020 8256 22159 8258
rect 22020 8200 22098 8256
rect 22154 8200 22159 8256
rect 22020 8198 22159 8200
rect 22020 8196 22026 8198
rect 22093 8195 22159 8198
rect 22502 8196 22508 8260
rect 22572 8258 22578 8260
rect 22645 8258 22711 8261
rect 23289 8260 23355 8261
rect 22572 8256 22711 8258
rect 22572 8200 22650 8256
rect 22706 8200 22711 8256
rect 22572 8198 22711 8200
rect 22572 8196 22578 8198
rect 22645 8195 22711 8198
rect 23238 8196 23244 8260
rect 23308 8258 23355 8260
rect 24025 8258 24091 8261
rect 25957 8258 26023 8261
rect 23308 8256 23400 8258
rect 23350 8200 23400 8256
rect 23308 8198 23400 8200
rect 24025 8256 26023 8258
rect 24025 8200 24030 8256
rect 24086 8200 25962 8256
rect 26018 8200 26023 8256
rect 24025 8198 26023 8200
rect 23308 8196 23355 8198
rect 23289 8195 23355 8196
rect 24025 8195 24091 8198
rect 25957 8195 26023 8198
rect 26233 8258 26299 8261
rect 27061 8258 27127 8261
rect 26233 8256 27127 8258
rect 26233 8200 26238 8256
rect 26294 8200 27066 8256
rect 27122 8200 27127 8256
rect 26233 8198 27127 8200
rect 26233 8195 26299 8198
rect 27061 8195 27127 8198
rect 29269 8258 29335 8261
rect 31017 8258 31083 8261
rect 29269 8256 31083 8258
rect 29269 8200 29274 8256
rect 29330 8200 31022 8256
rect 31078 8200 31083 8256
rect 29269 8198 31083 8200
rect 29269 8195 29335 8198
rect 31017 8195 31083 8198
rect 8342 8122 8402 8195
rect 12092 8192 12408 8193
rect 12092 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12408 8192
rect 12092 8127 12408 8128
rect 19866 8192 20182 8193
rect 19866 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20182 8192
rect 19866 8127 20182 8128
rect 27640 8192 27956 8193
rect 27640 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27956 8192
rect 27640 8127 27956 8128
rect 9581 8122 9647 8125
rect 8342 8120 9647 8122
rect 8342 8064 9586 8120
rect 9642 8064 9647 8120
rect 8342 8062 9647 8064
rect 9581 8059 9647 8062
rect 10685 8122 10751 8125
rect 11881 8122 11947 8125
rect 10685 8120 11947 8122
rect 10685 8064 10690 8120
rect 10746 8064 11886 8120
rect 11942 8064 11947 8120
rect 10685 8062 11947 8064
rect 10685 8059 10751 8062
rect 11881 8059 11947 8062
rect 13445 8122 13511 8125
rect 14457 8122 14523 8125
rect 16389 8122 16455 8125
rect 13445 8120 14523 8122
rect 13445 8064 13450 8120
rect 13506 8064 14462 8120
rect 14518 8064 14523 8120
rect 13445 8062 14523 8064
rect 13445 8059 13511 8062
rect 14457 8059 14523 8062
rect 14598 8120 16455 8122
rect 14598 8064 16394 8120
rect 16450 8064 16455 8120
rect 14598 8062 16455 8064
rect 14598 7986 14658 8062
rect 16389 8059 16455 8062
rect 16665 8122 16731 8125
rect 17217 8122 17283 8125
rect 16665 8120 17283 8122
rect 16665 8064 16670 8120
rect 16726 8064 17222 8120
rect 17278 8064 17283 8120
rect 16665 8062 17283 8064
rect 16665 8059 16731 8062
rect 17217 8059 17283 8062
rect 17350 8060 17356 8124
rect 17420 8122 17426 8124
rect 17861 8122 17927 8125
rect 17420 8120 17927 8122
rect 17420 8064 17866 8120
rect 17922 8064 17927 8120
rect 17420 8062 17927 8064
rect 17420 8060 17426 8062
rect 17861 8059 17927 8062
rect 18086 8060 18092 8124
rect 18156 8122 18162 8124
rect 18229 8122 18295 8125
rect 18156 8120 18295 8122
rect 18156 8064 18234 8120
rect 18290 8064 18295 8120
rect 18156 8062 18295 8064
rect 18156 8060 18162 8062
rect 18229 8059 18295 8062
rect 18454 8060 18460 8124
rect 18524 8122 18530 8124
rect 18781 8122 18847 8125
rect 18965 8124 19031 8125
rect 18965 8122 19012 8124
rect 18524 8120 18847 8122
rect 18524 8064 18786 8120
rect 18842 8064 18847 8120
rect 18524 8062 18847 8064
rect 18920 8120 19012 8122
rect 18920 8064 18970 8120
rect 18920 8062 19012 8064
rect 18524 8060 18530 8062
rect 18781 8059 18847 8062
rect 18965 8060 19012 8062
rect 19076 8060 19082 8124
rect 21725 8122 21791 8125
rect 22318 8122 22324 8124
rect 21725 8120 22324 8122
rect 21725 8064 21730 8120
rect 21786 8064 22324 8120
rect 21725 8062 22324 8064
rect 18965 8059 19031 8060
rect 21725 8059 21791 8062
rect 22318 8060 22324 8062
rect 22388 8060 22394 8124
rect 22921 8122 22987 8125
rect 24485 8122 24551 8125
rect 22921 8120 24551 8122
rect 22921 8064 22926 8120
rect 22982 8064 24490 8120
rect 24546 8064 24551 8120
rect 22921 8062 24551 8064
rect 22921 8059 22987 8062
rect 24485 8059 24551 8062
rect 25129 8122 25195 8125
rect 25814 8122 25820 8124
rect 25129 8120 25820 8122
rect 25129 8064 25134 8120
rect 25190 8064 25820 8120
rect 25129 8062 25820 8064
rect 25129 8059 25195 8062
rect 25814 8060 25820 8062
rect 25884 8060 25890 8124
rect 26550 8060 26556 8124
rect 26620 8122 26626 8124
rect 26693 8122 26759 8125
rect 26620 8120 26759 8122
rect 26620 8064 26698 8120
rect 26754 8064 26759 8120
rect 26620 8062 26759 8064
rect 26620 8060 26626 8062
rect 26693 8059 26759 8062
rect 7054 7926 14658 7986
rect 14733 7986 14799 7989
rect 18781 7986 18847 7989
rect 24117 7986 24183 7989
rect 24577 7986 24643 7989
rect 14733 7984 24643 7986
rect 14733 7928 14738 7984
rect 14794 7928 18786 7984
rect 18842 7928 24122 7984
rect 24178 7928 24582 7984
rect 24638 7928 24643 7984
rect 14733 7926 24643 7928
rect 749 7923 815 7926
rect 6913 7923 6979 7926
rect 14733 7923 14799 7926
rect 18781 7923 18847 7926
rect 24117 7923 24183 7926
rect 24577 7923 24643 7926
rect 24710 7924 24716 7988
rect 24780 7986 24786 7988
rect 28625 7986 28691 7989
rect 24780 7984 28691 7986
rect 24780 7928 28630 7984
rect 28686 7928 28691 7984
rect 24780 7926 28691 7928
rect 24780 7924 24786 7926
rect 28625 7923 28691 7926
rect 4889 7850 4955 7853
rect 5993 7850 6059 7853
rect 16430 7850 16436 7852
rect 4889 7848 16436 7850
rect 4889 7792 4894 7848
rect 4950 7792 5998 7848
rect 6054 7792 16436 7848
rect 4889 7790 16436 7792
rect 4889 7787 4955 7790
rect 5993 7787 6059 7790
rect 16430 7788 16436 7790
rect 16500 7788 16506 7852
rect 26233 7850 26299 7853
rect 16622 7848 26299 7850
rect 16622 7792 26238 7848
rect 26294 7792 26299 7848
rect 16622 7790 26299 7792
rect 5073 7714 5139 7717
rect 9029 7714 9095 7717
rect 5073 7712 9095 7714
rect 5073 7656 5078 7712
rect 5134 7656 9034 7712
rect 9090 7656 9095 7712
rect 5073 7654 9095 7656
rect 5073 7651 5139 7654
rect 9029 7651 9095 7654
rect 11973 7714 12039 7717
rect 13813 7714 13879 7717
rect 11973 7712 13879 7714
rect 11973 7656 11978 7712
rect 12034 7656 13818 7712
rect 13874 7656 13879 7712
rect 11973 7654 13879 7656
rect 11973 7651 12039 7654
rect 13813 7651 13879 7654
rect 14089 7714 14155 7717
rect 14917 7714 14983 7717
rect 14089 7712 14983 7714
rect 14089 7656 14094 7712
rect 14150 7656 14922 7712
rect 14978 7656 14983 7712
rect 14089 7654 14983 7656
rect 14089 7651 14155 7654
rect 14917 7651 14983 7654
rect 15101 7714 15167 7717
rect 15837 7714 15903 7717
rect 15101 7712 15903 7714
rect 15101 7656 15106 7712
rect 15162 7656 15842 7712
rect 15898 7656 15903 7712
rect 15101 7654 15903 7656
rect 15101 7651 15167 7654
rect 15837 7651 15903 7654
rect 16021 7714 16087 7717
rect 16622 7714 16682 7790
rect 26233 7787 26299 7790
rect 27470 7788 27476 7852
rect 27540 7850 27546 7852
rect 27981 7850 28047 7853
rect 27540 7848 28047 7850
rect 27540 7792 27986 7848
rect 28042 7792 28047 7848
rect 27540 7790 28047 7792
rect 27540 7788 27546 7790
rect 27981 7787 28047 7790
rect 16021 7712 16682 7714
rect 16021 7656 16026 7712
rect 16082 7656 16682 7712
rect 16021 7654 16682 7656
rect 19793 7714 19859 7717
rect 24894 7714 24900 7716
rect 19793 7712 24900 7714
rect 19793 7656 19798 7712
rect 19854 7656 24900 7712
rect 19793 7654 24900 7656
rect 16021 7651 16087 7654
rect 19793 7651 19859 7654
rect 24894 7652 24900 7654
rect 24964 7652 24970 7716
rect 25037 7714 25103 7717
rect 26509 7714 26575 7717
rect 25037 7712 26575 7714
rect 25037 7656 25042 7712
rect 25098 7656 26514 7712
rect 26570 7656 26575 7712
rect 25037 7654 26575 7656
rect 25037 7651 25103 7654
rect 26509 7651 26575 7654
rect 28165 7716 28231 7717
rect 28165 7712 28212 7716
rect 28276 7714 28282 7716
rect 28165 7656 28170 7712
rect 28165 7652 28212 7656
rect 28276 7654 28322 7714
rect 28276 7652 28282 7654
rect 28165 7651 28231 7652
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 11432 7648 11748 7649
rect 11432 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11748 7648
rect 11432 7583 11748 7584
rect 19206 7648 19522 7649
rect 19206 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19522 7648
rect 19206 7583 19522 7584
rect 26980 7648 27296 7649
rect 26980 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27296 7648
rect 26980 7583 27296 7584
rect 4889 7578 4955 7581
rect 5022 7578 5028 7580
rect 4889 7576 5028 7578
rect 4889 7520 4894 7576
rect 4950 7520 5028 7576
rect 4889 7518 5028 7520
rect 4889 7515 4955 7518
rect 5022 7516 5028 7518
rect 5092 7516 5098 7580
rect 8702 7516 8708 7580
rect 8772 7578 8778 7580
rect 8845 7578 8911 7581
rect 8772 7576 8911 7578
rect 8772 7520 8850 7576
rect 8906 7520 8911 7576
rect 8772 7518 8911 7520
rect 8772 7516 8778 7518
rect 8845 7515 8911 7518
rect 9438 7516 9444 7580
rect 9508 7578 9514 7580
rect 9949 7578 10015 7581
rect 20345 7580 20411 7581
rect 18270 7578 18276 7580
rect 9508 7576 10015 7578
rect 9508 7520 9954 7576
rect 10010 7520 10015 7576
rect 9508 7518 10015 7520
rect 9508 7516 9514 7518
rect 9949 7515 10015 7518
rect 12436 7518 18276 7578
rect 12436 7445 12496 7518
rect 18270 7516 18276 7518
rect 18340 7516 18346 7580
rect 20294 7516 20300 7580
rect 20364 7578 20411 7580
rect 21449 7578 21515 7581
rect 22553 7578 22619 7581
rect 20364 7576 20456 7578
rect 20406 7520 20456 7576
rect 20364 7518 20456 7520
rect 21449 7576 22619 7578
rect 21449 7520 21454 7576
rect 21510 7520 22558 7576
rect 22614 7520 22619 7576
rect 21449 7518 22619 7520
rect 20364 7516 20411 7518
rect 20345 7515 20411 7516
rect 21449 7515 21515 7518
rect 22553 7515 22619 7518
rect 23013 7578 23079 7581
rect 25497 7578 25563 7581
rect 23013 7576 25563 7578
rect 23013 7520 23018 7576
rect 23074 7520 25502 7576
rect 25558 7520 25563 7576
rect 23013 7518 25563 7520
rect 23013 7515 23079 7518
rect 25497 7515 25563 7518
rect 2221 7442 2287 7445
rect 6821 7442 6887 7445
rect 8753 7442 8819 7445
rect 2221 7440 6887 7442
rect 2221 7384 2226 7440
rect 2282 7384 6826 7440
rect 6882 7384 6887 7440
rect 2221 7382 6887 7384
rect 2221 7379 2287 7382
rect 6821 7379 6887 7382
rect 7054 7440 8819 7442
rect 7054 7384 8758 7440
rect 8814 7384 8819 7440
rect 7054 7382 8819 7384
rect 3969 7306 4035 7309
rect 7054 7306 7114 7382
rect 8753 7379 8819 7382
rect 9581 7442 9647 7445
rect 12433 7442 12499 7445
rect 9581 7440 12499 7442
rect 9581 7384 9586 7440
rect 9642 7384 12438 7440
rect 12494 7384 12499 7440
rect 9581 7382 12499 7384
rect 9581 7379 9647 7382
rect 12433 7379 12499 7382
rect 13537 7442 13603 7445
rect 24669 7442 24735 7445
rect 25313 7442 25379 7445
rect 30557 7442 30623 7445
rect 13537 7440 30623 7442
rect 13537 7384 13542 7440
rect 13598 7384 24674 7440
rect 24730 7384 25318 7440
rect 25374 7384 30562 7440
rect 30618 7384 30623 7440
rect 13537 7382 30623 7384
rect 13537 7379 13603 7382
rect 24669 7379 24735 7382
rect 25313 7379 25379 7382
rect 30557 7379 30623 7382
rect 3969 7304 7114 7306
rect 3969 7248 3974 7304
rect 4030 7248 7114 7304
rect 3969 7246 7114 7248
rect 7649 7306 7715 7309
rect 7649 7304 14658 7306
rect 7649 7248 7654 7304
rect 7710 7248 14658 7304
rect 7649 7246 14658 7248
rect 3969 7243 4035 7246
rect 7649 7243 7715 7246
rect 5349 7170 5415 7173
rect 6177 7170 6243 7173
rect 7925 7170 7991 7173
rect 5349 7168 7991 7170
rect 5349 7112 5354 7168
rect 5410 7112 6182 7168
rect 6238 7112 7930 7168
rect 7986 7112 7991 7168
rect 5349 7110 7991 7112
rect 5349 7107 5415 7110
rect 6177 7107 6243 7110
rect 7925 7107 7991 7110
rect 8661 7170 8727 7173
rect 9029 7170 9095 7173
rect 8661 7168 9095 7170
rect 8661 7112 8666 7168
rect 8722 7112 9034 7168
rect 9090 7112 9095 7168
rect 8661 7110 9095 7112
rect 8661 7107 8727 7110
rect 9029 7107 9095 7110
rect 12525 7170 12591 7173
rect 13905 7170 13971 7173
rect 12525 7168 13971 7170
rect 12525 7112 12530 7168
rect 12586 7112 13910 7168
rect 13966 7112 13971 7168
rect 12525 7110 13971 7112
rect 14598 7170 14658 7246
rect 14774 7244 14780 7308
rect 14844 7306 14850 7308
rect 18965 7306 19031 7309
rect 14844 7304 19031 7306
rect 14844 7248 18970 7304
rect 19026 7248 19031 7304
rect 14844 7246 19031 7248
rect 14844 7244 14850 7246
rect 18965 7243 19031 7246
rect 19566 7246 20500 7306
rect 16481 7170 16547 7173
rect 19566 7170 19626 7246
rect 14598 7110 16314 7170
rect 12525 7107 12591 7110
rect 13905 7107 13971 7110
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 12092 7104 12408 7105
rect 12092 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12408 7104
rect 12092 7039 12408 7040
rect 7097 7034 7163 7037
rect 9622 7034 9628 7036
rect 7097 7032 9628 7034
rect 7097 6976 7102 7032
rect 7158 6976 9628 7032
rect 7097 6974 9628 6976
rect 7097 6971 7163 6974
rect 9622 6972 9628 6974
rect 9692 6972 9698 7036
rect 12617 7034 12683 7037
rect 15469 7034 15535 7037
rect 12617 7032 15535 7034
rect 12617 6976 12622 7032
rect 12678 6976 15474 7032
rect 15530 6976 15535 7032
rect 12617 6974 15535 6976
rect 12617 6971 12683 6974
rect 15469 6971 15535 6974
rect 657 6898 723 6901
rect 13537 6898 13603 6901
rect 16113 6898 16179 6901
rect 657 6896 13603 6898
rect 657 6840 662 6896
rect 718 6840 13542 6896
rect 13598 6840 13603 6896
rect 657 6838 13603 6840
rect 657 6835 723 6838
rect 13537 6835 13603 6838
rect 13678 6896 16179 6898
rect 13678 6840 16118 6896
rect 16174 6840 16179 6896
rect 13678 6838 16179 6840
rect 16254 6898 16314 7110
rect 16481 7168 19626 7170
rect 16481 7112 16486 7168
rect 16542 7112 19626 7168
rect 16481 7110 19626 7112
rect 16481 7107 16547 7110
rect 19866 7104 20182 7105
rect 19866 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20182 7104
rect 19866 7039 20182 7040
rect 16941 7036 17007 7037
rect 16941 7032 16988 7036
rect 17052 7034 17058 7036
rect 16941 6976 16946 7032
rect 16941 6972 16988 6976
rect 17052 6974 17098 7034
rect 17861 7032 17927 7037
rect 17861 6976 17866 7032
rect 17922 6976 17927 7032
rect 17052 6972 17058 6974
rect 16941 6971 17007 6972
rect 17861 6971 17927 6976
rect 20440 7034 20500 7246
rect 20621 7304 20687 7309
rect 20621 7248 20626 7304
rect 20682 7248 20687 7304
rect 20621 7243 20687 7248
rect 20805 7306 20871 7309
rect 27429 7306 27495 7309
rect 20805 7304 27495 7306
rect 20805 7248 20810 7304
rect 20866 7248 27434 7304
rect 27490 7248 27495 7304
rect 20805 7246 27495 7248
rect 20805 7243 20871 7246
rect 27429 7243 27495 7246
rect 20624 7170 20684 7243
rect 24209 7170 24275 7173
rect 20624 7168 24275 7170
rect 20624 7112 24214 7168
rect 24270 7112 24275 7168
rect 20624 7110 24275 7112
rect 24209 7107 24275 7110
rect 24393 7170 24459 7173
rect 24853 7170 24919 7173
rect 25773 7170 25839 7173
rect 24393 7168 25839 7170
rect 24393 7112 24398 7168
rect 24454 7112 24858 7168
rect 24914 7112 25778 7168
rect 25834 7112 25839 7168
rect 24393 7110 25839 7112
rect 24393 7107 24459 7110
rect 24853 7107 24919 7110
rect 25773 7107 25839 7110
rect 27640 7104 27956 7105
rect 27640 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27956 7104
rect 27640 7039 27956 7040
rect 21725 7034 21791 7037
rect 20440 7032 21791 7034
rect 20440 6976 21730 7032
rect 21786 6976 21791 7032
rect 20440 6974 21791 6976
rect 21725 6971 21791 6974
rect 22553 7034 22619 7037
rect 24577 7034 24643 7037
rect 27470 7034 27476 7036
rect 22553 7032 27476 7034
rect 22553 6976 22558 7032
rect 22614 6976 24582 7032
rect 24638 6976 27476 7032
rect 22553 6974 27476 6976
rect 22553 6971 22619 6974
rect 24577 6971 24643 6974
rect 27470 6972 27476 6974
rect 27540 6972 27546 7036
rect 17864 6898 17924 6971
rect 19885 6898 19951 6901
rect 16254 6896 19951 6898
rect 16254 6840 19890 6896
rect 19946 6840 19951 6896
rect 16254 6838 19951 6840
rect 3969 6762 4035 6765
rect 8293 6762 8359 6765
rect 12433 6762 12499 6765
rect 3969 6760 4952 6762
rect 3969 6704 3974 6760
rect 4030 6704 4952 6760
rect 3969 6702 4952 6704
rect 3969 6699 4035 6702
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 4892 6490 4952 6702
rect 8293 6760 12499 6762
rect 8293 6704 8298 6760
rect 8354 6704 12438 6760
rect 12494 6704 12499 6760
rect 8293 6702 12499 6704
rect 8293 6699 8359 6702
rect 12433 6699 12499 6702
rect 12985 6762 13051 6765
rect 13678 6762 13738 6838
rect 16113 6835 16179 6838
rect 19885 6835 19951 6838
rect 20161 6898 20227 6901
rect 20478 6898 20484 6900
rect 20161 6896 20484 6898
rect 20161 6840 20166 6896
rect 20222 6840 20484 6896
rect 20161 6838 20484 6840
rect 20161 6835 20227 6838
rect 20478 6836 20484 6838
rect 20548 6836 20554 6900
rect 20897 6898 20963 6901
rect 22737 6898 22803 6901
rect 20897 6896 22803 6898
rect 20897 6840 20902 6896
rect 20958 6840 22742 6896
rect 22798 6840 22803 6896
rect 20897 6838 22803 6840
rect 20897 6835 20963 6838
rect 22737 6835 22803 6838
rect 24526 6836 24532 6900
rect 24596 6898 24602 6900
rect 24853 6898 24919 6901
rect 24596 6896 24919 6898
rect 24596 6840 24858 6896
rect 24914 6840 24919 6896
rect 24596 6838 24919 6840
rect 24596 6836 24602 6838
rect 24853 6835 24919 6838
rect 12985 6760 13738 6762
rect 12985 6704 12990 6760
rect 13046 6704 13738 6760
rect 12985 6702 13738 6704
rect 15101 6762 15167 6765
rect 23749 6762 23815 6765
rect 25681 6762 25747 6765
rect 28717 6762 28783 6765
rect 15101 6760 23815 6762
rect 15101 6704 15106 6760
rect 15162 6704 23754 6760
rect 23810 6704 23815 6760
rect 15101 6702 23815 6704
rect 12985 6699 13051 6702
rect 15101 6699 15167 6702
rect 23749 6699 23815 6702
rect 23982 6760 28783 6762
rect 23982 6704 25686 6760
rect 25742 6704 28722 6760
rect 28778 6704 28783 6760
rect 23982 6702 28783 6704
rect 10225 6626 10291 6629
rect 10726 6626 10732 6628
rect 10225 6624 10732 6626
rect 10225 6568 10230 6624
rect 10286 6568 10732 6624
rect 10225 6566 10732 6568
rect 10225 6563 10291 6566
rect 10726 6564 10732 6566
rect 10796 6564 10802 6628
rect 11973 6626 12039 6629
rect 12566 6626 12572 6628
rect 11973 6624 12572 6626
rect 11973 6568 11978 6624
rect 12034 6568 12572 6624
rect 11973 6566 12572 6568
rect 11973 6563 12039 6566
rect 12566 6564 12572 6566
rect 12636 6564 12642 6628
rect 19885 6626 19951 6629
rect 20897 6626 20963 6629
rect 19885 6624 20963 6626
rect 19885 6568 19890 6624
rect 19946 6568 20902 6624
rect 20958 6568 20963 6624
rect 19885 6566 20963 6568
rect 19885 6563 19951 6566
rect 20897 6563 20963 6566
rect 23657 6626 23723 6629
rect 23982 6626 24042 6702
rect 25681 6699 25747 6702
rect 28717 6699 28783 6702
rect 23657 6624 24042 6626
rect 23657 6568 23662 6624
rect 23718 6568 24042 6624
rect 23657 6566 24042 6568
rect 23657 6563 23723 6566
rect 11432 6560 11748 6561
rect 11432 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11748 6560
rect 11432 6495 11748 6496
rect 19206 6560 19522 6561
rect 19206 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19522 6560
rect 19206 6495 19522 6496
rect 26980 6560 27296 6561
rect 26980 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27296 6560
rect 26980 6495 27296 6496
rect 10685 6490 10751 6493
rect 4892 6488 10751 6490
rect 4892 6432 10690 6488
rect 10746 6432 10751 6488
rect 4892 6430 10751 6432
rect 10685 6427 10751 6430
rect 11881 6490 11947 6493
rect 12934 6490 12940 6492
rect 11881 6488 12940 6490
rect 11881 6432 11886 6488
rect 11942 6432 12940 6488
rect 11881 6430 12940 6432
rect 11881 6427 11947 6430
rect 12934 6428 12940 6430
rect 13004 6490 13010 6492
rect 18137 6490 18203 6493
rect 13004 6488 18203 6490
rect 13004 6432 18142 6488
rect 18198 6432 18203 6488
rect 13004 6430 18203 6432
rect 13004 6428 13010 6430
rect 18137 6427 18203 6430
rect 18638 6428 18644 6492
rect 18708 6490 18714 6492
rect 18873 6490 18939 6493
rect 18708 6488 18939 6490
rect 18708 6432 18878 6488
rect 18934 6432 18939 6488
rect 18708 6430 18939 6432
rect 18708 6428 18714 6430
rect 18873 6427 18939 6430
rect 22369 6490 22435 6493
rect 25589 6490 25655 6493
rect 22369 6488 25655 6490
rect 22369 6432 22374 6488
rect 22430 6432 25594 6488
rect 25650 6432 25655 6488
rect 22369 6430 25655 6432
rect 22369 6427 22435 6430
rect 25589 6427 25655 6430
rect 4797 6354 4863 6357
rect 5390 6354 5396 6356
rect 4797 6352 5396 6354
rect 4797 6296 4802 6352
rect 4858 6296 5396 6352
rect 4797 6294 5396 6296
rect 4797 6291 4863 6294
rect 5390 6292 5396 6294
rect 5460 6354 5466 6356
rect 5809 6354 5875 6357
rect 11053 6356 11119 6357
rect 11053 6354 11100 6356
rect 5460 6352 10426 6354
rect 5460 6296 5814 6352
rect 5870 6296 10426 6352
rect 5460 6294 10426 6296
rect 11008 6352 11100 6354
rect 11008 6296 11058 6352
rect 11008 6294 11100 6296
rect 5460 6292 5466 6294
rect 5809 6291 5875 6294
rect 841 6218 907 6221
rect 9397 6218 9463 6221
rect 10366 6220 10426 6294
rect 11053 6292 11100 6294
rect 11164 6292 11170 6356
rect 12249 6354 12315 6357
rect 16614 6354 16620 6356
rect 12249 6352 16620 6354
rect 12249 6296 12254 6352
rect 12310 6296 16620 6352
rect 12249 6294 16620 6296
rect 11053 6291 11119 6292
rect 12249 6291 12315 6294
rect 16614 6292 16620 6294
rect 16684 6292 16690 6356
rect 17677 6354 17743 6357
rect 21030 6354 21036 6356
rect 17677 6352 21036 6354
rect 17677 6296 17682 6352
rect 17738 6296 21036 6352
rect 17677 6294 21036 6296
rect 17677 6291 17743 6294
rect 21030 6292 21036 6294
rect 21100 6292 21106 6356
rect 21265 6354 21331 6357
rect 23657 6354 23723 6357
rect 21265 6352 23723 6354
rect 21265 6296 21270 6352
rect 21326 6296 23662 6352
rect 23718 6296 23723 6352
rect 21265 6294 23723 6296
rect 21265 6291 21331 6294
rect 23657 6291 23723 6294
rect 24025 6354 24091 6357
rect 30925 6354 30991 6357
rect 24025 6352 30991 6354
rect 24025 6296 24030 6352
rect 24086 6296 30930 6352
rect 30986 6296 30991 6352
rect 24025 6294 30991 6296
rect 24025 6291 24091 6294
rect 30925 6291 30991 6294
rect 841 6216 9463 6218
rect 841 6160 846 6216
rect 902 6160 9402 6216
rect 9458 6160 9463 6216
rect 841 6158 9463 6160
rect 841 6155 907 6158
rect 9397 6155 9463 6158
rect 10358 6156 10364 6220
rect 10428 6218 10434 6220
rect 17861 6218 17927 6221
rect 21817 6218 21883 6221
rect 29453 6218 29519 6221
rect 10428 6216 21883 6218
rect 10428 6160 17866 6216
rect 17922 6160 21822 6216
rect 21878 6160 21883 6216
rect 10428 6158 21883 6160
rect 10428 6156 10434 6158
rect 17861 6155 17927 6158
rect 21817 6155 21883 6158
rect 23430 6216 29519 6218
rect 23430 6160 29458 6216
rect 29514 6160 29519 6216
rect 23430 6158 29519 6160
rect 5257 6082 5323 6085
rect 8017 6084 8083 6085
rect 7966 6082 7972 6084
rect 5257 6080 7972 6082
rect 8036 6082 8083 6084
rect 9489 6082 9555 6085
rect 11789 6082 11855 6085
rect 8036 6080 8128 6082
rect 5257 6024 5262 6080
rect 5318 6024 7972 6080
rect 8078 6024 8128 6080
rect 5257 6022 7972 6024
rect 5257 6019 5323 6022
rect 7966 6020 7972 6022
rect 8036 6022 8128 6024
rect 9489 6080 11855 6082
rect 9489 6024 9494 6080
rect 9550 6024 11794 6080
rect 11850 6024 11855 6080
rect 9489 6022 11855 6024
rect 8036 6020 8083 6022
rect 8017 6019 8083 6020
rect 9489 6019 9555 6022
rect 11789 6019 11855 6022
rect 14733 6082 14799 6085
rect 18413 6082 18479 6085
rect 14733 6080 18479 6082
rect 14733 6024 14738 6080
rect 14794 6024 18418 6080
rect 18474 6024 18479 6080
rect 14733 6022 18479 6024
rect 14733 6019 14799 6022
rect 18413 6019 18479 6022
rect 18965 6082 19031 6085
rect 19425 6082 19491 6085
rect 18965 6080 19491 6082
rect 18965 6024 18970 6080
rect 19026 6024 19430 6080
rect 19486 6024 19491 6080
rect 18965 6022 19491 6024
rect 18965 6019 19031 6022
rect 19425 6019 19491 6022
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 12092 6016 12408 6017
rect 12092 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12408 6016
rect 12092 5951 12408 5952
rect 19866 6016 20182 6017
rect 19866 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20182 6016
rect 19866 5951 20182 5952
rect 6545 5946 6611 5949
rect 9857 5946 9923 5949
rect 6545 5944 9923 5946
rect 6545 5888 6550 5944
rect 6606 5888 9862 5944
rect 9918 5888 9923 5944
rect 6545 5886 9923 5888
rect 6545 5883 6611 5886
rect 9857 5883 9923 5886
rect 10542 5884 10548 5948
rect 10612 5946 10618 5948
rect 11329 5946 11395 5949
rect 10612 5944 11395 5946
rect 10612 5888 11334 5944
rect 11390 5888 11395 5944
rect 10612 5886 11395 5888
rect 10612 5884 10618 5886
rect 11329 5883 11395 5886
rect 14457 5946 14523 5949
rect 15510 5946 15516 5948
rect 14457 5944 15516 5946
rect 14457 5888 14462 5944
rect 14518 5888 15516 5944
rect 14457 5886 15516 5888
rect 14457 5883 14523 5886
rect 15510 5884 15516 5886
rect 15580 5946 15586 5948
rect 23430 5946 23490 6158
rect 29453 6155 29519 6158
rect 27640 6016 27956 6017
rect 27640 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27956 6016
rect 27640 5951 27956 5952
rect 15580 5886 16682 5946
rect 15580 5884 15586 5886
rect 8150 5748 8156 5812
rect 8220 5810 8226 5812
rect 10869 5810 10935 5813
rect 12985 5810 13051 5813
rect 16481 5810 16547 5813
rect 8220 5750 8402 5810
rect 8220 5748 8226 5750
rect 2497 5676 2563 5677
rect 2446 5612 2452 5676
rect 2516 5674 2563 5676
rect 7649 5674 7715 5677
rect 8150 5674 8156 5676
rect 2516 5672 2608 5674
rect 2558 5616 2608 5672
rect 2516 5614 2608 5616
rect 7649 5672 8156 5674
rect 7649 5616 7654 5672
rect 7710 5616 8156 5672
rect 7649 5614 8156 5616
rect 2516 5612 2563 5614
rect 2497 5611 2563 5612
rect 7649 5611 7715 5614
rect 8150 5612 8156 5614
rect 8220 5612 8226 5676
rect 8342 5674 8402 5750
rect 10869 5808 12220 5810
rect 10869 5752 10874 5808
rect 10930 5752 12220 5808
rect 10869 5750 12220 5752
rect 10869 5747 10935 5750
rect 10869 5674 10935 5677
rect 12160 5674 12220 5750
rect 12985 5808 16547 5810
rect 12985 5752 12990 5808
rect 13046 5752 16486 5808
rect 16542 5752 16547 5808
rect 12985 5750 16547 5752
rect 16622 5810 16682 5886
rect 20256 5886 23490 5946
rect 23657 5946 23723 5949
rect 23657 5944 27538 5946
rect 23657 5888 23662 5944
rect 23718 5888 27538 5944
rect 23657 5886 27538 5888
rect 20256 5810 20316 5886
rect 23657 5883 23723 5886
rect 16622 5750 20316 5810
rect 20897 5810 20963 5813
rect 24025 5810 24091 5813
rect 20897 5808 24091 5810
rect 20897 5752 20902 5808
rect 20958 5752 24030 5808
rect 24086 5752 24091 5808
rect 20897 5750 24091 5752
rect 27478 5810 27538 5886
rect 29637 5810 29703 5813
rect 27478 5808 29703 5810
rect 27478 5752 29642 5808
rect 29698 5752 29703 5808
rect 27478 5750 29703 5752
rect 12985 5747 13051 5750
rect 16481 5747 16547 5750
rect 20897 5747 20963 5750
rect 24025 5747 24091 5750
rect 29637 5747 29703 5750
rect 19333 5674 19399 5677
rect 25078 5674 25084 5676
rect 8342 5672 10935 5674
rect 8342 5616 10874 5672
rect 10930 5616 10935 5672
rect 8342 5614 10935 5616
rect 10869 5611 10935 5614
rect 11286 5614 12082 5674
rect 12160 5614 18752 5674
rect 4102 5476 4108 5540
rect 4172 5538 4178 5540
rect 4245 5538 4311 5541
rect 4172 5536 4311 5538
rect 4172 5480 4250 5536
rect 4306 5480 4311 5536
rect 4172 5478 4311 5480
rect 4172 5476 4178 5478
rect 4245 5475 4311 5478
rect 7465 5538 7531 5541
rect 7782 5538 7788 5540
rect 7465 5536 7788 5538
rect 7465 5480 7470 5536
rect 7526 5480 7788 5536
rect 7465 5478 7788 5480
rect 7465 5475 7531 5478
rect 7782 5476 7788 5478
rect 7852 5538 7858 5540
rect 11286 5538 11346 5614
rect 7852 5478 11346 5538
rect 7852 5476 7858 5478
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 11432 5472 11748 5473
rect 11432 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11748 5472
rect 11432 5407 11748 5408
rect 12022 5402 12082 5614
rect 18692 5541 18752 5614
rect 19333 5672 25084 5674
rect 19333 5616 19338 5672
rect 19394 5616 25084 5672
rect 19333 5614 25084 5616
rect 19333 5611 19399 5614
rect 25078 5612 25084 5614
rect 25148 5674 25154 5676
rect 26877 5674 26943 5677
rect 25148 5672 26943 5674
rect 25148 5616 26882 5672
rect 26938 5616 26943 5672
rect 25148 5614 26943 5616
rect 25148 5612 25154 5614
rect 26877 5611 26943 5614
rect 12709 5538 12775 5541
rect 15142 5538 15148 5540
rect 12709 5536 15148 5538
rect 12709 5480 12714 5536
rect 12770 5480 15148 5536
rect 12709 5478 15148 5480
rect 12709 5475 12775 5478
rect 15142 5476 15148 5478
rect 15212 5476 15218 5540
rect 18689 5538 18755 5541
rect 18822 5538 18828 5540
rect 18689 5536 18828 5538
rect 18689 5480 18694 5536
rect 18750 5480 18828 5536
rect 18689 5478 18828 5480
rect 18689 5475 18755 5478
rect 18822 5476 18828 5478
rect 18892 5476 18898 5540
rect 19206 5472 19522 5473
rect 19206 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19522 5472
rect 19206 5407 19522 5408
rect 26980 5472 27296 5473
rect 26980 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27296 5472
rect 26980 5407 27296 5408
rect 14917 5402 14983 5405
rect 12022 5400 14983 5402
rect 12022 5344 14922 5400
rect 14978 5344 14983 5400
rect 12022 5342 14983 5344
rect 14917 5339 14983 5342
rect 15101 5402 15167 5405
rect 18873 5402 18939 5405
rect 15101 5400 18939 5402
rect 15101 5344 15106 5400
rect 15162 5344 18878 5400
rect 18934 5344 18939 5400
rect 15101 5342 18939 5344
rect 15101 5339 15167 5342
rect 18873 5339 18939 5342
rect 20294 5340 20300 5404
rect 20364 5402 20370 5404
rect 20897 5402 20963 5405
rect 20364 5400 20963 5402
rect 20364 5344 20902 5400
rect 20958 5344 20963 5400
rect 20364 5342 20963 5344
rect 20364 5340 20370 5342
rect 20897 5339 20963 5342
rect 1853 5266 1919 5269
rect 16021 5266 16087 5269
rect 25405 5266 25471 5269
rect 1853 5264 25471 5266
rect 1853 5208 1858 5264
rect 1914 5208 16026 5264
rect 16082 5208 25410 5264
rect 25466 5208 25471 5264
rect 1853 5206 25471 5208
rect 1853 5203 1919 5206
rect 16021 5203 16087 5206
rect 25405 5203 25471 5206
rect 2497 5130 2563 5133
rect 12709 5130 12775 5133
rect 2497 5128 12775 5130
rect 2497 5072 2502 5128
rect 2558 5072 12714 5128
rect 12770 5072 12775 5128
rect 2497 5070 12775 5072
rect 2497 5067 2563 5070
rect 12709 5067 12775 5070
rect 14917 5130 14983 5133
rect 20989 5130 21055 5133
rect 28533 5132 28599 5133
rect 28533 5130 28580 5132
rect 14917 5128 21055 5130
rect 14917 5072 14922 5128
rect 14978 5072 20994 5128
rect 21050 5072 21055 5128
rect 14917 5070 21055 5072
rect 28488 5128 28580 5130
rect 28488 5072 28538 5128
rect 28488 5070 28580 5072
rect 14917 5067 14983 5070
rect 20989 5067 21055 5070
rect 28533 5068 28580 5070
rect 28644 5068 28650 5132
rect 28533 5067 28599 5068
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 12092 4928 12408 4929
rect 12092 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12408 4928
rect 12092 4863 12408 4864
rect 19866 4928 20182 4929
rect 19866 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20182 4928
rect 19866 4863 20182 4864
rect 27640 4928 27956 4929
rect 27640 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27956 4928
rect 27640 4863 27956 4864
rect 10041 4858 10107 4861
rect 15745 4860 15811 4861
rect 10174 4858 10180 4860
rect 10041 4856 10180 4858
rect 10041 4800 10046 4856
rect 10102 4800 10180 4856
rect 10041 4798 10180 4800
rect 10041 4795 10107 4798
rect 10174 4796 10180 4798
rect 10244 4796 10250 4860
rect 15694 4796 15700 4860
rect 15764 4858 15811 4860
rect 19057 4858 19123 4861
rect 20805 4860 20871 4861
rect 20805 4858 20852 4860
rect 15764 4856 19123 4858
rect 15806 4800 19062 4856
rect 19118 4800 19123 4856
rect 15764 4798 19123 4800
rect 20760 4856 20852 4858
rect 20760 4800 20810 4856
rect 20760 4798 20852 4800
rect 15764 4796 15811 4798
rect 15745 4795 15811 4796
rect 19057 4795 19123 4798
rect 20805 4796 20852 4798
rect 20916 4796 20922 4860
rect 20805 4795 20871 4796
rect 3182 4660 3188 4724
rect 3252 4722 3258 4724
rect 11973 4722 12039 4725
rect 3252 4720 12039 4722
rect 3252 4664 11978 4720
rect 12034 4664 12039 4720
rect 3252 4662 12039 4664
rect 3252 4660 3258 4662
rect 11973 4659 12039 4662
rect 15142 4660 15148 4724
rect 15212 4722 15218 4724
rect 21449 4722 21515 4725
rect 15212 4720 21515 4722
rect 15212 4664 21454 4720
rect 21510 4664 21515 4720
rect 15212 4662 21515 4664
rect 15212 4660 15218 4662
rect 21449 4659 21515 4662
rect 9673 4586 9739 4589
rect 10409 4586 10475 4589
rect 9673 4584 10475 4586
rect 9673 4528 9678 4584
rect 9734 4528 10414 4584
rect 10470 4528 10475 4584
rect 9673 4526 10475 4528
rect 9673 4523 9739 4526
rect 10409 4523 10475 4526
rect 10910 4524 10916 4588
rect 10980 4586 10986 4588
rect 12617 4586 12683 4589
rect 10980 4584 12683 4586
rect 10980 4528 12622 4584
rect 12678 4528 12683 4584
rect 10980 4526 12683 4528
rect 10980 4524 10986 4526
rect 12617 4523 12683 4526
rect 11973 4450 12039 4453
rect 17401 4450 17467 4453
rect 11973 4448 17467 4450
rect 11973 4392 11978 4448
rect 12034 4392 17406 4448
rect 17462 4392 17467 4448
rect 11973 4390 17467 4392
rect 11973 4387 12039 4390
rect 17401 4387 17467 4390
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 11432 4384 11748 4385
rect 11432 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11748 4384
rect 11432 4319 11748 4320
rect 19206 4384 19522 4385
rect 19206 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19522 4384
rect 19206 4319 19522 4320
rect 26980 4384 27296 4385
rect 26980 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27296 4384
rect 26980 4319 27296 4320
rect 3182 4116 3188 4180
rect 3252 4178 3258 4180
rect 3601 4178 3667 4181
rect 3252 4176 3667 4178
rect 3252 4120 3606 4176
rect 3662 4120 3667 4176
rect 3252 4118 3667 4120
rect 3252 4116 3258 4118
rect 3601 4115 3667 4118
rect 9397 4178 9463 4181
rect 9949 4178 10015 4181
rect 18321 4178 18387 4181
rect 21817 4180 21883 4181
rect 9397 4176 18387 4178
rect 9397 4120 9402 4176
rect 9458 4120 9954 4176
rect 10010 4120 18326 4176
rect 18382 4120 18387 4176
rect 9397 4118 18387 4120
rect 9397 4115 9463 4118
rect 9949 4115 10015 4118
rect 18321 4115 18387 4118
rect 21766 4116 21772 4180
rect 21836 4178 21883 4180
rect 21836 4176 21928 4178
rect 21878 4120 21928 4176
rect 21836 4118 21928 4120
rect 21836 4116 21883 4118
rect 21817 4115 21883 4116
rect 2630 3980 2636 4044
rect 2700 4042 2706 4044
rect 11605 4042 11671 4045
rect 26182 4042 26188 4044
rect 2700 4040 11671 4042
rect 2700 3984 11610 4040
rect 11666 3984 11671 4040
rect 2700 3982 11671 3984
rect 2700 3980 2706 3982
rect 11605 3979 11671 3982
rect 11884 3982 26188 4042
rect 11278 3844 11284 3908
rect 11348 3906 11354 3908
rect 11884 3906 11944 3982
rect 26182 3980 26188 3982
rect 26252 3980 26258 4044
rect 11348 3846 11944 3906
rect 13445 3906 13511 3909
rect 16062 3906 16068 3908
rect 13445 3904 16068 3906
rect 13445 3848 13450 3904
rect 13506 3848 16068 3904
rect 13445 3846 16068 3848
rect 11348 3844 11354 3846
rect 13445 3843 13511 3846
rect 16062 3844 16068 3846
rect 16132 3906 16138 3908
rect 16481 3906 16547 3909
rect 16132 3904 16547 3906
rect 16132 3848 16486 3904
rect 16542 3848 16547 3904
rect 16132 3846 16547 3848
rect 16132 3844 16138 3846
rect 16481 3843 16547 3846
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 12092 3840 12408 3841
rect 12092 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12408 3840
rect 12092 3775 12408 3776
rect 19866 3840 20182 3841
rect 19866 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20182 3840
rect 19866 3775 20182 3776
rect 27640 3840 27956 3841
rect 27640 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27956 3840
rect 27640 3775 27956 3776
rect 12750 3708 12756 3772
rect 12820 3770 12826 3772
rect 12893 3770 12959 3773
rect 14273 3770 14339 3773
rect 12820 3768 14339 3770
rect 12820 3712 12898 3768
rect 12954 3712 14278 3768
rect 14334 3712 14339 3768
rect 12820 3710 14339 3712
rect 12820 3708 12826 3710
rect 12893 3707 12959 3710
rect 14273 3707 14339 3710
rect 2446 3572 2452 3636
rect 2516 3634 2522 3636
rect 10593 3634 10659 3637
rect 13813 3634 13879 3637
rect 2516 3574 2790 3634
rect 2516 3572 2522 3574
rect 2730 2954 2790 3574
rect 10593 3632 13879 3634
rect 10593 3576 10598 3632
rect 10654 3576 13818 3632
rect 13874 3576 13879 3632
rect 10593 3574 13879 3576
rect 10593 3571 10659 3574
rect 13813 3571 13879 3574
rect 13997 3634 14063 3637
rect 14365 3636 14431 3637
rect 14365 3634 14412 3636
rect 13997 3632 14412 3634
rect 13997 3576 14002 3632
rect 14058 3576 14370 3632
rect 13997 3574 14412 3576
rect 13997 3571 14063 3574
rect 14365 3572 14412 3574
rect 14476 3572 14482 3636
rect 14365 3571 14431 3572
rect 8150 3436 8156 3500
rect 8220 3498 8226 3500
rect 23841 3498 23907 3501
rect 8220 3496 23907 3498
rect 8220 3440 23846 3496
rect 23902 3440 23907 3496
rect 8220 3438 23907 3440
rect 8220 3436 8226 3438
rect 23841 3435 23907 3438
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 11432 3296 11748 3297
rect 11432 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11748 3296
rect 11432 3231 11748 3232
rect 19206 3296 19522 3297
rect 19206 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19522 3296
rect 19206 3231 19522 3232
rect 26980 3296 27296 3297
rect 26980 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27296 3296
rect 26980 3231 27296 3232
rect 7966 3028 7972 3092
rect 8036 3090 8042 3092
rect 28993 3090 29059 3093
rect 8036 3088 29059 3090
rect 8036 3032 28998 3088
rect 29054 3032 29059 3088
rect 8036 3030 29059 3032
rect 8036 3028 8042 3030
rect 28993 3027 29059 3030
rect 13854 2954 13860 2956
rect 2730 2894 13860 2954
rect 13854 2892 13860 2894
rect 13924 2954 13930 2956
rect 21265 2954 21331 2957
rect 13924 2952 21331 2954
rect 13924 2896 21270 2952
rect 21326 2896 21331 2952
rect 13924 2894 21331 2896
rect 13924 2892 13930 2894
rect 21265 2891 21331 2894
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 12092 2752 12408 2753
rect 12092 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12408 2752
rect 12092 2687 12408 2688
rect 19866 2752 20182 2753
rect 19866 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20182 2752
rect 19866 2687 20182 2688
rect 27640 2752 27956 2753
rect 27640 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27956 2752
rect 27640 2687 27956 2688
rect 19701 2682 19767 2685
rect 12574 2680 19767 2682
rect 12574 2624 19706 2680
rect 19762 2624 19767 2680
rect 12574 2622 19767 2624
rect 8845 2546 8911 2549
rect 12574 2546 12634 2622
rect 19701 2619 19767 2622
rect 24853 2682 24919 2685
rect 25630 2682 25636 2684
rect 24853 2680 25636 2682
rect 24853 2624 24858 2680
rect 24914 2624 25636 2680
rect 24853 2622 25636 2624
rect 24853 2619 24919 2622
rect 25630 2620 25636 2622
rect 25700 2620 25706 2684
rect 21214 2546 21220 2548
rect 8845 2544 12634 2546
rect 8845 2488 8850 2544
rect 8906 2488 12634 2544
rect 8845 2486 12634 2488
rect 12758 2486 21220 2546
rect 8845 2483 8911 2486
rect 10869 2410 10935 2413
rect 12758 2410 12818 2486
rect 21214 2484 21220 2486
rect 21284 2484 21290 2548
rect 10869 2408 12818 2410
rect 10869 2352 10874 2408
rect 10930 2352 12818 2408
rect 10869 2350 12818 2352
rect 10869 2347 10935 2350
rect 13118 2348 13124 2412
rect 13188 2410 13194 2412
rect 20662 2410 20668 2412
rect 13188 2350 20668 2410
rect 13188 2348 13194 2350
rect 20662 2348 20668 2350
rect 20732 2348 20738 2412
rect 19701 2274 19767 2277
rect 23606 2274 23612 2276
rect 19701 2272 23612 2274
rect 19701 2216 19706 2272
rect 19762 2216 23612 2272
rect 19701 2214 23612 2216
rect 19701 2211 19767 2214
rect 23606 2212 23612 2214
rect 23676 2212 23682 2276
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 11432 2208 11748 2209
rect 11432 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11748 2208
rect 11432 2143 11748 2144
rect 19206 2208 19522 2209
rect 19206 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19522 2208
rect 19206 2143 19522 2144
rect 26980 2208 27296 2209
rect 26980 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27296 2208
rect 26980 2143 27296 2144
rect 13302 1940 13308 2004
rect 13372 2002 13378 2004
rect 26417 2002 26483 2005
rect 13372 2000 26483 2002
rect 13372 1944 26422 2000
rect 26478 1944 26483 2000
rect 13372 1942 26483 1944
rect 13372 1940 13378 1942
rect 26417 1939 26483 1942
rect 1158 1804 1164 1868
rect 1228 1866 1234 1868
rect 21582 1866 21588 1868
rect 1228 1806 21588 1866
rect 1228 1804 1234 1806
rect 21582 1804 21588 1806
rect 21652 1804 21658 1868
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 12092 1664 12408 1665
rect 12092 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12408 1664
rect 12092 1599 12408 1600
rect 19866 1664 20182 1665
rect 19866 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20182 1664
rect 19866 1599 20182 1600
rect 27640 1664 27956 1665
rect 27640 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27956 1664
rect 27640 1599 27956 1600
rect 1117 1458 1183 1461
rect 15878 1458 15884 1460
rect 1117 1456 15884 1458
rect 1117 1400 1122 1456
rect 1178 1400 15884 1456
rect 1117 1398 15884 1400
rect 1117 1395 1183 1398
rect 15878 1396 15884 1398
rect 15948 1396 15954 1460
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 11432 1120 11748 1121
rect 11432 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11748 1120
rect 11432 1055 11748 1056
rect 19206 1120 19522 1121
rect 19206 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19522 1120
rect 19206 1055 19522 1056
rect 26980 1120 27296 1121
rect 26980 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27296 1120
rect 26980 1055 27296 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 12092 576 12408 577
rect 12092 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12408 576
rect 12092 511 12408 512
rect 19866 576 20182 577
rect 19866 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20182 576
rect 19866 511 20182 512
rect 27640 576 27956 577
rect 27640 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27956 576
rect 27640 511 27956 512
<< via3 >>
rect 20300 22068 20364 22132
rect 11652 21932 11716 21996
rect 12204 21992 12268 21996
rect 12204 21936 12254 21992
rect 12254 21936 12268 21992
rect 12204 21932 12268 21936
rect 8892 21796 8956 21860
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 11438 21788 11502 21792
rect 11438 21732 11442 21788
rect 11442 21732 11498 21788
rect 11498 21732 11502 21788
rect 11438 21728 11502 21732
rect 11518 21788 11582 21792
rect 11518 21732 11522 21788
rect 11522 21732 11578 21788
rect 11578 21732 11582 21788
rect 11518 21728 11582 21732
rect 11598 21788 11662 21792
rect 11598 21732 11602 21788
rect 11602 21732 11658 21788
rect 11658 21732 11662 21788
rect 11598 21728 11662 21732
rect 11678 21788 11742 21792
rect 11678 21732 11682 21788
rect 11682 21732 11738 21788
rect 11738 21732 11742 21788
rect 11678 21728 11742 21732
rect 6132 21720 6196 21724
rect 6132 21664 6182 21720
rect 6182 21664 6196 21720
rect 6132 21660 6196 21664
rect 6684 21720 6748 21724
rect 6684 21664 6734 21720
rect 6734 21664 6748 21720
rect 6684 21660 6748 21664
rect 7236 21720 7300 21724
rect 7236 21664 7286 21720
rect 7286 21664 7300 21720
rect 7236 21660 7300 21664
rect 7788 21720 7852 21724
rect 7788 21664 7838 21720
rect 7838 21664 7852 21720
rect 7788 21660 7852 21664
rect 8340 21720 8404 21724
rect 8340 21664 8390 21720
rect 8390 21664 8404 21720
rect 8340 21660 8404 21664
rect 9444 21720 9508 21724
rect 9444 21664 9494 21720
rect 9494 21664 9508 21720
rect 9444 21660 9508 21664
rect 9996 21720 10060 21724
rect 9996 21664 10046 21720
rect 10046 21664 10060 21720
rect 9996 21660 10060 21664
rect 10548 21720 10612 21724
rect 10548 21664 10598 21720
rect 10598 21664 10612 21720
rect 10548 21660 10612 21664
rect 11100 21720 11164 21724
rect 11100 21664 11150 21720
rect 11150 21664 11164 21720
rect 11100 21660 11164 21664
rect 12756 21720 12820 21724
rect 12756 21664 12806 21720
rect 12806 21664 12820 21720
rect 12756 21660 12820 21664
rect 13308 21720 13372 21724
rect 13308 21664 13358 21720
rect 13358 21664 13372 21720
rect 13308 21660 13372 21664
rect 13860 21720 13924 21724
rect 13860 21664 13910 21720
rect 13910 21664 13924 21720
rect 13860 21660 13924 21664
rect 16620 21720 16684 21724
rect 16620 21664 16670 21720
rect 16670 21664 16684 21720
rect 16620 21660 16684 21664
rect 8156 21524 8220 21588
rect 24348 21932 24412 21996
rect 19212 21788 19276 21792
rect 19212 21732 19216 21788
rect 19216 21732 19272 21788
rect 19272 21732 19276 21788
rect 19212 21728 19276 21732
rect 19292 21788 19356 21792
rect 19292 21732 19296 21788
rect 19296 21732 19352 21788
rect 19352 21732 19356 21788
rect 19292 21728 19356 21732
rect 19372 21788 19436 21792
rect 19372 21732 19376 21788
rect 19376 21732 19432 21788
rect 19432 21732 19436 21788
rect 19372 21728 19436 21732
rect 19452 21788 19516 21792
rect 19452 21732 19456 21788
rect 19456 21732 19512 21788
rect 19512 21732 19516 21788
rect 19452 21728 19516 21732
rect 26986 21788 27050 21792
rect 26986 21732 26990 21788
rect 26990 21732 27046 21788
rect 27046 21732 27050 21788
rect 26986 21728 27050 21732
rect 27066 21788 27130 21792
rect 27066 21732 27070 21788
rect 27070 21732 27126 21788
rect 27126 21732 27130 21788
rect 27066 21728 27130 21732
rect 27146 21788 27210 21792
rect 27146 21732 27150 21788
rect 27150 21732 27206 21788
rect 27206 21732 27210 21788
rect 27146 21728 27210 21732
rect 27226 21788 27290 21792
rect 27226 21732 27230 21788
rect 27230 21732 27286 21788
rect 27286 21732 27290 21788
rect 27226 21728 27290 21732
rect 18828 21524 18892 21588
rect 25820 21524 25884 21588
rect 18276 21388 18340 21452
rect 26556 21388 26620 21452
rect 21036 21252 21100 21316
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 12098 21244 12162 21248
rect 12098 21188 12102 21244
rect 12102 21188 12158 21244
rect 12158 21188 12162 21244
rect 12098 21184 12162 21188
rect 12178 21244 12242 21248
rect 12178 21188 12182 21244
rect 12182 21188 12238 21244
rect 12238 21188 12242 21244
rect 12178 21184 12242 21188
rect 12258 21244 12322 21248
rect 12258 21188 12262 21244
rect 12262 21188 12318 21244
rect 12318 21188 12322 21244
rect 12258 21184 12322 21188
rect 12338 21244 12402 21248
rect 12338 21188 12342 21244
rect 12342 21188 12398 21244
rect 12398 21188 12402 21244
rect 12338 21184 12402 21188
rect 19872 21244 19936 21248
rect 19872 21188 19876 21244
rect 19876 21188 19932 21244
rect 19932 21188 19936 21244
rect 19872 21184 19936 21188
rect 19952 21244 20016 21248
rect 19952 21188 19956 21244
rect 19956 21188 20012 21244
rect 20012 21188 20016 21244
rect 19952 21184 20016 21188
rect 20032 21244 20096 21248
rect 20032 21188 20036 21244
rect 20036 21188 20092 21244
rect 20092 21188 20096 21244
rect 20032 21184 20096 21188
rect 20112 21244 20176 21248
rect 20112 21188 20116 21244
rect 20116 21188 20172 21244
rect 20172 21188 20176 21244
rect 20112 21184 20176 21188
rect 27646 21244 27710 21248
rect 27646 21188 27650 21244
rect 27650 21188 27706 21244
rect 27706 21188 27710 21244
rect 27646 21184 27710 21188
rect 27726 21244 27790 21248
rect 27726 21188 27730 21244
rect 27730 21188 27786 21244
rect 27786 21188 27790 21244
rect 27726 21184 27790 21188
rect 27806 21244 27870 21248
rect 27806 21188 27810 21244
rect 27810 21188 27866 21244
rect 27866 21188 27870 21244
rect 27806 21184 27870 21188
rect 27886 21244 27950 21248
rect 27886 21188 27890 21244
rect 27890 21188 27946 21244
rect 27946 21188 27950 21244
rect 27886 21184 27950 21188
rect 17172 21116 17236 21180
rect 15516 21040 15580 21044
rect 15516 20984 15530 21040
rect 15530 20984 15580 21040
rect 15516 20980 15580 20984
rect 27476 20980 27540 21044
rect 24164 20844 24228 20908
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 11438 20700 11502 20704
rect 11438 20644 11442 20700
rect 11442 20644 11498 20700
rect 11498 20644 11502 20700
rect 11438 20640 11502 20644
rect 11518 20700 11582 20704
rect 11518 20644 11522 20700
rect 11522 20644 11578 20700
rect 11578 20644 11582 20700
rect 11518 20640 11582 20644
rect 11598 20700 11662 20704
rect 11598 20644 11602 20700
rect 11602 20644 11658 20700
rect 11658 20644 11662 20700
rect 11598 20640 11662 20644
rect 11678 20700 11742 20704
rect 11678 20644 11682 20700
rect 11682 20644 11738 20700
rect 11738 20644 11742 20700
rect 11678 20640 11742 20644
rect 19212 20700 19276 20704
rect 19212 20644 19216 20700
rect 19216 20644 19272 20700
rect 19272 20644 19276 20700
rect 19212 20640 19276 20644
rect 19292 20700 19356 20704
rect 19292 20644 19296 20700
rect 19296 20644 19352 20700
rect 19352 20644 19356 20700
rect 19292 20640 19356 20644
rect 19372 20700 19436 20704
rect 19372 20644 19376 20700
rect 19376 20644 19432 20700
rect 19432 20644 19436 20700
rect 19372 20640 19436 20644
rect 19452 20700 19516 20704
rect 19452 20644 19456 20700
rect 19456 20644 19512 20700
rect 19512 20644 19516 20700
rect 19452 20640 19516 20644
rect 26986 20700 27050 20704
rect 26986 20644 26990 20700
rect 26990 20644 27046 20700
rect 27046 20644 27050 20700
rect 26986 20640 27050 20644
rect 27066 20700 27130 20704
rect 27066 20644 27070 20700
rect 27070 20644 27126 20700
rect 27126 20644 27130 20700
rect 27066 20640 27130 20644
rect 27146 20700 27210 20704
rect 27146 20644 27150 20700
rect 27150 20644 27206 20700
rect 27206 20644 27210 20700
rect 27146 20640 27210 20644
rect 27226 20700 27290 20704
rect 27226 20644 27230 20700
rect 27230 20644 27286 20700
rect 27286 20644 27290 20700
rect 27226 20640 27290 20644
rect 14412 20632 14476 20636
rect 14412 20576 14462 20632
rect 14462 20576 14476 20632
rect 14412 20572 14476 20576
rect 16068 20572 16132 20636
rect 17724 20572 17788 20636
rect 980 20436 1044 20500
rect 26188 20436 26252 20500
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 12098 20156 12162 20160
rect 12098 20100 12102 20156
rect 12102 20100 12158 20156
rect 12158 20100 12162 20156
rect 12098 20096 12162 20100
rect 12178 20156 12242 20160
rect 12178 20100 12182 20156
rect 12182 20100 12238 20156
rect 12238 20100 12242 20156
rect 12178 20096 12242 20100
rect 12258 20156 12322 20160
rect 12258 20100 12262 20156
rect 12262 20100 12318 20156
rect 12318 20100 12322 20156
rect 12258 20096 12322 20100
rect 12338 20156 12402 20160
rect 12338 20100 12342 20156
rect 12342 20100 12398 20156
rect 12398 20100 12402 20156
rect 12338 20096 12402 20100
rect 19872 20156 19936 20160
rect 19872 20100 19876 20156
rect 19876 20100 19932 20156
rect 19932 20100 19936 20156
rect 19872 20096 19936 20100
rect 19952 20156 20016 20160
rect 19952 20100 19956 20156
rect 19956 20100 20012 20156
rect 20012 20100 20016 20156
rect 19952 20096 20016 20100
rect 20032 20156 20096 20160
rect 20032 20100 20036 20156
rect 20036 20100 20092 20156
rect 20092 20100 20096 20156
rect 20032 20096 20096 20100
rect 20112 20156 20176 20160
rect 20112 20100 20116 20156
rect 20116 20100 20172 20156
rect 20172 20100 20176 20156
rect 20112 20096 20176 20100
rect 27646 20156 27710 20160
rect 27646 20100 27650 20156
rect 27650 20100 27706 20156
rect 27706 20100 27710 20156
rect 27646 20096 27710 20100
rect 27726 20156 27790 20160
rect 27726 20100 27730 20156
rect 27730 20100 27786 20156
rect 27786 20100 27790 20156
rect 27726 20096 27790 20100
rect 27806 20156 27870 20160
rect 27806 20100 27810 20156
rect 27810 20100 27866 20156
rect 27866 20100 27870 20156
rect 27806 20096 27870 20100
rect 27886 20156 27950 20160
rect 27886 20100 27890 20156
rect 27890 20100 27946 20156
rect 27946 20100 27950 20156
rect 27886 20096 27950 20100
rect 21036 20028 21100 20092
rect 14964 19952 15028 19956
rect 14964 19896 15014 19952
rect 15014 19896 15028 19952
rect 14964 19892 15028 19896
rect 24716 19756 24780 19820
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 11438 19612 11502 19616
rect 11438 19556 11442 19612
rect 11442 19556 11498 19612
rect 11498 19556 11502 19612
rect 11438 19552 11502 19556
rect 11518 19612 11582 19616
rect 11518 19556 11522 19612
rect 11522 19556 11578 19612
rect 11578 19556 11582 19612
rect 11518 19552 11582 19556
rect 11598 19612 11662 19616
rect 11598 19556 11602 19612
rect 11602 19556 11658 19612
rect 11658 19556 11662 19612
rect 11598 19552 11662 19556
rect 11678 19612 11742 19616
rect 11678 19556 11682 19612
rect 11682 19556 11738 19612
rect 11738 19556 11742 19612
rect 11678 19552 11742 19556
rect 16436 19348 16500 19412
rect 19212 19612 19276 19616
rect 19212 19556 19216 19612
rect 19216 19556 19272 19612
rect 19272 19556 19276 19612
rect 19212 19552 19276 19556
rect 19292 19612 19356 19616
rect 19292 19556 19296 19612
rect 19296 19556 19352 19612
rect 19352 19556 19356 19612
rect 19292 19552 19356 19556
rect 19372 19612 19436 19616
rect 19372 19556 19376 19612
rect 19376 19556 19432 19612
rect 19432 19556 19436 19612
rect 19372 19552 19436 19556
rect 19452 19612 19516 19616
rect 19452 19556 19456 19612
rect 19456 19556 19512 19612
rect 19512 19556 19516 19612
rect 19452 19552 19516 19556
rect 26986 19612 27050 19616
rect 26986 19556 26990 19612
rect 26990 19556 27046 19612
rect 27046 19556 27050 19612
rect 26986 19552 27050 19556
rect 27066 19612 27130 19616
rect 27066 19556 27070 19612
rect 27070 19556 27126 19612
rect 27126 19556 27130 19612
rect 27066 19552 27130 19556
rect 27146 19612 27210 19616
rect 27146 19556 27150 19612
rect 27150 19556 27206 19612
rect 27206 19556 27210 19612
rect 27146 19552 27210 19556
rect 27226 19612 27290 19616
rect 27226 19556 27230 19612
rect 27230 19556 27286 19612
rect 27286 19556 27290 19612
rect 27226 19552 27290 19556
rect 22508 19484 22572 19548
rect 26004 19484 26068 19548
rect 14044 19212 14108 19276
rect 20668 19212 20732 19276
rect 28764 19212 28828 19276
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 12098 19068 12162 19072
rect 12098 19012 12102 19068
rect 12102 19012 12158 19068
rect 12158 19012 12162 19068
rect 12098 19008 12162 19012
rect 12178 19068 12242 19072
rect 12178 19012 12182 19068
rect 12182 19012 12238 19068
rect 12238 19012 12242 19068
rect 12178 19008 12242 19012
rect 12258 19068 12322 19072
rect 12258 19012 12262 19068
rect 12262 19012 12318 19068
rect 12318 19012 12322 19068
rect 12258 19008 12322 19012
rect 12338 19068 12402 19072
rect 12338 19012 12342 19068
rect 12342 19012 12398 19068
rect 12398 19012 12402 19068
rect 12338 19008 12402 19012
rect 19872 19068 19936 19072
rect 19872 19012 19876 19068
rect 19876 19012 19932 19068
rect 19932 19012 19936 19068
rect 19872 19008 19936 19012
rect 19952 19068 20016 19072
rect 19952 19012 19956 19068
rect 19956 19012 20012 19068
rect 20012 19012 20016 19068
rect 19952 19008 20016 19012
rect 20032 19068 20096 19072
rect 20032 19012 20036 19068
rect 20036 19012 20092 19068
rect 20092 19012 20096 19068
rect 20032 19008 20096 19012
rect 20112 19068 20176 19072
rect 20112 19012 20116 19068
rect 20116 19012 20172 19068
rect 20172 19012 20176 19068
rect 20112 19008 20176 19012
rect 27646 19068 27710 19072
rect 27646 19012 27650 19068
rect 27650 19012 27706 19068
rect 27706 19012 27710 19068
rect 27646 19008 27710 19012
rect 27726 19068 27790 19072
rect 27726 19012 27730 19068
rect 27730 19012 27786 19068
rect 27786 19012 27790 19068
rect 27726 19008 27790 19012
rect 27806 19068 27870 19072
rect 27806 19012 27810 19068
rect 27810 19012 27866 19068
rect 27866 19012 27870 19068
rect 27806 19008 27870 19012
rect 27886 19068 27950 19072
rect 27886 19012 27890 19068
rect 27890 19012 27946 19068
rect 27946 19012 27950 19068
rect 27886 19008 27950 19012
rect 24716 18804 24780 18868
rect 5764 18532 5828 18596
rect 6684 18592 6748 18596
rect 6684 18536 6698 18592
rect 6698 18536 6748 18592
rect 6684 18532 6748 18536
rect 20300 18532 20364 18596
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 11438 18524 11502 18528
rect 11438 18468 11442 18524
rect 11442 18468 11498 18524
rect 11498 18468 11502 18524
rect 11438 18464 11502 18468
rect 11518 18524 11582 18528
rect 11518 18468 11522 18524
rect 11522 18468 11578 18524
rect 11578 18468 11582 18524
rect 11518 18464 11582 18468
rect 11598 18524 11662 18528
rect 11598 18468 11602 18524
rect 11602 18468 11658 18524
rect 11658 18468 11662 18524
rect 11598 18464 11662 18468
rect 11678 18524 11742 18528
rect 11678 18468 11682 18524
rect 11682 18468 11738 18524
rect 11738 18468 11742 18524
rect 11678 18464 11742 18468
rect 19212 18524 19276 18528
rect 19212 18468 19216 18524
rect 19216 18468 19272 18524
rect 19272 18468 19276 18524
rect 19212 18464 19276 18468
rect 19292 18524 19356 18528
rect 19292 18468 19296 18524
rect 19296 18468 19352 18524
rect 19352 18468 19356 18524
rect 19292 18464 19356 18468
rect 19372 18524 19436 18528
rect 19372 18468 19376 18524
rect 19376 18468 19432 18524
rect 19432 18468 19436 18524
rect 19372 18464 19436 18468
rect 19452 18524 19516 18528
rect 19452 18468 19456 18524
rect 19456 18468 19512 18524
rect 19512 18468 19516 18524
rect 19452 18464 19516 18468
rect 26986 18524 27050 18528
rect 26986 18468 26990 18524
rect 26990 18468 27046 18524
rect 27046 18468 27050 18524
rect 26986 18464 27050 18468
rect 27066 18524 27130 18528
rect 27066 18468 27070 18524
rect 27070 18468 27126 18524
rect 27126 18468 27130 18524
rect 27066 18464 27130 18468
rect 27146 18524 27210 18528
rect 27146 18468 27150 18524
rect 27150 18468 27206 18524
rect 27206 18468 27210 18524
rect 27146 18464 27210 18468
rect 27226 18524 27290 18528
rect 27226 18468 27230 18524
rect 27230 18468 27286 18524
rect 27286 18468 27290 18524
rect 27226 18464 27290 18468
rect 11836 18396 11900 18460
rect 29868 18396 29932 18460
rect 2636 18260 2700 18324
rect 4108 18124 4172 18188
rect 10180 18048 10244 18052
rect 10180 17992 10230 18048
rect 10230 17992 10244 18048
rect 10180 17988 10244 17992
rect 15516 17988 15580 18052
rect 26740 18124 26804 18188
rect 21956 17988 22020 18052
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 12098 17980 12162 17984
rect 12098 17924 12102 17980
rect 12102 17924 12158 17980
rect 12158 17924 12162 17980
rect 12098 17920 12162 17924
rect 12178 17980 12242 17984
rect 12178 17924 12182 17980
rect 12182 17924 12238 17980
rect 12238 17924 12242 17980
rect 12178 17920 12242 17924
rect 12258 17980 12322 17984
rect 12258 17924 12262 17980
rect 12262 17924 12318 17980
rect 12318 17924 12322 17980
rect 12258 17920 12322 17924
rect 12338 17980 12402 17984
rect 12338 17924 12342 17980
rect 12342 17924 12398 17980
rect 12398 17924 12402 17980
rect 12338 17920 12402 17924
rect 19872 17980 19936 17984
rect 19872 17924 19876 17980
rect 19876 17924 19932 17980
rect 19932 17924 19936 17980
rect 19872 17920 19936 17924
rect 19952 17980 20016 17984
rect 19952 17924 19956 17980
rect 19956 17924 20012 17980
rect 20012 17924 20016 17980
rect 19952 17920 20016 17924
rect 20032 17980 20096 17984
rect 20032 17924 20036 17980
rect 20036 17924 20092 17980
rect 20092 17924 20096 17980
rect 20032 17920 20096 17924
rect 20112 17980 20176 17984
rect 20112 17924 20116 17980
rect 20116 17924 20172 17980
rect 20172 17924 20176 17980
rect 20112 17920 20176 17924
rect 27646 17980 27710 17984
rect 27646 17924 27650 17980
rect 27650 17924 27706 17980
rect 27706 17924 27710 17980
rect 27646 17920 27710 17924
rect 27726 17980 27790 17984
rect 27726 17924 27730 17980
rect 27730 17924 27786 17980
rect 27786 17924 27790 17980
rect 27726 17920 27790 17924
rect 27806 17980 27870 17984
rect 27806 17924 27810 17980
rect 27810 17924 27866 17980
rect 27866 17924 27870 17980
rect 27806 17920 27870 17924
rect 27886 17980 27950 17984
rect 27886 17924 27890 17980
rect 27890 17924 27946 17980
rect 27946 17924 27950 17980
rect 27886 17920 27950 17924
rect 6316 17852 6380 17916
rect 11100 17852 11164 17916
rect 11836 17852 11900 17916
rect 26004 17852 26068 17916
rect 28396 17716 28460 17780
rect 8892 17580 8956 17644
rect 13860 17580 13924 17644
rect 14044 17580 14108 17644
rect 11836 17444 11900 17508
rect 12940 17444 13004 17508
rect 14412 17444 14476 17508
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 11438 17436 11502 17440
rect 11438 17380 11442 17436
rect 11442 17380 11498 17436
rect 11498 17380 11502 17436
rect 11438 17376 11502 17380
rect 11518 17436 11582 17440
rect 11518 17380 11522 17436
rect 11522 17380 11578 17436
rect 11578 17380 11582 17436
rect 11518 17376 11582 17380
rect 11598 17436 11662 17440
rect 11598 17380 11602 17436
rect 11602 17380 11658 17436
rect 11658 17380 11662 17436
rect 11598 17376 11662 17380
rect 11678 17436 11742 17440
rect 11678 17380 11682 17436
rect 11682 17380 11738 17436
rect 11738 17380 11742 17436
rect 11678 17376 11742 17380
rect 19212 17436 19276 17440
rect 19212 17380 19216 17436
rect 19216 17380 19272 17436
rect 19272 17380 19276 17436
rect 19212 17376 19276 17380
rect 19292 17436 19356 17440
rect 19292 17380 19296 17436
rect 19296 17380 19352 17436
rect 19352 17380 19356 17436
rect 19292 17376 19356 17380
rect 19372 17436 19436 17440
rect 19372 17380 19376 17436
rect 19376 17380 19432 17436
rect 19432 17380 19436 17436
rect 19372 17376 19436 17380
rect 19452 17436 19516 17440
rect 19452 17380 19456 17436
rect 19456 17380 19512 17436
rect 19512 17380 19516 17436
rect 19452 17376 19516 17380
rect 10548 17308 10612 17372
rect 14044 17172 14108 17236
rect 25820 17444 25884 17508
rect 26986 17436 27050 17440
rect 26986 17380 26990 17436
rect 26990 17380 27046 17436
rect 27046 17380 27050 17436
rect 26986 17376 27050 17380
rect 27066 17436 27130 17440
rect 27066 17380 27070 17436
rect 27070 17380 27126 17436
rect 27126 17380 27130 17436
rect 27066 17376 27130 17380
rect 27146 17436 27210 17440
rect 27146 17380 27150 17436
rect 27150 17380 27206 17436
rect 27206 17380 27210 17436
rect 27146 17376 27210 17380
rect 27226 17436 27290 17440
rect 27226 17380 27230 17436
rect 27230 17380 27286 17436
rect 27286 17380 27290 17436
rect 27226 17376 27290 17380
rect 28028 17308 28092 17372
rect 11100 17036 11164 17100
rect 12756 16960 12820 16964
rect 12756 16904 12770 16960
rect 12770 16904 12820 16960
rect 12756 16900 12820 16904
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 12098 16892 12162 16896
rect 12098 16836 12102 16892
rect 12102 16836 12158 16892
rect 12158 16836 12162 16892
rect 12098 16832 12162 16836
rect 12178 16892 12242 16896
rect 12178 16836 12182 16892
rect 12182 16836 12238 16892
rect 12238 16836 12242 16892
rect 12178 16832 12242 16836
rect 12258 16892 12322 16896
rect 12258 16836 12262 16892
rect 12262 16836 12318 16892
rect 12318 16836 12322 16892
rect 12258 16832 12322 16836
rect 12338 16892 12402 16896
rect 12338 16836 12342 16892
rect 12342 16836 12398 16892
rect 12398 16836 12402 16892
rect 12338 16832 12402 16836
rect 10916 16824 10980 16828
rect 10916 16768 10930 16824
rect 10930 16768 10980 16824
rect 10916 16764 10980 16768
rect 11836 16764 11900 16828
rect 5212 16628 5276 16692
rect 15148 16900 15212 16964
rect 19872 16892 19936 16896
rect 19872 16836 19876 16892
rect 19876 16836 19932 16892
rect 19932 16836 19936 16892
rect 19872 16832 19936 16836
rect 19952 16892 20016 16896
rect 19952 16836 19956 16892
rect 19956 16836 20012 16892
rect 20012 16836 20016 16892
rect 19952 16832 20016 16836
rect 20032 16892 20096 16896
rect 20032 16836 20036 16892
rect 20036 16836 20092 16892
rect 20092 16836 20096 16892
rect 20032 16832 20096 16836
rect 20112 16892 20176 16896
rect 20112 16836 20116 16892
rect 20116 16836 20172 16892
rect 20172 16836 20176 16892
rect 20112 16832 20176 16836
rect 15332 16628 15396 16692
rect 15884 16628 15948 16692
rect 16252 16628 16316 16692
rect 16804 16628 16868 16692
rect 18644 16764 18708 16828
rect 22692 17096 22756 17100
rect 22692 17040 22742 17096
rect 22742 17040 22756 17096
rect 22692 17036 22756 17040
rect 29500 17036 29564 17100
rect 22324 16764 22388 16828
rect 27646 16892 27710 16896
rect 27646 16836 27650 16892
rect 27650 16836 27706 16892
rect 27706 16836 27710 16892
rect 27646 16832 27710 16836
rect 27726 16892 27790 16896
rect 27726 16836 27730 16892
rect 27730 16836 27786 16892
rect 27786 16836 27790 16892
rect 27726 16832 27790 16836
rect 27806 16892 27870 16896
rect 27806 16836 27810 16892
rect 27810 16836 27866 16892
rect 27866 16836 27870 16892
rect 27806 16832 27870 16836
rect 27886 16892 27950 16896
rect 27886 16836 27890 16892
rect 27890 16836 27946 16892
rect 27946 16836 27950 16892
rect 27886 16832 27950 16836
rect 14596 16492 14660 16556
rect 22140 16552 22204 16556
rect 22140 16496 22154 16552
rect 22154 16496 22204 16552
rect 22140 16492 22204 16496
rect 22508 16492 22572 16556
rect 28396 16628 28460 16692
rect 26188 16552 26252 16556
rect 26188 16496 26238 16552
rect 26238 16496 26252 16552
rect 26188 16492 26252 16496
rect 29316 16552 29380 16556
rect 29316 16496 29330 16552
rect 29330 16496 29380 16552
rect 29316 16492 29380 16496
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 11438 16348 11502 16352
rect 11438 16292 11442 16348
rect 11442 16292 11498 16348
rect 11498 16292 11502 16348
rect 11438 16288 11502 16292
rect 11518 16348 11582 16352
rect 11518 16292 11522 16348
rect 11522 16292 11578 16348
rect 11578 16292 11582 16348
rect 11518 16288 11582 16292
rect 11598 16348 11662 16352
rect 11598 16292 11602 16348
rect 11602 16292 11658 16348
rect 11658 16292 11662 16348
rect 11598 16288 11662 16292
rect 11678 16348 11742 16352
rect 11678 16292 11682 16348
rect 11682 16292 11738 16348
rect 11738 16292 11742 16348
rect 11678 16288 11742 16292
rect 19212 16348 19276 16352
rect 19212 16292 19216 16348
rect 19216 16292 19272 16348
rect 19272 16292 19276 16348
rect 19212 16288 19276 16292
rect 19292 16348 19356 16352
rect 19292 16292 19296 16348
rect 19296 16292 19352 16348
rect 19352 16292 19356 16348
rect 19292 16288 19356 16292
rect 19372 16348 19436 16352
rect 19372 16292 19376 16348
rect 19376 16292 19432 16348
rect 19432 16292 19436 16348
rect 19372 16288 19436 16292
rect 19452 16348 19516 16352
rect 19452 16292 19456 16348
rect 19456 16292 19512 16348
rect 19512 16292 19516 16348
rect 19452 16288 19516 16292
rect 7236 16220 7300 16284
rect 10548 16220 10612 16284
rect 7420 16084 7484 16148
rect 21220 16220 21284 16284
rect 26188 16356 26252 16420
rect 28212 16356 28276 16420
rect 26986 16348 27050 16352
rect 26986 16292 26990 16348
rect 26990 16292 27046 16348
rect 27046 16292 27050 16348
rect 26986 16288 27050 16292
rect 27066 16348 27130 16352
rect 27066 16292 27070 16348
rect 27070 16292 27126 16348
rect 27126 16292 27130 16348
rect 27066 16288 27130 16292
rect 27146 16348 27210 16352
rect 27146 16292 27150 16348
rect 27150 16292 27206 16348
rect 27206 16292 27210 16348
rect 27146 16288 27210 16292
rect 27226 16348 27290 16352
rect 27226 16292 27230 16348
rect 27230 16292 27286 16348
rect 27286 16292 27290 16348
rect 27226 16288 27290 16292
rect 22324 16220 22388 16284
rect 8524 15812 8588 15876
rect 21772 15948 21836 16012
rect 22508 15948 22572 16012
rect 12572 15872 12636 15876
rect 12572 15816 12586 15872
rect 12586 15816 12636 15872
rect 12572 15812 12636 15816
rect 13124 15812 13188 15876
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 12098 15804 12162 15808
rect 12098 15748 12102 15804
rect 12102 15748 12158 15804
rect 12158 15748 12162 15804
rect 12098 15744 12162 15748
rect 12178 15804 12242 15808
rect 12178 15748 12182 15804
rect 12182 15748 12238 15804
rect 12238 15748 12242 15804
rect 12178 15744 12242 15748
rect 12258 15804 12322 15808
rect 12258 15748 12262 15804
rect 12262 15748 12318 15804
rect 12318 15748 12322 15804
rect 12258 15744 12322 15748
rect 12338 15804 12402 15808
rect 12338 15748 12342 15804
rect 12342 15748 12398 15804
rect 12398 15748 12402 15804
rect 12338 15744 12402 15748
rect 9260 15676 9324 15740
rect 19872 15804 19936 15808
rect 19872 15748 19876 15804
rect 19876 15748 19932 15804
rect 19932 15748 19936 15804
rect 19872 15744 19936 15748
rect 19952 15804 20016 15808
rect 19952 15748 19956 15804
rect 19956 15748 20012 15804
rect 20012 15748 20016 15804
rect 19952 15744 20016 15748
rect 20032 15804 20096 15808
rect 20032 15748 20036 15804
rect 20036 15748 20092 15804
rect 20092 15748 20096 15804
rect 20032 15744 20096 15748
rect 20112 15804 20176 15808
rect 20112 15748 20116 15804
rect 20116 15748 20172 15804
rect 20172 15748 20176 15804
rect 20112 15744 20176 15748
rect 8340 15600 8404 15604
rect 8340 15544 8390 15600
rect 8390 15544 8404 15600
rect 8340 15540 8404 15544
rect 8708 15540 8772 15604
rect 28028 15812 28092 15876
rect 27646 15804 27710 15808
rect 27646 15748 27650 15804
rect 27650 15748 27706 15804
rect 27706 15748 27710 15804
rect 27646 15744 27710 15748
rect 27726 15804 27790 15808
rect 27726 15748 27730 15804
rect 27730 15748 27786 15804
rect 27786 15748 27790 15804
rect 27726 15744 27790 15748
rect 27806 15804 27870 15808
rect 27806 15748 27810 15804
rect 27810 15748 27866 15804
rect 27866 15748 27870 15804
rect 27806 15744 27870 15748
rect 27886 15804 27950 15808
rect 27886 15748 27890 15804
rect 27890 15748 27946 15804
rect 27946 15748 27950 15804
rect 27886 15744 27950 15748
rect 26188 15676 26252 15740
rect 26372 15676 26436 15740
rect 21956 15540 22020 15604
rect 23060 15600 23124 15604
rect 23060 15544 23074 15600
rect 23074 15544 23124 15600
rect 23060 15540 23124 15544
rect 23244 15540 23308 15604
rect 28580 15540 28644 15604
rect 29132 15540 29196 15604
rect 21404 15404 21468 15468
rect 28028 15404 28092 15468
rect 28212 15404 28276 15468
rect 1164 15268 1228 15332
rect 11100 15268 11164 15332
rect 11836 15268 11900 15332
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 11438 15260 11502 15264
rect 11438 15204 11442 15260
rect 11442 15204 11498 15260
rect 11498 15204 11502 15260
rect 11438 15200 11502 15204
rect 11518 15260 11582 15264
rect 11518 15204 11522 15260
rect 11522 15204 11578 15260
rect 11578 15204 11582 15260
rect 11518 15200 11582 15204
rect 11598 15260 11662 15264
rect 11598 15204 11602 15260
rect 11602 15204 11658 15260
rect 11658 15204 11662 15260
rect 11598 15200 11662 15204
rect 11678 15260 11742 15264
rect 11678 15204 11682 15260
rect 11682 15204 11738 15260
rect 11738 15204 11742 15260
rect 11678 15200 11742 15204
rect 5764 15132 5828 15196
rect 7972 14996 8036 15060
rect 11284 15132 11348 15196
rect 13676 15268 13740 15332
rect 15700 15268 15764 15332
rect 27476 15268 27540 15332
rect 30236 15328 30300 15332
rect 30236 15272 30286 15328
rect 30286 15272 30300 15328
rect 30236 15268 30300 15272
rect 19212 15260 19276 15264
rect 19212 15204 19216 15260
rect 19216 15204 19272 15260
rect 19272 15204 19276 15260
rect 19212 15200 19276 15204
rect 19292 15260 19356 15264
rect 19292 15204 19296 15260
rect 19296 15204 19352 15260
rect 19352 15204 19356 15260
rect 19292 15200 19356 15204
rect 19372 15260 19436 15264
rect 19372 15204 19376 15260
rect 19376 15204 19432 15260
rect 19432 15204 19436 15260
rect 19372 15200 19436 15204
rect 19452 15260 19516 15264
rect 19452 15204 19456 15260
rect 19456 15204 19512 15260
rect 19512 15204 19516 15260
rect 19452 15200 19516 15204
rect 26986 15260 27050 15264
rect 26986 15204 26990 15260
rect 26990 15204 27046 15260
rect 27046 15204 27050 15260
rect 26986 15200 27050 15204
rect 27066 15260 27130 15264
rect 27066 15204 27070 15260
rect 27070 15204 27126 15260
rect 27126 15204 27130 15260
rect 27066 15200 27130 15204
rect 27146 15260 27210 15264
rect 27146 15204 27150 15260
rect 27150 15204 27206 15260
rect 27206 15204 27210 15260
rect 27146 15200 27210 15204
rect 27226 15260 27290 15264
rect 27226 15204 27230 15260
rect 27230 15204 27286 15260
rect 27286 15204 27290 15260
rect 27226 15200 27290 15204
rect 16436 15132 16500 15196
rect 25820 15192 25884 15196
rect 25820 15136 25870 15192
rect 25870 15136 25884 15192
rect 25820 15132 25884 15136
rect 7604 14860 7668 14924
rect 9812 14724 9876 14788
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 7604 14588 7668 14652
rect 12098 14716 12162 14720
rect 12098 14660 12102 14716
rect 12102 14660 12158 14716
rect 12158 14660 12162 14716
rect 12098 14656 12162 14660
rect 12178 14716 12242 14720
rect 12178 14660 12182 14716
rect 12182 14660 12238 14716
rect 12238 14660 12242 14716
rect 12178 14656 12242 14660
rect 12258 14716 12322 14720
rect 12258 14660 12262 14716
rect 12262 14660 12318 14716
rect 12318 14660 12322 14716
rect 12258 14656 12322 14660
rect 12338 14716 12402 14720
rect 12338 14660 12342 14716
rect 12342 14660 12398 14716
rect 12398 14660 12402 14716
rect 12338 14656 12402 14660
rect 8340 14512 8404 14516
rect 8340 14456 8390 14512
rect 8390 14456 8404 14512
rect 8340 14452 8404 14456
rect 20852 14724 20916 14788
rect 29868 14784 29932 14788
rect 29868 14728 29918 14784
rect 29918 14728 29932 14784
rect 29868 14724 29932 14728
rect 19872 14716 19936 14720
rect 19872 14660 19876 14716
rect 19876 14660 19932 14716
rect 19932 14660 19936 14716
rect 19872 14656 19936 14660
rect 19952 14716 20016 14720
rect 19952 14660 19956 14716
rect 19956 14660 20012 14716
rect 20012 14660 20016 14716
rect 19952 14656 20016 14660
rect 20032 14716 20096 14720
rect 20032 14660 20036 14716
rect 20036 14660 20092 14716
rect 20092 14660 20096 14716
rect 20032 14656 20096 14660
rect 20112 14716 20176 14720
rect 20112 14660 20116 14716
rect 20116 14660 20172 14716
rect 20172 14660 20176 14716
rect 20112 14656 20176 14660
rect 27646 14716 27710 14720
rect 27646 14660 27650 14716
rect 27650 14660 27706 14716
rect 27706 14660 27710 14716
rect 27646 14656 27710 14660
rect 27726 14716 27790 14720
rect 27726 14660 27730 14716
rect 27730 14660 27786 14716
rect 27786 14660 27790 14716
rect 27726 14656 27790 14660
rect 27806 14716 27870 14720
rect 27806 14660 27810 14716
rect 27810 14660 27866 14716
rect 27866 14660 27870 14716
rect 27806 14656 27870 14660
rect 27886 14716 27950 14720
rect 27886 14660 27890 14716
rect 27890 14660 27946 14716
rect 27946 14660 27950 14716
rect 27886 14656 27950 14660
rect 14044 14588 14108 14652
rect 18092 14588 18156 14652
rect 18828 14588 18892 14652
rect 20668 14588 20732 14652
rect 7236 14316 7300 14380
rect 8524 14376 8588 14380
rect 8524 14320 8574 14376
rect 8574 14320 8588 14376
rect 8524 14316 8588 14320
rect 24164 14452 24228 14516
rect 14964 14316 15028 14380
rect 26004 14316 26068 14380
rect 10732 14180 10796 14244
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 11438 14172 11502 14176
rect 11438 14116 11442 14172
rect 11442 14116 11498 14172
rect 11498 14116 11502 14172
rect 11438 14112 11502 14116
rect 11518 14172 11582 14176
rect 11518 14116 11522 14172
rect 11522 14116 11578 14172
rect 11578 14116 11582 14172
rect 11518 14112 11582 14116
rect 11598 14172 11662 14176
rect 11598 14116 11602 14172
rect 11602 14116 11658 14172
rect 11658 14116 11662 14172
rect 11598 14112 11662 14116
rect 11678 14172 11742 14176
rect 11678 14116 11682 14172
rect 11682 14116 11738 14172
rect 11738 14116 11742 14172
rect 11678 14112 11742 14116
rect 19212 14172 19276 14176
rect 19212 14116 19216 14172
rect 19216 14116 19272 14172
rect 19272 14116 19276 14172
rect 19212 14112 19276 14116
rect 19292 14172 19356 14176
rect 19292 14116 19296 14172
rect 19296 14116 19352 14172
rect 19352 14116 19356 14172
rect 19292 14112 19356 14116
rect 19372 14172 19436 14176
rect 19372 14116 19376 14172
rect 19376 14116 19432 14172
rect 19432 14116 19436 14172
rect 19372 14112 19436 14116
rect 19452 14172 19516 14176
rect 19452 14116 19456 14172
rect 19456 14116 19512 14172
rect 19512 14116 19516 14172
rect 19452 14112 19516 14116
rect 26986 14172 27050 14176
rect 26986 14116 26990 14172
rect 26990 14116 27046 14172
rect 27046 14116 27050 14172
rect 26986 14112 27050 14116
rect 27066 14172 27130 14176
rect 27066 14116 27070 14172
rect 27070 14116 27126 14172
rect 27126 14116 27130 14172
rect 27066 14112 27130 14116
rect 27146 14172 27210 14176
rect 27146 14116 27150 14172
rect 27150 14116 27206 14172
rect 27206 14116 27210 14172
rect 27146 14112 27210 14116
rect 27226 14172 27290 14176
rect 27226 14116 27230 14172
rect 27230 14116 27286 14172
rect 27286 14116 27290 14172
rect 27226 14112 27290 14116
rect 5764 13772 5828 13836
rect 6132 13636 6196 13700
rect 8708 13832 8772 13836
rect 8708 13776 8758 13832
rect 8758 13776 8772 13832
rect 8708 13772 8772 13776
rect 21772 13968 21836 13972
rect 21772 13912 21822 13968
rect 21822 13912 21836 13968
rect 21772 13908 21836 13912
rect 26740 13968 26804 13972
rect 26740 13912 26754 13968
rect 26754 13912 26804 13968
rect 26740 13908 26804 13912
rect 28764 13968 28828 13972
rect 28764 13912 28814 13968
rect 28814 13912 28828 13968
rect 28764 13908 28828 13912
rect 22140 13772 22204 13836
rect 24532 13832 24596 13836
rect 24532 13776 24546 13832
rect 24546 13776 24596 13832
rect 24532 13772 24596 13776
rect 29500 13772 29564 13836
rect 7972 13636 8036 13700
rect 10916 13636 10980 13700
rect 11836 13636 11900 13700
rect 12940 13636 13004 13700
rect 26740 13696 26804 13700
rect 26740 13640 26790 13696
rect 26790 13640 26804 13696
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 12098 13628 12162 13632
rect 12098 13572 12102 13628
rect 12102 13572 12158 13628
rect 12158 13572 12162 13628
rect 12098 13568 12162 13572
rect 12178 13628 12242 13632
rect 12178 13572 12182 13628
rect 12182 13572 12238 13628
rect 12238 13572 12242 13628
rect 12178 13568 12242 13572
rect 12258 13628 12322 13632
rect 12258 13572 12262 13628
rect 12262 13572 12318 13628
rect 12318 13572 12322 13628
rect 12258 13568 12322 13572
rect 12338 13628 12402 13632
rect 12338 13572 12342 13628
rect 12342 13572 12398 13628
rect 12398 13572 12402 13628
rect 12338 13568 12402 13572
rect 19872 13628 19936 13632
rect 19872 13572 19876 13628
rect 19876 13572 19932 13628
rect 19932 13572 19936 13628
rect 19872 13568 19936 13572
rect 19952 13628 20016 13632
rect 19952 13572 19956 13628
rect 19956 13572 20012 13628
rect 20012 13572 20016 13628
rect 19952 13568 20016 13572
rect 20032 13628 20096 13632
rect 20032 13572 20036 13628
rect 20036 13572 20092 13628
rect 20092 13572 20096 13628
rect 20032 13568 20096 13572
rect 20112 13628 20176 13632
rect 20112 13572 20116 13628
rect 20116 13572 20172 13628
rect 20172 13572 20176 13628
rect 20112 13568 20176 13572
rect 9444 13500 9508 13564
rect 10732 13500 10796 13564
rect 12940 13500 13004 13564
rect 13860 13500 13924 13564
rect 22324 13500 22388 13564
rect 24348 13500 24412 13564
rect 26740 13636 26804 13640
rect 27646 13628 27710 13632
rect 27646 13572 27650 13628
rect 27650 13572 27706 13628
rect 27706 13572 27710 13628
rect 27646 13568 27710 13572
rect 27726 13628 27790 13632
rect 27726 13572 27730 13628
rect 27730 13572 27786 13628
rect 27786 13572 27790 13628
rect 27726 13568 27790 13572
rect 27806 13628 27870 13632
rect 27806 13572 27810 13628
rect 27810 13572 27866 13628
rect 27866 13572 27870 13628
rect 27806 13568 27870 13572
rect 27886 13628 27950 13632
rect 27886 13572 27890 13628
rect 27890 13572 27946 13628
rect 27946 13572 27950 13628
rect 27886 13568 27950 13572
rect 8156 13092 8220 13156
rect 9628 13152 9692 13156
rect 19012 13228 19076 13292
rect 28212 13364 28276 13428
rect 9628 13096 9642 13152
rect 9642 13096 9692 13152
rect 9628 13092 9692 13096
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 11438 13084 11502 13088
rect 11438 13028 11442 13084
rect 11442 13028 11498 13084
rect 11498 13028 11502 13084
rect 11438 13024 11502 13028
rect 11518 13084 11582 13088
rect 11518 13028 11522 13084
rect 11522 13028 11578 13084
rect 11578 13028 11582 13084
rect 11518 13024 11582 13028
rect 11598 13084 11662 13088
rect 11598 13028 11602 13084
rect 11602 13028 11658 13084
rect 11658 13028 11662 13084
rect 11598 13024 11662 13028
rect 11678 13084 11742 13088
rect 11678 13028 11682 13084
rect 11682 13028 11738 13084
rect 11738 13028 11742 13084
rect 11678 13024 11742 13028
rect 5028 13016 5092 13020
rect 5028 12960 5078 13016
rect 5078 12960 5092 13016
rect 5028 12956 5092 12960
rect 3004 12820 3068 12884
rect 4844 12820 4908 12884
rect 17356 13092 17420 13156
rect 19212 13084 19276 13088
rect 19212 13028 19216 13084
rect 19216 13028 19272 13084
rect 19272 13028 19276 13084
rect 19212 13024 19276 13028
rect 19292 13084 19356 13088
rect 19292 13028 19296 13084
rect 19296 13028 19352 13084
rect 19352 13028 19356 13084
rect 19292 13024 19356 13028
rect 19372 13084 19436 13088
rect 19372 13028 19376 13084
rect 19376 13028 19432 13084
rect 19432 13028 19436 13084
rect 19372 13024 19436 13028
rect 19452 13084 19516 13088
rect 19452 13028 19456 13084
rect 19456 13028 19512 13084
rect 19512 13028 19516 13084
rect 19452 13024 19516 13028
rect 16620 12820 16684 12884
rect 18276 12820 18340 12884
rect 26986 13084 27050 13088
rect 26986 13028 26990 13084
rect 26990 13028 27046 13084
rect 27046 13028 27050 13084
rect 26986 13024 27050 13028
rect 27066 13084 27130 13088
rect 27066 13028 27070 13084
rect 27070 13028 27126 13084
rect 27126 13028 27130 13084
rect 27066 13024 27130 13028
rect 27146 13084 27210 13088
rect 27146 13028 27150 13084
rect 27150 13028 27206 13084
rect 27206 13028 27210 13084
rect 27146 13024 27210 13028
rect 27226 13084 27290 13088
rect 27226 13028 27230 13084
rect 27230 13028 27286 13084
rect 27286 13028 27290 13084
rect 27226 13024 27290 13028
rect 20668 12956 20732 13020
rect 25268 12956 25332 13020
rect 21036 12880 21100 12884
rect 21036 12824 21086 12880
rect 21086 12824 21100 12880
rect 21036 12820 21100 12824
rect 21956 12820 22020 12884
rect 22140 12880 22204 12884
rect 22140 12824 22190 12880
rect 22190 12824 22204 12880
rect 22140 12820 22204 12824
rect 26740 12820 26804 12884
rect 6500 12744 6564 12748
rect 6500 12688 6550 12744
rect 6550 12688 6564 12744
rect 6500 12684 6564 12688
rect 7788 12548 7852 12612
rect 13492 12744 13556 12748
rect 13492 12688 13542 12744
rect 13542 12688 13556 12744
rect 13492 12684 13556 12688
rect 14964 12684 15028 12748
rect 15884 12684 15948 12748
rect 11284 12608 11348 12612
rect 11284 12552 11334 12608
rect 11334 12552 11348 12608
rect 11284 12548 11348 12552
rect 16068 12548 16132 12612
rect 18460 12684 18524 12748
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 12098 12540 12162 12544
rect 12098 12484 12102 12540
rect 12102 12484 12158 12540
rect 12158 12484 12162 12540
rect 12098 12480 12162 12484
rect 12178 12540 12242 12544
rect 12178 12484 12182 12540
rect 12182 12484 12238 12540
rect 12238 12484 12242 12540
rect 12178 12480 12242 12484
rect 12258 12540 12322 12544
rect 12258 12484 12262 12540
rect 12262 12484 12318 12540
rect 12318 12484 12322 12540
rect 12258 12480 12322 12484
rect 12338 12540 12402 12544
rect 12338 12484 12342 12540
rect 12342 12484 12398 12540
rect 12398 12484 12402 12540
rect 12338 12480 12402 12484
rect 19872 12540 19936 12544
rect 19872 12484 19876 12540
rect 19876 12484 19932 12540
rect 19932 12484 19936 12540
rect 19872 12480 19936 12484
rect 19952 12540 20016 12544
rect 19952 12484 19956 12540
rect 19956 12484 20012 12540
rect 20012 12484 20016 12540
rect 19952 12480 20016 12484
rect 20032 12540 20096 12544
rect 20032 12484 20036 12540
rect 20036 12484 20092 12540
rect 20092 12484 20096 12540
rect 20032 12480 20096 12484
rect 20112 12540 20176 12544
rect 20112 12484 20116 12540
rect 20116 12484 20172 12540
rect 20172 12484 20176 12540
rect 20112 12480 20176 12484
rect 27646 12540 27710 12544
rect 27646 12484 27650 12540
rect 27650 12484 27706 12540
rect 27706 12484 27710 12540
rect 27646 12480 27710 12484
rect 27726 12540 27790 12544
rect 27726 12484 27730 12540
rect 27730 12484 27786 12540
rect 27786 12484 27790 12540
rect 27726 12480 27790 12484
rect 27806 12540 27870 12544
rect 27806 12484 27810 12540
rect 27810 12484 27866 12540
rect 27866 12484 27870 12540
rect 27806 12480 27870 12484
rect 27886 12540 27950 12544
rect 27886 12484 27890 12540
rect 27890 12484 27946 12540
rect 27946 12484 27950 12540
rect 27886 12480 27950 12484
rect 12940 12412 13004 12476
rect 14964 12276 15028 12340
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 7420 12140 7484 12204
rect 8892 12140 8956 12204
rect 9996 12140 10060 12204
rect 8156 12004 8220 12068
rect 9076 12064 9140 12068
rect 9076 12008 9126 12064
rect 9126 12008 9140 12064
rect 9076 12004 9140 12008
rect 10548 12004 10612 12068
rect 10916 12064 10980 12068
rect 14964 12140 15028 12204
rect 26004 12276 26068 12340
rect 29500 12412 29564 12476
rect 29132 12336 29196 12340
rect 29132 12280 29146 12336
rect 29146 12280 29196 12336
rect 29132 12276 29196 12280
rect 10916 12008 10930 12064
rect 10930 12008 10980 12064
rect 10916 12004 10980 12008
rect 11438 11996 11502 12000
rect 11438 11940 11442 11996
rect 11442 11940 11498 11996
rect 11498 11940 11502 11996
rect 11438 11936 11502 11940
rect 11518 11996 11582 12000
rect 11518 11940 11522 11996
rect 11522 11940 11578 11996
rect 11578 11940 11582 11996
rect 11518 11936 11582 11940
rect 11598 11996 11662 12000
rect 11598 11940 11602 11996
rect 11602 11940 11658 11996
rect 11658 11940 11662 11996
rect 11598 11936 11662 11940
rect 11678 11996 11742 12000
rect 11678 11940 11682 11996
rect 11682 11940 11738 11996
rect 11738 11940 11742 11996
rect 11678 11936 11742 11940
rect 7420 11868 7484 11932
rect 7788 11868 7852 11932
rect 17908 12140 17972 12204
rect 25636 12004 25700 12068
rect 19212 11996 19276 12000
rect 19212 11940 19216 11996
rect 19216 11940 19272 11996
rect 19272 11940 19276 11996
rect 19212 11936 19276 11940
rect 19292 11996 19356 12000
rect 19292 11940 19296 11996
rect 19296 11940 19352 11996
rect 19352 11940 19356 11996
rect 19292 11936 19356 11940
rect 19372 11996 19436 12000
rect 19372 11940 19376 11996
rect 19376 11940 19432 11996
rect 19432 11940 19436 11996
rect 19372 11936 19436 11940
rect 19452 11996 19516 12000
rect 19452 11940 19456 11996
rect 19456 11940 19512 11996
rect 19512 11940 19516 11996
rect 19452 11936 19516 11940
rect 20484 11928 20548 11932
rect 20484 11872 20534 11928
rect 20534 11872 20548 11928
rect 20484 11868 20548 11872
rect 21956 11868 22020 11932
rect 15516 11732 15580 11796
rect 18828 11732 18892 11796
rect 21220 11732 21284 11796
rect 26986 11996 27050 12000
rect 26986 11940 26990 11996
rect 26990 11940 27046 11996
rect 27046 11940 27050 11996
rect 26986 11936 27050 11940
rect 27066 11996 27130 12000
rect 27066 11940 27070 11996
rect 27070 11940 27126 11996
rect 27126 11940 27130 11996
rect 27066 11936 27130 11940
rect 27146 11996 27210 12000
rect 27146 11940 27150 11996
rect 27150 11940 27206 11996
rect 27206 11940 27210 11996
rect 27146 11936 27210 11940
rect 27226 11996 27290 12000
rect 27226 11940 27230 11996
rect 27230 11940 27286 11996
rect 27286 11940 27290 11996
rect 27226 11936 27290 11940
rect 28028 11868 28092 11932
rect 28396 11732 28460 11796
rect 8524 11460 8588 11524
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 12098 11452 12162 11456
rect 12098 11396 12102 11452
rect 12102 11396 12158 11452
rect 12158 11396 12162 11452
rect 12098 11392 12162 11396
rect 12178 11452 12242 11456
rect 12178 11396 12182 11452
rect 12182 11396 12238 11452
rect 12238 11396 12242 11452
rect 12178 11392 12242 11396
rect 12258 11452 12322 11456
rect 12258 11396 12262 11452
rect 12262 11396 12318 11452
rect 12318 11396 12322 11452
rect 12258 11392 12322 11396
rect 12338 11452 12402 11456
rect 12338 11396 12342 11452
rect 12342 11396 12398 11452
rect 12398 11396 12402 11452
rect 12338 11392 12402 11396
rect 3004 11248 3068 11252
rect 3004 11192 3018 11248
rect 3018 11192 3068 11248
rect 3004 11188 3068 11192
rect 3372 11188 3436 11252
rect 10548 11188 10612 11252
rect 11100 11188 11164 11252
rect 12572 11188 12636 11252
rect 14044 11460 14108 11524
rect 19702 11460 19766 11524
rect 20668 11460 20732 11524
rect 22876 11460 22940 11524
rect 26188 11460 26252 11524
rect 19872 11452 19936 11456
rect 19872 11396 19876 11452
rect 19876 11396 19932 11452
rect 19932 11396 19936 11452
rect 19872 11392 19936 11396
rect 19952 11452 20016 11456
rect 19952 11396 19956 11452
rect 19956 11396 20012 11452
rect 20012 11396 20016 11452
rect 19952 11392 20016 11396
rect 20032 11452 20096 11456
rect 20032 11396 20036 11452
rect 20036 11396 20092 11452
rect 20092 11396 20096 11452
rect 20032 11392 20096 11396
rect 20112 11452 20176 11456
rect 20112 11396 20116 11452
rect 20116 11396 20172 11452
rect 20172 11396 20176 11452
rect 20112 11392 20176 11396
rect 27646 11452 27710 11456
rect 27646 11396 27650 11452
rect 27650 11396 27706 11452
rect 27706 11396 27710 11452
rect 27646 11392 27710 11396
rect 27726 11452 27790 11456
rect 27726 11396 27730 11452
rect 27730 11396 27786 11452
rect 27786 11396 27790 11452
rect 27726 11392 27790 11396
rect 27806 11452 27870 11456
rect 27806 11396 27810 11452
rect 27810 11396 27866 11452
rect 27866 11396 27870 11452
rect 27806 11392 27870 11396
rect 27886 11452 27950 11456
rect 27886 11396 27890 11452
rect 27890 11396 27946 11452
rect 27946 11396 27950 11452
rect 27886 11392 27950 11396
rect 15516 11324 15580 11388
rect 16436 11324 16500 11388
rect 6684 11112 6748 11116
rect 6684 11056 6698 11112
rect 6698 11056 6748 11112
rect 6684 11052 6748 11056
rect 9076 11112 9140 11116
rect 9076 11056 9126 11112
rect 9126 11056 9140 11112
rect 9076 11052 9140 11056
rect 4844 10916 4908 10980
rect 12940 11112 13004 11116
rect 14596 11188 14660 11252
rect 26372 11324 26436 11388
rect 12940 11056 12954 11112
rect 12954 11056 13004 11112
rect 12940 11052 13004 11056
rect 26556 11052 26620 11116
rect 10548 10916 10612 10980
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 11438 10908 11502 10912
rect 11438 10852 11442 10908
rect 11442 10852 11498 10908
rect 11498 10852 11502 10908
rect 11438 10848 11502 10852
rect 11518 10908 11582 10912
rect 11518 10852 11522 10908
rect 11522 10852 11578 10908
rect 11578 10852 11582 10908
rect 11518 10848 11582 10852
rect 11598 10908 11662 10912
rect 11598 10852 11602 10908
rect 11602 10852 11658 10908
rect 11658 10852 11662 10908
rect 11598 10848 11662 10852
rect 11678 10908 11742 10912
rect 11678 10852 11682 10908
rect 11682 10852 11738 10908
rect 11738 10852 11742 10908
rect 11678 10848 11742 10852
rect 4844 10780 4908 10844
rect 9628 10780 9692 10844
rect 9444 10644 9508 10708
rect 13124 10916 13188 10980
rect 14044 10916 14108 10980
rect 14228 10916 14292 10980
rect 19702 10916 19766 10980
rect 19212 10908 19276 10912
rect 19212 10852 19216 10908
rect 19216 10852 19272 10908
rect 19272 10852 19276 10908
rect 19212 10848 19276 10852
rect 19292 10908 19356 10912
rect 19292 10852 19296 10908
rect 19296 10852 19352 10908
rect 19352 10852 19356 10908
rect 19292 10848 19356 10852
rect 19372 10908 19436 10912
rect 19372 10852 19376 10908
rect 19376 10852 19432 10908
rect 19432 10852 19436 10908
rect 19372 10848 19436 10852
rect 19452 10908 19516 10912
rect 19452 10852 19456 10908
rect 19456 10852 19512 10908
rect 19512 10852 19516 10908
rect 19452 10848 19516 10852
rect 26986 10908 27050 10912
rect 26986 10852 26990 10908
rect 26990 10852 27046 10908
rect 27046 10852 27050 10908
rect 26986 10848 27050 10852
rect 27066 10908 27130 10912
rect 27066 10852 27070 10908
rect 27070 10852 27126 10908
rect 27126 10852 27130 10908
rect 27066 10848 27130 10852
rect 27146 10908 27210 10912
rect 27146 10852 27150 10908
rect 27150 10852 27206 10908
rect 27206 10852 27210 10908
rect 27146 10848 27210 10852
rect 27226 10908 27290 10912
rect 27226 10852 27230 10908
rect 27230 10852 27286 10908
rect 27286 10852 27290 10908
rect 27226 10848 27290 10852
rect 2452 10508 2516 10572
rect 6132 10508 6196 10572
rect 5396 10372 5460 10436
rect 7788 10432 7852 10436
rect 7788 10376 7802 10432
rect 7802 10376 7852 10432
rect 7788 10372 7852 10376
rect 9996 10508 10060 10572
rect 20300 10780 20364 10844
rect 25084 10780 25148 10844
rect 18460 10644 18524 10708
rect 21588 10508 21652 10572
rect 14780 10372 14844 10436
rect 15884 10372 15948 10436
rect 20300 10372 20364 10436
rect 21036 10372 21100 10436
rect 30236 10508 30300 10572
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 12098 10364 12162 10368
rect 12098 10308 12102 10364
rect 12102 10308 12158 10364
rect 12158 10308 12162 10364
rect 12098 10304 12162 10308
rect 12178 10364 12242 10368
rect 12178 10308 12182 10364
rect 12182 10308 12238 10364
rect 12238 10308 12242 10364
rect 12178 10304 12242 10308
rect 12258 10364 12322 10368
rect 12258 10308 12262 10364
rect 12262 10308 12318 10364
rect 12318 10308 12322 10364
rect 12258 10304 12322 10308
rect 12338 10364 12402 10368
rect 12338 10308 12342 10364
rect 12342 10308 12398 10364
rect 12398 10308 12402 10364
rect 12338 10304 12402 10308
rect 19872 10364 19936 10368
rect 19872 10308 19876 10364
rect 19876 10308 19932 10364
rect 19932 10308 19936 10364
rect 19872 10304 19936 10308
rect 19952 10364 20016 10368
rect 19952 10308 19956 10364
rect 19956 10308 20012 10364
rect 20012 10308 20016 10364
rect 19952 10304 20016 10308
rect 20032 10364 20096 10368
rect 20032 10308 20036 10364
rect 20036 10308 20092 10364
rect 20092 10308 20096 10364
rect 20032 10304 20096 10308
rect 20112 10364 20176 10368
rect 20112 10308 20116 10364
rect 20116 10308 20172 10364
rect 20172 10308 20176 10364
rect 20112 10304 20176 10308
rect 27646 10364 27710 10368
rect 27646 10308 27650 10364
rect 27650 10308 27706 10364
rect 27706 10308 27710 10364
rect 27646 10304 27710 10308
rect 27726 10364 27790 10368
rect 27726 10308 27730 10364
rect 27730 10308 27786 10364
rect 27786 10308 27790 10364
rect 27726 10304 27790 10308
rect 27806 10364 27870 10368
rect 27806 10308 27810 10364
rect 27810 10308 27866 10364
rect 27866 10308 27870 10364
rect 27806 10304 27870 10308
rect 27886 10364 27950 10368
rect 27886 10308 27890 10364
rect 27890 10308 27946 10364
rect 27946 10308 27950 10364
rect 27886 10304 27950 10308
rect 4108 10236 4172 10300
rect 6316 10236 6380 10300
rect 9996 10236 10060 10300
rect 11284 10236 11348 10300
rect 17540 10236 17604 10300
rect 18828 10236 18892 10300
rect 21404 10236 21468 10300
rect 24900 10236 24964 10300
rect 14228 10100 14292 10164
rect 15148 10100 15212 10164
rect 9260 9828 9324 9892
rect 9812 9828 9876 9892
rect 10364 9828 10428 9892
rect 11100 9828 11164 9892
rect 12572 9828 12636 9892
rect 13860 9828 13924 9892
rect 14596 9828 14660 9892
rect 15516 9828 15580 9892
rect 16620 9828 16684 9892
rect 16988 9828 17052 9892
rect 18276 9888 18340 9892
rect 18276 9832 18290 9888
rect 18290 9832 18340 9888
rect 18276 9828 18340 9832
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 11438 9820 11502 9824
rect 11438 9764 11442 9820
rect 11442 9764 11498 9820
rect 11498 9764 11502 9820
rect 11438 9760 11502 9764
rect 11518 9820 11582 9824
rect 11518 9764 11522 9820
rect 11522 9764 11578 9820
rect 11578 9764 11582 9820
rect 11518 9760 11582 9764
rect 11598 9820 11662 9824
rect 11598 9764 11602 9820
rect 11602 9764 11658 9820
rect 11658 9764 11662 9820
rect 11598 9760 11662 9764
rect 11678 9820 11742 9824
rect 11678 9764 11682 9820
rect 11682 9764 11738 9820
rect 11738 9764 11742 9820
rect 11678 9760 11742 9764
rect 19212 9820 19276 9824
rect 19212 9764 19216 9820
rect 19216 9764 19272 9820
rect 19272 9764 19276 9820
rect 19212 9760 19276 9764
rect 19292 9820 19356 9824
rect 19292 9764 19296 9820
rect 19296 9764 19352 9820
rect 19352 9764 19356 9820
rect 19292 9760 19356 9764
rect 19372 9820 19436 9824
rect 19372 9764 19376 9820
rect 19376 9764 19432 9820
rect 19432 9764 19436 9820
rect 19372 9760 19436 9764
rect 19452 9820 19516 9824
rect 19452 9764 19456 9820
rect 19456 9764 19512 9820
rect 19512 9764 19516 9820
rect 19452 9760 19516 9764
rect 5764 9692 5828 9756
rect 11100 9692 11164 9756
rect 22692 9828 22756 9892
rect 24716 9828 24780 9892
rect 26986 9820 27050 9824
rect 26986 9764 26990 9820
rect 26990 9764 27046 9820
rect 27046 9764 27050 9820
rect 26986 9760 27050 9764
rect 27066 9820 27130 9824
rect 27066 9764 27070 9820
rect 27070 9764 27126 9820
rect 27126 9764 27130 9820
rect 27066 9760 27130 9764
rect 27146 9820 27210 9824
rect 27146 9764 27150 9820
rect 27150 9764 27206 9820
rect 27206 9764 27210 9820
rect 27146 9760 27210 9764
rect 27226 9820 27290 9824
rect 27226 9764 27230 9820
rect 27230 9764 27286 9820
rect 27286 9764 27290 9820
rect 27226 9760 27290 9764
rect 3004 9556 3068 9620
rect 6500 9556 6564 9620
rect 13492 9556 13556 9620
rect 3188 9284 3252 9348
rect 13124 9420 13188 9484
rect 12572 9344 12636 9348
rect 18644 9556 18708 9620
rect 22876 9556 22940 9620
rect 26556 9692 26620 9756
rect 25452 9556 25516 9620
rect 16804 9420 16868 9484
rect 29132 9420 29196 9484
rect 12572 9288 12622 9344
rect 12622 9288 12636 9344
rect 12572 9284 12636 9288
rect 13860 9284 13924 9348
rect 16620 9284 16684 9348
rect 17908 9284 17972 9348
rect 18460 9284 18524 9348
rect 29500 9284 29564 9348
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 12098 9276 12162 9280
rect 12098 9220 12102 9276
rect 12102 9220 12158 9276
rect 12158 9220 12162 9276
rect 12098 9216 12162 9220
rect 12178 9276 12242 9280
rect 12178 9220 12182 9276
rect 12182 9220 12238 9276
rect 12238 9220 12242 9276
rect 12178 9216 12242 9220
rect 12258 9276 12322 9280
rect 12258 9220 12262 9276
rect 12262 9220 12318 9276
rect 12318 9220 12322 9276
rect 12258 9216 12322 9220
rect 12338 9276 12402 9280
rect 12338 9220 12342 9276
rect 12342 9220 12398 9276
rect 12398 9220 12402 9276
rect 12338 9216 12402 9220
rect 19872 9276 19936 9280
rect 19872 9220 19876 9276
rect 19876 9220 19932 9276
rect 19932 9220 19936 9276
rect 19872 9216 19936 9220
rect 19952 9276 20016 9280
rect 19952 9220 19956 9276
rect 19956 9220 20012 9276
rect 20012 9220 20016 9276
rect 19952 9216 20016 9220
rect 20032 9276 20096 9280
rect 20032 9220 20036 9276
rect 20036 9220 20092 9276
rect 20092 9220 20096 9276
rect 20032 9216 20096 9220
rect 20112 9276 20176 9280
rect 20112 9220 20116 9276
rect 20116 9220 20172 9276
rect 20172 9220 20176 9276
rect 20112 9216 20176 9220
rect 27646 9276 27710 9280
rect 27646 9220 27650 9276
rect 27650 9220 27706 9276
rect 27706 9220 27710 9276
rect 27646 9216 27710 9220
rect 27726 9276 27790 9280
rect 27726 9220 27730 9276
rect 27730 9220 27786 9276
rect 27786 9220 27790 9276
rect 27726 9216 27790 9220
rect 27806 9276 27870 9280
rect 27806 9220 27810 9276
rect 27810 9220 27866 9276
rect 27866 9220 27870 9276
rect 27806 9216 27870 9220
rect 27886 9276 27950 9280
rect 27886 9220 27890 9276
rect 27890 9220 27946 9276
rect 27946 9220 27950 9276
rect 27886 9216 27950 9220
rect 26188 9148 26252 9212
rect 28396 9208 28460 9212
rect 28396 9152 28446 9208
rect 28446 9152 28460 9208
rect 28396 9148 28460 9152
rect 9260 9012 9324 9076
rect 11284 9012 11348 9076
rect 11836 9012 11900 9076
rect 13308 9012 13372 9076
rect 13860 9012 13924 9076
rect 16252 9012 16316 9076
rect 4108 8876 4172 8940
rect 4844 8876 4908 8940
rect 5212 8876 5276 8940
rect 14044 8876 14108 8940
rect 23060 9012 23124 9076
rect 25452 9012 25516 9076
rect 26740 9012 26804 9076
rect 30236 8876 30300 8940
rect 7604 8740 7668 8804
rect 8892 8740 8956 8804
rect 18644 8800 18708 8804
rect 18644 8744 18694 8800
rect 18694 8744 18708 8800
rect 18644 8740 18708 8744
rect 21036 8740 21100 8804
rect 22140 8740 22204 8804
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 11438 8732 11502 8736
rect 11438 8676 11442 8732
rect 11442 8676 11498 8732
rect 11498 8676 11502 8732
rect 11438 8672 11502 8676
rect 11518 8732 11582 8736
rect 11518 8676 11522 8732
rect 11522 8676 11578 8732
rect 11578 8676 11582 8732
rect 11518 8672 11582 8676
rect 11598 8732 11662 8736
rect 11598 8676 11602 8732
rect 11602 8676 11658 8732
rect 11658 8676 11662 8732
rect 11598 8672 11662 8676
rect 11678 8732 11742 8736
rect 11678 8676 11682 8732
rect 11682 8676 11738 8732
rect 11738 8676 11742 8732
rect 11678 8672 11742 8676
rect 19212 8732 19276 8736
rect 19212 8676 19216 8732
rect 19216 8676 19272 8732
rect 19272 8676 19276 8732
rect 19212 8672 19276 8676
rect 19292 8732 19356 8736
rect 19292 8676 19296 8732
rect 19296 8676 19352 8732
rect 19352 8676 19356 8732
rect 19292 8672 19356 8676
rect 19372 8732 19436 8736
rect 19372 8676 19376 8732
rect 19376 8676 19432 8732
rect 19432 8676 19436 8732
rect 19372 8672 19436 8676
rect 19452 8732 19516 8736
rect 19452 8676 19456 8732
rect 19456 8676 19512 8732
rect 19512 8676 19516 8732
rect 19452 8672 19516 8676
rect 5396 8468 5460 8532
rect 8524 8468 8588 8532
rect 13676 8604 13740 8668
rect 15332 8664 15396 8668
rect 15332 8608 15382 8664
rect 15382 8608 15396 8664
rect 15332 8604 15396 8608
rect 17540 8468 17604 8532
rect 25820 8604 25884 8668
rect 980 8392 1044 8396
rect 980 8336 1030 8392
rect 1030 8336 1044 8392
rect 980 8332 1044 8336
rect 5212 8332 5276 8396
rect 8340 8256 8404 8260
rect 8340 8200 8354 8256
rect 8354 8200 8404 8256
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 8340 8196 8404 8200
rect 26986 8732 27050 8736
rect 26986 8676 26990 8732
rect 26990 8676 27046 8732
rect 27046 8676 27050 8732
rect 26986 8672 27050 8676
rect 27066 8732 27130 8736
rect 27066 8676 27070 8732
rect 27070 8676 27126 8732
rect 27126 8676 27130 8732
rect 27066 8672 27130 8676
rect 27146 8732 27210 8736
rect 27146 8676 27150 8732
rect 27150 8676 27206 8732
rect 27206 8676 27210 8732
rect 27146 8672 27210 8676
rect 27226 8732 27290 8736
rect 27226 8676 27230 8732
rect 27230 8676 27286 8732
rect 27286 8676 27290 8732
rect 27226 8672 27290 8676
rect 23612 8332 23676 8396
rect 27476 8332 27540 8396
rect 29132 8332 29196 8396
rect 14596 8196 14660 8260
rect 14964 8256 15028 8260
rect 14964 8200 15014 8256
rect 15014 8200 15028 8256
rect 14964 8196 15028 8200
rect 21956 8196 22020 8260
rect 22508 8196 22572 8260
rect 23244 8256 23308 8260
rect 23244 8200 23294 8256
rect 23294 8200 23308 8256
rect 23244 8196 23308 8200
rect 12098 8188 12162 8192
rect 12098 8132 12102 8188
rect 12102 8132 12158 8188
rect 12158 8132 12162 8188
rect 12098 8128 12162 8132
rect 12178 8188 12242 8192
rect 12178 8132 12182 8188
rect 12182 8132 12238 8188
rect 12238 8132 12242 8188
rect 12178 8128 12242 8132
rect 12258 8188 12322 8192
rect 12258 8132 12262 8188
rect 12262 8132 12318 8188
rect 12318 8132 12322 8188
rect 12258 8128 12322 8132
rect 12338 8188 12402 8192
rect 12338 8132 12342 8188
rect 12342 8132 12398 8188
rect 12398 8132 12402 8188
rect 12338 8128 12402 8132
rect 19872 8188 19936 8192
rect 19872 8132 19876 8188
rect 19876 8132 19932 8188
rect 19932 8132 19936 8188
rect 19872 8128 19936 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 27646 8188 27710 8192
rect 27646 8132 27650 8188
rect 27650 8132 27706 8188
rect 27706 8132 27710 8188
rect 27646 8128 27710 8132
rect 27726 8188 27790 8192
rect 27726 8132 27730 8188
rect 27730 8132 27786 8188
rect 27786 8132 27790 8188
rect 27726 8128 27790 8132
rect 27806 8188 27870 8192
rect 27806 8132 27810 8188
rect 27810 8132 27866 8188
rect 27866 8132 27870 8188
rect 27806 8128 27870 8132
rect 27886 8188 27950 8192
rect 27886 8132 27890 8188
rect 27890 8132 27946 8188
rect 27946 8132 27950 8188
rect 27886 8128 27950 8132
rect 17356 8060 17420 8124
rect 18092 8060 18156 8124
rect 18460 8060 18524 8124
rect 19012 8120 19076 8124
rect 19012 8064 19026 8120
rect 19026 8064 19076 8120
rect 19012 8060 19076 8064
rect 22324 8060 22388 8124
rect 25820 8060 25884 8124
rect 26556 8060 26620 8124
rect 24716 7924 24780 7988
rect 16436 7788 16500 7852
rect 27476 7788 27540 7852
rect 24900 7652 24964 7716
rect 28212 7712 28276 7716
rect 28212 7656 28226 7712
rect 28226 7656 28276 7712
rect 28212 7652 28276 7656
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 11438 7644 11502 7648
rect 11438 7588 11442 7644
rect 11442 7588 11498 7644
rect 11498 7588 11502 7644
rect 11438 7584 11502 7588
rect 11518 7644 11582 7648
rect 11518 7588 11522 7644
rect 11522 7588 11578 7644
rect 11578 7588 11582 7644
rect 11518 7584 11582 7588
rect 11598 7644 11662 7648
rect 11598 7588 11602 7644
rect 11602 7588 11658 7644
rect 11658 7588 11662 7644
rect 11598 7584 11662 7588
rect 11678 7644 11742 7648
rect 11678 7588 11682 7644
rect 11682 7588 11738 7644
rect 11738 7588 11742 7644
rect 11678 7584 11742 7588
rect 19212 7644 19276 7648
rect 19212 7588 19216 7644
rect 19216 7588 19272 7644
rect 19272 7588 19276 7644
rect 19212 7584 19276 7588
rect 19292 7644 19356 7648
rect 19292 7588 19296 7644
rect 19296 7588 19352 7644
rect 19352 7588 19356 7644
rect 19292 7584 19356 7588
rect 19372 7644 19436 7648
rect 19372 7588 19376 7644
rect 19376 7588 19432 7644
rect 19432 7588 19436 7644
rect 19372 7584 19436 7588
rect 19452 7644 19516 7648
rect 19452 7588 19456 7644
rect 19456 7588 19512 7644
rect 19512 7588 19516 7644
rect 19452 7584 19516 7588
rect 26986 7644 27050 7648
rect 26986 7588 26990 7644
rect 26990 7588 27046 7644
rect 27046 7588 27050 7644
rect 26986 7584 27050 7588
rect 27066 7644 27130 7648
rect 27066 7588 27070 7644
rect 27070 7588 27126 7644
rect 27126 7588 27130 7644
rect 27066 7584 27130 7588
rect 27146 7644 27210 7648
rect 27146 7588 27150 7644
rect 27150 7588 27206 7644
rect 27206 7588 27210 7644
rect 27146 7584 27210 7588
rect 27226 7644 27290 7648
rect 27226 7588 27230 7644
rect 27230 7588 27286 7644
rect 27286 7588 27290 7644
rect 27226 7584 27290 7588
rect 5028 7516 5092 7580
rect 8708 7516 8772 7580
rect 9444 7516 9508 7580
rect 18276 7516 18340 7580
rect 20300 7576 20364 7580
rect 20300 7520 20350 7576
rect 20350 7520 20364 7576
rect 20300 7516 20364 7520
rect 14780 7244 14844 7308
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 12098 7100 12162 7104
rect 12098 7044 12102 7100
rect 12102 7044 12158 7100
rect 12158 7044 12162 7100
rect 12098 7040 12162 7044
rect 12178 7100 12242 7104
rect 12178 7044 12182 7100
rect 12182 7044 12238 7100
rect 12238 7044 12242 7100
rect 12178 7040 12242 7044
rect 12258 7100 12322 7104
rect 12258 7044 12262 7100
rect 12262 7044 12318 7100
rect 12318 7044 12322 7100
rect 12258 7040 12322 7044
rect 12338 7100 12402 7104
rect 12338 7044 12342 7100
rect 12342 7044 12398 7100
rect 12398 7044 12402 7100
rect 12338 7040 12402 7044
rect 9628 6972 9692 7036
rect 19872 7100 19936 7104
rect 19872 7044 19876 7100
rect 19876 7044 19932 7100
rect 19932 7044 19936 7100
rect 19872 7040 19936 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 16988 7032 17052 7036
rect 16988 6976 17002 7032
rect 17002 6976 17052 7032
rect 16988 6972 17052 6976
rect 27646 7100 27710 7104
rect 27646 7044 27650 7100
rect 27650 7044 27706 7100
rect 27706 7044 27710 7100
rect 27646 7040 27710 7044
rect 27726 7100 27790 7104
rect 27726 7044 27730 7100
rect 27730 7044 27786 7100
rect 27786 7044 27790 7100
rect 27726 7040 27790 7044
rect 27806 7100 27870 7104
rect 27806 7044 27810 7100
rect 27810 7044 27866 7100
rect 27866 7044 27870 7100
rect 27806 7040 27870 7044
rect 27886 7100 27950 7104
rect 27886 7044 27890 7100
rect 27890 7044 27946 7100
rect 27946 7044 27950 7100
rect 27886 7040 27950 7044
rect 27476 6972 27540 7036
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 20484 6836 20548 6900
rect 24532 6836 24596 6900
rect 10732 6564 10796 6628
rect 12572 6564 12636 6628
rect 11438 6556 11502 6560
rect 11438 6500 11442 6556
rect 11442 6500 11498 6556
rect 11498 6500 11502 6556
rect 11438 6496 11502 6500
rect 11518 6556 11582 6560
rect 11518 6500 11522 6556
rect 11522 6500 11578 6556
rect 11578 6500 11582 6556
rect 11518 6496 11582 6500
rect 11598 6556 11662 6560
rect 11598 6500 11602 6556
rect 11602 6500 11658 6556
rect 11658 6500 11662 6556
rect 11598 6496 11662 6500
rect 11678 6556 11742 6560
rect 11678 6500 11682 6556
rect 11682 6500 11738 6556
rect 11738 6500 11742 6556
rect 11678 6496 11742 6500
rect 19212 6556 19276 6560
rect 19212 6500 19216 6556
rect 19216 6500 19272 6556
rect 19272 6500 19276 6556
rect 19212 6496 19276 6500
rect 19292 6556 19356 6560
rect 19292 6500 19296 6556
rect 19296 6500 19352 6556
rect 19352 6500 19356 6556
rect 19292 6496 19356 6500
rect 19372 6556 19436 6560
rect 19372 6500 19376 6556
rect 19376 6500 19432 6556
rect 19432 6500 19436 6556
rect 19372 6496 19436 6500
rect 19452 6556 19516 6560
rect 19452 6500 19456 6556
rect 19456 6500 19512 6556
rect 19512 6500 19516 6556
rect 19452 6496 19516 6500
rect 26986 6556 27050 6560
rect 26986 6500 26990 6556
rect 26990 6500 27046 6556
rect 27046 6500 27050 6556
rect 26986 6496 27050 6500
rect 27066 6556 27130 6560
rect 27066 6500 27070 6556
rect 27070 6500 27126 6556
rect 27126 6500 27130 6556
rect 27066 6496 27130 6500
rect 27146 6556 27210 6560
rect 27146 6500 27150 6556
rect 27150 6500 27206 6556
rect 27206 6500 27210 6556
rect 27146 6496 27210 6500
rect 27226 6556 27290 6560
rect 27226 6500 27230 6556
rect 27230 6500 27286 6556
rect 27286 6500 27290 6556
rect 27226 6496 27290 6500
rect 12940 6428 13004 6492
rect 18644 6428 18708 6492
rect 5396 6292 5460 6356
rect 11100 6352 11164 6356
rect 11100 6296 11114 6352
rect 11114 6296 11164 6352
rect 11100 6292 11164 6296
rect 16620 6292 16684 6356
rect 21036 6292 21100 6356
rect 10364 6156 10428 6220
rect 7972 6080 8036 6084
rect 7972 6024 8022 6080
rect 8022 6024 8036 6080
rect 7972 6020 8036 6024
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 12098 6012 12162 6016
rect 12098 5956 12102 6012
rect 12102 5956 12158 6012
rect 12158 5956 12162 6012
rect 12098 5952 12162 5956
rect 12178 6012 12242 6016
rect 12178 5956 12182 6012
rect 12182 5956 12238 6012
rect 12238 5956 12242 6012
rect 12178 5952 12242 5956
rect 12258 6012 12322 6016
rect 12258 5956 12262 6012
rect 12262 5956 12318 6012
rect 12318 5956 12322 6012
rect 12258 5952 12322 5956
rect 12338 6012 12402 6016
rect 12338 5956 12342 6012
rect 12342 5956 12398 6012
rect 12398 5956 12402 6012
rect 12338 5952 12402 5956
rect 19872 6012 19936 6016
rect 19872 5956 19876 6012
rect 19876 5956 19932 6012
rect 19932 5956 19936 6012
rect 19872 5952 19936 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 10548 5884 10612 5948
rect 15516 5884 15580 5948
rect 27646 6012 27710 6016
rect 27646 5956 27650 6012
rect 27650 5956 27706 6012
rect 27706 5956 27710 6012
rect 27646 5952 27710 5956
rect 27726 6012 27790 6016
rect 27726 5956 27730 6012
rect 27730 5956 27786 6012
rect 27786 5956 27790 6012
rect 27726 5952 27790 5956
rect 27806 6012 27870 6016
rect 27806 5956 27810 6012
rect 27810 5956 27866 6012
rect 27866 5956 27870 6012
rect 27806 5952 27870 5956
rect 27886 6012 27950 6016
rect 27886 5956 27890 6012
rect 27890 5956 27946 6012
rect 27946 5956 27950 6012
rect 27886 5952 27950 5956
rect 8156 5748 8220 5812
rect 2452 5672 2516 5676
rect 2452 5616 2502 5672
rect 2502 5616 2516 5672
rect 2452 5612 2516 5616
rect 8156 5612 8220 5676
rect 4108 5476 4172 5540
rect 7788 5476 7852 5540
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 11438 5468 11502 5472
rect 11438 5412 11442 5468
rect 11442 5412 11498 5468
rect 11498 5412 11502 5468
rect 11438 5408 11502 5412
rect 11518 5468 11582 5472
rect 11518 5412 11522 5468
rect 11522 5412 11578 5468
rect 11578 5412 11582 5468
rect 11518 5408 11582 5412
rect 11598 5468 11662 5472
rect 11598 5412 11602 5468
rect 11602 5412 11658 5468
rect 11658 5412 11662 5468
rect 11598 5408 11662 5412
rect 11678 5468 11742 5472
rect 11678 5412 11682 5468
rect 11682 5412 11738 5468
rect 11738 5412 11742 5468
rect 11678 5408 11742 5412
rect 25084 5612 25148 5676
rect 15148 5476 15212 5540
rect 18828 5476 18892 5540
rect 19212 5468 19276 5472
rect 19212 5412 19216 5468
rect 19216 5412 19272 5468
rect 19272 5412 19276 5468
rect 19212 5408 19276 5412
rect 19292 5468 19356 5472
rect 19292 5412 19296 5468
rect 19296 5412 19352 5468
rect 19352 5412 19356 5468
rect 19292 5408 19356 5412
rect 19372 5468 19436 5472
rect 19372 5412 19376 5468
rect 19376 5412 19432 5468
rect 19432 5412 19436 5468
rect 19372 5408 19436 5412
rect 19452 5468 19516 5472
rect 19452 5412 19456 5468
rect 19456 5412 19512 5468
rect 19512 5412 19516 5468
rect 19452 5408 19516 5412
rect 26986 5468 27050 5472
rect 26986 5412 26990 5468
rect 26990 5412 27046 5468
rect 27046 5412 27050 5468
rect 26986 5408 27050 5412
rect 27066 5468 27130 5472
rect 27066 5412 27070 5468
rect 27070 5412 27126 5468
rect 27126 5412 27130 5468
rect 27066 5408 27130 5412
rect 27146 5468 27210 5472
rect 27146 5412 27150 5468
rect 27150 5412 27206 5468
rect 27206 5412 27210 5468
rect 27146 5408 27210 5412
rect 27226 5468 27290 5472
rect 27226 5412 27230 5468
rect 27230 5412 27286 5468
rect 27286 5412 27290 5468
rect 27226 5408 27290 5412
rect 20300 5340 20364 5404
rect 28580 5128 28644 5132
rect 28580 5072 28594 5128
rect 28594 5072 28644 5128
rect 28580 5068 28644 5072
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 12098 4924 12162 4928
rect 12098 4868 12102 4924
rect 12102 4868 12158 4924
rect 12158 4868 12162 4924
rect 12098 4864 12162 4868
rect 12178 4924 12242 4928
rect 12178 4868 12182 4924
rect 12182 4868 12238 4924
rect 12238 4868 12242 4924
rect 12178 4864 12242 4868
rect 12258 4924 12322 4928
rect 12258 4868 12262 4924
rect 12262 4868 12318 4924
rect 12318 4868 12322 4924
rect 12258 4864 12322 4868
rect 12338 4924 12402 4928
rect 12338 4868 12342 4924
rect 12342 4868 12398 4924
rect 12398 4868 12402 4924
rect 12338 4864 12402 4868
rect 19872 4924 19936 4928
rect 19872 4868 19876 4924
rect 19876 4868 19932 4924
rect 19932 4868 19936 4924
rect 19872 4864 19936 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 27646 4924 27710 4928
rect 27646 4868 27650 4924
rect 27650 4868 27706 4924
rect 27706 4868 27710 4924
rect 27646 4864 27710 4868
rect 27726 4924 27790 4928
rect 27726 4868 27730 4924
rect 27730 4868 27786 4924
rect 27786 4868 27790 4924
rect 27726 4864 27790 4868
rect 27806 4924 27870 4928
rect 27806 4868 27810 4924
rect 27810 4868 27866 4924
rect 27866 4868 27870 4924
rect 27806 4864 27870 4868
rect 27886 4924 27950 4928
rect 27886 4868 27890 4924
rect 27890 4868 27946 4924
rect 27946 4868 27950 4924
rect 27886 4864 27950 4868
rect 10180 4796 10244 4860
rect 15700 4856 15764 4860
rect 15700 4800 15750 4856
rect 15750 4800 15764 4856
rect 15700 4796 15764 4800
rect 20852 4856 20916 4860
rect 20852 4800 20866 4856
rect 20866 4800 20916 4856
rect 20852 4796 20916 4800
rect 3188 4660 3252 4724
rect 15148 4660 15212 4724
rect 10916 4524 10980 4588
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 11438 4380 11502 4384
rect 11438 4324 11442 4380
rect 11442 4324 11498 4380
rect 11498 4324 11502 4380
rect 11438 4320 11502 4324
rect 11518 4380 11582 4384
rect 11518 4324 11522 4380
rect 11522 4324 11578 4380
rect 11578 4324 11582 4380
rect 11518 4320 11582 4324
rect 11598 4380 11662 4384
rect 11598 4324 11602 4380
rect 11602 4324 11658 4380
rect 11658 4324 11662 4380
rect 11598 4320 11662 4324
rect 11678 4380 11742 4384
rect 11678 4324 11682 4380
rect 11682 4324 11738 4380
rect 11738 4324 11742 4380
rect 11678 4320 11742 4324
rect 19212 4380 19276 4384
rect 19212 4324 19216 4380
rect 19216 4324 19272 4380
rect 19272 4324 19276 4380
rect 19212 4320 19276 4324
rect 19292 4380 19356 4384
rect 19292 4324 19296 4380
rect 19296 4324 19352 4380
rect 19352 4324 19356 4380
rect 19292 4320 19356 4324
rect 19372 4380 19436 4384
rect 19372 4324 19376 4380
rect 19376 4324 19432 4380
rect 19432 4324 19436 4380
rect 19372 4320 19436 4324
rect 19452 4380 19516 4384
rect 19452 4324 19456 4380
rect 19456 4324 19512 4380
rect 19512 4324 19516 4380
rect 19452 4320 19516 4324
rect 26986 4380 27050 4384
rect 26986 4324 26990 4380
rect 26990 4324 27046 4380
rect 27046 4324 27050 4380
rect 26986 4320 27050 4324
rect 27066 4380 27130 4384
rect 27066 4324 27070 4380
rect 27070 4324 27126 4380
rect 27126 4324 27130 4380
rect 27066 4320 27130 4324
rect 27146 4380 27210 4384
rect 27146 4324 27150 4380
rect 27150 4324 27206 4380
rect 27206 4324 27210 4380
rect 27146 4320 27210 4324
rect 27226 4380 27290 4384
rect 27226 4324 27230 4380
rect 27230 4324 27286 4380
rect 27286 4324 27290 4380
rect 27226 4320 27290 4324
rect 3188 4116 3252 4180
rect 21772 4176 21836 4180
rect 21772 4120 21822 4176
rect 21822 4120 21836 4176
rect 21772 4116 21836 4120
rect 2636 3980 2700 4044
rect 11284 3844 11348 3908
rect 26188 3980 26252 4044
rect 16068 3844 16132 3908
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 12098 3836 12162 3840
rect 12098 3780 12102 3836
rect 12102 3780 12158 3836
rect 12158 3780 12162 3836
rect 12098 3776 12162 3780
rect 12178 3836 12242 3840
rect 12178 3780 12182 3836
rect 12182 3780 12238 3836
rect 12238 3780 12242 3836
rect 12178 3776 12242 3780
rect 12258 3836 12322 3840
rect 12258 3780 12262 3836
rect 12262 3780 12318 3836
rect 12318 3780 12322 3836
rect 12258 3776 12322 3780
rect 12338 3836 12402 3840
rect 12338 3780 12342 3836
rect 12342 3780 12398 3836
rect 12398 3780 12402 3836
rect 12338 3776 12402 3780
rect 19872 3836 19936 3840
rect 19872 3780 19876 3836
rect 19876 3780 19932 3836
rect 19932 3780 19936 3836
rect 19872 3776 19936 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 27646 3836 27710 3840
rect 27646 3780 27650 3836
rect 27650 3780 27706 3836
rect 27706 3780 27710 3836
rect 27646 3776 27710 3780
rect 27726 3836 27790 3840
rect 27726 3780 27730 3836
rect 27730 3780 27786 3836
rect 27786 3780 27790 3836
rect 27726 3776 27790 3780
rect 27806 3836 27870 3840
rect 27806 3780 27810 3836
rect 27810 3780 27866 3836
rect 27866 3780 27870 3836
rect 27806 3776 27870 3780
rect 27886 3836 27950 3840
rect 27886 3780 27890 3836
rect 27890 3780 27946 3836
rect 27946 3780 27950 3836
rect 27886 3776 27950 3780
rect 12756 3708 12820 3772
rect 2452 3572 2516 3636
rect 14412 3632 14476 3636
rect 14412 3576 14426 3632
rect 14426 3576 14476 3632
rect 14412 3572 14476 3576
rect 8156 3436 8220 3500
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 11438 3292 11502 3296
rect 11438 3236 11442 3292
rect 11442 3236 11498 3292
rect 11498 3236 11502 3292
rect 11438 3232 11502 3236
rect 11518 3292 11582 3296
rect 11518 3236 11522 3292
rect 11522 3236 11578 3292
rect 11578 3236 11582 3292
rect 11518 3232 11582 3236
rect 11598 3292 11662 3296
rect 11598 3236 11602 3292
rect 11602 3236 11658 3292
rect 11658 3236 11662 3292
rect 11598 3232 11662 3236
rect 11678 3292 11742 3296
rect 11678 3236 11682 3292
rect 11682 3236 11738 3292
rect 11738 3236 11742 3292
rect 11678 3232 11742 3236
rect 19212 3292 19276 3296
rect 19212 3236 19216 3292
rect 19216 3236 19272 3292
rect 19272 3236 19276 3292
rect 19212 3232 19276 3236
rect 19292 3292 19356 3296
rect 19292 3236 19296 3292
rect 19296 3236 19352 3292
rect 19352 3236 19356 3292
rect 19292 3232 19356 3236
rect 19372 3292 19436 3296
rect 19372 3236 19376 3292
rect 19376 3236 19432 3292
rect 19432 3236 19436 3292
rect 19372 3232 19436 3236
rect 19452 3292 19516 3296
rect 19452 3236 19456 3292
rect 19456 3236 19512 3292
rect 19512 3236 19516 3292
rect 19452 3232 19516 3236
rect 26986 3292 27050 3296
rect 26986 3236 26990 3292
rect 26990 3236 27046 3292
rect 27046 3236 27050 3292
rect 26986 3232 27050 3236
rect 27066 3292 27130 3296
rect 27066 3236 27070 3292
rect 27070 3236 27126 3292
rect 27126 3236 27130 3292
rect 27066 3232 27130 3236
rect 27146 3292 27210 3296
rect 27146 3236 27150 3292
rect 27150 3236 27206 3292
rect 27206 3236 27210 3292
rect 27146 3232 27210 3236
rect 27226 3292 27290 3296
rect 27226 3236 27230 3292
rect 27230 3236 27286 3292
rect 27286 3236 27290 3292
rect 27226 3232 27290 3236
rect 7972 3028 8036 3092
rect 13860 2892 13924 2956
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 12098 2748 12162 2752
rect 12098 2692 12102 2748
rect 12102 2692 12158 2748
rect 12158 2692 12162 2748
rect 12098 2688 12162 2692
rect 12178 2748 12242 2752
rect 12178 2692 12182 2748
rect 12182 2692 12238 2748
rect 12238 2692 12242 2748
rect 12178 2688 12242 2692
rect 12258 2748 12322 2752
rect 12258 2692 12262 2748
rect 12262 2692 12318 2748
rect 12318 2692 12322 2748
rect 12258 2688 12322 2692
rect 12338 2748 12402 2752
rect 12338 2692 12342 2748
rect 12342 2692 12398 2748
rect 12398 2692 12402 2748
rect 12338 2688 12402 2692
rect 19872 2748 19936 2752
rect 19872 2692 19876 2748
rect 19876 2692 19932 2748
rect 19932 2692 19936 2748
rect 19872 2688 19936 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 27646 2748 27710 2752
rect 27646 2692 27650 2748
rect 27650 2692 27706 2748
rect 27706 2692 27710 2748
rect 27646 2688 27710 2692
rect 27726 2748 27790 2752
rect 27726 2692 27730 2748
rect 27730 2692 27786 2748
rect 27786 2692 27790 2748
rect 27726 2688 27790 2692
rect 27806 2748 27870 2752
rect 27806 2692 27810 2748
rect 27810 2692 27866 2748
rect 27866 2692 27870 2748
rect 27806 2688 27870 2692
rect 27886 2748 27950 2752
rect 27886 2692 27890 2748
rect 27890 2692 27946 2748
rect 27946 2692 27950 2748
rect 27886 2688 27950 2692
rect 25636 2620 25700 2684
rect 21220 2484 21284 2548
rect 13124 2348 13188 2412
rect 20668 2348 20732 2412
rect 23612 2212 23676 2276
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 11438 2204 11502 2208
rect 11438 2148 11442 2204
rect 11442 2148 11498 2204
rect 11498 2148 11502 2204
rect 11438 2144 11502 2148
rect 11518 2204 11582 2208
rect 11518 2148 11522 2204
rect 11522 2148 11578 2204
rect 11578 2148 11582 2204
rect 11518 2144 11582 2148
rect 11598 2204 11662 2208
rect 11598 2148 11602 2204
rect 11602 2148 11658 2204
rect 11658 2148 11662 2204
rect 11598 2144 11662 2148
rect 11678 2204 11742 2208
rect 11678 2148 11682 2204
rect 11682 2148 11738 2204
rect 11738 2148 11742 2204
rect 11678 2144 11742 2148
rect 19212 2204 19276 2208
rect 19212 2148 19216 2204
rect 19216 2148 19272 2204
rect 19272 2148 19276 2204
rect 19212 2144 19276 2148
rect 19292 2204 19356 2208
rect 19292 2148 19296 2204
rect 19296 2148 19352 2204
rect 19352 2148 19356 2204
rect 19292 2144 19356 2148
rect 19372 2204 19436 2208
rect 19372 2148 19376 2204
rect 19376 2148 19432 2204
rect 19432 2148 19436 2204
rect 19372 2144 19436 2148
rect 19452 2204 19516 2208
rect 19452 2148 19456 2204
rect 19456 2148 19512 2204
rect 19512 2148 19516 2204
rect 19452 2144 19516 2148
rect 26986 2204 27050 2208
rect 26986 2148 26990 2204
rect 26990 2148 27046 2204
rect 27046 2148 27050 2204
rect 26986 2144 27050 2148
rect 27066 2204 27130 2208
rect 27066 2148 27070 2204
rect 27070 2148 27126 2204
rect 27126 2148 27130 2204
rect 27066 2144 27130 2148
rect 27146 2204 27210 2208
rect 27146 2148 27150 2204
rect 27150 2148 27206 2204
rect 27206 2148 27210 2204
rect 27146 2144 27210 2148
rect 27226 2204 27290 2208
rect 27226 2148 27230 2204
rect 27230 2148 27286 2204
rect 27286 2148 27290 2204
rect 27226 2144 27290 2148
rect 13308 1940 13372 2004
rect 1164 1804 1228 1868
rect 21588 1804 21652 1868
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 12098 1660 12162 1664
rect 12098 1604 12102 1660
rect 12102 1604 12158 1660
rect 12158 1604 12162 1660
rect 12098 1600 12162 1604
rect 12178 1660 12242 1664
rect 12178 1604 12182 1660
rect 12182 1604 12238 1660
rect 12238 1604 12242 1660
rect 12178 1600 12242 1604
rect 12258 1660 12322 1664
rect 12258 1604 12262 1660
rect 12262 1604 12318 1660
rect 12318 1604 12322 1660
rect 12258 1600 12322 1604
rect 12338 1660 12402 1664
rect 12338 1604 12342 1660
rect 12342 1604 12398 1660
rect 12398 1604 12402 1660
rect 12338 1600 12402 1604
rect 19872 1660 19936 1664
rect 19872 1604 19876 1660
rect 19876 1604 19932 1660
rect 19932 1604 19936 1660
rect 19872 1600 19936 1604
rect 19952 1660 20016 1664
rect 19952 1604 19956 1660
rect 19956 1604 20012 1660
rect 20012 1604 20016 1660
rect 19952 1600 20016 1604
rect 20032 1660 20096 1664
rect 20032 1604 20036 1660
rect 20036 1604 20092 1660
rect 20092 1604 20096 1660
rect 20032 1600 20096 1604
rect 20112 1660 20176 1664
rect 20112 1604 20116 1660
rect 20116 1604 20172 1660
rect 20172 1604 20176 1660
rect 20112 1600 20176 1604
rect 27646 1660 27710 1664
rect 27646 1604 27650 1660
rect 27650 1604 27706 1660
rect 27706 1604 27710 1660
rect 27646 1600 27710 1604
rect 27726 1660 27790 1664
rect 27726 1604 27730 1660
rect 27730 1604 27786 1660
rect 27786 1604 27790 1660
rect 27726 1600 27790 1604
rect 27806 1660 27870 1664
rect 27806 1604 27810 1660
rect 27810 1604 27866 1660
rect 27866 1604 27870 1660
rect 27806 1600 27870 1604
rect 27886 1660 27950 1664
rect 27886 1604 27890 1660
rect 27890 1604 27946 1660
rect 27946 1604 27950 1660
rect 27886 1600 27950 1604
rect 15884 1396 15948 1460
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 11438 1116 11502 1120
rect 11438 1060 11442 1116
rect 11442 1060 11498 1116
rect 11498 1060 11502 1116
rect 11438 1056 11502 1060
rect 11518 1116 11582 1120
rect 11518 1060 11522 1116
rect 11522 1060 11578 1116
rect 11578 1060 11582 1116
rect 11518 1056 11582 1060
rect 11598 1116 11662 1120
rect 11598 1060 11602 1116
rect 11602 1060 11658 1116
rect 11658 1060 11662 1116
rect 11598 1056 11662 1060
rect 11678 1116 11742 1120
rect 11678 1060 11682 1116
rect 11682 1060 11738 1116
rect 11738 1060 11742 1116
rect 11678 1056 11742 1060
rect 19212 1116 19276 1120
rect 19212 1060 19216 1116
rect 19216 1060 19272 1116
rect 19272 1060 19276 1116
rect 19212 1056 19276 1060
rect 19292 1116 19356 1120
rect 19292 1060 19296 1116
rect 19296 1060 19352 1116
rect 19352 1060 19356 1116
rect 19292 1056 19356 1060
rect 19372 1116 19436 1120
rect 19372 1060 19376 1116
rect 19376 1060 19432 1116
rect 19432 1060 19436 1116
rect 19372 1056 19436 1060
rect 19452 1116 19516 1120
rect 19452 1060 19456 1116
rect 19456 1060 19512 1116
rect 19512 1060 19516 1116
rect 19452 1056 19516 1060
rect 26986 1116 27050 1120
rect 26986 1060 26990 1116
rect 26990 1060 27046 1116
rect 27046 1060 27050 1116
rect 26986 1056 27050 1060
rect 27066 1116 27130 1120
rect 27066 1060 27070 1116
rect 27070 1060 27126 1116
rect 27126 1060 27130 1116
rect 27066 1056 27130 1060
rect 27146 1116 27210 1120
rect 27146 1060 27150 1116
rect 27150 1060 27206 1116
rect 27206 1060 27210 1116
rect 27146 1056 27210 1060
rect 27226 1116 27290 1120
rect 27226 1060 27230 1116
rect 27230 1060 27286 1116
rect 27286 1060 27290 1116
rect 27226 1056 27290 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 12098 572 12162 576
rect 12098 516 12102 572
rect 12102 516 12158 572
rect 12158 516 12162 572
rect 12098 512 12162 516
rect 12178 572 12242 576
rect 12178 516 12182 572
rect 12182 516 12238 572
rect 12238 516 12242 572
rect 12178 512 12242 516
rect 12258 572 12322 576
rect 12258 516 12262 572
rect 12262 516 12318 572
rect 12318 516 12322 572
rect 12258 512 12322 516
rect 12338 572 12402 576
rect 12338 516 12342 572
rect 12342 516 12398 572
rect 12398 516 12402 572
rect 12338 512 12402 516
rect 19872 572 19936 576
rect 19872 516 19876 572
rect 19876 516 19932 572
rect 19932 516 19936 572
rect 19872 512 19936 516
rect 19952 572 20016 576
rect 19952 516 19956 572
rect 19956 516 20012 572
rect 20012 516 20016 572
rect 19952 512 20016 516
rect 20032 572 20096 576
rect 20032 516 20036 572
rect 20036 516 20092 572
rect 20092 516 20096 572
rect 20032 512 20096 516
rect 20112 572 20176 576
rect 20112 516 20116 572
rect 20116 516 20172 572
rect 20172 516 20176 572
rect 20112 512 20176 516
rect 27646 572 27710 576
rect 27646 516 27650 572
rect 27650 516 27706 572
rect 27706 516 27710 572
rect 27646 512 27710 516
rect 27726 572 27790 576
rect 27726 516 27730 572
rect 27730 516 27786 572
rect 27786 516 27790 572
rect 27726 512 27790 516
rect 27806 572 27870 576
rect 27806 516 27810 572
rect 27810 516 27866 572
rect 27866 516 27870 572
rect 27806 512 27870 516
rect 27886 572 27950 576
rect 27886 516 27890 572
rect 27890 516 27946 572
rect 27946 516 27950 572
rect 27886 512 27950 516
<< metal4 >>
rect 3656 21792 3976 21808
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 979 20500 1045 20501
rect 979 20436 980 20500
rect 1044 20436 1045 20500
rect 979 20435 1045 20436
rect 982 8397 1042 20435
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 2635 18324 2701 18325
rect 2635 18260 2636 18324
rect 2700 18260 2701 18324
rect 2635 18259 2701 18260
rect 1163 15332 1229 15333
rect 1163 15268 1164 15332
rect 1228 15268 1229 15332
rect 1163 15267 1229 15268
rect 979 8396 1045 8397
rect 979 8332 980 8396
rect 1044 8332 1045 8396
rect 979 8331 1045 8332
rect 1166 1869 1226 15267
rect 2451 10572 2517 10573
rect 2451 10508 2452 10572
rect 2516 10508 2517 10572
rect 2451 10507 2517 10508
rect 2454 5677 2514 10507
rect 2451 5676 2517 5677
rect 2451 5612 2452 5676
rect 2516 5612 2517 5676
rect 2451 5611 2517 5612
rect 2454 3637 2514 5611
rect 2638 4045 2698 18259
rect 3656 17440 3976 18464
rect 4316 21248 4636 21808
rect 6134 21725 6194 22304
rect 6686 21725 6746 22304
rect 7238 21725 7298 22304
rect 7790 21725 7850 22304
rect 8342 21725 8402 22304
rect 8894 21861 8954 22304
rect 8891 21860 8957 21861
rect 8891 21796 8892 21860
rect 8956 21796 8957 21860
rect 8891 21795 8957 21796
rect 9446 21725 9506 22304
rect 9998 21725 10058 22304
rect 10550 21725 10610 22304
rect 11102 21725 11162 22304
rect 11654 21997 11714 22304
rect 12206 21997 12266 22304
rect 11651 21996 11717 21997
rect 11651 21932 11652 21996
rect 11716 21932 11717 21996
rect 11651 21931 11717 21932
rect 12203 21996 12269 21997
rect 12203 21932 12204 21996
rect 12268 21932 12269 21996
rect 12203 21931 12269 21932
rect 11430 21792 11750 21808
rect 11430 21728 11438 21792
rect 11502 21728 11518 21792
rect 11582 21728 11598 21792
rect 11662 21728 11678 21792
rect 11742 21728 11750 21792
rect 6131 21724 6197 21725
rect 6131 21660 6132 21724
rect 6196 21660 6197 21724
rect 6131 21659 6197 21660
rect 6683 21724 6749 21725
rect 6683 21660 6684 21724
rect 6748 21660 6749 21724
rect 6683 21659 6749 21660
rect 7235 21724 7301 21725
rect 7235 21660 7236 21724
rect 7300 21660 7301 21724
rect 7235 21659 7301 21660
rect 7787 21724 7853 21725
rect 7787 21660 7788 21724
rect 7852 21660 7853 21724
rect 7787 21659 7853 21660
rect 8339 21724 8405 21725
rect 8339 21660 8340 21724
rect 8404 21660 8405 21724
rect 8339 21659 8405 21660
rect 9443 21724 9509 21725
rect 9443 21660 9444 21724
rect 9508 21660 9509 21724
rect 9443 21659 9509 21660
rect 9995 21724 10061 21725
rect 9995 21660 9996 21724
rect 10060 21660 10061 21724
rect 9995 21659 10061 21660
rect 10547 21724 10613 21725
rect 10547 21660 10548 21724
rect 10612 21660 10613 21724
rect 10547 21659 10613 21660
rect 11099 21724 11165 21725
rect 11099 21660 11100 21724
rect 11164 21660 11165 21724
rect 11099 21659 11165 21660
rect 8155 21588 8221 21589
rect 8155 21524 8156 21588
rect 8220 21524 8221 21588
rect 8155 21523 8221 21524
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4107 18188 4173 18189
rect 4107 18124 4108 18188
rect 4172 18124 4173 18188
rect 4107 18123 4173 18124
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3003 12884 3069 12885
rect 3003 12820 3004 12884
rect 3068 12820 3069 12884
rect 3003 12819 3069 12820
rect 3006 11253 3066 12819
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3003 11252 3069 11253
rect 3003 11188 3004 11252
rect 3068 11188 3069 11252
rect 3003 11187 3069 11188
rect 3371 11252 3437 11253
rect 3371 11188 3372 11252
rect 3436 11188 3437 11252
rect 3371 11187 3437 11188
rect 3006 9621 3066 11187
rect 3003 9620 3069 9621
rect 3003 9556 3004 9620
rect 3068 9556 3069 9620
rect 3003 9555 3069 9556
rect 3187 9348 3253 9349
rect 3187 9284 3188 9348
rect 3252 9346 3253 9348
rect 3374 9346 3434 11187
rect 3252 9286 3434 9346
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 4110 10301 4170 18123
rect 4316 17984 4636 19008
rect 5763 18596 5829 18597
rect 5763 18532 5764 18596
rect 5828 18532 5829 18596
rect 5763 18531 5829 18532
rect 6683 18596 6749 18597
rect 6683 18532 6684 18596
rect 6748 18532 6749 18596
rect 6683 18531 6749 18532
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 5211 16692 5277 16693
rect 5211 16628 5212 16692
rect 5276 16628 5277 16692
rect 5211 16627 5277 16628
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 5027 13020 5093 13021
rect 5027 12956 5028 13020
rect 5092 12956 5093 13020
rect 5027 12955 5093 12956
rect 4843 12884 4909 12885
rect 4843 12820 4844 12884
rect 4908 12820 4909 12884
rect 4843 12819 4909 12820
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4846 10981 4906 12819
rect 4843 10980 4909 10981
rect 4843 10916 4844 10980
rect 4908 10916 4909 10980
rect 4843 10915 4909 10916
rect 4843 10844 4909 10845
rect 4843 10780 4844 10844
rect 4908 10780 4909 10844
rect 4843 10779 4909 10780
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4107 10300 4173 10301
rect 4107 10236 4108 10300
rect 4172 10236 4173 10300
rect 4107 10235 4173 10236
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3252 9284 3253 9286
rect 3187 9283 3253 9284
rect 3190 4725 3250 9283
rect 3656 8736 3976 9760
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4107 8940 4173 8941
rect 4107 8876 4108 8940
rect 4172 8876 4173 8940
rect 4107 8875 4173 8876
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 4110 5541 4170 8875
rect 4316 8192 4636 9216
rect 4846 8941 4906 10779
rect 4843 8940 4909 8941
rect 4843 8876 4844 8940
rect 4908 8876 4909 8940
rect 4843 8875 4909 8876
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 5030 7581 5090 12955
rect 5214 10570 5274 16627
rect 5766 15197 5826 18531
rect 6315 17916 6381 17917
rect 6315 17852 6316 17916
rect 6380 17852 6381 17916
rect 6315 17851 6381 17852
rect 5763 15196 5829 15197
rect 5763 15132 5764 15196
rect 5828 15132 5829 15196
rect 5763 15131 5829 15132
rect 5763 13836 5829 13837
rect 5763 13772 5764 13836
rect 5828 13772 5829 13836
rect 5763 13771 5829 13772
rect 5214 10510 5458 10570
rect 5398 10437 5458 10510
rect 5395 10436 5461 10437
rect 5395 10372 5396 10436
rect 5460 10372 5461 10436
rect 5395 10371 5461 10372
rect 5211 8940 5277 8941
rect 5211 8876 5212 8940
rect 5276 8876 5277 8940
rect 5211 8875 5277 8876
rect 5214 8397 5274 8875
rect 5398 8533 5458 10371
rect 5766 9757 5826 13771
rect 6131 13700 6197 13701
rect 6131 13636 6132 13700
rect 6196 13636 6197 13700
rect 6131 13635 6197 13636
rect 6134 10573 6194 13635
rect 6131 10572 6197 10573
rect 6131 10508 6132 10572
rect 6196 10508 6197 10572
rect 6131 10507 6197 10508
rect 6318 10301 6378 17851
rect 6499 12748 6565 12749
rect 6499 12684 6500 12748
rect 6564 12684 6565 12748
rect 6499 12683 6565 12684
rect 6315 10300 6381 10301
rect 6315 10236 6316 10300
rect 6380 10236 6381 10300
rect 6315 10235 6381 10236
rect 5763 9756 5829 9757
rect 5763 9692 5764 9756
rect 5828 9692 5829 9756
rect 5763 9691 5829 9692
rect 6502 9621 6562 12683
rect 6686 11117 6746 18531
rect 7235 16284 7301 16285
rect 7235 16220 7236 16284
rect 7300 16220 7301 16284
rect 7235 16219 7301 16220
rect 7238 14381 7298 16219
rect 7419 16148 7485 16149
rect 7419 16084 7420 16148
rect 7484 16084 7485 16148
rect 7419 16083 7485 16084
rect 7235 14380 7301 14381
rect 7235 14316 7236 14380
rect 7300 14316 7301 14380
rect 7235 14315 7301 14316
rect 7422 12205 7482 16083
rect 7971 15060 8037 15061
rect 7971 14996 7972 15060
rect 8036 14996 8037 15060
rect 7971 14995 8037 14996
rect 7603 14924 7669 14925
rect 7603 14860 7604 14924
rect 7668 14860 7669 14924
rect 7603 14859 7669 14860
rect 7606 14653 7666 14859
rect 7603 14652 7669 14653
rect 7603 14588 7604 14652
rect 7668 14588 7669 14652
rect 7603 14587 7669 14588
rect 7974 13701 8034 14995
rect 7971 13700 8037 13701
rect 7971 13636 7972 13700
rect 8036 13636 8037 13700
rect 7971 13635 8037 13636
rect 8158 13157 8218 21523
rect 11430 20704 11750 21728
rect 11430 20640 11438 20704
rect 11502 20640 11518 20704
rect 11582 20640 11598 20704
rect 11662 20640 11678 20704
rect 11742 20640 11750 20704
rect 11430 19616 11750 20640
rect 11430 19552 11438 19616
rect 11502 19552 11518 19616
rect 11582 19552 11598 19616
rect 11662 19552 11678 19616
rect 11742 19552 11750 19616
rect 11430 18528 11750 19552
rect 11430 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11750 18528
rect 10179 18052 10245 18053
rect 10179 17988 10180 18052
rect 10244 17988 10245 18052
rect 10179 17987 10245 17988
rect 8891 17644 8957 17645
rect 8891 17580 8892 17644
rect 8956 17580 8957 17644
rect 8891 17579 8957 17580
rect 8894 16590 8954 17579
rect 8894 16530 9138 16590
rect 8523 15876 8589 15877
rect 8523 15812 8524 15876
rect 8588 15812 8589 15876
rect 8523 15811 8589 15812
rect 8339 15604 8405 15605
rect 8339 15540 8340 15604
rect 8404 15540 8405 15604
rect 8339 15539 8405 15540
rect 8342 14517 8402 15539
rect 8339 14516 8405 14517
rect 8339 14452 8340 14516
rect 8404 14452 8405 14516
rect 8339 14451 8405 14452
rect 8526 14381 8586 15811
rect 8707 15604 8773 15605
rect 8707 15540 8708 15604
rect 8772 15540 8773 15604
rect 8707 15539 8773 15540
rect 8523 14380 8589 14381
rect 8523 14316 8524 14380
rect 8588 14316 8589 14380
rect 8523 14315 8589 14316
rect 8710 13970 8770 15539
rect 8342 13910 8770 13970
rect 8155 13156 8221 13157
rect 8155 13092 8156 13156
rect 8220 13092 8221 13156
rect 8155 13091 8221 13092
rect 7787 12612 7853 12613
rect 7787 12548 7788 12612
rect 7852 12548 7853 12612
rect 7787 12547 7853 12548
rect 7419 12204 7485 12205
rect 7419 12140 7420 12204
rect 7484 12140 7485 12204
rect 7419 12139 7485 12140
rect 7422 11933 7482 12139
rect 7790 11933 7850 12547
rect 8155 12068 8221 12069
rect 8155 12004 8156 12068
rect 8220 12004 8221 12068
rect 8155 12003 8221 12004
rect 7419 11932 7485 11933
rect 7419 11868 7420 11932
rect 7484 11868 7485 11932
rect 7787 11932 7853 11933
rect 7787 11930 7788 11932
rect 7419 11867 7485 11868
rect 7606 11870 7788 11930
rect 6683 11116 6749 11117
rect 6683 11052 6684 11116
rect 6748 11052 6749 11116
rect 6683 11051 6749 11052
rect 6499 9620 6565 9621
rect 6499 9556 6500 9620
rect 6564 9556 6565 9620
rect 6499 9555 6565 9556
rect 7606 8805 7666 11870
rect 7787 11868 7788 11870
rect 7852 11868 7853 11932
rect 7787 11867 7853 11868
rect 7787 10436 7853 10437
rect 7787 10372 7788 10436
rect 7852 10372 7853 10436
rect 7787 10371 7853 10372
rect 7603 8804 7669 8805
rect 7603 8740 7604 8804
rect 7668 8740 7669 8804
rect 7603 8739 7669 8740
rect 5395 8532 5461 8533
rect 5395 8468 5396 8532
rect 5460 8468 5461 8532
rect 5395 8467 5461 8468
rect 5211 8396 5277 8397
rect 5211 8332 5212 8396
rect 5276 8332 5277 8396
rect 5211 8331 5277 8332
rect 5027 7580 5093 7581
rect 5027 7516 5028 7580
rect 5092 7516 5093 7580
rect 5027 7515 5093 7516
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 5398 6357 5458 8467
rect 5395 6356 5461 6357
rect 5395 6292 5396 6356
rect 5460 6292 5461 6356
rect 5395 6291 5461 6292
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4107 5540 4173 5541
rect 4107 5476 4108 5540
rect 4172 5476 4173 5540
rect 4107 5475 4173 5476
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3187 4724 3253 4725
rect 3187 4660 3188 4724
rect 3252 4660 3253 4724
rect 3187 4659 3253 4660
rect 3190 4181 3250 4659
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3187 4180 3253 4181
rect 3187 4116 3188 4180
rect 3252 4116 3253 4180
rect 3187 4115 3253 4116
rect 2635 4044 2701 4045
rect 2635 3980 2636 4044
rect 2700 3980 2701 4044
rect 2635 3979 2701 3980
rect 2451 3636 2517 3637
rect 2451 3572 2452 3636
rect 2516 3572 2517 3636
rect 2451 3571 2517 3572
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 1163 1868 1229 1869
rect 1163 1804 1164 1868
rect 1228 1804 1229 1868
rect 1163 1803 1229 1804
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 4928 4636 5952
rect 7790 5541 7850 10371
rect 7971 6084 8037 6085
rect 7971 6020 7972 6084
rect 8036 6020 8037 6084
rect 7971 6019 8037 6020
rect 7787 5540 7853 5541
rect 7787 5476 7788 5540
rect 7852 5476 7853 5540
rect 7787 5475 7853 5476
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 7974 3093 8034 6019
rect 8158 5813 8218 12003
rect 8342 8261 8402 13910
rect 8707 13836 8773 13837
rect 8707 13772 8708 13836
rect 8772 13772 8773 13836
rect 8707 13771 8773 13772
rect 8523 11524 8589 11525
rect 8523 11460 8524 11524
rect 8588 11460 8589 11524
rect 8523 11459 8589 11460
rect 8526 8533 8586 11459
rect 8523 8532 8589 8533
rect 8523 8468 8524 8532
rect 8588 8468 8589 8532
rect 8523 8467 8589 8468
rect 8339 8260 8405 8261
rect 8339 8196 8340 8260
rect 8404 8196 8405 8260
rect 8339 8195 8405 8196
rect 8710 7581 8770 13771
rect 8891 12204 8957 12205
rect 8891 12140 8892 12204
rect 8956 12140 8957 12204
rect 8891 12139 8957 12140
rect 8894 8805 8954 12139
rect 9078 12069 9138 16530
rect 9259 15740 9325 15741
rect 9259 15676 9260 15740
rect 9324 15676 9325 15740
rect 9259 15675 9325 15676
rect 9075 12068 9141 12069
rect 9075 12004 9076 12068
rect 9140 12004 9141 12068
rect 9075 12003 9141 12004
rect 9075 11116 9141 11117
rect 9075 11052 9076 11116
rect 9140 11052 9141 11116
rect 9075 11051 9141 11052
rect 8891 8804 8957 8805
rect 8891 8740 8892 8804
rect 8956 8740 8957 8804
rect 8891 8739 8957 8740
rect 9078 8310 9138 11051
rect 9262 9893 9322 15675
rect 9811 14788 9877 14789
rect 9811 14724 9812 14788
rect 9876 14724 9877 14788
rect 9811 14723 9877 14724
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 9446 10709 9506 13499
rect 9627 13156 9693 13157
rect 9627 13092 9628 13156
rect 9692 13092 9693 13156
rect 9627 13091 9693 13092
rect 9630 10845 9690 13091
rect 9627 10844 9693 10845
rect 9627 10780 9628 10844
rect 9692 10780 9693 10844
rect 9627 10779 9693 10780
rect 9443 10708 9509 10709
rect 9443 10644 9444 10708
rect 9508 10644 9509 10708
rect 9443 10643 9509 10644
rect 9814 9893 9874 14723
rect 9995 12204 10061 12205
rect 9995 12140 9996 12204
rect 10060 12140 10061 12204
rect 9995 12139 10061 12140
rect 9998 10573 10058 12139
rect 9995 10572 10061 10573
rect 9995 10508 9996 10572
rect 10060 10508 10061 10572
rect 9995 10507 10061 10508
rect 9995 10300 10061 10301
rect 9995 10236 9996 10300
rect 10060 10236 10061 10300
rect 9995 10235 10061 10236
rect 9259 9892 9325 9893
rect 9259 9828 9260 9892
rect 9324 9828 9325 9892
rect 9259 9827 9325 9828
rect 9811 9892 9877 9893
rect 9811 9828 9812 9892
rect 9876 9828 9877 9892
rect 9811 9827 9877 9828
rect 9262 9077 9322 9827
rect 9998 9690 10058 10235
rect 9630 9630 10058 9690
rect 9259 9076 9325 9077
rect 9259 9012 9260 9076
rect 9324 9012 9325 9076
rect 9259 9011 9325 9012
rect 9078 8250 9506 8310
rect 9446 7581 9506 8250
rect 8707 7580 8773 7581
rect 8707 7516 8708 7580
rect 8772 7516 8773 7580
rect 8707 7515 8773 7516
rect 9443 7580 9509 7581
rect 9443 7516 9444 7580
rect 9508 7516 9509 7580
rect 9443 7515 9509 7516
rect 9630 7037 9690 9630
rect 9627 7036 9693 7037
rect 9627 6972 9628 7036
rect 9692 6972 9693 7036
rect 9627 6971 9693 6972
rect 8155 5812 8221 5813
rect 8155 5748 8156 5812
rect 8220 5748 8221 5812
rect 8155 5747 8221 5748
rect 8155 5676 8221 5677
rect 8155 5612 8156 5676
rect 8220 5612 8221 5676
rect 8155 5611 8221 5612
rect 8158 3501 8218 5611
rect 10182 4861 10242 17987
rect 11099 17916 11165 17917
rect 11099 17852 11100 17916
rect 11164 17852 11165 17916
rect 11099 17851 11165 17852
rect 10547 17372 10613 17373
rect 10547 17308 10548 17372
rect 10612 17308 10613 17372
rect 10547 17307 10613 17308
rect 10550 16285 10610 17307
rect 11102 17101 11162 17851
rect 11430 17440 11750 18464
rect 12090 21248 12410 21808
rect 12758 21725 12818 22304
rect 13310 21725 13370 22304
rect 13862 21725 13922 22304
rect 12755 21724 12821 21725
rect 12755 21660 12756 21724
rect 12820 21660 12821 21724
rect 12755 21659 12821 21660
rect 13307 21724 13373 21725
rect 13307 21660 13308 21724
rect 13372 21660 13373 21724
rect 13307 21659 13373 21660
rect 13859 21724 13925 21725
rect 13859 21660 13860 21724
rect 13924 21660 13925 21724
rect 13859 21659 13925 21660
rect 12090 21184 12098 21248
rect 12162 21184 12178 21248
rect 12242 21184 12258 21248
rect 12322 21184 12338 21248
rect 12402 21184 12410 21248
rect 12090 20160 12410 21184
rect 14414 20637 14474 22304
rect 14411 20636 14477 20637
rect 14411 20572 14412 20636
rect 14476 20572 14477 20636
rect 14411 20571 14477 20572
rect 12090 20096 12098 20160
rect 12162 20096 12178 20160
rect 12242 20096 12258 20160
rect 12322 20096 12338 20160
rect 12402 20096 12410 20160
rect 12090 19072 12410 20096
rect 14966 19957 15026 22304
rect 15518 21045 15578 22304
rect 15515 21044 15581 21045
rect 15515 20980 15516 21044
rect 15580 20980 15581 21044
rect 15515 20979 15581 20980
rect 16070 20637 16130 22304
rect 16622 21725 16682 22304
rect 16619 21724 16685 21725
rect 16619 21660 16620 21724
rect 16684 21660 16685 21724
rect 16619 21659 16685 21660
rect 17174 21181 17234 22304
rect 17171 21180 17237 21181
rect 17171 21116 17172 21180
rect 17236 21116 17237 21180
rect 17171 21115 17237 21116
rect 17726 20637 17786 22304
rect 18278 21453 18338 22304
rect 18830 21589 18890 22304
rect 19382 22104 19442 22304
rect 19934 22104 19994 22304
rect 20299 22132 20365 22133
rect 20299 22068 20300 22132
rect 20364 22068 20365 22132
rect 20486 22104 20546 22304
rect 21038 22104 21098 22304
rect 21590 22104 21650 22304
rect 22142 22104 22202 22304
rect 22694 22104 22754 22304
rect 23246 22104 23306 22304
rect 23798 22104 23858 22304
rect 24350 22104 24410 22304
rect 24902 22104 24962 22304
rect 25454 22104 25514 22304
rect 26006 22104 26066 22304
rect 26558 22104 26618 22304
rect 27110 22104 27170 22304
rect 27662 22104 27722 22304
rect 20299 22067 20365 22068
rect 20302 21994 20362 22067
rect 24347 21996 24413 21997
rect 20302 21934 20546 21994
rect 19204 21792 19524 21808
rect 19204 21728 19212 21792
rect 19276 21728 19292 21792
rect 19356 21728 19372 21792
rect 19436 21728 19452 21792
rect 19516 21728 19524 21792
rect 18827 21588 18893 21589
rect 18827 21524 18828 21588
rect 18892 21524 18893 21588
rect 18827 21523 18893 21524
rect 18275 21452 18341 21453
rect 18275 21388 18276 21452
rect 18340 21388 18341 21452
rect 18275 21387 18341 21388
rect 19204 20704 19524 21728
rect 19204 20640 19212 20704
rect 19276 20640 19292 20704
rect 19356 20640 19372 20704
rect 19436 20640 19452 20704
rect 19516 20640 19524 20704
rect 16067 20636 16133 20637
rect 16067 20572 16068 20636
rect 16132 20572 16133 20636
rect 16067 20571 16133 20572
rect 17723 20636 17789 20637
rect 17723 20572 17724 20636
rect 17788 20572 17789 20636
rect 17723 20571 17789 20572
rect 14963 19956 15029 19957
rect 14963 19892 14964 19956
rect 15028 19892 15029 19956
rect 14963 19891 15029 19892
rect 19204 19616 19524 20640
rect 19204 19552 19212 19616
rect 19276 19552 19292 19616
rect 19356 19552 19372 19616
rect 19436 19552 19452 19616
rect 19516 19552 19524 19616
rect 16435 19412 16501 19413
rect 16435 19348 16436 19412
rect 16500 19348 16501 19412
rect 16435 19347 16501 19348
rect 14043 19276 14109 19277
rect 14043 19212 14044 19276
rect 14108 19212 14109 19276
rect 14043 19211 14109 19212
rect 12090 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12410 19072
rect 11835 18460 11901 18461
rect 11835 18396 11836 18460
rect 11900 18396 11901 18460
rect 11835 18395 11901 18396
rect 11838 17917 11898 18395
rect 12090 17984 12410 19008
rect 12090 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12410 17984
rect 11835 17916 11901 17917
rect 11835 17852 11836 17916
rect 11900 17852 11901 17916
rect 11835 17851 11901 17852
rect 11835 17508 11901 17509
rect 11835 17444 11836 17508
rect 11900 17444 11901 17508
rect 11835 17443 11901 17444
rect 11430 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11750 17440
rect 11099 17100 11165 17101
rect 11099 17036 11100 17100
rect 11164 17036 11165 17100
rect 11099 17035 11165 17036
rect 10915 16828 10981 16829
rect 10915 16764 10916 16828
rect 10980 16764 10981 16828
rect 10915 16763 10981 16764
rect 10547 16284 10613 16285
rect 10547 16220 10548 16284
rect 10612 16220 10613 16284
rect 10547 16219 10613 16220
rect 10731 14244 10797 14245
rect 10731 14180 10732 14244
rect 10796 14180 10797 14244
rect 10731 14179 10797 14180
rect 10734 13565 10794 14179
rect 10918 13701 10978 16763
rect 11430 16352 11750 17376
rect 11838 16829 11898 17443
rect 12090 16896 12410 17920
rect 14046 17645 14106 19211
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 13859 17644 13925 17645
rect 13859 17580 13860 17644
rect 13924 17580 13925 17644
rect 13859 17579 13925 17580
rect 14043 17644 14109 17645
rect 14043 17580 14044 17644
rect 14108 17580 14109 17644
rect 14043 17579 14109 17580
rect 12939 17508 13005 17509
rect 12939 17444 12940 17508
rect 13004 17444 13005 17508
rect 12939 17443 13005 17444
rect 12755 16964 12821 16965
rect 12755 16900 12756 16964
rect 12820 16900 12821 16964
rect 12755 16899 12821 16900
rect 12090 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12410 16896
rect 11835 16828 11901 16829
rect 11835 16764 11836 16828
rect 11900 16764 11901 16828
rect 11835 16763 11901 16764
rect 11430 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11750 16352
rect 11099 15332 11165 15333
rect 11099 15268 11100 15332
rect 11164 15268 11165 15332
rect 11099 15267 11165 15268
rect 10915 13700 10981 13701
rect 10915 13636 10916 13700
rect 10980 13636 10981 13700
rect 10915 13635 10981 13636
rect 10731 13564 10797 13565
rect 10731 13500 10732 13564
rect 10796 13500 10797 13564
rect 10731 13499 10797 13500
rect 10547 12068 10613 12069
rect 10547 12004 10548 12068
rect 10612 12004 10613 12068
rect 10547 12003 10613 12004
rect 10550 11253 10610 12003
rect 10547 11252 10613 11253
rect 10547 11188 10548 11252
rect 10612 11188 10613 11252
rect 10547 11187 10613 11188
rect 10547 10980 10613 10981
rect 10547 10916 10548 10980
rect 10612 10916 10613 10980
rect 10547 10915 10613 10916
rect 10363 9892 10429 9893
rect 10363 9828 10364 9892
rect 10428 9828 10429 9892
rect 10363 9827 10429 9828
rect 10366 6221 10426 9827
rect 10363 6220 10429 6221
rect 10363 6156 10364 6220
rect 10428 6156 10429 6220
rect 10363 6155 10429 6156
rect 10550 5949 10610 10915
rect 10734 6629 10794 13499
rect 11102 12474 11162 15267
rect 11430 15264 11750 16288
rect 12090 15808 12410 16832
rect 12571 15876 12637 15877
rect 12571 15812 12572 15876
rect 12636 15812 12637 15876
rect 12571 15811 12637 15812
rect 12090 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12410 15808
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11430 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11750 15264
rect 11283 15196 11349 15197
rect 11283 15132 11284 15196
rect 11348 15132 11349 15196
rect 11283 15131 11349 15132
rect 11286 12613 11346 15131
rect 11430 14176 11750 15200
rect 11430 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11750 14176
rect 11430 13088 11750 14112
rect 11838 13701 11898 15267
rect 12090 14720 12410 15744
rect 12090 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12410 14720
rect 11835 13700 11901 13701
rect 11835 13636 11836 13700
rect 11900 13636 11901 13700
rect 11835 13635 11901 13636
rect 11430 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11750 13088
rect 11283 12612 11349 12613
rect 11283 12548 11284 12612
rect 11348 12548 11349 12612
rect 11283 12547 11349 12548
rect 11102 12414 11346 12474
rect 10915 12068 10981 12069
rect 10915 12004 10916 12068
rect 10980 12004 10981 12068
rect 10915 12003 10981 12004
rect 10731 6628 10797 6629
rect 10731 6564 10732 6628
rect 10796 6564 10797 6628
rect 10731 6563 10797 6564
rect 10547 5948 10613 5949
rect 10547 5884 10548 5948
rect 10612 5884 10613 5948
rect 10547 5883 10613 5884
rect 10179 4860 10245 4861
rect 10179 4796 10180 4860
rect 10244 4796 10245 4860
rect 10179 4795 10245 4796
rect 10918 4589 10978 12003
rect 11099 11252 11165 11253
rect 11099 11188 11100 11252
rect 11164 11188 11165 11252
rect 11099 11187 11165 11188
rect 11102 9893 11162 11187
rect 11286 10301 11346 12414
rect 11430 12000 11750 13024
rect 11430 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11750 12000
rect 11430 10912 11750 11936
rect 11430 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11750 10912
rect 11283 10300 11349 10301
rect 11283 10236 11284 10300
rect 11348 10236 11349 10300
rect 11283 10235 11349 10236
rect 11099 9892 11165 9893
rect 11099 9828 11100 9892
rect 11164 9828 11165 9892
rect 11099 9827 11165 9828
rect 11430 9824 11750 10848
rect 11430 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11750 9824
rect 11099 9756 11165 9757
rect 11099 9692 11100 9756
rect 11164 9692 11165 9756
rect 11099 9691 11165 9692
rect 11102 6357 11162 9691
rect 11283 9076 11349 9077
rect 11283 9012 11284 9076
rect 11348 9012 11349 9076
rect 11283 9011 11349 9012
rect 11099 6356 11165 6357
rect 11099 6292 11100 6356
rect 11164 6292 11165 6356
rect 11099 6291 11165 6292
rect 10915 4588 10981 4589
rect 10915 4524 10916 4588
rect 10980 4524 10981 4588
rect 10915 4523 10981 4524
rect 11286 3909 11346 9011
rect 11430 8736 11750 9760
rect 11838 9077 11898 13635
rect 12090 13632 12410 14656
rect 12090 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12410 13632
rect 12090 12544 12410 13568
rect 12090 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12410 12544
rect 12090 11456 12410 12480
rect 12090 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12410 11456
rect 12090 10368 12410 11392
rect 12574 11253 12634 15811
rect 12571 11252 12637 11253
rect 12571 11188 12572 11252
rect 12636 11188 12637 11252
rect 12571 11187 12637 11188
rect 12090 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12410 10368
rect 12090 9280 12410 10304
rect 12571 9892 12637 9893
rect 12571 9828 12572 9892
rect 12636 9828 12637 9892
rect 12571 9827 12637 9828
rect 12574 9349 12634 9827
rect 12571 9348 12637 9349
rect 12571 9284 12572 9348
rect 12636 9284 12637 9348
rect 12571 9283 12637 9284
rect 12090 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12410 9280
rect 11835 9076 11901 9077
rect 11835 9012 11836 9076
rect 11900 9012 11901 9076
rect 11835 9011 11901 9012
rect 11430 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11750 8736
rect 11430 7648 11750 8672
rect 11430 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11750 7648
rect 11430 6560 11750 7584
rect 11430 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11750 6560
rect 11430 5472 11750 6496
rect 11430 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11750 5472
rect 11430 4384 11750 5408
rect 11430 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11750 4384
rect 11283 3908 11349 3909
rect 11283 3844 11284 3908
rect 11348 3844 11349 3908
rect 11283 3843 11349 3844
rect 8155 3500 8221 3501
rect 8155 3436 8156 3500
rect 8220 3436 8221 3500
rect 8155 3435 8221 3436
rect 11430 3296 11750 4320
rect 11430 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11750 3296
rect 7971 3092 8037 3093
rect 7971 3028 7972 3092
rect 8036 3028 8037 3092
rect 7971 3027 8037 3028
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 11430 2208 11750 3232
rect 11430 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11750 2208
rect 11430 1120 11750 2144
rect 11430 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11750 1120
rect 11430 496 11750 1056
rect 12090 8192 12410 9216
rect 12090 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12410 8192
rect 12090 7104 12410 8128
rect 12090 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12410 7104
rect 12090 6016 12410 7040
rect 12574 6629 12634 9283
rect 12571 6628 12637 6629
rect 12571 6564 12572 6628
rect 12636 6564 12637 6628
rect 12571 6563 12637 6564
rect 12090 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12410 6016
rect 12090 4928 12410 5952
rect 12090 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12410 4928
rect 12090 3840 12410 4864
rect 12090 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12410 3840
rect 12090 2752 12410 3776
rect 12758 3773 12818 16899
rect 12942 13701 13002 17443
rect 13123 15876 13189 15877
rect 13123 15812 13124 15876
rect 13188 15812 13189 15876
rect 13123 15811 13189 15812
rect 12939 13700 13005 13701
rect 12939 13636 12940 13700
rect 13004 13636 13005 13700
rect 12939 13635 13005 13636
rect 12939 13564 13005 13565
rect 12939 13500 12940 13564
rect 13004 13500 13005 13564
rect 12939 13499 13005 13500
rect 12942 12477 13002 13499
rect 12939 12476 13005 12477
rect 12939 12412 12940 12476
rect 13004 12412 13005 12476
rect 12939 12411 13005 12412
rect 12939 11116 13005 11117
rect 12939 11052 12940 11116
rect 13004 11052 13005 11116
rect 12939 11051 13005 11052
rect 12942 6493 13002 11051
rect 13126 10981 13186 15811
rect 13675 15332 13741 15333
rect 13675 15268 13676 15332
rect 13740 15268 13741 15332
rect 13675 15267 13741 15268
rect 13491 12748 13557 12749
rect 13491 12684 13492 12748
rect 13556 12684 13557 12748
rect 13491 12683 13557 12684
rect 13123 10980 13189 10981
rect 13123 10916 13124 10980
rect 13188 10916 13189 10980
rect 13123 10915 13189 10916
rect 13494 9621 13554 12683
rect 13491 9620 13557 9621
rect 13491 9556 13492 9620
rect 13556 9556 13557 9620
rect 13491 9555 13557 9556
rect 13123 9484 13189 9485
rect 13123 9420 13124 9484
rect 13188 9420 13189 9484
rect 13123 9419 13189 9420
rect 12939 6492 13005 6493
rect 12939 6428 12940 6492
rect 13004 6428 13005 6492
rect 12939 6427 13005 6428
rect 12755 3772 12821 3773
rect 12755 3708 12756 3772
rect 12820 3708 12821 3772
rect 12755 3707 12821 3708
rect 12090 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12410 2752
rect 12090 1664 12410 2688
rect 13126 2413 13186 9419
rect 13307 9076 13373 9077
rect 13307 9012 13308 9076
rect 13372 9012 13373 9076
rect 13307 9011 13373 9012
rect 13123 2412 13189 2413
rect 13123 2348 13124 2412
rect 13188 2348 13189 2412
rect 13123 2347 13189 2348
rect 13310 2005 13370 9011
rect 13678 8669 13738 15267
rect 13862 13565 13922 17579
rect 14411 17508 14477 17509
rect 14411 17444 14412 17508
rect 14476 17444 14477 17508
rect 14411 17443 14477 17444
rect 14043 17236 14109 17237
rect 14043 17172 14044 17236
rect 14108 17172 14109 17236
rect 14043 17171 14109 17172
rect 14046 14653 14106 17171
rect 14043 14652 14109 14653
rect 14043 14588 14044 14652
rect 14108 14588 14109 14652
rect 14043 14587 14109 14588
rect 13859 13564 13925 13565
rect 13859 13500 13860 13564
rect 13924 13500 13925 13564
rect 13859 13499 13925 13500
rect 14046 11525 14106 14587
rect 14043 11524 14109 11525
rect 14043 11460 14044 11524
rect 14108 11460 14109 11524
rect 14043 11459 14109 11460
rect 14043 10980 14109 10981
rect 14043 10916 14044 10980
rect 14108 10916 14109 10980
rect 14043 10915 14109 10916
rect 14227 10980 14293 10981
rect 14227 10916 14228 10980
rect 14292 10916 14293 10980
rect 14227 10915 14293 10916
rect 13859 9892 13925 9893
rect 13859 9828 13860 9892
rect 13924 9828 13925 9892
rect 13859 9827 13925 9828
rect 13862 9349 13922 9827
rect 13859 9348 13925 9349
rect 13859 9284 13860 9348
rect 13924 9284 13925 9348
rect 13859 9283 13925 9284
rect 13859 9076 13925 9077
rect 13859 9012 13860 9076
rect 13924 9012 13925 9076
rect 13859 9011 13925 9012
rect 13675 8668 13741 8669
rect 13675 8604 13676 8668
rect 13740 8604 13741 8668
rect 13675 8603 13741 8604
rect 13862 2957 13922 9011
rect 14046 8941 14106 10915
rect 14230 10165 14290 10915
rect 14227 10164 14293 10165
rect 14227 10100 14228 10164
rect 14292 10100 14293 10164
rect 14227 10099 14293 10100
rect 14043 8940 14109 8941
rect 14043 8876 14044 8940
rect 14108 8876 14109 8940
rect 14043 8875 14109 8876
rect 14414 7578 14474 17443
rect 15147 16964 15213 16965
rect 15147 16900 15148 16964
rect 15212 16900 15213 16964
rect 15147 16899 15213 16900
rect 14595 16556 14661 16557
rect 14595 16492 14596 16556
rect 14660 16492 14661 16556
rect 14595 16491 14661 16492
rect 14598 11253 14658 16491
rect 15150 15210 15210 16899
rect 15331 16692 15397 16693
rect 15331 16628 15332 16692
rect 15396 16628 15397 16692
rect 15331 16627 15397 16628
rect 14782 15150 15210 15210
rect 14782 12610 14842 15150
rect 14963 14380 15029 14381
rect 14963 14316 14964 14380
rect 15028 14316 15029 14380
rect 14963 14315 15029 14316
rect 14966 12749 15026 14315
rect 14963 12748 15029 12749
rect 14963 12684 14964 12748
rect 15028 12684 15029 12748
rect 14963 12683 15029 12684
rect 14782 12550 15210 12610
rect 14963 12340 15029 12341
rect 14963 12338 14964 12340
rect 14782 12278 14964 12338
rect 14595 11252 14661 11253
rect 14595 11188 14596 11252
rect 14660 11188 14661 11252
rect 14595 11187 14661 11188
rect 14782 10570 14842 12278
rect 14963 12276 14964 12278
rect 15028 12276 15029 12340
rect 14963 12275 15029 12276
rect 14963 12204 15029 12205
rect 14963 12140 14964 12204
rect 15028 12140 15029 12204
rect 14963 12139 15029 12140
rect 14598 10510 14842 10570
rect 14598 9893 14658 10510
rect 14779 10436 14845 10437
rect 14779 10372 14780 10436
rect 14844 10372 14845 10436
rect 14779 10371 14845 10372
rect 14595 9892 14661 9893
rect 14595 9828 14596 9892
rect 14660 9828 14661 9892
rect 14595 9827 14661 9828
rect 14782 8666 14842 10371
rect 14598 8606 14842 8666
rect 14966 8666 15026 12139
rect 15150 10165 15210 12550
rect 15147 10164 15213 10165
rect 15147 10100 15148 10164
rect 15212 10100 15213 10164
rect 15147 10099 15213 10100
rect 15334 9074 15394 16627
rect 15518 11797 15578 17987
rect 15883 16692 15949 16693
rect 15883 16628 15884 16692
rect 15948 16628 15949 16692
rect 15883 16627 15949 16628
rect 16251 16692 16317 16693
rect 16251 16628 16252 16692
rect 16316 16628 16317 16692
rect 16251 16627 16317 16628
rect 15699 15332 15765 15333
rect 15699 15268 15700 15332
rect 15764 15268 15765 15332
rect 15699 15267 15765 15268
rect 15515 11796 15581 11797
rect 15515 11732 15516 11796
rect 15580 11732 15581 11796
rect 15515 11731 15581 11732
rect 15515 11388 15581 11389
rect 15515 11324 15516 11388
rect 15580 11324 15581 11388
rect 15515 11323 15581 11324
rect 15518 9893 15578 11323
rect 15515 9892 15581 9893
rect 15515 9828 15516 9892
rect 15580 9828 15581 9892
rect 15515 9827 15581 9828
rect 15334 9014 15578 9074
rect 15331 8668 15397 8669
rect 15331 8666 15332 8668
rect 14966 8606 15332 8666
rect 14598 8261 14658 8606
rect 15331 8604 15332 8606
rect 15396 8604 15397 8668
rect 15331 8603 15397 8604
rect 14595 8260 14661 8261
rect 14595 8196 14596 8260
rect 14660 8196 14661 8260
rect 14595 8195 14661 8196
rect 14963 8260 15029 8261
rect 14963 8196 14964 8260
rect 15028 8196 15029 8260
rect 14963 8195 15029 8196
rect 14598 7850 14658 8195
rect 14598 7790 14842 7850
rect 14414 7518 14658 7578
rect 14598 6930 14658 7518
rect 14782 7309 14842 7790
rect 14779 7308 14845 7309
rect 14779 7244 14780 7308
rect 14844 7244 14845 7308
rect 14779 7243 14845 7244
rect 14414 6870 14658 6930
rect 14414 3637 14474 6870
rect 14966 5550 15026 8195
rect 15518 5949 15578 9014
rect 15515 5948 15581 5949
rect 15515 5884 15516 5948
rect 15580 5884 15581 5948
rect 15515 5883 15581 5884
rect 14966 5541 15210 5550
rect 14966 5540 15213 5541
rect 14966 5490 15148 5540
rect 15147 5476 15148 5490
rect 15212 5476 15213 5540
rect 15147 5475 15213 5476
rect 15150 4725 15210 5475
rect 15702 4861 15762 15267
rect 15886 12749 15946 16627
rect 15883 12748 15949 12749
rect 15883 12684 15884 12748
rect 15948 12684 15949 12748
rect 15883 12683 15949 12684
rect 16067 12612 16133 12613
rect 16067 12548 16068 12612
rect 16132 12548 16133 12612
rect 16067 12547 16133 12548
rect 15883 10436 15949 10437
rect 15883 10372 15884 10436
rect 15948 10372 15949 10436
rect 15883 10371 15949 10372
rect 15699 4860 15765 4861
rect 15699 4796 15700 4860
rect 15764 4796 15765 4860
rect 15699 4795 15765 4796
rect 15147 4724 15213 4725
rect 15147 4660 15148 4724
rect 15212 4660 15213 4724
rect 15147 4659 15213 4660
rect 14411 3636 14477 3637
rect 14411 3572 14412 3636
rect 14476 3572 14477 3636
rect 14411 3571 14477 3572
rect 13859 2956 13925 2957
rect 13859 2892 13860 2956
rect 13924 2892 13925 2956
rect 13859 2891 13925 2892
rect 13307 2004 13373 2005
rect 13307 1940 13308 2004
rect 13372 1940 13373 2004
rect 13307 1939 13373 1940
rect 12090 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12410 1664
rect 12090 576 12410 1600
rect 15886 1461 15946 10371
rect 16070 3909 16130 12547
rect 16254 9077 16314 16627
rect 16438 15197 16498 19347
rect 19204 18528 19524 19552
rect 19204 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19524 18528
rect 19204 17440 19524 18464
rect 19204 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19524 17440
rect 18643 16828 18709 16829
rect 18643 16764 18644 16828
rect 18708 16764 18709 16828
rect 18643 16763 18709 16764
rect 16803 16692 16869 16693
rect 16803 16628 16804 16692
rect 16868 16628 16869 16692
rect 16803 16627 16869 16628
rect 16435 15196 16501 15197
rect 16435 15132 16436 15196
rect 16500 15132 16501 15196
rect 16435 15131 16501 15132
rect 16619 12884 16685 12885
rect 16619 12820 16620 12884
rect 16684 12820 16685 12884
rect 16619 12819 16685 12820
rect 16435 11388 16501 11389
rect 16435 11324 16436 11388
rect 16500 11324 16501 11388
rect 16435 11323 16501 11324
rect 16251 9076 16317 9077
rect 16251 9012 16252 9076
rect 16316 9012 16317 9076
rect 16251 9011 16317 9012
rect 16438 7853 16498 11323
rect 16622 9893 16682 12819
rect 16619 9892 16685 9893
rect 16619 9828 16620 9892
rect 16684 9828 16685 9892
rect 16619 9827 16685 9828
rect 16806 9485 16866 16627
rect 18091 14652 18157 14653
rect 18091 14588 18092 14652
rect 18156 14588 18157 14652
rect 18091 14587 18157 14588
rect 17355 13156 17421 13157
rect 17355 13092 17356 13156
rect 17420 13092 17421 13156
rect 17355 13091 17421 13092
rect 16987 9892 17053 9893
rect 16987 9828 16988 9892
rect 17052 9828 17053 9892
rect 16987 9827 17053 9828
rect 16803 9484 16869 9485
rect 16803 9420 16804 9484
rect 16868 9420 16869 9484
rect 16803 9419 16869 9420
rect 16619 9348 16685 9349
rect 16619 9284 16620 9348
rect 16684 9284 16685 9348
rect 16619 9283 16685 9284
rect 16435 7852 16501 7853
rect 16435 7788 16436 7852
rect 16500 7788 16501 7852
rect 16435 7787 16501 7788
rect 16622 6357 16682 9283
rect 16990 7037 17050 9827
rect 17358 8125 17418 13091
rect 17907 12204 17973 12205
rect 17907 12140 17908 12204
rect 17972 12140 17973 12204
rect 17907 12139 17973 12140
rect 17539 10300 17605 10301
rect 17539 10236 17540 10300
rect 17604 10236 17605 10300
rect 17539 10235 17605 10236
rect 17542 8533 17602 10235
rect 17910 9349 17970 12139
rect 17907 9348 17973 9349
rect 17907 9284 17908 9348
rect 17972 9284 17973 9348
rect 17907 9283 17973 9284
rect 17539 8532 17605 8533
rect 17539 8468 17540 8532
rect 17604 8468 17605 8532
rect 17539 8467 17605 8468
rect 18094 8125 18154 14587
rect 18275 12884 18341 12885
rect 18275 12820 18276 12884
rect 18340 12820 18341 12884
rect 18275 12819 18341 12820
rect 18278 9893 18338 12819
rect 18459 12748 18525 12749
rect 18459 12684 18460 12748
rect 18524 12684 18525 12748
rect 18459 12683 18525 12684
rect 18462 10709 18522 12683
rect 18459 10708 18525 10709
rect 18459 10644 18460 10708
rect 18524 10644 18525 10708
rect 18459 10643 18525 10644
rect 18275 9892 18341 9893
rect 18275 9828 18276 9892
rect 18340 9828 18341 9892
rect 18275 9827 18341 9828
rect 18646 9621 18706 16763
rect 19204 16352 19524 17376
rect 19204 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19524 16352
rect 19204 15264 19524 16288
rect 19204 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19524 15264
rect 18827 14652 18893 14653
rect 18827 14588 18828 14652
rect 18892 14588 18893 14652
rect 18827 14587 18893 14588
rect 18830 11797 18890 14587
rect 19204 14176 19524 15200
rect 19204 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19524 14176
rect 19011 13292 19077 13293
rect 19011 13228 19012 13292
rect 19076 13228 19077 13292
rect 19011 13227 19077 13228
rect 18827 11796 18893 11797
rect 18827 11732 18828 11796
rect 18892 11732 18893 11796
rect 18827 11731 18893 11732
rect 18827 10300 18893 10301
rect 18827 10236 18828 10300
rect 18892 10236 18893 10300
rect 18827 10235 18893 10236
rect 18643 9620 18709 9621
rect 18643 9618 18644 9620
rect 18278 9558 18644 9618
rect 17355 8124 17421 8125
rect 17355 8060 17356 8124
rect 17420 8060 17421 8124
rect 17355 8059 17421 8060
rect 18091 8124 18157 8125
rect 18091 8060 18092 8124
rect 18156 8060 18157 8124
rect 18091 8059 18157 8060
rect 18278 7581 18338 9558
rect 18643 9556 18644 9558
rect 18708 9556 18709 9620
rect 18643 9555 18709 9556
rect 18646 9464 18706 9555
rect 18459 9348 18525 9349
rect 18459 9284 18460 9348
rect 18524 9284 18525 9348
rect 18459 9283 18525 9284
rect 18462 8125 18522 9283
rect 18643 8804 18709 8805
rect 18643 8740 18644 8804
rect 18708 8740 18709 8804
rect 18643 8739 18709 8740
rect 18459 8124 18525 8125
rect 18459 8060 18460 8124
rect 18524 8060 18525 8124
rect 18459 8059 18525 8060
rect 18275 7580 18341 7581
rect 18275 7516 18276 7580
rect 18340 7516 18341 7580
rect 18275 7515 18341 7516
rect 16987 7036 17053 7037
rect 16987 6972 16988 7036
rect 17052 6972 17053 7036
rect 16987 6971 17053 6972
rect 18646 6493 18706 8739
rect 18643 6492 18709 6493
rect 18643 6428 18644 6492
rect 18708 6428 18709 6492
rect 18643 6427 18709 6428
rect 16619 6356 16685 6357
rect 16619 6292 16620 6356
rect 16684 6292 16685 6356
rect 16619 6291 16685 6292
rect 18830 5541 18890 10235
rect 19014 8125 19074 13227
rect 19204 13088 19524 14112
rect 19204 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19524 13088
rect 19204 12000 19524 13024
rect 19204 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19524 12000
rect 19204 10912 19524 11936
rect 19864 21248 20184 21808
rect 19864 21184 19872 21248
rect 19936 21184 19952 21248
rect 20016 21184 20032 21248
rect 20096 21184 20112 21248
rect 20176 21184 20184 21248
rect 19864 20160 20184 21184
rect 19864 20096 19872 20160
rect 19936 20096 19952 20160
rect 20016 20096 20032 20160
rect 20096 20096 20112 20160
rect 20176 20096 20184 20160
rect 19864 19072 20184 20096
rect 19864 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20184 19072
rect 19864 17984 20184 19008
rect 20299 18596 20365 18597
rect 20299 18532 20300 18596
rect 20364 18532 20365 18596
rect 20299 18531 20365 18532
rect 19864 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20184 17984
rect 19864 16896 20184 17920
rect 19864 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20184 16896
rect 19864 15808 20184 16832
rect 19864 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20184 15808
rect 19864 14720 20184 15744
rect 19864 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20184 14720
rect 19864 13632 20184 14656
rect 19864 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20184 13632
rect 19864 12544 20184 13568
rect 19864 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20184 12544
rect 19701 11524 19767 11525
rect 19701 11460 19702 11524
rect 19766 11460 19767 11524
rect 19701 11459 19767 11460
rect 19704 10981 19764 11459
rect 19864 11456 20184 12480
rect 19864 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20184 11456
rect 19701 10980 19767 10981
rect 19701 10916 19702 10980
rect 19766 10916 19767 10980
rect 19701 10915 19767 10916
rect 19204 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19524 10912
rect 19204 9824 19524 10848
rect 19204 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19524 9824
rect 19204 8736 19524 9760
rect 19204 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19524 8736
rect 19011 8124 19077 8125
rect 19011 8060 19012 8124
rect 19076 8060 19077 8124
rect 19011 8059 19077 8060
rect 19204 7648 19524 8672
rect 19204 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19524 7648
rect 19204 6560 19524 7584
rect 19204 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19524 6560
rect 18827 5540 18893 5541
rect 18827 5476 18828 5540
rect 18892 5476 18893 5540
rect 18827 5475 18893 5476
rect 19204 5472 19524 6496
rect 19204 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19524 5472
rect 19204 4384 19524 5408
rect 19204 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19524 4384
rect 16067 3908 16133 3909
rect 16067 3844 16068 3908
rect 16132 3844 16133 3908
rect 16067 3843 16133 3844
rect 19204 3296 19524 4320
rect 19204 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19524 3296
rect 19204 2208 19524 3232
rect 19204 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19524 2208
rect 15883 1460 15949 1461
rect 15883 1396 15884 1460
rect 15948 1396 15949 1460
rect 15883 1395 15949 1396
rect 12090 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12410 576
rect 12090 496 12410 512
rect 19204 1120 19524 2144
rect 19204 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19524 1120
rect 19204 496 19524 1056
rect 19864 10368 20184 11392
rect 20302 10845 20362 18531
rect 20486 11933 20546 21934
rect 24347 21932 24348 21996
rect 24412 21932 24413 21996
rect 24347 21931 24413 21932
rect 21035 21316 21101 21317
rect 21035 21252 21036 21316
rect 21100 21252 21101 21316
rect 21035 21251 21101 21252
rect 21038 20093 21098 21251
rect 24163 20908 24229 20909
rect 24163 20844 24164 20908
rect 24228 20844 24229 20908
rect 24163 20843 24229 20844
rect 21035 20092 21101 20093
rect 21035 20028 21036 20092
rect 21100 20028 21101 20092
rect 21035 20027 21101 20028
rect 20667 19276 20733 19277
rect 20667 19212 20668 19276
rect 20732 19212 20733 19276
rect 20667 19211 20733 19212
rect 20670 14653 20730 19211
rect 20851 14788 20917 14789
rect 20851 14724 20852 14788
rect 20916 14724 20917 14788
rect 20851 14723 20917 14724
rect 20667 14652 20733 14653
rect 20667 14588 20668 14652
rect 20732 14588 20733 14652
rect 20667 14587 20733 14588
rect 20667 13020 20733 13021
rect 20667 12956 20668 13020
rect 20732 12956 20733 13020
rect 20667 12955 20733 12956
rect 20483 11932 20549 11933
rect 20483 11868 20484 11932
rect 20548 11868 20549 11932
rect 20483 11867 20549 11868
rect 20670 11794 20730 12955
rect 20486 11734 20730 11794
rect 20299 10844 20365 10845
rect 20299 10780 20300 10844
rect 20364 10780 20365 10844
rect 20299 10779 20365 10780
rect 20299 10436 20365 10437
rect 20299 10372 20300 10436
rect 20364 10372 20365 10436
rect 20299 10371 20365 10372
rect 19864 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20184 10368
rect 19864 9280 20184 10304
rect 19864 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20184 9280
rect 19864 8192 20184 9216
rect 19864 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20184 8192
rect 19864 7104 20184 8128
rect 20302 7581 20362 10371
rect 20299 7580 20365 7581
rect 20299 7516 20300 7580
rect 20364 7516 20365 7580
rect 20299 7515 20365 7516
rect 19864 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20184 7104
rect 19864 6016 20184 7040
rect 19864 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20184 6016
rect 19864 4928 20184 5952
rect 20302 5405 20362 7515
rect 20486 6901 20546 11734
rect 20667 11524 20733 11525
rect 20667 11460 20668 11524
rect 20732 11460 20733 11524
rect 20667 11459 20733 11460
rect 20483 6900 20549 6901
rect 20483 6836 20484 6900
rect 20548 6836 20549 6900
rect 20483 6835 20549 6836
rect 20299 5404 20365 5405
rect 20299 5340 20300 5404
rect 20364 5340 20365 5404
rect 20299 5339 20365 5340
rect 19864 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20184 4928
rect 19864 3840 20184 4864
rect 19864 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20184 3840
rect 19864 2752 20184 3776
rect 19864 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20184 2752
rect 19864 1664 20184 2688
rect 20670 2413 20730 11459
rect 20854 4861 20914 14723
rect 21038 12885 21098 20027
rect 22507 19548 22573 19549
rect 22507 19484 22508 19548
rect 22572 19484 22573 19548
rect 22507 19483 22573 19484
rect 21955 18052 22021 18053
rect 21955 17988 21956 18052
rect 22020 17988 22021 18052
rect 21955 17987 22021 17988
rect 21219 16284 21285 16285
rect 21219 16220 21220 16284
rect 21284 16220 21285 16284
rect 21219 16219 21285 16220
rect 21035 12884 21101 12885
rect 21035 12820 21036 12884
rect 21100 12820 21101 12884
rect 21035 12819 21101 12820
rect 21222 11930 21282 16219
rect 21771 16012 21837 16013
rect 21771 15948 21772 16012
rect 21836 15948 21837 16012
rect 21771 15947 21837 15948
rect 21403 15468 21469 15469
rect 21403 15404 21404 15468
rect 21468 15404 21469 15468
rect 21403 15403 21469 15404
rect 21038 11870 21282 11930
rect 21038 10437 21098 11870
rect 21219 11796 21285 11797
rect 21219 11732 21220 11796
rect 21284 11732 21285 11796
rect 21219 11731 21285 11732
rect 21035 10436 21101 10437
rect 21035 10372 21036 10436
rect 21100 10372 21101 10436
rect 21035 10371 21101 10372
rect 21035 8804 21101 8805
rect 21035 8740 21036 8804
rect 21100 8740 21101 8804
rect 21035 8739 21101 8740
rect 21038 6357 21098 8739
rect 21035 6356 21101 6357
rect 21035 6292 21036 6356
rect 21100 6292 21101 6356
rect 21035 6291 21101 6292
rect 20851 4860 20917 4861
rect 20851 4796 20852 4860
rect 20916 4796 20917 4860
rect 20851 4795 20917 4796
rect 21222 2549 21282 11731
rect 21406 10301 21466 15403
rect 21774 14378 21834 15947
rect 21958 15605 22018 17987
rect 22323 16828 22389 16829
rect 22323 16764 22324 16828
rect 22388 16764 22389 16828
rect 22323 16763 22389 16764
rect 22139 16556 22205 16557
rect 22139 16492 22140 16556
rect 22204 16492 22205 16556
rect 22139 16491 22205 16492
rect 21955 15604 22021 15605
rect 21955 15540 21956 15604
rect 22020 15540 22021 15604
rect 21955 15539 22021 15540
rect 21774 14318 22018 14378
rect 21771 13972 21837 13973
rect 21771 13908 21772 13972
rect 21836 13908 21837 13972
rect 21771 13907 21837 13908
rect 21587 10572 21653 10573
rect 21587 10508 21588 10572
rect 21652 10508 21653 10572
rect 21587 10507 21653 10508
rect 21403 10300 21469 10301
rect 21403 10236 21404 10300
rect 21468 10236 21469 10300
rect 21403 10235 21469 10236
rect 21219 2548 21285 2549
rect 21219 2484 21220 2548
rect 21284 2484 21285 2548
rect 21219 2483 21285 2484
rect 20667 2412 20733 2413
rect 20667 2348 20668 2412
rect 20732 2348 20733 2412
rect 20667 2347 20733 2348
rect 21590 1869 21650 10507
rect 21774 4181 21834 13907
rect 21958 13018 22018 14318
rect 22142 13837 22202 16491
rect 22326 16285 22386 16763
rect 22510 16557 22570 19483
rect 22691 17100 22757 17101
rect 22691 17036 22692 17100
rect 22756 17036 22757 17100
rect 22691 17035 22757 17036
rect 22507 16556 22573 16557
rect 22507 16492 22508 16556
rect 22572 16492 22573 16556
rect 22507 16491 22573 16492
rect 22323 16284 22389 16285
rect 22323 16220 22324 16284
rect 22388 16220 22389 16284
rect 22323 16219 22389 16220
rect 22139 13836 22205 13837
rect 22139 13772 22140 13836
rect 22204 13772 22205 13836
rect 22139 13771 22205 13772
rect 22326 13565 22386 16219
rect 22507 16012 22573 16013
rect 22507 15948 22508 16012
rect 22572 15948 22573 16012
rect 22507 15947 22573 15948
rect 22323 13564 22389 13565
rect 22323 13500 22324 13564
rect 22388 13500 22389 13564
rect 22323 13499 22389 13500
rect 21958 12958 22386 13018
rect 21955 12884 22021 12885
rect 21955 12820 21956 12884
rect 22020 12820 22021 12884
rect 21955 12819 22021 12820
rect 22139 12884 22205 12885
rect 22139 12820 22140 12884
rect 22204 12820 22205 12884
rect 22139 12819 22205 12820
rect 21958 11933 22018 12819
rect 21955 11932 22021 11933
rect 21955 11868 21956 11932
rect 22020 11868 22021 11932
rect 21955 11867 22021 11868
rect 21958 8261 22018 11867
rect 22142 8805 22202 12819
rect 22139 8804 22205 8805
rect 22139 8740 22140 8804
rect 22204 8740 22205 8804
rect 22139 8739 22205 8740
rect 21955 8260 22021 8261
rect 21955 8196 21956 8260
rect 22020 8196 22021 8260
rect 21955 8195 22021 8196
rect 22326 8125 22386 12958
rect 22510 8261 22570 15947
rect 22694 9893 22754 17035
rect 23059 15604 23125 15605
rect 23059 15540 23060 15604
rect 23124 15540 23125 15604
rect 23059 15539 23125 15540
rect 23243 15604 23309 15605
rect 23243 15540 23244 15604
rect 23308 15540 23309 15604
rect 23243 15539 23309 15540
rect 22875 11524 22941 11525
rect 22875 11460 22876 11524
rect 22940 11460 22941 11524
rect 22875 11459 22941 11460
rect 22691 9892 22757 9893
rect 22691 9828 22692 9892
rect 22756 9828 22757 9892
rect 22691 9827 22757 9828
rect 22878 9621 22938 11459
rect 22875 9620 22941 9621
rect 22875 9556 22876 9620
rect 22940 9556 22941 9620
rect 22875 9555 22941 9556
rect 23062 9077 23122 15539
rect 23059 9076 23125 9077
rect 23059 9012 23060 9076
rect 23124 9012 23125 9076
rect 23059 9011 23125 9012
rect 23246 8261 23306 15539
rect 24166 14517 24226 20843
rect 24163 14516 24229 14517
rect 24163 14452 24164 14516
rect 24228 14452 24229 14516
rect 24163 14451 24229 14452
rect 24350 13565 24410 21931
rect 26978 21792 27298 21808
rect 26978 21728 26986 21792
rect 27050 21728 27066 21792
rect 27130 21728 27146 21792
rect 27210 21728 27226 21792
rect 27290 21728 27298 21792
rect 25819 21588 25885 21589
rect 25819 21524 25820 21588
rect 25884 21524 25885 21588
rect 25819 21523 25885 21524
rect 24715 19820 24781 19821
rect 24715 19756 24716 19820
rect 24780 19756 24781 19820
rect 24715 19755 24781 19756
rect 24718 18869 24778 19755
rect 24715 18868 24781 18869
rect 24715 18804 24716 18868
rect 24780 18804 24781 18868
rect 24715 18803 24781 18804
rect 25822 17509 25882 21523
rect 26555 21452 26621 21453
rect 26555 21388 26556 21452
rect 26620 21388 26621 21452
rect 26555 21387 26621 21388
rect 26187 20500 26253 20501
rect 26187 20436 26188 20500
rect 26252 20436 26253 20500
rect 26187 20435 26253 20436
rect 26003 19548 26069 19549
rect 26003 19484 26004 19548
rect 26068 19484 26069 19548
rect 26003 19483 26069 19484
rect 26006 17917 26066 19483
rect 26003 17916 26069 17917
rect 26003 17852 26004 17916
rect 26068 17852 26069 17916
rect 26003 17851 26069 17852
rect 25819 17508 25885 17509
rect 25819 17444 25820 17508
rect 25884 17444 25885 17508
rect 25819 17443 25885 17444
rect 26190 16557 26250 20435
rect 26187 16556 26253 16557
rect 26187 16492 26188 16556
rect 26252 16492 26253 16556
rect 26187 16491 26253 16492
rect 26187 16420 26253 16421
rect 26187 16356 26188 16420
rect 26252 16356 26253 16420
rect 26187 16355 26253 16356
rect 26190 15741 26250 16355
rect 26187 15740 26253 15741
rect 26187 15676 26188 15740
rect 26252 15676 26253 15740
rect 26187 15675 26253 15676
rect 26371 15740 26437 15741
rect 26371 15676 26372 15740
rect 26436 15676 26437 15740
rect 26371 15675 26437 15676
rect 25819 15196 25885 15197
rect 25819 15132 25820 15196
rect 25884 15132 25885 15196
rect 25819 15131 25885 15132
rect 24531 13836 24597 13837
rect 24531 13772 24532 13836
rect 24596 13772 24597 13836
rect 24531 13771 24597 13772
rect 24347 13564 24413 13565
rect 24347 13500 24348 13564
rect 24412 13500 24413 13564
rect 24347 13499 24413 13500
rect 23611 8396 23677 8397
rect 23611 8332 23612 8396
rect 23676 8332 23677 8396
rect 23611 8331 23677 8332
rect 22507 8260 22573 8261
rect 22507 8196 22508 8260
rect 22572 8196 22573 8260
rect 22507 8195 22573 8196
rect 23243 8260 23309 8261
rect 23243 8196 23244 8260
rect 23308 8196 23309 8260
rect 23243 8195 23309 8196
rect 22323 8124 22389 8125
rect 22323 8060 22324 8124
rect 22388 8060 22389 8124
rect 22323 8059 22389 8060
rect 21771 4180 21837 4181
rect 21771 4116 21772 4180
rect 21836 4116 21837 4180
rect 21771 4115 21837 4116
rect 23614 2277 23674 8331
rect 24534 6901 24594 13771
rect 25267 13020 25333 13021
rect 25267 12956 25268 13020
rect 25332 12956 25333 13020
rect 25267 12955 25333 12956
rect 25083 10844 25149 10845
rect 25083 10780 25084 10844
rect 25148 10842 25149 10844
rect 25270 10842 25330 12955
rect 25635 12068 25701 12069
rect 25635 12004 25636 12068
rect 25700 12004 25701 12068
rect 25635 12003 25701 12004
rect 25148 10782 25330 10842
rect 25148 10780 25149 10782
rect 25083 10779 25149 10780
rect 24899 10300 24965 10301
rect 24899 10236 24900 10300
rect 24964 10236 24965 10300
rect 24899 10235 24965 10236
rect 24715 9892 24781 9893
rect 24715 9828 24716 9892
rect 24780 9828 24781 9892
rect 24715 9827 24781 9828
rect 24718 7989 24778 9827
rect 24715 7988 24781 7989
rect 24715 7924 24716 7988
rect 24780 7924 24781 7988
rect 24715 7923 24781 7924
rect 24902 7717 24962 10235
rect 24899 7716 24965 7717
rect 24899 7652 24900 7716
rect 24964 7652 24965 7716
rect 24899 7651 24965 7652
rect 24531 6900 24597 6901
rect 24531 6836 24532 6900
rect 24596 6836 24597 6900
rect 24531 6835 24597 6836
rect 25086 5677 25146 10779
rect 25451 9620 25517 9621
rect 25451 9556 25452 9620
rect 25516 9556 25517 9620
rect 25451 9555 25517 9556
rect 25454 9077 25514 9555
rect 25451 9076 25517 9077
rect 25451 9012 25452 9076
rect 25516 9012 25517 9076
rect 25451 9011 25517 9012
rect 25083 5676 25149 5677
rect 25083 5612 25084 5676
rect 25148 5612 25149 5676
rect 25083 5611 25149 5612
rect 25638 2685 25698 12003
rect 25822 8669 25882 15131
rect 26003 14380 26069 14381
rect 26003 14316 26004 14380
rect 26068 14316 26069 14380
rect 26003 14315 26069 14316
rect 26006 12341 26066 14315
rect 26003 12340 26069 12341
rect 26003 12276 26004 12340
rect 26068 12276 26069 12340
rect 26003 12275 26069 12276
rect 26190 11525 26250 15675
rect 26187 11524 26253 11525
rect 26187 11460 26188 11524
rect 26252 11460 26253 11524
rect 26187 11459 26253 11460
rect 26374 11389 26434 15675
rect 26371 11388 26437 11389
rect 26371 11324 26372 11388
rect 26436 11324 26437 11388
rect 26371 11323 26437 11324
rect 26558 11117 26618 21387
rect 26978 20704 27298 21728
rect 27638 21248 27958 21808
rect 27638 21184 27646 21248
rect 27710 21184 27726 21248
rect 27790 21184 27806 21248
rect 27870 21184 27886 21248
rect 27950 21184 27958 21248
rect 27475 21044 27541 21045
rect 27475 20980 27476 21044
rect 27540 20980 27541 21044
rect 27475 20979 27541 20980
rect 26978 20640 26986 20704
rect 27050 20640 27066 20704
rect 27130 20640 27146 20704
rect 27210 20640 27226 20704
rect 27290 20640 27298 20704
rect 26978 19616 27298 20640
rect 26978 19552 26986 19616
rect 27050 19552 27066 19616
rect 27130 19552 27146 19616
rect 27210 19552 27226 19616
rect 27290 19552 27298 19616
rect 26978 18528 27298 19552
rect 26978 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27298 18528
rect 26739 18188 26805 18189
rect 26739 18124 26740 18188
rect 26804 18124 26805 18188
rect 26739 18123 26805 18124
rect 26742 13973 26802 18123
rect 26978 17440 27298 18464
rect 26978 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27298 17440
rect 26978 16352 27298 17376
rect 26978 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27298 16352
rect 26978 15264 27298 16288
rect 27478 15333 27538 20979
rect 27638 20160 27958 21184
rect 27638 20096 27646 20160
rect 27710 20096 27726 20160
rect 27790 20096 27806 20160
rect 27870 20096 27886 20160
rect 27950 20096 27958 20160
rect 27638 19072 27958 20096
rect 27638 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27958 19072
rect 27638 17984 27958 19008
rect 27638 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27958 17984
rect 27638 16896 27958 17920
rect 28027 17372 28093 17373
rect 28027 17308 28028 17372
rect 28092 17308 28093 17372
rect 28027 17307 28093 17308
rect 27638 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27958 16896
rect 27638 15808 27958 16832
rect 28030 15877 28090 17307
rect 28214 16421 28274 22304
rect 28766 19277 28826 22304
rect 28763 19276 28829 19277
rect 28763 19212 28764 19276
rect 28828 19212 28829 19276
rect 28763 19211 28829 19212
rect 28395 17780 28461 17781
rect 28395 17716 28396 17780
rect 28460 17716 28461 17780
rect 28395 17715 28461 17716
rect 28398 16693 28458 17715
rect 28395 16692 28461 16693
rect 28395 16628 28396 16692
rect 28460 16628 28461 16692
rect 28395 16627 28461 16628
rect 29318 16557 29378 22304
rect 29867 18460 29933 18461
rect 29867 18396 29868 18460
rect 29932 18396 29933 18460
rect 29867 18395 29933 18396
rect 29499 17100 29565 17101
rect 29499 17036 29500 17100
rect 29564 17036 29565 17100
rect 29499 17035 29565 17036
rect 29315 16556 29381 16557
rect 29315 16492 29316 16556
rect 29380 16492 29381 16556
rect 29315 16491 29381 16492
rect 28211 16420 28277 16421
rect 28211 16356 28212 16420
rect 28276 16356 28277 16420
rect 28211 16355 28277 16356
rect 28027 15876 28093 15877
rect 28027 15812 28028 15876
rect 28092 15812 28093 15876
rect 28027 15811 28093 15812
rect 27638 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27958 15808
rect 27475 15332 27541 15333
rect 27475 15268 27476 15332
rect 27540 15268 27541 15332
rect 27475 15267 27541 15268
rect 26978 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27298 15264
rect 26978 14176 27298 15200
rect 26978 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27298 14176
rect 26739 13972 26805 13973
rect 26739 13908 26740 13972
rect 26804 13908 26805 13972
rect 26739 13907 26805 13908
rect 26739 13700 26805 13701
rect 26739 13636 26740 13700
rect 26804 13636 26805 13700
rect 26739 13635 26805 13636
rect 26742 12885 26802 13635
rect 26978 13088 27298 14112
rect 26978 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27298 13088
rect 26739 12884 26805 12885
rect 26739 12820 26740 12884
rect 26804 12820 26805 12884
rect 26739 12819 26805 12820
rect 26555 11116 26621 11117
rect 26555 11052 26556 11116
rect 26620 11052 26621 11116
rect 26555 11051 26621 11052
rect 26555 9756 26621 9757
rect 26555 9692 26556 9756
rect 26620 9692 26621 9756
rect 26555 9691 26621 9692
rect 26187 9212 26253 9213
rect 26187 9148 26188 9212
rect 26252 9148 26253 9212
rect 26187 9147 26253 9148
rect 25819 8668 25885 8669
rect 25819 8604 25820 8668
rect 25884 8604 25885 8668
rect 25819 8603 25885 8604
rect 25822 8125 25882 8603
rect 25819 8124 25885 8125
rect 25819 8060 25820 8124
rect 25884 8060 25885 8124
rect 25819 8059 25885 8060
rect 26190 4045 26250 9147
rect 26558 8125 26618 9691
rect 26742 9077 26802 12819
rect 26978 12000 27298 13024
rect 26978 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27298 12000
rect 26978 10912 27298 11936
rect 26978 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27298 10912
rect 26978 9824 27298 10848
rect 26978 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27298 9824
rect 26739 9076 26805 9077
rect 26739 9012 26740 9076
rect 26804 9012 26805 9076
rect 26739 9011 26805 9012
rect 26978 8736 27298 9760
rect 26978 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27298 8736
rect 26555 8124 26621 8125
rect 26555 8060 26556 8124
rect 26620 8060 26621 8124
rect 26555 8059 26621 8060
rect 26978 7648 27298 8672
rect 27638 14720 27958 15744
rect 28579 15604 28645 15605
rect 28579 15540 28580 15604
rect 28644 15540 28645 15604
rect 28579 15539 28645 15540
rect 29131 15604 29197 15605
rect 29131 15540 29132 15604
rect 29196 15540 29197 15604
rect 29131 15539 29197 15540
rect 28027 15468 28093 15469
rect 28027 15404 28028 15468
rect 28092 15404 28093 15468
rect 28027 15403 28093 15404
rect 28211 15468 28277 15469
rect 28211 15404 28212 15468
rect 28276 15404 28277 15468
rect 28211 15403 28277 15404
rect 27638 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27958 14720
rect 27638 13632 27958 14656
rect 27638 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27958 13632
rect 27638 12544 27958 13568
rect 27638 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27958 12544
rect 27638 11456 27958 12480
rect 28030 11933 28090 15403
rect 28214 13429 28274 15403
rect 28211 13428 28277 13429
rect 28211 13364 28212 13428
rect 28276 13364 28277 13428
rect 28211 13363 28277 13364
rect 28027 11932 28093 11933
rect 28027 11868 28028 11932
rect 28092 11868 28093 11932
rect 28027 11867 28093 11868
rect 27638 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27958 11456
rect 27638 10368 27958 11392
rect 27638 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27958 10368
rect 27638 9280 27958 10304
rect 27638 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27958 9280
rect 27475 8396 27541 8397
rect 27475 8332 27476 8396
rect 27540 8332 27541 8396
rect 27475 8331 27541 8332
rect 27478 7853 27538 8331
rect 27638 8192 27958 9216
rect 27638 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27958 8192
rect 27475 7852 27541 7853
rect 27475 7788 27476 7852
rect 27540 7788 27541 7852
rect 27475 7787 27541 7788
rect 26978 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27298 7648
rect 26978 6560 27298 7584
rect 27478 7037 27538 7787
rect 27638 7104 27958 8128
rect 28214 7717 28274 13363
rect 28395 11796 28461 11797
rect 28395 11732 28396 11796
rect 28460 11732 28461 11796
rect 28395 11731 28461 11732
rect 28398 9213 28458 11731
rect 28395 9212 28461 9213
rect 28395 9148 28396 9212
rect 28460 9148 28461 9212
rect 28395 9147 28461 9148
rect 28211 7716 28277 7717
rect 28211 7652 28212 7716
rect 28276 7652 28277 7716
rect 28211 7651 28277 7652
rect 27638 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27958 7104
rect 27475 7036 27541 7037
rect 27475 6972 27476 7036
rect 27540 6972 27541 7036
rect 27475 6971 27541 6972
rect 26978 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27298 6560
rect 26978 5472 27298 6496
rect 26978 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27298 5472
rect 26978 4384 27298 5408
rect 26978 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27298 4384
rect 26187 4044 26253 4045
rect 26187 3980 26188 4044
rect 26252 3980 26253 4044
rect 26187 3979 26253 3980
rect 26978 3296 27298 4320
rect 26978 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27298 3296
rect 25635 2684 25701 2685
rect 25635 2620 25636 2684
rect 25700 2620 25701 2684
rect 25635 2619 25701 2620
rect 23611 2276 23677 2277
rect 23611 2212 23612 2276
rect 23676 2212 23677 2276
rect 23611 2211 23677 2212
rect 26978 2208 27298 3232
rect 26978 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27298 2208
rect 21587 1868 21653 1869
rect 21587 1804 21588 1868
rect 21652 1804 21653 1868
rect 21587 1803 21653 1804
rect 19864 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20184 1664
rect 19864 576 20184 1600
rect 19864 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20184 576
rect 19864 496 20184 512
rect 26978 1120 27298 2144
rect 26978 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27298 1120
rect 26978 496 27298 1056
rect 27638 6016 27958 7040
rect 27638 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27958 6016
rect 27638 4928 27958 5952
rect 28582 5133 28642 15539
rect 28763 13972 28829 13973
rect 28763 13908 28764 13972
rect 28828 13908 28829 13972
rect 28763 13907 28829 13908
rect 28766 9690 28826 13907
rect 29134 12341 29194 15539
rect 29502 13837 29562 17035
rect 29870 14789 29930 18395
rect 30235 15332 30301 15333
rect 30235 15268 30236 15332
rect 30300 15268 30301 15332
rect 30235 15267 30301 15268
rect 29867 14788 29933 14789
rect 29867 14724 29868 14788
rect 29932 14724 29933 14788
rect 29867 14723 29933 14724
rect 29499 13836 29565 13837
rect 29499 13772 29500 13836
rect 29564 13772 29565 13836
rect 29499 13771 29565 13772
rect 29499 12476 29565 12477
rect 29499 12412 29500 12476
rect 29564 12412 29565 12476
rect 29499 12411 29565 12412
rect 29131 12340 29197 12341
rect 29131 12276 29132 12340
rect 29196 12276 29197 12340
rect 29131 12275 29197 12276
rect 28766 9630 29194 9690
rect 29134 9485 29194 9630
rect 29131 9484 29197 9485
rect 29131 9420 29132 9484
rect 29196 9420 29197 9484
rect 29131 9419 29197 9420
rect 29134 8397 29194 9419
rect 29502 9349 29562 12411
rect 30238 10573 30298 15267
rect 30235 10572 30301 10573
rect 30235 10508 30236 10572
rect 30300 10508 30301 10572
rect 30235 10507 30301 10508
rect 29499 9348 29565 9349
rect 29499 9284 29500 9348
rect 29564 9284 29565 9348
rect 29499 9283 29565 9284
rect 30238 8941 30298 10507
rect 30235 8940 30301 8941
rect 30235 8876 30236 8940
rect 30300 8876 30301 8940
rect 30235 8875 30301 8876
rect 29131 8396 29197 8397
rect 29131 8332 29132 8396
rect 29196 8332 29197 8396
rect 29131 8331 29197 8332
rect 28579 5132 28645 5133
rect 28579 5068 28580 5132
rect 28644 5068 28645 5132
rect 28579 5067 28645 5068
rect 27638 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27958 4928
rect 27638 3840 27958 4864
rect 27638 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27958 3840
rect 27638 2752 27958 3776
rect 27638 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27958 2752
rect 27638 1664 27958 2688
rect 27638 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27958 1664
rect 27638 576 27958 1600
rect 27638 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27958 576
rect 27638 496 27958 512
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 0
transform 1 0 31096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 0
transform 1 0 14260 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 0
transform -1 0 13800 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 0
transform 1 0 3864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 0
transform -1 0 4508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 0
transform 1 0 5796 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 0
transform -1 0 6532 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 0
transform -1 0 25576 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 0
transform -1 0 30912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 0
transform -1 0 23644 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 0
transform 1 0 30636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 0
transform -1 0 29532 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 0
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 0
transform 1 0 26772 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 0
transform -1 0 11040 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 0
transform -1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0803_
timestamp 0
transform 1 0 7912 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0804_
timestamp 0
transform 1 0 8372 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0805_
timestamp 0
transform -1 0 11500 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0806_
timestamp 0
transform -1 0 10856 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0807_
timestamp 0
transform 1 0 11408 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0808_
timestamp 0
transform -1 0 11776 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0809_
timestamp 0
transform 1 0 10120 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0810_
timestamp 0
transform -1 0 9292 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0811_
timestamp 0
transform -1 0 25944 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0812_
timestamp 0
transform 1 0 15272 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0813_
timestamp 0
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0814_
timestamp 0
transform -1 0 7084 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0815_
timestamp 0
transform 1 0 17020 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0816_
timestamp 0
transform -1 0 10856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 0
transform -1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 0
transform 1 0 1564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 0
transform 1 0 19044 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 0
transform 1 0 24288 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _0821_
timestamp 0
transform 1 0 29348 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0822_
timestamp 0
transform -1 0 18584 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _0823_
timestamp 0
transform 1 0 1748 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0824_
timestamp 0
transform -1 0 5612 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_2  _0825_
timestamp 0
transform 1 0 3220 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0826_
timestamp 0
transform -1 0 20424 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _0827_
timestamp 0
transform 1 0 19596 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0828_
timestamp 0
transform 1 0 23828 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0829_
timestamp 0
transform -1 0 2668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0830_
timestamp 0
transform -1 0 10580 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0831_
timestamp 0
transform -1 0 28888 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0832_
timestamp 0
transform -1 0 19596 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0833_
timestamp 0
transform -1 0 19228 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0834_
timestamp 0
transform 1 0 9200 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0835_
timestamp 0
transform -1 0 30544 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0836_
timestamp 0
transform -1 0 28520 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 0
transform 1 0 23184 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _0838_
timestamp 0
transform 1 0 24932 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__o211a_2  _0839_
timestamp 0
transform 1 0 2392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _0840_
timestamp 0
transform 1 0 29624 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0841_
timestamp 0
transform -1 0 22080 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0842_
timestamp 0
transform 1 0 26772 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0843_
timestamp 0
transform -1 0 6256 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _0844_
timestamp 0
transform 1 0 18676 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0845_
timestamp 0
transform 1 0 1288 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0846_
timestamp 0
transform 1 0 6532 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _0847_
timestamp 0
transform -1 0 26312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0848_
timestamp 0
transform -1 0 30360 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0849_
timestamp 0
transform -1 0 26128 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 0
transform -1 0 16284 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0851_
timestamp 0
transform -1 0 28060 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_4  _0852_
timestamp 0
transform 1 0 29532 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _0853_
timestamp 0
transform -1 0 23184 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 0
transform -1 0 25944 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0855_
timestamp 0
transform 1 0 25484 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _0856_
timestamp 0
transform 1 0 2944 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__a311oi_4  _0857_
timestamp 0
transform 1 0 26680 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_2  _0858_
timestamp 0
transform 1 0 18676 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0859_
timestamp 0
transform 1 0 27508 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0860_
timestamp 0
transform -1 0 28060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0861_
timestamp 0
transform -1 0 27508 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 0
transform -1 0 13892 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _0863_
timestamp 0
transform -1 0 27324 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0864_
timestamp 0
transform 1 0 26036 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0865_
timestamp 0
transform -1 0 17940 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_4  _0866_
timestamp 0
transform 1 0 1564 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_1  _0867_
timestamp 0
transform 1 0 28980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0868_
timestamp 0
transform 1 0 26772 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0869_
timestamp 0
transform 1 0 24748 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 0
transform -1 0 28980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0871_
timestamp 0
transform 1 0 29072 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0872_
timestamp 0
transform -1 0 24748 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0873_
timestamp 0
transform 1 0 3220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _0874_
timestamp 0
transform -1 0 19596 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _0875_
timestamp 0
transform -1 0 31280 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 0
transform -1 0 15732 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 0
transform 1 0 20240 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 0
transform 1 0 17020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0879_
timestamp 0
transform -1 0 23460 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0880_
timestamp 0
transform 1 0 27140 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0881_
timestamp 0
transform -1 0 24472 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0882_
timestamp 0
transform -1 0 29164 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0883_
timestamp 0
transform -1 0 19136 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _0884_
timestamp 0
transform -1 0 30636 0 -1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 0
transform -1 0 24288 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0886_
timestamp 0
transform 1 0 23460 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0887_
timestamp 0
transform -1 0 23552 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0888_
timestamp 0
transform -1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 0
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0890_
timestamp 0
transform -1 0 15180 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0891_
timestamp 0
transform -1 0 12052 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _0892_
timestamp 0
transform -1 0 26036 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 0
transform 1 0 12788 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0894_
timestamp 0
transform 1 0 4784 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0895_
timestamp 0
transform -1 0 4600 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0896_
timestamp 0
transform -1 0 16008 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0897_
timestamp 0
transform -1 0 15088 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 0
transform 1 0 18032 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _0899_
timestamp 0
transform -1 0 30544 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0900_
timestamp 0
transform 1 0 29808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 0
transform 1 0 29072 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 0
transform -1 0 12328 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0903_
timestamp 0
transform 1 0 19228 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _0904_
timestamp 0
transform -1 0 2116 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _0905_
timestamp 0
transform 1 0 25116 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__a211oi_1  _0906_
timestamp 0
transform 1 0 1288 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0907_
timestamp 0
transform -1 0 2484 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0908_
timestamp 0
transform 1 0 4968 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0909_
timestamp 0
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _0910_
timestamp 0
transform -1 0 22080 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _0911_
timestamp 0
transform 1 0 29808 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__o2111a_1  _0912_
timestamp 0
transform 1 0 24104 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_4  _0913_
timestamp 0
transform 1 0 1104 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 0
transform 1 0 7912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 0
transform -1 0 18676 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _0916_
timestamp 0
transform -1 0 28704 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0917_
timestamp 0
transform -1 0 20148 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 0
transform -1 0 21988 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0919_
timestamp 0
transform 1 0 21068 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0920_
timestamp 0
transform -1 0 20056 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 0
transform 1 0 19228 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0922_
timestamp 0
transform -1 0 14996 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0923_
timestamp 0
transform 1 0 3864 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0924_
timestamp 0
transform 1 0 10120 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0925_
timestamp 0
transform 1 0 3220 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0926_
timestamp 0
transform 1 0 7544 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 0
transform 1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0928_
timestamp 0
transform 1 0 21344 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0929_
timestamp 0
transform -1 0 28796 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _0930_
timestamp 0
transform -1 0 5980 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0931_
timestamp 0
transform -1 0 29624 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 0
transform -1 0 23092 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0933_
timestamp 0
transform -1 0 18400 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0934_
timestamp 0
transform -1 0 11592 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0935_
timestamp 0
transform -1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _0936_
timestamp 0
transform -1 0 2760 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0937_
timestamp 0
transform 1 0 5244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0938_
timestamp 0
transform 1 0 8372 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0939_
timestamp 0
transform -1 0 11960 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0940_
timestamp 0
transform -1 0 23368 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0941_
timestamp 0
transform -1 0 11960 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0942_
timestamp 0
transform -1 0 18124 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0943_
timestamp 0
transform -1 0 18216 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0944_
timestamp 0
transform 1 0 5060 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_4  _0945_
timestamp 0
transform -1 0 2852 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 0
transform 1 0 26956 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 0
transform -1 0 7820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _0948_
timestamp 0
transform 1 0 15272 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _0949_
timestamp 0
transform 1 0 22356 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0950_
timestamp 0
transform -1 0 17940 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0951_
timestamp 0
transform -1 0 4416 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0952_
timestamp 0
transform 1 0 2392 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0953_
timestamp 0
transform -1 0 24196 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0954_
timestamp 0
transform 1 0 14536 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0955_
timestamp 0
transform 1 0 28980 0 1 15776
box -38 -48 1050 592
use sky130_fd_sc_hd__a22o_1  _0956_
timestamp 0
transform 1 0 16652 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0957_
timestamp 0
transform -1 0 29808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0958_
timestamp 0
transform 1 0 27968 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0959_
timestamp 0
transform 1 0 19320 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0960_
timestamp 0
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0961_
timestamp 0
transform -1 0 5244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0962_
timestamp 0
transform 1 0 4232 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0963_
timestamp 0
transform -1 0 5704 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0964_
timestamp 0
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0965_
timestamp 0
transform -1 0 20148 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0966_
timestamp 0
transform 1 0 18676 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0967_
timestamp 0
transform 1 0 17020 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 0
transform 1 0 24380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0969_
timestamp 0
transform 1 0 3772 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o311ai_4  _0970_
timestamp 0
transform -1 0 30912 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _0971_
timestamp 0
transform -1 0 25208 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0972_
timestamp 0
transform 1 0 23920 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0973_
timestamp 0
transform 1 0 12328 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0974_
timestamp 0
transform -1 0 13432 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_4  _0975_
timestamp 0
transform -1 0 2852 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__o211ai_1  _0976_
timestamp 0
transform 1 0 16468 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0977_
timestamp 0
transform 1 0 17112 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0978_
timestamp 0
transform -1 0 21160 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 0
transform -1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0980_
timestamp 0
transform -1 0 1564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0981_
timestamp 0
transform 1 0 21896 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0982_
timestamp 0
transform -1 0 21712 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0983_
timestamp 0
transform 1 0 20424 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0984_
timestamp 0
transform 1 0 22448 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _0985_
timestamp 0
transform -1 0 27508 0 -1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0986_
timestamp 0
transform -1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0987_
timestamp 0
transform 1 0 1196 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0988_
timestamp 0
transform 1 0 30636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 0
transform -1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0990_
timestamp 0
transform -1 0 11684 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0991_
timestamp 0
transform -1 0 18860 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0992_
timestamp 0
transform 1 0 16836 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0993_
timestamp 0
transform 1 0 16836 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0994_
timestamp 0
transform -1 0 4416 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0995_
timestamp 0
transform -1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 0
transform -1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0997_
timestamp 0
transform 1 0 12236 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0998_
timestamp 0
transform 1 0 12512 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0999_
timestamp 0
transform 1 0 23920 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1000_
timestamp 0
transform -1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1001_
timestamp 0
transform 1 0 19688 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1002_
timestamp 0
transform 1 0 10212 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1003_
timestamp 0
transform -1 0 11868 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1004_
timestamp 0
transform 1 0 4416 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1005_
timestamp 0
transform -1 0 6992 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1006_
timestamp 0
transform 1 0 4600 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 0
transform 1 0 10764 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1008_
timestamp 0
transform -1 0 6900 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1009_
timestamp 0
transform -1 0 3588 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _1010_
timestamp 0
transform 1 0 3496 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _1011_
timestamp 0
transform 1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1012_
timestamp 0
transform -1 0 10212 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 0
transform -1 0 9200 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1014_
timestamp 0
transform 1 0 8280 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1015_
timestamp 0
transform 1 0 4600 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 0
transform 1 0 3588 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1017_
timestamp 0
transform -1 0 1472 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 0
transform 1 0 4508 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1019_
timestamp 0
transform -1 0 5428 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1020_
timestamp 0
transform 1 0 7360 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 0
transform -1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1022_
timestamp 0
transform -1 0 7820 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1023_
timestamp 0
transform -1 0 7268 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _1024_
timestamp 0
transform 1 0 12604 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_2  _1025_
timestamp 0
transform -1 0 13984 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _1026_
timestamp 0
transform -1 0 3772 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1027_
timestamp 0
transform -1 0 5152 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1028_
timestamp 0
transform 1 0 4968 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1029_
timestamp 0
transform -1 0 6624 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_1  _1030_
timestamp 0
transform 1 0 7360 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1031_
timestamp 0
transform -1 0 6624 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1032_
timestamp 0
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1033_
timestamp 0
transform 1 0 12420 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 0
transform -1 0 19504 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1035_
timestamp 0
transform -1 0 24288 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1036_
timestamp 0
transform 1 0 3956 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1037_
timestamp 0
transform 1 0 2852 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1038_
timestamp 0
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 0
transform -1 0 29900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1040_
timestamp 0
transform 1 0 14260 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_4  _1041_
timestamp 0
transform -1 0 31280 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__a21bo_1  _1042_
timestamp 0
transform -1 0 29992 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1043_
timestamp 0
transform -1 0 25668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1044_
timestamp 0
transform -1 0 29072 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1045_
timestamp 0
transform 1 0 29624 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1046_
timestamp 0
transform 1 0 28980 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1047_
timestamp 0
transform -1 0 20792 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 0
transform -1 0 18216 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1049_
timestamp 0
transform -1 0 7820 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1050_
timestamp 0
transform 1 0 5060 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1051_
timestamp 0
transform 1 0 4600 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1052_
timestamp 0
transform -1 0 4876 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1053_
timestamp 0
transform -1 0 19228 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 0
transform -1 0 18124 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1055_
timestamp 0
transform 1 0 1288 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1056_
timestamp 0
transform -1 0 1748 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1057_
timestamp 0
transform -1 0 24104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1058_
timestamp 0
transform 1 0 1656 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1059_
timestamp 0
transform -1 0 7452 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1060_
timestamp 0
transform -1 0 3680 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1061_
timestamp 0
transform 1 0 3220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1062_
timestamp 0
transform -1 0 4232 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1063_
timestamp 0
transform 1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1064_
timestamp 0
transform 1 0 20240 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1065_
timestamp 0
transform 1 0 25668 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1066_
timestamp 0
transform 1 0 7636 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 0
transform -1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 0
transform 1 0 20148 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1069_
timestamp 0
transform 1 0 19780 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 0
transform 1 0 3128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1071_
timestamp 0
transform 1 0 3128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1072_
timestamp 0
transform -1 0 5980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1073_
timestamp 0
transform -1 0 5520 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1074_
timestamp 0
transform -1 0 5520 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1075_
timestamp 0
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 0
transform 1 0 17848 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1077_
timestamp 0
transform 1 0 4508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 0
transform -1 0 4416 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1079_
timestamp 0
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1080_
timestamp 0
transform 1 0 3312 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1081_
timestamp 0
transform 1 0 5888 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1082_
timestamp 0
transform 1 0 4968 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1083_
timestamp 0
transform 1 0 5152 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1084_
timestamp 0
transform 1 0 26128 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1085_
timestamp 0
transform -1 0 20792 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1086_
timestamp 0
transform -1 0 25300 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1087_
timestamp 0
transform 1 0 5060 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1088_
timestamp 0
transform 1 0 4876 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1089_
timestamp 0
transform -1 0 6164 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1090_
timestamp 0
transform -1 0 5704 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1091_
timestamp 0
transform -1 0 6440 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 0
transform -1 0 14076 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _1093_
timestamp 0
transform 1 0 20516 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1094_
timestamp 0
transform 1 0 20700 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1095_
timestamp 0
transform 1 0 26496 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1096_
timestamp 0
transform 1 0 21528 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1097_
timestamp 0
transform -1 0 21896 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 0
transform 1 0 28060 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1099_
timestamp 0
transform -1 0 27692 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _1100_
timestamp 0
transform 1 0 29992 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1101_
timestamp 0
transform 1 0 29808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1102_
timestamp 0
transform -1 0 30544 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1103_
timestamp 0
transform 1 0 28704 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1104_
timestamp 0
transform 1 0 27048 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1105_
timestamp 0
transform 1 0 26404 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1106_
timestamp 0
transform 1 0 25392 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1107_
timestamp 0
transform -1 0 26680 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1108_
timestamp 0
transform 1 0 12512 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1109_
timestamp 0
transform 1 0 12512 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1110_
timestamp 0
transform -1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 0
transform -1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1112_
timestamp 0
transform 1 0 10948 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1113_
timestamp 0
transform 1 0 12052 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 0
transform -1 0 24840 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1115_
timestamp 0
transform 1 0 11592 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1116_
timestamp 0
transform 1 0 2024 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _1117_
timestamp 0
transform 1 0 7452 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1118_
timestamp 0
transform 1 0 6532 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_1  _1119_
timestamp 0
transform -1 0 8924 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1120_
timestamp 0
transform 1 0 7544 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1121_
timestamp 0
transform 1 0 6808 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1122_
timestamp 0
transform -1 0 25024 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1123_
timestamp 0
transform 1 0 24656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1124_
timestamp 0
transform -1 0 25300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1125_
timestamp 0
transform -1 0 7728 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1126_
timestamp 0
transform -1 0 8832 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _1127_
timestamp 0
transform 1 0 14444 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1128_
timestamp 0
transform -1 0 9568 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1129_
timestamp 0
transform 1 0 8372 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1130_
timestamp 0
transform -1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1131_
timestamp 0
transform 1 0 18676 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1132_
timestamp 0
transform 1 0 1932 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1133_
timestamp 0
transform -1 0 3220 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1134_
timestamp 0
transform 1 0 12696 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1135_
timestamp 0
transform -1 0 16744 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1136_
timestamp 0
transform 1 0 9660 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1137_
timestamp 0
transform -1 0 7452 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1138_
timestamp 0
transform -1 0 26312 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1139_
timestamp 0
transform 1 0 27968 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1140_
timestamp 0
transform 1 0 11316 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1141_
timestamp 0
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1142_
timestamp 0
transform -1 0 11500 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1143_
timestamp 0
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a32oi_1  _1144_
timestamp 0
transform 1 0 11316 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1145_
timestamp 0
transform -1 0 13984 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 0
transform 1 0 18308 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1147_
timestamp 0
transform -1 0 27692 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1148_
timestamp 0
transform 1 0 13708 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1149_
timestamp 0
transform 1 0 12972 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1150_
timestamp 0
transform 1 0 12972 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1151_
timestamp 0
transform 1 0 17204 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1152_
timestamp 0
transform 1 0 17480 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1153_
timestamp 0
transform 1 0 12696 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1154_
timestamp 0
transform 1 0 28152 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1155_
timestamp 0
transform -1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1156_
timestamp 0
transform 1 0 26588 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1157_
timestamp 0
transform 1 0 19872 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1158_
timestamp 0
transform 1 0 18676 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1159_
timestamp 0
transform -1 0 19872 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1160_
timestamp 0
transform 1 0 11500 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1161_
timestamp 0
transform 1 0 17204 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1162_
timestamp 0
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1163_
timestamp 0
transform -1 0 17296 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1164_
timestamp 0
transform -1 0 17204 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1165_
timestamp 0
transform 1 0 16376 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1166_
timestamp 0
transform 1 0 14260 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1167_
timestamp 0
transform -1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1168_
timestamp 0
transform 1 0 17112 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1169_
timestamp 0
transform 1 0 17020 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1170_
timestamp 0
transform -1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1171_
timestamp 0
transform -1 0 17940 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1172_
timestamp 0
transform -1 0 17112 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1173_
timestamp 0
transform -1 0 17388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1174_
timestamp 0
transform 1 0 16100 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1175_
timestamp 0
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1176_
timestamp 0
transform 1 0 13800 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1177_
timestamp 0
transform -1 0 15640 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1178_
timestamp 0
transform 1 0 12236 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1179_
timestamp 0
transform 1 0 12144 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1180_
timestamp 0
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1181_
timestamp 0
transform -1 0 22356 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1182_
timestamp 0
transform 1 0 12144 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1183_
timestamp 0
transform 1 0 26128 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1184_
timestamp 0
transform -1 0 25668 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1185_
timestamp 0
transform 1 0 24564 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1186_
timestamp 0
transform 1 0 11500 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1187_
timestamp 0
transform 1 0 11684 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1188_
timestamp 0
transform 1 0 6900 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1189_
timestamp 0
transform -1 0 7452 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1190_
timestamp 0
transform 1 0 6440 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1191_
timestamp 0
transform -1 0 7728 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1192_
timestamp 0
transform 1 0 8280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1193_
timestamp 0
transform -1 0 9200 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1194_
timestamp 0
transform -1 0 9108 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1195_
timestamp 0
transform 1 0 18860 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1196_
timestamp 0
transform 1 0 16284 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 0
transform 1 0 11592 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1198_
timestamp 0
transform 1 0 11592 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1199_
timestamp 0
transform -1 0 21344 0 1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1200_
timestamp 0
transform 1 0 11500 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1201_
timestamp 0
transform -1 0 10028 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1202_
timestamp 0
transform 1 0 9752 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1203_
timestamp 0
transform -1 0 11684 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1204_
timestamp 0
transform 1 0 11040 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1205_
timestamp 0
transform -1 0 8188 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1206_
timestamp 0
transform 1 0 10120 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1207_
timestamp 0
transform -1 0 9844 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1208_
timestamp 0
transform -1 0 16652 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1209_
timestamp 0
transform 1 0 16928 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1210_
timestamp 0
transform -1 0 16928 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1211_
timestamp 0
transform 1 0 14628 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 0
transform -1 0 21160 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1213_
timestamp 0
transform 1 0 16284 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1214_
timestamp 0
transform 1 0 15824 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1215_
timestamp 0
transform -1 0 7084 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1216_
timestamp 0
transform -1 0 8924 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1217_
timestamp 0
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1218_
timestamp 0
transform -1 0 10396 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1219_
timestamp 0
transform 1 0 9108 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 0
transform -1 0 9476 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1221_
timestamp 0
transform -1 0 25116 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_2  _1222_
timestamp 0
transform 1 0 24472 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1223_
timestamp 0
transform 1 0 28888 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1224_
timestamp 0
transform 1 0 27600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1225_
timestamp 0
transform -1 0 16560 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1226_
timestamp 0
transform 1 0 15272 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1227_
timestamp 0
transform -1 0 31372 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1228_
timestamp 0
transform 1 0 29900 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1229_
timestamp 0
transform 1 0 22356 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1230_
timestamp 0
transform 1 0 29808 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1231_
timestamp 0
transform 1 0 29348 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1232_
timestamp 0
transform 1 0 29256 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 0
transform 1 0 18308 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1234_
timestamp 0
transform 1 0 18860 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1235_
timestamp 0
transform 1 0 25760 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1236_
timestamp 0
transform -1 0 26956 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1237_
timestamp 0
transform -1 0 26312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1238_
timestamp 0
transform 1 0 26404 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 0
transform -1 0 24840 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1240_
timestamp 0
transform -1 0 26128 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1241_
timestamp 0
transform -1 0 21712 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1242_
timestamp 0
transform -1 0 20516 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1243_
timestamp 0
transform -1 0 21252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1244_
timestamp 0
transform 1 0 21712 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1245_
timestamp 0
transform 1 0 22356 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1246_
timestamp 0
transform 1 0 22724 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1247_
timestamp 0
transform 1 0 22356 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1248_
timestamp 0
transform -1 0 19872 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1249_
timestamp 0
transform 1 0 19504 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1250_
timestamp 0
transform 1 0 19872 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1251_
timestamp 0
transform -1 0 22908 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1252_
timestamp 0
transform -1 0 16560 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1253_
timestamp 0
transform -1 0 16008 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1254_
timestamp 0
transform -1 0 16008 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_2  _1255_
timestamp 0
transform 1 0 13800 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1256_
timestamp 0
transform -1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1257_
timestamp 0
transform 1 0 18492 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 0
transform 1 0 18676 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1259_
timestamp 0
transform 1 0 6440 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1260_
timestamp 0
transform 1 0 8648 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1261_
timestamp 0
transform 1 0 8556 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1262_
timestamp 0
transform 1 0 7544 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1263_
timestamp 0
transform -1 0 7544 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1264_
timestamp 0
transform -1 0 14444 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1265_
timestamp 0
transform 1 0 15088 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1266_
timestamp 0
transform 1 0 15180 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1267_
timestamp 0
transform 1 0 19504 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1268_
timestamp 0
transform 1 0 15364 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1269_
timestamp 0
transform 1 0 24932 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1270_
timestamp 0
transform 1 0 24288 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1271_
timestamp 0
transform 1 0 14444 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1272_
timestamp 0
transform -1 0 14444 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1273_
timestamp 0
transform 1 0 17388 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1274_
timestamp 0
transform 1 0 16100 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1275_
timestamp 0
transform 1 0 14996 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1276_
timestamp 0
transform 1 0 13892 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1277_
timestamp 0
transform 1 0 14444 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1278_
timestamp 0
transform 1 0 13892 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1279_
timestamp 0
transform -1 0 28796 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1280_
timestamp 0
transform -1 0 28888 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1281_
timestamp 0
transform -1 0 29716 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1282_
timestamp 0
transform -1 0 29256 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1283_
timestamp 0
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_2  _1284_
timestamp 0
transform -1 0 21528 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1285_
timestamp 0
transform -1 0 27416 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1286_
timestamp 0
transform -1 0 26128 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1287_
timestamp 0
transform -1 0 24012 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1288_
timestamp 0
transform -1 0 25484 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1289_
timestamp 0
transform -1 0 25024 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1290_
timestamp 0
transform -1 0 25392 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1291_
timestamp 0
transform -1 0 19412 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1292_
timestamp 0
transform 1 0 20700 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1293_
timestamp 0
transform -1 0 25668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1294_
timestamp 0
transform -1 0 25760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1295_
timestamp 0
transform -1 0 25760 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1296_
timestamp 0
transform 1 0 24932 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1297_
timestamp 0
transform 1 0 24104 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1298_
timestamp 0
transform -1 0 20240 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1299_
timestamp 0
transform -1 0 22172 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1300_
timestamp 0
transform 1 0 21804 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1301_
timestamp 0
transform 1 0 22356 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1302_
timestamp 0
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1303_
timestamp 0
transform -1 0 20792 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1304_
timestamp 0
transform 1 0 23828 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_1  _1305_
timestamp 0
transform -1 0 25668 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1306_
timestamp 0
transform 1 0 23644 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1307_
timestamp 0
transform 1 0 23000 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1308_
timestamp 0
transform 1 0 30360 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1309_
timestamp 0
transform -1 0 30360 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1310_
timestamp 0
transform -1 0 23000 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1311_
timestamp 0
transform 1 0 22724 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1312_
timestamp 0
transform -1 0 22724 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1313_
timestamp 0
transform -1 0 22724 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1314_
timestamp 0
transform 1 0 23276 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1315_
timestamp 0
transform 1 0 22724 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1316_
timestamp 0
transform 1 0 22356 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1317_
timestamp 0
transform 1 0 13064 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1318_
timestamp 0
transform 1 0 21712 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1319_
timestamp 0
transform -1 0 27508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1320_
timestamp 0
transform -1 0 27876 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1321_
timestamp 0
transform 1 0 21896 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1322_
timestamp 0
transform 1 0 21988 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1323_
timestamp 0
transform 1 0 25668 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1324_
timestamp 0
transform 1 0 25668 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1325_
timestamp 0
transform -1 0 26588 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1326_
timestamp 0
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _1327_
timestamp 0
transform -1 0 19780 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1328_
timestamp 0
transform 1 0 28980 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1329_
timestamp 0
transform 1 0 28060 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1330_
timestamp 0
transform 1 0 25576 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1331_
timestamp 0
transform 1 0 21620 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1332_
timestamp 0
transform -1 0 21160 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1333_
timestamp 0
transform -1 0 21528 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 0
transform -1 0 22264 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1335_
timestamp 0
transform 1 0 18032 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1336_
timestamp 0
transform -1 0 19504 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1337_
timestamp 0
transform 1 0 21344 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1338_
timestamp 0
transform 1 0 20424 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1339_
timestamp 0
transform -1 0 22356 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1340_
timestamp 0
transform -1 0 21804 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1341_
timestamp 0
transform -1 0 20700 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1342_
timestamp 0
transform 1 0 24012 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 0
transform 1 0 23276 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1344_
timestamp 0
transform 1 0 23828 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1345_
timestamp 0
transform -1 0 21804 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1346_
timestamp 0
transform 1 0 21252 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1347_
timestamp 0
transform 1 0 21252 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1348_
timestamp 0
transform 1 0 1564 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1349_
timestamp 0
transform 1 0 3220 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1350_
timestamp 0
transform -1 0 26588 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1351_
timestamp 0
transform 1 0 9936 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1352_
timestamp 0
transform -1 0 4968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1353_
timestamp 0
transform 1 0 1564 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1354_
timestamp 0
transform 1 0 1012 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1355_
timestamp 0
transform 1 0 1288 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1356_
timestamp 0
transform 1 0 3220 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 0
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1358_
timestamp 0
transform 1 0 14720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1359_
timestamp 0
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1360_
timestamp 0
transform 1 0 8832 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1361_
timestamp 0
transform 1 0 26220 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1362_
timestamp 0
transform 1 0 26588 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1363_
timestamp 0
transform 1 0 26404 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 0
transform -1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1365_
timestamp 0
transform 1 0 23092 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1366_
timestamp 0
transform 1 0 23000 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1367_
timestamp 0
transform 1 0 22816 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1368_
timestamp 0
transform 1 0 22356 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1369_
timestamp 0
transform -1 0 8832 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1370_
timestamp 0
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1371_
timestamp 0
transform -1 0 14904 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1372_
timestamp 0
transform 1 0 14812 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1373_
timestamp 0
transform 1 0 14996 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1374_
timestamp 0
transform 1 0 14352 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _1375_
timestamp 0
transform 1 0 13616 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__o41a_1  _1376_
timestamp 0
transform -1 0 14076 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1377_
timestamp 0
transform 1 0 13892 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1378_
timestamp 0
transform -1 0 6808 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1379_
timestamp 0
transform 1 0 6808 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1380_
timestamp 0
transform -1 0 5520 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1381_
timestamp 0
transform 1 0 2576 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1382_
timestamp 0
transform 1 0 3404 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1383_
timestamp 0
transform -1 0 4416 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1384_
timestamp 0
transform -1 0 23368 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1385_
timestamp 0
transform -1 0 22816 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _1386_
timestamp 0
transform -1 0 23460 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1387_
timestamp 0
transform 1 0 9752 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1388_
timestamp 0
transform 1 0 4784 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1389_
timestamp 0
transform 1 0 13340 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1390_
timestamp 0
transform 1 0 13064 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1391_
timestamp 0
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1392_
timestamp 0
transform 1 0 13064 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1393_
timestamp 0
transform -1 0 17940 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1394_
timestamp 0
transform 1 0 16744 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1395_
timestamp 0
transform 1 0 17848 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1396_
timestamp 0
transform 1 0 16652 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1397_
timestamp 0
transform 1 0 2300 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1398_
timestamp 0
transform -1 0 17848 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1399_
timestamp 0
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1400_
timestamp 0
transform -1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 0
transform -1 0 16008 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1402_
timestamp 0
transform 1 0 15364 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1403_
timestamp 0
transform -1 0 16928 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1404_
timestamp 0
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1405_
timestamp 0
transform -1 0 18676 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1406_
timestamp 0
transform 1 0 13064 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1407_
timestamp 0
transform 1 0 12420 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1408_
timestamp 0
transform 1 0 1840 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1409_
timestamp 0
transform -1 0 3956 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1410_
timestamp 0
transform 1 0 2760 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1411_
timestamp 0
transform -1 0 24288 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1412_
timestamp 0
transform 1 0 7176 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1413_
timestamp 0
transform -1 0 6716 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _1414_
timestamp 0
transform 1 0 6256 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1415_
timestamp 0
transform 1 0 6624 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1416_
timestamp 0
transform 1 0 9016 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1417_
timestamp 0
transform -1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1418_
timestamp 0
transform -1 0 6072 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1419_
timestamp 0
transform 1 0 6072 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1420_
timestamp 0
transform -1 0 8464 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1421_
timestamp 0
transform 1 0 6532 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1422_
timestamp 0
transform -1 0 6348 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1423_
timestamp 0
transform 1 0 6532 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1424_
timestamp 0
transform 1 0 7820 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1425_
timestamp 0
transform 1 0 828 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1426_
timestamp 0
transform -1 0 2116 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1427_
timestamp 0
transform -1 0 7360 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 0
transform -1 0 4324 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1429_
timestamp 0
transform -1 0 4048 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1430_
timestamp 0
transform 1 0 5520 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1431_
timestamp 0
transform 1 0 13524 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1432_
timestamp 0
transform 1 0 13248 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1433_
timestamp 0
transform -1 0 24748 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1434_
timestamp 0
transform -1 0 15088 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1435_
timestamp 0
transform -1 0 28428 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1436_
timestamp 0
transform -1 0 27232 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1437_
timestamp 0
transform 1 0 24288 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or4bb_1  _1438_
timestamp 0
transform 1 0 13708 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1439_
timestamp 0
transform -1 0 6716 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1440_
timestamp 0
transform 1 0 5888 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1441_
timestamp 0
transform 1 0 9936 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1442_
timestamp 0
transform -1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1443_
timestamp 0
transform 1 0 4416 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1444_
timestamp 0
transform 1 0 9292 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1445_
timestamp 0
transform 1 0 3864 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a41oi_2  _1446_
timestamp 0
transform -1 0 6808 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _1447_
timestamp 0
transform -1 0 12880 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1448_
timestamp 0
transform 1 0 11960 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1449_
timestamp 0
transform -1 0 8280 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1450_
timestamp 0
transform 1 0 7360 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1451_
timestamp 0
transform -1 0 8004 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1452_
timestamp 0
transform 1 0 8648 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _1453_
timestamp 0
transform -1 0 9200 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1454_
timestamp 0
transform -1 0 9844 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1455_
timestamp 0
transform -1 0 9108 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1456_
timestamp 0
transform 1 0 15088 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1457_
timestamp 0
transform 1 0 12052 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1458_
timestamp 0
transform -1 0 9568 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 0
transform 1 0 29440 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1460_
timestamp 0
transform -1 0 28704 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1461_
timestamp 0
transform 1 0 26956 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1462_
timestamp 0
transform -1 0 27876 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1463_
timestamp 0
transform 1 0 12604 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1464_
timestamp 0
transform 1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1465_
timestamp 0
transform -1 0 10212 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1466_
timestamp 0
transform -1 0 10764 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1467_
timestamp 0
transform -1 0 8280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1468_
timestamp 0
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _1469_
timestamp 0
transform 1 0 10212 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1470_
timestamp 0
transform 1 0 10948 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1471_
timestamp 0
transform 1 0 10212 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1472_
timestamp 0
transform 1 0 10028 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1473_
timestamp 0
transform -1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1474_
timestamp 0
transform 1 0 12328 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1475_
timestamp 0
transform 1 0 11592 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1476_
timestamp 0
transform 1 0 11500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1477_
timestamp 0
transform -1 0 10580 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1478_
timestamp 0
transform 1 0 7912 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1479_
timestamp 0
transform -1 0 9476 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1480_
timestamp 0
transform 1 0 8556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1481_
timestamp 0
transform 1 0 8924 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_1  _1482_
timestamp 0
transform 1 0 10028 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1483_
timestamp 0
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1484_
timestamp 0
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1485_
timestamp 0
transform -1 0 15364 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1486_
timestamp 0
transform 1 0 14444 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1487_
timestamp 0
transform 1 0 11132 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1488_
timestamp 0
transform 1 0 11316 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _1489_
timestamp 0
transform 1 0 11500 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_1  _1490_
timestamp 0
transform 1 0 11960 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1491_
timestamp 0
transform 1 0 12604 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1492_
timestamp 0
transform -1 0 14260 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1493_
timestamp 0
transform -1 0 14352 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1494_
timestamp 0
transform -1 0 28888 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1495_
timestamp 0
transform 1 0 25944 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1496_
timestamp 0
transform 1 0 23092 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1497_
timestamp 0
transform 1 0 23368 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _1498_
timestamp 0
transform 1 0 23828 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 0
transform -1 0 26864 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 0
transform -1 0 31280 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1501_
timestamp 0
transform -1 0 28152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1502_
timestamp 0
transform 1 0 27140 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1503_
timestamp 0
transform 1 0 30452 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1504_
timestamp 0
transform -1 0 29808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1505_
timestamp 0
transform -1 0 29624 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1506_
timestamp 0
transform 1 0 29808 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1507_
timestamp 0
transform 1 0 28244 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1508_
timestamp 0
transform -1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1509_
timestamp 0
transform 1 0 29624 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1510_
timestamp 0
transform -1 0 31188 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 0
transform 1 0 25116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1512_
timestamp 0
transform 1 0 29348 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1513_
timestamp 0
transform -1 0 31280 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1514_
timestamp 0
transform -1 0 24104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1515_
timestamp 0
transform 1 0 30820 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1516_
timestamp 0
transform 1 0 28612 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1517_
timestamp 0
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1518_
timestamp 0
transform -1 0 29808 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1519_
timestamp 0
transform 1 0 27140 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1520_
timestamp 0
transform -1 0 31372 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1521_
timestamp 0
transform 1 0 25392 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1522_
timestamp 0
transform -1 0 23920 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 0
transform -1 0 24748 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1524_
timestamp 0
transform 1 0 17940 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1525_
timestamp 0
transform -1 0 19412 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1526_
timestamp 0
transform 1 0 18860 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1527_
timestamp 0
transform 1 0 18860 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1528_
timestamp 0
transform 1 0 18400 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1529_
timestamp 0
transform 1 0 19780 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp 0
transform -1 0 20792 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1531_
timestamp 0
transform -1 0 25116 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1532_
timestamp 0
transform 1 0 24932 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1533_
timestamp 0
transform 1 0 31096 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 0
transform -1 0 26220 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _1535_
timestamp 0
transform 1 0 19504 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1536_
timestamp 0
transform -1 0 28704 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1537_
timestamp 0
transform 1 0 24932 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 0
transform 1 0 25668 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 0
transform -1 0 29624 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1540_
timestamp 0
transform 1 0 27692 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1541_
timestamp 0
transform -1 0 31372 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1542_
timestamp 0
transform 1 0 31096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1543_
timestamp 0
transform -1 0 28796 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1544_
timestamp 0
transform 1 0 28704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 0
transform 1 0 27692 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1546_
timestamp 0
transform -1 0 21436 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1547_
timestamp 0
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1548_
timestamp 0
transform -1 0 23552 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1549_
timestamp 0
transform 1 0 22356 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1550_
timestamp 0
transform -1 0 21160 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1551_
timestamp 0
transform -1 0 21160 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1552_
timestamp 0
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1553_
timestamp 0
transform -1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1554_
timestamp 0
transform 1 0 23828 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1555_
timestamp 0
transform -1 0 27140 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1556_
timestamp 0
transform 1 0 22264 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1557_
timestamp 0
transform -1 0 20424 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1558_
timestamp 0
transform 1 0 17020 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1559_
timestamp 0
transform -1 0 16836 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1560_
timestamp 0
transform -1 0 21712 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1561_
timestamp 0
transform 1 0 17112 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1562_
timestamp 0
transform -1 0 16560 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 0
transform 1 0 15180 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1564_
timestamp 0
transform 1 0 17020 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1565_
timestamp 0
transform 1 0 15548 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1566_
timestamp 0
transform -1 0 17940 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1567_
timestamp 0
transform 1 0 15548 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1568_
timestamp 0
transform 1 0 16284 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1569_
timestamp 0
transform 1 0 16100 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1570_
timestamp 0
transform 1 0 18860 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1571_
timestamp 0
transform 1 0 20792 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1572_
timestamp 0
transform -1 0 21252 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1573_
timestamp 0
transform -1 0 20056 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _1574_
timestamp 0
transform 1 0 23552 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1575_
timestamp 0
transform 1 0 16376 0 1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1576_
timestamp 0
transform 1 0 26404 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1577_
timestamp 0
transform 1 0 26956 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1578_
timestamp 0
transform 1 0 28980 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1579_
timestamp 0
transform 1 0 28980 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1580_
timestamp 0
transform 1 0 28980 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1581_
timestamp 0
transform 1 0 26404 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1582_
timestamp 0
transform 1 0 23920 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1583_
timestamp 0
transform 1 0 24104 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1584_
timestamp 0
transform 1 0 21528 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1585_
timestamp 0
transform -1 0 23552 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1586_
timestamp 0
transform 1 0 21252 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1587_
timestamp 0
transform 1 0 18676 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1588_
timestamp 0
transform -1 0 28244 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1589_
timestamp 0
transform 1 0 24288 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1590_
timestamp 0
transform -1 0 27140 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1591_
timestamp 0
transform 1 0 29348 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1592_
timestamp 0
transform -1 0 30084 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1593_
timestamp 0
transform 1 0 28980 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1594_
timestamp 0
transform 1 0 23092 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1595_
timestamp 0
transform -1 0 23092 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1596_
timestamp 0
transform -1 0 24932 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1597_
timestamp 0
transform -1 0 23736 0 1 19040
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1598_
timestamp 0
transform 1 0 16836 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1599_
timestamp 0
transform 1 0 14628 0 1 17952
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1600_
timestamp 0
transform 1 0 16468 0 1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1601_
timestamp 0
transform -1 0 16468 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1602_
timestamp 0
transform -1 0 22080 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1603_
timestamp 0
transform 1 0 19320 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1604_
timestamp 0
transform 1 0 7912 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1605_
timestamp 0
transform 1 0 7176 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1606_
timestamp 0
transform 1 0 11500 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1607_
timestamp 0
transform 1 0 9016 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1608_
timestamp 0
transform 1 0 13984 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 26864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 0
transform 1 0 15088 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 0
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 0
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 0
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 0
transform -1 0 11684 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 0
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 0
transform -1 0 9844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 0
transform -1 0 11408 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 0
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 0
transform -1 0 12880 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 0
transform -1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 20516 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 13432 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform -1 0 18676 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform 1 0 26404 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform -1 0 26312 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinvlp_4  clkload0
timestamp 0
transform 1 0 11040 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp 0
transform 1 0 15180 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 0
transform 1 0 24748 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout4
timestamp 0
transform -1 0 4232 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout5
timestamp 0
transform -1 0 6164 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout6
timestamp 0
transform -1 0 3772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 0
transform 1 0 28336 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 0
transform -1 0 27968 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 0
transform 1 0 27600 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 0
transform 1 0 12236 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 0
transform -1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 0
transform 1 0 15456 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 0
transform -1 0 24932 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout20
timestamp 0
transform 1 0 24748 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 0
transform 1 0 2300 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout22
timestamp 0
transform 1 0 25668 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 0
transform -1 0 17848 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 0
transform 1 0 27232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 0
transform -1 0 7912 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 0
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout27
timestamp 0
transform 1 0 7452 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 0
transform -1 0 13064 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 0
transform 1 0 28520 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 0
transform -1 0 29624 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 0
transform 1 0 13064 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 0
transform -1 0 30728 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 0
transform -1 0 30912 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 0
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 0
transform 1 0 6072 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 0
transform -1 0 18216 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 0
transform 1 0 9384 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 0
transform 1 0 21252 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 0
transform 1 0 20608 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 0
transform 1 0 8556 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 0
transform -1 0 14628 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 0
transform -1 0 26680 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 0
transform -1 0 27692 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 0
transform -1 0 16008 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 0
transform -1 0 24656 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 0
transform -1 0 24288 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 0
transform -1 0 21988 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 0
transform -1 0 22540 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 0
transform 1 0 14904 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 0
transform 1 0 14168 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 0
transform -1 0 8280 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 0
transform -1 0 13156 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 0
transform 1 0 26680 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 0
transform 1 0 24840 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 0
transform -1 0 23736 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 0
transform 1 0 23368 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 0
transform -1 0 24196 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 0
transform 1 0 6072 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 0
transform -1 0 3588 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 0
transform -1 0 7728 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp 0
transform -1 0 10764 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp 0
transform -1 0 15548 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 0
transform -1 0 10212 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 0
transform 1 0 18952 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 0
transform -1 0 24288 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout66
timestamp 0
transform 1 0 30820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 0
transform 1 0 30728 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 0
transform -1 0 30176 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout69
timestamp 0
transform -1 0 9844 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 0
transform 1 0 14720 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 0
transform -1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 0
transform -1 0 8556 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 0
transform -1 0 16008 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout74
timestamp 0
transform -1 0 30636 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 0
transform 1 0 30544 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 0
transform -1 0 29532 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout77
timestamp 0
transform -1 0 29348 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 0
transform 1 0 30912 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 0
transform -1 0 28060 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout80
timestamp 0
transform -1 0 7084 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout81
timestamp 0
transform 1 0 7544 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 0
transform -1 0 7084 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 0
transform -1 0 13892 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 0
transform -1 0 22724 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout85
timestamp 0
transform -1 0 22356 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout86
timestamp 0
transform -1 0 27416 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout87
timestamp 0
transform -1 0 30084 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout88
timestamp 0
transform -1 0 29532 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout89
timestamp 0
transform -1 0 30636 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout90
timestamp 0
transform 1 0 30636 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 0
transform -1 0 30544 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout92
timestamp 0
transform 1 0 6256 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout93
timestamp 0
transform -1 0 3680 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout94
timestamp 0
transform 1 0 12880 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout95
timestamp 0
transform 1 0 27508 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout96
timestamp 0
transform 1 0 28612 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 0
transform -1 0 28520 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout98
timestamp 0
transform 1 0 28336 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 0
transform -1 0 29348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout100
timestamp 0
transform 1 0 30176 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout101
timestamp 0
transform 1 0 5980 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 0
transform -1 0 2392 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout103
timestamp 0
transform -1 0 14260 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout104
timestamp 0
transform 1 0 28704 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout105
timestamp 0
transform -1 0 24472 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout106
timestamp 0
transform -1 0 27692 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 0
transform 1 0 26404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 0
transform 1 0 28060 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout109
timestamp 0
transform -1 0 2116 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 0
transform -1 0 13432 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout111
timestamp 0
transform 1 0 25576 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 0
transform -1 0 29072 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout113
timestamp 0
transform 1 0 28980 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout114
timestamp 0
transform -1 0 21988 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 0
transform 1 0 30820 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout116
timestamp 0
transform -1 0 29072 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout117
timestamp 0
transform -1 0 26312 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout118
timestamp 0
transform 1 0 30820 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp 0
transform 1 0 30728 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout120
timestamp 0
transform -1 0 19228 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_3
timestamp 0
transform 1 0 828 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_6
timestamp 0
transform 1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_9
timestamp 0
transform 1 0 1380 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_12
timestamp 0
transform 1 0 1656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_15
timestamp 0
transform 1 0 1932 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_18
timestamp 0
transform 1 0 2208 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_21
timestamp 0
transform 1 0 2484 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_24
timestamp 0
transform 1 0 2760 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29
timestamp 0
transform 1 0 3220 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_32
timestamp 0
transform 1 0 3496 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_35
timestamp 0
transform 1 0 3772 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_38
timestamp 0
transform 1 0 4048 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_41
timestamp 0
transform 1 0 4324 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_44
timestamp 0
transform 1 0 4600 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_47
timestamp 0
transform 1 0 4876 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_50
timestamp 0
transform 1 0 5152 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57
timestamp 0
transform 1 0 5796 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_60
timestamp 0
transform 1 0 6072 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63
timestamp 0
transform 1 0 6348 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_66
timestamp 0
transform 1 0 6624 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69
timestamp 0
transform 1 0 6900 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_72
timestamp 0
transform 1 0 7176 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_75
timestamp 0
transform 1 0 7452 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_78
timestamp 0
transform 1 0 7728 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_85
timestamp 0
transform 1 0 8372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_88
timestamp 0
transform 1 0 8648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_91
timestamp 0
transform 1 0 8924 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_94
timestamp 0
transform 1 0 9200 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_97
timestamp 0
transform 1 0 9476 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_100
timestamp 0
transform 1 0 9752 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_103
timestamp 0
transform 1 0 10028 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_106
timestamp 0
transform 1 0 10304 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 0
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_116
timestamp 0
transform 1 0 11224 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_119
timestamp 0
transform 1 0 11500 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_122
timestamp 0
transform 1 0 11776 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_125
timestamp 0
transform 1 0 12052 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_128
timestamp 0
transform 1 0 12328 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_131
timestamp 0
transform 1 0 12604 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_134
timestamp 0
transform 1 0 12880 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_141
timestamp 0
transform 1 0 13524 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_144
timestamp 0
transform 1 0 13800 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_147
timestamp 0
transform 1 0 14076 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_150
timestamp 0
transform 1 0 14352 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_153
timestamp 0
transform 1 0 14628 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_156
timestamp 0
transform 1 0 14904 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_159
timestamp 0
transform 1 0 15180 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_162
timestamp 0
transform 1 0 15456 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_169
timestamp 0
transform 1 0 16100 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_172
timestamp 0
transform 1 0 16376 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_175
timestamp 0
transform 1 0 16652 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_178
timestamp 0
transform 1 0 16928 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_181
timestamp 0
transform 1 0 17204 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_184
timestamp 0
transform 1 0 17480 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_187
timestamp 0
transform 1 0 17756 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_190
timestamp 0
transform 1 0 18032 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 0
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_197
timestamp 0
transform 1 0 18676 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_200
timestamp 0
transform 1 0 18952 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_203
timestamp 0
transform 1 0 19228 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_206
timestamp 0
transform 1 0 19504 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_209
timestamp 0
transform 1 0 19780 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_212
timestamp 0
transform 1 0 20056 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_215
timestamp 0
transform 1 0 20332 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_218
timestamp 0
transform 1 0 20608 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 0
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_228
timestamp 0
transform 1 0 21528 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_231
timestamp 0
transform 1 0 21804 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_234
timestamp 0
transform 1 0 22080 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_237
timestamp 0
transform 1 0 22356 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_240
timestamp 0
transform 1 0 22632 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_243
timestamp 0
transform 1 0 22908 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_246
timestamp 0
transform 1 0 23184 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 0
transform 1 0 23828 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_256
timestamp 0
transform 1 0 24104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_259
timestamp 0
transform 1 0 24380 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_262
timestamp 0
transform 1 0 24656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_265
timestamp 0
transform 1 0 24932 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_268
timestamp 0
transform 1 0 25208 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_271
timestamp 0
transform 1 0 25484 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_274
timestamp 0
transform 1 0 25760 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 0
transform 1 0 26404 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_284
timestamp 0
transform 1 0 26680 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_287
timestamp 0
transform 1 0 26956 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_290
timestamp 0
transform 1 0 27232 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_293
timestamp 0
transform 1 0 27508 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_296
timestamp 0
transform 1 0 27784 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_299
timestamp 0
transform 1 0 28060 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_302
timestamp 0
transform 1 0 28336 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 0
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_309
timestamp 0
transform 1 0 28980 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_312
timestamp 0
transform 1 0 29256 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_315
timestamp 0
transform 1 0 29532 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_318
timestamp 0
transform 1 0 29808 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_321
timestamp 0
transform 1 0 30084 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_324
timestamp 0
transform 1 0 30360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_327
timestamp 0
transform 1 0 30636 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_330
timestamp 0
transform 1 0 30912 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 0
transform 1 0 31188 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_3
timestamp 0
transform 1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_6
timestamp 0
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_9
timestamp 0
transform 1 0 1380 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_12
timestamp 0
transform 1 0 1656 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_15
timestamp 0
transform 1 0 1932 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_18
timestamp 0
transform 1 0 2208 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_21
timestamp 0
transform 1 0 2484 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_24
timestamp 0
transform 1 0 2760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_27
timestamp 0
transform 1 0 3036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_30
timestamp 0
transform 1 0 3312 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_33
timestamp 0
transform 1 0 3588 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_36
timestamp 0
transform 1 0 3864 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_39
timestamp 0
transform 1 0 4140 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_42
timestamp 0
transform 1 0 4416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_45
timestamp 0
transform 1 0 4692 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_48
timestamp 0
transform 1 0 4968 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_51
timestamp 0
transform 1 0 5244 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 0
transform 1 0 5520 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 0
transform 1 0 5796 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_60
timestamp 0
transform 1 0 6072 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_63
timestamp 0
transform 1 0 6348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_66
timestamp 0
transform 1 0 6624 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_69
timestamp 0
transform 1 0 6900 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_72
timestamp 0
transform 1 0 7176 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_75
timestamp 0
transform 1 0 7452 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_78
timestamp 0
transform 1 0 7728 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_81
timestamp 0
transform 1 0 8004 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_84
timestamp 0
transform 1 0 8280 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_87
timestamp 0
transform 1 0 8556 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_90
timestamp 0
transform 1 0 8832 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_93
timestamp 0
transform 1 0 9108 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_96
timestamp 0
transform 1 0 9384 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_99
timestamp 0
transform 1 0 9660 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_102
timestamp 0
transform 1 0 9936 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_105
timestamp 0
transform 1 0 10212 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_108
timestamp 0
transform 1 0 10488 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_113
timestamp 0
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_116
timestamp 0
transform 1 0 11224 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_119
timestamp 0
transform 1 0 11500 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_122
timestamp 0
transform 1 0 11776 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_125
timestamp 0
transform 1 0 12052 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_128
timestamp 0
transform 1 0 12328 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_131
timestamp 0
transform 1 0 12604 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_134
timestamp 0
transform 1 0 12880 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_137
timestamp 0
transform 1 0 13156 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_140
timestamp 0
transform 1 0 13432 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_143
timestamp 0
transform 1 0 13708 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_146
timestamp 0
transform 1 0 13984 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_149
timestamp 0
transform 1 0 14260 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_152
timestamp 0
transform 1 0 14536 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_155
timestamp 0
transform 1 0 14812 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_158
timestamp 0
transform 1 0 15088 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_161
timestamp 0
transform 1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_164
timestamp 0
transform 1 0 15640 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_169
timestamp 0
transform 1 0 16100 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_172
timestamp 0
transform 1 0 16376 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_175
timestamp 0
transform 1 0 16652 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_178
timestamp 0
transform 1 0 16928 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_181
timestamp 0
transform 1 0 17204 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_184
timestamp 0
transform 1 0 17480 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_187
timestamp 0
transform 1 0 17756 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_190
timestamp 0
transform 1 0 18032 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_193
timestamp 0
transform 1 0 18308 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_196
timestamp 0
transform 1 0 18584 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_199
timestamp 0
transform 1 0 18860 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_202
timestamp 0
transform 1 0 19136 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_205
timestamp 0
transform 1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_208
timestamp 0
transform 1 0 19688 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_211
timestamp 0
transform 1 0 19964 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_214
timestamp 0
transform 1 0 20240 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_217
timestamp 0
transform 1 0 20516 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_220
timestamp 0
transform 1 0 20792 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 0
transform 1 0 21252 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_228
timestamp 0
transform 1 0 21528 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_231
timestamp 0
transform 1 0 21804 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_234
timestamp 0
transform 1 0 22080 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_237
timestamp 0
transform 1 0 22356 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_240
timestamp 0
transform 1 0 22632 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_243
timestamp 0
transform 1 0 22908 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_246
timestamp 0
transform 1 0 23184 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_249
timestamp 0
transform 1 0 23460 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_252
timestamp 0
transform 1 0 23736 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_255
timestamp 0
transform 1 0 24012 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_258
timestamp 0
transform 1 0 24288 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_261
timestamp 0
transform 1 0 24564 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_264
timestamp 0
transform 1 0 24840 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_267
timestamp 0
transform 1 0 25116 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_270
timestamp 0
transform 1 0 25392 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_273
timestamp 0
transform 1 0 25668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_276
timestamp 0
transform 1 0 25944 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_281
timestamp 0
transform 1 0 26404 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_284
timestamp 0
transform 1 0 26680 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_287
timestamp 0
transform 1 0 26956 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_290
timestamp 0
transform 1 0 27232 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_293
timestamp 0
transform 1 0 27508 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_296
timestamp 0
transform 1 0 27784 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_299
timestamp 0
transform 1 0 28060 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_302
timestamp 0
transform 1 0 28336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_305
timestamp 0
transform 1 0 28612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_308
timestamp 0
transform 1 0 28888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_311
timestamp 0
transform 1 0 29164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_314
timestamp 0
transform 1 0 29440 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_317
timestamp 0
transform 1 0 29716 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_320
timestamp 0
transform 1 0 29992 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_323
timestamp 0
transform 1 0 30268 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_326
timestamp 0
transform 1 0 30544 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_329
timestamp 0
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_332
timestamp 0
transform 1 0 31096 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_3
timestamp 0
transform 1 0 828 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_6
timestamp 0
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_9
timestamp 0
transform 1 0 1380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_12
timestamp 0
transform 1 0 1656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_15
timestamp 0
transform 1 0 1932 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_18
timestamp 0
transform 1 0 2208 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_21
timestamp 0
transform 1 0 2484 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_24
timestamp 0
transform 1 0 2760 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_29
timestamp 0
transform 1 0 3220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_32
timestamp 0
transform 1 0 3496 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_35
timestamp 0
transform 1 0 3772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_38
timestamp 0
transform 1 0 4048 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_41
timestamp 0
transform 1 0 4324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_44
timestamp 0
transform 1 0 4600 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_47
timestamp 0
transform 1 0 4876 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_50
timestamp 0
transform 1 0 5152 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_53
timestamp 0
transform 1 0 5428 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_56
timestamp 0
transform 1 0 5704 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_59
timestamp 0
transform 1 0 5980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_62
timestamp 0
transform 1 0 6256 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_65
timestamp 0
transform 1 0 6532 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_68
timestamp 0
transform 1 0 6808 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_71
timestamp 0
transform 1 0 7084 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_74
timestamp 0
transform 1 0 7360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_77
timestamp 0
transform 1 0 7636 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_80
timestamp 0
transform 1 0 7912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 0
transform 1 0 8372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_88
timestamp 0
transform 1 0 8648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_91
timestamp 0
transform 1 0 8924 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_94
timestamp 0
transform 1 0 9200 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_97
timestamp 0
transform 1 0 9476 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_100
timestamp 0
transform 1 0 9752 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_103
timestamp 0
transform 1 0 10028 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_106
timestamp 0
transform 1 0 10304 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_109
timestamp 0
transform 1 0 10580 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_112
timestamp 0
transform 1 0 10856 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_115
timestamp 0
transform 1 0 11132 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_118
timestamp 0
transform 1 0 11408 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_121
timestamp 0
transform 1 0 11684 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_124
timestamp 0
transform 1 0 11960 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_127
timestamp 0
transform 1 0 12236 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_130
timestamp 0
transform 1 0 12512 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_133
timestamp 0
transform 1 0 12788 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_136
timestamp 0
transform 1 0 13064 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 0
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_144
timestamp 0
transform 1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_147
timestamp 0
transform 1 0 14076 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_150
timestamp 0
transform 1 0 14352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_153
timestamp 0
transform 1 0 14628 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_156
timestamp 0
transform 1 0 14904 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_159
timestamp 0
transform 1 0 15180 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_162
timestamp 0
transform 1 0 15456 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_165
timestamp 0
transform 1 0 15732 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_168
timestamp 0
transform 1 0 16008 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_171
timestamp 0
transform 1 0 16284 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_174
timestamp 0
transform 1 0 16560 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_177
timestamp 0
transform 1 0 16836 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_180
timestamp 0
transform 1 0 17112 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_183
timestamp 0
transform 1 0 17388 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_186
timestamp 0
transform 1 0 17664 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_189
timestamp 0
transform 1 0 17940 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_192
timestamp 0
transform 1 0 18216 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_197
timestamp 0
transform 1 0 18676 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_200
timestamp 0
transform 1 0 18952 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_203
timestamp 0
transform 1 0 19228 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_206
timestamp 0
transform 1 0 19504 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_209
timestamp 0
transform 1 0 19780 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_212
timestamp 0
transform 1 0 20056 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_215
timestamp 0
transform 1 0 20332 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_218
timestamp 0
transform 1 0 20608 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_221
timestamp 0
transform 1 0 20884 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_224
timestamp 0
transform 1 0 21160 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_227
timestamp 0
transform 1 0 21436 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_230
timestamp 0
transform 1 0 21712 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_233
timestamp 0
transform 1 0 21988 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_236
timestamp 0
transform 1 0 22264 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_239
timestamp 0
transform 1 0 22540 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_242
timestamp 0
transform 1 0 22816 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_245
timestamp 0
transform 1 0 23092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_248
timestamp 0
transform 1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 0
transform 1 0 23828 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_256
timestamp 0
transform 1 0 24104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_259
timestamp 0
transform 1 0 24380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_262
timestamp 0
transform 1 0 24656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_265
timestamp 0
transform 1 0 24932 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_268
timestamp 0
transform 1 0 25208 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_271
timestamp 0
transform 1 0 25484 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_274
timestamp 0
transform 1 0 25760 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_277
timestamp 0
transform 1 0 26036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_280
timestamp 0
transform 1 0 26312 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_283
timestamp 0
transform 1 0 26588 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_286
timestamp 0
transform 1 0 26864 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_289
timestamp 0
transform 1 0 27140 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_292
timestamp 0
transform 1 0 27416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_295
timestamp 0
transform 1 0 27692 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_298
timestamp 0
transform 1 0 27968 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_301
timestamp 0
transform 1 0 28244 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_304
timestamp 0
transform 1 0 28520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_309
timestamp 0
transform 1 0 28980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_312
timestamp 0
transform 1 0 29256 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_315
timestamp 0
transform 1 0 29532 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_318
timestamp 0
transform 1 0 29808 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_321
timestamp 0
transform 1 0 30084 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_324
timestamp 0
transform 1 0 30360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_327
timestamp 0
transform 1 0 30636 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_330
timestamp 0
transform 1 0 30912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 0
transform 1 0 31188 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_3
timestamp 0
transform 1 0 828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_6
timestamp 0
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_9
timestamp 0
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_12
timestamp 0
transform 1 0 1656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_15
timestamp 0
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_18
timestamp 0
transform 1 0 2208 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_21
timestamp 0
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_24
timestamp 0
transform 1 0 2760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_27
timestamp 0
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_30
timestamp 0
transform 1 0 3312 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_33
timestamp 0
transform 1 0 3588 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_36
timestamp 0
transform 1 0 3864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_39
timestamp 0
transform 1 0 4140 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_42
timestamp 0
transform 1 0 4416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_45
timestamp 0
transform 1 0 4692 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_48
timestamp 0
transform 1 0 4968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_51
timestamp 0
transform 1 0 5244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 0
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_57
timestamp 0
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_60
timestamp 0
transform 1 0 6072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_63
timestamp 0
transform 1 0 6348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_66
timestamp 0
transform 1 0 6624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_69
timestamp 0
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_72
timestamp 0
transform 1 0 7176 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_75
timestamp 0
transform 1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_78
timestamp 0
transform 1 0 7728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_81
timestamp 0
transform 1 0 8004 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_84
timestamp 0
transform 1 0 8280 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_87
timestamp 0
transform 1 0 8556 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_90
timestamp 0
transform 1 0 8832 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_93
timestamp 0
transform 1 0 9108 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_96
timestamp 0
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_99
timestamp 0
transform 1 0 9660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_102
timestamp 0
transform 1 0 9936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_105
timestamp 0
transform 1 0 10212 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_108
timestamp 0
transform 1 0 10488 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 0
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_116
timestamp 0
transform 1 0 11224 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_119
timestamp 0
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_122
timestamp 0
transform 1 0 11776 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_125
timestamp 0
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_128
timestamp 0
transform 1 0 12328 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_131
timestamp 0
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_134
timestamp 0
transform 1 0 12880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_137
timestamp 0
transform 1 0 13156 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_140
timestamp 0
transform 1 0 13432 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_143
timestamp 0
transform 1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_146
timestamp 0
transform 1 0 13984 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_149
timestamp 0
transform 1 0 14260 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_152
timestamp 0
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_155
timestamp 0
transform 1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_158
timestamp 0
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_161
timestamp 0
transform 1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_164
timestamp 0
transform 1 0 15640 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_169
timestamp 0
transform 1 0 16100 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_172
timestamp 0
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_175
timestamp 0
transform 1 0 16652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_178
timestamp 0
transform 1 0 16928 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_181
timestamp 0
transform 1 0 17204 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_184
timestamp 0
transform 1 0 17480 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_187
timestamp 0
transform 1 0 17756 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_190
timestamp 0
transform 1 0 18032 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_193
timestamp 0
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_196
timestamp 0
transform 1 0 18584 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_199
timestamp 0
transform 1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_202
timestamp 0
transform 1 0 19136 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_205
timestamp 0
transform 1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_208
timestamp 0
transform 1 0 19688 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_211
timestamp 0
transform 1 0 19964 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_214
timestamp 0
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_217
timestamp 0
transform 1 0 20516 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_220
timestamp 0
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_225
timestamp 0
transform 1 0 21252 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_228
timestamp 0
transform 1 0 21528 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_231
timestamp 0
transform 1 0 21804 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_234
timestamp 0
transform 1 0 22080 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_237
timestamp 0
transform 1 0 22356 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_240
timestamp 0
transform 1 0 22632 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_243
timestamp 0
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_246
timestamp 0
transform 1 0 23184 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_249
timestamp 0
transform 1 0 23460 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_252
timestamp 0
transform 1 0 23736 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_255
timestamp 0
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_258
timestamp 0
transform 1 0 24288 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_261
timestamp 0
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_264
timestamp 0
transform 1 0 24840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_267
timestamp 0
transform 1 0 25116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_270
timestamp 0
transform 1 0 25392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_273
timestamp 0
transform 1 0 25668 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_276
timestamp 0
transform 1 0 25944 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_281
timestamp 0
transform 1 0 26404 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_284
timestamp 0
transform 1 0 26680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_287
timestamp 0
transform 1 0 26956 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_290
timestamp 0
transform 1 0 27232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_293
timestamp 0
transform 1 0 27508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_296
timestamp 0
transform 1 0 27784 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_299
timestamp 0
transform 1 0 28060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_302
timestamp 0
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_305
timestamp 0
transform 1 0 28612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_308
timestamp 0
transform 1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_311
timestamp 0
transform 1 0 29164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_314
timestamp 0
transform 1 0 29440 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_317
timestamp 0
transform 1 0 29716 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_320
timestamp 0
transform 1 0 29992 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_323
timestamp 0
transform 1 0 30268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_326
timestamp 0
transform 1 0 30544 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_329
timestamp 0
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_332
timestamp 0
transform 1 0 31096 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_3
timestamp 0
transform 1 0 828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_6
timestamp 0
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_9
timestamp 0
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_12
timestamp 0
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_15
timestamp 0
transform 1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_18
timestamp 0
transform 1 0 2208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_21
timestamp 0
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_24
timestamp 0
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_29
timestamp 0
transform 1 0 3220 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_32
timestamp 0
transform 1 0 3496 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_35
timestamp 0
transform 1 0 3772 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_38
timestamp 0
transform 1 0 4048 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_41
timestamp 0
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_44
timestamp 0
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_47
timestamp 0
transform 1 0 4876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_50
timestamp 0
transform 1 0 5152 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_53
timestamp 0
transform 1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_56
timestamp 0
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_59
timestamp 0
transform 1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_62
timestamp 0
transform 1 0 6256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_65
timestamp 0
transform 1 0 6532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_68
timestamp 0
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_71
timestamp 0
transform 1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_74
timestamp 0
transform 1 0 7360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_77
timestamp 0
transform 1 0 7636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_80
timestamp 0
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 0
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_88
timestamp 0
transform 1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_91
timestamp 0
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_94
timestamp 0
transform 1 0 9200 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_97
timestamp 0
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_100
timestamp 0
transform 1 0 9752 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_103
timestamp 0
transform 1 0 10028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_106
timestamp 0
transform 1 0 10304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_109
timestamp 0
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_112
timestamp 0
transform 1 0 10856 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_115
timestamp 0
transform 1 0 11132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_118
timestamp 0
transform 1 0 11408 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_121
timestamp 0
transform 1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_124
timestamp 0
transform 1 0 11960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_127
timestamp 0
transform 1 0 12236 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_130
timestamp 0
transform 1 0 12512 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_133
timestamp 0
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_136
timestamp 0
transform 1 0 13064 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_141
timestamp 0
transform 1 0 13524 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_144
timestamp 0
transform 1 0 13800 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_147
timestamp 0
transform 1 0 14076 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_150
timestamp 0
transform 1 0 14352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_153
timestamp 0
transform 1 0 14628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_156
timestamp 0
transform 1 0 14904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_159
timestamp 0
transform 1 0 15180 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_162
timestamp 0
transform 1 0 15456 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_165
timestamp 0
transform 1 0 15732 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_168
timestamp 0
transform 1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_171
timestamp 0
transform 1 0 16284 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_174
timestamp 0
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_177
timestamp 0
transform 1 0 16836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_180
timestamp 0
transform 1 0 17112 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_183
timestamp 0
transform 1 0 17388 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_186
timestamp 0
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_189
timestamp 0
transform 1 0 17940 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_192
timestamp 0
transform 1 0 18216 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_197
timestamp 0
transform 1 0 18676 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_200
timestamp 0
transform 1 0 18952 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_203
timestamp 0
transform 1 0 19228 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_206
timestamp 0
transform 1 0 19504 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_209
timestamp 0
transform 1 0 19780 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_212
timestamp 0
transform 1 0 20056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_215
timestamp 0
transform 1 0 20332 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_218
timestamp 0
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_221
timestamp 0
transform 1 0 20884 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_224
timestamp 0
transform 1 0 21160 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_227
timestamp 0
transform 1 0 21436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_230
timestamp 0
transform 1 0 21712 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_233
timestamp 0
transform 1 0 21988 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_236
timestamp 0
transform 1 0 22264 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_239
timestamp 0
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_242
timestamp 0
transform 1 0 22816 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_245
timestamp 0
transform 1 0 23092 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_248
timestamp 0
transform 1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_253
timestamp 0
transform 1 0 23828 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_256
timestamp 0
transform 1 0 24104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_259
timestamp 0
transform 1 0 24380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_262
timestamp 0
transform 1 0 24656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_265
timestamp 0
transform 1 0 24932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_268
timestamp 0
transform 1 0 25208 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_271
timestamp 0
transform 1 0 25484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_274
timestamp 0
transform 1 0 25760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_277
timestamp 0
transform 1 0 26036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_280
timestamp 0
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_283
timestamp 0
transform 1 0 26588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_286
timestamp 0
transform 1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_289
timestamp 0
transform 1 0 27140 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_292
timestamp 0
transform 1 0 27416 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_295
timestamp 0
transform 1 0 27692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_298
timestamp 0
transform 1 0 27968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_301
timestamp 0
transform 1 0 28244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_304
timestamp 0
transform 1 0 28520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_309
timestamp 0
transform 1 0 28980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_312
timestamp 0
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_315
timestamp 0
transform 1 0 29532 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_318
timestamp 0
transform 1 0 29808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_321
timestamp 0
transform 1 0 30084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_324
timestamp 0
transform 1 0 30360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_327
timestamp 0
transform 1 0 30636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_330
timestamp 0
transform 1 0 30912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_333
timestamp 0
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 0
transform 1 0 828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_6
timestamp 0
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_9
timestamp 0
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_12
timestamp 0
transform 1 0 1656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_15
timestamp 0
transform 1 0 1932 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_18
timestamp 0
transform 1 0 2208 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_21
timestamp 0
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_24
timestamp 0
transform 1 0 2760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_35
timestamp 0
transform 1 0 3772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_38
timestamp 0
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_41
timestamp 0
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_44
timestamp 0
transform 1 0 4600 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_47
timestamp 0
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_50
timestamp 0
transform 1 0 5152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 0
transform 1 0 5428 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 0
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_60
timestamp 0
transform 1 0 6072 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_63
timestamp 0
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_87
timestamp 0
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_90
timestamp 0
transform 1 0 8832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_93
timestamp 0
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_96
timestamp 0
transform 1 0 9384 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_99
timestamp 0
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_102
timestamp 0
transform 1 0 9936 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_105
timestamp 0
transform 1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 0
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_116
timestamp 0
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_119
timestamp 0
transform 1 0 11500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_122
timestamp 0
transform 1 0 11776 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_125
timestamp 0
transform 1 0 12052 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_128
timestamp 0
transform 1 0 12328 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_148
timestamp 0
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_154
timestamp 0
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_157
timestamp 0
transform 1 0 14996 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_160
timestamp 0
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_163
timestamp 0
transform 1 0 15548 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 0
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_169
timestamp 0
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_172
timestamp 0
transform 1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_175
timestamp 0
transform 1 0 16652 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_178
timestamp 0
transform 1 0 16928 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_181
timestamp 0
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_184
timestamp 0
transform 1 0 17480 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_187
timestamp 0
transform 1 0 17756 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_190
timestamp 0
transform 1 0 18032 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_193
timestamp 0
transform 1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_196
timestamp 0
transform 1 0 18584 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_199
timestamp 0
transform 1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_202
timestamp 0
transform 1 0 19136 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_205
timestamp 0
transform 1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_208
timestamp 0
transform 1 0 19688 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_211
timestamp 0
transform 1 0 19964 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_214
timestamp 0
transform 1 0 20240 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_217
timestamp 0
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_220
timestamp 0
transform 1 0 20792 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_225
timestamp 0
transform 1 0 21252 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_228
timestamp 0
transform 1 0 21528 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_231
timestamp 0
transform 1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_234
timestamp 0
transform 1 0 22080 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_237
timestamp 0
transform 1 0 22356 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_240
timestamp 0
transform 1 0 22632 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_243
timestamp 0
transform 1 0 22908 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_246
timestamp 0
transform 1 0 23184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_249
timestamp 0
transform 1 0 23460 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_252
timestamp 0
transform 1 0 23736 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_255
timestamp 0
transform 1 0 24012 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_258
timestamp 0
transform 1 0 24288 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_261
timestamp 0
transform 1 0 24564 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_264
timestamp 0
transform 1 0 24840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_267
timestamp 0
transform 1 0 25116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_270
timestamp 0
transform 1 0 25392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_273
timestamp 0
transform 1 0 25668 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_276
timestamp 0
transform 1 0 25944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 0
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_281
timestamp 0
transform 1 0 26404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_284
timestamp 0
transform 1 0 26680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_287
timestamp 0
transform 1 0 26956 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_290
timestamp 0
transform 1 0 27232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_293
timestamp 0
transform 1 0 27508 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_296
timestamp 0
transform 1 0 27784 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_299
timestamp 0
transform 1 0 28060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_302
timestamp 0
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_305
timestamp 0
transform 1 0 28612 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_308
timestamp 0
transform 1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_311
timestamp 0
transform 1 0 29164 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_314
timestamp 0
transform 1 0 29440 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_317
timestamp 0
transform 1 0 29716 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_320
timestamp 0
transform 1 0 29992 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_323
timestamp 0
transform 1 0 30268 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_326
timestamp 0
transform 1 0 30544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_329
timestamp 0
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_332
timestamp 0
transform 1 0 31096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 0
transform 1 0 828 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_6
timestamp 0
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_9
timestamp 0
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_12
timestamp 0
transform 1 0 1656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_15
timestamp 0
transform 1 0 1932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_18
timestamp 0
transform 1 0 2208 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_21
timestamp 0
transform 1 0 2484 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_24
timestamp 0
transform 1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 0
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_32
timestamp 0
transform 1 0 3496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_42
timestamp 0
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_45
timestamp 0
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_53
timestamp 0
transform 1 0 5428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_56
timestamp 0
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_59
timestamp 0
transform 1 0 5980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_62
timestamp 0
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_74
timestamp 0
transform 1 0 7360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 0
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_93
timestamp 0
transform 1 0 9108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_96
timestamp 0
transform 1 0 9384 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_99
timestamp 0
transform 1 0 9660 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_112
timestamp 0
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_121
timestamp 0
transform 1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_124
timestamp 0
transform 1 0 11960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_127
timestamp 0
transform 1 0 12236 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_130
timestamp 0
transform 1 0 12512 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 0
transform 1 0 13156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_146
timestamp 0
transform 1 0 13984 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_149
timestamp 0
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_157
timestamp 0
transform 1 0 14996 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_168
timestamp 0
transform 1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_171
timestamp 0
transform 1 0 16284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_174
timestamp 0
transform 1 0 16560 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_177
timestamp 0
transform 1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_180
timestamp 0
transform 1 0 17112 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_183
timestamp 0
transform 1 0 17388 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_189
timestamp 0
transform 1 0 17940 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_192
timestamp 0
transform 1 0 18216 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 0
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_197
timestamp 0
transform 1 0 18676 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_200
timestamp 0
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_207
timestamp 0
transform 1 0 19596 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_234
timestamp 0
transform 1 0 22080 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_248
timestamp 0
transform 1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_253
timestamp 0
transform 1 0 23828 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_265
timestamp 0
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_280
timestamp 0
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_283
timestamp 0
transform 1 0 26588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_286
timestamp 0
transform 1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_289
timestamp 0
transform 1 0 27140 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_292
timestamp 0
transform 1 0 27416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_295
timestamp 0
transform 1 0 27692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_298
timestamp 0
transform 1 0 27968 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_301
timestamp 0
transform 1 0 28244 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_304
timestamp 0
transform 1 0 28520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 0
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_309
timestamp 0
transform 1 0 28980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_312
timestamp 0
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_315
timestamp 0
transform 1 0 29532 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_318
timestamp 0
transform 1 0 29808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_321
timestamp 0
transform 1 0 30084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_324
timestamp 0
transform 1 0 30360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_327
timestamp 0
transform 1 0 30636 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_330
timestamp 0
transform 1 0 30912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_333
timestamp 0
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 0
transform 1 0 828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_6
timestamp 0
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_9
timestamp 0
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_12
timestamp 0
transform 1 0 1656 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_23
timestamp 0
transform 1 0 2668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_26
timestamp 0
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_44
timestamp 0
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_50
timestamp 0
transform 1 0 5152 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 0
transform 1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_66
timestamp 0
transform 1 0 6624 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_69
timestamp 0
transform 1 0 6900 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_72
timestamp 0
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_84
timestamp 0
transform 1 0 8280 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_87
timestamp 0
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_90
timestamp 0
transform 1 0 8832 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_93
timestamp 0
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_96
timestamp 0
transform 1 0 9384 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 0
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 0
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_116
timestamp 0
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_126
timestamp 0
transform 1 0 12144 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_129
timestamp 0
transform 1 0 12420 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_132
timestamp 0
transform 1 0 12696 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_135
timestamp 0
transform 1 0 12972 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_138
timestamp 0
transform 1 0 13248 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_141
timestamp 0
transform 1 0 13524 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_144
timestamp 0
transform 1 0 13800 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_147
timestamp 0
transform 1 0 14076 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_150
timestamp 0
transform 1 0 14352 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_153
timestamp 0
transform 1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_156
timestamp 0
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_159
timestamp 0
transform 1 0 15180 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 0
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_169
timestamp 0
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_172
timestamp 0
transform 1 0 16376 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_182
timestamp 0
transform 1 0 17296 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_185
timestamp 0
transform 1 0 17572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_188
timestamp 0
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_206
timestamp 0
transform 1 0 19504 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_209
timestamp 0
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_212
timestamp 0
transform 1 0 20056 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_220
timestamp 0
transform 1 0 20792 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_225
timestamp 0
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_228
timestamp 0
transform 1 0 21528 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_231
timestamp 0
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_234
timestamp 0
transform 1 0 22080 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_245
timestamp 0
transform 1 0 23092 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_248
timestamp 0
transform 1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_251
timestamp 0
transform 1 0 23644 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_254
timestamp 0
transform 1 0 23920 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_257
timestamp 0
transform 1 0 24196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_260
timestamp 0
transform 1 0 24472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_263
timestamp 0
transform 1 0 24748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_269
timestamp 0
transform 1 0 25300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_272
timestamp 0
transform 1 0 25576 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_275
timestamp 0
transform 1 0 25852 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_278
timestamp 0
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_281
timestamp 0
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_293
timestamp 0
transform 1 0 27508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_296
timestamp 0
transform 1 0 27784 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_299
timestamp 0
transform 1 0 28060 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_302
timestamp 0
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_305
timestamp 0
transform 1 0 28612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_308
timestamp 0
transform 1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_311
timestamp 0
transform 1 0 29164 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_315
timestamp 0
transform 1 0 29532 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_318
timestamp 0
transform 1 0 29808 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_321
timestamp 0
transform 1 0 30084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_324
timestamp 0
transform 1 0 30360 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_327
timestamp 0
transform 1 0 30636 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_330
timestamp 0
transform 1 0 30912 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_333
timestamp 0
transform 1 0 31188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_3
timestamp 0
transform 1 0 828 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_6
timestamp 0
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_9
timestamp 0
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_12
timestamp 0
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 0
transform 1 0 2852 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_34
timestamp 0
transform 1 0 3680 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_37
timestamp 0
transform 1 0 3956 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_40
timestamp 0
transform 1 0 4232 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_43
timestamp 0
transform 1 0 4508 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_46
timestamp 0
transform 1 0 4784 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_49
timestamp 0
transform 1 0 5060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_52
timestamp 0
transform 1 0 5336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_55
timestamp 0
transform 1 0 5612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_67
timestamp 0
transform 1 0 6716 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_70
timestamp 0
transform 1 0 6992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_73
timestamp 0
transform 1 0 7268 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 0
transform 1 0 8004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_85
timestamp 0
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_88
timestamp 0
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_91
timestamp 0
transform 1 0 8924 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_94
timestamp 0
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_97
timestamp 0
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_100
timestamp 0
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_103
timestamp 0
transform 1 0 10028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_106
timestamp 0
transform 1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_109
timestamp 0
transform 1 0 10580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_112
timestamp 0
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_115
timestamp 0
transform 1 0 11132 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_118
timestamp 0
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_127
timestamp 0
transform 1 0 12236 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_136
timestamp 0
transform 1 0 13064 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_149
timestamp 0
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_171
timestamp 0
transform 1 0 16284 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_174
timestamp 0
transform 1 0 16560 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_177
timestamp 0
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_183
timestamp 0
transform 1 0 17388 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_186
timestamp 0
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_189
timestamp 0
transform 1 0 17940 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_192
timestamp 0
transform 1 0 18216 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_203
timestamp 0
transform 1 0 19228 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_206
timestamp 0
transform 1 0 19504 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_209
timestamp 0
transform 1 0 19780 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_212
timestamp 0
transform 1 0 20056 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_215
timestamp 0
transform 1 0 20332 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_228
timestamp 0
transform 1 0 21528 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_231
timestamp 0
transform 1 0 21804 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_234
timestamp 0
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_237
timestamp 0
transform 1 0 22356 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_240
timestamp 0
transform 1 0 22632 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_243
timestamp 0
transform 1 0 22908 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_260
timestamp 0
transform 1 0 24472 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_267
timestamp 0
transform 1 0 25116 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_273
timestamp 0
transform 1 0 25668 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_276
timestamp 0
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_305
timestamp 0
transform 1 0 28612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_330
timestamp 0
transform 1 0 30912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_333
timestamp 0
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 0
transform 1 0 828 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_6
timestamp 0
transform 1 0 1104 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_25
timestamp 0
transform 1 0 2852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_43
timestamp 0
transform 1 0 4508 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_52
timestamp 0
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 0
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 0
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_66
timestamp 0
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_69
timestamp 0
transform 1 0 6900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_72
timestamp 0
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_81
timestamp 0
transform 1 0 8004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 0
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_105
timestamp 0
transform 1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_108
timestamp 0
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_125
timestamp 0
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_128
timestamp 0
transform 1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_131
timestamp 0
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_134
timestamp 0
transform 1 0 12880 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_137
timestamp 0
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_140
timestamp 0
transform 1 0 13432 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_143
timestamp 0
transform 1 0 13708 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_146
timestamp 0
transform 1 0 13984 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_149
timestamp 0
transform 1 0 14260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_152
timestamp 0
transform 1 0 14536 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_155
timestamp 0
transform 1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_158
timestamp 0
transform 1 0 15088 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_161
timestamp 0
transform 1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_164
timestamp 0
transform 1 0 15640 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 0
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_177
timestamp 0
transform 1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_180
timestamp 0
transform 1 0 17112 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_190
timestamp 0
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_198
timestamp 0
transform 1 0 18768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_201
timestamp 0
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_216
timestamp 0
transform 1 0 20424 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_219
timestamp 0
transform 1 0 20700 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 0
transform 1 0 20976 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 0
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_236
timestamp 0
transform 1 0 22264 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_240
timestamp 0
transform 1 0 22632 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_243
timestamp 0
transform 1 0 22908 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_246
timestamp 0
transform 1 0 23184 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_249
timestamp 0
transform 1 0 23460 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_257
timestamp 0
transform 1 0 24196 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_260
timestamp 0
transform 1 0 24472 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_263
timestamp 0
transform 1 0 24748 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_266
timestamp 0
transform 1 0 25024 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_272
timestamp 0
transform 1 0 25576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 0
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_281
timestamp 0
transform 1 0 26404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_292
timestamp 0
transform 1 0 27416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_295
timestamp 0
transform 1 0 27692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_319
timestamp 0
transform 1 0 29900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_322
timestamp 0
transform 1 0 30176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_325
timestamp 0
transform 1 0 30452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_328
timestamp 0
transform 1 0 30728 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_331
timestamp 0
transform 1 0 31004 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_334
timestamp 0
transform 1 0 31280 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_3
timestamp 0
transform 1 0 828 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_6
timestamp 0
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_15
timestamp 0
transform 1 0 1932 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_18
timestamp 0
transform 1 0 2208 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_21
timestamp 0
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 0
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_44
timestamp 0
transform 1 0 4600 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_47
timestamp 0
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_61
timestamp 0
transform 1 0 6164 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_64
timestamp 0
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_80
timestamp 0
transform 1 0 7912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 0
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_88
timestamp 0
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_91
timestamp 0
transform 1 0 8924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_94
timestamp 0
transform 1 0 9200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_97
timestamp 0
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_100
timestamp 0
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_103
timestamp 0
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_112
timestamp 0
transform 1 0 10856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_115
timestamp 0
transform 1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_118
timestamp 0
transform 1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_121
timestamp 0
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_124
timestamp 0
transform 1 0 11960 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_127
timestamp 0
transform 1 0 12236 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_141
timestamp 0
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_163
timestamp 0
transform 1 0 15548 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_166
timestamp 0
transform 1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_175
timestamp 0
transform 1 0 16652 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_178
timestamp 0
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_181
timestamp 0
transform 1 0 17204 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_184
timestamp 0
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_187
timestamp 0
transform 1 0 17756 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_190
timestamp 0
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 0
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_197
timestamp 0
transform 1 0 18676 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_200
timestamp 0
transform 1 0 18952 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_207
timestamp 0
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_210
timestamp 0
transform 1 0 19872 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_213
timestamp 0
transform 1 0 20148 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_216
timestamp 0
transform 1 0 20424 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_219
timestamp 0
transform 1 0 20700 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_222
timestamp 0
transform 1 0 20976 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_225
timestamp 0
transform 1 0 21252 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_228
timestamp 0
transform 1 0 21528 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_231
timestamp 0
transform 1 0 21804 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_235
timestamp 0
transform 1 0 22172 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_238
timestamp 0
transform 1 0 22448 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_241
timestamp 0
transform 1 0 22724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_244
timestamp 0
transform 1 0 23000 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_247
timestamp 0
transform 1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 0
transform 1 0 23552 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_261
timestamp 0
transform 1 0 24564 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_264
timestamp 0
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_269
timestamp 0
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_276
timestamp 0
transform 1 0 25944 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_279
timestamp 0
transform 1 0 26220 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_282
timestamp 0
transform 1 0 26496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_285
timestamp 0
transform 1 0 26772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_288
timestamp 0
transform 1 0 27048 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_292
timestamp 0
transform 1 0 27416 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_295
timestamp 0
transform 1 0 27692 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_298
timestamp 0
transform 1 0 27968 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_301
timestamp 0
transform 1 0 28244 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_304
timestamp 0
transform 1 0 28520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_326
timestamp 0
transform 1 0 30544 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_329
timestamp 0
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_332
timestamp 0
transform 1 0 31096 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 0
transform 1 0 828 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_6
timestamp 0
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_9
timestamp 0
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_25
timestamp 0
transform 1 0 2852 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_28
timestamp 0
transform 1 0 3128 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 0
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_60
timestamp 0
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_79
timestamp 0
transform 1 0 7820 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_82
timestamp 0
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_100
timestamp 0
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_103
timestamp 0
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_108
timestamp 0
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_126
timestamp 0
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_142
timestamp 0
transform 1 0 13616 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_145
timestamp 0
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_148
timestamp 0
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_163
timestamp 0
transform 1 0 15548 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 0
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 0
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_202
timestamp 0
transform 1 0 19136 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_205
timestamp 0
transform 1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_208
timestamp 0
transform 1 0 19688 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_220
timestamp 0
transform 1 0 20792 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 0
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 0
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_240
timestamp 0
transform 1 0 22632 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_243
timestamp 0
transform 1 0 22908 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_246
timestamp 0
transform 1 0 23184 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_264
timestamp 0
transform 1 0 24840 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_276
timestamp 0
transform 1 0 25944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_281
timestamp 0
transform 1 0 26404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_284
timestamp 0
transform 1 0 26680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_287
timestamp 0
transform 1 0 26956 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_290
timestamp 0
transform 1 0 27232 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_297
timestamp 0
transform 1 0 27876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_300
timestamp 0
transform 1 0 28152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_303
timestamp 0
transform 1 0 28428 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_316
timestamp 0
transform 1 0 29624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_334
timestamp 0
transform 1 0 31280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_3
timestamp 0
transform 1 0 828 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_6
timestamp 0
transform 1 0 1104 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 0
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 0
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_32
timestamp 0
transform 1 0 3496 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_56
timestamp 0
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_59
timestamp 0
transform 1 0 5980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_62
timestamp 0
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_71
timestamp 0
transform 1 0 7084 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_74
timestamp 0
transform 1 0 7360 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_77
timestamp 0
transform 1 0 7636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_80
timestamp 0
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_95
timestamp 0
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_98
timestamp 0
transform 1 0 9568 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_101
timestamp 0
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_108
timestamp 0
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_111
timestamp 0
transform 1 0 10764 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_114
timestamp 0
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_117
timestamp 0
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_120
timestamp 0
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_123
timestamp 0
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_126
timestamp 0
transform 1 0 12144 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_129
timestamp 0
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_136
timestamp 0
transform 1 0 13064 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_141
timestamp 0
transform 1 0 13524 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_144
timestamp 0
transform 1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_147
timestamp 0
transform 1 0 14076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_150
timestamp 0
transform 1 0 14352 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_166
timestamp 0
transform 1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_181
timestamp 0
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_184
timestamp 0
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_187
timestamp 0
transform 1 0 17756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_190
timestamp 0
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 0
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_197
timestamp 0
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_200
timestamp 0
transform 1 0 18952 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_203
timestamp 0
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_206
timestamp 0
transform 1 0 19504 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_209
timestamp 0
transform 1 0 19780 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_212
timestamp 0
transform 1 0 20056 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_220
timestamp 0
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_244
timestamp 0
transform 1 0 23000 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_247
timestamp 0
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 0
transform 1 0 23552 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_266
timestamp 0
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_279
timestamp 0
transform 1 0 26220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_282
timestamp 0
transform 1 0 26496 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_285
timestamp 0
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_309
timestamp 0
transform 1 0 28980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_330
timestamp 0
transform 1 0 30912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 0
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 0
transform 1 0 828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_6
timestamp 0
transform 1 0 1104 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_21
timestamp 0
transform 1 0 2484 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_24
timestamp 0
transform 1 0 2760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_27
timestamp 0
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_30
timestamp 0
transform 1 0 3312 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_33
timestamp 0
transform 1 0 3588 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_36
timestamp 0
transform 1 0 3864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_39
timestamp 0
transform 1 0 4140 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_42
timestamp 0
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_49
timestamp 0
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 0
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 0
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_60
timestamp 0
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_63
timestamp 0
transform 1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_66
timestamp 0
transform 1 0 6624 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_69
timestamp 0
transform 1 0 6900 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_72
timestamp 0
transform 1 0 7176 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_75
timestamp 0
transform 1 0 7452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_78
timestamp 0
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 0
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_84
timestamp 0
transform 1 0 8280 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_100
timestamp 0
transform 1 0 9752 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_103
timestamp 0
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_106
timestamp 0
transform 1 0 10304 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 0
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_133
timestamp 0
transform 1 0 12788 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 0
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 0
transform 1 0 16100 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_183
timestamp 0
transform 1 0 17388 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_186
timestamp 0
transform 1 0 17664 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_189
timestamp 0
transform 1 0 17940 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_192
timestamp 0
transform 1 0 18216 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_209
timestamp 0
transform 1 0 19780 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_212
timestamp 0
transform 1 0 20056 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_219
timestamp 0
transform 1 0 20700 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 0
transform 1 0 20976 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 0
transform 1 0 21252 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_228
timestamp 0
transform 1 0 21528 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_241
timestamp 0
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_252
timestamp 0
transform 1 0 23736 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_255
timestamp 0
transform 1 0 24012 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_272
timestamp 0
transform 1 0 25576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 0
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_311
timestamp 0
transform 1 0 29164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_330
timestamp 0
transform 1 0 30912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_333
timestamp 0
transform 1 0 31188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_3
timestamp 0
transform 1 0 828 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_6
timestamp 0
transform 1 0 1104 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_19
timestamp 0
transform 1 0 2300 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_22
timestamp 0
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 0
transform 1 0 2852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_44
timestamp 0
transform 1 0 4600 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_59
timestamp 0
transform 1 0 5980 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_62
timestamp 0
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 0
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_93
timestamp 0
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_96
timestamp 0
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_99
timestamp 0
transform 1 0 9660 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_102
timestamp 0
transform 1 0 9936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_105
timestamp 0
transform 1 0 10212 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_109
timestamp 0
transform 1 0 10580 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_112
timestamp 0
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_122
timestamp 0
transform 1 0 11776 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 0
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 0
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_162
timestamp 0
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_165
timestamp 0
transform 1 0 15732 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_168
timestamp 0
transform 1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_171
timestamp 0
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_174
timestamp 0
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_177
timestamp 0
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_190
timestamp 0
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 0
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_202
timestamp 0
transform 1 0 19136 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_205
timestamp 0
transform 1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_208
timestamp 0
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_214
timestamp 0
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_258
timestamp 0
transform 1 0 24288 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_262
timestamp 0
transform 1 0 24656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_265
timestamp 0
transform 1 0 24932 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_283
timestamp 0
transform 1 0 26588 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_286
timestamp 0
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_293
timestamp 0
transform 1 0 27508 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_316
timestamp 0
transform 1 0 29624 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_324
timestamp 0
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_330
timestamp 0
transform 1 0 30912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_333
timestamp 0
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 0
transform 1 0 828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_24
timestamp 0
transform 1 0 2760 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_34
timestamp 0
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_37
timestamp 0
transform 1 0 3956 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_40
timestamp 0
transform 1 0 4232 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_46
timestamp 0
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_51
timestamp 0
transform 1 0 5244 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 0
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_57
timestamp 0
transform 1 0 5796 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_60
timestamp 0
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_68
timestamp 0
transform 1 0 6808 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_72
timestamp 0
transform 1 0 7176 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_75
timestamp 0
transform 1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_78
timestamp 0
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_81
timestamp 0
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_84
timestamp 0
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_87
timestamp 0
transform 1 0 8556 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_100
timestamp 0
transform 1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_103
timestamp 0
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_106
timestamp 0
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 0
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_118
timestamp 0
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_121
timestamp 0
transform 1 0 11684 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_124
timestamp 0
transform 1 0 11960 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_128
timestamp 0
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_136
timestamp 0
transform 1 0 13064 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_139
timestamp 0
transform 1 0 13340 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_142
timestamp 0
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_174
timestamp 0
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_177
timestamp 0
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_188
timestamp 0
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_191
timestamp 0
transform 1 0 18124 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_197
timestamp 0
transform 1 0 18676 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_204
timestamp 0
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_207
timestamp 0
transform 1 0 19596 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_217
timestamp 0
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_220
timestamp 0
transform 1 0 20792 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 0
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_232
timestamp 0
transform 1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_235
timestamp 0
transform 1 0 22172 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_238
timestamp 0
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_241
timestamp 0
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_251
timestamp 0
transform 1 0 23644 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_268
timestamp 0
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_276
timestamp 0
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 0
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_281
timestamp 0
transform 1 0 26404 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_284
timestamp 0
transform 1 0 26680 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_295
timestamp 0
transform 1 0 27692 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_298
timestamp 0
transform 1 0 27968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_315
timestamp 0
transform 1 0 29532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_332
timestamp 0
transform 1 0 31096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_3
timestamp 0
transform 1 0 828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_6
timestamp 0
transform 1 0 1104 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_15
timestamp 0
transform 1 0 1932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_18
timestamp 0
transform 1 0 2208 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_21
timestamp 0
transform 1 0 2484 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_24
timestamp 0
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_36
timestamp 0
transform 1 0 3864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_39
timestamp 0
transform 1 0 4140 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_42
timestamp 0
transform 1 0 4416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_71
timestamp 0
transform 1 0 7084 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_78
timestamp 0
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 0
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_101
timestamp 0
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_110
timestamp 0
transform 1 0 10672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_113
timestamp 0
transform 1 0 10948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_116
timestamp 0
transform 1 0 11224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_123
timestamp 0
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_126
timestamp 0
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 0
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_144
timestamp 0
transform 1 0 13800 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_187
timestamp 0
transform 1 0 17756 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_191
timestamp 0
transform 1 0 18124 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 0
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_213
timestamp 0
transform 1 0 20148 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_221
timestamp 0
transform 1 0 20884 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_224
timestamp 0
transform 1 0 21160 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_227
timestamp 0
transform 1 0 21436 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_240
timestamp 0
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_248
timestamp 0
transform 1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 0
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_253
timestamp 0
transform 1 0 23828 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_278
timestamp 0
transform 1 0 26128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_304
timestamp 0
transform 1 0 28520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 0
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_309
timestamp 0
transform 1 0 28980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_333
timestamp 0
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 0
transform 1 0 828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_6
timestamp 0
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_9
timestamp 0
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_12
timestamp 0
transform 1 0 1656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_15
timestamp 0
transform 1 0 1932 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_18
timestamp 0
transform 1 0 2208 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_21
timestamp 0
transform 1 0 2484 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_24
timestamp 0
transform 1 0 2760 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_27
timestamp 0
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_41
timestamp 0
transform 1 0 4324 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_44
timestamp 0
transform 1 0 4600 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_47
timestamp 0
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_50
timestamp 0
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 0
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_57
timestamp 0
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_71
timestamp 0
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_74
timestamp 0
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_80
timestamp 0
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_83
timestamp 0
transform 1 0 8188 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_90
timestamp 0
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_106
timestamp 0
transform 1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 0
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_119
timestamp 0
transform 1 0 11500 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_122
timestamp 0
transform 1 0 11776 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 0
transform 1 0 12052 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_128
timestamp 0
transform 1 0 12328 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_131
timestamp 0
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_139
timestamp 0
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_142
timestamp 0
transform 1 0 13616 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_145
timestamp 0
transform 1 0 13892 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_156
timestamp 0
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_159
timestamp 0
transform 1 0 15180 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_162
timestamp 0
transform 1 0 15456 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 0
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 0
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_172
timestamp 0
transform 1 0 16376 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_182
timestamp 0
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_185
timestamp 0
transform 1 0 17572 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_188
timestamp 0
transform 1 0 17848 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_191
timestamp 0
transform 1 0 18124 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_194
timestamp 0
transform 1 0 18400 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_197
timestamp 0
transform 1 0 18676 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_209
timestamp 0
transform 1 0 19780 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_212
timestamp 0
transform 1 0 20056 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_215
timestamp 0
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_218
timestamp 0
transform 1 0 20608 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_225
timestamp 0
transform 1 0 21252 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_228
timestamp 0
transform 1 0 21528 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_236
timestamp 0
transform 1 0 22264 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_239
timestamp 0
transform 1 0 22540 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_242
timestamp 0
transform 1 0 22816 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_248
timestamp 0
transform 1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_251
timestamp 0
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_258
timestamp 0
transform 1 0 24288 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_267
timestamp 0
transform 1 0 25116 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_270
timestamp 0
transform 1 0 25392 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_295
timestamp 0
transform 1 0 27692 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_305
timestamp 0
transform 1 0 28612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_312
timestamp 0
transform 1 0 29256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_3
timestamp 0
transform 1 0 828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_6
timestamp 0
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_9
timestamp 0
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_17
timestamp 0
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_20
timestamp 0
transform 1 0 2392 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_23
timestamp 0
transform 1 0 2668 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 0
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_42
timestamp 0
transform 1 0 4416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_45
timestamp 0
transform 1 0 4692 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 0
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_105
timestamp 0
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_124
timestamp 0
transform 1 0 11960 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_127
timestamp 0
transform 1 0 12236 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_130
timestamp 0
transform 1 0 12512 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_133
timestamp 0
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_136
timestamp 0
transform 1 0 13064 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 0
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_155
timestamp 0
transform 1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_158
timestamp 0
transform 1 0 15088 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_167
timestamp 0
transform 1 0 15916 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_170
timestamp 0
transform 1 0 16192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_173
timestamp 0
transform 1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_176
timestamp 0
transform 1 0 16744 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_179
timestamp 0
transform 1 0 17020 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_191
timestamp 0
transform 1 0 18124 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_206
timestamp 0
transform 1 0 19504 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_217
timestamp 0
transform 1 0 20516 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_220
timestamp 0
transform 1 0 20792 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_223
timestamp 0
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_232
timestamp 0
transform 1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_235
timestamp 0
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_246
timestamp 0
transform 1 0 23184 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 0
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 0
transform 1 0 23828 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_268
timestamp 0
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_271
timestamp 0
transform 1 0 25484 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_297
timestamp 0
transform 1 0 27876 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_300
timestamp 0
transform 1 0 28152 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_303
timestamp 0
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_309
timestamp 0
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_334
timestamp 0
transform 1 0 31280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_3
timestamp 0
transform 1 0 828 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_40
timestamp 0
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_49
timestamp 0
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_52
timestamp 0
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_57
timestamp 0
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_60
timestamp 0
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_63
timestamp 0
transform 1 0 6348 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 0
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_73
timestamp 0
transform 1 0 7268 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_76
timestamp 0
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_79
timestamp 0
transform 1 0 7820 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_83
timestamp 0
transform 1 0 8188 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_86
timestamp 0
transform 1 0 8464 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_89
timestamp 0
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_94
timestamp 0
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_99
timestamp 0
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_102
timestamp 0
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_105
timestamp 0
transform 1 0 10212 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_108
timestamp 0
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_123
timestamp 0
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_126
timestamp 0
transform 1 0 12144 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_140
timestamp 0
transform 1 0 13432 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_143
timestamp 0
transform 1 0 13708 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_146
timestamp 0
transform 1 0 13984 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_161
timestamp 0
transform 1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_164
timestamp 0
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 0
transform 1 0 16100 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_178
timestamp 0
transform 1 0 16928 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_181
timestamp 0
transform 1 0 17204 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_184
timestamp 0
transform 1 0 17480 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_187
timestamp 0
transform 1 0 17756 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_190
timestamp 0
transform 1 0 18032 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_193
timestamp 0
transform 1 0 18308 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_196
timestamp 0
transform 1 0 18584 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_199
timestamp 0
transform 1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_202
timestamp 0
transform 1 0 19136 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_205
timestamp 0
transform 1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_208
timestamp 0
transform 1 0 19688 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_211
timestamp 0
transform 1 0 19964 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_217
timestamp 0
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_220
timestamp 0
transform 1 0 20792 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 0
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_225
timestamp 0
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_228
timestamp 0
transform 1 0 21528 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_231
timestamp 0
transform 1 0 21804 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_234
timestamp 0
transform 1 0 22080 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 0
transform 1 0 22356 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_240
timestamp 0
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_245
timestamp 0
transform 1 0 23092 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_248
timestamp 0
transform 1 0 23368 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_256
timestamp 0
transform 1 0 24104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_265
timestamp 0
transform 1 0 24932 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_274
timestamp 0
transform 1 0 25760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_277
timestamp 0
transform 1 0 26036 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_281
timestamp 0
transform 1 0 26404 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_284
timestamp 0
transform 1 0 26680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_334
timestamp 0
transform 1 0 31280 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 0
transform 1 0 828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_6
timestamp 0
transform 1 0 1104 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_21
timestamp 0
transform 1 0 2484 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_40
timestamp 0
transform 1 0 4232 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_43
timestamp 0
transform 1 0 4508 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_50
timestamp 0
transform 1 0 5152 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 0
transform 1 0 5428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_56
timestamp 0
transform 1 0 5704 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_69
timestamp 0
transform 1 0 6900 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_72
timestamp 0
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_75
timestamp 0
transform 1 0 7452 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_91
timestamp 0
transform 1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_94
timestamp 0
transform 1 0 9200 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_97
timestamp 0
transform 1 0 9476 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_100
timestamp 0
transform 1 0 9752 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_103
timestamp 0
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_125
timestamp 0
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_128
timestamp 0
transform 1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_131
timestamp 0
transform 1 0 12604 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_134
timestamp 0
transform 1 0 12880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 0
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_141
timestamp 0
transform 1 0 13524 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_144
timestamp 0
transform 1 0 13800 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_147
timestamp 0
transform 1 0 14076 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_150
timestamp 0
transform 1 0 14352 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_163
timestamp 0
transform 1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_166
timestamp 0
transform 1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_169
timestamp 0
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_172
timestamp 0
transform 1 0 16376 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_175
timestamp 0
transform 1 0 16652 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_188
timestamp 0
transform 1 0 17848 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_191
timestamp 0
transform 1 0 18124 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 0
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_203
timestamp 0
transform 1 0 19228 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_206
timestamp 0
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_219
timestamp 0
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_222
timestamp 0
transform 1 0 20976 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_231
timestamp 0
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_242
timestamp 0
transform 1 0 22816 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_245
timestamp 0
transform 1 0 23092 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_248
timestamp 0
transform 1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 0
transform 1 0 23828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_262
timestamp 0
transform 1 0 24656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_265
timestamp 0
transform 1 0 24932 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_268
timestamp 0
transform 1 0 25208 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_287
timestamp 0
transform 1 0 26956 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_292
timestamp 0
transform 1 0 27416 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_295
timestamp 0
transform 1 0 27692 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_298
timestamp 0
transform 1 0 27968 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 0
transform 1 0 28704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_309
timestamp 0
transform 1 0 28980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_3
timestamp 0
transform 1 0 828 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_6
timestamp 0
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_9
timestamp 0
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_15
timestamp 0
transform 1 0 1932 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_18
timestamp 0
transform 1 0 2208 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_21
timestamp 0
transform 1 0 2484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_24
timestamp 0
transform 1 0 2760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_27
timestamp 0
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_37
timestamp 0
transform 1 0 3956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_40
timestamp 0
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_43
timestamp 0
transform 1 0 4508 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_50
timestamp 0
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 0
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_57
timestamp 0
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_60
timestamp 0
transform 1 0 6072 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_63
timestamp 0
transform 1 0 6348 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_66
timestamp 0
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_75
timestamp 0
transform 1 0 7452 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_78
timestamp 0
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_81
timestamp 0
transform 1 0 8004 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_84
timestamp 0
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_87
timestamp 0
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_90
timestamp 0
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 0
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 0
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_116
timestamp 0
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_119
timestamp 0
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_122
timestamp 0
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_125
timestamp 0
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_130
timestamp 0
transform 1 0 12512 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_133
timestamp 0
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 0
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_169
timestamp 0
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_172
timestamp 0
transform 1 0 16376 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_194
timestamp 0
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_204
timestamp 0
transform 1 0 19320 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_207
timestamp 0
transform 1 0 19596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_210
timestamp 0
transform 1 0 19872 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_213
timestamp 0
transform 1 0 20148 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_216
timestamp 0
transform 1 0 20424 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_219
timestamp 0
transform 1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 0
transform 1 0 20976 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_225
timestamp 0
transform 1 0 21252 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_228
timestamp 0
transform 1 0 21528 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_231
timestamp 0
transform 1 0 21804 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_252
timestamp 0
transform 1 0 23736 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_255
timestamp 0
transform 1 0 24012 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_274
timestamp 0
transform 1 0 25760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_296
timestamp 0
transform 1 0 27784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_304
timestamp 0
transform 1 0 28520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_312
timestamp 0
transform 1 0 29256 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_315
timestamp 0
transform 1 0 29532 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_318
timestamp 0
transform 1 0 29808 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_326
timestamp 0
transform 1 0 30544 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_329
timestamp 0
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_332
timestamp 0
transform 1 0 31096 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_3
timestamp 0
transform 1 0 828 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_6
timestamp 0
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_9
timestamp 0
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_12
timestamp 0
transform 1 0 1656 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_15
timestamp 0
transform 1 0 1932 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_18
timestamp 0
transform 1 0 2208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_21
timestamp 0
transform 1 0 2484 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_24
timestamp 0
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 0
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_32
timestamp 0
transform 1 0 3496 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_35
timestamp 0
transform 1 0 3772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_38
timestamp 0
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_56
timestamp 0
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_59
timestamp 0
transform 1 0 5980 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_75
timestamp 0
transform 1 0 7452 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_78
timestamp 0
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_92
timestamp 0
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_95
timestamp 0
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_98
timestamp 0
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_107
timestamp 0
transform 1 0 10396 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_110
timestamp 0
transform 1 0 10672 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_113
timestamp 0
transform 1 0 10948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_116
timestamp 0
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_121
timestamp 0
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_124
timestamp 0
transform 1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 0
transform 1 0 13524 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_146
timestamp 0
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_149
timestamp 0
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_152
timestamp 0
transform 1 0 14536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_164
timestamp 0
transform 1 0 15640 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_167
timestamp 0
transform 1 0 15916 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_170
timestamp 0
transform 1 0 16192 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_173
timestamp 0
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_197
timestamp 0
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_212
timestamp 0
transform 1 0 20056 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_215
timestamp 0
transform 1 0 20332 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_224
timestamp 0
transform 1 0 21160 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_227
timestamp 0
transform 1 0 21436 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_230
timestamp 0
transform 1 0 21712 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_233
timestamp 0
transform 1 0 21988 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_236
timestamp 0
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_244
timestamp 0
transform 1 0 23000 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_247
timestamp 0
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 0
transform 1 0 23552 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_261
timestamp 0
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_266
timestamp 0
transform 1 0 25024 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_269
timestamp 0
transform 1 0 25300 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_272
timestamp 0
transform 1 0 25576 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_275
timestamp 0
transform 1 0 25852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_278
timestamp 0
transform 1 0 26128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_286
timestamp 0
transform 1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_289
timestamp 0
transform 1 0 27140 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_292
timestamp 0
transform 1 0 27416 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_295
timestamp 0
transform 1 0 27692 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_298
timestamp 0
transform 1 0 27968 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_301
timestamp 0
transform 1 0 28244 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_304
timestamp 0
transform 1 0 28520 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_317
timestamp 0
transform 1 0 29716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_330
timestamp 0
transform 1 0 30912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_333
timestamp 0
transform 1 0 31188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_17
timestamp 0
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_30
timestamp 0
transform 1 0 3312 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_33
timestamp 0
transform 1 0 3588 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_36
timestamp 0
transform 1 0 3864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_39
timestamp 0
transform 1 0 4140 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_42
timestamp 0
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_45
timestamp 0
transform 1 0 4692 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_48
timestamp 0
transform 1 0 4968 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_51
timestamp 0
transform 1 0 5244 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 0
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 0
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_60
timestamp 0
transform 1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_63
timestamp 0
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_70
timestamp 0
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_73
timestamp 0
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_79
timestamp 0
transform 1 0 7820 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_82
timestamp 0
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_91
timestamp 0
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_94
timestamp 0
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_97
timestamp 0
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_100
timestamp 0
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_103
timestamp 0
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_121
timestamp 0
transform 1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_124
timestamp 0
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_133
timestamp 0
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_143
timestamp 0
transform 1 0 13708 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_146
timestamp 0
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_149
timestamp 0
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_152
timestamp 0
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_174
timestamp 0
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_177
timestamp 0
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_186
timestamp 0
transform 1 0 17664 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_189
timestamp 0
transform 1 0 17940 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_192
timestamp 0
transform 1 0 18216 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_195
timestamp 0
transform 1 0 18492 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_206
timestamp 0
transform 1 0 19504 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_209
timestamp 0
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_212
timestamp 0
transform 1 0 20056 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_215
timestamp 0
transform 1 0 20332 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_218
timestamp 0
transform 1 0 20608 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_237
timestamp 0
transform 1 0 22356 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_240
timestamp 0
transform 1 0 22632 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_247
timestamp 0
transform 1 0 23276 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_250
timestamp 0
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_253
timestamp 0
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_273
timestamp 0
transform 1 0 25668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_290
timestamp 0
transform 1 0 27232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_293
timestamp 0
transform 1 0 27508 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_296
timestamp 0
transform 1 0 27784 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_312
timestamp 0
transform 1 0 29256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_315
timestamp 0
transform 1 0 29532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_321
timestamp 0
transform 1 0 30084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_324
timestamp 0
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_327
timestamp 0
transform 1 0 30636 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_330
timestamp 0
transform 1 0 30912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_333
timestamp 0
transform 1 0 31188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_3
timestamp 0
transform 1 0 828 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_6
timestamp 0
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_9
timestamp 0
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_12
timestamp 0
transform 1 0 1656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_15
timestamp 0
transform 1 0 1932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_18
timestamp 0
transform 1 0 2208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_21
timestamp 0
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_24
timestamp 0
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 0
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_36
timestamp 0
transform 1 0 3864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_39
timestamp 0
transform 1 0 4140 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_42
timestamp 0
transform 1 0 4416 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_57
timestamp 0
transform 1 0 5796 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_60
timestamp 0
transform 1 0 6072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_75
timestamp 0
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_88
timestamp 0
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_105
timestamp 0
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_108
timestamp 0
transform 1 0 10488 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_111
timestamp 0
transform 1 0 10764 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_114
timestamp 0
transform 1 0 11040 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_117
timestamp 0
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_120
timestamp 0
transform 1 0 11592 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_123
timestamp 0
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_126
timestamp 0
transform 1 0 12144 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_129
timestamp 0
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_132
timestamp 0
transform 1 0 12696 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_135
timestamp 0
transform 1 0 12972 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 0
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_149
timestamp 0
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_152
timestamp 0
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_155
timestamp 0
transform 1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_161
timestamp 0
transform 1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_164
timestamp 0
transform 1 0 15640 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_167
timestamp 0
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_170
timestamp 0
transform 1 0 16192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_173
timestamp 0
transform 1 0 16468 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_176
timestamp 0
transform 1 0 16744 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_191
timestamp 0
transform 1 0 18124 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 0
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_206
timestamp 0
transform 1 0 19504 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_209
timestamp 0
transform 1 0 19780 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_212
timestamp 0
transform 1 0 20056 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_215
timestamp 0
transform 1 0 20332 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_244
timestamp 0
transform 1 0 23000 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_247
timestamp 0
transform 1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 0
transform 1 0 23552 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_253
timestamp 0
transform 1 0 23828 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_256
timestamp 0
transform 1 0 24104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_259
timestamp 0
transform 1 0 24380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_262
timestamp 0
transform 1 0 24656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_265
timestamp 0
transform 1 0 24932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_268
timestamp 0
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_271
timestamp 0
transform 1 0 25484 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_278
timestamp 0
transform 1 0 26128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_281
timestamp 0
transform 1 0 26404 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_284
timestamp 0
transform 1 0 26680 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_287
timestamp 0
transform 1 0 26956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_290
timestamp 0
transform 1 0 27232 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_293
timestamp 0
transform 1 0 27508 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_296
timestamp 0
transform 1 0 27784 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_299
timestamp 0
transform 1 0 28060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_309
timestamp 0
transform 1 0 28980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_312
timestamp 0
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_315
timestamp 0
transform 1 0 29532 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_325
timestamp 0
transform 1 0 30452 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_328
timestamp 0
transform 1 0 30728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_334
timestamp 0
transform 1 0 31280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_3
timestamp 0
transform 1 0 828 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_6
timestamp 0
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_9
timestamp 0
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_21
timestamp 0
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_24
timestamp 0
transform 1 0 2760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_27
timestamp 0
transform 1 0 3036 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_34
timestamp 0
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_37
timestamp 0
transform 1 0 3956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_40
timestamp 0
transform 1 0 4232 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_43
timestamp 0
transform 1 0 4508 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_46
timestamp 0
transform 1 0 4784 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_64
timestamp 0
transform 1 0 6440 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_75
timestamp 0
transform 1 0 7452 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_79
timestamp 0
transform 1 0 7820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_82
timestamp 0
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_85
timestamp 0
transform 1 0 8372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_97
timestamp 0
transform 1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_100
timestamp 0
transform 1 0 9752 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_103
timestamp 0
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_106
timestamp 0
transform 1 0 10304 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_124
timestamp 0
transform 1 0 11960 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_127
timestamp 0
transform 1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_130
timestamp 0
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_137
timestamp 0
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_147
timestamp 0
transform 1 0 14076 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_150
timestamp 0
transform 1 0 14352 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_153
timestamp 0
transform 1 0 14628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_177
timestamp 0
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_180
timestamp 0
transform 1 0 17112 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_183
timestamp 0
transform 1 0 17388 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_186
timestamp 0
transform 1 0 17664 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_189
timestamp 0
transform 1 0 17940 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_196
timestamp 0
transform 1 0 18584 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_199
timestamp 0
transform 1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_202
timestamp 0
transform 1 0 19136 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_214
timestamp 0
transform 1 0 20240 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_217
timestamp 0
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_220
timestamp 0
transform 1 0 20792 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_225
timestamp 0
transform 1 0 21252 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_228
timestamp 0
transform 1 0 21528 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_231
timestamp 0
transform 1 0 21804 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_234
timestamp 0
transform 1 0 22080 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_237
timestamp 0
transform 1 0 22356 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_250
timestamp 0
transform 1 0 23552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_270
timestamp 0
transform 1 0 25392 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_276
timestamp 0
transform 1 0 25944 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_281
timestamp 0
transform 1 0 26404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_284
timestamp 0
transform 1 0 26680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_303
timestamp 0
transform 1 0 28428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_309
timestamp 0
transform 1 0 28980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_312
timestamp 0
transform 1 0 29256 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_333
timestamp 0
transform 1 0 31188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_3
timestamp 0
transform 1 0 828 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_6
timestamp 0
transform 1 0 1104 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_13
timestamp 0
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_16
timestamp 0
transform 1 0 2024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_19
timestamp 0
transform 1 0 2300 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_22
timestamp 0
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 0
transform 1 0 2852 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 0
transform 1 0 3220 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_41
timestamp 0
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_44
timestamp 0
transform 1 0 4600 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_52
timestamp 0
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_61
timestamp 0
transform 1 0 6164 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_64
timestamp 0
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_67
timestamp 0
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_77
timestamp 0
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 0
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_101
timestamp 0
transform 1 0 9844 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_104
timestamp 0
transform 1 0 10120 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_107
timestamp 0
transform 1 0 10396 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_110
timestamp 0
transform 1 0 10672 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_113
timestamp 0
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_124
timestamp 0
transform 1 0 11960 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_127
timestamp 0
transform 1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_130
timestamp 0
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_133
timestamp 0
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_136
timestamp 0
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13340 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_150
timestamp 0
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_158
timestamp 0
transform 1 0 15088 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_161
timestamp 0
transform 1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_164
timestamp 0
transform 1 0 15640 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_167
timestamp 0
transform 1 0 15916 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_170
timestamp 0
transform 1 0 16192 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_173
timestamp 0
transform 1 0 16468 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_176
timestamp 0
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_192
timestamp 0
transform 1 0 18216 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_197
timestamp 0
transform 1 0 18676 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_200
timestamp 0
transform 1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_203
timestamp 0
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_214
timestamp 0
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_223
timestamp 0
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_230
timestamp 0
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_240
timestamp 0
transform 1 0 22632 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_243
timestamp 0
transform 1 0 22908 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 0
transform 1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_253
timestamp 0
transform 1 0 23828 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_256
timestamp 0
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_266
timestamp 0
transform 1 0 25024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_269
timestamp 0
transform 1 0 25300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_284
timestamp 0
transform 1 0 26680 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_287
timestamp 0
transform 1 0 26956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_290
timestamp 0
transform 1 0 27232 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_293
timestamp 0
transform 1 0 27508 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_296
timestamp 0
transform 1 0 27784 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_300
timestamp 0
transform 1 0 28152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_303
timestamp 0
transform 1 0 28428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 0
transform 1 0 28704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_313
timestamp 0
transform 1 0 29348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_333
timestamp 0
transform 1 0 31188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 0
transform 1 0 828 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_6
timestamp 0
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_9
timestamp 0
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_13
timestamp 0
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_16
timestamp 0
transform 1 0 2024 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_19
timestamp 0
transform 1 0 2300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_22
timestamp 0
transform 1 0 2576 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_25
timestamp 0
transform 1 0 2852 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_38
timestamp 0
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_41
timestamp 0
transform 1 0 4324 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_44
timestamp 0
transform 1 0 4600 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_47
timestamp 0
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 0
transform 1 0 5796 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_64
timestamp 0
transform 1 0 6440 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_67
timestamp 0
transform 1 0 6716 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_70
timestamp 0
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_73
timestamp 0
transform 1 0 7268 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_87
timestamp 0
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_90
timestamp 0
transform 1 0 8832 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_98
timestamp 0
transform 1 0 9568 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_101
timestamp 0
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_113
timestamp 0
transform 1 0 10948 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_116
timestamp 0
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_119
timestamp 0
transform 1 0 11500 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_122
timestamp 0
transform 1 0 11776 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_128
timestamp 0
transform 1 0 12328 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_131
timestamp 0
transform 1 0 12604 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_134
timestamp 0
transform 1 0 12880 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_137
timestamp 0
transform 1 0 13156 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_153
timestamp 0
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_162
timestamp 0
transform 1 0 15456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 0
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_179
timestamp 0
transform 1 0 17020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_182
timestamp 0
transform 1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_185
timestamp 0
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_191
timestamp 0
transform 1 0 18124 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_194
timestamp 0
transform 1 0 18400 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_197
timestamp 0
transform 1 0 18676 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_200
timestamp 0
transform 1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_203
timestamp 0
transform 1 0 19228 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_206
timestamp 0
transform 1 0 19504 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_209
timestamp 0
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_212
timestamp 0
transform 1 0 20056 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_215
timestamp 0
transform 1 0 20332 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_218
timestamp 0
transform 1 0 20608 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_228
timestamp 0
transform 1 0 21528 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_231
timestamp 0
transform 1 0 21804 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_234
timestamp 0
transform 1 0 22080 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_237
timestamp 0
transform 1 0 22356 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_244
timestamp 0
transform 1 0 23000 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_247
timestamp 0
transform 1 0 23276 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 0
transform 1 0 26128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_281
timestamp 0
transform 1 0 26404 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_284
timestamp 0
transform 1 0 26680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_300
timestamp 0
transform 1 0 28152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_316
timestamp 0
transform 1 0 29624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_327
timestamp 0
transform 1 0 30636 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_3
timestamp 0
transform 1 0 828 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_6
timestamp 0
transform 1 0 1104 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_24
timestamp 0
transform 1 0 2760 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_29
timestamp 0
transform 1 0 3220 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_41
timestamp 0
transform 1 0 4324 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_44
timestamp 0
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_47
timestamp 0
transform 1 0 4876 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_52
timestamp 0
transform 1 0 5336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_55
timestamp 0
transform 1 0 5612 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_58
timestamp 0
transform 1 0 5888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_61
timestamp 0
transform 1 0 6164 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_67
timestamp 0
transform 1 0 6716 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_70
timestamp 0
transform 1 0 6992 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_73
timestamp 0
transform 1 0 7268 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_76
timestamp 0
transform 1 0 7544 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_93
timestamp 0
transform 1 0 9108 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_102
timestamp 0
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_110
timestamp 0
transform 1 0 10672 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_113
timestamp 0
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_116
timestamp 0
transform 1 0 11224 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 0
transform 1 0 13156 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 0
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_152
timestamp 0
transform 1 0 14536 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_155
timestamp 0
transform 1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_166
timestamp 0
transform 1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_169
timestamp 0
transform 1 0 16100 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_172
timestamp 0
transform 1 0 16376 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_175
timestamp 0
transform 1 0 16652 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_178
timestamp 0
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_181
timestamp 0
transform 1 0 17204 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_184
timestamp 0
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_187
timestamp 0
transform 1 0 17756 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_190
timestamp 0
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_193
timestamp 0
transform 1 0 18308 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_202
timestamp 0
transform 1 0 19136 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_212
timestamp 0
transform 1 0 20056 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_215
timestamp 0
transform 1 0 20332 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_218
timestamp 0
transform 1 0 20608 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_221
timestamp 0
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_233
timestamp 0
transform 1 0 21988 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_257
timestamp 0
transform 1 0 24196 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_281
timestamp 0
transform 1 0 26404 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_284
timestamp 0
transform 1 0 26680 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_288
timestamp 0
transform 1 0 27048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_294
timestamp 0
transform 1 0 27600 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_320
timestamp 0
transform 1 0 29992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_326
timestamp 0
transform 1 0 30544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_333
timestamp 0
transform 1 0 31188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_3
timestamp 0
transform 1 0 828 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_6
timestamp 0
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_9
timestamp 0
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_12
timestamp 0
transform 1 0 1656 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_15
timestamp 0
transform 1 0 1932 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_18
timestamp 0
transform 1 0 2208 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_21
timestamp 0
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_29
timestamp 0
transform 1 0 3220 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_32
timestamp 0
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_35
timestamp 0
transform 1 0 3772 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_38
timestamp 0
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_41
timestamp 0
transform 1 0 4324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_44
timestamp 0
transform 1 0 4600 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 0
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 0
transform 1 0 5796 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_64
timestamp 0
transform 1 0 6440 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_72
timestamp 0
transform 1 0 7176 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_75
timestamp 0
transform 1 0 7452 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_78
timestamp 0
transform 1 0 7728 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_86
timestamp 0
transform 1 0 8464 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_89
timestamp 0
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_92
timestamp 0
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_101
timestamp 0
transform 1 0 9844 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_104
timestamp 0
transform 1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_107
timestamp 0
transform 1 0 10396 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 0
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_113
timestamp 0
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_116
timestamp 0
transform 1 0 11224 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_134
timestamp 0
transform 1 0 12880 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_137
timestamp 0
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_146
timestamp 0
transform 1 0 13984 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_149
timestamp 0
transform 1 0 14260 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_152
timestamp 0
transform 1 0 14536 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_155
timestamp 0
transform 1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_158
timestamp 0
transform 1 0 15088 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_161
timestamp 0
transform 1 0 15364 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_186
timestamp 0
transform 1 0 17664 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_189
timestamp 0
transform 1 0 17940 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_192
timestamp 0
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_195
timestamp 0
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_200
timestamp 0
transform 1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_203
timestamp 0
transform 1 0 19228 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_206
timestamp 0
transform 1 0 19504 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_209
timestamp 0
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_212
timestamp 0
transform 1 0 20056 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_215
timestamp 0
transform 1 0 20332 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_3
timestamp 0
transform 1 0 828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_6
timestamp 0
transform 1 0 1104 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_11
timestamp 0
transform 1 0 1564 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_14
timestamp 0
transform 1 0 1840 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_23
timestamp 0
transform 1 0 2668 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 0
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_35
timestamp 0
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_42
timestamp 0
transform 1 0 4416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_45
timestamp 0
transform 1 0 4692 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_54
timestamp 0
transform 1 0 5520 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_57
timestamp 0
transform 1 0 5796 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_60
timestamp 0
transform 1 0 6072 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_63
timestamp 0
transform 1 0 6348 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_66
timestamp 0
transform 1 0 6624 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_75
timestamp 0
transform 1 0 7452 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_78
timestamp 0
transform 1 0 7728 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 0
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_90
timestamp 0
transform 1 0 8832 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_93
timestamp 0
transform 1 0 9108 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_96
timestamp 0
transform 1 0 9384 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_99
timestamp 0
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_109
timestamp 0
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_112
timestamp 0
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_115
timestamp 0
transform 1 0 11132 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_118
timestamp 0
transform 1 0 11408 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_127
timestamp 0
transform 1 0 12236 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_130
timestamp 0
transform 1 0 12512 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 0
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_144
timestamp 0
transform 1 0 13800 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_160
timestamp 0
transform 1 0 15272 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_163
timestamp 0
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_173
timestamp 0
transform 1 0 16468 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_176
timestamp 0
transform 1 0 16744 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_179
timestamp 0
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_186
timestamp 0
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_189
timestamp 0
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 0
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_215
timestamp 0
transform 1 0 20332 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_218
timestamp 0
transform 1 0 20608 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_221
timestamp 0
transform 1 0 20884 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_224
timestamp 0
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_333
timestamp 0
transform 1 0 31188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_3
timestamp 0
transform 1 0 828 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_6
timestamp 0
transform 1 0 1104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_34
timestamp 0
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_51
timestamp 0
transform 1 0 5244 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 0
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_64
timestamp 0
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_75
timestamp 0
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_113
timestamp 0
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_116
timestamp 0
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_119
timestamp 0
transform 1 0 11500 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_126
timestamp 0
transform 1 0 12144 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_129
timestamp 0
transform 1 0 12420 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_152
timestamp 0
transform 1 0 14536 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_155
timestamp 0
transform 1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_158
timestamp 0
transform 1 0 15088 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 15916 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_169
timestamp 0
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_172
timestamp 0
transform 1 0 16376 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_175
timestamp 0
transform 1 0 16652 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_178
timestamp 0
transform 1 0 16928 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_199
timestamp 0
transform 1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_202
timestamp 0
transform 1 0 19136 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_205
timestamp 0
transform 1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_208
timestamp 0
transform 1 0 19688 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_333
timestamp 0
transform 1 0 31188 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_3
timestamp 0
transform 1 0 828 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_6
timestamp 0
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_9
timestamp 0
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_17
timestamp 0
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 0
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_33
timestamp 0
transform 1 0 3588 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_36
timestamp 0
transform 1 0 3864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_39
timestamp 0
transform 1 0 4140 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_42
timestamp 0
transform 1 0 4416 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_45
timestamp 0
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_48
timestamp 0
transform 1 0 4968 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_51
timestamp 0
transform 1 0 5244 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_54
timestamp 0
transform 1 0 5520 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_78
timestamp 0
transform 1 0 7728 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 0
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 0
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_93
timestamp 0
transform 1 0 9108 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_96
timestamp 0
transform 1 0 9384 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_111
timestamp 0
transform 1 0 10764 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_124
timestamp 0
transform 1 0 11960 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_127
timestamp 0
transform 1 0 12236 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_130
timestamp 0
transform 1 0 12512 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_133
timestamp 0
transform 1 0 12788 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_144
timestamp 0
transform 1 0 13800 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_151
timestamp 0
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_176
timestamp 0
transform 1 0 16744 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_185
timestamp 0
transform 1 0 17572 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_188
timestamp 0
transform 1 0 17848 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_191
timestamp 0
transform 1 0 18124 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 0
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 0
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_220
timestamp 0
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 0
transform 1 0 23552 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_306
timestamp 0
transform 1 0 28704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_334
timestamp 0
transform 1 0 31280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_3
timestamp 0
transform 1 0 828 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_6
timestamp 0
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_9
timestamp 0
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_12
timestamp 0
transform 1 0 1656 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_15
timestamp 0
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_18
timestamp 0
transform 1 0 2208 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_21
timestamp 0
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_24
timestamp 0
transform 1 0 2760 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_27
timestamp 0
transform 1 0 3036 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_39
timestamp 0
transform 1 0 4140 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_43
timestamp 0
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_46
timestamp 0
transform 1 0 4784 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_52
timestamp 0
transform 1 0 5336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_62
timestamp 0
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_78
timestamp 0
transform 1 0 7728 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_81
timestamp 0
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_96
timestamp 0
transform 1 0 9384 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_99
timestamp 0
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 0
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 0
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_116
timestamp 0
transform 1 0 11224 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_122
timestamp 0
transform 1 0 11776 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_125
timestamp 0
transform 1 0 12052 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_134
timestamp 0
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_140
timestamp 0
transform 1 0 13432 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_143
timestamp 0
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_146
timestamp 0
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_149
timestamp 0
transform 1 0 14260 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_152
timestamp 0
transform 1 0 14536 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_155
timestamp 0
transform 1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_158
timestamp 0
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_197
timestamp 0
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_225
timestamp 0
transform 1 0 21252 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_243
timestamp 0
transform 1 0 22908 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26220 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_3
timestamp 0
transform 1 0 828 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_6
timestamp 0
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_9
timestamp 0
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_12
timestamp 0
transform 1 0 1656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_15
timestamp 0
transform 1 0 1932 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_18
timestamp 0
transform 1 0 2208 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_21
timestamp 0
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_24
timestamp 0
transform 1 0 2760 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3036 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_29
timestamp 0
transform 1 0 3220 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_32
timestamp 0
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_35
timestamp 0
transform 1 0 3772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_38
timestamp 0
transform 1 0 4048 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_41
timestamp 0
transform 1 0 4324 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_44
timestamp 0
transform 1 0 4600 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_47
timestamp 0
transform 1 0 4876 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_50
timestamp 0
transform 1 0 5152 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_53
timestamp 0
transform 1 0 5428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_56
timestamp 0
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_59
timestamp 0
transform 1 0 5980 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_65
timestamp 0
transform 1 0 6532 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_68
timestamp 0
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_71
timestamp 0
transform 1 0 7084 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_74
timestamp 0
transform 1 0 7360 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_77
timestamp 0
transform 1 0 7636 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_80
timestamp 0
transform 1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_91
timestamp 0
transform 1 0 8924 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_94
timestamp 0
transform 1 0 9200 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_97
timestamp 0
transform 1 0 9476 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_100
timestamp 0
transform 1 0 9752 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_103
timestamp 0
transform 1 0 10028 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_106
timestamp 0
transform 1 0 10304 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_109
timestamp 0
transform 1 0 10580 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_112
timestamp 0
transform 1 0 10856 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_115
timestamp 0
transform 1 0 11132 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_118
timestamp 0
transform 1 0 11408 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_121
timestamp 0
transform 1 0 11684 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_130
timestamp 0
transform 1 0 12512 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_133
timestamp 0
transform 1 0 12788 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_149
timestamp 0
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_152
timestamp 0
transform 1 0 14536 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_155
timestamp 0
transform 1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_158
timestamp 0
transform 1 0 15088 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_161
timestamp 0
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_164
timestamp 0
transform 1 0 15640 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_167
timestamp 0
transform 1 0 15916 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_170
timestamp 0
transform 1 0 16192 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_176
timestamp 0
transform 1 0 16744 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_179
timestamp 0
transform 1 0 17020 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_192
timestamp 0
transform 1 0 18216 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 18492 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_286
timestamp 0
transform 1 0 26864 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_334
timestamp 0
transform 1 0 31280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_3
timestamp 0
transform 1 0 828 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_6
timestamp 0
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_9
timestamp 0
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_12
timestamp 0
transform 1 0 1656 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_15
timestamp 0
transform 1 0 1932 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_18
timestamp 0
transform 1 0 2208 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_21
timestamp 0
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_24
timestamp 0
transform 1 0 2760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_27
timestamp 0
transform 1 0 3036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_30
timestamp 0
transform 1 0 3312 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_33
timestamp 0
transform 1 0 3588 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_36
timestamp 0
transform 1 0 3864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_39
timestamp 0
transform 1 0 4140 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_42
timestamp 0
transform 1 0 4416 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_45
timestamp 0
transform 1 0 4692 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_48
timestamp 0
transform 1 0 4968 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_51
timestamp 0
transform 1 0 5244 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 0
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_57
timestamp 0
transform 1 0 5796 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_60
timestamp 0
transform 1 0 6072 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_63
timestamp 0
transform 1 0 6348 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_66
timestamp 0
transform 1 0 6624 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_69
timestamp 0
transform 1 0 6900 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_113
timestamp 0
transform 1 0 10948 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_116
timestamp 0
transform 1 0 11224 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_122
timestamp 0
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_136
timestamp 0
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_152
timestamp 0
transform 1 0 14536 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_158
timestamp 0
transform 1 0 15088 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_161
timestamp 0
transform 1 0 15364 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_176
timestamp 0
transform 1 0 16744 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 0
transform 1 0 26128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_3
timestamp 0
transform 1 0 828 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_6
timestamp 0
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_9
timestamp 0
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_12
timestamp 0
transform 1 0 1656 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_15
timestamp 0
transform 1 0 1932 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_18
timestamp 0
transform 1 0 2208 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_21
timestamp 0
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_24
timestamp 0
transform 1 0 2760 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_29
timestamp 0
transform 1 0 3220 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_32
timestamp 0
transform 1 0 3496 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_35
timestamp 0
transform 1 0 3772 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_38
timestamp 0
transform 1 0 4048 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_41
timestamp 0
transform 1 0 4324 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_44
timestamp 0
transform 1 0 4600 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_47
timestamp 0
transform 1 0 4876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_50
timestamp 0
transform 1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_53
timestamp 0
transform 1 0 5428 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_56
timestamp 0
transform 1 0 5704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_59
timestamp 0
transform 1 0 5980 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_62
timestamp 0
transform 1 0 6256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_65
timestamp 0
transform 1 0 6532 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_68
timestamp 0
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_71
timestamp 0
transform 1 0 7084 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_74
timestamp 0
transform 1 0 7360 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_77
timestamp 0
transform 1 0 7636 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_85
timestamp 0
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_88
timestamp 0
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_103
timestamp 0
transform 1 0 10028 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_110
timestamp 0
transform 1 0 10672 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_141
timestamp 0
transform 1 0 13524 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_212
timestamp 0
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 0
transform 1 0 23552 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_3
timestamp 0
transform 1 0 828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_6
timestamp 0
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_9
timestamp 0
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_12
timestamp 0
transform 1 0 1656 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_15
timestamp 0
transform 1 0 1932 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_18
timestamp 0
transform 1 0 2208 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_21
timestamp 0
transform 1 0 2484 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_24
timestamp 0
transform 1 0 2760 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_27
timestamp 0
transform 1 0 3036 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_30
timestamp 0
transform 1 0 3312 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_33
timestamp 0
transform 1 0 3588 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_36
timestamp 0
transform 1 0 3864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_39
timestamp 0
transform 1 0 4140 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_42
timestamp 0
transform 1 0 4416 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_45
timestamp 0
transform 1 0 4692 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_48
timestamp 0
transform 1 0 4968 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_51
timestamp 0
transform 1 0 5244 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 0
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_57
timestamp 0
transform 1 0 5796 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_60
timestamp 0
transform 1 0 6072 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_63
timestamp 0
transform 1 0 6348 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_66
timestamp 0
transform 1 0 6624 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_69
timestamp 0
transform 1 0 6900 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_72
timestamp 0
transform 1 0 7176 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_75
timestamp 0
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_101
timestamp 0
transform 1 0 9844 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_104
timestamp 0
transform 1 0 10120 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_107
timestamp 0
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_139
timestamp 0
transform 1 0 13340 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_203
timestamp 0
transform 1 0 19228 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_258
timestamp 0
transform 1 0 24288 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_3
timestamp 0
transform 1 0 828 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_6
timestamp 0
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_9
timestamp 0
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_12
timestamp 0
transform 1 0 1656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_15
timestamp 0
transform 1 0 1932 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_18
timestamp 0
transform 1 0 2208 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_21
timestamp 0
transform 1 0 2484 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_24
timestamp 0
transform 1 0 2760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_29
timestamp 0
transform 1 0 3220 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_32
timestamp 0
transform 1 0 3496 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_35
timestamp 0
transform 1 0 3772 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_38
timestamp 0
transform 1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_41
timestamp 0
transform 1 0 4324 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_44
timestamp 0
transform 1 0 4600 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_47
timestamp 0
transform 1 0 4876 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_50
timestamp 0
transform 1 0 5152 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_53
timestamp 0
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_57
timestamp 0
transform 1 0 5796 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_60
timestamp 0
transform 1 0 6072 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_64
timestamp 0
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_70
timestamp 0
transform 1 0 6992 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_76
timestamp 0
transform 1 0 7544 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 0
transform 1 0 8096 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_88
timestamp 0
transform 1 0 8648 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_106
timestamp 0
transform 1 0 10304 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_126
timestamp 0
transform 1 0 12144 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_130
timestamp 0
transform 1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_136
timestamp 0
transform 1 0 13064 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 0
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_166
timestamp 0
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 18492 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_217
timestamp 0
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 0
transform 1 0 23552 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_253
timestamp 0
transform 1 0 23828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 20792 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 20056 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 9476 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 27140 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 30820 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 31096 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 26128 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 28612 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 22264 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform 1 0 27876 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 10028 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform -1 0 28704 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 30544 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap3
timestamp 0
transform 1 0 21988 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap7
timestamp 0
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap8
timestamp 0
transform -1 0 25024 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  max_cap9
timestamp 0
transform 1 0 6900 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap11
timestamp 0
transform -1 0 28060 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap13
timestamp 0
transform 1 0 3956 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 0
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 31648 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 0
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 31648 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 0
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 31648 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 0
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 31648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 0
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 0
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 31648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 0
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 0
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 31648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 0
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 31648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 0
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 31648 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 0
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 31648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 0
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 31648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 0
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 31648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 0
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 31648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 0
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 31648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 0
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 0
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 31648 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 0
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 0
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 31648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 0
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 31648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 0
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 31648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 0
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 31648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 0
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 31648 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 0
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 0
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 31648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 0
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 31648 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 0
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 31648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 0
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 31648 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 0
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 31648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 0
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 31648 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 0
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 31648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 0
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 31648 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 0
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 31648 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 0
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 31648 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 0
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 31648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 0
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 31648 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 0
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 31648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 0
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 31648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 0
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 0
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 0
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 0
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 0
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 0
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 0
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 0
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 0
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 0
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 0
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 0
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 0
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 0
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 0
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 0
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 0
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 0
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 0
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 0
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 0
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 0
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 0
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 0
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 0
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 0
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 0
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 0
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 0
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 0
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 0
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 0
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 0
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 0
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 0
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 0
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 0
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 0
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 0
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 0
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 0
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 0
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 0
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 0
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 0
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 0
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 0
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 0
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 0
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 0
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 0
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 0
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 0
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 0
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 0
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 0
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 0
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 0
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 0
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 0
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 0
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 0
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 0
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 0
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 0
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 0
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 0
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 0
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 0
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 0
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 0
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 0
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 0
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 0
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 0
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 0
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 0
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 0
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 0
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 0
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 0
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 0
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 0
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 0
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 0
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 0
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 0
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 0
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 0
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 0
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 0
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 0
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 0
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 0
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 0
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 0
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 0
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 0
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 0
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 0
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 0
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 0
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 0
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 0
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 0
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 0
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 0
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 0
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 0
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 0
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 0
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 0
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 0
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 0
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 0
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 0
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 0
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 0
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 0
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 0
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 0
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 0
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 0
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 0
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 0
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 0
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 0
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 0
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 0
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 0
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 0
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 0
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 0
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 0
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 0
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 0
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 0
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 0
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 0
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 0
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 0
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 0
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 0
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 0
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 0
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 0
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 0
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 0
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 0
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 0
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 0
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 0
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 0
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 0
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 0
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 0
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 0
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 0
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 0
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 0
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 0
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 0
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 0
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 0
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 0
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 0
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 0
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 0
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 0
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 0
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 0
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 0
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 0
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 0
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 0
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 0
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 0
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 0
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 0
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 0
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 0
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 0
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 0
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 0
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 0
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 0
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 0
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 0
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 0
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 0
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 0
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 0
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 0
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 0
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 0
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 0
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 0
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 0
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 0
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 0
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 0
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 0
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 0
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 0
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 0
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 0
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 0
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 0
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 0
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 0
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 0
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 0
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 0
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 0
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 0
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 0
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 0
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 0
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 0
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 0
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 0
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 0
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 0
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 0
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 0
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 0
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_121
timestamp 0
transform -1 0 10304 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_122
timestamp 0
transform -1 0 9752 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_123
timestamp 0
transform -1 0 10028 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_124
timestamp 0
transform -1 0 8648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_125
timestamp 0
transform -1 0 8096 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_126
timestamp 0
transform -1 0 7544 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_127
timestamp 0
transform -1 0 6992 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_128
timestamp 0
transform -1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_129
timestamp 0
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_130
timestamp 0
transform 1 0 13708 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_131
timestamp 0
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_132
timestamp 0
transform -1 0 13064 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_133
timestamp 0
transform -1 0 12512 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_134
timestamp 0
transform -1 0 12144 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_135
timestamp 0
transform 1 0 10948 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_136
timestamp 0
transform -1 0 10856 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_137
timestamp 0
transform -1 0 21528 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_138
timestamp 0
transform -1 0 18952 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_139
timestamp 0
transform 1 0 14628 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_140
timestamp 0
transform 1 0 16100 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_141
timestamp 0
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_142
timestamp 0
transform 1 0 14352 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_audio_player_143
timestamp 0
transform 1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  wire10
timestamp 0
transform 1 0 3036 0 -1 9248
box -38 -48 406 592
<< labels >>
flabel metal4 s 27638 496 27958 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 19864 496 20184 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12090 496 12410 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4316 496 4636 21808 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 26978 496 27298 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 19204 496 19524 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 11430 496 11750 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3656 496 3976 21808 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 28766 22104 28826 22304 0 FreeSans 600 90 0 0 clk
port 3 nsew
flabel metal4 s 29318 22104 29378 22304 0 FreeSans 600 90 0 0 ena
port 4 nsew
flabel metal4 s 28214 22104 28274 22304 0 FreeSans 600 90 0 0 rst_n
port 5 nsew
flabel metal4 s 27662 22104 27722 22304 0 FreeSans 600 90 0 0 ui_in[0]
port 6 nsew
flabel metal4 s 27110 22104 27170 22304 0 FreeSans 600 90 0 0 ui_in[1]
port 7 nsew
flabel metal4 s 26558 22104 26618 22304 0 FreeSans 600 90 0 0 ui_in[2]
port 8 nsew
flabel metal4 s 26006 22104 26066 22304 0 FreeSans 600 90 0 0 ui_in[3]
port 9 nsew
flabel metal4 s 25454 22104 25514 22304 0 FreeSans 600 90 0 0 ui_in[4]
port 10 nsew
flabel metal4 s 24902 22104 24962 22304 0 FreeSans 600 90 0 0 ui_in[5]
port 11 nsew
flabel metal4 s 24350 22104 24410 22304 0 FreeSans 600 90 0 0 ui_in[6]
port 12 nsew
flabel metal4 s 23798 22104 23858 22304 0 FreeSans 600 90 0 0 ui_in[7]
port 13 nsew
flabel metal4 s 23246 22104 23306 22304 0 FreeSans 600 90 0 0 uio_in[0]
port 14 nsew
flabel metal4 s 22694 22104 22754 22304 0 FreeSans 600 90 0 0 uio_in[1]
port 15 nsew
flabel metal4 s 22142 22104 22202 22304 0 FreeSans 600 90 0 0 uio_in[2]
port 16 nsew
flabel metal4 s 21590 22104 21650 22304 0 FreeSans 600 90 0 0 uio_in[3]
port 17 nsew
flabel metal4 s 21038 22104 21098 22304 0 FreeSans 600 90 0 0 uio_in[4]
port 18 nsew
flabel metal4 s 20486 22104 20546 22304 0 FreeSans 600 90 0 0 uio_in[5]
port 19 nsew
flabel metal4 s 19934 22104 19994 22304 0 FreeSans 600 90 0 0 uio_in[6]
port 20 nsew
flabel metal4 s 19382 22104 19442 22304 0 FreeSans 600 90 0 0 uio_in[7]
port 21 nsew
flabel metal4 s 9998 22104 10058 22304 0 FreeSans 600 90 0 0 uio_oe[0]
port 22 nsew
flabel metal4 s 9446 22104 9506 22304 0 FreeSans 600 90 0 0 uio_oe[1]
port 23 nsew
flabel metal4 s 8894 22104 8954 22304 0 FreeSans 600 90 0 0 uio_oe[2]
port 24 nsew
flabel metal4 s 8342 22104 8402 22304 0 FreeSans 600 90 0 0 uio_oe[3]
port 25 nsew
flabel metal4 s 7790 22104 7850 22304 0 FreeSans 600 90 0 0 uio_oe[4]
port 26 nsew
flabel metal4 s 7238 22104 7298 22304 0 FreeSans 600 90 0 0 uio_oe[5]
port 27 nsew
flabel metal4 s 6686 22104 6746 22304 0 FreeSans 600 90 0 0 uio_oe[6]
port 28 nsew
flabel metal4 s 6134 22104 6194 22304 0 FreeSans 600 90 0 0 uio_oe[7]
port 29 nsew
flabel metal4 s 14414 22104 14474 22304 0 FreeSans 600 90 0 0 uio_out[0]
port 30 nsew
flabel metal4 s 13862 22104 13922 22304 0 FreeSans 600 90 0 0 uio_out[1]
port 31 nsew
flabel metal4 s 13310 22104 13370 22304 0 FreeSans 600 90 0 0 uio_out[2]
port 32 nsew
flabel metal4 s 12758 22104 12818 22304 0 FreeSans 600 90 0 0 uio_out[3]
port 33 nsew
flabel metal4 s 12206 22104 12266 22304 0 FreeSans 600 90 0 0 uio_out[4]
port 34 nsew
flabel metal4 s 11654 22104 11714 22304 0 FreeSans 600 90 0 0 uio_out[5]
port 35 nsew
flabel metal4 s 11102 22104 11162 22304 0 FreeSans 600 90 0 0 uio_out[6]
port 36 nsew
flabel metal4 s 10550 22104 10610 22304 0 FreeSans 600 90 0 0 uio_out[7]
port 37 nsew
flabel metal4 s 18830 22104 18890 22304 0 FreeSans 600 90 0 0 uo_out[0]
port 38 nsew
flabel metal4 s 18278 22104 18338 22304 0 FreeSans 600 90 0 0 uo_out[1]
port 39 nsew
flabel metal4 s 17726 22104 17786 22304 0 FreeSans 600 90 0 0 uo_out[2]
port 40 nsew
flabel metal4 s 17174 22104 17234 22304 0 FreeSans 600 90 0 0 uo_out[3]
port 41 nsew
flabel metal4 s 16622 22104 16682 22304 0 FreeSans 600 90 0 0 uo_out[4]
port 42 nsew
flabel metal4 s 16070 22104 16130 22304 0 FreeSans 600 90 0 0 uo_out[5]
port 43 nsew
flabel metal4 s 15518 22104 15578 22304 0 FreeSans 600 90 0 0 uo_out[6]
port 44 nsew
flabel metal4 s 14966 22104 15026 22304 0 FreeSans 600 90 0 0 uo_out[7]
port 45 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 22304
<< end >>
