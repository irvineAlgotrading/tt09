magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -116 -66 219 666
<< mvpmos >>
rect 0 0 100 600
<< mvpdiff >>
rect -50 0 0 600
rect 100 0 150 600
<< poly >>
rect 0 600 100 626
rect 0 -26 100 0
<< locali >>
rect 111 -4 145 538
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_0
timestamp 1704896540
transform 1 0 100 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -25 300 -25 300 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87873666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87872782
<< end >>
