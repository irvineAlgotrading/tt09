magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 1900 9490 8579 39520
rect 1900 3303 7883 9490
<< nwell >>
rect 1820 39246 8659 39600
rect 1820 9764 2174 39246
rect 8305 9764 8659 39246
rect 1820 9528 8659 9764
rect 1820 3577 2174 9528
rect 7609 9410 8659 9528
rect 7609 3577 7963 9410
rect 1820 3223 7963 3577
rect 1734 797 5106 2083
<< pwell >>
rect 2248 38946 8245 39168
rect 2248 9945 2470 38946
rect 2678 17098 4718 29008
rect 8023 17098 8245 38946
rect 2678 15886 8245 17098
rect 8023 9945 8245 15886
rect 2248 9859 8245 9945
rect 2254 9370 7547 9456
rect 2254 7707 2360 9370
rect 7461 7707 7547 9370
rect 2254 7621 7547 7707
rect 2254 5867 2360 7621
rect 7461 5867 7547 7621
rect 2254 5781 7547 5867
rect 2254 3956 2360 5781
rect 7461 3956 7547 5781
rect 2254 3824 7547 3956
rect 1805 2369 7930 3153
rect 5314 326 7620 2369
<< psubdiff >>
rect 2274 39108 2405 39142
rect 2439 39108 2473 39142
rect 2274 39074 2473 39108
rect 2376 39040 2473 39074
rect 8151 39040 8219 39142
rect 2376 39006 2541 39040
rect 2444 38972 2541 39006
rect 8083 39023 8219 39040
rect 8083 38989 8185 39023
rect 8083 38972 8219 38989
rect 8049 38955 8219 38972
rect 8049 38887 8117 38955
rect 2704 28958 4692 28982
rect 2704 28924 2715 28958
rect 2749 28924 2853 28958
rect 2887 28924 2991 28958
rect 3025 28924 3129 28958
rect 3163 28924 3267 28958
rect 3301 28924 3405 28958
rect 3439 28924 3543 28958
rect 3577 28924 3681 28958
rect 3715 28924 3819 28958
rect 3853 28924 3957 28958
rect 3991 28924 4095 28958
rect 4129 28924 4233 28958
rect 4267 28924 4371 28958
rect 4405 28924 4509 28958
rect 4543 28924 4647 28958
rect 4681 28924 4692 28958
rect 2704 28822 4692 28924
rect 2704 28788 2715 28822
rect 2749 28788 2853 28822
rect 2887 28788 2991 28822
rect 3025 28788 3129 28822
rect 3163 28788 3267 28822
rect 3301 28788 3405 28822
rect 3439 28788 3543 28822
rect 3577 28788 3681 28822
rect 3715 28788 3819 28822
rect 3853 28788 3957 28822
rect 3991 28788 4095 28822
rect 4129 28788 4233 28822
rect 4267 28788 4371 28822
rect 4405 28788 4509 28822
rect 4543 28788 4647 28822
rect 4681 28788 4692 28822
rect 2704 28686 4692 28788
rect 2704 28652 2715 28686
rect 2749 28652 2853 28686
rect 2887 28652 2991 28686
rect 3025 28652 3129 28686
rect 3163 28652 3267 28686
rect 3301 28652 3405 28686
rect 3439 28652 3543 28686
rect 3577 28652 3681 28686
rect 3715 28652 3819 28686
rect 3853 28652 3957 28686
rect 3991 28652 4095 28686
rect 4129 28652 4233 28686
rect 4267 28652 4371 28686
rect 4405 28652 4509 28686
rect 4543 28652 4647 28686
rect 4681 28652 4692 28686
rect 2704 28550 4692 28652
rect 2704 28516 2715 28550
rect 2749 28516 2853 28550
rect 2887 28516 2991 28550
rect 3025 28516 3129 28550
rect 3163 28516 3267 28550
rect 3301 28516 3405 28550
rect 3439 28516 3543 28550
rect 3577 28516 3681 28550
rect 3715 28516 3819 28550
rect 3853 28516 3957 28550
rect 3991 28516 4095 28550
rect 4129 28516 4233 28550
rect 4267 28516 4371 28550
rect 4405 28516 4509 28550
rect 4543 28516 4647 28550
rect 4681 28516 4692 28550
rect 2704 28414 4692 28516
rect 2704 28380 2715 28414
rect 2749 28380 2853 28414
rect 2887 28380 2991 28414
rect 3025 28380 3129 28414
rect 3163 28380 3267 28414
rect 3301 28380 3405 28414
rect 3439 28380 3543 28414
rect 3577 28380 3681 28414
rect 3715 28380 3819 28414
rect 3853 28380 3957 28414
rect 3991 28380 4095 28414
rect 4129 28380 4233 28414
rect 4267 28380 4371 28414
rect 4405 28380 4509 28414
rect 4543 28380 4647 28414
rect 4681 28380 4692 28414
rect 2704 28278 4692 28380
rect 2704 28244 2715 28278
rect 2749 28244 2853 28278
rect 2887 28244 2991 28278
rect 3025 28244 3129 28278
rect 3163 28244 3267 28278
rect 3301 28244 3405 28278
rect 3439 28244 3543 28278
rect 3577 28244 3681 28278
rect 3715 28244 3819 28278
rect 3853 28244 3957 28278
rect 3991 28244 4095 28278
rect 4129 28244 4233 28278
rect 4267 28244 4371 28278
rect 4405 28244 4509 28278
rect 4543 28244 4647 28278
rect 4681 28244 4692 28278
rect 2704 28142 4692 28244
rect 2704 28108 2715 28142
rect 2749 28108 2853 28142
rect 2887 28108 2991 28142
rect 3025 28108 3129 28142
rect 3163 28108 3267 28142
rect 3301 28108 3405 28142
rect 3439 28108 3543 28142
rect 3577 28108 3681 28142
rect 3715 28108 3819 28142
rect 3853 28108 3957 28142
rect 3991 28108 4095 28142
rect 4129 28108 4233 28142
rect 4267 28108 4371 28142
rect 4405 28108 4509 28142
rect 4543 28108 4647 28142
rect 4681 28108 4692 28142
rect 2704 28006 4692 28108
rect 2704 27972 2715 28006
rect 2749 27972 2853 28006
rect 2887 27972 2991 28006
rect 3025 27972 3129 28006
rect 3163 27972 3267 28006
rect 3301 27972 3405 28006
rect 3439 27972 3543 28006
rect 3577 27972 3681 28006
rect 3715 27972 3819 28006
rect 3853 27972 3957 28006
rect 3991 27972 4095 28006
rect 4129 27972 4233 28006
rect 4267 27972 4371 28006
rect 4405 27972 4509 28006
rect 4543 27972 4647 28006
rect 4681 27972 4692 28006
rect 2704 27870 4692 27972
rect 2704 27836 2715 27870
rect 2749 27836 2853 27870
rect 2887 27836 2991 27870
rect 3025 27836 3129 27870
rect 3163 27836 3267 27870
rect 3301 27836 3405 27870
rect 3439 27836 3543 27870
rect 3577 27836 3681 27870
rect 3715 27836 3819 27870
rect 3853 27836 3957 27870
rect 3991 27836 4095 27870
rect 4129 27836 4233 27870
rect 4267 27836 4371 27870
rect 4405 27836 4509 27870
rect 4543 27836 4647 27870
rect 4681 27836 4692 27870
rect 2704 27734 4692 27836
rect 2704 27700 2715 27734
rect 2749 27700 2853 27734
rect 2887 27700 2991 27734
rect 3025 27700 3129 27734
rect 3163 27700 3267 27734
rect 3301 27700 3405 27734
rect 3439 27700 3543 27734
rect 3577 27700 3681 27734
rect 3715 27700 3819 27734
rect 3853 27700 3957 27734
rect 3991 27700 4095 27734
rect 4129 27700 4233 27734
rect 4267 27700 4371 27734
rect 4405 27700 4509 27734
rect 4543 27700 4647 27734
rect 4681 27700 4692 27734
rect 2704 27598 4692 27700
rect 2704 27564 2715 27598
rect 2749 27564 2853 27598
rect 2887 27564 2991 27598
rect 3025 27564 3129 27598
rect 3163 27564 3267 27598
rect 3301 27564 3405 27598
rect 3439 27564 3543 27598
rect 3577 27564 3681 27598
rect 3715 27564 3819 27598
rect 3853 27564 3957 27598
rect 3991 27564 4095 27598
rect 4129 27564 4233 27598
rect 4267 27564 4371 27598
rect 4405 27564 4509 27598
rect 4543 27564 4647 27598
rect 4681 27564 4692 27598
rect 2704 27462 4692 27564
rect 2704 27428 2715 27462
rect 2749 27428 2853 27462
rect 2887 27428 2991 27462
rect 3025 27428 3129 27462
rect 3163 27428 3267 27462
rect 3301 27428 3405 27462
rect 3439 27428 3543 27462
rect 3577 27428 3681 27462
rect 3715 27428 3819 27462
rect 3853 27428 3957 27462
rect 3991 27428 4095 27462
rect 4129 27428 4233 27462
rect 4267 27428 4371 27462
rect 4405 27428 4509 27462
rect 4543 27428 4647 27462
rect 4681 27428 4692 27462
rect 2704 27326 4692 27428
rect 2704 27292 2715 27326
rect 2749 27292 2853 27326
rect 2887 27292 2991 27326
rect 3025 27292 3129 27326
rect 3163 27292 3267 27326
rect 3301 27292 3405 27326
rect 3439 27292 3543 27326
rect 3577 27292 3681 27326
rect 3715 27292 3819 27326
rect 3853 27292 3957 27326
rect 3991 27292 4095 27326
rect 4129 27292 4233 27326
rect 4267 27292 4371 27326
rect 4405 27292 4509 27326
rect 4543 27292 4647 27326
rect 4681 27292 4692 27326
rect 2704 27190 4692 27292
rect 2704 27156 2715 27190
rect 2749 27156 2853 27190
rect 2887 27156 2991 27190
rect 3025 27156 3129 27190
rect 3163 27156 3267 27190
rect 3301 27156 3405 27190
rect 3439 27156 3543 27190
rect 3577 27156 3681 27190
rect 3715 27156 3819 27190
rect 3853 27156 3957 27190
rect 3991 27156 4095 27190
rect 4129 27156 4233 27190
rect 4267 27156 4371 27190
rect 4405 27156 4509 27190
rect 4543 27156 4647 27190
rect 4681 27156 4692 27190
rect 2704 27054 4692 27156
rect 2704 27020 2715 27054
rect 2749 27020 2853 27054
rect 2887 27020 2991 27054
rect 3025 27020 3129 27054
rect 3163 27020 3267 27054
rect 3301 27020 3405 27054
rect 3439 27020 3543 27054
rect 3577 27020 3681 27054
rect 3715 27020 3819 27054
rect 3853 27020 3957 27054
rect 3991 27020 4095 27054
rect 4129 27020 4233 27054
rect 4267 27020 4371 27054
rect 4405 27020 4509 27054
rect 4543 27020 4647 27054
rect 4681 27020 4692 27054
rect 2704 26918 4692 27020
rect 2704 26884 2715 26918
rect 2749 26884 2853 26918
rect 2887 26884 2991 26918
rect 3025 26884 3129 26918
rect 3163 26884 3267 26918
rect 3301 26884 3405 26918
rect 3439 26884 3543 26918
rect 3577 26884 3681 26918
rect 3715 26884 3819 26918
rect 3853 26884 3957 26918
rect 3991 26884 4095 26918
rect 4129 26884 4233 26918
rect 4267 26884 4371 26918
rect 4405 26884 4509 26918
rect 4543 26884 4647 26918
rect 4681 26884 4692 26918
rect 2704 26782 4692 26884
rect 2704 26748 2715 26782
rect 2749 26748 2853 26782
rect 2887 26748 2991 26782
rect 3025 26748 3129 26782
rect 3163 26748 3267 26782
rect 3301 26748 3405 26782
rect 3439 26748 3543 26782
rect 3577 26748 3681 26782
rect 3715 26748 3819 26782
rect 3853 26748 3957 26782
rect 3991 26748 4095 26782
rect 4129 26748 4233 26782
rect 4267 26748 4371 26782
rect 4405 26748 4509 26782
rect 4543 26748 4647 26782
rect 4681 26748 4692 26782
rect 2704 26646 4692 26748
rect 2704 26612 2715 26646
rect 2749 26612 2853 26646
rect 2887 26612 2991 26646
rect 3025 26612 3129 26646
rect 3163 26612 3267 26646
rect 3301 26612 3405 26646
rect 3439 26612 3543 26646
rect 3577 26612 3681 26646
rect 3715 26612 3819 26646
rect 3853 26612 3957 26646
rect 3991 26612 4095 26646
rect 4129 26612 4233 26646
rect 4267 26612 4371 26646
rect 4405 26612 4509 26646
rect 4543 26612 4647 26646
rect 4681 26612 4692 26646
rect 2704 26510 4692 26612
rect 2704 26476 2715 26510
rect 2749 26476 2853 26510
rect 2887 26476 2991 26510
rect 3025 26476 3129 26510
rect 3163 26476 3267 26510
rect 3301 26476 3405 26510
rect 3439 26476 3543 26510
rect 3577 26476 3681 26510
rect 3715 26476 3819 26510
rect 3853 26476 3957 26510
rect 3991 26476 4095 26510
rect 4129 26476 4233 26510
rect 4267 26476 4371 26510
rect 4405 26476 4509 26510
rect 4543 26476 4647 26510
rect 4681 26476 4692 26510
rect 2704 26374 4692 26476
rect 2704 26340 2715 26374
rect 2749 26340 2853 26374
rect 2887 26340 2991 26374
rect 3025 26340 3129 26374
rect 3163 26340 3267 26374
rect 3301 26340 3405 26374
rect 3439 26340 3543 26374
rect 3577 26340 3681 26374
rect 3715 26340 3819 26374
rect 3853 26340 3957 26374
rect 3991 26340 4095 26374
rect 4129 26340 4233 26374
rect 4267 26340 4371 26374
rect 4405 26340 4509 26374
rect 4543 26340 4647 26374
rect 4681 26340 4692 26374
rect 2704 26238 4692 26340
rect 2704 26204 2715 26238
rect 2749 26204 2853 26238
rect 2887 26204 2991 26238
rect 3025 26204 3129 26238
rect 3163 26204 3267 26238
rect 3301 26204 3405 26238
rect 3439 26204 3543 26238
rect 3577 26204 3681 26238
rect 3715 26204 3819 26238
rect 3853 26204 3957 26238
rect 3991 26204 4095 26238
rect 4129 26204 4233 26238
rect 4267 26204 4371 26238
rect 4405 26204 4509 26238
rect 4543 26204 4647 26238
rect 4681 26204 4692 26238
rect 2704 26102 4692 26204
rect 2704 26068 2715 26102
rect 2749 26068 2853 26102
rect 2887 26068 2991 26102
rect 3025 26068 3129 26102
rect 3163 26068 3267 26102
rect 3301 26068 3405 26102
rect 3439 26068 3543 26102
rect 3577 26068 3681 26102
rect 3715 26068 3819 26102
rect 3853 26068 3957 26102
rect 3991 26068 4095 26102
rect 4129 26068 4233 26102
rect 4267 26068 4371 26102
rect 4405 26068 4509 26102
rect 4543 26068 4647 26102
rect 4681 26068 4692 26102
rect 2704 25966 4692 26068
rect 2704 25932 2715 25966
rect 2749 25932 2853 25966
rect 2887 25932 2991 25966
rect 3025 25932 3129 25966
rect 3163 25932 3267 25966
rect 3301 25932 3405 25966
rect 3439 25932 3543 25966
rect 3577 25932 3681 25966
rect 3715 25932 3819 25966
rect 3853 25932 3957 25966
rect 3991 25932 4095 25966
rect 4129 25932 4233 25966
rect 4267 25932 4371 25966
rect 4405 25932 4509 25966
rect 4543 25932 4647 25966
rect 4681 25932 4692 25966
rect 2704 25830 4692 25932
rect 2704 25796 2715 25830
rect 2749 25796 2853 25830
rect 2887 25796 2991 25830
rect 3025 25796 3129 25830
rect 3163 25796 3267 25830
rect 3301 25796 3405 25830
rect 3439 25796 3543 25830
rect 3577 25796 3681 25830
rect 3715 25796 3819 25830
rect 3853 25796 3957 25830
rect 3991 25796 4095 25830
rect 4129 25796 4233 25830
rect 4267 25796 4371 25830
rect 4405 25796 4509 25830
rect 4543 25796 4647 25830
rect 4681 25796 4692 25830
rect 2704 25694 4692 25796
rect 2704 25660 2715 25694
rect 2749 25660 2853 25694
rect 2887 25660 2991 25694
rect 3025 25660 3129 25694
rect 3163 25660 3267 25694
rect 3301 25660 3405 25694
rect 3439 25660 3543 25694
rect 3577 25660 3681 25694
rect 3715 25660 3819 25694
rect 3853 25660 3957 25694
rect 3991 25660 4095 25694
rect 4129 25660 4233 25694
rect 4267 25660 4371 25694
rect 4405 25660 4509 25694
rect 4543 25660 4647 25694
rect 4681 25660 4692 25694
rect 2704 25558 4692 25660
rect 2704 25524 2715 25558
rect 2749 25524 2853 25558
rect 2887 25524 2991 25558
rect 3025 25524 3129 25558
rect 3163 25524 3267 25558
rect 3301 25524 3405 25558
rect 3439 25524 3543 25558
rect 3577 25524 3681 25558
rect 3715 25524 3819 25558
rect 3853 25524 3957 25558
rect 3991 25524 4095 25558
rect 4129 25524 4233 25558
rect 4267 25524 4371 25558
rect 4405 25524 4509 25558
rect 4543 25524 4647 25558
rect 4681 25524 4692 25558
rect 2704 25422 4692 25524
rect 2704 25388 2715 25422
rect 2749 25388 2853 25422
rect 2887 25388 2991 25422
rect 3025 25388 3129 25422
rect 3163 25388 3267 25422
rect 3301 25388 3405 25422
rect 3439 25388 3543 25422
rect 3577 25388 3681 25422
rect 3715 25388 3819 25422
rect 3853 25388 3957 25422
rect 3991 25388 4095 25422
rect 4129 25388 4233 25422
rect 4267 25388 4371 25422
rect 4405 25388 4509 25422
rect 4543 25388 4647 25422
rect 4681 25388 4692 25422
rect 2704 25286 4692 25388
rect 2704 25252 2715 25286
rect 2749 25252 2853 25286
rect 2887 25252 2991 25286
rect 3025 25252 3129 25286
rect 3163 25252 3267 25286
rect 3301 25252 3405 25286
rect 3439 25252 3543 25286
rect 3577 25252 3681 25286
rect 3715 25252 3819 25286
rect 3853 25252 3957 25286
rect 3991 25252 4095 25286
rect 4129 25252 4233 25286
rect 4267 25252 4371 25286
rect 4405 25252 4509 25286
rect 4543 25252 4647 25286
rect 4681 25252 4692 25286
rect 2704 25149 4692 25252
rect 2704 25115 2715 25149
rect 2749 25115 2853 25149
rect 2887 25115 2991 25149
rect 3025 25115 3129 25149
rect 3163 25115 3267 25149
rect 3301 25115 3405 25149
rect 3439 25115 3543 25149
rect 3577 25115 3681 25149
rect 3715 25115 3819 25149
rect 3853 25115 3957 25149
rect 3991 25115 4095 25149
rect 4129 25115 4233 25149
rect 4267 25115 4371 25149
rect 4405 25115 4509 25149
rect 4543 25115 4647 25149
rect 4681 25115 4692 25149
rect 2704 25012 4692 25115
rect 2704 24978 2715 25012
rect 2749 24978 2853 25012
rect 2887 24978 2991 25012
rect 3025 24978 3129 25012
rect 3163 24978 3267 25012
rect 3301 24978 3405 25012
rect 3439 24978 3543 25012
rect 3577 24978 3681 25012
rect 3715 24978 3819 25012
rect 3853 24978 3957 25012
rect 3991 24978 4095 25012
rect 4129 24978 4233 25012
rect 4267 24978 4371 25012
rect 4405 24978 4509 25012
rect 4543 24978 4647 25012
rect 4681 24978 4692 25012
rect 2704 24875 4692 24978
rect 2704 24841 2715 24875
rect 2749 24841 2853 24875
rect 2887 24841 2991 24875
rect 3025 24841 3129 24875
rect 3163 24841 3267 24875
rect 3301 24841 3405 24875
rect 3439 24841 3543 24875
rect 3577 24841 3681 24875
rect 3715 24841 3819 24875
rect 3853 24841 3957 24875
rect 3991 24841 4095 24875
rect 4129 24841 4233 24875
rect 4267 24841 4371 24875
rect 4405 24841 4509 24875
rect 4543 24841 4647 24875
rect 4681 24841 4692 24875
rect 2704 24738 4692 24841
rect 2704 24704 2715 24738
rect 2749 24704 2853 24738
rect 2887 24704 2991 24738
rect 3025 24704 3129 24738
rect 3163 24704 3267 24738
rect 3301 24704 3405 24738
rect 3439 24704 3543 24738
rect 3577 24704 3681 24738
rect 3715 24704 3819 24738
rect 3853 24704 3957 24738
rect 3991 24704 4095 24738
rect 4129 24704 4233 24738
rect 4267 24704 4371 24738
rect 4405 24704 4509 24738
rect 4543 24704 4647 24738
rect 4681 24704 4692 24738
rect 2704 24601 4692 24704
rect 2704 24567 2715 24601
rect 2749 24567 2853 24601
rect 2887 24567 2991 24601
rect 3025 24567 3129 24601
rect 3163 24567 3267 24601
rect 3301 24567 3405 24601
rect 3439 24567 3543 24601
rect 3577 24567 3681 24601
rect 3715 24567 3819 24601
rect 3853 24567 3957 24601
rect 3991 24567 4095 24601
rect 4129 24567 4233 24601
rect 4267 24567 4371 24601
rect 4405 24567 4509 24601
rect 4543 24567 4647 24601
rect 4681 24567 4692 24601
rect 2704 24464 4692 24567
rect 2704 24430 2715 24464
rect 2749 24430 2853 24464
rect 2887 24430 2991 24464
rect 3025 24430 3129 24464
rect 3163 24430 3267 24464
rect 3301 24430 3405 24464
rect 3439 24430 3543 24464
rect 3577 24430 3681 24464
rect 3715 24430 3819 24464
rect 3853 24430 3957 24464
rect 3991 24430 4095 24464
rect 4129 24430 4233 24464
rect 4267 24430 4371 24464
rect 4405 24430 4509 24464
rect 4543 24430 4647 24464
rect 4681 24430 4692 24464
rect 2704 24327 4692 24430
rect 2704 24293 2715 24327
rect 2749 24293 2853 24327
rect 2887 24293 2991 24327
rect 3025 24293 3129 24327
rect 3163 24293 3267 24327
rect 3301 24293 3405 24327
rect 3439 24293 3543 24327
rect 3577 24293 3681 24327
rect 3715 24293 3819 24327
rect 3853 24293 3957 24327
rect 3991 24293 4095 24327
rect 4129 24293 4233 24327
rect 4267 24293 4371 24327
rect 4405 24293 4509 24327
rect 4543 24293 4647 24327
rect 4681 24293 4692 24327
rect 2704 24190 4692 24293
rect 2704 24156 2715 24190
rect 2749 24156 2853 24190
rect 2887 24156 2991 24190
rect 3025 24156 3129 24190
rect 3163 24156 3267 24190
rect 3301 24156 3405 24190
rect 3439 24156 3543 24190
rect 3577 24156 3681 24190
rect 3715 24156 3819 24190
rect 3853 24156 3957 24190
rect 3991 24156 4095 24190
rect 4129 24156 4233 24190
rect 4267 24156 4371 24190
rect 4405 24156 4509 24190
rect 4543 24156 4647 24190
rect 4681 24156 4692 24190
rect 2704 24053 4692 24156
rect 2704 24019 2715 24053
rect 2749 24019 2853 24053
rect 2887 24019 2991 24053
rect 3025 24019 3129 24053
rect 3163 24019 3267 24053
rect 3301 24019 3405 24053
rect 3439 24019 3543 24053
rect 3577 24019 3681 24053
rect 3715 24019 3819 24053
rect 3853 24019 3957 24053
rect 3991 24019 4095 24053
rect 4129 24019 4233 24053
rect 4267 24019 4371 24053
rect 4405 24019 4509 24053
rect 4543 24019 4647 24053
rect 4681 24019 4692 24053
rect 2704 23916 4692 24019
rect 2704 23882 2715 23916
rect 2749 23882 2853 23916
rect 2887 23882 2991 23916
rect 3025 23882 3129 23916
rect 3163 23882 3267 23916
rect 3301 23882 3405 23916
rect 3439 23882 3543 23916
rect 3577 23882 3681 23916
rect 3715 23882 3819 23916
rect 3853 23882 3957 23916
rect 3991 23882 4095 23916
rect 4129 23882 4233 23916
rect 4267 23882 4371 23916
rect 4405 23882 4509 23916
rect 4543 23882 4647 23916
rect 4681 23882 4692 23916
rect 2704 23779 4692 23882
rect 2704 23745 2715 23779
rect 2749 23745 2853 23779
rect 2887 23745 2991 23779
rect 3025 23745 3129 23779
rect 3163 23745 3267 23779
rect 3301 23745 3405 23779
rect 3439 23745 3543 23779
rect 3577 23745 3681 23779
rect 3715 23745 3819 23779
rect 3853 23745 3957 23779
rect 3991 23745 4095 23779
rect 4129 23745 4233 23779
rect 4267 23745 4371 23779
rect 4405 23745 4509 23779
rect 4543 23745 4647 23779
rect 4681 23745 4692 23779
rect 2704 23642 4692 23745
rect 2704 23608 2715 23642
rect 2749 23608 2853 23642
rect 2887 23608 2991 23642
rect 3025 23608 3129 23642
rect 3163 23608 3267 23642
rect 3301 23608 3405 23642
rect 3439 23608 3543 23642
rect 3577 23608 3681 23642
rect 3715 23608 3819 23642
rect 3853 23608 3957 23642
rect 3991 23608 4095 23642
rect 4129 23608 4233 23642
rect 4267 23608 4371 23642
rect 4405 23608 4509 23642
rect 4543 23608 4647 23642
rect 4681 23608 4692 23642
rect 2704 23505 4692 23608
rect 2704 23471 2715 23505
rect 2749 23471 2853 23505
rect 2887 23471 2991 23505
rect 3025 23471 3129 23505
rect 3163 23471 3267 23505
rect 3301 23471 3405 23505
rect 3439 23471 3543 23505
rect 3577 23471 3681 23505
rect 3715 23471 3819 23505
rect 3853 23471 3957 23505
rect 3991 23471 4095 23505
rect 4129 23471 4233 23505
rect 4267 23471 4371 23505
rect 4405 23471 4509 23505
rect 4543 23471 4647 23505
rect 4681 23471 4692 23505
rect 2704 23368 4692 23471
rect 2704 23334 2715 23368
rect 2749 23334 2853 23368
rect 2887 23334 2991 23368
rect 3025 23334 3129 23368
rect 3163 23334 3267 23368
rect 3301 23334 3405 23368
rect 3439 23334 3543 23368
rect 3577 23334 3681 23368
rect 3715 23334 3819 23368
rect 3853 23334 3957 23368
rect 3991 23334 4095 23368
rect 4129 23334 4233 23368
rect 4267 23334 4371 23368
rect 4405 23334 4509 23368
rect 4543 23334 4647 23368
rect 4681 23334 4692 23368
rect 2704 23231 4692 23334
rect 2704 23197 2715 23231
rect 2749 23197 2853 23231
rect 2887 23197 2991 23231
rect 3025 23197 3129 23231
rect 3163 23197 3267 23231
rect 3301 23197 3405 23231
rect 3439 23197 3543 23231
rect 3577 23197 3681 23231
rect 3715 23197 3819 23231
rect 3853 23197 3957 23231
rect 3991 23197 4095 23231
rect 4129 23197 4233 23231
rect 4267 23197 4371 23231
rect 4405 23197 4509 23231
rect 4543 23197 4647 23231
rect 4681 23197 4692 23231
rect 2704 23094 4692 23197
rect 2704 23060 2715 23094
rect 2749 23060 2853 23094
rect 2887 23060 2991 23094
rect 3025 23060 3129 23094
rect 3163 23060 3267 23094
rect 3301 23060 3405 23094
rect 3439 23060 3543 23094
rect 3577 23060 3681 23094
rect 3715 23060 3819 23094
rect 3853 23060 3957 23094
rect 3991 23060 4095 23094
rect 4129 23060 4233 23094
rect 4267 23060 4371 23094
rect 4405 23060 4509 23094
rect 4543 23060 4647 23094
rect 4681 23060 4692 23094
rect 2704 22957 4692 23060
rect 2704 22923 2715 22957
rect 2749 22923 2853 22957
rect 2887 22923 2991 22957
rect 3025 22923 3129 22957
rect 3163 22923 3267 22957
rect 3301 22923 3405 22957
rect 3439 22923 3543 22957
rect 3577 22923 3681 22957
rect 3715 22923 3819 22957
rect 3853 22923 3957 22957
rect 3991 22923 4095 22957
rect 4129 22923 4233 22957
rect 4267 22923 4371 22957
rect 4405 22923 4509 22957
rect 4543 22923 4647 22957
rect 4681 22923 4692 22957
rect 2704 22820 4692 22923
rect 2704 22786 2715 22820
rect 2749 22786 2853 22820
rect 2887 22786 2991 22820
rect 3025 22786 3129 22820
rect 3163 22786 3267 22820
rect 3301 22786 3405 22820
rect 3439 22786 3543 22820
rect 3577 22786 3681 22820
rect 3715 22786 3819 22820
rect 3853 22786 3957 22820
rect 3991 22786 4095 22820
rect 4129 22786 4233 22820
rect 4267 22786 4371 22820
rect 4405 22786 4509 22820
rect 4543 22786 4647 22820
rect 4681 22786 4692 22820
rect 2704 22683 4692 22786
rect 2704 22649 2715 22683
rect 2749 22649 2853 22683
rect 2887 22649 2991 22683
rect 3025 22649 3129 22683
rect 3163 22649 3267 22683
rect 3301 22649 3405 22683
rect 3439 22649 3543 22683
rect 3577 22649 3681 22683
rect 3715 22649 3819 22683
rect 3853 22649 3957 22683
rect 3991 22649 4095 22683
rect 4129 22649 4233 22683
rect 4267 22649 4371 22683
rect 4405 22649 4509 22683
rect 4543 22649 4647 22683
rect 4681 22649 4692 22683
rect 2704 22546 4692 22649
rect 2704 22512 2715 22546
rect 2749 22512 2853 22546
rect 2887 22512 2991 22546
rect 3025 22512 3129 22546
rect 3163 22512 3267 22546
rect 3301 22512 3405 22546
rect 3439 22512 3543 22546
rect 3577 22512 3681 22546
rect 3715 22512 3819 22546
rect 3853 22512 3957 22546
rect 3991 22512 4095 22546
rect 4129 22512 4233 22546
rect 4267 22512 4371 22546
rect 4405 22512 4509 22546
rect 4543 22512 4647 22546
rect 4681 22512 4692 22546
rect 2704 22409 4692 22512
rect 2704 22375 2715 22409
rect 2749 22375 2853 22409
rect 2887 22375 2991 22409
rect 3025 22375 3129 22409
rect 3163 22375 3267 22409
rect 3301 22375 3405 22409
rect 3439 22375 3543 22409
rect 3577 22375 3681 22409
rect 3715 22375 3819 22409
rect 3853 22375 3957 22409
rect 3991 22375 4095 22409
rect 4129 22375 4233 22409
rect 4267 22375 4371 22409
rect 4405 22375 4509 22409
rect 4543 22375 4647 22409
rect 4681 22375 4692 22409
rect 2704 22272 4692 22375
rect 2704 22238 2715 22272
rect 2749 22238 2853 22272
rect 2887 22238 2991 22272
rect 3025 22238 3129 22272
rect 3163 22238 3267 22272
rect 3301 22238 3405 22272
rect 3439 22238 3543 22272
rect 3577 22238 3681 22272
rect 3715 22238 3819 22272
rect 3853 22238 3957 22272
rect 3991 22238 4095 22272
rect 4129 22238 4233 22272
rect 4267 22238 4371 22272
rect 4405 22238 4509 22272
rect 4543 22238 4647 22272
rect 4681 22238 4692 22272
rect 2704 22135 4692 22238
rect 2704 22101 2715 22135
rect 2749 22101 2853 22135
rect 2887 22101 2991 22135
rect 3025 22101 3129 22135
rect 3163 22101 3267 22135
rect 3301 22101 3405 22135
rect 3439 22101 3543 22135
rect 3577 22101 3681 22135
rect 3715 22101 3819 22135
rect 3853 22101 3957 22135
rect 3991 22101 4095 22135
rect 4129 22101 4233 22135
rect 4267 22101 4371 22135
rect 4405 22101 4509 22135
rect 4543 22101 4647 22135
rect 4681 22101 4692 22135
rect 2704 21998 4692 22101
rect 2704 21964 2715 21998
rect 2749 21964 2853 21998
rect 2887 21964 2991 21998
rect 3025 21964 3129 21998
rect 3163 21964 3267 21998
rect 3301 21964 3405 21998
rect 3439 21964 3543 21998
rect 3577 21964 3681 21998
rect 3715 21964 3819 21998
rect 3853 21964 3957 21998
rect 3991 21964 4095 21998
rect 4129 21964 4233 21998
rect 4267 21964 4371 21998
rect 4405 21964 4509 21998
rect 4543 21964 4647 21998
rect 4681 21964 4692 21998
rect 2704 21861 4692 21964
rect 2704 21827 2715 21861
rect 2749 21827 2853 21861
rect 2887 21827 2991 21861
rect 3025 21827 3129 21861
rect 3163 21827 3267 21861
rect 3301 21827 3405 21861
rect 3439 21827 3543 21861
rect 3577 21827 3681 21861
rect 3715 21827 3819 21861
rect 3853 21827 3957 21861
rect 3991 21827 4095 21861
rect 4129 21827 4233 21861
rect 4267 21827 4371 21861
rect 4405 21827 4509 21861
rect 4543 21827 4647 21861
rect 4681 21827 4692 21861
rect 2704 21724 4692 21827
rect 2704 21690 2715 21724
rect 2749 21690 2853 21724
rect 2887 21690 2991 21724
rect 3025 21690 3129 21724
rect 3163 21690 3267 21724
rect 3301 21690 3405 21724
rect 3439 21690 3543 21724
rect 3577 21690 3681 21724
rect 3715 21690 3819 21724
rect 3853 21690 3957 21724
rect 3991 21690 4095 21724
rect 4129 21690 4233 21724
rect 4267 21690 4371 21724
rect 4405 21690 4509 21724
rect 4543 21690 4647 21724
rect 4681 21690 4692 21724
rect 2704 21587 4692 21690
rect 2704 21553 2715 21587
rect 2749 21553 2853 21587
rect 2887 21553 2991 21587
rect 3025 21553 3129 21587
rect 3163 21553 3267 21587
rect 3301 21553 3405 21587
rect 3439 21553 3543 21587
rect 3577 21553 3681 21587
rect 3715 21553 3819 21587
rect 3853 21553 3957 21587
rect 3991 21553 4095 21587
rect 4129 21553 4233 21587
rect 4267 21553 4371 21587
rect 4405 21553 4509 21587
rect 4543 21553 4647 21587
rect 4681 21553 4692 21587
rect 2704 21450 4692 21553
rect 2704 21416 2715 21450
rect 2749 21416 2853 21450
rect 2887 21416 2991 21450
rect 3025 21416 3129 21450
rect 3163 21416 3267 21450
rect 3301 21416 3405 21450
rect 3439 21416 3543 21450
rect 3577 21416 3681 21450
rect 3715 21416 3819 21450
rect 3853 21416 3957 21450
rect 3991 21416 4095 21450
rect 4129 21416 4233 21450
rect 4267 21416 4371 21450
rect 4405 21416 4509 21450
rect 4543 21416 4647 21450
rect 4681 21416 4692 21450
rect 2704 21313 4692 21416
rect 2704 21279 2715 21313
rect 2749 21279 2853 21313
rect 2887 21279 2991 21313
rect 3025 21279 3129 21313
rect 3163 21279 3267 21313
rect 3301 21279 3405 21313
rect 3439 21279 3543 21313
rect 3577 21279 3681 21313
rect 3715 21279 3819 21313
rect 3853 21279 3957 21313
rect 3991 21279 4095 21313
rect 4129 21279 4233 21313
rect 4267 21279 4371 21313
rect 4405 21279 4509 21313
rect 4543 21279 4647 21313
rect 4681 21279 4692 21313
rect 2704 21176 4692 21279
rect 2704 21142 2715 21176
rect 2749 21142 2853 21176
rect 2887 21142 2991 21176
rect 3025 21142 3129 21176
rect 3163 21142 3267 21176
rect 3301 21142 3405 21176
rect 3439 21142 3543 21176
rect 3577 21142 3681 21176
rect 3715 21142 3819 21176
rect 3853 21142 3957 21176
rect 3991 21142 4095 21176
rect 4129 21142 4233 21176
rect 4267 21142 4371 21176
rect 4405 21142 4509 21176
rect 4543 21142 4647 21176
rect 4681 21142 4692 21176
rect 2704 21039 4692 21142
rect 2704 21005 2715 21039
rect 2749 21005 2853 21039
rect 2887 21005 2991 21039
rect 3025 21005 3129 21039
rect 3163 21005 3267 21039
rect 3301 21005 3405 21039
rect 3439 21005 3543 21039
rect 3577 21005 3681 21039
rect 3715 21005 3819 21039
rect 3853 21005 3957 21039
rect 3991 21005 4095 21039
rect 4129 21005 4233 21039
rect 4267 21005 4371 21039
rect 4405 21005 4509 21039
rect 4543 21005 4647 21039
rect 4681 21005 4692 21039
rect 2704 20902 4692 21005
rect 2704 20868 2715 20902
rect 2749 20868 2853 20902
rect 2887 20868 2991 20902
rect 3025 20868 3129 20902
rect 3163 20868 3267 20902
rect 3301 20868 3405 20902
rect 3439 20868 3543 20902
rect 3577 20868 3681 20902
rect 3715 20868 3819 20902
rect 3853 20868 3957 20902
rect 3991 20868 4095 20902
rect 4129 20868 4233 20902
rect 4267 20868 4371 20902
rect 4405 20868 4509 20902
rect 4543 20868 4647 20902
rect 4681 20868 4692 20902
rect 2704 20765 4692 20868
rect 2704 20731 2715 20765
rect 2749 20731 2853 20765
rect 2887 20731 2991 20765
rect 3025 20731 3129 20765
rect 3163 20731 3267 20765
rect 3301 20731 3405 20765
rect 3439 20731 3543 20765
rect 3577 20731 3681 20765
rect 3715 20731 3819 20765
rect 3853 20731 3957 20765
rect 3991 20731 4095 20765
rect 4129 20731 4233 20765
rect 4267 20731 4371 20765
rect 4405 20731 4509 20765
rect 4543 20731 4647 20765
rect 4681 20731 4692 20765
rect 2704 20628 4692 20731
rect 2704 20594 2715 20628
rect 2749 20594 2853 20628
rect 2887 20594 2991 20628
rect 3025 20594 3129 20628
rect 3163 20594 3267 20628
rect 3301 20594 3405 20628
rect 3439 20594 3543 20628
rect 3577 20594 3681 20628
rect 3715 20594 3819 20628
rect 3853 20594 3957 20628
rect 3991 20594 4095 20628
rect 4129 20594 4233 20628
rect 4267 20594 4371 20628
rect 4405 20594 4509 20628
rect 4543 20594 4647 20628
rect 4681 20594 4692 20628
rect 2704 20491 4692 20594
rect 2704 20457 2715 20491
rect 2749 20457 2853 20491
rect 2887 20457 2991 20491
rect 3025 20457 3129 20491
rect 3163 20457 3267 20491
rect 3301 20457 3405 20491
rect 3439 20457 3543 20491
rect 3577 20457 3681 20491
rect 3715 20457 3819 20491
rect 3853 20457 3957 20491
rect 3991 20457 4095 20491
rect 4129 20457 4233 20491
rect 4267 20457 4371 20491
rect 4405 20457 4509 20491
rect 4543 20457 4647 20491
rect 4681 20457 4692 20491
rect 2704 20354 4692 20457
rect 2704 20320 2715 20354
rect 2749 20320 2853 20354
rect 2887 20320 2991 20354
rect 3025 20320 3129 20354
rect 3163 20320 3267 20354
rect 3301 20320 3405 20354
rect 3439 20320 3543 20354
rect 3577 20320 3681 20354
rect 3715 20320 3819 20354
rect 3853 20320 3957 20354
rect 3991 20320 4095 20354
rect 4129 20320 4233 20354
rect 4267 20320 4371 20354
rect 4405 20320 4509 20354
rect 4543 20320 4647 20354
rect 4681 20320 4692 20354
rect 2704 20217 4692 20320
rect 2704 20183 2715 20217
rect 2749 20183 2853 20217
rect 2887 20183 2991 20217
rect 3025 20183 3129 20217
rect 3163 20183 3267 20217
rect 3301 20183 3405 20217
rect 3439 20183 3543 20217
rect 3577 20183 3681 20217
rect 3715 20183 3819 20217
rect 3853 20183 3957 20217
rect 3991 20183 4095 20217
rect 4129 20183 4233 20217
rect 4267 20183 4371 20217
rect 4405 20183 4509 20217
rect 4543 20183 4647 20217
rect 4681 20183 4692 20217
rect 2704 20080 4692 20183
rect 2704 20046 2715 20080
rect 2749 20046 2853 20080
rect 2887 20046 2991 20080
rect 3025 20046 3129 20080
rect 3163 20046 3267 20080
rect 3301 20046 3405 20080
rect 3439 20046 3543 20080
rect 3577 20046 3681 20080
rect 3715 20046 3819 20080
rect 3853 20046 3957 20080
rect 3991 20046 4095 20080
rect 4129 20046 4233 20080
rect 4267 20046 4371 20080
rect 4405 20046 4509 20080
rect 4543 20046 4647 20080
rect 4681 20046 4692 20080
rect 2704 19943 4692 20046
rect 2704 19909 2715 19943
rect 2749 19909 2853 19943
rect 2887 19909 2991 19943
rect 3025 19909 3129 19943
rect 3163 19909 3267 19943
rect 3301 19909 3405 19943
rect 3439 19909 3543 19943
rect 3577 19909 3681 19943
rect 3715 19909 3819 19943
rect 3853 19909 3957 19943
rect 3991 19909 4095 19943
rect 4129 19909 4233 19943
rect 4267 19909 4371 19943
rect 4405 19909 4509 19943
rect 4543 19909 4647 19943
rect 4681 19909 4692 19943
rect 2704 19806 4692 19909
rect 2704 19772 2715 19806
rect 2749 19772 2853 19806
rect 2887 19772 2991 19806
rect 3025 19772 3129 19806
rect 3163 19772 3267 19806
rect 3301 19772 3405 19806
rect 3439 19772 3543 19806
rect 3577 19772 3681 19806
rect 3715 19772 3819 19806
rect 3853 19772 3957 19806
rect 3991 19772 4095 19806
rect 4129 19772 4233 19806
rect 4267 19772 4371 19806
rect 4405 19772 4509 19806
rect 4543 19772 4647 19806
rect 4681 19772 4692 19806
rect 2704 19669 4692 19772
rect 2704 19635 2715 19669
rect 2749 19635 2853 19669
rect 2887 19635 2991 19669
rect 3025 19635 3129 19669
rect 3163 19635 3267 19669
rect 3301 19635 3405 19669
rect 3439 19635 3543 19669
rect 3577 19635 3681 19669
rect 3715 19635 3819 19669
rect 3853 19635 3957 19669
rect 3991 19635 4095 19669
rect 4129 19635 4233 19669
rect 4267 19635 4371 19669
rect 4405 19635 4509 19669
rect 4543 19635 4647 19669
rect 4681 19635 4692 19669
rect 2704 19532 4692 19635
rect 2704 19498 2715 19532
rect 2749 19498 2853 19532
rect 2887 19498 2991 19532
rect 3025 19498 3129 19532
rect 3163 19498 3267 19532
rect 3301 19498 3405 19532
rect 3439 19498 3543 19532
rect 3577 19498 3681 19532
rect 3715 19498 3819 19532
rect 3853 19498 3957 19532
rect 3991 19498 4095 19532
rect 4129 19498 4233 19532
rect 4267 19498 4371 19532
rect 4405 19498 4509 19532
rect 4543 19498 4647 19532
rect 4681 19498 4692 19532
rect 2704 19395 4692 19498
rect 2704 19361 2715 19395
rect 2749 19361 2853 19395
rect 2887 19361 2991 19395
rect 3025 19361 3129 19395
rect 3163 19361 3267 19395
rect 3301 19361 3405 19395
rect 3439 19361 3543 19395
rect 3577 19361 3681 19395
rect 3715 19361 3819 19395
rect 3853 19361 3957 19395
rect 3991 19361 4095 19395
rect 4129 19361 4233 19395
rect 4267 19361 4371 19395
rect 4405 19361 4509 19395
rect 4543 19361 4647 19395
rect 4681 19361 4692 19395
rect 2704 19258 4692 19361
rect 2704 19224 2715 19258
rect 2749 19224 2853 19258
rect 2887 19224 2991 19258
rect 3025 19224 3129 19258
rect 3163 19224 3267 19258
rect 3301 19224 3405 19258
rect 3439 19224 3543 19258
rect 3577 19224 3681 19258
rect 3715 19224 3819 19258
rect 3853 19224 3957 19258
rect 3991 19224 4095 19258
rect 4129 19224 4233 19258
rect 4267 19224 4371 19258
rect 4405 19224 4509 19258
rect 4543 19224 4647 19258
rect 4681 19224 4692 19258
rect 2704 19121 4692 19224
rect 2704 19087 2715 19121
rect 2749 19087 2853 19121
rect 2887 19087 2991 19121
rect 3025 19087 3129 19121
rect 3163 19087 3267 19121
rect 3301 19087 3405 19121
rect 3439 19087 3543 19121
rect 3577 19087 3681 19121
rect 3715 19087 3819 19121
rect 3853 19087 3957 19121
rect 3991 19087 4095 19121
rect 4129 19087 4233 19121
rect 4267 19087 4371 19121
rect 4405 19087 4509 19121
rect 4543 19087 4647 19121
rect 4681 19087 4692 19121
rect 2704 18984 4692 19087
rect 2704 18950 2715 18984
rect 2749 18950 2853 18984
rect 2887 18950 2991 18984
rect 3025 18950 3129 18984
rect 3163 18950 3267 18984
rect 3301 18950 3405 18984
rect 3439 18950 3543 18984
rect 3577 18950 3681 18984
rect 3715 18950 3819 18984
rect 3853 18950 3957 18984
rect 3991 18950 4095 18984
rect 4129 18950 4233 18984
rect 4267 18950 4371 18984
rect 4405 18950 4509 18984
rect 4543 18950 4647 18984
rect 4681 18950 4692 18984
rect 2704 18847 4692 18950
rect 2704 18813 2715 18847
rect 2749 18813 2853 18847
rect 2887 18813 2991 18847
rect 3025 18813 3129 18847
rect 3163 18813 3267 18847
rect 3301 18813 3405 18847
rect 3439 18813 3543 18847
rect 3577 18813 3681 18847
rect 3715 18813 3819 18847
rect 3853 18813 3957 18847
rect 3991 18813 4095 18847
rect 4129 18813 4233 18847
rect 4267 18813 4371 18847
rect 4405 18813 4509 18847
rect 4543 18813 4647 18847
rect 4681 18813 4692 18847
rect 2704 18710 4692 18813
rect 2704 18676 2715 18710
rect 2749 18676 2853 18710
rect 2887 18676 2991 18710
rect 3025 18676 3129 18710
rect 3163 18676 3267 18710
rect 3301 18676 3405 18710
rect 3439 18676 3543 18710
rect 3577 18676 3681 18710
rect 3715 18676 3819 18710
rect 3853 18676 3957 18710
rect 3991 18676 4095 18710
rect 4129 18676 4233 18710
rect 4267 18676 4371 18710
rect 4405 18676 4509 18710
rect 4543 18676 4647 18710
rect 4681 18676 4692 18710
rect 2704 18573 4692 18676
rect 2704 18539 2715 18573
rect 2749 18539 2853 18573
rect 2887 18539 2991 18573
rect 3025 18539 3129 18573
rect 3163 18539 3267 18573
rect 3301 18539 3405 18573
rect 3439 18539 3543 18573
rect 3577 18539 3681 18573
rect 3715 18539 3819 18573
rect 3853 18539 3957 18573
rect 3991 18539 4095 18573
rect 4129 18539 4233 18573
rect 4267 18539 4371 18573
rect 4405 18539 4509 18573
rect 4543 18539 4647 18573
rect 4681 18539 4692 18573
rect 2704 18436 4692 18539
rect 2704 18402 2715 18436
rect 2749 18402 2853 18436
rect 2887 18402 2991 18436
rect 3025 18402 3129 18436
rect 3163 18402 3267 18436
rect 3301 18402 3405 18436
rect 3439 18402 3543 18436
rect 3577 18402 3681 18436
rect 3715 18402 3819 18436
rect 3853 18402 3957 18436
rect 3991 18402 4095 18436
rect 4129 18402 4233 18436
rect 4267 18402 4371 18436
rect 4405 18402 4509 18436
rect 4543 18402 4647 18436
rect 4681 18402 4692 18436
rect 2704 18299 4692 18402
rect 2704 18265 2715 18299
rect 2749 18265 2853 18299
rect 2887 18265 2991 18299
rect 3025 18265 3129 18299
rect 3163 18265 3267 18299
rect 3301 18265 3405 18299
rect 3439 18265 3543 18299
rect 3577 18265 3681 18299
rect 3715 18265 3819 18299
rect 3853 18265 3957 18299
rect 3991 18265 4095 18299
rect 4129 18265 4233 18299
rect 4267 18265 4371 18299
rect 4405 18265 4509 18299
rect 4543 18265 4647 18299
rect 4681 18265 4692 18299
rect 2704 18162 4692 18265
rect 2704 18128 2715 18162
rect 2749 18128 2853 18162
rect 2887 18128 2991 18162
rect 3025 18128 3129 18162
rect 3163 18128 3267 18162
rect 3301 18128 3405 18162
rect 3439 18128 3543 18162
rect 3577 18128 3681 18162
rect 3715 18128 3819 18162
rect 3853 18128 3957 18162
rect 3991 18128 4095 18162
rect 4129 18128 4233 18162
rect 4267 18128 4371 18162
rect 4405 18128 4509 18162
rect 4543 18128 4647 18162
rect 4681 18128 4692 18162
rect 2704 18025 4692 18128
rect 2704 17991 2715 18025
rect 2749 17991 2853 18025
rect 2887 17991 2991 18025
rect 3025 17991 3129 18025
rect 3163 17991 3267 18025
rect 3301 17991 3405 18025
rect 3439 17991 3543 18025
rect 3577 17991 3681 18025
rect 3715 17991 3819 18025
rect 3853 17991 3957 18025
rect 3991 17991 4095 18025
rect 4129 17991 4233 18025
rect 4267 17991 4371 18025
rect 4405 17991 4509 18025
rect 4543 17991 4647 18025
rect 4681 17991 4692 18025
rect 2704 17888 4692 17991
rect 2704 17854 2715 17888
rect 2749 17854 2853 17888
rect 2887 17854 2991 17888
rect 3025 17854 3129 17888
rect 3163 17854 3267 17888
rect 3301 17854 3405 17888
rect 3439 17854 3543 17888
rect 3577 17854 3681 17888
rect 3715 17854 3819 17888
rect 3853 17854 3957 17888
rect 3991 17854 4095 17888
rect 4129 17854 4233 17888
rect 4267 17854 4371 17888
rect 4405 17854 4509 17888
rect 4543 17854 4647 17888
rect 4681 17854 4692 17888
rect 2704 17751 4692 17854
rect 2704 17717 2715 17751
rect 2749 17717 2853 17751
rect 2887 17717 2991 17751
rect 3025 17717 3129 17751
rect 3163 17717 3267 17751
rect 3301 17717 3405 17751
rect 3439 17717 3543 17751
rect 3577 17717 3681 17751
rect 3715 17717 3819 17751
rect 3853 17717 3957 17751
rect 3991 17717 4095 17751
rect 4129 17717 4233 17751
rect 4267 17717 4371 17751
rect 4405 17717 4509 17751
rect 4543 17717 4647 17751
rect 4681 17717 4692 17751
rect 2704 17614 4692 17717
rect 2704 17580 2715 17614
rect 2749 17580 2853 17614
rect 2887 17580 2991 17614
rect 3025 17580 3129 17614
rect 3163 17580 3267 17614
rect 3301 17580 3405 17614
rect 3439 17580 3543 17614
rect 3577 17580 3681 17614
rect 3715 17580 3819 17614
rect 3853 17580 3957 17614
rect 3991 17580 4095 17614
rect 4129 17580 4233 17614
rect 4267 17580 4371 17614
rect 4405 17580 4509 17614
rect 4543 17580 4647 17614
rect 4681 17580 4692 17614
rect 2704 17477 4692 17580
rect 2704 17443 2715 17477
rect 2749 17443 2853 17477
rect 2887 17443 2991 17477
rect 3025 17443 3129 17477
rect 3163 17443 3267 17477
rect 3301 17443 3405 17477
rect 3439 17443 3543 17477
rect 3577 17443 3681 17477
rect 3715 17443 3819 17477
rect 3853 17443 3957 17477
rect 3991 17443 4095 17477
rect 4129 17443 4233 17477
rect 4267 17443 4371 17477
rect 4405 17443 4509 17477
rect 4543 17443 4647 17477
rect 4681 17443 4692 17477
rect 2704 17340 4692 17443
rect 2704 17306 2715 17340
rect 2749 17306 2853 17340
rect 2887 17306 2991 17340
rect 3025 17306 3129 17340
rect 3163 17306 3267 17340
rect 3301 17306 3405 17340
rect 3439 17306 3543 17340
rect 3577 17306 3681 17340
rect 3715 17306 3819 17340
rect 3853 17306 3957 17340
rect 3991 17306 4095 17340
rect 4129 17306 4233 17340
rect 4267 17306 4371 17340
rect 4405 17306 4509 17340
rect 4543 17306 4647 17340
rect 4681 17306 4692 17340
rect 2704 17203 4692 17306
rect 2704 17169 2715 17203
rect 2749 17169 2853 17203
rect 2887 17169 2991 17203
rect 3025 17169 3129 17203
rect 3163 17169 3267 17203
rect 3301 17169 3405 17203
rect 3439 17169 3543 17203
rect 3577 17169 3681 17203
rect 3715 17169 3819 17203
rect 3853 17169 3957 17203
rect 3991 17169 4095 17203
rect 4129 17169 4233 17203
rect 4267 17169 4371 17203
rect 4405 17169 4509 17203
rect 4543 17169 4647 17203
rect 4681 17169 4692 17203
rect 2704 17072 4692 17169
rect 2704 17066 7908 17072
rect 2704 17032 2715 17066
rect 2749 17032 2853 17066
rect 2887 17032 2991 17066
rect 3025 17032 3129 17066
rect 3163 17032 3267 17066
rect 3301 17032 3405 17066
rect 3439 17032 3543 17066
rect 3577 17032 3681 17066
rect 3715 17032 3819 17066
rect 3853 17032 3957 17066
rect 3991 17032 4095 17066
rect 4129 17032 4233 17066
rect 4267 17032 4371 17066
rect 4405 17032 4509 17066
rect 4543 17032 4647 17066
rect 4681 17034 7908 17066
rect 4681 17032 4740 17034
rect 2704 17000 4740 17032
rect 4774 17000 4809 17034
rect 4843 17000 4878 17034
rect 4912 17000 4947 17034
rect 4981 17000 5016 17034
rect 5050 17000 5085 17034
rect 5119 17000 5154 17034
rect 5188 17000 5223 17034
rect 5257 17000 5292 17034
rect 5326 17000 5361 17034
rect 5395 17000 5430 17034
rect 5464 17000 5499 17034
rect 5533 17000 5568 17034
rect 5602 17000 5637 17034
rect 5671 17000 5706 17034
rect 5740 17000 5775 17034
rect 5809 17000 5844 17034
rect 5878 17000 5913 17034
rect 5947 17000 5982 17034
rect 6016 17000 6051 17034
rect 6085 17000 6120 17034
rect 6154 17000 6189 17034
rect 6223 17000 6258 17034
rect 6292 17000 6327 17034
rect 6361 17000 6396 17034
rect 6430 17000 6465 17034
rect 6499 17000 6534 17034
rect 6568 17000 6603 17034
rect 6637 17000 6672 17034
rect 6706 17000 6741 17034
rect 6775 17000 6810 17034
rect 6844 17000 6879 17034
rect 6913 17000 6948 17034
rect 6982 17000 7017 17034
rect 7051 17000 7086 17034
rect 7120 17000 7155 17034
rect 7189 17000 7224 17034
rect 7258 17000 7293 17034
rect 7327 17000 7362 17034
rect 7396 17000 7431 17034
rect 7465 17000 7500 17034
rect 7534 17000 7568 17034
rect 7602 17000 7636 17034
rect 7670 17000 7704 17034
rect 7738 17000 7772 17034
rect 7806 17000 7840 17034
rect 7874 17000 7908 17034
rect 2704 16964 7908 17000
rect 2704 16930 4740 16964
rect 4774 16930 4809 16964
rect 4843 16930 4878 16964
rect 4912 16930 4947 16964
rect 4981 16930 5016 16964
rect 5050 16930 5085 16964
rect 5119 16930 5154 16964
rect 5188 16930 5223 16964
rect 5257 16930 5292 16964
rect 5326 16930 5361 16964
rect 5395 16930 5430 16964
rect 5464 16930 5499 16964
rect 5533 16930 5568 16964
rect 5602 16930 5637 16964
rect 5671 16930 5706 16964
rect 5740 16930 5775 16964
rect 5809 16930 5844 16964
rect 5878 16930 5913 16964
rect 5947 16930 5982 16964
rect 6016 16930 6051 16964
rect 6085 16930 6120 16964
rect 6154 16930 6189 16964
rect 6223 16930 6258 16964
rect 6292 16930 6327 16964
rect 6361 16930 6396 16964
rect 6430 16930 6465 16964
rect 6499 16930 6534 16964
rect 6568 16930 6603 16964
rect 6637 16930 6672 16964
rect 6706 16930 6741 16964
rect 6775 16930 6810 16964
rect 6844 16930 6879 16964
rect 6913 16930 6948 16964
rect 6982 16930 7017 16964
rect 7051 16930 7086 16964
rect 7120 16930 7155 16964
rect 7189 16930 7224 16964
rect 7258 16930 7293 16964
rect 7327 16930 7362 16964
rect 7396 16930 7431 16964
rect 7465 16930 7500 16964
rect 7534 16930 7568 16964
rect 7602 16930 7636 16964
rect 7670 16930 7704 16964
rect 7738 16930 7772 16964
rect 7806 16930 7840 16964
rect 7874 16930 7908 16964
rect 2704 16929 7908 16930
rect 2704 16895 2715 16929
rect 2749 16895 2853 16929
rect 2887 16895 2991 16929
rect 3025 16895 3129 16929
rect 3163 16895 3267 16929
rect 3301 16895 3405 16929
rect 3439 16895 3543 16929
rect 3577 16895 3681 16929
rect 3715 16895 3819 16929
rect 3853 16895 3957 16929
rect 3991 16895 4095 16929
rect 4129 16895 4233 16929
rect 4267 16895 4371 16929
rect 4405 16895 4509 16929
rect 4543 16895 4647 16929
rect 4681 16895 7908 16929
rect 2704 16894 7908 16895
rect 2704 16860 4740 16894
rect 4774 16860 4809 16894
rect 4843 16860 4878 16894
rect 4912 16860 4947 16894
rect 4981 16860 5016 16894
rect 5050 16860 5085 16894
rect 5119 16860 5154 16894
rect 5188 16860 5223 16894
rect 5257 16860 5292 16894
rect 5326 16860 5361 16894
rect 5395 16860 5430 16894
rect 5464 16860 5499 16894
rect 5533 16860 5568 16894
rect 5602 16860 5637 16894
rect 5671 16860 5706 16894
rect 5740 16860 5775 16894
rect 5809 16860 5844 16894
rect 5878 16860 5913 16894
rect 5947 16860 5982 16894
rect 6016 16860 6051 16894
rect 6085 16860 6120 16894
rect 6154 16860 6189 16894
rect 6223 16860 6258 16894
rect 6292 16860 6327 16894
rect 6361 16860 6396 16894
rect 6430 16860 6465 16894
rect 6499 16860 6534 16894
rect 6568 16860 6603 16894
rect 6637 16860 6672 16894
rect 6706 16860 6741 16894
rect 6775 16860 6810 16894
rect 6844 16860 6879 16894
rect 6913 16860 6948 16894
rect 6982 16860 7017 16894
rect 7051 16860 7086 16894
rect 7120 16860 7155 16894
rect 7189 16860 7224 16894
rect 7258 16860 7293 16894
rect 7327 16860 7362 16894
rect 7396 16860 7431 16894
rect 7465 16860 7500 16894
rect 7534 16860 7568 16894
rect 7602 16860 7636 16894
rect 7670 16860 7704 16894
rect 7738 16860 7772 16894
rect 7806 16860 7840 16894
rect 7874 16860 7908 16894
rect 2704 16824 7908 16860
rect 2704 16792 4740 16824
rect 2704 16758 2715 16792
rect 2749 16758 2853 16792
rect 2887 16758 2991 16792
rect 3025 16758 3129 16792
rect 3163 16758 3267 16792
rect 3301 16758 3405 16792
rect 3439 16758 3543 16792
rect 3577 16758 3681 16792
rect 3715 16758 3819 16792
rect 3853 16758 3957 16792
rect 3991 16758 4095 16792
rect 4129 16758 4233 16792
rect 4267 16758 4371 16792
rect 4405 16758 4509 16792
rect 4543 16758 4647 16792
rect 4681 16790 4740 16792
rect 4774 16790 4809 16824
rect 4843 16790 4878 16824
rect 4912 16790 4947 16824
rect 4981 16790 5016 16824
rect 5050 16790 5085 16824
rect 5119 16790 5154 16824
rect 5188 16790 5223 16824
rect 5257 16790 5292 16824
rect 5326 16790 5361 16824
rect 5395 16790 5430 16824
rect 5464 16790 5499 16824
rect 5533 16790 5568 16824
rect 5602 16790 5637 16824
rect 5671 16790 5706 16824
rect 5740 16790 5775 16824
rect 5809 16790 5844 16824
rect 5878 16790 5913 16824
rect 5947 16790 5982 16824
rect 6016 16790 6051 16824
rect 6085 16790 6120 16824
rect 6154 16790 6189 16824
rect 6223 16790 6258 16824
rect 6292 16790 6327 16824
rect 6361 16790 6396 16824
rect 6430 16790 6465 16824
rect 6499 16790 6534 16824
rect 6568 16790 6603 16824
rect 6637 16790 6672 16824
rect 6706 16790 6741 16824
rect 6775 16790 6810 16824
rect 6844 16790 6879 16824
rect 6913 16790 6948 16824
rect 6982 16790 7017 16824
rect 7051 16790 7086 16824
rect 7120 16790 7155 16824
rect 7189 16790 7224 16824
rect 7258 16790 7293 16824
rect 7327 16790 7362 16824
rect 7396 16790 7431 16824
rect 7465 16790 7500 16824
rect 7534 16790 7568 16824
rect 7602 16790 7636 16824
rect 7670 16790 7704 16824
rect 7738 16790 7772 16824
rect 7806 16790 7840 16824
rect 7874 16790 7908 16824
rect 4681 16758 7908 16790
rect 2704 16754 7908 16758
rect 2704 16720 4740 16754
rect 4774 16720 4809 16754
rect 4843 16720 4878 16754
rect 4912 16720 4947 16754
rect 4981 16720 5016 16754
rect 5050 16720 5085 16754
rect 5119 16720 5154 16754
rect 5188 16720 5223 16754
rect 5257 16720 5292 16754
rect 5326 16720 5361 16754
rect 5395 16720 5430 16754
rect 5464 16720 5499 16754
rect 5533 16720 5568 16754
rect 5602 16720 5637 16754
rect 5671 16720 5706 16754
rect 5740 16720 5775 16754
rect 5809 16720 5844 16754
rect 5878 16720 5913 16754
rect 5947 16720 5982 16754
rect 6016 16720 6051 16754
rect 6085 16720 6120 16754
rect 6154 16720 6189 16754
rect 6223 16720 6258 16754
rect 6292 16720 6327 16754
rect 6361 16720 6396 16754
rect 6430 16720 6465 16754
rect 6499 16720 6534 16754
rect 6568 16720 6603 16754
rect 6637 16720 6672 16754
rect 6706 16720 6741 16754
rect 6775 16720 6810 16754
rect 6844 16720 6879 16754
rect 6913 16720 6948 16754
rect 6982 16720 7017 16754
rect 7051 16720 7086 16754
rect 7120 16720 7155 16754
rect 7189 16720 7224 16754
rect 7258 16720 7293 16754
rect 7327 16720 7362 16754
rect 7396 16720 7431 16754
rect 7465 16720 7500 16754
rect 7534 16720 7568 16754
rect 7602 16720 7636 16754
rect 7670 16720 7704 16754
rect 7738 16720 7772 16754
rect 7806 16720 7840 16754
rect 7874 16720 7908 16754
rect 2704 16684 7908 16720
rect 2704 16655 4740 16684
rect 2704 16621 2715 16655
rect 2749 16621 2853 16655
rect 2887 16621 2991 16655
rect 3025 16621 3129 16655
rect 3163 16621 3267 16655
rect 3301 16621 3405 16655
rect 3439 16621 3543 16655
rect 3577 16621 3681 16655
rect 3715 16621 3819 16655
rect 3853 16621 3957 16655
rect 3991 16621 4095 16655
rect 4129 16621 4233 16655
rect 4267 16621 4371 16655
rect 4405 16621 4509 16655
rect 4543 16621 4647 16655
rect 4681 16650 4740 16655
rect 4774 16650 4809 16684
rect 4843 16650 4878 16684
rect 4912 16650 4947 16684
rect 4981 16650 5016 16684
rect 5050 16650 5085 16684
rect 5119 16650 5154 16684
rect 5188 16650 5223 16684
rect 5257 16650 5292 16684
rect 5326 16650 5361 16684
rect 5395 16650 5430 16684
rect 5464 16650 5499 16684
rect 5533 16650 5568 16684
rect 5602 16650 5637 16684
rect 5671 16650 5706 16684
rect 5740 16650 5775 16684
rect 5809 16650 5844 16684
rect 5878 16650 5913 16684
rect 5947 16650 5982 16684
rect 6016 16650 6051 16684
rect 6085 16650 6120 16684
rect 6154 16650 6189 16684
rect 6223 16650 6258 16684
rect 6292 16650 6327 16684
rect 6361 16650 6396 16684
rect 6430 16650 6465 16684
rect 6499 16650 6534 16684
rect 6568 16650 6603 16684
rect 6637 16650 6672 16684
rect 6706 16650 6741 16684
rect 6775 16650 6810 16684
rect 6844 16650 6879 16684
rect 6913 16650 6948 16684
rect 6982 16650 7017 16684
rect 7051 16650 7086 16684
rect 7120 16650 7155 16684
rect 7189 16650 7224 16684
rect 7258 16650 7293 16684
rect 7327 16650 7362 16684
rect 7396 16650 7431 16684
rect 7465 16650 7500 16684
rect 7534 16650 7568 16684
rect 7602 16650 7636 16684
rect 7670 16650 7704 16684
rect 7738 16650 7772 16684
rect 7806 16650 7840 16684
rect 7874 16650 7908 16684
rect 4681 16621 7908 16650
rect 2704 16614 7908 16621
rect 2704 16580 4740 16614
rect 4774 16580 4809 16614
rect 4843 16580 4878 16614
rect 4912 16580 4947 16614
rect 4981 16580 5016 16614
rect 5050 16580 5085 16614
rect 5119 16580 5154 16614
rect 5188 16580 5223 16614
rect 5257 16580 5292 16614
rect 5326 16580 5361 16614
rect 5395 16580 5430 16614
rect 5464 16580 5499 16614
rect 5533 16580 5568 16614
rect 5602 16580 5637 16614
rect 5671 16580 5706 16614
rect 5740 16580 5775 16614
rect 5809 16580 5844 16614
rect 5878 16580 5913 16614
rect 5947 16580 5982 16614
rect 6016 16580 6051 16614
rect 6085 16580 6120 16614
rect 6154 16580 6189 16614
rect 6223 16580 6258 16614
rect 6292 16580 6327 16614
rect 6361 16580 6396 16614
rect 6430 16580 6465 16614
rect 6499 16580 6534 16614
rect 6568 16580 6603 16614
rect 6637 16580 6672 16614
rect 6706 16580 6741 16614
rect 6775 16580 6810 16614
rect 6844 16580 6879 16614
rect 6913 16580 6948 16614
rect 6982 16580 7017 16614
rect 7051 16580 7086 16614
rect 7120 16580 7155 16614
rect 7189 16580 7224 16614
rect 7258 16580 7293 16614
rect 7327 16580 7362 16614
rect 7396 16580 7431 16614
rect 7465 16580 7500 16614
rect 7534 16580 7568 16614
rect 7602 16580 7636 16614
rect 7670 16580 7704 16614
rect 7738 16580 7772 16614
rect 7806 16580 7840 16614
rect 7874 16580 7908 16614
rect 2704 16544 7908 16580
rect 2704 16518 4740 16544
rect 2704 16484 2715 16518
rect 2749 16484 2853 16518
rect 2887 16484 2991 16518
rect 3025 16484 3129 16518
rect 3163 16484 3267 16518
rect 3301 16484 3405 16518
rect 3439 16484 3543 16518
rect 3577 16484 3681 16518
rect 3715 16484 3819 16518
rect 3853 16484 3957 16518
rect 3991 16484 4095 16518
rect 4129 16484 4233 16518
rect 4267 16484 4371 16518
rect 4405 16484 4509 16518
rect 4543 16484 4647 16518
rect 4681 16510 4740 16518
rect 4774 16510 4809 16544
rect 4843 16510 4878 16544
rect 4912 16510 4947 16544
rect 4981 16510 5016 16544
rect 5050 16510 5085 16544
rect 5119 16510 5154 16544
rect 5188 16510 5223 16544
rect 5257 16510 5292 16544
rect 5326 16510 5361 16544
rect 5395 16510 5430 16544
rect 5464 16510 5499 16544
rect 5533 16510 5568 16544
rect 5602 16510 5637 16544
rect 5671 16510 5706 16544
rect 5740 16510 5775 16544
rect 5809 16510 5844 16544
rect 5878 16510 5913 16544
rect 5947 16510 5982 16544
rect 6016 16510 6051 16544
rect 6085 16510 6120 16544
rect 6154 16510 6189 16544
rect 6223 16510 6258 16544
rect 6292 16510 6327 16544
rect 6361 16510 6396 16544
rect 6430 16510 6465 16544
rect 6499 16510 6534 16544
rect 6568 16510 6603 16544
rect 6637 16510 6672 16544
rect 6706 16510 6741 16544
rect 6775 16510 6810 16544
rect 6844 16510 6879 16544
rect 6913 16510 6948 16544
rect 6982 16510 7017 16544
rect 7051 16510 7086 16544
rect 7120 16510 7155 16544
rect 7189 16510 7224 16544
rect 7258 16510 7293 16544
rect 7327 16510 7362 16544
rect 7396 16510 7431 16544
rect 7465 16510 7500 16544
rect 7534 16510 7568 16544
rect 7602 16510 7636 16544
rect 7670 16510 7704 16544
rect 7738 16510 7772 16544
rect 7806 16510 7840 16544
rect 7874 16510 7908 16544
rect 4681 16484 7908 16510
rect 2704 16474 7908 16484
rect 2704 16440 4740 16474
rect 4774 16440 4809 16474
rect 4843 16440 4878 16474
rect 4912 16440 4947 16474
rect 4981 16440 5016 16474
rect 5050 16440 5085 16474
rect 5119 16440 5154 16474
rect 5188 16440 5223 16474
rect 5257 16440 5292 16474
rect 5326 16440 5361 16474
rect 5395 16440 5430 16474
rect 5464 16440 5499 16474
rect 5533 16440 5568 16474
rect 5602 16440 5637 16474
rect 5671 16440 5706 16474
rect 5740 16440 5775 16474
rect 5809 16440 5844 16474
rect 5878 16440 5913 16474
rect 5947 16440 5982 16474
rect 6016 16440 6051 16474
rect 6085 16440 6120 16474
rect 6154 16440 6189 16474
rect 6223 16440 6258 16474
rect 6292 16440 6327 16474
rect 6361 16440 6396 16474
rect 6430 16440 6465 16474
rect 6499 16440 6534 16474
rect 6568 16440 6603 16474
rect 6637 16440 6672 16474
rect 6706 16440 6741 16474
rect 6775 16440 6810 16474
rect 6844 16440 6879 16474
rect 6913 16440 6948 16474
rect 6982 16440 7017 16474
rect 7051 16440 7086 16474
rect 7120 16440 7155 16474
rect 7189 16440 7224 16474
rect 7258 16440 7293 16474
rect 7327 16440 7362 16474
rect 7396 16440 7431 16474
rect 7465 16440 7500 16474
rect 7534 16440 7568 16474
rect 7602 16440 7636 16474
rect 7670 16440 7704 16474
rect 7738 16440 7772 16474
rect 7806 16440 7840 16474
rect 7874 16440 7908 16474
rect 2704 16404 7908 16440
rect 2704 16381 4740 16404
rect 2704 16347 2715 16381
rect 2749 16347 2853 16381
rect 2887 16347 2991 16381
rect 3025 16347 3129 16381
rect 3163 16347 3267 16381
rect 3301 16347 3405 16381
rect 3439 16347 3543 16381
rect 3577 16347 3681 16381
rect 3715 16347 3819 16381
rect 3853 16347 3957 16381
rect 3991 16347 4095 16381
rect 4129 16347 4233 16381
rect 4267 16347 4371 16381
rect 4405 16347 4509 16381
rect 4543 16347 4647 16381
rect 4681 16370 4740 16381
rect 4774 16370 4809 16404
rect 4843 16370 4878 16404
rect 4912 16370 4947 16404
rect 4981 16370 5016 16404
rect 5050 16370 5085 16404
rect 5119 16370 5154 16404
rect 5188 16370 5223 16404
rect 5257 16370 5292 16404
rect 5326 16370 5361 16404
rect 5395 16370 5430 16404
rect 5464 16370 5499 16404
rect 5533 16370 5568 16404
rect 5602 16370 5637 16404
rect 5671 16370 5706 16404
rect 5740 16370 5775 16404
rect 5809 16370 5844 16404
rect 5878 16370 5913 16404
rect 5947 16370 5982 16404
rect 6016 16370 6051 16404
rect 6085 16370 6120 16404
rect 6154 16370 6189 16404
rect 6223 16370 6258 16404
rect 6292 16370 6327 16404
rect 6361 16370 6396 16404
rect 6430 16370 6465 16404
rect 6499 16370 6534 16404
rect 6568 16370 6603 16404
rect 6637 16370 6672 16404
rect 6706 16370 6741 16404
rect 6775 16370 6810 16404
rect 6844 16370 6879 16404
rect 6913 16370 6948 16404
rect 6982 16370 7017 16404
rect 7051 16370 7086 16404
rect 7120 16370 7155 16404
rect 7189 16370 7224 16404
rect 7258 16370 7293 16404
rect 7327 16370 7362 16404
rect 7396 16370 7431 16404
rect 7465 16370 7500 16404
rect 7534 16370 7568 16404
rect 7602 16370 7636 16404
rect 7670 16370 7704 16404
rect 7738 16370 7772 16404
rect 7806 16370 7840 16404
rect 7874 16370 7908 16404
rect 4681 16347 7908 16370
rect 2704 16334 7908 16347
rect 2704 16300 4740 16334
rect 4774 16300 4809 16334
rect 4843 16300 4878 16334
rect 4912 16300 4947 16334
rect 4981 16300 5016 16334
rect 5050 16300 5085 16334
rect 5119 16300 5154 16334
rect 5188 16300 5223 16334
rect 5257 16300 5292 16334
rect 5326 16300 5361 16334
rect 5395 16300 5430 16334
rect 5464 16300 5499 16334
rect 5533 16300 5568 16334
rect 5602 16300 5637 16334
rect 5671 16300 5706 16334
rect 5740 16300 5775 16334
rect 5809 16300 5844 16334
rect 5878 16300 5913 16334
rect 5947 16300 5982 16334
rect 6016 16300 6051 16334
rect 6085 16300 6120 16334
rect 6154 16300 6189 16334
rect 6223 16300 6258 16334
rect 6292 16300 6327 16334
rect 6361 16300 6396 16334
rect 6430 16300 6465 16334
rect 6499 16300 6534 16334
rect 6568 16300 6603 16334
rect 6637 16300 6672 16334
rect 6706 16300 6741 16334
rect 6775 16300 6810 16334
rect 6844 16300 6879 16334
rect 6913 16300 6948 16334
rect 6982 16300 7017 16334
rect 7051 16300 7086 16334
rect 7120 16300 7155 16334
rect 7189 16300 7224 16334
rect 7258 16300 7293 16334
rect 7327 16300 7362 16334
rect 7396 16300 7431 16334
rect 7465 16300 7500 16334
rect 7534 16300 7568 16334
rect 7602 16300 7636 16334
rect 7670 16300 7704 16334
rect 7738 16300 7772 16334
rect 7806 16300 7840 16334
rect 7874 16300 7908 16334
rect 2704 16264 7908 16300
rect 2704 16244 4740 16264
rect 2704 16210 2715 16244
rect 2749 16210 2853 16244
rect 2887 16210 2991 16244
rect 3025 16210 3129 16244
rect 3163 16210 3267 16244
rect 3301 16210 3405 16244
rect 3439 16210 3543 16244
rect 3577 16210 3681 16244
rect 3715 16210 3819 16244
rect 3853 16210 3957 16244
rect 3991 16210 4095 16244
rect 4129 16210 4233 16244
rect 4267 16210 4371 16244
rect 4405 16210 4509 16244
rect 4543 16210 4647 16244
rect 4681 16230 4740 16244
rect 4774 16230 4809 16264
rect 4843 16230 4878 16264
rect 4912 16230 4947 16264
rect 4981 16230 5016 16264
rect 5050 16230 5085 16264
rect 5119 16230 5154 16264
rect 5188 16230 5223 16264
rect 5257 16230 5292 16264
rect 5326 16230 5361 16264
rect 5395 16230 5430 16264
rect 5464 16230 5499 16264
rect 5533 16230 5568 16264
rect 5602 16230 5637 16264
rect 5671 16230 5706 16264
rect 5740 16230 5775 16264
rect 5809 16230 5844 16264
rect 5878 16230 5913 16264
rect 5947 16230 5982 16264
rect 6016 16230 6051 16264
rect 6085 16230 6120 16264
rect 6154 16230 6189 16264
rect 6223 16230 6258 16264
rect 6292 16230 6327 16264
rect 6361 16230 6396 16264
rect 6430 16230 6465 16264
rect 6499 16230 6534 16264
rect 6568 16230 6603 16264
rect 6637 16230 6672 16264
rect 6706 16230 6741 16264
rect 6775 16230 6810 16264
rect 6844 16230 6879 16264
rect 6913 16230 6948 16264
rect 6982 16230 7017 16264
rect 7051 16230 7086 16264
rect 7120 16230 7155 16264
rect 7189 16230 7224 16264
rect 7258 16230 7293 16264
rect 7327 16230 7362 16264
rect 7396 16230 7431 16264
rect 7465 16230 7500 16264
rect 7534 16230 7568 16264
rect 7602 16230 7636 16264
rect 7670 16230 7704 16264
rect 7738 16230 7772 16264
rect 7806 16230 7840 16264
rect 7874 16230 7908 16264
rect 4681 16210 7908 16230
rect 2704 16194 7908 16210
rect 2704 16160 4740 16194
rect 4774 16160 4809 16194
rect 4843 16160 4878 16194
rect 4912 16160 4947 16194
rect 4981 16160 5016 16194
rect 5050 16160 5085 16194
rect 5119 16160 5154 16194
rect 5188 16160 5223 16194
rect 5257 16160 5292 16194
rect 5326 16160 5361 16194
rect 5395 16160 5430 16194
rect 5464 16160 5499 16194
rect 5533 16160 5568 16194
rect 5602 16160 5637 16194
rect 5671 16160 5706 16194
rect 5740 16160 5775 16194
rect 5809 16160 5844 16194
rect 5878 16160 5913 16194
rect 5947 16160 5982 16194
rect 6016 16160 6051 16194
rect 6085 16160 6120 16194
rect 6154 16160 6189 16194
rect 6223 16160 6258 16194
rect 6292 16160 6327 16194
rect 6361 16160 6396 16194
rect 6430 16160 6465 16194
rect 6499 16160 6534 16194
rect 6568 16160 6603 16194
rect 6637 16160 6672 16194
rect 6706 16160 6741 16194
rect 6775 16160 6810 16194
rect 6844 16160 6879 16194
rect 6913 16160 6948 16194
rect 6982 16160 7017 16194
rect 7051 16160 7086 16194
rect 7120 16160 7155 16194
rect 7189 16160 7224 16194
rect 7258 16160 7293 16194
rect 7327 16160 7362 16194
rect 7396 16160 7431 16194
rect 7465 16160 7500 16194
rect 7534 16160 7568 16194
rect 7602 16160 7636 16194
rect 7670 16160 7704 16194
rect 7738 16160 7772 16194
rect 7806 16160 7840 16194
rect 7874 16160 7908 16194
rect 2704 16124 7908 16160
rect 2704 16107 4740 16124
rect 2704 16073 2715 16107
rect 2749 16073 2853 16107
rect 2887 16073 2991 16107
rect 3025 16073 3129 16107
rect 3163 16073 3267 16107
rect 3301 16073 3405 16107
rect 3439 16073 3543 16107
rect 3577 16073 3681 16107
rect 3715 16073 3819 16107
rect 3853 16073 3957 16107
rect 3991 16073 4095 16107
rect 4129 16073 4233 16107
rect 4267 16073 4371 16107
rect 4405 16073 4509 16107
rect 4543 16073 4647 16107
rect 4681 16090 4740 16107
rect 4774 16090 4809 16124
rect 4843 16090 4878 16124
rect 4912 16090 4947 16124
rect 4981 16090 5016 16124
rect 5050 16090 5085 16124
rect 5119 16090 5154 16124
rect 5188 16090 5223 16124
rect 5257 16090 5292 16124
rect 5326 16090 5361 16124
rect 5395 16090 5430 16124
rect 5464 16090 5499 16124
rect 5533 16090 5568 16124
rect 5602 16090 5637 16124
rect 5671 16090 5706 16124
rect 5740 16090 5775 16124
rect 5809 16090 5844 16124
rect 5878 16090 5913 16124
rect 5947 16090 5982 16124
rect 6016 16090 6051 16124
rect 6085 16090 6120 16124
rect 6154 16090 6189 16124
rect 6223 16090 6258 16124
rect 6292 16090 6327 16124
rect 6361 16090 6396 16124
rect 6430 16090 6465 16124
rect 6499 16090 6534 16124
rect 6568 16090 6603 16124
rect 6637 16090 6672 16124
rect 6706 16090 6741 16124
rect 6775 16090 6810 16124
rect 6844 16090 6879 16124
rect 6913 16090 6948 16124
rect 6982 16090 7017 16124
rect 7051 16090 7086 16124
rect 7120 16090 7155 16124
rect 7189 16090 7224 16124
rect 7258 16090 7293 16124
rect 7327 16090 7362 16124
rect 7396 16090 7431 16124
rect 7465 16090 7500 16124
rect 7534 16090 7568 16124
rect 7602 16090 7636 16124
rect 7670 16090 7704 16124
rect 7738 16090 7772 16124
rect 7806 16090 7840 16124
rect 7874 16090 7908 16124
rect 4681 16073 7908 16090
rect 2704 16054 7908 16073
rect 2704 16020 4740 16054
rect 4774 16020 4809 16054
rect 4843 16020 4878 16054
rect 4912 16020 4947 16054
rect 4981 16020 5016 16054
rect 5050 16020 5085 16054
rect 5119 16020 5154 16054
rect 5188 16020 5223 16054
rect 5257 16020 5292 16054
rect 5326 16020 5361 16054
rect 5395 16020 5430 16054
rect 5464 16020 5499 16054
rect 5533 16020 5568 16054
rect 5602 16020 5637 16054
rect 5671 16020 5706 16054
rect 5740 16020 5775 16054
rect 5809 16020 5844 16054
rect 5878 16020 5913 16054
rect 5947 16020 5982 16054
rect 6016 16020 6051 16054
rect 6085 16020 6120 16054
rect 6154 16020 6189 16054
rect 6223 16020 6258 16054
rect 6292 16020 6327 16054
rect 6361 16020 6396 16054
rect 6430 16020 6465 16054
rect 6499 16020 6534 16054
rect 6568 16020 6603 16054
rect 6637 16020 6672 16054
rect 6706 16020 6741 16054
rect 6775 16020 6810 16054
rect 6844 16020 6879 16054
rect 6913 16020 6948 16054
rect 6982 16020 7017 16054
rect 7051 16020 7086 16054
rect 7120 16020 7155 16054
rect 7189 16020 7224 16054
rect 7258 16020 7293 16054
rect 7327 16020 7362 16054
rect 7396 16020 7431 16054
rect 7465 16020 7500 16054
rect 7534 16020 7568 16054
rect 7602 16020 7636 16054
rect 7670 16020 7704 16054
rect 7738 16020 7772 16054
rect 7806 16020 7840 16054
rect 7874 16020 7908 16054
rect 2704 15984 7908 16020
rect 2704 15970 4740 15984
rect 2704 15936 2715 15970
rect 2749 15936 2853 15970
rect 2887 15936 2991 15970
rect 3025 15936 3129 15970
rect 3163 15936 3267 15970
rect 3301 15936 3405 15970
rect 3439 15936 3543 15970
rect 3577 15936 3681 15970
rect 3715 15936 3819 15970
rect 3853 15936 3957 15970
rect 3991 15936 4095 15970
rect 4129 15936 4233 15970
rect 4267 15936 4371 15970
rect 4405 15936 4509 15970
rect 4543 15936 4647 15970
rect 4681 15950 4740 15970
rect 4774 15950 4809 15984
rect 4843 15950 4878 15984
rect 4912 15950 4947 15984
rect 4981 15950 5016 15984
rect 5050 15950 5085 15984
rect 5119 15950 5154 15984
rect 5188 15950 5223 15984
rect 5257 15950 5292 15984
rect 5326 15950 5361 15984
rect 5395 15950 5430 15984
rect 5464 15950 5499 15984
rect 5533 15950 5568 15984
rect 5602 15950 5637 15984
rect 5671 15950 5706 15984
rect 5740 15950 5775 15984
rect 5809 15950 5844 15984
rect 5878 15950 5913 15984
rect 5947 15950 5982 15984
rect 6016 15950 6051 15984
rect 6085 15950 6120 15984
rect 6154 15950 6189 15984
rect 6223 15950 6258 15984
rect 6292 15950 6327 15984
rect 6361 15950 6396 15984
rect 6430 15950 6465 15984
rect 6499 15950 6534 15984
rect 6568 15950 6603 15984
rect 6637 15950 6672 15984
rect 6706 15950 6741 15984
rect 6775 15950 6810 15984
rect 6844 15950 6879 15984
rect 6913 15950 6948 15984
rect 6982 15950 7017 15984
rect 7051 15950 7086 15984
rect 7120 15950 7155 15984
rect 7189 15950 7224 15984
rect 7258 15950 7293 15984
rect 7327 15950 7362 15984
rect 7396 15950 7431 15984
rect 7465 15950 7500 15984
rect 7534 15950 7568 15984
rect 7602 15950 7636 15984
rect 7670 15950 7704 15984
rect 7738 15950 7772 15984
rect 7806 15950 7840 15984
rect 7874 15950 7908 15984
rect 4681 15936 7908 15950
rect 2704 15912 7908 15936
rect 2274 9919 2444 10004
rect 2274 9885 2298 9919
rect 2332 9885 2367 9919
rect 2401 9885 2436 9919
rect 2470 9885 2505 9919
rect 2539 9885 2574 9919
rect 2608 9885 2643 9919
rect 2677 9885 2712 9919
rect 2746 9885 2781 9919
rect 2815 9885 2850 9919
rect 2884 9885 2919 9919
rect 2953 9885 2988 9919
rect 3022 9885 3057 9919
rect 3091 9885 3126 9919
rect 3160 9885 3195 9919
rect 3229 9885 3264 9919
rect 3298 9885 3333 9919
rect 3367 9885 3401 9919
rect 3435 9885 3469 9919
rect 3503 9885 3537 9919
rect 3571 9885 3605 9919
rect 3639 9885 3673 9919
rect 3707 9885 3741 9919
rect 3775 9885 3809 9919
rect 3843 9885 3877 9919
rect 3911 9885 3945 9919
rect 3979 9885 4013 9919
rect 4047 9885 4081 9919
rect 4115 9885 4149 9919
rect 4183 9885 4217 9919
rect 4251 9885 4285 9919
rect 4319 9885 4353 9919
rect 4387 9885 4421 9919
rect 4455 9885 4489 9919
rect 4523 9885 4557 9919
rect 4591 9885 4625 9919
rect 4659 9885 4693 9919
rect 4727 9885 4761 9919
rect 4795 9885 4829 9919
rect 4863 9885 4897 9919
rect 4931 9885 4965 9919
rect 4999 9885 5033 9919
rect 5067 9885 5101 9919
rect 5135 9885 5169 9919
rect 5203 9885 5237 9919
rect 5271 9885 5305 9919
rect 5339 9885 5373 9919
rect 5407 9885 5441 9919
rect 5475 9885 5509 9919
rect 5543 9885 5577 9919
rect 5611 9885 5645 9919
rect 5679 9885 5713 9919
rect 5747 9885 5781 9919
rect 5815 9885 5849 9919
rect 5883 9885 5917 9919
rect 5951 9885 5985 9919
rect 6019 9885 6053 9919
rect 6087 9885 6121 9919
rect 6155 9885 6189 9919
rect 6223 9885 6257 9919
rect 6291 9885 6325 9919
rect 6359 9885 6393 9919
rect 6427 9885 6461 9919
rect 6495 9885 6529 9919
rect 6563 9885 6597 9919
rect 6631 9885 6665 9919
rect 6699 9885 6733 9919
rect 6767 9885 6801 9919
rect 6835 9885 6869 9919
rect 6903 9885 6937 9919
rect 6971 9885 7005 9919
rect 7039 9885 7073 9919
rect 7107 9885 7141 9919
rect 7175 9885 7209 9919
rect 7243 9885 7277 9919
rect 7311 9885 7345 9919
rect 7379 9885 7413 9919
rect 7447 9885 7481 9919
rect 7515 9885 7549 9919
rect 7583 9885 7617 9919
rect 7651 9885 7685 9919
rect 7719 9885 7753 9919
rect 7787 9885 7821 9919
rect 7855 9885 7889 9919
rect 7923 9885 7957 9919
rect 7991 9885 8025 9919
rect 8195 9885 8219 9953
rect 2280 9396 2304 9430
rect 2338 9396 2373 9430
rect 2407 9396 2442 9430
rect 2476 9396 2511 9430
rect 2545 9396 2580 9430
rect 2614 9396 2649 9430
rect 2683 9396 2718 9430
rect 2752 9396 2787 9430
rect 2821 9396 2856 9430
rect 2890 9396 2925 9430
rect 2959 9396 2994 9430
rect 3028 9396 3062 9430
rect 3096 9396 3130 9430
rect 3164 9396 3198 9430
rect 3232 9396 3266 9430
rect 3300 9396 3334 9430
rect 3368 9396 3402 9430
rect 3436 9396 3470 9430
rect 3504 9396 3538 9430
rect 3572 9396 3606 9430
rect 3640 9396 3674 9430
rect 3708 9396 3742 9430
rect 3776 9396 3810 9430
rect 3844 9396 3878 9430
rect 3912 9396 3946 9430
rect 3980 9396 4014 9430
rect 4048 9396 4082 9430
rect 4116 9396 4150 9430
rect 4184 9396 4218 9430
rect 4252 9396 4286 9430
rect 4320 9396 4354 9430
rect 4388 9396 4422 9430
rect 4456 9396 4490 9430
rect 4524 9396 4558 9430
rect 4592 9396 4626 9430
rect 4660 9396 4694 9430
rect 4728 9396 4762 9430
rect 4796 9396 4830 9430
rect 4864 9396 4898 9430
rect 4932 9396 4966 9430
rect 5000 9396 5034 9430
rect 5068 9396 5102 9430
rect 5136 9396 5170 9430
rect 5204 9396 5238 9430
rect 5272 9396 5306 9430
rect 5340 9396 5374 9430
rect 5408 9396 5442 9430
rect 5476 9396 5510 9430
rect 5544 9396 5578 9430
rect 5612 9396 5646 9430
rect 5680 9396 5714 9430
rect 5748 9396 5782 9430
rect 5816 9396 5850 9430
rect 5884 9396 5918 9430
rect 5952 9396 5986 9430
rect 6020 9396 6054 9430
rect 6088 9396 6122 9430
rect 6156 9396 6190 9430
rect 6224 9396 6258 9430
rect 6292 9396 6326 9430
rect 6360 9396 6394 9430
rect 6428 9396 6462 9430
rect 6496 9396 6530 9430
rect 6564 9396 6598 9430
rect 6632 9396 6666 9430
rect 6700 9396 6734 9430
rect 6768 9396 6802 9430
rect 6836 9396 6870 9430
rect 6904 9396 6938 9430
rect 6972 9396 7006 9430
rect 7040 9396 7074 9430
rect 7108 9396 7142 9430
rect 7176 9396 7210 9430
rect 7244 9396 7278 9430
rect 7312 9396 7346 9430
rect 7380 9396 7414 9430
rect 7448 9396 7521 9430
rect 2280 9362 2334 9396
rect 2280 9328 2290 9362
rect 2324 9328 2334 9362
rect 7487 9370 7521 9396
rect 2280 9294 2334 9328
rect 2280 9260 2290 9294
rect 2324 9260 2334 9294
rect 7487 9302 7521 9336
rect 2280 9226 2334 9260
rect 2280 9192 2290 9226
rect 2324 9192 2334 9226
rect 2280 9158 2334 9192
rect 2280 9124 2290 9158
rect 2324 9124 2334 9158
rect 2280 9090 2334 9124
rect 2280 9056 2290 9090
rect 2324 9056 2334 9090
rect 2280 9022 2334 9056
rect 2280 8988 2290 9022
rect 2324 8988 2334 9022
rect 2280 8954 2334 8988
rect 2280 8920 2290 8954
rect 2324 8920 2334 8954
rect 2280 8886 2334 8920
rect 2280 8852 2290 8886
rect 2324 8852 2334 8886
rect 2280 8818 2334 8852
rect 2280 8784 2290 8818
rect 2324 8784 2334 8818
rect 2280 8750 2334 8784
rect 2280 8716 2290 8750
rect 2324 8716 2334 8750
rect 2280 8682 2334 8716
rect 2280 8648 2290 8682
rect 2324 8648 2334 8682
rect 2280 8614 2334 8648
rect 2280 8580 2290 8614
rect 2324 8580 2334 8614
rect 2280 8546 2334 8580
rect 2280 8512 2290 8546
rect 2324 8512 2334 8546
rect 2280 8478 2334 8512
rect 2280 8444 2290 8478
rect 2324 8444 2334 8478
rect 2280 8410 2334 8444
rect 2280 8376 2290 8410
rect 2324 8376 2334 8410
rect 2280 8342 2334 8376
rect 2280 8308 2290 8342
rect 2324 8308 2334 8342
rect 2280 8274 2334 8308
rect 2280 8240 2290 8274
rect 2324 8240 2334 8274
rect 2280 8206 2334 8240
rect 2280 8172 2290 8206
rect 2324 8172 2334 8206
rect 2280 8138 2334 8172
rect 2280 8104 2290 8138
rect 2324 8104 2334 8138
rect 2280 8070 2334 8104
rect 2280 8036 2290 8070
rect 2324 8036 2334 8070
rect 2280 8002 2334 8036
rect 2280 7968 2290 8002
rect 2324 7968 2334 8002
rect 2280 7934 2334 7968
rect 2280 7900 2290 7934
rect 2324 7900 2334 7934
rect 2280 7866 2334 7900
rect 2280 7832 2290 7866
rect 2324 7832 2334 7866
rect 2280 7798 2334 7832
rect 2280 7764 2290 7798
rect 2324 7764 2334 7798
rect 2280 7730 2334 7764
rect 2280 7696 2290 7730
rect 2324 7696 2334 7730
rect 2280 7681 2334 7696
rect 7487 9234 7521 9268
rect 7487 9166 7521 9200
rect 7487 9098 7521 9132
rect 7487 9030 7521 9064
rect 7487 8962 7521 8996
rect 7487 8894 7521 8928
rect 7487 8826 7521 8860
rect 7487 8758 7521 8792
rect 7487 8690 7521 8724
rect 7487 8622 7521 8656
rect 7487 8554 7521 8588
rect 7487 8486 7521 8520
rect 7487 8418 7521 8452
rect 7487 8350 7521 8384
rect 7487 8282 7521 8316
rect 7487 8214 7521 8248
rect 7487 8146 7521 8180
rect 7487 8078 7521 8112
rect 7487 8010 7521 8044
rect 7487 7942 7521 7976
rect 7487 7874 7521 7908
rect 7487 7806 7521 7840
rect 7487 7738 7521 7772
rect 7487 7681 7521 7704
rect 2280 7662 2358 7681
rect 2280 7628 2290 7662
rect 2324 7647 2358 7662
rect 2392 7647 2427 7681
rect 2461 7647 2496 7681
rect 2530 7647 2565 7681
rect 2599 7647 2634 7681
rect 2668 7647 2703 7681
rect 2737 7647 2772 7681
rect 2806 7647 2841 7681
rect 2875 7647 2910 7681
rect 2944 7647 2979 7681
rect 3013 7647 3048 7681
rect 3082 7647 3117 7681
rect 3151 7647 3186 7681
rect 3220 7647 3255 7681
rect 3289 7647 3324 7681
rect 3358 7647 3393 7681
rect 3427 7647 3462 7681
rect 3496 7647 3531 7681
rect 3565 7647 3600 7681
rect 3634 7647 3669 7681
rect 3703 7647 3738 7681
rect 3772 7647 3807 7681
rect 3841 7647 3875 7681
rect 3909 7647 3943 7681
rect 3977 7647 4011 7681
rect 4045 7647 4079 7681
rect 4113 7647 4147 7681
rect 4181 7647 4215 7681
rect 4249 7647 4283 7681
rect 4317 7647 4351 7681
rect 4385 7647 4419 7681
rect 4453 7647 4487 7681
rect 4521 7647 4555 7681
rect 4589 7647 4623 7681
rect 4657 7647 4691 7681
rect 4725 7647 4759 7681
rect 4793 7647 4827 7681
rect 4861 7647 4895 7681
rect 4929 7647 4963 7681
rect 4997 7647 5031 7681
rect 5065 7647 5099 7681
rect 5133 7647 5167 7681
rect 5201 7647 5235 7681
rect 5269 7647 5303 7681
rect 5337 7647 5371 7681
rect 5405 7647 5439 7681
rect 5473 7647 5507 7681
rect 5541 7647 5575 7681
rect 5609 7647 5643 7681
rect 5677 7647 5711 7681
rect 5745 7647 5779 7681
rect 5813 7647 5847 7681
rect 5881 7647 5915 7681
rect 5949 7647 5983 7681
rect 6017 7647 6051 7681
rect 6085 7647 6119 7681
rect 6153 7647 6187 7681
rect 6221 7647 6255 7681
rect 6289 7647 6323 7681
rect 6357 7647 6391 7681
rect 6425 7647 6459 7681
rect 6493 7647 6527 7681
rect 6561 7647 6595 7681
rect 6629 7647 6663 7681
rect 6697 7647 6731 7681
rect 6765 7647 6799 7681
rect 6833 7647 6867 7681
rect 6901 7647 6935 7681
rect 6969 7647 7003 7681
rect 7037 7647 7071 7681
rect 7105 7647 7139 7681
rect 7173 7647 7207 7681
rect 7241 7647 7275 7681
rect 7309 7647 7343 7681
rect 7377 7647 7411 7681
rect 7445 7670 7521 7681
rect 7445 7647 7487 7670
rect 2324 7628 2334 7647
rect 2280 7594 2334 7628
rect 2280 7560 2290 7594
rect 2324 7560 2334 7594
rect 2280 7526 2334 7560
rect 7487 7602 7521 7636
rect 2280 7492 2290 7526
rect 2324 7492 2334 7526
rect 2280 7458 2334 7492
rect 7487 7534 7521 7568
rect 2280 7424 2290 7458
rect 2324 7424 2334 7458
rect 2280 7390 2334 7424
rect 2280 7356 2290 7390
rect 2324 7356 2334 7390
rect 2280 7322 2334 7356
rect 2280 7288 2290 7322
rect 2324 7288 2334 7322
rect 2280 7254 2334 7288
rect 2280 7220 2290 7254
rect 2324 7220 2334 7254
rect 2280 7186 2334 7220
rect 2280 7152 2290 7186
rect 2324 7152 2334 7186
rect 2280 7118 2334 7152
rect 2280 7084 2290 7118
rect 2324 7084 2334 7118
rect 2280 7050 2334 7084
rect 2280 7016 2290 7050
rect 2324 7016 2334 7050
rect 2280 6982 2334 7016
rect 2280 6948 2290 6982
rect 2324 6948 2334 6982
rect 2280 6914 2334 6948
rect 2280 6880 2290 6914
rect 2324 6880 2334 6914
rect 2280 6846 2334 6880
rect 2280 6812 2290 6846
rect 2324 6812 2334 6846
rect 2280 6778 2334 6812
rect 2280 6744 2290 6778
rect 2324 6744 2334 6778
rect 2280 6710 2334 6744
rect 2280 6676 2290 6710
rect 2324 6676 2334 6710
rect 2280 6642 2334 6676
rect 2280 6608 2290 6642
rect 2324 6608 2334 6642
rect 2280 6574 2334 6608
rect 2280 6540 2290 6574
rect 2324 6540 2334 6574
rect 2280 6506 2334 6540
rect 2280 6472 2290 6506
rect 2324 6472 2334 6506
rect 2280 6438 2334 6472
rect 2280 6404 2290 6438
rect 2324 6404 2334 6438
rect 2280 6370 2334 6404
rect 2280 6336 2290 6370
rect 2324 6336 2334 6370
rect 2280 6302 2334 6336
rect 2280 6268 2290 6302
rect 2324 6268 2334 6302
rect 2280 6234 2334 6268
rect 2280 6200 2290 6234
rect 2324 6200 2334 6234
rect 2280 6166 2334 6200
rect 2280 6132 2290 6166
rect 2324 6132 2334 6166
rect 2280 6098 2334 6132
rect 2280 6064 2290 6098
rect 2324 6064 2334 6098
rect 2280 6030 2334 6064
rect 2280 5996 2290 6030
rect 2324 5996 2334 6030
rect 2280 5962 2334 5996
rect 2280 5928 2290 5962
rect 2324 5928 2334 5962
rect 2280 5894 2334 5928
rect 2280 5860 2290 5894
rect 2324 5860 2334 5894
rect 2280 5841 2334 5860
rect 7487 7466 7521 7500
rect 7487 7398 7521 7432
rect 7487 7330 7521 7364
rect 7487 7262 7521 7296
rect 7487 7194 7521 7228
rect 7487 7126 7521 7160
rect 7487 7058 7521 7092
rect 7487 6990 7521 7024
rect 7487 6922 7521 6956
rect 7487 6854 7521 6888
rect 7487 6786 7521 6820
rect 7487 6718 7521 6752
rect 7487 6650 7521 6684
rect 7487 6582 7521 6616
rect 7487 6514 7521 6548
rect 7487 6446 7521 6480
rect 7487 6378 7521 6412
rect 7487 6310 7521 6344
rect 7487 6242 7521 6276
rect 7487 6174 7521 6208
rect 7487 6106 7521 6140
rect 7487 6038 7521 6072
rect 7487 5970 7521 6004
rect 7487 5902 7521 5936
rect 7487 5841 7521 5868
rect 2280 5826 2358 5841
rect 2280 5792 2290 5826
rect 2324 5807 2358 5826
rect 2392 5807 2427 5841
rect 2461 5807 2496 5841
rect 2530 5807 2565 5841
rect 2599 5807 2634 5841
rect 2668 5807 2703 5841
rect 2737 5807 2772 5841
rect 2806 5807 2841 5841
rect 2875 5807 2910 5841
rect 2944 5807 2979 5841
rect 3013 5807 3048 5841
rect 3082 5807 3117 5841
rect 3151 5807 3186 5841
rect 3220 5807 3255 5841
rect 3289 5807 3324 5841
rect 3358 5807 3393 5841
rect 3427 5807 3462 5841
rect 3496 5807 3531 5841
rect 3565 5807 3600 5841
rect 3634 5807 3669 5841
rect 3703 5807 3737 5841
rect 3771 5807 3805 5841
rect 3839 5807 3873 5841
rect 3907 5807 3941 5841
rect 3975 5807 4009 5841
rect 4043 5807 4077 5841
rect 4111 5807 4145 5841
rect 4179 5807 4213 5841
rect 4247 5807 4281 5841
rect 4315 5807 4349 5841
rect 4383 5807 4417 5841
rect 4451 5807 4485 5841
rect 4519 5807 4553 5841
rect 4587 5807 4621 5841
rect 4655 5807 4689 5841
rect 4723 5807 4757 5841
rect 4791 5807 4825 5841
rect 4859 5807 4893 5841
rect 4927 5807 4961 5841
rect 4995 5807 5029 5841
rect 5063 5807 5097 5841
rect 5131 5807 5165 5841
rect 5199 5807 5233 5841
rect 5267 5807 5301 5841
rect 5335 5807 5369 5841
rect 5403 5807 5437 5841
rect 5471 5807 5505 5841
rect 5539 5807 5573 5841
rect 5607 5807 5641 5841
rect 5675 5807 5709 5841
rect 5743 5807 5777 5841
rect 5811 5807 5845 5841
rect 5879 5807 5913 5841
rect 5947 5807 5981 5841
rect 6015 5807 6049 5841
rect 6083 5807 6117 5841
rect 6151 5807 6185 5841
rect 6219 5807 6253 5841
rect 6287 5807 6321 5841
rect 6355 5807 6389 5841
rect 6423 5807 6457 5841
rect 6491 5807 6525 5841
rect 6559 5807 6593 5841
rect 6627 5807 6661 5841
rect 6695 5807 6729 5841
rect 6763 5807 6797 5841
rect 6831 5807 6865 5841
rect 6899 5807 6933 5841
rect 6967 5807 7001 5841
rect 7035 5807 7069 5841
rect 7103 5807 7137 5841
rect 7171 5807 7205 5841
rect 7239 5807 7273 5841
rect 7307 5807 7341 5841
rect 7375 5807 7409 5841
rect 7443 5834 7521 5841
rect 7443 5807 7487 5834
rect 2324 5792 2334 5807
rect 2280 5758 2334 5792
rect 2280 5724 2290 5758
rect 2324 5724 2334 5758
rect 2280 5690 2334 5724
rect 2280 5656 2290 5690
rect 2324 5656 2334 5690
rect 7487 5766 7521 5800
rect 7487 5698 7521 5732
rect 2280 5622 2334 5656
rect 2280 5588 2290 5622
rect 2324 5588 2334 5622
rect 7487 5630 7521 5664
rect 2280 5554 2334 5588
rect 2280 5520 2290 5554
rect 2324 5520 2334 5554
rect 2280 5486 2334 5520
rect 2280 5452 2290 5486
rect 2324 5452 2334 5486
rect 2280 5418 2334 5452
rect 2280 5384 2290 5418
rect 2324 5384 2334 5418
rect 2280 5350 2334 5384
rect 2280 5316 2290 5350
rect 2324 5316 2334 5350
rect 2280 5282 2334 5316
rect 2280 5248 2290 5282
rect 2324 5248 2334 5282
rect 2280 5214 2334 5248
rect 2280 5180 2290 5214
rect 2324 5180 2334 5214
rect 2280 5146 2334 5180
rect 2280 5112 2290 5146
rect 2324 5112 2334 5146
rect 2280 5078 2334 5112
rect 2280 5044 2290 5078
rect 2324 5044 2334 5078
rect 2280 5010 2334 5044
rect 2280 4976 2290 5010
rect 2324 4976 2334 5010
rect 2280 4942 2334 4976
rect 2280 4908 2290 4942
rect 2324 4908 2334 4942
rect 2280 4874 2334 4908
rect 2280 4840 2290 4874
rect 2324 4840 2334 4874
rect 2280 4806 2334 4840
rect 2280 4772 2290 4806
rect 2324 4772 2334 4806
rect 2280 4738 2334 4772
rect 2280 4704 2290 4738
rect 2324 4704 2334 4738
rect 2280 4670 2334 4704
rect 2280 4636 2290 4670
rect 2324 4636 2334 4670
rect 2280 4602 2334 4636
rect 2280 4568 2290 4602
rect 2324 4568 2334 4602
rect 2280 4534 2334 4568
rect 2280 4500 2290 4534
rect 2324 4500 2334 4534
rect 2280 4466 2334 4500
rect 2280 4432 2290 4466
rect 2324 4432 2334 4466
rect 2280 4398 2334 4432
rect 2280 4364 2290 4398
rect 2324 4364 2334 4398
rect 2280 4330 2334 4364
rect 2280 4296 2290 4330
rect 2324 4296 2334 4330
rect 2280 4262 2334 4296
rect 2280 4228 2290 4262
rect 2324 4228 2334 4262
rect 2280 4194 2334 4228
rect 2280 4160 2290 4194
rect 2324 4160 2334 4194
rect 2280 4126 2334 4160
rect 2280 4092 2290 4126
rect 2324 4092 2334 4126
rect 2280 4058 2334 4092
rect 2280 4024 2290 4058
rect 2324 4024 2334 4058
rect 2280 3930 2334 4024
rect 7487 5562 7521 5596
rect 7487 5494 7521 5528
rect 7487 5426 7521 5460
rect 7487 5358 7521 5392
rect 7487 5290 7521 5324
rect 7487 5222 7521 5256
rect 7487 5154 7521 5188
rect 7487 5086 7521 5120
rect 7487 5018 7521 5052
rect 7487 4950 7521 4984
rect 7487 4882 7521 4916
rect 7487 4814 7521 4848
rect 7487 4746 7521 4780
rect 7487 4678 7521 4712
rect 7487 4610 7521 4644
rect 7487 4542 7521 4576
rect 7487 4474 7521 4508
rect 7487 4406 7521 4440
rect 7487 4338 7521 4372
rect 7487 4270 7521 4304
rect 7487 4202 7521 4236
rect 7487 4134 7521 4168
rect 7487 4066 7521 4100
rect 7487 3998 7521 4032
rect 7487 3930 7521 3964
rect 2280 3907 7521 3930
rect 2280 3873 2314 3907
rect 2348 3873 2382 3907
rect 2416 3873 2450 3907
rect 2484 3873 2518 3907
rect 2552 3873 2586 3907
rect 2620 3873 2654 3907
rect 2688 3873 2722 3907
rect 2756 3873 2790 3907
rect 2824 3873 2858 3907
rect 2892 3873 2926 3907
rect 2960 3873 2994 3907
rect 3028 3873 3062 3907
rect 3096 3873 3130 3907
rect 3164 3873 3198 3907
rect 3232 3873 3266 3907
rect 3300 3873 3334 3907
rect 3368 3873 3402 3907
rect 3436 3873 3470 3907
rect 3504 3873 3538 3907
rect 3572 3873 3606 3907
rect 3640 3873 3674 3907
rect 3708 3873 3742 3907
rect 3776 3873 3810 3907
rect 3844 3873 3878 3907
rect 3912 3873 3946 3907
rect 3980 3873 4014 3907
rect 4048 3873 4082 3907
rect 4116 3873 4150 3907
rect 4184 3873 4218 3907
rect 4252 3873 4286 3907
rect 4320 3873 4354 3907
rect 4388 3873 4422 3907
rect 4456 3873 4490 3907
rect 4524 3873 4558 3907
rect 4592 3873 4626 3907
rect 4660 3873 4694 3907
rect 4728 3873 4762 3907
rect 4796 3873 4830 3907
rect 4864 3873 4898 3907
rect 4932 3873 4966 3907
rect 5000 3873 5034 3907
rect 5068 3873 5102 3907
rect 5136 3873 5170 3907
rect 5204 3873 5238 3907
rect 5272 3873 5306 3907
rect 5340 3873 5374 3907
rect 5408 3873 5442 3907
rect 5476 3873 5510 3907
rect 5544 3873 5578 3907
rect 5612 3873 5646 3907
rect 5680 3873 5714 3907
rect 5748 3873 5782 3907
rect 5816 3873 5850 3907
rect 5884 3873 5918 3907
rect 5952 3873 5986 3907
rect 6020 3873 6054 3907
rect 6088 3873 6122 3907
rect 6156 3873 6190 3907
rect 6224 3873 6258 3907
rect 6292 3873 6326 3907
rect 6360 3873 6394 3907
rect 6428 3873 6462 3907
rect 6496 3873 6530 3907
rect 6564 3873 6598 3907
rect 6632 3873 6666 3907
rect 6700 3873 6734 3907
rect 6768 3873 6802 3907
rect 6836 3873 6870 3907
rect 6904 3873 6938 3907
rect 6972 3873 7006 3907
rect 7040 3873 7074 3907
rect 7108 3873 7142 3907
rect 7176 3873 7210 3907
rect 7244 3873 7278 3907
rect 7312 3873 7346 3907
rect 7380 3873 7414 3907
rect 7448 3873 7521 3907
rect 2280 3850 7521 3873
rect 1831 3126 7904 3127
rect 1831 3092 1855 3126
rect 1889 3092 1992 3126
rect 2026 3092 2129 3126
rect 2163 3092 2266 3126
rect 2300 3092 2403 3126
rect 2437 3092 2540 3126
rect 2574 3092 2677 3126
rect 2711 3092 2814 3126
rect 2848 3092 2950 3126
rect 2984 3092 3086 3126
rect 3120 3092 3222 3126
rect 3256 3092 3358 3126
rect 3392 3092 3494 3126
rect 3528 3092 3630 3126
rect 3664 3092 3766 3126
rect 3800 3092 3902 3126
rect 3936 3092 4038 3126
rect 4072 3092 4174 3126
rect 4208 3092 4310 3126
rect 4344 3092 4446 3126
rect 4480 3092 4582 3126
rect 4616 3092 4718 3126
rect 4752 3092 4854 3126
rect 4888 3092 4990 3126
rect 5024 3092 5126 3126
rect 5160 3092 5262 3126
rect 5296 3092 5398 3126
rect 5432 3092 5534 3126
rect 5568 3092 5670 3126
rect 5704 3092 5806 3126
rect 5840 3092 5942 3126
rect 5976 3092 6078 3126
rect 6112 3092 6214 3126
rect 6248 3092 6350 3126
rect 6384 3092 6486 3126
rect 6520 3092 6622 3126
rect 6656 3092 6758 3126
rect 6792 3092 6894 3126
rect 6928 3092 7030 3126
rect 7064 3092 7166 3126
rect 7200 3092 7302 3126
rect 7336 3092 7438 3126
rect 7472 3092 7574 3126
rect 7608 3092 7710 3126
rect 7744 3092 7846 3126
rect 7880 3092 7904 3126
rect 1831 3010 7904 3092
rect 1831 2976 1855 3010
rect 1889 2976 1992 3010
rect 2026 2976 2129 3010
rect 2163 2976 2266 3010
rect 2300 2976 2403 3010
rect 2437 2976 2540 3010
rect 2574 2976 2677 3010
rect 2711 2976 2814 3010
rect 2848 2976 2950 3010
rect 2984 2976 3086 3010
rect 3120 2976 3222 3010
rect 3256 2976 3358 3010
rect 3392 2976 3494 3010
rect 3528 2976 3630 3010
rect 3664 2976 3766 3010
rect 3800 2976 3902 3010
rect 3936 2976 4038 3010
rect 4072 2976 4174 3010
rect 4208 2976 4310 3010
rect 4344 2976 4446 3010
rect 4480 2976 4582 3010
rect 4616 2976 4718 3010
rect 4752 2976 4854 3010
rect 4888 2976 4990 3010
rect 5024 2976 5126 3010
rect 5160 2976 5262 3010
rect 5296 2976 5398 3010
rect 5432 2976 5534 3010
rect 5568 2976 5670 3010
rect 5704 2976 5806 3010
rect 5840 2976 5942 3010
rect 5976 2976 6078 3010
rect 6112 2976 6214 3010
rect 6248 2976 6350 3010
rect 6384 2976 6486 3010
rect 6520 2976 6622 3010
rect 6656 2976 6758 3010
rect 6792 2976 6894 3010
rect 6928 2976 7030 3010
rect 7064 2976 7166 3010
rect 7200 2976 7302 3010
rect 7336 2976 7438 3010
rect 7472 2976 7574 3010
rect 7608 2976 7710 3010
rect 7744 2976 7846 3010
rect 7880 2976 7904 3010
rect 1831 2894 7904 2976
rect 1831 2860 1855 2894
rect 1889 2860 1992 2894
rect 2026 2860 2129 2894
rect 2163 2860 2266 2894
rect 2300 2860 2403 2894
rect 2437 2860 2540 2894
rect 2574 2860 2677 2894
rect 2711 2860 2814 2894
rect 2848 2860 2950 2894
rect 2984 2860 3086 2894
rect 3120 2860 3222 2894
rect 3256 2860 3358 2894
rect 3392 2860 3494 2894
rect 3528 2860 3630 2894
rect 3664 2860 3766 2894
rect 3800 2860 3902 2894
rect 3936 2860 4038 2894
rect 4072 2860 4174 2894
rect 4208 2860 4310 2894
rect 4344 2860 4446 2894
rect 4480 2860 4582 2894
rect 4616 2860 4718 2894
rect 4752 2860 4854 2894
rect 4888 2860 4990 2894
rect 5024 2860 5126 2894
rect 5160 2860 5262 2894
rect 5296 2860 5398 2894
rect 5432 2860 5534 2894
rect 5568 2860 5670 2894
rect 5704 2860 5806 2894
rect 5840 2860 5942 2894
rect 5976 2860 6078 2894
rect 6112 2860 6214 2894
rect 6248 2860 6350 2894
rect 6384 2860 6486 2894
rect 6520 2860 6622 2894
rect 6656 2860 6758 2894
rect 6792 2860 6894 2894
rect 6928 2860 7030 2894
rect 7064 2860 7166 2894
rect 7200 2860 7302 2894
rect 7336 2860 7438 2894
rect 7472 2860 7574 2894
rect 7608 2860 7710 2894
rect 7744 2860 7846 2894
rect 7880 2860 7904 2894
rect 1831 2778 7904 2860
rect 1831 2744 1855 2778
rect 1889 2744 1992 2778
rect 2026 2744 2129 2778
rect 2163 2744 2266 2778
rect 2300 2744 2403 2778
rect 2437 2744 2540 2778
rect 2574 2744 2677 2778
rect 2711 2744 2814 2778
rect 2848 2744 2950 2778
rect 2984 2744 3086 2778
rect 3120 2744 3222 2778
rect 3256 2744 3358 2778
rect 3392 2744 3494 2778
rect 3528 2744 3630 2778
rect 3664 2744 3766 2778
rect 3800 2744 3902 2778
rect 3936 2744 4038 2778
rect 4072 2744 4174 2778
rect 4208 2744 4310 2778
rect 4344 2744 4446 2778
rect 4480 2744 4582 2778
rect 4616 2744 4718 2778
rect 4752 2744 4854 2778
rect 4888 2744 4990 2778
rect 5024 2744 5126 2778
rect 5160 2744 5262 2778
rect 5296 2744 5398 2778
rect 5432 2744 5534 2778
rect 5568 2744 5670 2778
rect 5704 2744 5806 2778
rect 5840 2744 5942 2778
rect 5976 2744 6078 2778
rect 6112 2744 6214 2778
rect 6248 2744 6350 2778
rect 6384 2744 6486 2778
rect 6520 2744 6622 2778
rect 6656 2744 6758 2778
rect 6792 2744 6894 2778
rect 6928 2744 7030 2778
rect 7064 2744 7166 2778
rect 7200 2744 7302 2778
rect 7336 2744 7438 2778
rect 7472 2744 7574 2778
rect 7608 2744 7710 2778
rect 7744 2744 7846 2778
rect 7880 2744 7904 2778
rect 1831 2662 7904 2744
rect 1831 2628 1855 2662
rect 1889 2628 1992 2662
rect 2026 2628 2129 2662
rect 2163 2628 2266 2662
rect 2300 2628 2403 2662
rect 2437 2628 2540 2662
rect 2574 2628 2677 2662
rect 2711 2628 2814 2662
rect 2848 2628 2950 2662
rect 2984 2628 3086 2662
rect 3120 2628 3222 2662
rect 3256 2628 3358 2662
rect 3392 2628 3494 2662
rect 3528 2628 3630 2662
rect 3664 2628 3766 2662
rect 3800 2628 3902 2662
rect 3936 2628 4038 2662
rect 4072 2628 4174 2662
rect 4208 2628 4310 2662
rect 4344 2628 4446 2662
rect 4480 2628 4582 2662
rect 4616 2628 4718 2662
rect 4752 2628 4854 2662
rect 4888 2628 4990 2662
rect 5024 2628 5126 2662
rect 5160 2628 5262 2662
rect 5296 2628 5398 2662
rect 5432 2628 5534 2662
rect 5568 2628 5670 2662
rect 5704 2628 5806 2662
rect 5840 2628 5942 2662
rect 5976 2628 6078 2662
rect 6112 2628 6214 2662
rect 6248 2628 6350 2662
rect 6384 2628 6486 2662
rect 6520 2628 6622 2662
rect 6656 2628 6758 2662
rect 6792 2628 6894 2662
rect 6928 2628 7030 2662
rect 7064 2628 7166 2662
rect 7200 2628 7302 2662
rect 7336 2628 7438 2662
rect 7472 2628 7574 2662
rect 7608 2628 7710 2662
rect 7744 2628 7846 2662
rect 7880 2628 7904 2662
rect 1831 2546 7904 2628
rect 1831 2512 1855 2546
rect 1889 2512 1992 2546
rect 2026 2512 2129 2546
rect 2163 2512 2266 2546
rect 2300 2512 2403 2546
rect 2437 2512 2540 2546
rect 2574 2512 2677 2546
rect 2711 2512 2814 2546
rect 2848 2512 2950 2546
rect 2984 2512 3086 2546
rect 3120 2512 3222 2546
rect 3256 2512 3358 2546
rect 3392 2512 3494 2546
rect 3528 2512 3630 2546
rect 3664 2512 3766 2546
rect 3800 2512 3902 2546
rect 3936 2512 4038 2546
rect 4072 2512 4174 2546
rect 4208 2512 4310 2546
rect 4344 2512 4446 2546
rect 4480 2512 4582 2546
rect 4616 2512 4718 2546
rect 4752 2512 4854 2546
rect 4888 2512 4990 2546
rect 5024 2512 5126 2546
rect 5160 2512 5262 2546
rect 5296 2512 5398 2546
rect 5432 2512 5534 2546
rect 5568 2512 5670 2546
rect 5704 2512 5806 2546
rect 5840 2512 5942 2546
rect 5976 2512 6078 2546
rect 6112 2512 6214 2546
rect 6248 2512 6350 2546
rect 6384 2512 6486 2546
rect 6520 2512 6622 2546
rect 6656 2512 6758 2546
rect 6792 2512 6894 2546
rect 6928 2512 7030 2546
rect 7064 2512 7166 2546
rect 7200 2512 7302 2546
rect 7336 2512 7438 2546
rect 7472 2512 7574 2546
rect 7608 2512 7710 2546
rect 7744 2512 7846 2546
rect 7880 2512 7904 2546
rect 1831 2430 7904 2512
rect 1831 2396 1855 2430
rect 1889 2396 1992 2430
rect 2026 2396 2129 2430
rect 2163 2396 2266 2430
rect 2300 2396 2403 2430
rect 2437 2396 2540 2430
rect 2574 2396 2677 2430
rect 2711 2396 2814 2430
rect 2848 2396 2950 2430
rect 2984 2396 3086 2430
rect 3120 2396 3222 2430
rect 3256 2396 3358 2430
rect 3392 2396 3494 2430
rect 3528 2396 3630 2430
rect 3664 2396 3766 2430
rect 3800 2396 3902 2430
rect 3936 2396 4038 2430
rect 4072 2396 4174 2430
rect 4208 2396 4310 2430
rect 4344 2396 4446 2430
rect 4480 2396 4582 2430
rect 4616 2396 4718 2430
rect 4752 2396 4854 2430
rect 4888 2396 4990 2430
rect 5024 2396 5126 2430
rect 5160 2396 5262 2430
rect 5296 2396 5398 2430
rect 5432 2396 5534 2430
rect 5568 2396 5670 2430
rect 5704 2396 5806 2430
rect 5840 2396 5942 2430
rect 5976 2396 6078 2430
rect 6112 2396 6214 2430
rect 6248 2396 6350 2430
rect 6384 2396 6486 2430
rect 6520 2396 6622 2430
rect 6656 2396 6758 2430
rect 6792 2396 6894 2430
rect 6928 2396 7030 2430
rect 7064 2396 7166 2430
rect 7200 2396 7302 2430
rect 7336 2396 7438 2430
rect 7472 2396 7574 2430
rect 7608 2396 7710 2430
rect 7744 2396 7846 2430
rect 7880 2396 7904 2430
rect 1831 2395 7904 2396
rect 5340 2361 7594 2395
rect 5340 2327 5346 2361
rect 5380 2327 5484 2361
rect 5518 2327 5622 2361
rect 5656 2327 5760 2361
rect 5794 2327 5898 2361
rect 5932 2327 6036 2361
rect 6070 2327 6174 2361
rect 6208 2327 6312 2361
rect 6346 2327 6450 2361
rect 6484 2327 6588 2361
rect 6622 2327 6726 2361
rect 6760 2327 6864 2361
rect 6898 2327 7002 2361
rect 7036 2327 7140 2361
rect 7174 2327 7278 2361
rect 7312 2327 7416 2361
rect 7450 2327 7554 2361
rect 7588 2327 7594 2361
rect 5340 2223 7594 2327
rect 5340 2189 5346 2223
rect 5380 2189 5484 2223
rect 5518 2189 5622 2223
rect 5656 2189 5760 2223
rect 5794 2189 5898 2223
rect 5932 2189 6036 2223
rect 6070 2189 6174 2223
rect 6208 2189 6312 2223
rect 6346 2189 6450 2223
rect 6484 2189 6588 2223
rect 6622 2189 6726 2223
rect 6760 2189 6864 2223
rect 6898 2189 7002 2223
rect 7036 2189 7140 2223
rect 7174 2189 7278 2223
rect 7312 2189 7416 2223
rect 7450 2189 7554 2223
rect 7588 2189 7594 2223
rect 5340 2085 7594 2189
rect 5340 2051 5346 2085
rect 5380 2051 5484 2085
rect 5518 2051 5622 2085
rect 5656 2051 5760 2085
rect 5794 2051 5898 2085
rect 5932 2051 6036 2085
rect 6070 2051 6174 2085
rect 6208 2051 6312 2085
rect 6346 2051 6450 2085
rect 6484 2051 6588 2085
rect 6622 2051 6726 2085
rect 6760 2051 6864 2085
rect 6898 2051 7002 2085
rect 7036 2051 7140 2085
rect 7174 2051 7278 2085
rect 7312 2051 7416 2085
rect 7450 2051 7554 2085
rect 7588 2051 7594 2085
rect 5340 1947 7594 2051
rect 5340 1913 5346 1947
rect 5380 1913 5484 1947
rect 5518 1913 5622 1947
rect 5656 1913 5760 1947
rect 5794 1913 5898 1947
rect 5932 1913 6036 1947
rect 6070 1913 6174 1947
rect 6208 1913 6312 1947
rect 6346 1913 6450 1947
rect 6484 1913 6588 1947
rect 6622 1913 6726 1947
rect 6760 1913 6864 1947
rect 6898 1913 7002 1947
rect 7036 1913 7140 1947
rect 7174 1913 7278 1947
rect 7312 1913 7416 1947
rect 7450 1913 7554 1947
rect 7588 1913 7594 1947
rect 5340 1809 7594 1913
rect 5340 1775 5346 1809
rect 5380 1775 5484 1809
rect 5518 1775 5622 1809
rect 5656 1775 5760 1809
rect 5794 1775 5898 1809
rect 5932 1775 6036 1809
rect 6070 1775 6174 1809
rect 6208 1775 6312 1809
rect 6346 1775 6450 1809
rect 6484 1775 6588 1809
rect 6622 1775 6726 1809
rect 6760 1775 6864 1809
rect 6898 1775 7002 1809
rect 7036 1775 7140 1809
rect 7174 1775 7278 1809
rect 7312 1775 7416 1809
rect 7450 1775 7554 1809
rect 7588 1775 7594 1809
rect 5340 1671 7594 1775
rect 5340 1637 5346 1671
rect 5380 1637 5484 1671
rect 5518 1637 5622 1671
rect 5656 1637 5760 1671
rect 5794 1637 5898 1671
rect 5932 1637 6036 1671
rect 6070 1637 6174 1671
rect 6208 1637 6312 1671
rect 6346 1637 6450 1671
rect 6484 1637 6588 1671
rect 6622 1637 6726 1671
rect 6760 1637 6864 1671
rect 6898 1637 7002 1671
rect 7036 1637 7140 1671
rect 7174 1637 7278 1671
rect 7312 1637 7416 1671
rect 7450 1637 7554 1671
rect 7588 1637 7594 1671
rect 5340 1532 7594 1637
rect 5340 1498 5346 1532
rect 5380 1498 5484 1532
rect 5518 1498 5622 1532
rect 5656 1498 5760 1532
rect 5794 1498 5898 1532
rect 5932 1498 6036 1532
rect 6070 1498 6174 1532
rect 6208 1498 6312 1532
rect 6346 1498 6450 1532
rect 6484 1498 6588 1532
rect 6622 1498 6726 1532
rect 6760 1498 6864 1532
rect 6898 1498 7002 1532
rect 7036 1498 7140 1532
rect 7174 1498 7278 1532
rect 7312 1498 7416 1532
rect 7450 1498 7554 1532
rect 7588 1498 7594 1532
rect 5340 1393 7594 1498
rect 5340 1359 5346 1393
rect 5380 1359 5484 1393
rect 5518 1359 5622 1393
rect 5656 1359 5760 1393
rect 5794 1359 5898 1393
rect 5932 1359 6036 1393
rect 6070 1359 6174 1393
rect 6208 1359 6312 1393
rect 6346 1359 6450 1393
rect 6484 1359 6588 1393
rect 6622 1359 6726 1393
rect 6760 1359 6864 1393
rect 6898 1359 7002 1393
rect 7036 1359 7140 1393
rect 7174 1359 7278 1393
rect 7312 1359 7416 1393
rect 7450 1359 7554 1393
rect 7588 1359 7594 1393
rect 5340 1254 7594 1359
rect 5340 1220 5346 1254
rect 5380 1220 5484 1254
rect 5518 1220 5622 1254
rect 5656 1220 5760 1254
rect 5794 1220 5898 1254
rect 5932 1220 6036 1254
rect 6070 1220 6174 1254
rect 6208 1220 6312 1254
rect 6346 1220 6450 1254
rect 6484 1220 6588 1254
rect 6622 1220 6726 1254
rect 6760 1220 6864 1254
rect 6898 1220 7002 1254
rect 7036 1220 7140 1254
rect 7174 1220 7278 1254
rect 7312 1220 7416 1254
rect 7450 1220 7554 1254
rect 7588 1220 7594 1254
rect 5340 1115 7594 1220
rect 5340 1081 5346 1115
rect 5380 1081 5484 1115
rect 5518 1081 5622 1115
rect 5656 1081 5760 1115
rect 5794 1081 5898 1115
rect 5932 1081 6036 1115
rect 6070 1081 6174 1115
rect 6208 1081 6312 1115
rect 6346 1081 6450 1115
rect 6484 1081 6588 1115
rect 6622 1081 6726 1115
rect 6760 1081 6864 1115
rect 6898 1081 7002 1115
rect 7036 1081 7140 1115
rect 7174 1081 7278 1115
rect 7312 1081 7416 1115
rect 7450 1081 7554 1115
rect 7588 1081 7594 1115
rect 5340 976 7594 1081
rect 5340 942 5346 976
rect 5380 942 5484 976
rect 5518 942 5622 976
rect 5656 942 5760 976
rect 5794 942 5898 976
rect 5932 942 6036 976
rect 6070 942 6174 976
rect 6208 942 6312 976
rect 6346 942 6450 976
rect 6484 942 6588 976
rect 6622 942 6726 976
rect 6760 942 6864 976
rect 6898 942 7002 976
rect 7036 942 7140 976
rect 7174 942 7278 976
rect 7312 942 7416 976
rect 7450 942 7554 976
rect 7588 942 7594 976
rect 5340 837 7594 942
rect 5340 803 5346 837
rect 5380 803 5484 837
rect 5518 803 5622 837
rect 5656 803 5760 837
rect 5794 803 5898 837
rect 5932 803 6036 837
rect 6070 803 6174 837
rect 6208 803 6312 837
rect 6346 803 6450 837
rect 6484 803 6588 837
rect 6622 803 6726 837
rect 6760 803 6864 837
rect 6898 803 7002 837
rect 7036 803 7140 837
rect 7174 803 7278 837
rect 7312 803 7416 837
rect 7450 803 7554 837
rect 7588 803 7594 837
rect 5340 698 7594 803
rect 5340 664 5346 698
rect 5380 664 5484 698
rect 5518 664 5622 698
rect 5656 664 5760 698
rect 5794 664 5898 698
rect 5932 664 6036 698
rect 6070 664 6174 698
rect 6208 664 6312 698
rect 6346 664 6450 698
rect 6484 664 6588 698
rect 6622 664 6726 698
rect 6760 664 6864 698
rect 6898 664 7002 698
rect 7036 664 7140 698
rect 7174 664 7278 698
rect 7312 664 7416 698
rect 7450 664 7554 698
rect 7588 664 7594 698
rect 5340 559 7594 664
rect 5340 525 5346 559
rect 5380 525 5484 559
rect 5518 525 5622 559
rect 5656 525 5760 559
rect 5794 525 5898 559
rect 5932 525 6036 559
rect 6070 525 6174 559
rect 6208 525 6312 559
rect 6346 525 6450 559
rect 6484 525 6588 559
rect 6622 525 6726 559
rect 6760 525 6864 559
rect 6898 525 7002 559
rect 7036 525 7140 559
rect 7174 525 7278 559
rect 7312 525 7416 559
rect 7450 525 7554 559
rect 7588 525 7594 559
rect 5340 420 7594 525
rect 5340 386 5346 420
rect 5380 386 5484 420
rect 5518 386 5622 420
rect 5656 386 5760 420
rect 5794 386 5898 420
rect 5932 386 6036 420
rect 6070 386 6174 420
rect 6208 386 6312 420
rect 6346 386 6450 420
rect 6484 386 6588 420
rect 6622 386 6726 420
rect 6760 386 6864 420
rect 6898 386 7002 420
rect 7036 386 7140 420
rect 7174 386 7278 420
rect 7312 386 7416 420
rect 7450 386 7554 420
rect 7588 386 7594 420
rect 5340 352 7594 386
<< nsubdiff >>
rect 1801 1982 1869 2016
rect 1903 1982 1937 2016
rect 1971 1982 2005 2016
rect 2039 1982 2073 2016
rect 2107 1982 2141 2016
rect 2175 1982 2209 2016
rect 2243 1982 2277 2016
rect 2311 1982 2345 2016
rect 2379 1982 2413 2016
rect 2447 1982 2481 2016
rect 2515 1982 2549 2016
rect 2583 1982 2617 2016
rect 2651 1982 2685 2016
rect 2719 1982 2753 2016
rect 2787 1982 2821 2016
rect 2855 1982 2889 2016
rect 2923 1982 2957 2016
rect 2991 1982 3025 2016
rect 3059 1982 3093 2016
rect 3127 1982 3161 2016
rect 3195 1982 3229 2016
rect 3263 1982 3297 2016
rect 3331 1982 3365 2016
rect 3399 1982 3433 2016
rect 3467 1982 3501 2016
rect 3535 1982 3569 2016
rect 3603 1982 3637 2016
rect 3671 1982 3705 2016
rect 3739 1982 3773 2016
rect 3807 1982 3841 2016
rect 3875 1982 3909 2016
rect 3943 1982 3977 2016
rect 4011 1982 4045 2016
rect 4079 1982 4113 2016
rect 4147 1982 4181 2016
rect 4215 1982 4249 2016
rect 4283 1982 4317 2016
rect 4351 1982 4385 2016
rect 4419 1982 4453 2016
rect 4487 1982 4521 2016
rect 4555 1982 4589 2016
rect 4623 1982 4657 2016
rect 4691 1982 4725 2016
rect 4759 1982 4793 2016
rect 4827 1982 4861 2016
rect 4895 1982 4929 2016
rect 4963 1982 5039 2016
rect 1801 1918 1835 1982
rect 1801 1850 1835 1884
rect 5005 1948 5039 1982
rect 5005 1880 5039 1914
rect 1801 1782 1835 1816
rect 1801 1714 1835 1748
rect 1801 1646 1835 1680
rect 1801 1578 1835 1612
rect 1801 1510 1835 1544
rect 1801 1442 1835 1476
rect 1801 1374 1835 1408
rect 1801 1306 1835 1340
rect 1801 1238 1835 1272
rect 1801 1170 1835 1204
rect 1801 1102 1835 1136
rect 1801 1034 1835 1068
rect 5005 1812 5039 1846
rect 5005 1744 5039 1778
rect 5005 1676 5039 1710
rect 5005 1608 5039 1642
rect 5005 1540 5039 1574
rect 5005 1472 5039 1506
rect 5005 1404 5039 1438
rect 5005 1336 5039 1370
rect 5005 1268 5039 1302
rect 5005 1200 5039 1234
rect 5005 1132 5039 1166
rect 5005 1064 5039 1098
rect 1801 966 1835 1000
rect 1801 898 1835 932
rect 5005 996 5039 1030
rect 5005 898 5039 962
rect 1801 864 1945 898
rect 1979 864 2013 898
rect 2047 864 2081 898
rect 2115 864 2149 898
rect 2183 864 2217 898
rect 2251 864 2285 898
rect 2319 864 2353 898
rect 2387 864 2421 898
rect 2455 864 2489 898
rect 2523 864 2557 898
rect 2591 864 2625 898
rect 2659 864 2693 898
rect 2727 864 2761 898
rect 2795 864 2829 898
rect 2863 864 2897 898
rect 2931 864 2965 898
rect 2999 864 3033 898
rect 3067 864 3101 898
rect 3135 864 3169 898
rect 3203 864 3237 898
rect 3271 864 3305 898
rect 3339 864 3373 898
rect 3407 864 3441 898
rect 3475 864 3509 898
rect 3543 864 3577 898
rect 3611 864 3645 898
rect 3679 864 3713 898
rect 3747 864 3781 898
rect 3815 864 3849 898
rect 3883 864 3917 898
rect 3951 864 3985 898
rect 4019 864 4053 898
rect 4087 864 4121 898
rect 4155 864 4189 898
rect 4223 864 4257 898
rect 4291 864 4325 898
rect 4359 864 4393 898
rect 4427 864 4461 898
rect 4495 864 4529 898
rect 4563 864 4597 898
rect 4631 864 4665 898
rect 4699 864 4733 898
rect 4767 864 4801 898
rect 4835 864 4869 898
rect 4903 864 4937 898
rect 4971 864 5039 898
<< mvnsubdiff >>
rect 1946 39440 2039 39474
rect 2073 39440 2107 39474
rect 1946 39406 2107 39440
rect 2048 39372 2107 39406
rect 8465 39372 8533 39474
rect 8431 39354 8533 39372
rect 8431 39320 8499 39354
rect 8431 39286 8533 39320
rect 2048 9595 2208 9697
rect 7546 9638 8431 9697
rect 7546 9595 7803 9638
rect 7735 9536 7803 9595
rect 8381 9604 8431 9638
rect 8381 9570 8533 9604
rect 8381 9536 8415 9570
rect 8449 9536 8533 9570
rect 7735 9513 7837 9536
rect 7769 9479 7837 9513
rect 7735 9445 7837 9479
rect 1946 3927 2048 4080
rect 7735 4063 7837 4175
rect 2048 3417 2088 3451
rect 1946 3383 2088 3417
rect 1946 3349 2020 3383
rect 2054 3349 2088 3383
rect 2598 3349 2666 3451
rect 7120 3349 7235 3451
rect 7677 3417 7735 3451
rect 7677 3383 7837 3417
rect 7677 3349 7711 3383
rect 7745 3349 7837 3383
<< psubdiffcont >>
rect 2405 39108 2439 39142
rect 2274 39006 2376 39074
rect 2473 39040 8151 39142
rect 2274 10004 2444 39006
rect 2541 38972 8083 39040
rect 8185 38989 8219 39023
rect 8117 38887 8219 38955
rect 2715 28924 2749 28958
rect 2853 28924 2887 28958
rect 2991 28924 3025 28958
rect 3129 28924 3163 28958
rect 3267 28924 3301 28958
rect 3405 28924 3439 28958
rect 3543 28924 3577 28958
rect 3681 28924 3715 28958
rect 3819 28924 3853 28958
rect 3957 28924 3991 28958
rect 4095 28924 4129 28958
rect 4233 28924 4267 28958
rect 4371 28924 4405 28958
rect 4509 28924 4543 28958
rect 4647 28924 4681 28958
rect 2715 28788 2749 28822
rect 2853 28788 2887 28822
rect 2991 28788 3025 28822
rect 3129 28788 3163 28822
rect 3267 28788 3301 28822
rect 3405 28788 3439 28822
rect 3543 28788 3577 28822
rect 3681 28788 3715 28822
rect 3819 28788 3853 28822
rect 3957 28788 3991 28822
rect 4095 28788 4129 28822
rect 4233 28788 4267 28822
rect 4371 28788 4405 28822
rect 4509 28788 4543 28822
rect 4647 28788 4681 28822
rect 2715 28652 2749 28686
rect 2853 28652 2887 28686
rect 2991 28652 3025 28686
rect 3129 28652 3163 28686
rect 3267 28652 3301 28686
rect 3405 28652 3439 28686
rect 3543 28652 3577 28686
rect 3681 28652 3715 28686
rect 3819 28652 3853 28686
rect 3957 28652 3991 28686
rect 4095 28652 4129 28686
rect 4233 28652 4267 28686
rect 4371 28652 4405 28686
rect 4509 28652 4543 28686
rect 4647 28652 4681 28686
rect 2715 28516 2749 28550
rect 2853 28516 2887 28550
rect 2991 28516 3025 28550
rect 3129 28516 3163 28550
rect 3267 28516 3301 28550
rect 3405 28516 3439 28550
rect 3543 28516 3577 28550
rect 3681 28516 3715 28550
rect 3819 28516 3853 28550
rect 3957 28516 3991 28550
rect 4095 28516 4129 28550
rect 4233 28516 4267 28550
rect 4371 28516 4405 28550
rect 4509 28516 4543 28550
rect 4647 28516 4681 28550
rect 2715 28380 2749 28414
rect 2853 28380 2887 28414
rect 2991 28380 3025 28414
rect 3129 28380 3163 28414
rect 3267 28380 3301 28414
rect 3405 28380 3439 28414
rect 3543 28380 3577 28414
rect 3681 28380 3715 28414
rect 3819 28380 3853 28414
rect 3957 28380 3991 28414
rect 4095 28380 4129 28414
rect 4233 28380 4267 28414
rect 4371 28380 4405 28414
rect 4509 28380 4543 28414
rect 4647 28380 4681 28414
rect 2715 28244 2749 28278
rect 2853 28244 2887 28278
rect 2991 28244 3025 28278
rect 3129 28244 3163 28278
rect 3267 28244 3301 28278
rect 3405 28244 3439 28278
rect 3543 28244 3577 28278
rect 3681 28244 3715 28278
rect 3819 28244 3853 28278
rect 3957 28244 3991 28278
rect 4095 28244 4129 28278
rect 4233 28244 4267 28278
rect 4371 28244 4405 28278
rect 4509 28244 4543 28278
rect 4647 28244 4681 28278
rect 2715 28108 2749 28142
rect 2853 28108 2887 28142
rect 2991 28108 3025 28142
rect 3129 28108 3163 28142
rect 3267 28108 3301 28142
rect 3405 28108 3439 28142
rect 3543 28108 3577 28142
rect 3681 28108 3715 28142
rect 3819 28108 3853 28142
rect 3957 28108 3991 28142
rect 4095 28108 4129 28142
rect 4233 28108 4267 28142
rect 4371 28108 4405 28142
rect 4509 28108 4543 28142
rect 4647 28108 4681 28142
rect 2715 27972 2749 28006
rect 2853 27972 2887 28006
rect 2991 27972 3025 28006
rect 3129 27972 3163 28006
rect 3267 27972 3301 28006
rect 3405 27972 3439 28006
rect 3543 27972 3577 28006
rect 3681 27972 3715 28006
rect 3819 27972 3853 28006
rect 3957 27972 3991 28006
rect 4095 27972 4129 28006
rect 4233 27972 4267 28006
rect 4371 27972 4405 28006
rect 4509 27972 4543 28006
rect 4647 27972 4681 28006
rect 2715 27836 2749 27870
rect 2853 27836 2887 27870
rect 2991 27836 3025 27870
rect 3129 27836 3163 27870
rect 3267 27836 3301 27870
rect 3405 27836 3439 27870
rect 3543 27836 3577 27870
rect 3681 27836 3715 27870
rect 3819 27836 3853 27870
rect 3957 27836 3991 27870
rect 4095 27836 4129 27870
rect 4233 27836 4267 27870
rect 4371 27836 4405 27870
rect 4509 27836 4543 27870
rect 4647 27836 4681 27870
rect 2715 27700 2749 27734
rect 2853 27700 2887 27734
rect 2991 27700 3025 27734
rect 3129 27700 3163 27734
rect 3267 27700 3301 27734
rect 3405 27700 3439 27734
rect 3543 27700 3577 27734
rect 3681 27700 3715 27734
rect 3819 27700 3853 27734
rect 3957 27700 3991 27734
rect 4095 27700 4129 27734
rect 4233 27700 4267 27734
rect 4371 27700 4405 27734
rect 4509 27700 4543 27734
rect 4647 27700 4681 27734
rect 2715 27564 2749 27598
rect 2853 27564 2887 27598
rect 2991 27564 3025 27598
rect 3129 27564 3163 27598
rect 3267 27564 3301 27598
rect 3405 27564 3439 27598
rect 3543 27564 3577 27598
rect 3681 27564 3715 27598
rect 3819 27564 3853 27598
rect 3957 27564 3991 27598
rect 4095 27564 4129 27598
rect 4233 27564 4267 27598
rect 4371 27564 4405 27598
rect 4509 27564 4543 27598
rect 4647 27564 4681 27598
rect 2715 27428 2749 27462
rect 2853 27428 2887 27462
rect 2991 27428 3025 27462
rect 3129 27428 3163 27462
rect 3267 27428 3301 27462
rect 3405 27428 3439 27462
rect 3543 27428 3577 27462
rect 3681 27428 3715 27462
rect 3819 27428 3853 27462
rect 3957 27428 3991 27462
rect 4095 27428 4129 27462
rect 4233 27428 4267 27462
rect 4371 27428 4405 27462
rect 4509 27428 4543 27462
rect 4647 27428 4681 27462
rect 2715 27292 2749 27326
rect 2853 27292 2887 27326
rect 2991 27292 3025 27326
rect 3129 27292 3163 27326
rect 3267 27292 3301 27326
rect 3405 27292 3439 27326
rect 3543 27292 3577 27326
rect 3681 27292 3715 27326
rect 3819 27292 3853 27326
rect 3957 27292 3991 27326
rect 4095 27292 4129 27326
rect 4233 27292 4267 27326
rect 4371 27292 4405 27326
rect 4509 27292 4543 27326
rect 4647 27292 4681 27326
rect 2715 27156 2749 27190
rect 2853 27156 2887 27190
rect 2991 27156 3025 27190
rect 3129 27156 3163 27190
rect 3267 27156 3301 27190
rect 3405 27156 3439 27190
rect 3543 27156 3577 27190
rect 3681 27156 3715 27190
rect 3819 27156 3853 27190
rect 3957 27156 3991 27190
rect 4095 27156 4129 27190
rect 4233 27156 4267 27190
rect 4371 27156 4405 27190
rect 4509 27156 4543 27190
rect 4647 27156 4681 27190
rect 2715 27020 2749 27054
rect 2853 27020 2887 27054
rect 2991 27020 3025 27054
rect 3129 27020 3163 27054
rect 3267 27020 3301 27054
rect 3405 27020 3439 27054
rect 3543 27020 3577 27054
rect 3681 27020 3715 27054
rect 3819 27020 3853 27054
rect 3957 27020 3991 27054
rect 4095 27020 4129 27054
rect 4233 27020 4267 27054
rect 4371 27020 4405 27054
rect 4509 27020 4543 27054
rect 4647 27020 4681 27054
rect 2715 26884 2749 26918
rect 2853 26884 2887 26918
rect 2991 26884 3025 26918
rect 3129 26884 3163 26918
rect 3267 26884 3301 26918
rect 3405 26884 3439 26918
rect 3543 26884 3577 26918
rect 3681 26884 3715 26918
rect 3819 26884 3853 26918
rect 3957 26884 3991 26918
rect 4095 26884 4129 26918
rect 4233 26884 4267 26918
rect 4371 26884 4405 26918
rect 4509 26884 4543 26918
rect 4647 26884 4681 26918
rect 2715 26748 2749 26782
rect 2853 26748 2887 26782
rect 2991 26748 3025 26782
rect 3129 26748 3163 26782
rect 3267 26748 3301 26782
rect 3405 26748 3439 26782
rect 3543 26748 3577 26782
rect 3681 26748 3715 26782
rect 3819 26748 3853 26782
rect 3957 26748 3991 26782
rect 4095 26748 4129 26782
rect 4233 26748 4267 26782
rect 4371 26748 4405 26782
rect 4509 26748 4543 26782
rect 4647 26748 4681 26782
rect 2715 26612 2749 26646
rect 2853 26612 2887 26646
rect 2991 26612 3025 26646
rect 3129 26612 3163 26646
rect 3267 26612 3301 26646
rect 3405 26612 3439 26646
rect 3543 26612 3577 26646
rect 3681 26612 3715 26646
rect 3819 26612 3853 26646
rect 3957 26612 3991 26646
rect 4095 26612 4129 26646
rect 4233 26612 4267 26646
rect 4371 26612 4405 26646
rect 4509 26612 4543 26646
rect 4647 26612 4681 26646
rect 2715 26476 2749 26510
rect 2853 26476 2887 26510
rect 2991 26476 3025 26510
rect 3129 26476 3163 26510
rect 3267 26476 3301 26510
rect 3405 26476 3439 26510
rect 3543 26476 3577 26510
rect 3681 26476 3715 26510
rect 3819 26476 3853 26510
rect 3957 26476 3991 26510
rect 4095 26476 4129 26510
rect 4233 26476 4267 26510
rect 4371 26476 4405 26510
rect 4509 26476 4543 26510
rect 4647 26476 4681 26510
rect 2715 26340 2749 26374
rect 2853 26340 2887 26374
rect 2991 26340 3025 26374
rect 3129 26340 3163 26374
rect 3267 26340 3301 26374
rect 3405 26340 3439 26374
rect 3543 26340 3577 26374
rect 3681 26340 3715 26374
rect 3819 26340 3853 26374
rect 3957 26340 3991 26374
rect 4095 26340 4129 26374
rect 4233 26340 4267 26374
rect 4371 26340 4405 26374
rect 4509 26340 4543 26374
rect 4647 26340 4681 26374
rect 2715 26204 2749 26238
rect 2853 26204 2887 26238
rect 2991 26204 3025 26238
rect 3129 26204 3163 26238
rect 3267 26204 3301 26238
rect 3405 26204 3439 26238
rect 3543 26204 3577 26238
rect 3681 26204 3715 26238
rect 3819 26204 3853 26238
rect 3957 26204 3991 26238
rect 4095 26204 4129 26238
rect 4233 26204 4267 26238
rect 4371 26204 4405 26238
rect 4509 26204 4543 26238
rect 4647 26204 4681 26238
rect 2715 26068 2749 26102
rect 2853 26068 2887 26102
rect 2991 26068 3025 26102
rect 3129 26068 3163 26102
rect 3267 26068 3301 26102
rect 3405 26068 3439 26102
rect 3543 26068 3577 26102
rect 3681 26068 3715 26102
rect 3819 26068 3853 26102
rect 3957 26068 3991 26102
rect 4095 26068 4129 26102
rect 4233 26068 4267 26102
rect 4371 26068 4405 26102
rect 4509 26068 4543 26102
rect 4647 26068 4681 26102
rect 2715 25932 2749 25966
rect 2853 25932 2887 25966
rect 2991 25932 3025 25966
rect 3129 25932 3163 25966
rect 3267 25932 3301 25966
rect 3405 25932 3439 25966
rect 3543 25932 3577 25966
rect 3681 25932 3715 25966
rect 3819 25932 3853 25966
rect 3957 25932 3991 25966
rect 4095 25932 4129 25966
rect 4233 25932 4267 25966
rect 4371 25932 4405 25966
rect 4509 25932 4543 25966
rect 4647 25932 4681 25966
rect 2715 25796 2749 25830
rect 2853 25796 2887 25830
rect 2991 25796 3025 25830
rect 3129 25796 3163 25830
rect 3267 25796 3301 25830
rect 3405 25796 3439 25830
rect 3543 25796 3577 25830
rect 3681 25796 3715 25830
rect 3819 25796 3853 25830
rect 3957 25796 3991 25830
rect 4095 25796 4129 25830
rect 4233 25796 4267 25830
rect 4371 25796 4405 25830
rect 4509 25796 4543 25830
rect 4647 25796 4681 25830
rect 2715 25660 2749 25694
rect 2853 25660 2887 25694
rect 2991 25660 3025 25694
rect 3129 25660 3163 25694
rect 3267 25660 3301 25694
rect 3405 25660 3439 25694
rect 3543 25660 3577 25694
rect 3681 25660 3715 25694
rect 3819 25660 3853 25694
rect 3957 25660 3991 25694
rect 4095 25660 4129 25694
rect 4233 25660 4267 25694
rect 4371 25660 4405 25694
rect 4509 25660 4543 25694
rect 4647 25660 4681 25694
rect 2715 25524 2749 25558
rect 2853 25524 2887 25558
rect 2991 25524 3025 25558
rect 3129 25524 3163 25558
rect 3267 25524 3301 25558
rect 3405 25524 3439 25558
rect 3543 25524 3577 25558
rect 3681 25524 3715 25558
rect 3819 25524 3853 25558
rect 3957 25524 3991 25558
rect 4095 25524 4129 25558
rect 4233 25524 4267 25558
rect 4371 25524 4405 25558
rect 4509 25524 4543 25558
rect 4647 25524 4681 25558
rect 2715 25388 2749 25422
rect 2853 25388 2887 25422
rect 2991 25388 3025 25422
rect 3129 25388 3163 25422
rect 3267 25388 3301 25422
rect 3405 25388 3439 25422
rect 3543 25388 3577 25422
rect 3681 25388 3715 25422
rect 3819 25388 3853 25422
rect 3957 25388 3991 25422
rect 4095 25388 4129 25422
rect 4233 25388 4267 25422
rect 4371 25388 4405 25422
rect 4509 25388 4543 25422
rect 4647 25388 4681 25422
rect 2715 25252 2749 25286
rect 2853 25252 2887 25286
rect 2991 25252 3025 25286
rect 3129 25252 3163 25286
rect 3267 25252 3301 25286
rect 3405 25252 3439 25286
rect 3543 25252 3577 25286
rect 3681 25252 3715 25286
rect 3819 25252 3853 25286
rect 3957 25252 3991 25286
rect 4095 25252 4129 25286
rect 4233 25252 4267 25286
rect 4371 25252 4405 25286
rect 4509 25252 4543 25286
rect 4647 25252 4681 25286
rect 2715 25115 2749 25149
rect 2853 25115 2887 25149
rect 2991 25115 3025 25149
rect 3129 25115 3163 25149
rect 3267 25115 3301 25149
rect 3405 25115 3439 25149
rect 3543 25115 3577 25149
rect 3681 25115 3715 25149
rect 3819 25115 3853 25149
rect 3957 25115 3991 25149
rect 4095 25115 4129 25149
rect 4233 25115 4267 25149
rect 4371 25115 4405 25149
rect 4509 25115 4543 25149
rect 4647 25115 4681 25149
rect 2715 24978 2749 25012
rect 2853 24978 2887 25012
rect 2991 24978 3025 25012
rect 3129 24978 3163 25012
rect 3267 24978 3301 25012
rect 3405 24978 3439 25012
rect 3543 24978 3577 25012
rect 3681 24978 3715 25012
rect 3819 24978 3853 25012
rect 3957 24978 3991 25012
rect 4095 24978 4129 25012
rect 4233 24978 4267 25012
rect 4371 24978 4405 25012
rect 4509 24978 4543 25012
rect 4647 24978 4681 25012
rect 2715 24841 2749 24875
rect 2853 24841 2887 24875
rect 2991 24841 3025 24875
rect 3129 24841 3163 24875
rect 3267 24841 3301 24875
rect 3405 24841 3439 24875
rect 3543 24841 3577 24875
rect 3681 24841 3715 24875
rect 3819 24841 3853 24875
rect 3957 24841 3991 24875
rect 4095 24841 4129 24875
rect 4233 24841 4267 24875
rect 4371 24841 4405 24875
rect 4509 24841 4543 24875
rect 4647 24841 4681 24875
rect 2715 24704 2749 24738
rect 2853 24704 2887 24738
rect 2991 24704 3025 24738
rect 3129 24704 3163 24738
rect 3267 24704 3301 24738
rect 3405 24704 3439 24738
rect 3543 24704 3577 24738
rect 3681 24704 3715 24738
rect 3819 24704 3853 24738
rect 3957 24704 3991 24738
rect 4095 24704 4129 24738
rect 4233 24704 4267 24738
rect 4371 24704 4405 24738
rect 4509 24704 4543 24738
rect 4647 24704 4681 24738
rect 2715 24567 2749 24601
rect 2853 24567 2887 24601
rect 2991 24567 3025 24601
rect 3129 24567 3163 24601
rect 3267 24567 3301 24601
rect 3405 24567 3439 24601
rect 3543 24567 3577 24601
rect 3681 24567 3715 24601
rect 3819 24567 3853 24601
rect 3957 24567 3991 24601
rect 4095 24567 4129 24601
rect 4233 24567 4267 24601
rect 4371 24567 4405 24601
rect 4509 24567 4543 24601
rect 4647 24567 4681 24601
rect 2715 24430 2749 24464
rect 2853 24430 2887 24464
rect 2991 24430 3025 24464
rect 3129 24430 3163 24464
rect 3267 24430 3301 24464
rect 3405 24430 3439 24464
rect 3543 24430 3577 24464
rect 3681 24430 3715 24464
rect 3819 24430 3853 24464
rect 3957 24430 3991 24464
rect 4095 24430 4129 24464
rect 4233 24430 4267 24464
rect 4371 24430 4405 24464
rect 4509 24430 4543 24464
rect 4647 24430 4681 24464
rect 2715 24293 2749 24327
rect 2853 24293 2887 24327
rect 2991 24293 3025 24327
rect 3129 24293 3163 24327
rect 3267 24293 3301 24327
rect 3405 24293 3439 24327
rect 3543 24293 3577 24327
rect 3681 24293 3715 24327
rect 3819 24293 3853 24327
rect 3957 24293 3991 24327
rect 4095 24293 4129 24327
rect 4233 24293 4267 24327
rect 4371 24293 4405 24327
rect 4509 24293 4543 24327
rect 4647 24293 4681 24327
rect 2715 24156 2749 24190
rect 2853 24156 2887 24190
rect 2991 24156 3025 24190
rect 3129 24156 3163 24190
rect 3267 24156 3301 24190
rect 3405 24156 3439 24190
rect 3543 24156 3577 24190
rect 3681 24156 3715 24190
rect 3819 24156 3853 24190
rect 3957 24156 3991 24190
rect 4095 24156 4129 24190
rect 4233 24156 4267 24190
rect 4371 24156 4405 24190
rect 4509 24156 4543 24190
rect 4647 24156 4681 24190
rect 2715 24019 2749 24053
rect 2853 24019 2887 24053
rect 2991 24019 3025 24053
rect 3129 24019 3163 24053
rect 3267 24019 3301 24053
rect 3405 24019 3439 24053
rect 3543 24019 3577 24053
rect 3681 24019 3715 24053
rect 3819 24019 3853 24053
rect 3957 24019 3991 24053
rect 4095 24019 4129 24053
rect 4233 24019 4267 24053
rect 4371 24019 4405 24053
rect 4509 24019 4543 24053
rect 4647 24019 4681 24053
rect 2715 23882 2749 23916
rect 2853 23882 2887 23916
rect 2991 23882 3025 23916
rect 3129 23882 3163 23916
rect 3267 23882 3301 23916
rect 3405 23882 3439 23916
rect 3543 23882 3577 23916
rect 3681 23882 3715 23916
rect 3819 23882 3853 23916
rect 3957 23882 3991 23916
rect 4095 23882 4129 23916
rect 4233 23882 4267 23916
rect 4371 23882 4405 23916
rect 4509 23882 4543 23916
rect 4647 23882 4681 23916
rect 2715 23745 2749 23779
rect 2853 23745 2887 23779
rect 2991 23745 3025 23779
rect 3129 23745 3163 23779
rect 3267 23745 3301 23779
rect 3405 23745 3439 23779
rect 3543 23745 3577 23779
rect 3681 23745 3715 23779
rect 3819 23745 3853 23779
rect 3957 23745 3991 23779
rect 4095 23745 4129 23779
rect 4233 23745 4267 23779
rect 4371 23745 4405 23779
rect 4509 23745 4543 23779
rect 4647 23745 4681 23779
rect 2715 23608 2749 23642
rect 2853 23608 2887 23642
rect 2991 23608 3025 23642
rect 3129 23608 3163 23642
rect 3267 23608 3301 23642
rect 3405 23608 3439 23642
rect 3543 23608 3577 23642
rect 3681 23608 3715 23642
rect 3819 23608 3853 23642
rect 3957 23608 3991 23642
rect 4095 23608 4129 23642
rect 4233 23608 4267 23642
rect 4371 23608 4405 23642
rect 4509 23608 4543 23642
rect 4647 23608 4681 23642
rect 2715 23471 2749 23505
rect 2853 23471 2887 23505
rect 2991 23471 3025 23505
rect 3129 23471 3163 23505
rect 3267 23471 3301 23505
rect 3405 23471 3439 23505
rect 3543 23471 3577 23505
rect 3681 23471 3715 23505
rect 3819 23471 3853 23505
rect 3957 23471 3991 23505
rect 4095 23471 4129 23505
rect 4233 23471 4267 23505
rect 4371 23471 4405 23505
rect 4509 23471 4543 23505
rect 4647 23471 4681 23505
rect 2715 23334 2749 23368
rect 2853 23334 2887 23368
rect 2991 23334 3025 23368
rect 3129 23334 3163 23368
rect 3267 23334 3301 23368
rect 3405 23334 3439 23368
rect 3543 23334 3577 23368
rect 3681 23334 3715 23368
rect 3819 23334 3853 23368
rect 3957 23334 3991 23368
rect 4095 23334 4129 23368
rect 4233 23334 4267 23368
rect 4371 23334 4405 23368
rect 4509 23334 4543 23368
rect 4647 23334 4681 23368
rect 2715 23197 2749 23231
rect 2853 23197 2887 23231
rect 2991 23197 3025 23231
rect 3129 23197 3163 23231
rect 3267 23197 3301 23231
rect 3405 23197 3439 23231
rect 3543 23197 3577 23231
rect 3681 23197 3715 23231
rect 3819 23197 3853 23231
rect 3957 23197 3991 23231
rect 4095 23197 4129 23231
rect 4233 23197 4267 23231
rect 4371 23197 4405 23231
rect 4509 23197 4543 23231
rect 4647 23197 4681 23231
rect 2715 23060 2749 23094
rect 2853 23060 2887 23094
rect 2991 23060 3025 23094
rect 3129 23060 3163 23094
rect 3267 23060 3301 23094
rect 3405 23060 3439 23094
rect 3543 23060 3577 23094
rect 3681 23060 3715 23094
rect 3819 23060 3853 23094
rect 3957 23060 3991 23094
rect 4095 23060 4129 23094
rect 4233 23060 4267 23094
rect 4371 23060 4405 23094
rect 4509 23060 4543 23094
rect 4647 23060 4681 23094
rect 2715 22923 2749 22957
rect 2853 22923 2887 22957
rect 2991 22923 3025 22957
rect 3129 22923 3163 22957
rect 3267 22923 3301 22957
rect 3405 22923 3439 22957
rect 3543 22923 3577 22957
rect 3681 22923 3715 22957
rect 3819 22923 3853 22957
rect 3957 22923 3991 22957
rect 4095 22923 4129 22957
rect 4233 22923 4267 22957
rect 4371 22923 4405 22957
rect 4509 22923 4543 22957
rect 4647 22923 4681 22957
rect 2715 22786 2749 22820
rect 2853 22786 2887 22820
rect 2991 22786 3025 22820
rect 3129 22786 3163 22820
rect 3267 22786 3301 22820
rect 3405 22786 3439 22820
rect 3543 22786 3577 22820
rect 3681 22786 3715 22820
rect 3819 22786 3853 22820
rect 3957 22786 3991 22820
rect 4095 22786 4129 22820
rect 4233 22786 4267 22820
rect 4371 22786 4405 22820
rect 4509 22786 4543 22820
rect 4647 22786 4681 22820
rect 2715 22649 2749 22683
rect 2853 22649 2887 22683
rect 2991 22649 3025 22683
rect 3129 22649 3163 22683
rect 3267 22649 3301 22683
rect 3405 22649 3439 22683
rect 3543 22649 3577 22683
rect 3681 22649 3715 22683
rect 3819 22649 3853 22683
rect 3957 22649 3991 22683
rect 4095 22649 4129 22683
rect 4233 22649 4267 22683
rect 4371 22649 4405 22683
rect 4509 22649 4543 22683
rect 4647 22649 4681 22683
rect 2715 22512 2749 22546
rect 2853 22512 2887 22546
rect 2991 22512 3025 22546
rect 3129 22512 3163 22546
rect 3267 22512 3301 22546
rect 3405 22512 3439 22546
rect 3543 22512 3577 22546
rect 3681 22512 3715 22546
rect 3819 22512 3853 22546
rect 3957 22512 3991 22546
rect 4095 22512 4129 22546
rect 4233 22512 4267 22546
rect 4371 22512 4405 22546
rect 4509 22512 4543 22546
rect 4647 22512 4681 22546
rect 2715 22375 2749 22409
rect 2853 22375 2887 22409
rect 2991 22375 3025 22409
rect 3129 22375 3163 22409
rect 3267 22375 3301 22409
rect 3405 22375 3439 22409
rect 3543 22375 3577 22409
rect 3681 22375 3715 22409
rect 3819 22375 3853 22409
rect 3957 22375 3991 22409
rect 4095 22375 4129 22409
rect 4233 22375 4267 22409
rect 4371 22375 4405 22409
rect 4509 22375 4543 22409
rect 4647 22375 4681 22409
rect 2715 22238 2749 22272
rect 2853 22238 2887 22272
rect 2991 22238 3025 22272
rect 3129 22238 3163 22272
rect 3267 22238 3301 22272
rect 3405 22238 3439 22272
rect 3543 22238 3577 22272
rect 3681 22238 3715 22272
rect 3819 22238 3853 22272
rect 3957 22238 3991 22272
rect 4095 22238 4129 22272
rect 4233 22238 4267 22272
rect 4371 22238 4405 22272
rect 4509 22238 4543 22272
rect 4647 22238 4681 22272
rect 2715 22101 2749 22135
rect 2853 22101 2887 22135
rect 2991 22101 3025 22135
rect 3129 22101 3163 22135
rect 3267 22101 3301 22135
rect 3405 22101 3439 22135
rect 3543 22101 3577 22135
rect 3681 22101 3715 22135
rect 3819 22101 3853 22135
rect 3957 22101 3991 22135
rect 4095 22101 4129 22135
rect 4233 22101 4267 22135
rect 4371 22101 4405 22135
rect 4509 22101 4543 22135
rect 4647 22101 4681 22135
rect 2715 21964 2749 21998
rect 2853 21964 2887 21998
rect 2991 21964 3025 21998
rect 3129 21964 3163 21998
rect 3267 21964 3301 21998
rect 3405 21964 3439 21998
rect 3543 21964 3577 21998
rect 3681 21964 3715 21998
rect 3819 21964 3853 21998
rect 3957 21964 3991 21998
rect 4095 21964 4129 21998
rect 4233 21964 4267 21998
rect 4371 21964 4405 21998
rect 4509 21964 4543 21998
rect 4647 21964 4681 21998
rect 2715 21827 2749 21861
rect 2853 21827 2887 21861
rect 2991 21827 3025 21861
rect 3129 21827 3163 21861
rect 3267 21827 3301 21861
rect 3405 21827 3439 21861
rect 3543 21827 3577 21861
rect 3681 21827 3715 21861
rect 3819 21827 3853 21861
rect 3957 21827 3991 21861
rect 4095 21827 4129 21861
rect 4233 21827 4267 21861
rect 4371 21827 4405 21861
rect 4509 21827 4543 21861
rect 4647 21827 4681 21861
rect 2715 21690 2749 21724
rect 2853 21690 2887 21724
rect 2991 21690 3025 21724
rect 3129 21690 3163 21724
rect 3267 21690 3301 21724
rect 3405 21690 3439 21724
rect 3543 21690 3577 21724
rect 3681 21690 3715 21724
rect 3819 21690 3853 21724
rect 3957 21690 3991 21724
rect 4095 21690 4129 21724
rect 4233 21690 4267 21724
rect 4371 21690 4405 21724
rect 4509 21690 4543 21724
rect 4647 21690 4681 21724
rect 2715 21553 2749 21587
rect 2853 21553 2887 21587
rect 2991 21553 3025 21587
rect 3129 21553 3163 21587
rect 3267 21553 3301 21587
rect 3405 21553 3439 21587
rect 3543 21553 3577 21587
rect 3681 21553 3715 21587
rect 3819 21553 3853 21587
rect 3957 21553 3991 21587
rect 4095 21553 4129 21587
rect 4233 21553 4267 21587
rect 4371 21553 4405 21587
rect 4509 21553 4543 21587
rect 4647 21553 4681 21587
rect 2715 21416 2749 21450
rect 2853 21416 2887 21450
rect 2991 21416 3025 21450
rect 3129 21416 3163 21450
rect 3267 21416 3301 21450
rect 3405 21416 3439 21450
rect 3543 21416 3577 21450
rect 3681 21416 3715 21450
rect 3819 21416 3853 21450
rect 3957 21416 3991 21450
rect 4095 21416 4129 21450
rect 4233 21416 4267 21450
rect 4371 21416 4405 21450
rect 4509 21416 4543 21450
rect 4647 21416 4681 21450
rect 2715 21279 2749 21313
rect 2853 21279 2887 21313
rect 2991 21279 3025 21313
rect 3129 21279 3163 21313
rect 3267 21279 3301 21313
rect 3405 21279 3439 21313
rect 3543 21279 3577 21313
rect 3681 21279 3715 21313
rect 3819 21279 3853 21313
rect 3957 21279 3991 21313
rect 4095 21279 4129 21313
rect 4233 21279 4267 21313
rect 4371 21279 4405 21313
rect 4509 21279 4543 21313
rect 4647 21279 4681 21313
rect 2715 21142 2749 21176
rect 2853 21142 2887 21176
rect 2991 21142 3025 21176
rect 3129 21142 3163 21176
rect 3267 21142 3301 21176
rect 3405 21142 3439 21176
rect 3543 21142 3577 21176
rect 3681 21142 3715 21176
rect 3819 21142 3853 21176
rect 3957 21142 3991 21176
rect 4095 21142 4129 21176
rect 4233 21142 4267 21176
rect 4371 21142 4405 21176
rect 4509 21142 4543 21176
rect 4647 21142 4681 21176
rect 2715 21005 2749 21039
rect 2853 21005 2887 21039
rect 2991 21005 3025 21039
rect 3129 21005 3163 21039
rect 3267 21005 3301 21039
rect 3405 21005 3439 21039
rect 3543 21005 3577 21039
rect 3681 21005 3715 21039
rect 3819 21005 3853 21039
rect 3957 21005 3991 21039
rect 4095 21005 4129 21039
rect 4233 21005 4267 21039
rect 4371 21005 4405 21039
rect 4509 21005 4543 21039
rect 4647 21005 4681 21039
rect 2715 20868 2749 20902
rect 2853 20868 2887 20902
rect 2991 20868 3025 20902
rect 3129 20868 3163 20902
rect 3267 20868 3301 20902
rect 3405 20868 3439 20902
rect 3543 20868 3577 20902
rect 3681 20868 3715 20902
rect 3819 20868 3853 20902
rect 3957 20868 3991 20902
rect 4095 20868 4129 20902
rect 4233 20868 4267 20902
rect 4371 20868 4405 20902
rect 4509 20868 4543 20902
rect 4647 20868 4681 20902
rect 2715 20731 2749 20765
rect 2853 20731 2887 20765
rect 2991 20731 3025 20765
rect 3129 20731 3163 20765
rect 3267 20731 3301 20765
rect 3405 20731 3439 20765
rect 3543 20731 3577 20765
rect 3681 20731 3715 20765
rect 3819 20731 3853 20765
rect 3957 20731 3991 20765
rect 4095 20731 4129 20765
rect 4233 20731 4267 20765
rect 4371 20731 4405 20765
rect 4509 20731 4543 20765
rect 4647 20731 4681 20765
rect 2715 20594 2749 20628
rect 2853 20594 2887 20628
rect 2991 20594 3025 20628
rect 3129 20594 3163 20628
rect 3267 20594 3301 20628
rect 3405 20594 3439 20628
rect 3543 20594 3577 20628
rect 3681 20594 3715 20628
rect 3819 20594 3853 20628
rect 3957 20594 3991 20628
rect 4095 20594 4129 20628
rect 4233 20594 4267 20628
rect 4371 20594 4405 20628
rect 4509 20594 4543 20628
rect 4647 20594 4681 20628
rect 2715 20457 2749 20491
rect 2853 20457 2887 20491
rect 2991 20457 3025 20491
rect 3129 20457 3163 20491
rect 3267 20457 3301 20491
rect 3405 20457 3439 20491
rect 3543 20457 3577 20491
rect 3681 20457 3715 20491
rect 3819 20457 3853 20491
rect 3957 20457 3991 20491
rect 4095 20457 4129 20491
rect 4233 20457 4267 20491
rect 4371 20457 4405 20491
rect 4509 20457 4543 20491
rect 4647 20457 4681 20491
rect 2715 20320 2749 20354
rect 2853 20320 2887 20354
rect 2991 20320 3025 20354
rect 3129 20320 3163 20354
rect 3267 20320 3301 20354
rect 3405 20320 3439 20354
rect 3543 20320 3577 20354
rect 3681 20320 3715 20354
rect 3819 20320 3853 20354
rect 3957 20320 3991 20354
rect 4095 20320 4129 20354
rect 4233 20320 4267 20354
rect 4371 20320 4405 20354
rect 4509 20320 4543 20354
rect 4647 20320 4681 20354
rect 2715 20183 2749 20217
rect 2853 20183 2887 20217
rect 2991 20183 3025 20217
rect 3129 20183 3163 20217
rect 3267 20183 3301 20217
rect 3405 20183 3439 20217
rect 3543 20183 3577 20217
rect 3681 20183 3715 20217
rect 3819 20183 3853 20217
rect 3957 20183 3991 20217
rect 4095 20183 4129 20217
rect 4233 20183 4267 20217
rect 4371 20183 4405 20217
rect 4509 20183 4543 20217
rect 4647 20183 4681 20217
rect 2715 20046 2749 20080
rect 2853 20046 2887 20080
rect 2991 20046 3025 20080
rect 3129 20046 3163 20080
rect 3267 20046 3301 20080
rect 3405 20046 3439 20080
rect 3543 20046 3577 20080
rect 3681 20046 3715 20080
rect 3819 20046 3853 20080
rect 3957 20046 3991 20080
rect 4095 20046 4129 20080
rect 4233 20046 4267 20080
rect 4371 20046 4405 20080
rect 4509 20046 4543 20080
rect 4647 20046 4681 20080
rect 2715 19909 2749 19943
rect 2853 19909 2887 19943
rect 2991 19909 3025 19943
rect 3129 19909 3163 19943
rect 3267 19909 3301 19943
rect 3405 19909 3439 19943
rect 3543 19909 3577 19943
rect 3681 19909 3715 19943
rect 3819 19909 3853 19943
rect 3957 19909 3991 19943
rect 4095 19909 4129 19943
rect 4233 19909 4267 19943
rect 4371 19909 4405 19943
rect 4509 19909 4543 19943
rect 4647 19909 4681 19943
rect 2715 19772 2749 19806
rect 2853 19772 2887 19806
rect 2991 19772 3025 19806
rect 3129 19772 3163 19806
rect 3267 19772 3301 19806
rect 3405 19772 3439 19806
rect 3543 19772 3577 19806
rect 3681 19772 3715 19806
rect 3819 19772 3853 19806
rect 3957 19772 3991 19806
rect 4095 19772 4129 19806
rect 4233 19772 4267 19806
rect 4371 19772 4405 19806
rect 4509 19772 4543 19806
rect 4647 19772 4681 19806
rect 2715 19635 2749 19669
rect 2853 19635 2887 19669
rect 2991 19635 3025 19669
rect 3129 19635 3163 19669
rect 3267 19635 3301 19669
rect 3405 19635 3439 19669
rect 3543 19635 3577 19669
rect 3681 19635 3715 19669
rect 3819 19635 3853 19669
rect 3957 19635 3991 19669
rect 4095 19635 4129 19669
rect 4233 19635 4267 19669
rect 4371 19635 4405 19669
rect 4509 19635 4543 19669
rect 4647 19635 4681 19669
rect 2715 19498 2749 19532
rect 2853 19498 2887 19532
rect 2991 19498 3025 19532
rect 3129 19498 3163 19532
rect 3267 19498 3301 19532
rect 3405 19498 3439 19532
rect 3543 19498 3577 19532
rect 3681 19498 3715 19532
rect 3819 19498 3853 19532
rect 3957 19498 3991 19532
rect 4095 19498 4129 19532
rect 4233 19498 4267 19532
rect 4371 19498 4405 19532
rect 4509 19498 4543 19532
rect 4647 19498 4681 19532
rect 2715 19361 2749 19395
rect 2853 19361 2887 19395
rect 2991 19361 3025 19395
rect 3129 19361 3163 19395
rect 3267 19361 3301 19395
rect 3405 19361 3439 19395
rect 3543 19361 3577 19395
rect 3681 19361 3715 19395
rect 3819 19361 3853 19395
rect 3957 19361 3991 19395
rect 4095 19361 4129 19395
rect 4233 19361 4267 19395
rect 4371 19361 4405 19395
rect 4509 19361 4543 19395
rect 4647 19361 4681 19395
rect 2715 19224 2749 19258
rect 2853 19224 2887 19258
rect 2991 19224 3025 19258
rect 3129 19224 3163 19258
rect 3267 19224 3301 19258
rect 3405 19224 3439 19258
rect 3543 19224 3577 19258
rect 3681 19224 3715 19258
rect 3819 19224 3853 19258
rect 3957 19224 3991 19258
rect 4095 19224 4129 19258
rect 4233 19224 4267 19258
rect 4371 19224 4405 19258
rect 4509 19224 4543 19258
rect 4647 19224 4681 19258
rect 2715 19087 2749 19121
rect 2853 19087 2887 19121
rect 2991 19087 3025 19121
rect 3129 19087 3163 19121
rect 3267 19087 3301 19121
rect 3405 19087 3439 19121
rect 3543 19087 3577 19121
rect 3681 19087 3715 19121
rect 3819 19087 3853 19121
rect 3957 19087 3991 19121
rect 4095 19087 4129 19121
rect 4233 19087 4267 19121
rect 4371 19087 4405 19121
rect 4509 19087 4543 19121
rect 4647 19087 4681 19121
rect 2715 18950 2749 18984
rect 2853 18950 2887 18984
rect 2991 18950 3025 18984
rect 3129 18950 3163 18984
rect 3267 18950 3301 18984
rect 3405 18950 3439 18984
rect 3543 18950 3577 18984
rect 3681 18950 3715 18984
rect 3819 18950 3853 18984
rect 3957 18950 3991 18984
rect 4095 18950 4129 18984
rect 4233 18950 4267 18984
rect 4371 18950 4405 18984
rect 4509 18950 4543 18984
rect 4647 18950 4681 18984
rect 2715 18813 2749 18847
rect 2853 18813 2887 18847
rect 2991 18813 3025 18847
rect 3129 18813 3163 18847
rect 3267 18813 3301 18847
rect 3405 18813 3439 18847
rect 3543 18813 3577 18847
rect 3681 18813 3715 18847
rect 3819 18813 3853 18847
rect 3957 18813 3991 18847
rect 4095 18813 4129 18847
rect 4233 18813 4267 18847
rect 4371 18813 4405 18847
rect 4509 18813 4543 18847
rect 4647 18813 4681 18847
rect 2715 18676 2749 18710
rect 2853 18676 2887 18710
rect 2991 18676 3025 18710
rect 3129 18676 3163 18710
rect 3267 18676 3301 18710
rect 3405 18676 3439 18710
rect 3543 18676 3577 18710
rect 3681 18676 3715 18710
rect 3819 18676 3853 18710
rect 3957 18676 3991 18710
rect 4095 18676 4129 18710
rect 4233 18676 4267 18710
rect 4371 18676 4405 18710
rect 4509 18676 4543 18710
rect 4647 18676 4681 18710
rect 2715 18539 2749 18573
rect 2853 18539 2887 18573
rect 2991 18539 3025 18573
rect 3129 18539 3163 18573
rect 3267 18539 3301 18573
rect 3405 18539 3439 18573
rect 3543 18539 3577 18573
rect 3681 18539 3715 18573
rect 3819 18539 3853 18573
rect 3957 18539 3991 18573
rect 4095 18539 4129 18573
rect 4233 18539 4267 18573
rect 4371 18539 4405 18573
rect 4509 18539 4543 18573
rect 4647 18539 4681 18573
rect 2715 18402 2749 18436
rect 2853 18402 2887 18436
rect 2991 18402 3025 18436
rect 3129 18402 3163 18436
rect 3267 18402 3301 18436
rect 3405 18402 3439 18436
rect 3543 18402 3577 18436
rect 3681 18402 3715 18436
rect 3819 18402 3853 18436
rect 3957 18402 3991 18436
rect 4095 18402 4129 18436
rect 4233 18402 4267 18436
rect 4371 18402 4405 18436
rect 4509 18402 4543 18436
rect 4647 18402 4681 18436
rect 2715 18265 2749 18299
rect 2853 18265 2887 18299
rect 2991 18265 3025 18299
rect 3129 18265 3163 18299
rect 3267 18265 3301 18299
rect 3405 18265 3439 18299
rect 3543 18265 3577 18299
rect 3681 18265 3715 18299
rect 3819 18265 3853 18299
rect 3957 18265 3991 18299
rect 4095 18265 4129 18299
rect 4233 18265 4267 18299
rect 4371 18265 4405 18299
rect 4509 18265 4543 18299
rect 4647 18265 4681 18299
rect 2715 18128 2749 18162
rect 2853 18128 2887 18162
rect 2991 18128 3025 18162
rect 3129 18128 3163 18162
rect 3267 18128 3301 18162
rect 3405 18128 3439 18162
rect 3543 18128 3577 18162
rect 3681 18128 3715 18162
rect 3819 18128 3853 18162
rect 3957 18128 3991 18162
rect 4095 18128 4129 18162
rect 4233 18128 4267 18162
rect 4371 18128 4405 18162
rect 4509 18128 4543 18162
rect 4647 18128 4681 18162
rect 2715 17991 2749 18025
rect 2853 17991 2887 18025
rect 2991 17991 3025 18025
rect 3129 17991 3163 18025
rect 3267 17991 3301 18025
rect 3405 17991 3439 18025
rect 3543 17991 3577 18025
rect 3681 17991 3715 18025
rect 3819 17991 3853 18025
rect 3957 17991 3991 18025
rect 4095 17991 4129 18025
rect 4233 17991 4267 18025
rect 4371 17991 4405 18025
rect 4509 17991 4543 18025
rect 4647 17991 4681 18025
rect 2715 17854 2749 17888
rect 2853 17854 2887 17888
rect 2991 17854 3025 17888
rect 3129 17854 3163 17888
rect 3267 17854 3301 17888
rect 3405 17854 3439 17888
rect 3543 17854 3577 17888
rect 3681 17854 3715 17888
rect 3819 17854 3853 17888
rect 3957 17854 3991 17888
rect 4095 17854 4129 17888
rect 4233 17854 4267 17888
rect 4371 17854 4405 17888
rect 4509 17854 4543 17888
rect 4647 17854 4681 17888
rect 2715 17717 2749 17751
rect 2853 17717 2887 17751
rect 2991 17717 3025 17751
rect 3129 17717 3163 17751
rect 3267 17717 3301 17751
rect 3405 17717 3439 17751
rect 3543 17717 3577 17751
rect 3681 17717 3715 17751
rect 3819 17717 3853 17751
rect 3957 17717 3991 17751
rect 4095 17717 4129 17751
rect 4233 17717 4267 17751
rect 4371 17717 4405 17751
rect 4509 17717 4543 17751
rect 4647 17717 4681 17751
rect 2715 17580 2749 17614
rect 2853 17580 2887 17614
rect 2991 17580 3025 17614
rect 3129 17580 3163 17614
rect 3267 17580 3301 17614
rect 3405 17580 3439 17614
rect 3543 17580 3577 17614
rect 3681 17580 3715 17614
rect 3819 17580 3853 17614
rect 3957 17580 3991 17614
rect 4095 17580 4129 17614
rect 4233 17580 4267 17614
rect 4371 17580 4405 17614
rect 4509 17580 4543 17614
rect 4647 17580 4681 17614
rect 2715 17443 2749 17477
rect 2853 17443 2887 17477
rect 2991 17443 3025 17477
rect 3129 17443 3163 17477
rect 3267 17443 3301 17477
rect 3405 17443 3439 17477
rect 3543 17443 3577 17477
rect 3681 17443 3715 17477
rect 3819 17443 3853 17477
rect 3957 17443 3991 17477
rect 4095 17443 4129 17477
rect 4233 17443 4267 17477
rect 4371 17443 4405 17477
rect 4509 17443 4543 17477
rect 4647 17443 4681 17477
rect 2715 17306 2749 17340
rect 2853 17306 2887 17340
rect 2991 17306 3025 17340
rect 3129 17306 3163 17340
rect 3267 17306 3301 17340
rect 3405 17306 3439 17340
rect 3543 17306 3577 17340
rect 3681 17306 3715 17340
rect 3819 17306 3853 17340
rect 3957 17306 3991 17340
rect 4095 17306 4129 17340
rect 4233 17306 4267 17340
rect 4371 17306 4405 17340
rect 4509 17306 4543 17340
rect 4647 17306 4681 17340
rect 2715 17169 2749 17203
rect 2853 17169 2887 17203
rect 2991 17169 3025 17203
rect 3129 17169 3163 17203
rect 3267 17169 3301 17203
rect 3405 17169 3439 17203
rect 3543 17169 3577 17203
rect 3681 17169 3715 17203
rect 3819 17169 3853 17203
rect 3957 17169 3991 17203
rect 4095 17169 4129 17203
rect 4233 17169 4267 17203
rect 4371 17169 4405 17203
rect 4509 17169 4543 17203
rect 4647 17169 4681 17203
rect 2715 17032 2749 17066
rect 2853 17032 2887 17066
rect 2991 17032 3025 17066
rect 3129 17032 3163 17066
rect 3267 17032 3301 17066
rect 3405 17032 3439 17066
rect 3543 17032 3577 17066
rect 3681 17032 3715 17066
rect 3819 17032 3853 17066
rect 3957 17032 3991 17066
rect 4095 17032 4129 17066
rect 4233 17032 4267 17066
rect 4371 17032 4405 17066
rect 4509 17032 4543 17066
rect 4647 17032 4681 17066
rect 4740 17000 4774 17034
rect 4809 17000 4843 17034
rect 4878 17000 4912 17034
rect 4947 17000 4981 17034
rect 5016 17000 5050 17034
rect 5085 17000 5119 17034
rect 5154 17000 5188 17034
rect 5223 17000 5257 17034
rect 5292 17000 5326 17034
rect 5361 17000 5395 17034
rect 5430 17000 5464 17034
rect 5499 17000 5533 17034
rect 5568 17000 5602 17034
rect 5637 17000 5671 17034
rect 5706 17000 5740 17034
rect 5775 17000 5809 17034
rect 5844 17000 5878 17034
rect 5913 17000 5947 17034
rect 5982 17000 6016 17034
rect 6051 17000 6085 17034
rect 6120 17000 6154 17034
rect 6189 17000 6223 17034
rect 6258 17000 6292 17034
rect 6327 17000 6361 17034
rect 6396 17000 6430 17034
rect 6465 17000 6499 17034
rect 6534 17000 6568 17034
rect 6603 17000 6637 17034
rect 6672 17000 6706 17034
rect 6741 17000 6775 17034
rect 6810 17000 6844 17034
rect 6879 17000 6913 17034
rect 6948 17000 6982 17034
rect 7017 17000 7051 17034
rect 7086 17000 7120 17034
rect 7155 17000 7189 17034
rect 7224 17000 7258 17034
rect 7293 17000 7327 17034
rect 7362 17000 7396 17034
rect 7431 17000 7465 17034
rect 7500 17000 7534 17034
rect 7568 17000 7602 17034
rect 7636 17000 7670 17034
rect 7704 17000 7738 17034
rect 7772 17000 7806 17034
rect 7840 17000 7874 17034
rect 4740 16930 4774 16964
rect 4809 16930 4843 16964
rect 4878 16930 4912 16964
rect 4947 16930 4981 16964
rect 5016 16930 5050 16964
rect 5085 16930 5119 16964
rect 5154 16930 5188 16964
rect 5223 16930 5257 16964
rect 5292 16930 5326 16964
rect 5361 16930 5395 16964
rect 5430 16930 5464 16964
rect 5499 16930 5533 16964
rect 5568 16930 5602 16964
rect 5637 16930 5671 16964
rect 5706 16930 5740 16964
rect 5775 16930 5809 16964
rect 5844 16930 5878 16964
rect 5913 16930 5947 16964
rect 5982 16930 6016 16964
rect 6051 16930 6085 16964
rect 6120 16930 6154 16964
rect 6189 16930 6223 16964
rect 6258 16930 6292 16964
rect 6327 16930 6361 16964
rect 6396 16930 6430 16964
rect 6465 16930 6499 16964
rect 6534 16930 6568 16964
rect 6603 16930 6637 16964
rect 6672 16930 6706 16964
rect 6741 16930 6775 16964
rect 6810 16930 6844 16964
rect 6879 16930 6913 16964
rect 6948 16930 6982 16964
rect 7017 16930 7051 16964
rect 7086 16930 7120 16964
rect 7155 16930 7189 16964
rect 7224 16930 7258 16964
rect 7293 16930 7327 16964
rect 7362 16930 7396 16964
rect 7431 16930 7465 16964
rect 7500 16930 7534 16964
rect 7568 16930 7602 16964
rect 7636 16930 7670 16964
rect 7704 16930 7738 16964
rect 7772 16930 7806 16964
rect 7840 16930 7874 16964
rect 2715 16895 2749 16929
rect 2853 16895 2887 16929
rect 2991 16895 3025 16929
rect 3129 16895 3163 16929
rect 3267 16895 3301 16929
rect 3405 16895 3439 16929
rect 3543 16895 3577 16929
rect 3681 16895 3715 16929
rect 3819 16895 3853 16929
rect 3957 16895 3991 16929
rect 4095 16895 4129 16929
rect 4233 16895 4267 16929
rect 4371 16895 4405 16929
rect 4509 16895 4543 16929
rect 4647 16895 4681 16929
rect 4740 16860 4774 16894
rect 4809 16860 4843 16894
rect 4878 16860 4912 16894
rect 4947 16860 4981 16894
rect 5016 16860 5050 16894
rect 5085 16860 5119 16894
rect 5154 16860 5188 16894
rect 5223 16860 5257 16894
rect 5292 16860 5326 16894
rect 5361 16860 5395 16894
rect 5430 16860 5464 16894
rect 5499 16860 5533 16894
rect 5568 16860 5602 16894
rect 5637 16860 5671 16894
rect 5706 16860 5740 16894
rect 5775 16860 5809 16894
rect 5844 16860 5878 16894
rect 5913 16860 5947 16894
rect 5982 16860 6016 16894
rect 6051 16860 6085 16894
rect 6120 16860 6154 16894
rect 6189 16860 6223 16894
rect 6258 16860 6292 16894
rect 6327 16860 6361 16894
rect 6396 16860 6430 16894
rect 6465 16860 6499 16894
rect 6534 16860 6568 16894
rect 6603 16860 6637 16894
rect 6672 16860 6706 16894
rect 6741 16860 6775 16894
rect 6810 16860 6844 16894
rect 6879 16860 6913 16894
rect 6948 16860 6982 16894
rect 7017 16860 7051 16894
rect 7086 16860 7120 16894
rect 7155 16860 7189 16894
rect 7224 16860 7258 16894
rect 7293 16860 7327 16894
rect 7362 16860 7396 16894
rect 7431 16860 7465 16894
rect 7500 16860 7534 16894
rect 7568 16860 7602 16894
rect 7636 16860 7670 16894
rect 7704 16860 7738 16894
rect 7772 16860 7806 16894
rect 7840 16860 7874 16894
rect 2715 16758 2749 16792
rect 2853 16758 2887 16792
rect 2991 16758 3025 16792
rect 3129 16758 3163 16792
rect 3267 16758 3301 16792
rect 3405 16758 3439 16792
rect 3543 16758 3577 16792
rect 3681 16758 3715 16792
rect 3819 16758 3853 16792
rect 3957 16758 3991 16792
rect 4095 16758 4129 16792
rect 4233 16758 4267 16792
rect 4371 16758 4405 16792
rect 4509 16758 4543 16792
rect 4647 16758 4681 16792
rect 4740 16790 4774 16824
rect 4809 16790 4843 16824
rect 4878 16790 4912 16824
rect 4947 16790 4981 16824
rect 5016 16790 5050 16824
rect 5085 16790 5119 16824
rect 5154 16790 5188 16824
rect 5223 16790 5257 16824
rect 5292 16790 5326 16824
rect 5361 16790 5395 16824
rect 5430 16790 5464 16824
rect 5499 16790 5533 16824
rect 5568 16790 5602 16824
rect 5637 16790 5671 16824
rect 5706 16790 5740 16824
rect 5775 16790 5809 16824
rect 5844 16790 5878 16824
rect 5913 16790 5947 16824
rect 5982 16790 6016 16824
rect 6051 16790 6085 16824
rect 6120 16790 6154 16824
rect 6189 16790 6223 16824
rect 6258 16790 6292 16824
rect 6327 16790 6361 16824
rect 6396 16790 6430 16824
rect 6465 16790 6499 16824
rect 6534 16790 6568 16824
rect 6603 16790 6637 16824
rect 6672 16790 6706 16824
rect 6741 16790 6775 16824
rect 6810 16790 6844 16824
rect 6879 16790 6913 16824
rect 6948 16790 6982 16824
rect 7017 16790 7051 16824
rect 7086 16790 7120 16824
rect 7155 16790 7189 16824
rect 7224 16790 7258 16824
rect 7293 16790 7327 16824
rect 7362 16790 7396 16824
rect 7431 16790 7465 16824
rect 7500 16790 7534 16824
rect 7568 16790 7602 16824
rect 7636 16790 7670 16824
rect 7704 16790 7738 16824
rect 7772 16790 7806 16824
rect 7840 16790 7874 16824
rect 4740 16720 4774 16754
rect 4809 16720 4843 16754
rect 4878 16720 4912 16754
rect 4947 16720 4981 16754
rect 5016 16720 5050 16754
rect 5085 16720 5119 16754
rect 5154 16720 5188 16754
rect 5223 16720 5257 16754
rect 5292 16720 5326 16754
rect 5361 16720 5395 16754
rect 5430 16720 5464 16754
rect 5499 16720 5533 16754
rect 5568 16720 5602 16754
rect 5637 16720 5671 16754
rect 5706 16720 5740 16754
rect 5775 16720 5809 16754
rect 5844 16720 5878 16754
rect 5913 16720 5947 16754
rect 5982 16720 6016 16754
rect 6051 16720 6085 16754
rect 6120 16720 6154 16754
rect 6189 16720 6223 16754
rect 6258 16720 6292 16754
rect 6327 16720 6361 16754
rect 6396 16720 6430 16754
rect 6465 16720 6499 16754
rect 6534 16720 6568 16754
rect 6603 16720 6637 16754
rect 6672 16720 6706 16754
rect 6741 16720 6775 16754
rect 6810 16720 6844 16754
rect 6879 16720 6913 16754
rect 6948 16720 6982 16754
rect 7017 16720 7051 16754
rect 7086 16720 7120 16754
rect 7155 16720 7189 16754
rect 7224 16720 7258 16754
rect 7293 16720 7327 16754
rect 7362 16720 7396 16754
rect 7431 16720 7465 16754
rect 7500 16720 7534 16754
rect 7568 16720 7602 16754
rect 7636 16720 7670 16754
rect 7704 16720 7738 16754
rect 7772 16720 7806 16754
rect 7840 16720 7874 16754
rect 2715 16621 2749 16655
rect 2853 16621 2887 16655
rect 2991 16621 3025 16655
rect 3129 16621 3163 16655
rect 3267 16621 3301 16655
rect 3405 16621 3439 16655
rect 3543 16621 3577 16655
rect 3681 16621 3715 16655
rect 3819 16621 3853 16655
rect 3957 16621 3991 16655
rect 4095 16621 4129 16655
rect 4233 16621 4267 16655
rect 4371 16621 4405 16655
rect 4509 16621 4543 16655
rect 4647 16621 4681 16655
rect 4740 16650 4774 16684
rect 4809 16650 4843 16684
rect 4878 16650 4912 16684
rect 4947 16650 4981 16684
rect 5016 16650 5050 16684
rect 5085 16650 5119 16684
rect 5154 16650 5188 16684
rect 5223 16650 5257 16684
rect 5292 16650 5326 16684
rect 5361 16650 5395 16684
rect 5430 16650 5464 16684
rect 5499 16650 5533 16684
rect 5568 16650 5602 16684
rect 5637 16650 5671 16684
rect 5706 16650 5740 16684
rect 5775 16650 5809 16684
rect 5844 16650 5878 16684
rect 5913 16650 5947 16684
rect 5982 16650 6016 16684
rect 6051 16650 6085 16684
rect 6120 16650 6154 16684
rect 6189 16650 6223 16684
rect 6258 16650 6292 16684
rect 6327 16650 6361 16684
rect 6396 16650 6430 16684
rect 6465 16650 6499 16684
rect 6534 16650 6568 16684
rect 6603 16650 6637 16684
rect 6672 16650 6706 16684
rect 6741 16650 6775 16684
rect 6810 16650 6844 16684
rect 6879 16650 6913 16684
rect 6948 16650 6982 16684
rect 7017 16650 7051 16684
rect 7086 16650 7120 16684
rect 7155 16650 7189 16684
rect 7224 16650 7258 16684
rect 7293 16650 7327 16684
rect 7362 16650 7396 16684
rect 7431 16650 7465 16684
rect 7500 16650 7534 16684
rect 7568 16650 7602 16684
rect 7636 16650 7670 16684
rect 7704 16650 7738 16684
rect 7772 16650 7806 16684
rect 7840 16650 7874 16684
rect 4740 16580 4774 16614
rect 4809 16580 4843 16614
rect 4878 16580 4912 16614
rect 4947 16580 4981 16614
rect 5016 16580 5050 16614
rect 5085 16580 5119 16614
rect 5154 16580 5188 16614
rect 5223 16580 5257 16614
rect 5292 16580 5326 16614
rect 5361 16580 5395 16614
rect 5430 16580 5464 16614
rect 5499 16580 5533 16614
rect 5568 16580 5602 16614
rect 5637 16580 5671 16614
rect 5706 16580 5740 16614
rect 5775 16580 5809 16614
rect 5844 16580 5878 16614
rect 5913 16580 5947 16614
rect 5982 16580 6016 16614
rect 6051 16580 6085 16614
rect 6120 16580 6154 16614
rect 6189 16580 6223 16614
rect 6258 16580 6292 16614
rect 6327 16580 6361 16614
rect 6396 16580 6430 16614
rect 6465 16580 6499 16614
rect 6534 16580 6568 16614
rect 6603 16580 6637 16614
rect 6672 16580 6706 16614
rect 6741 16580 6775 16614
rect 6810 16580 6844 16614
rect 6879 16580 6913 16614
rect 6948 16580 6982 16614
rect 7017 16580 7051 16614
rect 7086 16580 7120 16614
rect 7155 16580 7189 16614
rect 7224 16580 7258 16614
rect 7293 16580 7327 16614
rect 7362 16580 7396 16614
rect 7431 16580 7465 16614
rect 7500 16580 7534 16614
rect 7568 16580 7602 16614
rect 7636 16580 7670 16614
rect 7704 16580 7738 16614
rect 7772 16580 7806 16614
rect 7840 16580 7874 16614
rect 2715 16484 2749 16518
rect 2853 16484 2887 16518
rect 2991 16484 3025 16518
rect 3129 16484 3163 16518
rect 3267 16484 3301 16518
rect 3405 16484 3439 16518
rect 3543 16484 3577 16518
rect 3681 16484 3715 16518
rect 3819 16484 3853 16518
rect 3957 16484 3991 16518
rect 4095 16484 4129 16518
rect 4233 16484 4267 16518
rect 4371 16484 4405 16518
rect 4509 16484 4543 16518
rect 4647 16484 4681 16518
rect 4740 16510 4774 16544
rect 4809 16510 4843 16544
rect 4878 16510 4912 16544
rect 4947 16510 4981 16544
rect 5016 16510 5050 16544
rect 5085 16510 5119 16544
rect 5154 16510 5188 16544
rect 5223 16510 5257 16544
rect 5292 16510 5326 16544
rect 5361 16510 5395 16544
rect 5430 16510 5464 16544
rect 5499 16510 5533 16544
rect 5568 16510 5602 16544
rect 5637 16510 5671 16544
rect 5706 16510 5740 16544
rect 5775 16510 5809 16544
rect 5844 16510 5878 16544
rect 5913 16510 5947 16544
rect 5982 16510 6016 16544
rect 6051 16510 6085 16544
rect 6120 16510 6154 16544
rect 6189 16510 6223 16544
rect 6258 16510 6292 16544
rect 6327 16510 6361 16544
rect 6396 16510 6430 16544
rect 6465 16510 6499 16544
rect 6534 16510 6568 16544
rect 6603 16510 6637 16544
rect 6672 16510 6706 16544
rect 6741 16510 6775 16544
rect 6810 16510 6844 16544
rect 6879 16510 6913 16544
rect 6948 16510 6982 16544
rect 7017 16510 7051 16544
rect 7086 16510 7120 16544
rect 7155 16510 7189 16544
rect 7224 16510 7258 16544
rect 7293 16510 7327 16544
rect 7362 16510 7396 16544
rect 7431 16510 7465 16544
rect 7500 16510 7534 16544
rect 7568 16510 7602 16544
rect 7636 16510 7670 16544
rect 7704 16510 7738 16544
rect 7772 16510 7806 16544
rect 7840 16510 7874 16544
rect 4740 16440 4774 16474
rect 4809 16440 4843 16474
rect 4878 16440 4912 16474
rect 4947 16440 4981 16474
rect 5016 16440 5050 16474
rect 5085 16440 5119 16474
rect 5154 16440 5188 16474
rect 5223 16440 5257 16474
rect 5292 16440 5326 16474
rect 5361 16440 5395 16474
rect 5430 16440 5464 16474
rect 5499 16440 5533 16474
rect 5568 16440 5602 16474
rect 5637 16440 5671 16474
rect 5706 16440 5740 16474
rect 5775 16440 5809 16474
rect 5844 16440 5878 16474
rect 5913 16440 5947 16474
rect 5982 16440 6016 16474
rect 6051 16440 6085 16474
rect 6120 16440 6154 16474
rect 6189 16440 6223 16474
rect 6258 16440 6292 16474
rect 6327 16440 6361 16474
rect 6396 16440 6430 16474
rect 6465 16440 6499 16474
rect 6534 16440 6568 16474
rect 6603 16440 6637 16474
rect 6672 16440 6706 16474
rect 6741 16440 6775 16474
rect 6810 16440 6844 16474
rect 6879 16440 6913 16474
rect 6948 16440 6982 16474
rect 7017 16440 7051 16474
rect 7086 16440 7120 16474
rect 7155 16440 7189 16474
rect 7224 16440 7258 16474
rect 7293 16440 7327 16474
rect 7362 16440 7396 16474
rect 7431 16440 7465 16474
rect 7500 16440 7534 16474
rect 7568 16440 7602 16474
rect 7636 16440 7670 16474
rect 7704 16440 7738 16474
rect 7772 16440 7806 16474
rect 7840 16440 7874 16474
rect 2715 16347 2749 16381
rect 2853 16347 2887 16381
rect 2991 16347 3025 16381
rect 3129 16347 3163 16381
rect 3267 16347 3301 16381
rect 3405 16347 3439 16381
rect 3543 16347 3577 16381
rect 3681 16347 3715 16381
rect 3819 16347 3853 16381
rect 3957 16347 3991 16381
rect 4095 16347 4129 16381
rect 4233 16347 4267 16381
rect 4371 16347 4405 16381
rect 4509 16347 4543 16381
rect 4647 16347 4681 16381
rect 4740 16370 4774 16404
rect 4809 16370 4843 16404
rect 4878 16370 4912 16404
rect 4947 16370 4981 16404
rect 5016 16370 5050 16404
rect 5085 16370 5119 16404
rect 5154 16370 5188 16404
rect 5223 16370 5257 16404
rect 5292 16370 5326 16404
rect 5361 16370 5395 16404
rect 5430 16370 5464 16404
rect 5499 16370 5533 16404
rect 5568 16370 5602 16404
rect 5637 16370 5671 16404
rect 5706 16370 5740 16404
rect 5775 16370 5809 16404
rect 5844 16370 5878 16404
rect 5913 16370 5947 16404
rect 5982 16370 6016 16404
rect 6051 16370 6085 16404
rect 6120 16370 6154 16404
rect 6189 16370 6223 16404
rect 6258 16370 6292 16404
rect 6327 16370 6361 16404
rect 6396 16370 6430 16404
rect 6465 16370 6499 16404
rect 6534 16370 6568 16404
rect 6603 16370 6637 16404
rect 6672 16370 6706 16404
rect 6741 16370 6775 16404
rect 6810 16370 6844 16404
rect 6879 16370 6913 16404
rect 6948 16370 6982 16404
rect 7017 16370 7051 16404
rect 7086 16370 7120 16404
rect 7155 16370 7189 16404
rect 7224 16370 7258 16404
rect 7293 16370 7327 16404
rect 7362 16370 7396 16404
rect 7431 16370 7465 16404
rect 7500 16370 7534 16404
rect 7568 16370 7602 16404
rect 7636 16370 7670 16404
rect 7704 16370 7738 16404
rect 7772 16370 7806 16404
rect 7840 16370 7874 16404
rect 4740 16300 4774 16334
rect 4809 16300 4843 16334
rect 4878 16300 4912 16334
rect 4947 16300 4981 16334
rect 5016 16300 5050 16334
rect 5085 16300 5119 16334
rect 5154 16300 5188 16334
rect 5223 16300 5257 16334
rect 5292 16300 5326 16334
rect 5361 16300 5395 16334
rect 5430 16300 5464 16334
rect 5499 16300 5533 16334
rect 5568 16300 5602 16334
rect 5637 16300 5671 16334
rect 5706 16300 5740 16334
rect 5775 16300 5809 16334
rect 5844 16300 5878 16334
rect 5913 16300 5947 16334
rect 5982 16300 6016 16334
rect 6051 16300 6085 16334
rect 6120 16300 6154 16334
rect 6189 16300 6223 16334
rect 6258 16300 6292 16334
rect 6327 16300 6361 16334
rect 6396 16300 6430 16334
rect 6465 16300 6499 16334
rect 6534 16300 6568 16334
rect 6603 16300 6637 16334
rect 6672 16300 6706 16334
rect 6741 16300 6775 16334
rect 6810 16300 6844 16334
rect 6879 16300 6913 16334
rect 6948 16300 6982 16334
rect 7017 16300 7051 16334
rect 7086 16300 7120 16334
rect 7155 16300 7189 16334
rect 7224 16300 7258 16334
rect 7293 16300 7327 16334
rect 7362 16300 7396 16334
rect 7431 16300 7465 16334
rect 7500 16300 7534 16334
rect 7568 16300 7602 16334
rect 7636 16300 7670 16334
rect 7704 16300 7738 16334
rect 7772 16300 7806 16334
rect 7840 16300 7874 16334
rect 2715 16210 2749 16244
rect 2853 16210 2887 16244
rect 2991 16210 3025 16244
rect 3129 16210 3163 16244
rect 3267 16210 3301 16244
rect 3405 16210 3439 16244
rect 3543 16210 3577 16244
rect 3681 16210 3715 16244
rect 3819 16210 3853 16244
rect 3957 16210 3991 16244
rect 4095 16210 4129 16244
rect 4233 16210 4267 16244
rect 4371 16210 4405 16244
rect 4509 16210 4543 16244
rect 4647 16210 4681 16244
rect 4740 16230 4774 16264
rect 4809 16230 4843 16264
rect 4878 16230 4912 16264
rect 4947 16230 4981 16264
rect 5016 16230 5050 16264
rect 5085 16230 5119 16264
rect 5154 16230 5188 16264
rect 5223 16230 5257 16264
rect 5292 16230 5326 16264
rect 5361 16230 5395 16264
rect 5430 16230 5464 16264
rect 5499 16230 5533 16264
rect 5568 16230 5602 16264
rect 5637 16230 5671 16264
rect 5706 16230 5740 16264
rect 5775 16230 5809 16264
rect 5844 16230 5878 16264
rect 5913 16230 5947 16264
rect 5982 16230 6016 16264
rect 6051 16230 6085 16264
rect 6120 16230 6154 16264
rect 6189 16230 6223 16264
rect 6258 16230 6292 16264
rect 6327 16230 6361 16264
rect 6396 16230 6430 16264
rect 6465 16230 6499 16264
rect 6534 16230 6568 16264
rect 6603 16230 6637 16264
rect 6672 16230 6706 16264
rect 6741 16230 6775 16264
rect 6810 16230 6844 16264
rect 6879 16230 6913 16264
rect 6948 16230 6982 16264
rect 7017 16230 7051 16264
rect 7086 16230 7120 16264
rect 7155 16230 7189 16264
rect 7224 16230 7258 16264
rect 7293 16230 7327 16264
rect 7362 16230 7396 16264
rect 7431 16230 7465 16264
rect 7500 16230 7534 16264
rect 7568 16230 7602 16264
rect 7636 16230 7670 16264
rect 7704 16230 7738 16264
rect 7772 16230 7806 16264
rect 7840 16230 7874 16264
rect 4740 16160 4774 16194
rect 4809 16160 4843 16194
rect 4878 16160 4912 16194
rect 4947 16160 4981 16194
rect 5016 16160 5050 16194
rect 5085 16160 5119 16194
rect 5154 16160 5188 16194
rect 5223 16160 5257 16194
rect 5292 16160 5326 16194
rect 5361 16160 5395 16194
rect 5430 16160 5464 16194
rect 5499 16160 5533 16194
rect 5568 16160 5602 16194
rect 5637 16160 5671 16194
rect 5706 16160 5740 16194
rect 5775 16160 5809 16194
rect 5844 16160 5878 16194
rect 5913 16160 5947 16194
rect 5982 16160 6016 16194
rect 6051 16160 6085 16194
rect 6120 16160 6154 16194
rect 6189 16160 6223 16194
rect 6258 16160 6292 16194
rect 6327 16160 6361 16194
rect 6396 16160 6430 16194
rect 6465 16160 6499 16194
rect 6534 16160 6568 16194
rect 6603 16160 6637 16194
rect 6672 16160 6706 16194
rect 6741 16160 6775 16194
rect 6810 16160 6844 16194
rect 6879 16160 6913 16194
rect 6948 16160 6982 16194
rect 7017 16160 7051 16194
rect 7086 16160 7120 16194
rect 7155 16160 7189 16194
rect 7224 16160 7258 16194
rect 7293 16160 7327 16194
rect 7362 16160 7396 16194
rect 7431 16160 7465 16194
rect 7500 16160 7534 16194
rect 7568 16160 7602 16194
rect 7636 16160 7670 16194
rect 7704 16160 7738 16194
rect 7772 16160 7806 16194
rect 7840 16160 7874 16194
rect 2715 16073 2749 16107
rect 2853 16073 2887 16107
rect 2991 16073 3025 16107
rect 3129 16073 3163 16107
rect 3267 16073 3301 16107
rect 3405 16073 3439 16107
rect 3543 16073 3577 16107
rect 3681 16073 3715 16107
rect 3819 16073 3853 16107
rect 3957 16073 3991 16107
rect 4095 16073 4129 16107
rect 4233 16073 4267 16107
rect 4371 16073 4405 16107
rect 4509 16073 4543 16107
rect 4647 16073 4681 16107
rect 4740 16090 4774 16124
rect 4809 16090 4843 16124
rect 4878 16090 4912 16124
rect 4947 16090 4981 16124
rect 5016 16090 5050 16124
rect 5085 16090 5119 16124
rect 5154 16090 5188 16124
rect 5223 16090 5257 16124
rect 5292 16090 5326 16124
rect 5361 16090 5395 16124
rect 5430 16090 5464 16124
rect 5499 16090 5533 16124
rect 5568 16090 5602 16124
rect 5637 16090 5671 16124
rect 5706 16090 5740 16124
rect 5775 16090 5809 16124
rect 5844 16090 5878 16124
rect 5913 16090 5947 16124
rect 5982 16090 6016 16124
rect 6051 16090 6085 16124
rect 6120 16090 6154 16124
rect 6189 16090 6223 16124
rect 6258 16090 6292 16124
rect 6327 16090 6361 16124
rect 6396 16090 6430 16124
rect 6465 16090 6499 16124
rect 6534 16090 6568 16124
rect 6603 16090 6637 16124
rect 6672 16090 6706 16124
rect 6741 16090 6775 16124
rect 6810 16090 6844 16124
rect 6879 16090 6913 16124
rect 6948 16090 6982 16124
rect 7017 16090 7051 16124
rect 7086 16090 7120 16124
rect 7155 16090 7189 16124
rect 7224 16090 7258 16124
rect 7293 16090 7327 16124
rect 7362 16090 7396 16124
rect 7431 16090 7465 16124
rect 7500 16090 7534 16124
rect 7568 16090 7602 16124
rect 7636 16090 7670 16124
rect 7704 16090 7738 16124
rect 7772 16090 7806 16124
rect 7840 16090 7874 16124
rect 4740 16020 4774 16054
rect 4809 16020 4843 16054
rect 4878 16020 4912 16054
rect 4947 16020 4981 16054
rect 5016 16020 5050 16054
rect 5085 16020 5119 16054
rect 5154 16020 5188 16054
rect 5223 16020 5257 16054
rect 5292 16020 5326 16054
rect 5361 16020 5395 16054
rect 5430 16020 5464 16054
rect 5499 16020 5533 16054
rect 5568 16020 5602 16054
rect 5637 16020 5671 16054
rect 5706 16020 5740 16054
rect 5775 16020 5809 16054
rect 5844 16020 5878 16054
rect 5913 16020 5947 16054
rect 5982 16020 6016 16054
rect 6051 16020 6085 16054
rect 6120 16020 6154 16054
rect 6189 16020 6223 16054
rect 6258 16020 6292 16054
rect 6327 16020 6361 16054
rect 6396 16020 6430 16054
rect 6465 16020 6499 16054
rect 6534 16020 6568 16054
rect 6603 16020 6637 16054
rect 6672 16020 6706 16054
rect 6741 16020 6775 16054
rect 6810 16020 6844 16054
rect 6879 16020 6913 16054
rect 6948 16020 6982 16054
rect 7017 16020 7051 16054
rect 7086 16020 7120 16054
rect 7155 16020 7189 16054
rect 7224 16020 7258 16054
rect 7293 16020 7327 16054
rect 7362 16020 7396 16054
rect 7431 16020 7465 16054
rect 7500 16020 7534 16054
rect 7568 16020 7602 16054
rect 7636 16020 7670 16054
rect 7704 16020 7738 16054
rect 7772 16020 7806 16054
rect 7840 16020 7874 16054
rect 2715 15936 2749 15970
rect 2853 15936 2887 15970
rect 2991 15936 3025 15970
rect 3129 15936 3163 15970
rect 3267 15936 3301 15970
rect 3405 15936 3439 15970
rect 3543 15936 3577 15970
rect 3681 15936 3715 15970
rect 3819 15936 3853 15970
rect 3957 15936 3991 15970
rect 4095 15936 4129 15970
rect 4233 15936 4267 15970
rect 4371 15936 4405 15970
rect 4509 15936 4543 15970
rect 4647 15936 4681 15970
rect 4740 15950 4774 15984
rect 4809 15950 4843 15984
rect 4878 15950 4912 15984
rect 4947 15950 4981 15984
rect 5016 15950 5050 15984
rect 5085 15950 5119 15984
rect 5154 15950 5188 15984
rect 5223 15950 5257 15984
rect 5292 15950 5326 15984
rect 5361 15950 5395 15984
rect 5430 15950 5464 15984
rect 5499 15950 5533 15984
rect 5568 15950 5602 15984
rect 5637 15950 5671 15984
rect 5706 15950 5740 15984
rect 5775 15950 5809 15984
rect 5844 15950 5878 15984
rect 5913 15950 5947 15984
rect 5982 15950 6016 15984
rect 6051 15950 6085 15984
rect 6120 15950 6154 15984
rect 6189 15950 6223 15984
rect 6258 15950 6292 15984
rect 6327 15950 6361 15984
rect 6396 15950 6430 15984
rect 6465 15950 6499 15984
rect 6534 15950 6568 15984
rect 6603 15950 6637 15984
rect 6672 15950 6706 15984
rect 6741 15950 6775 15984
rect 6810 15950 6844 15984
rect 6879 15950 6913 15984
rect 6948 15950 6982 15984
rect 7017 15950 7051 15984
rect 7086 15950 7120 15984
rect 7155 15950 7189 15984
rect 7224 15950 7258 15984
rect 7293 15950 7327 15984
rect 7362 15950 7396 15984
rect 7431 15950 7465 15984
rect 7500 15950 7534 15984
rect 7568 15950 7602 15984
rect 7636 15950 7670 15984
rect 7704 15950 7738 15984
rect 7772 15950 7806 15984
rect 7840 15950 7874 15984
rect 8049 9953 8219 38887
rect 8049 9919 8195 9953
rect 2298 9885 2332 9919
rect 2367 9885 2401 9919
rect 2436 9885 2470 9919
rect 2505 9885 2539 9919
rect 2574 9885 2608 9919
rect 2643 9885 2677 9919
rect 2712 9885 2746 9919
rect 2781 9885 2815 9919
rect 2850 9885 2884 9919
rect 2919 9885 2953 9919
rect 2988 9885 3022 9919
rect 3057 9885 3091 9919
rect 3126 9885 3160 9919
rect 3195 9885 3229 9919
rect 3264 9885 3298 9919
rect 3333 9885 3367 9919
rect 3401 9885 3435 9919
rect 3469 9885 3503 9919
rect 3537 9885 3571 9919
rect 3605 9885 3639 9919
rect 3673 9885 3707 9919
rect 3741 9885 3775 9919
rect 3809 9885 3843 9919
rect 3877 9885 3911 9919
rect 3945 9885 3979 9919
rect 4013 9885 4047 9919
rect 4081 9885 4115 9919
rect 4149 9885 4183 9919
rect 4217 9885 4251 9919
rect 4285 9885 4319 9919
rect 4353 9885 4387 9919
rect 4421 9885 4455 9919
rect 4489 9885 4523 9919
rect 4557 9885 4591 9919
rect 4625 9885 4659 9919
rect 4693 9885 4727 9919
rect 4761 9885 4795 9919
rect 4829 9885 4863 9919
rect 4897 9885 4931 9919
rect 4965 9885 4999 9919
rect 5033 9885 5067 9919
rect 5101 9885 5135 9919
rect 5169 9885 5203 9919
rect 5237 9885 5271 9919
rect 5305 9885 5339 9919
rect 5373 9885 5407 9919
rect 5441 9885 5475 9919
rect 5509 9885 5543 9919
rect 5577 9885 5611 9919
rect 5645 9885 5679 9919
rect 5713 9885 5747 9919
rect 5781 9885 5815 9919
rect 5849 9885 5883 9919
rect 5917 9885 5951 9919
rect 5985 9885 6019 9919
rect 6053 9885 6087 9919
rect 6121 9885 6155 9919
rect 6189 9885 6223 9919
rect 6257 9885 6291 9919
rect 6325 9885 6359 9919
rect 6393 9885 6427 9919
rect 6461 9885 6495 9919
rect 6529 9885 6563 9919
rect 6597 9885 6631 9919
rect 6665 9885 6699 9919
rect 6733 9885 6767 9919
rect 6801 9885 6835 9919
rect 6869 9885 6903 9919
rect 6937 9885 6971 9919
rect 7005 9885 7039 9919
rect 7073 9885 7107 9919
rect 7141 9885 7175 9919
rect 7209 9885 7243 9919
rect 7277 9885 7311 9919
rect 7345 9885 7379 9919
rect 7413 9885 7447 9919
rect 7481 9885 7515 9919
rect 7549 9885 7583 9919
rect 7617 9885 7651 9919
rect 7685 9885 7719 9919
rect 7753 9885 7787 9919
rect 7821 9885 7855 9919
rect 7889 9885 7923 9919
rect 7957 9885 7991 9919
rect 8025 9885 8195 9919
rect 2304 9396 2338 9430
rect 2373 9396 2407 9430
rect 2442 9396 2476 9430
rect 2511 9396 2545 9430
rect 2580 9396 2614 9430
rect 2649 9396 2683 9430
rect 2718 9396 2752 9430
rect 2787 9396 2821 9430
rect 2856 9396 2890 9430
rect 2925 9396 2959 9430
rect 2994 9396 3028 9430
rect 3062 9396 3096 9430
rect 3130 9396 3164 9430
rect 3198 9396 3232 9430
rect 3266 9396 3300 9430
rect 3334 9396 3368 9430
rect 3402 9396 3436 9430
rect 3470 9396 3504 9430
rect 3538 9396 3572 9430
rect 3606 9396 3640 9430
rect 3674 9396 3708 9430
rect 3742 9396 3776 9430
rect 3810 9396 3844 9430
rect 3878 9396 3912 9430
rect 3946 9396 3980 9430
rect 4014 9396 4048 9430
rect 4082 9396 4116 9430
rect 4150 9396 4184 9430
rect 4218 9396 4252 9430
rect 4286 9396 4320 9430
rect 4354 9396 4388 9430
rect 4422 9396 4456 9430
rect 4490 9396 4524 9430
rect 4558 9396 4592 9430
rect 4626 9396 4660 9430
rect 4694 9396 4728 9430
rect 4762 9396 4796 9430
rect 4830 9396 4864 9430
rect 4898 9396 4932 9430
rect 4966 9396 5000 9430
rect 5034 9396 5068 9430
rect 5102 9396 5136 9430
rect 5170 9396 5204 9430
rect 5238 9396 5272 9430
rect 5306 9396 5340 9430
rect 5374 9396 5408 9430
rect 5442 9396 5476 9430
rect 5510 9396 5544 9430
rect 5578 9396 5612 9430
rect 5646 9396 5680 9430
rect 5714 9396 5748 9430
rect 5782 9396 5816 9430
rect 5850 9396 5884 9430
rect 5918 9396 5952 9430
rect 5986 9396 6020 9430
rect 6054 9396 6088 9430
rect 6122 9396 6156 9430
rect 6190 9396 6224 9430
rect 6258 9396 6292 9430
rect 6326 9396 6360 9430
rect 6394 9396 6428 9430
rect 6462 9396 6496 9430
rect 6530 9396 6564 9430
rect 6598 9396 6632 9430
rect 6666 9396 6700 9430
rect 6734 9396 6768 9430
rect 6802 9396 6836 9430
rect 6870 9396 6904 9430
rect 6938 9396 6972 9430
rect 7006 9396 7040 9430
rect 7074 9396 7108 9430
rect 7142 9396 7176 9430
rect 7210 9396 7244 9430
rect 7278 9396 7312 9430
rect 7346 9396 7380 9430
rect 7414 9396 7448 9430
rect 2290 9328 2324 9362
rect 2290 9260 2324 9294
rect 7487 9336 7521 9370
rect 2290 9192 2324 9226
rect 2290 9124 2324 9158
rect 2290 9056 2324 9090
rect 2290 8988 2324 9022
rect 2290 8920 2324 8954
rect 2290 8852 2324 8886
rect 2290 8784 2324 8818
rect 2290 8716 2324 8750
rect 2290 8648 2324 8682
rect 2290 8580 2324 8614
rect 2290 8512 2324 8546
rect 2290 8444 2324 8478
rect 2290 8376 2324 8410
rect 2290 8308 2324 8342
rect 2290 8240 2324 8274
rect 2290 8172 2324 8206
rect 2290 8104 2324 8138
rect 2290 8036 2324 8070
rect 2290 7968 2324 8002
rect 2290 7900 2324 7934
rect 2290 7832 2324 7866
rect 2290 7764 2324 7798
rect 2290 7696 2324 7730
rect 7487 9268 7521 9302
rect 7487 9200 7521 9234
rect 7487 9132 7521 9166
rect 7487 9064 7521 9098
rect 7487 8996 7521 9030
rect 7487 8928 7521 8962
rect 7487 8860 7521 8894
rect 7487 8792 7521 8826
rect 7487 8724 7521 8758
rect 7487 8656 7521 8690
rect 7487 8588 7521 8622
rect 7487 8520 7521 8554
rect 7487 8452 7521 8486
rect 7487 8384 7521 8418
rect 7487 8316 7521 8350
rect 7487 8248 7521 8282
rect 7487 8180 7521 8214
rect 7487 8112 7521 8146
rect 7487 8044 7521 8078
rect 7487 7976 7521 8010
rect 7487 7908 7521 7942
rect 7487 7840 7521 7874
rect 7487 7772 7521 7806
rect 7487 7704 7521 7738
rect 2290 7628 2324 7662
rect 2358 7647 2392 7681
rect 2427 7647 2461 7681
rect 2496 7647 2530 7681
rect 2565 7647 2599 7681
rect 2634 7647 2668 7681
rect 2703 7647 2737 7681
rect 2772 7647 2806 7681
rect 2841 7647 2875 7681
rect 2910 7647 2944 7681
rect 2979 7647 3013 7681
rect 3048 7647 3082 7681
rect 3117 7647 3151 7681
rect 3186 7647 3220 7681
rect 3255 7647 3289 7681
rect 3324 7647 3358 7681
rect 3393 7647 3427 7681
rect 3462 7647 3496 7681
rect 3531 7647 3565 7681
rect 3600 7647 3634 7681
rect 3669 7647 3703 7681
rect 3738 7647 3772 7681
rect 3807 7647 3841 7681
rect 3875 7647 3909 7681
rect 3943 7647 3977 7681
rect 4011 7647 4045 7681
rect 4079 7647 4113 7681
rect 4147 7647 4181 7681
rect 4215 7647 4249 7681
rect 4283 7647 4317 7681
rect 4351 7647 4385 7681
rect 4419 7647 4453 7681
rect 4487 7647 4521 7681
rect 4555 7647 4589 7681
rect 4623 7647 4657 7681
rect 4691 7647 4725 7681
rect 4759 7647 4793 7681
rect 4827 7647 4861 7681
rect 4895 7647 4929 7681
rect 4963 7647 4997 7681
rect 5031 7647 5065 7681
rect 5099 7647 5133 7681
rect 5167 7647 5201 7681
rect 5235 7647 5269 7681
rect 5303 7647 5337 7681
rect 5371 7647 5405 7681
rect 5439 7647 5473 7681
rect 5507 7647 5541 7681
rect 5575 7647 5609 7681
rect 5643 7647 5677 7681
rect 5711 7647 5745 7681
rect 5779 7647 5813 7681
rect 5847 7647 5881 7681
rect 5915 7647 5949 7681
rect 5983 7647 6017 7681
rect 6051 7647 6085 7681
rect 6119 7647 6153 7681
rect 6187 7647 6221 7681
rect 6255 7647 6289 7681
rect 6323 7647 6357 7681
rect 6391 7647 6425 7681
rect 6459 7647 6493 7681
rect 6527 7647 6561 7681
rect 6595 7647 6629 7681
rect 6663 7647 6697 7681
rect 6731 7647 6765 7681
rect 6799 7647 6833 7681
rect 6867 7647 6901 7681
rect 6935 7647 6969 7681
rect 7003 7647 7037 7681
rect 7071 7647 7105 7681
rect 7139 7647 7173 7681
rect 7207 7647 7241 7681
rect 7275 7647 7309 7681
rect 7343 7647 7377 7681
rect 7411 7647 7445 7681
rect 2290 7560 2324 7594
rect 7487 7636 7521 7670
rect 7487 7568 7521 7602
rect 2290 7492 2324 7526
rect 7487 7500 7521 7534
rect 2290 7424 2324 7458
rect 2290 7356 2324 7390
rect 2290 7288 2324 7322
rect 2290 7220 2324 7254
rect 2290 7152 2324 7186
rect 2290 7084 2324 7118
rect 2290 7016 2324 7050
rect 2290 6948 2324 6982
rect 2290 6880 2324 6914
rect 2290 6812 2324 6846
rect 2290 6744 2324 6778
rect 2290 6676 2324 6710
rect 2290 6608 2324 6642
rect 2290 6540 2324 6574
rect 2290 6472 2324 6506
rect 2290 6404 2324 6438
rect 2290 6336 2324 6370
rect 2290 6268 2324 6302
rect 2290 6200 2324 6234
rect 2290 6132 2324 6166
rect 2290 6064 2324 6098
rect 2290 5996 2324 6030
rect 2290 5928 2324 5962
rect 2290 5860 2324 5894
rect 7487 7432 7521 7466
rect 7487 7364 7521 7398
rect 7487 7296 7521 7330
rect 7487 7228 7521 7262
rect 7487 7160 7521 7194
rect 7487 7092 7521 7126
rect 7487 7024 7521 7058
rect 7487 6956 7521 6990
rect 7487 6888 7521 6922
rect 7487 6820 7521 6854
rect 7487 6752 7521 6786
rect 7487 6684 7521 6718
rect 7487 6616 7521 6650
rect 7487 6548 7521 6582
rect 7487 6480 7521 6514
rect 7487 6412 7521 6446
rect 7487 6344 7521 6378
rect 7487 6276 7521 6310
rect 7487 6208 7521 6242
rect 7487 6140 7521 6174
rect 7487 6072 7521 6106
rect 7487 6004 7521 6038
rect 7487 5936 7521 5970
rect 7487 5868 7521 5902
rect 2290 5792 2324 5826
rect 2358 5807 2392 5841
rect 2427 5807 2461 5841
rect 2496 5807 2530 5841
rect 2565 5807 2599 5841
rect 2634 5807 2668 5841
rect 2703 5807 2737 5841
rect 2772 5807 2806 5841
rect 2841 5807 2875 5841
rect 2910 5807 2944 5841
rect 2979 5807 3013 5841
rect 3048 5807 3082 5841
rect 3117 5807 3151 5841
rect 3186 5807 3220 5841
rect 3255 5807 3289 5841
rect 3324 5807 3358 5841
rect 3393 5807 3427 5841
rect 3462 5807 3496 5841
rect 3531 5807 3565 5841
rect 3600 5807 3634 5841
rect 3669 5807 3703 5841
rect 3737 5807 3771 5841
rect 3805 5807 3839 5841
rect 3873 5807 3907 5841
rect 3941 5807 3975 5841
rect 4009 5807 4043 5841
rect 4077 5807 4111 5841
rect 4145 5807 4179 5841
rect 4213 5807 4247 5841
rect 4281 5807 4315 5841
rect 4349 5807 4383 5841
rect 4417 5807 4451 5841
rect 4485 5807 4519 5841
rect 4553 5807 4587 5841
rect 4621 5807 4655 5841
rect 4689 5807 4723 5841
rect 4757 5807 4791 5841
rect 4825 5807 4859 5841
rect 4893 5807 4927 5841
rect 4961 5807 4995 5841
rect 5029 5807 5063 5841
rect 5097 5807 5131 5841
rect 5165 5807 5199 5841
rect 5233 5807 5267 5841
rect 5301 5807 5335 5841
rect 5369 5807 5403 5841
rect 5437 5807 5471 5841
rect 5505 5807 5539 5841
rect 5573 5807 5607 5841
rect 5641 5807 5675 5841
rect 5709 5807 5743 5841
rect 5777 5807 5811 5841
rect 5845 5807 5879 5841
rect 5913 5807 5947 5841
rect 5981 5807 6015 5841
rect 6049 5807 6083 5841
rect 6117 5807 6151 5841
rect 6185 5807 6219 5841
rect 6253 5807 6287 5841
rect 6321 5807 6355 5841
rect 6389 5807 6423 5841
rect 6457 5807 6491 5841
rect 6525 5807 6559 5841
rect 6593 5807 6627 5841
rect 6661 5807 6695 5841
rect 6729 5807 6763 5841
rect 6797 5807 6831 5841
rect 6865 5807 6899 5841
rect 6933 5807 6967 5841
rect 7001 5807 7035 5841
rect 7069 5807 7103 5841
rect 7137 5807 7171 5841
rect 7205 5807 7239 5841
rect 7273 5807 7307 5841
rect 7341 5807 7375 5841
rect 7409 5807 7443 5841
rect 2290 5724 2324 5758
rect 2290 5656 2324 5690
rect 7487 5800 7521 5834
rect 7487 5732 7521 5766
rect 7487 5664 7521 5698
rect 2290 5588 2324 5622
rect 7487 5596 7521 5630
rect 2290 5520 2324 5554
rect 2290 5452 2324 5486
rect 2290 5384 2324 5418
rect 2290 5316 2324 5350
rect 2290 5248 2324 5282
rect 2290 5180 2324 5214
rect 2290 5112 2324 5146
rect 2290 5044 2324 5078
rect 2290 4976 2324 5010
rect 2290 4908 2324 4942
rect 2290 4840 2324 4874
rect 2290 4772 2324 4806
rect 2290 4704 2324 4738
rect 2290 4636 2324 4670
rect 2290 4568 2324 4602
rect 2290 4500 2324 4534
rect 2290 4432 2324 4466
rect 2290 4364 2324 4398
rect 2290 4296 2324 4330
rect 2290 4228 2324 4262
rect 2290 4160 2324 4194
rect 2290 4092 2324 4126
rect 2290 4024 2324 4058
rect 7487 5528 7521 5562
rect 7487 5460 7521 5494
rect 7487 5392 7521 5426
rect 7487 5324 7521 5358
rect 7487 5256 7521 5290
rect 7487 5188 7521 5222
rect 7487 5120 7521 5154
rect 7487 5052 7521 5086
rect 7487 4984 7521 5018
rect 7487 4916 7521 4950
rect 7487 4848 7521 4882
rect 7487 4780 7521 4814
rect 7487 4712 7521 4746
rect 7487 4644 7521 4678
rect 7487 4576 7521 4610
rect 7487 4508 7521 4542
rect 7487 4440 7521 4474
rect 7487 4372 7521 4406
rect 7487 4304 7521 4338
rect 7487 4236 7521 4270
rect 7487 4168 7521 4202
rect 7487 4100 7521 4134
rect 7487 4032 7521 4066
rect 7487 3964 7521 3998
rect 2314 3873 2348 3907
rect 2382 3873 2416 3907
rect 2450 3873 2484 3907
rect 2518 3873 2552 3907
rect 2586 3873 2620 3907
rect 2654 3873 2688 3907
rect 2722 3873 2756 3907
rect 2790 3873 2824 3907
rect 2858 3873 2892 3907
rect 2926 3873 2960 3907
rect 2994 3873 3028 3907
rect 3062 3873 3096 3907
rect 3130 3873 3164 3907
rect 3198 3873 3232 3907
rect 3266 3873 3300 3907
rect 3334 3873 3368 3907
rect 3402 3873 3436 3907
rect 3470 3873 3504 3907
rect 3538 3873 3572 3907
rect 3606 3873 3640 3907
rect 3674 3873 3708 3907
rect 3742 3873 3776 3907
rect 3810 3873 3844 3907
rect 3878 3873 3912 3907
rect 3946 3873 3980 3907
rect 4014 3873 4048 3907
rect 4082 3873 4116 3907
rect 4150 3873 4184 3907
rect 4218 3873 4252 3907
rect 4286 3873 4320 3907
rect 4354 3873 4388 3907
rect 4422 3873 4456 3907
rect 4490 3873 4524 3907
rect 4558 3873 4592 3907
rect 4626 3873 4660 3907
rect 4694 3873 4728 3907
rect 4762 3873 4796 3907
rect 4830 3873 4864 3907
rect 4898 3873 4932 3907
rect 4966 3873 5000 3907
rect 5034 3873 5068 3907
rect 5102 3873 5136 3907
rect 5170 3873 5204 3907
rect 5238 3873 5272 3907
rect 5306 3873 5340 3907
rect 5374 3873 5408 3907
rect 5442 3873 5476 3907
rect 5510 3873 5544 3907
rect 5578 3873 5612 3907
rect 5646 3873 5680 3907
rect 5714 3873 5748 3907
rect 5782 3873 5816 3907
rect 5850 3873 5884 3907
rect 5918 3873 5952 3907
rect 5986 3873 6020 3907
rect 6054 3873 6088 3907
rect 6122 3873 6156 3907
rect 6190 3873 6224 3907
rect 6258 3873 6292 3907
rect 6326 3873 6360 3907
rect 6394 3873 6428 3907
rect 6462 3873 6496 3907
rect 6530 3873 6564 3907
rect 6598 3873 6632 3907
rect 6666 3873 6700 3907
rect 6734 3873 6768 3907
rect 6802 3873 6836 3907
rect 6870 3873 6904 3907
rect 6938 3873 6972 3907
rect 7006 3873 7040 3907
rect 7074 3873 7108 3907
rect 7142 3873 7176 3907
rect 7210 3873 7244 3907
rect 7278 3873 7312 3907
rect 7346 3873 7380 3907
rect 7414 3873 7448 3907
rect 1855 3092 1889 3126
rect 1992 3092 2026 3126
rect 2129 3092 2163 3126
rect 2266 3092 2300 3126
rect 2403 3092 2437 3126
rect 2540 3092 2574 3126
rect 2677 3092 2711 3126
rect 2814 3092 2848 3126
rect 2950 3092 2984 3126
rect 3086 3092 3120 3126
rect 3222 3092 3256 3126
rect 3358 3092 3392 3126
rect 3494 3092 3528 3126
rect 3630 3092 3664 3126
rect 3766 3092 3800 3126
rect 3902 3092 3936 3126
rect 4038 3092 4072 3126
rect 4174 3092 4208 3126
rect 4310 3092 4344 3126
rect 4446 3092 4480 3126
rect 4582 3092 4616 3126
rect 4718 3092 4752 3126
rect 4854 3092 4888 3126
rect 4990 3092 5024 3126
rect 5126 3092 5160 3126
rect 5262 3092 5296 3126
rect 5398 3092 5432 3126
rect 5534 3092 5568 3126
rect 5670 3092 5704 3126
rect 5806 3092 5840 3126
rect 5942 3092 5976 3126
rect 6078 3092 6112 3126
rect 6214 3092 6248 3126
rect 6350 3092 6384 3126
rect 6486 3092 6520 3126
rect 6622 3092 6656 3126
rect 6758 3092 6792 3126
rect 6894 3092 6928 3126
rect 7030 3092 7064 3126
rect 7166 3092 7200 3126
rect 7302 3092 7336 3126
rect 7438 3092 7472 3126
rect 7574 3092 7608 3126
rect 7710 3092 7744 3126
rect 7846 3092 7880 3126
rect 1855 2976 1889 3010
rect 1992 2976 2026 3010
rect 2129 2976 2163 3010
rect 2266 2976 2300 3010
rect 2403 2976 2437 3010
rect 2540 2976 2574 3010
rect 2677 2976 2711 3010
rect 2814 2976 2848 3010
rect 2950 2976 2984 3010
rect 3086 2976 3120 3010
rect 3222 2976 3256 3010
rect 3358 2976 3392 3010
rect 3494 2976 3528 3010
rect 3630 2976 3664 3010
rect 3766 2976 3800 3010
rect 3902 2976 3936 3010
rect 4038 2976 4072 3010
rect 4174 2976 4208 3010
rect 4310 2976 4344 3010
rect 4446 2976 4480 3010
rect 4582 2976 4616 3010
rect 4718 2976 4752 3010
rect 4854 2976 4888 3010
rect 4990 2976 5024 3010
rect 5126 2976 5160 3010
rect 5262 2976 5296 3010
rect 5398 2976 5432 3010
rect 5534 2976 5568 3010
rect 5670 2976 5704 3010
rect 5806 2976 5840 3010
rect 5942 2976 5976 3010
rect 6078 2976 6112 3010
rect 6214 2976 6248 3010
rect 6350 2976 6384 3010
rect 6486 2976 6520 3010
rect 6622 2976 6656 3010
rect 6758 2976 6792 3010
rect 6894 2976 6928 3010
rect 7030 2976 7064 3010
rect 7166 2976 7200 3010
rect 7302 2976 7336 3010
rect 7438 2976 7472 3010
rect 7574 2976 7608 3010
rect 7710 2976 7744 3010
rect 7846 2976 7880 3010
rect 1855 2860 1889 2894
rect 1992 2860 2026 2894
rect 2129 2860 2163 2894
rect 2266 2860 2300 2894
rect 2403 2860 2437 2894
rect 2540 2860 2574 2894
rect 2677 2860 2711 2894
rect 2814 2860 2848 2894
rect 2950 2860 2984 2894
rect 3086 2860 3120 2894
rect 3222 2860 3256 2894
rect 3358 2860 3392 2894
rect 3494 2860 3528 2894
rect 3630 2860 3664 2894
rect 3766 2860 3800 2894
rect 3902 2860 3936 2894
rect 4038 2860 4072 2894
rect 4174 2860 4208 2894
rect 4310 2860 4344 2894
rect 4446 2860 4480 2894
rect 4582 2860 4616 2894
rect 4718 2860 4752 2894
rect 4854 2860 4888 2894
rect 4990 2860 5024 2894
rect 5126 2860 5160 2894
rect 5262 2860 5296 2894
rect 5398 2860 5432 2894
rect 5534 2860 5568 2894
rect 5670 2860 5704 2894
rect 5806 2860 5840 2894
rect 5942 2860 5976 2894
rect 6078 2860 6112 2894
rect 6214 2860 6248 2894
rect 6350 2860 6384 2894
rect 6486 2860 6520 2894
rect 6622 2860 6656 2894
rect 6758 2860 6792 2894
rect 6894 2860 6928 2894
rect 7030 2860 7064 2894
rect 7166 2860 7200 2894
rect 7302 2860 7336 2894
rect 7438 2860 7472 2894
rect 7574 2860 7608 2894
rect 7710 2860 7744 2894
rect 7846 2860 7880 2894
rect 1855 2744 1889 2778
rect 1992 2744 2026 2778
rect 2129 2744 2163 2778
rect 2266 2744 2300 2778
rect 2403 2744 2437 2778
rect 2540 2744 2574 2778
rect 2677 2744 2711 2778
rect 2814 2744 2848 2778
rect 2950 2744 2984 2778
rect 3086 2744 3120 2778
rect 3222 2744 3256 2778
rect 3358 2744 3392 2778
rect 3494 2744 3528 2778
rect 3630 2744 3664 2778
rect 3766 2744 3800 2778
rect 3902 2744 3936 2778
rect 4038 2744 4072 2778
rect 4174 2744 4208 2778
rect 4310 2744 4344 2778
rect 4446 2744 4480 2778
rect 4582 2744 4616 2778
rect 4718 2744 4752 2778
rect 4854 2744 4888 2778
rect 4990 2744 5024 2778
rect 5126 2744 5160 2778
rect 5262 2744 5296 2778
rect 5398 2744 5432 2778
rect 5534 2744 5568 2778
rect 5670 2744 5704 2778
rect 5806 2744 5840 2778
rect 5942 2744 5976 2778
rect 6078 2744 6112 2778
rect 6214 2744 6248 2778
rect 6350 2744 6384 2778
rect 6486 2744 6520 2778
rect 6622 2744 6656 2778
rect 6758 2744 6792 2778
rect 6894 2744 6928 2778
rect 7030 2744 7064 2778
rect 7166 2744 7200 2778
rect 7302 2744 7336 2778
rect 7438 2744 7472 2778
rect 7574 2744 7608 2778
rect 7710 2744 7744 2778
rect 7846 2744 7880 2778
rect 1855 2628 1889 2662
rect 1992 2628 2026 2662
rect 2129 2628 2163 2662
rect 2266 2628 2300 2662
rect 2403 2628 2437 2662
rect 2540 2628 2574 2662
rect 2677 2628 2711 2662
rect 2814 2628 2848 2662
rect 2950 2628 2984 2662
rect 3086 2628 3120 2662
rect 3222 2628 3256 2662
rect 3358 2628 3392 2662
rect 3494 2628 3528 2662
rect 3630 2628 3664 2662
rect 3766 2628 3800 2662
rect 3902 2628 3936 2662
rect 4038 2628 4072 2662
rect 4174 2628 4208 2662
rect 4310 2628 4344 2662
rect 4446 2628 4480 2662
rect 4582 2628 4616 2662
rect 4718 2628 4752 2662
rect 4854 2628 4888 2662
rect 4990 2628 5024 2662
rect 5126 2628 5160 2662
rect 5262 2628 5296 2662
rect 5398 2628 5432 2662
rect 5534 2628 5568 2662
rect 5670 2628 5704 2662
rect 5806 2628 5840 2662
rect 5942 2628 5976 2662
rect 6078 2628 6112 2662
rect 6214 2628 6248 2662
rect 6350 2628 6384 2662
rect 6486 2628 6520 2662
rect 6622 2628 6656 2662
rect 6758 2628 6792 2662
rect 6894 2628 6928 2662
rect 7030 2628 7064 2662
rect 7166 2628 7200 2662
rect 7302 2628 7336 2662
rect 7438 2628 7472 2662
rect 7574 2628 7608 2662
rect 7710 2628 7744 2662
rect 7846 2628 7880 2662
rect 1855 2512 1889 2546
rect 1992 2512 2026 2546
rect 2129 2512 2163 2546
rect 2266 2512 2300 2546
rect 2403 2512 2437 2546
rect 2540 2512 2574 2546
rect 2677 2512 2711 2546
rect 2814 2512 2848 2546
rect 2950 2512 2984 2546
rect 3086 2512 3120 2546
rect 3222 2512 3256 2546
rect 3358 2512 3392 2546
rect 3494 2512 3528 2546
rect 3630 2512 3664 2546
rect 3766 2512 3800 2546
rect 3902 2512 3936 2546
rect 4038 2512 4072 2546
rect 4174 2512 4208 2546
rect 4310 2512 4344 2546
rect 4446 2512 4480 2546
rect 4582 2512 4616 2546
rect 4718 2512 4752 2546
rect 4854 2512 4888 2546
rect 4990 2512 5024 2546
rect 5126 2512 5160 2546
rect 5262 2512 5296 2546
rect 5398 2512 5432 2546
rect 5534 2512 5568 2546
rect 5670 2512 5704 2546
rect 5806 2512 5840 2546
rect 5942 2512 5976 2546
rect 6078 2512 6112 2546
rect 6214 2512 6248 2546
rect 6350 2512 6384 2546
rect 6486 2512 6520 2546
rect 6622 2512 6656 2546
rect 6758 2512 6792 2546
rect 6894 2512 6928 2546
rect 7030 2512 7064 2546
rect 7166 2512 7200 2546
rect 7302 2512 7336 2546
rect 7438 2512 7472 2546
rect 7574 2512 7608 2546
rect 7710 2512 7744 2546
rect 7846 2512 7880 2546
rect 1855 2396 1889 2430
rect 1992 2396 2026 2430
rect 2129 2396 2163 2430
rect 2266 2396 2300 2430
rect 2403 2396 2437 2430
rect 2540 2396 2574 2430
rect 2677 2396 2711 2430
rect 2814 2396 2848 2430
rect 2950 2396 2984 2430
rect 3086 2396 3120 2430
rect 3222 2396 3256 2430
rect 3358 2396 3392 2430
rect 3494 2396 3528 2430
rect 3630 2396 3664 2430
rect 3766 2396 3800 2430
rect 3902 2396 3936 2430
rect 4038 2396 4072 2430
rect 4174 2396 4208 2430
rect 4310 2396 4344 2430
rect 4446 2396 4480 2430
rect 4582 2396 4616 2430
rect 4718 2396 4752 2430
rect 4854 2396 4888 2430
rect 4990 2396 5024 2430
rect 5126 2396 5160 2430
rect 5262 2396 5296 2430
rect 5398 2396 5432 2430
rect 5534 2396 5568 2430
rect 5670 2396 5704 2430
rect 5806 2396 5840 2430
rect 5942 2396 5976 2430
rect 6078 2396 6112 2430
rect 6214 2396 6248 2430
rect 6350 2396 6384 2430
rect 6486 2396 6520 2430
rect 6622 2396 6656 2430
rect 6758 2396 6792 2430
rect 6894 2396 6928 2430
rect 7030 2396 7064 2430
rect 7166 2396 7200 2430
rect 7302 2396 7336 2430
rect 7438 2396 7472 2430
rect 7574 2396 7608 2430
rect 7710 2396 7744 2430
rect 7846 2396 7880 2430
rect 5346 2327 5380 2361
rect 5484 2327 5518 2361
rect 5622 2327 5656 2361
rect 5760 2327 5794 2361
rect 5898 2327 5932 2361
rect 6036 2327 6070 2361
rect 6174 2327 6208 2361
rect 6312 2327 6346 2361
rect 6450 2327 6484 2361
rect 6588 2327 6622 2361
rect 6726 2327 6760 2361
rect 6864 2327 6898 2361
rect 7002 2327 7036 2361
rect 7140 2327 7174 2361
rect 7278 2327 7312 2361
rect 7416 2327 7450 2361
rect 7554 2327 7588 2361
rect 5346 2189 5380 2223
rect 5484 2189 5518 2223
rect 5622 2189 5656 2223
rect 5760 2189 5794 2223
rect 5898 2189 5932 2223
rect 6036 2189 6070 2223
rect 6174 2189 6208 2223
rect 6312 2189 6346 2223
rect 6450 2189 6484 2223
rect 6588 2189 6622 2223
rect 6726 2189 6760 2223
rect 6864 2189 6898 2223
rect 7002 2189 7036 2223
rect 7140 2189 7174 2223
rect 7278 2189 7312 2223
rect 7416 2189 7450 2223
rect 7554 2189 7588 2223
rect 5346 2051 5380 2085
rect 5484 2051 5518 2085
rect 5622 2051 5656 2085
rect 5760 2051 5794 2085
rect 5898 2051 5932 2085
rect 6036 2051 6070 2085
rect 6174 2051 6208 2085
rect 6312 2051 6346 2085
rect 6450 2051 6484 2085
rect 6588 2051 6622 2085
rect 6726 2051 6760 2085
rect 6864 2051 6898 2085
rect 7002 2051 7036 2085
rect 7140 2051 7174 2085
rect 7278 2051 7312 2085
rect 7416 2051 7450 2085
rect 7554 2051 7588 2085
rect 5346 1913 5380 1947
rect 5484 1913 5518 1947
rect 5622 1913 5656 1947
rect 5760 1913 5794 1947
rect 5898 1913 5932 1947
rect 6036 1913 6070 1947
rect 6174 1913 6208 1947
rect 6312 1913 6346 1947
rect 6450 1913 6484 1947
rect 6588 1913 6622 1947
rect 6726 1913 6760 1947
rect 6864 1913 6898 1947
rect 7002 1913 7036 1947
rect 7140 1913 7174 1947
rect 7278 1913 7312 1947
rect 7416 1913 7450 1947
rect 7554 1913 7588 1947
rect 5346 1775 5380 1809
rect 5484 1775 5518 1809
rect 5622 1775 5656 1809
rect 5760 1775 5794 1809
rect 5898 1775 5932 1809
rect 6036 1775 6070 1809
rect 6174 1775 6208 1809
rect 6312 1775 6346 1809
rect 6450 1775 6484 1809
rect 6588 1775 6622 1809
rect 6726 1775 6760 1809
rect 6864 1775 6898 1809
rect 7002 1775 7036 1809
rect 7140 1775 7174 1809
rect 7278 1775 7312 1809
rect 7416 1775 7450 1809
rect 7554 1775 7588 1809
rect 5346 1637 5380 1671
rect 5484 1637 5518 1671
rect 5622 1637 5656 1671
rect 5760 1637 5794 1671
rect 5898 1637 5932 1671
rect 6036 1637 6070 1671
rect 6174 1637 6208 1671
rect 6312 1637 6346 1671
rect 6450 1637 6484 1671
rect 6588 1637 6622 1671
rect 6726 1637 6760 1671
rect 6864 1637 6898 1671
rect 7002 1637 7036 1671
rect 7140 1637 7174 1671
rect 7278 1637 7312 1671
rect 7416 1637 7450 1671
rect 7554 1637 7588 1671
rect 5346 1498 5380 1532
rect 5484 1498 5518 1532
rect 5622 1498 5656 1532
rect 5760 1498 5794 1532
rect 5898 1498 5932 1532
rect 6036 1498 6070 1532
rect 6174 1498 6208 1532
rect 6312 1498 6346 1532
rect 6450 1498 6484 1532
rect 6588 1498 6622 1532
rect 6726 1498 6760 1532
rect 6864 1498 6898 1532
rect 7002 1498 7036 1532
rect 7140 1498 7174 1532
rect 7278 1498 7312 1532
rect 7416 1498 7450 1532
rect 7554 1498 7588 1532
rect 5346 1359 5380 1393
rect 5484 1359 5518 1393
rect 5622 1359 5656 1393
rect 5760 1359 5794 1393
rect 5898 1359 5932 1393
rect 6036 1359 6070 1393
rect 6174 1359 6208 1393
rect 6312 1359 6346 1393
rect 6450 1359 6484 1393
rect 6588 1359 6622 1393
rect 6726 1359 6760 1393
rect 6864 1359 6898 1393
rect 7002 1359 7036 1393
rect 7140 1359 7174 1393
rect 7278 1359 7312 1393
rect 7416 1359 7450 1393
rect 7554 1359 7588 1393
rect 5346 1220 5380 1254
rect 5484 1220 5518 1254
rect 5622 1220 5656 1254
rect 5760 1220 5794 1254
rect 5898 1220 5932 1254
rect 6036 1220 6070 1254
rect 6174 1220 6208 1254
rect 6312 1220 6346 1254
rect 6450 1220 6484 1254
rect 6588 1220 6622 1254
rect 6726 1220 6760 1254
rect 6864 1220 6898 1254
rect 7002 1220 7036 1254
rect 7140 1220 7174 1254
rect 7278 1220 7312 1254
rect 7416 1220 7450 1254
rect 7554 1220 7588 1254
rect 5346 1081 5380 1115
rect 5484 1081 5518 1115
rect 5622 1081 5656 1115
rect 5760 1081 5794 1115
rect 5898 1081 5932 1115
rect 6036 1081 6070 1115
rect 6174 1081 6208 1115
rect 6312 1081 6346 1115
rect 6450 1081 6484 1115
rect 6588 1081 6622 1115
rect 6726 1081 6760 1115
rect 6864 1081 6898 1115
rect 7002 1081 7036 1115
rect 7140 1081 7174 1115
rect 7278 1081 7312 1115
rect 7416 1081 7450 1115
rect 7554 1081 7588 1115
rect 5346 942 5380 976
rect 5484 942 5518 976
rect 5622 942 5656 976
rect 5760 942 5794 976
rect 5898 942 5932 976
rect 6036 942 6070 976
rect 6174 942 6208 976
rect 6312 942 6346 976
rect 6450 942 6484 976
rect 6588 942 6622 976
rect 6726 942 6760 976
rect 6864 942 6898 976
rect 7002 942 7036 976
rect 7140 942 7174 976
rect 7278 942 7312 976
rect 7416 942 7450 976
rect 7554 942 7588 976
rect 5346 803 5380 837
rect 5484 803 5518 837
rect 5622 803 5656 837
rect 5760 803 5794 837
rect 5898 803 5932 837
rect 6036 803 6070 837
rect 6174 803 6208 837
rect 6312 803 6346 837
rect 6450 803 6484 837
rect 6588 803 6622 837
rect 6726 803 6760 837
rect 6864 803 6898 837
rect 7002 803 7036 837
rect 7140 803 7174 837
rect 7278 803 7312 837
rect 7416 803 7450 837
rect 7554 803 7588 837
rect 5346 664 5380 698
rect 5484 664 5518 698
rect 5622 664 5656 698
rect 5760 664 5794 698
rect 5898 664 5932 698
rect 6036 664 6070 698
rect 6174 664 6208 698
rect 6312 664 6346 698
rect 6450 664 6484 698
rect 6588 664 6622 698
rect 6726 664 6760 698
rect 6864 664 6898 698
rect 7002 664 7036 698
rect 7140 664 7174 698
rect 7278 664 7312 698
rect 7416 664 7450 698
rect 7554 664 7588 698
rect 5346 525 5380 559
rect 5484 525 5518 559
rect 5622 525 5656 559
rect 5760 525 5794 559
rect 5898 525 5932 559
rect 6036 525 6070 559
rect 6174 525 6208 559
rect 6312 525 6346 559
rect 6450 525 6484 559
rect 6588 525 6622 559
rect 6726 525 6760 559
rect 6864 525 6898 559
rect 7002 525 7036 559
rect 7140 525 7174 559
rect 7278 525 7312 559
rect 7416 525 7450 559
rect 7554 525 7588 559
rect 5346 386 5380 420
rect 5484 386 5518 420
rect 5622 386 5656 420
rect 5760 386 5794 420
rect 5898 386 5932 420
rect 6036 386 6070 420
rect 6174 386 6208 420
rect 6312 386 6346 420
rect 6450 386 6484 420
rect 6588 386 6622 420
rect 6726 386 6760 420
rect 6864 386 6898 420
rect 7002 386 7036 420
rect 7140 386 7174 420
rect 7278 386 7312 420
rect 7416 386 7450 420
rect 7554 386 7588 420
<< nsubdiffcont >>
rect 1869 1982 1903 2016
rect 1937 1982 1971 2016
rect 2005 1982 2039 2016
rect 2073 1982 2107 2016
rect 2141 1982 2175 2016
rect 2209 1982 2243 2016
rect 2277 1982 2311 2016
rect 2345 1982 2379 2016
rect 2413 1982 2447 2016
rect 2481 1982 2515 2016
rect 2549 1982 2583 2016
rect 2617 1982 2651 2016
rect 2685 1982 2719 2016
rect 2753 1982 2787 2016
rect 2821 1982 2855 2016
rect 2889 1982 2923 2016
rect 2957 1982 2991 2016
rect 3025 1982 3059 2016
rect 3093 1982 3127 2016
rect 3161 1982 3195 2016
rect 3229 1982 3263 2016
rect 3297 1982 3331 2016
rect 3365 1982 3399 2016
rect 3433 1982 3467 2016
rect 3501 1982 3535 2016
rect 3569 1982 3603 2016
rect 3637 1982 3671 2016
rect 3705 1982 3739 2016
rect 3773 1982 3807 2016
rect 3841 1982 3875 2016
rect 3909 1982 3943 2016
rect 3977 1982 4011 2016
rect 4045 1982 4079 2016
rect 4113 1982 4147 2016
rect 4181 1982 4215 2016
rect 4249 1982 4283 2016
rect 4317 1982 4351 2016
rect 4385 1982 4419 2016
rect 4453 1982 4487 2016
rect 4521 1982 4555 2016
rect 4589 1982 4623 2016
rect 4657 1982 4691 2016
rect 4725 1982 4759 2016
rect 4793 1982 4827 2016
rect 4861 1982 4895 2016
rect 4929 1982 4963 2016
rect 1801 1884 1835 1918
rect 5005 1914 5039 1948
rect 1801 1816 1835 1850
rect 1801 1748 1835 1782
rect 1801 1680 1835 1714
rect 1801 1612 1835 1646
rect 1801 1544 1835 1578
rect 1801 1476 1835 1510
rect 1801 1408 1835 1442
rect 1801 1340 1835 1374
rect 1801 1272 1835 1306
rect 1801 1204 1835 1238
rect 1801 1136 1835 1170
rect 1801 1068 1835 1102
rect 1801 1000 1835 1034
rect 5005 1846 5039 1880
rect 5005 1778 5039 1812
rect 5005 1710 5039 1744
rect 5005 1642 5039 1676
rect 5005 1574 5039 1608
rect 5005 1506 5039 1540
rect 5005 1438 5039 1472
rect 5005 1370 5039 1404
rect 5005 1302 5039 1336
rect 5005 1234 5039 1268
rect 5005 1166 5039 1200
rect 5005 1098 5039 1132
rect 5005 1030 5039 1064
rect 1801 932 1835 966
rect 5005 962 5039 996
rect 1945 864 1979 898
rect 2013 864 2047 898
rect 2081 864 2115 898
rect 2149 864 2183 898
rect 2217 864 2251 898
rect 2285 864 2319 898
rect 2353 864 2387 898
rect 2421 864 2455 898
rect 2489 864 2523 898
rect 2557 864 2591 898
rect 2625 864 2659 898
rect 2693 864 2727 898
rect 2761 864 2795 898
rect 2829 864 2863 898
rect 2897 864 2931 898
rect 2965 864 2999 898
rect 3033 864 3067 898
rect 3101 864 3135 898
rect 3169 864 3203 898
rect 3237 864 3271 898
rect 3305 864 3339 898
rect 3373 864 3407 898
rect 3441 864 3475 898
rect 3509 864 3543 898
rect 3577 864 3611 898
rect 3645 864 3679 898
rect 3713 864 3747 898
rect 3781 864 3815 898
rect 3849 864 3883 898
rect 3917 864 3951 898
rect 3985 864 4019 898
rect 4053 864 4087 898
rect 4121 864 4155 898
rect 4189 864 4223 898
rect 4257 864 4291 898
rect 4325 864 4359 898
rect 4393 864 4427 898
rect 4461 864 4495 898
rect 4529 864 4563 898
rect 4597 864 4631 898
rect 4665 864 4699 898
rect 4733 864 4767 898
rect 4801 864 4835 898
rect 4869 864 4903 898
rect 4937 864 4971 898
<< mvnsubdiffcont >>
rect 2039 39440 2073 39474
rect 1946 4080 2048 39406
rect 2107 39372 8465 39474
rect 8499 39320 8533 39354
rect 2208 9595 7546 9697
rect 7803 9536 8381 9638
rect 8431 9604 8533 39286
rect 8415 9536 8449 9570
rect 7735 9479 7769 9513
rect 1946 3417 2048 3927
rect 7735 4175 7837 9445
rect 2020 3349 2054 3383
rect 2088 3349 2598 3451
rect 2666 3349 7120 3451
rect 7235 3349 7677 3451
rect 7735 3417 7837 4063
rect 7711 3349 7745 3383
<< poly >>
rect 3023 38854 7729 38870
rect 3023 38820 3039 38854
rect 3073 38820 3108 38854
rect 3142 38820 3177 38854
rect 3211 38820 3246 38854
rect 3280 38820 3315 38854
rect 3349 38820 3384 38854
rect 3418 38820 3453 38854
rect 3487 38820 3522 38854
rect 3556 38820 3591 38854
rect 3625 38820 3660 38854
rect 3694 38820 3729 38854
rect 3763 38820 3798 38854
rect 3832 38820 3867 38854
rect 3901 38820 3936 38854
rect 3970 38820 4005 38854
rect 4039 38820 4074 38854
rect 4108 38820 4143 38854
rect 4177 38820 4211 38854
rect 4245 38820 4279 38854
rect 4313 38820 4347 38854
rect 4381 38820 4415 38854
rect 4449 38820 4483 38854
rect 4517 38820 4551 38854
rect 4585 38820 4619 38854
rect 4653 38820 4687 38854
rect 4721 38820 4755 38854
rect 4789 38820 4823 38854
rect 4857 38820 4891 38854
rect 4925 38820 4959 38854
rect 4993 38820 5027 38854
rect 5061 38820 5095 38854
rect 5129 38820 5163 38854
rect 5197 38820 5231 38854
rect 5265 38820 5299 38854
rect 5333 38820 5367 38854
rect 5401 38820 5435 38854
rect 5469 38820 5503 38854
rect 5537 38820 5571 38854
rect 5605 38820 5639 38854
rect 5673 38820 5707 38854
rect 5741 38820 5775 38854
rect 5809 38820 5843 38854
rect 5877 38820 5911 38854
rect 5945 38820 5979 38854
rect 6013 38820 6047 38854
rect 6081 38820 6115 38854
rect 6149 38820 6183 38854
rect 6217 38820 6251 38854
rect 6285 38820 6319 38854
rect 6353 38820 6387 38854
rect 6421 38820 6455 38854
rect 6489 38820 6523 38854
rect 6557 38820 6591 38854
rect 6625 38820 6659 38854
rect 6693 38820 6727 38854
rect 6761 38820 6795 38854
rect 6829 38820 6863 38854
rect 6897 38820 6931 38854
rect 6965 38820 6999 38854
rect 7033 38820 7067 38854
rect 7101 38820 7135 38854
rect 7169 38820 7203 38854
rect 7237 38820 7271 38854
rect 7305 38820 7339 38854
rect 7373 38820 7407 38854
rect 7441 38820 7475 38854
rect 7509 38820 7543 38854
rect 7577 38820 7611 38854
rect 7645 38820 7679 38854
rect 7713 38820 7729 38854
rect 3023 38804 7729 38820
rect 3023 37081 3059 37340
rect 3261 37081 3297 37340
rect 3577 37081 3613 37340
rect 3815 37081 3851 37340
rect 4131 37081 4167 37340
rect 4369 37081 4405 37340
rect 4685 37081 4721 37340
rect 4923 37081 4959 37340
rect 5239 37081 5275 37340
rect 5477 37081 5513 37340
rect 5793 37081 5829 37340
rect 6031 37081 6067 37340
rect 6347 37081 6383 37340
rect 6585 37081 6621 37340
rect 6901 37081 6937 37340
rect 7139 37081 7175 37340
rect 7455 37081 7491 37340
rect 7693 37081 7729 37340
rect 3023 37065 7729 37081
rect 3023 37031 3039 37065
rect 3073 37031 3108 37065
rect 3142 37031 3177 37065
rect 3211 37031 3246 37065
rect 3280 37031 3315 37065
rect 3349 37031 3384 37065
rect 3418 37031 3453 37065
rect 3487 37031 3522 37065
rect 3556 37031 3591 37065
rect 3625 37031 3660 37065
rect 3694 37031 3729 37065
rect 3763 37031 3798 37065
rect 3832 37031 3867 37065
rect 3901 37031 3936 37065
rect 3970 37031 4005 37065
rect 4039 37031 4074 37065
rect 4108 37031 4143 37065
rect 4177 37031 4211 37065
rect 4245 37031 4279 37065
rect 4313 37031 4347 37065
rect 4381 37031 4415 37065
rect 4449 37031 4483 37065
rect 4517 37031 4551 37065
rect 4585 37031 4619 37065
rect 4653 37031 4687 37065
rect 4721 37031 4755 37065
rect 4789 37031 4823 37065
rect 4857 37031 4891 37065
rect 4925 37031 4959 37065
rect 4993 37031 5027 37065
rect 5061 37031 5095 37065
rect 5129 37031 5163 37065
rect 5197 37031 5231 37065
rect 5265 37031 5299 37065
rect 5333 37031 5367 37065
rect 5401 37031 5435 37065
rect 5469 37031 5503 37065
rect 5537 37031 5571 37065
rect 5605 37031 5639 37065
rect 5673 37031 5707 37065
rect 5741 37031 5775 37065
rect 5809 37031 5843 37065
rect 5877 37031 5911 37065
rect 5945 37031 5979 37065
rect 6013 37031 6047 37065
rect 6081 37031 6115 37065
rect 6149 37031 6183 37065
rect 6217 37031 6251 37065
rect 6285 37031 6319 37065
rect 6353 37031 6387 37065
rect 6421 37031 6455 37065
rect 6489 37031 6523 37065
rect 6557 37031 6591 37065
rect 6625 37031 6659 37065
rect 6693 37031 6727 37065
rect 6761 37031 6795 37065
rect 6829 37031 6863 37065
rect 6897 37031 6931 37065
rect 6965 37031 6999 37065
rect 7033 37031 7067 37065
rect 7101 37031 7135 37065
rect 7169 37031 7203 37065
rect 7237 37031 7271 37065
rect 7305 37031 7339 37065
rect 7373 37031 7407 37065
rect 7441 37031 7475 37065
rect 7509 37031 7543 37065
rect 7577 37031 7611 37065
rect 7645 37031 7679 37065
rect 7713 37031 7729 37065
rect 3023 37015 7729 37031
rect 3023 36804 3059 37015
rect 3261 36804 3297 37015
rect 3577 36804 3613 37015
rect 3815 36804 3851 37015
rect 4131 36804 4167 37015
rect 4369 36804 4405 37015
rect 4685 36804 4721 37015
rect 4923 36804 4959 37015
rect 5239 36804 5275 37015
rect 5477 36804 5513 37015
rect 5793 36804 5829 37015
rect 6031 36804 6067 37015
rect 6347 36804 6383 37015
rect 6585 36804 6621 37015
rect 6901 36804 6937 37015
rect 7139 36804 7175 37015
rect 7455 36804 7491 37015
rect 7693 36804 7729 37015
rect 3023 35115 3059 35340
rect 3261 35115 3297 35340
rect 3577 35115 3613 35340
rect 3815 35115 3851 35340
rect 4131 35115 4167 35340
rect 4369 35115 4405 35340
rect 4685 35115 4721 35340
rect 4923 35115 4959 35340
rect 5239 35115 5275 35340
rect 5477 35115 5513 35340
rect 5793 35115 5829 35340
rect 6031 35115 6067 35340
rect 6347 35115 6383 35340
rect 6585 35115 6621 35340
rect 6901 35115 6937 35340
rect 7139 35115 7175 35340
rect 7455 35115 7491 35340
rect 7693 35115 7729 35340
rect 3023 35099 7729 35115
rect 3023 35065 3039 35099
rect 3073 35065 3108 35099
rect 3142 35065 3177 35099
rect 3211 35065 3246 35099
rect 3280 35065 3315 35099
rect 3349 35065 3384 35099
rect 3418 35065 3453 35099
rect 3487 35065 3522 35099
rect 3556 35065 3591 35099
rect 3625 35065 3660 35099
rect 3694 35065 3729 35099
rect 3763 35065 3798 35099
rect 3832 35065 3867 35099
rect 3901 35065 3936 35099
rect 3970 35065 4005 35099
rect 4039 35065 4074 35099
rect 4108 35065 4143 35099
rect 4177 35065 4211 35099
rect 4245 35065 4279 35099
rect 4313 35065 4347 35099
rect 4381 35065 4415 35099
rect 4449 35065 4483 35099
rect 4517 35065 4551 35099
rect 4585 35065 4619 35099
rect 4653 35065 4687 35099
rect 4721 35065 4755 35099
rect 4789 35065 4823 35099
rect 4857 35065 4891 35099
rect 4925 35065 4959 35099
rect 4993 35065 5027 35099
rect 5061 35065 5095 35099
rect 5129 35065 5163 35099
rect 5197 35065 5231 35099
rect 5265 35065 5299 35099
rect 5333 35065 5367 35099
rect 5401 35065 5435 35099
rect 5469 35065 5503 35099
rect 5537 35065 5571 35099
rect 5605 35065 5639 35099
rect 5673 35065 5707 35099
rect 5741 35065 5775 35099
rect 5809 35065 5843 35099
rect 5877 35065 5911 35099
rect 5945 35065 5979 35099
rect 6013 35065 6047 35099
rect 6081 35065 6115 35099
rect 6149 35065 6183 35099
rect 6217 35065 6251 35099
rect 6285 35065 6319 35099
rect 6353 35065 6387 35099
rect 6421 35065 6455 35099
rect 6489 35065 6523 35099
rect 6557 35065 6591 35099
rect 6625 35065 6659 35099
rect 6693 35065 6727 35099
rect 6761 35065 6795 35099
rect 6829 35065 6863 35099
rect 6897 35065 6931 35099
rect 6965 35065 6999 35099
rect 7033 35065 7067 35099
rect 7101 35065 7135 35099
rect 7169 35065 7203 35099
rect 7237 35065 7271 35099
rect 7305 35065 7339 35099
rect 7373 35065 7407 35099
rect 7441 35065 7475 35099
rect 7509 35065 7543 35099
rect 7577 35065 7611 35099
rect 7645 35065 7679 35099
rect 7713 35065 7729 35099
rect 3023 35049 7729 35065
rect 3023 34804 3059 35049
rect 3261 34804 3297 35049
rect 3577 34804 3613 35049
rect 3815 34804 3851 35049
rect 4131 34804 4167 35049
rect 4369 34804 4405 35049
rect 4685 34804 4721 35049
rect 4923 34804 4959 35049
rect 5239 34804 5275 35049
rect 5477 34804 5513 35049
rect 5793 34804 5829 35049
rect 6031 34804 6067 35049
rect 6347 34804 6383 35049
rect 6585 34804 6621 35049
rect 6901 34804 6937 35049
rect 7139 34804 7175 35049
rect 7455 34804 7491 35049
rect 7693 34804 7729 35049
rect 3023 33116 3059 33340
rect 3261 33116 3297 33340
rect 3577 33116 3613 33340
rect 3815 33116 3851 33340
rect 4131 33116 4167 33340
rect 4369 33116 4405 33340
rect 4685 33116 4721 33340
rect 4923 33116 4959 33340
rect 5239 33116 5275 33340
rect 5477 33116 5513 33340
rect 5793 33116 5829 33340
rect 6031 33116 6067 33340
rect 6347 33116 6383 33340
rect 6585 33116 6621 33340
rect 6901 33116 6937 33340
rect 7139 33116 7175 33340
rect 7455 33116 7491 33340
rect 7693 33116 7729 33340
rect 3023 33100 7729 33116
rect 3023 33066 3039 33100
rect 3073 33066 3108 33100
rect 3142 33066 3177 33100
rect 3211 33066 3246 33100
rect 3280 33066 3315 33100
rect 3349 33066 3384 33100
rect 3418 33066 3453 33100
rect 3487 33066 3522 33100
rect 3556 33066 3591 33100
rect 3625 33066 3660 33100
rect 3694 33066 3729 33100
rect 3763 33066 3798 33100
rect 3832 33066 3867 33100
rect 3901 33066 3936 33100
rect 3970 33066 4005 33100
rect 4039 33066 4074 33100
rect 4108 33066 4143 33100
rect 4177 33066 4211 33100
rect 4245 33066 4279 33100
rect 4313 33066 4347 33100
rect 4381 33066 4415 33100
rect 4449 33066 4483 33100
rect 4517 33066 4551 33100
rect 4585 33066 4619 33100
rect 4653 33066 4687 33100
rect 4721 33066 4755 33100
rect 4789 33066 4823 33100
rect 4857 33066 4891 33100
rect 4925 33066 4959 33100
rect 4993 33066 5027 33100
rect 5061 33066 5095 33100
rect 5129 33066 5163 33100
rect 5197 33066 5231 33100
rect 5265 33066 5299 33100
rect 5333 33066 5367 33100
rect 5401 33066 5435 33100
rect 5469 33066 5503 33100
rect 5537 33066 5571 33100
rect 5605 33066 5639 33100
rect 5673 33066 5707 33100
rect 5741 33066 5775 33100
rect 5809 33066 5843 33100
rect 5877 33066 5911 33100
rect 5945 33066 5979 33100
rect 6013 33066 6047 33100
rect 6081 33066 6115 33100
rect 6149 33066 6183 33100
rect 6217 33066 6251 33100
rect 6285 33066 6319 33100
rect 6353 33066 6387 33100
rect 6421 33066 6455 33100
rect 6489 33066 6523 33100
rect 6557 33066 6591 33100
rect 6625 33066 6659 33100
rect 6693 33066 6727 33100
rect 6761 33066 6795 33100
rect 6829 33066 6863 33100
rect 6897 33066 6931 33100
rect 6965 33066 6999 33100
rect 7033 33066 7067 33100
rect 7101 33066 7135 33100
rect 7169 33066 7203 33100
rect 7237 33066 7271 33100
rect 7305 33066 7339 33100
rect 7373 33066 7407 33100
rect 7441 33066 7475 33100
rect 7509 33066 7543 33100
rect 7577 33066 7611 33100
rect 7645 33066 7679 33100
rect 7713 33066 7729 33100
rect 3023 33050 7729 33066
rect 3023 32804 3059 33050
rect 3261 32804 3297 33050
rect 3577 32804 3613 33050
rect 3815 32804 3851 33050
rect 4131 32804 4167 33050
rect 4369 32804 4405 33050
rect 4685 32804 4721 33050
rect 4923 32804 4959 33050
rect 5239 32804 5275 33050
rect 5477 32804 5513 33050
rect 5793 32804 5829 33050
rect 6031 32804 6067 33050
rect 6347 32804 6383 33050
rect 6585 32804 6621 33050
rect 6901 32804 6937 33050
rect 7139 32804 7175 33050
rect 7455 32804 7491 33050
rect 7693 32804 7729 33050
rect 3023 31093 3059 31340
rect 3261 31093 3297 31340
rect 3577 31093 3613 31340
rect 3815 31093 3851 31340
rect 4131 31093 4167 31340
rect 4369 31093 4405 31340
rect 4685 31093 4721 31340
rect 4923 31093 4959 31340
rect 5239 31093 5275 31340
rect 5477 31093 5513 31340
rect 5793 31093 5829 31340
rect 6031 31093 6067 31340
rect 6347 31093 6383 31340
rect 6585 31093 6621 31340
rect 6901 31093 6937 31340
rect 7139 31093 7175 31340
rect 7455 31093 7491 31340
rect 7693 31093 7729 31340
rect 3023 31077 7729 31093
rect 3023 31043 3039 31077
rect 3073 31043 3108 31077
rect 3142 31043 3177 31077
rect 3211 31043 3246 31077
rect 3280 31043 3315 31077
rect 3349 31043 3384 31077
rect 3418 31043 3453 31077
rect 3487 31043 3522 31077
rect 3556 31043 3591 31077
rect 3625 31043 3660 31077
rect 3694 31043 3729 31077
rect 3763 31043 3798 31077
rect 3832 31043 3867 31077
rect 3901 31043 3936 31077
rect 3970 31043 4005 31077
rect 4039 31043 4074 31077
rect 4108 31043 4143 31077
rect 4177 31043 4211 31077
rect 4245 31043 4279 31077
rect 4313 31043 4347 31077
rect 4381 31043 4415 31077
rect 4449 31043 4483 31077
rect 4517 31043 4551 31077
rect 4585 31043 4619 31077
rect 4653 31043 4687 31077
rect 4721 31043 4755 31077
rect 4789 31043 4823 31077
rect 4857 31043 4891 31077
rect 4925 31043 4959 31077
rect 4993 31043 5027 31077
rect 5061 31043 5095 31077
rect 5129 31043 5163 31077
rect 5197 31043 5231 31077
rect 5265 31043 5299 31077
rect 5333 31043 5367 31077
rect 5401 31043 5435 31077
rect 5469 31043 5503 31077
rect 5537 31043 5571 31077
rect 5605 31043 5639 31077
rect 5673 31043 5707 31077
rect 5741 31043 5775 31077
rect 5809 31043 5843 31077
rect 5877 31043 5911 31077
rect 5945 31043 5979 31077
rect 6013 31043 6047 31077
rect 6081 31043 6115 31077
rect 6149 31043 6183 31077
rect 6217 31043 6251 31077
rect 6285 31043 6319 31077
rect 6353 31043 6387 31077
rect 6421 31043 6455 31077
rect 6489 31043 6523 31077
rect 6557 31043 6591 31077
rect 6625 31043 6659 31077
rect 6693 31043 6727 31077
rect 6761 31043 6795 31077
rect 6829 31043 6863 31077
rect 6897 31043 6931 31077
rect 6965 31043 6999 31077
rect 7033 31043 7067 31077
rect 7101 31043 7135 31077
rect 7169 31043 7203 31077
rect 7237 31043 7271 31077
rect 7305 31043 7339 31077
rect 7373 31043 7407 31077
rect 7441 31043 7475 31077
rect 7509 31043 7543 31077
rect 7577 31043 7611 31077
rect 7645 31043 7679 31077
rect 7713 31043 7729 31077
rect 3023 31027 7729 31043
rect 3023 30804 3059 31027
rect 3261 30804 3297 31027
rect 3577 30804 3613 31027
rect 3815 30804 3851 31027
rect 4131 30804 4167 31027
rect 4369 30804 4405 31027
rect 4685 30804 4721 31027
rect 4923 30804 4959 31027
rect 5239 30804 5275 31027
rect 5477 30804 5513 31027
rect 5793 30804 5829 31027
rect 6031 30804 6067 31027
rect 6347 30804 6383 31027
rect 6585 30804 6621 31027
rect 6901 30804 6937 31027
rect 7139 30804 7175 31027
rect 7455 30804 7491 31027
rect 7693 30804 7729 31027
rect 3023 29266 3059 29340
rect 3261 29266 3297 29340
rect 3577 29266 3613 29340
rect 3815 29266 3851 29340
rect 4131 29266 4167 29340
rect 4369 29266 4405 29340
rect 4685 29266 4721 29340
rect 4923 29266 4959 29340
rect 5239 29266 5275 29340
rect 5477 29266 5513 29340
rect 5793 29266 5829 29340
rect 6031 29266 6067 29340
rect 6347 29266 6383 29340
rect 6585 29266 6621 29340
rect 6901 29266 6937 29340
rect 7139 29266 7175 29340
rect 7455 29266 7491 29340
rect 7693 29266 7729 29340
rect 3023 29250 7729 29266
rect 3023 29216 3039 29250
rect 3073 29216 3108 29250
rect 3142 29216 3177 29250
rect 3211 29216 3246 29250
rect 3280 29216 3315 29250
rect 3349 29216 3384 29250
rect 3418 29216 3453 29250
rect 3487 29216 3522 29250
rect 3556 29216 3591 29250
rect 3625 29216 3660 29250
rect 3694 29216 3729 29250
rect 3763 29216 3798 29250
rect 3832 29216 3867 29250
rect 3901 29216 3936 29250
rect 3970 29216 4005 29250
rect 4039 29216 4074 29250
rect 4108 29216 4143 29250
rect 4177 29216 4211 29250
rect 4245 29216 4279 29250
rect 4313 29216 4347 29250
rect 4381 29216 4415 29250
rect 4449 29216 4483 29250
rect 4517 29216 4551 29250
rect 4585 29216 4619 29250
rect 4653 29216 4687 29250
rect 4721 29216 4755 29250
rect 4789 29216 4823 29250
rect 4857 29216 4891 29250
rect 4925 29216 4959 29250
rect 4993 29216 5027 29250
rect 5061 29216 5095 29250
rect 5129 29216 5163 29250
rect 5197 29216 5231 29250
rect 5265 29216 5299 29250
rect 5333 29216 5367 29250
rect 5401 29216 5435 29250
rect 5469 29216 5503 29250
rect 5537 29216 5571 29250
rect 5605 29216 5639 29250
rect 5673 29216 5707 29250
rect 5741 29216 5775 29250
rect 5809 29216 5843 29250
rect 5877 29216 5911 29250
rect 5945 29216 5979 29250
rect 6013 29216 6047 29250
rect 6081 29216 6115 29250
rect 6149 29216 6183 29250
rect 6217 29216 6251 29250
rect 6285 29216 6319 29250
rect 6353 29216 6387 29250
rect 6421 29216 6455 29250
rect 6489 29216 6523 29250
rect 6557 29216 6591 29250
rect 6625 29216 6659 29250
rect 6693 29216 6727 29250
rect 6761 29216 6795 29250
rect 6829 29216 6863 29250
rect 6897 29216 6931 29250
rect 6965 29216 6999 29250
rect 7033 29216 7067 29250
rect 7101 29216 7135 29250
rect 7169 29216 7203 29250
rect 7237 29216 7271 29250
rect 7305 29216 7339 29250
rect 7373 29216 7407 29250
rect 7441 29216 7475 29250
rect 7509 29216 7543 29250
rect 7577 29216 7611 29250
rect 7645 29216 7679 29250
rect 7713 29216 7729 29250
rect 3023 29200 7729 29216
rect 5239 28804 5275 29200
rect 5477 28804 5513 29200
rect 5793 28804 5829 29200
rect 6031 28804 6067 29200
rect 6347 28804 6383 29200
rect 6585 28804 6621 29200
rect 6901 28804 6937 29200
rect 7139 28804 7175 29200
rect 7455 28804 7491 29200
rect 7693 28804 7729 29200
rect 5239 27121 5275 27340
rect 5477 27121 5513 27340
rect 5793 27121 5829 27340
rect 6031 27121 6067 27340
rect 6347 27121 6383 27340
rect 6585 27121 6621 27340
rect 6901 27121 6937 27340
rect 7139 27121 7175 27340
rect 7455 27121 7491 27340
rect 7693 27121 7729 27340
rect 5239 27105 7729 27121
rect 5239 27071 5255 27105
rect 5289 27071 5325 27105
rect 5359 27071 5395 27105
rect 5429 27071 5465 27105
rect 5499 27071 5535 27105
rect 5569 27071 5605 27105
rect 5639 27071 5675 27105
rect 5709 27071 5745 27105
rect 5779 27071 5815 27105
rect 5849 27071 5885 27105
rect 5919 27071 5954 27105
rect 5988 27071 6023 27105
rect 6057 27071 6092 27105
rect 6126 27071 6161 27105
rect 6195 27071 6230 27105
rect 6264 27071 6299 27105
rect 6333 27071 6368 27105
rect 6402 27071 6437 27105
rect 6471 27071 6506 27105
rect 6540 27071 6575 27105
rect 6609 27071 6644 27105
rect 6678 27071 6713 27105
rect 6747 27071 6782 27105
rect 6816 27071 6851 27105
rect 6885 27071 6920 27105
rect 6954 27071 6989 27105
rect 7023 27071 7058 27105
rect 7092 27071 7127 27105
rect 7161 27071 7196 27105
rect 7230 27071 7265 27105
rect 7299 27071 7334 27105
rect 7368 27071 7403 27105
rect 7437 27071 7472 27105
rect 7506 27071 7541 27105
rect 7575 27071 7610 27105
rect 7644 27071 7679 27105
rect 7713 27071 7729 27105
rect 5239 27055 7729 27071
rect 5239 26804 5275 27055
rect 5477 26804 5513 27055
rect 5793 26804 5829 27055
rect 6031 26804 6067 27055
rect 6347 26804 6383 27055
rect 6585 26804 6621 27055
rect 6901 26804 6937 27055
rect 7139 26804 7175 27055
rect 7455 26804 7491 27055
rect 7693 26804 7729 27055
rect 5239 25128 5275 25340
rect 5477 25128 5513 25340
rect 5793 25128 5829 25340
rect 6031 25128 6067 25340
rect 6347 25128 6383 25340
rect 6585 25128 6621 25340
rect 6901 25128 6937 25340
rect 7139 25128 7175 25340
rect 7455 25128 7491 25340
rect 7693 25128 7729 25340
rect 5239 25112 7729 25128
rect 5239 25078 5255 25112
rect 5289 25078 5325 25112
rect 5359 25078 5395 25112
rect 5429 25078 5465 25112
rect 5499 25078 5535 25112
rect 5569 25078 5605 25112
rect 5639 25078 5675 25112
rect 5709 25078 5745 25112
rect 5779 25078 5815 25112
rect 5849 25078 5885 25112
rect 5919 25078 5954 25112
rect 5988 25078 6023 25112
rect 6057 25078 6092 25112
rect 6126 25078 6161 25112
rect 6195 25078 6230 25112
rect 6264 25078 6299 25112
rect 6333 25078 6368 25112
rect 6402 25078 6437 25112
rect 6471 25078 6506 25112
rect 6540 25078 6575 25112
rect 6609 25078 6644 25112
rect 6678 25078 6713 25112
rect 6747 25078 6782 25112
rect 6816 25078 6851 25112
rect 6885 25078 6920 25112
rect 6954 25078 6989 25112
rect 7023 25078 7058 25112
rect 7092 25078 7127 25112
rect 7161 25078 7196 25112
rect 7230 25078 7265 25112
rect 7299 25078 7334 25112
rect 7368 25078 7403 25112
rect 7437 25078 7472 25112
rect 7506 25078 7541 25112
rect 7575 25078 7610 25112
rect 7644 25078 7679 25112
rect 7713 25078 7729 25112
rect 5239 25062 7729 25078
rect 5239 24804 5275 25062
rect 5477 24804 5513 25062
rect 5793 24804 5829 25062
rect 6031 24804 6067 25062
rect 6347 24804 6383 25062
rect 6585 24804 6621 25062
rect 6901 24804 6937 25062
rect 7139 24804 7175 25062
rect 7455 24804 7491 25062
rect 7693 24804 7729 25062
rect 5239 23140 5275 23340
rect 5477 23140 5513 23340
rect 5793 23140 5829 23340
rect 6031 23140 6067 23340
rect 6347 23140 6383 23340
rect 6585 23140 6621 23340
rect 6901 23140 6937 23340
rect 7139 23140 7175 23340
rect 7455 23140 7491 23340
rect 7693 23140 7729 23340
rect 5239 23124 7729 23140
rect 5239 23090 5255 23124
rect 5289 23090 5325 23124
rect 5359 23090 5395 23124
rect 5429 23090 5465 23124
rect 5499 23090 5535 23124
rect 5569 23090 5605 23124
rect 5639 23090 5675 23124
rect 5709 23090 5745 23124
rect 5779 23090 5815 23124
rect 5849 23090 5885 23124
rect 5919 23090 5954 23124
rect 5988 23090 6023 23124
rect 6057 23090 6092 23124
rect 6126 23090 6161 23124
rect 6195 23090 6230 23124
rect 6264 23090 6299 23124
rect 6333 23090 6368 23124
rect 6402 23090 6437 23124
rect 6471 23090 6506 23124
rect 6540 23090 6575 23124
rect 6609 23090 6644 23124
rect 6678 23090 6713 23124
rect 6747 23090 6782 23124
rect 6816 23090 6851 23124
rect 6885 23090 6920 23124
rect 6954 23090 6989 23124
rect 7023 23090 7058 23124
rect 7092 23090 7127 23124
rect 7161 23090 7196 23124
rect 7230 23090 7265 23124
rect 7299 23090 7334 23124
rect 7368 23090 7403 23124
rect 7437 23090 7472 23124
rect 7506 23090 7541 23124
rect 7575 23090 7610 23124
rect 7644 23090 7679 23124
rect 7713 23090 7729 23124
rect 5239 23074 7729 23090
rect 5239 22804 5275 23074
rect 5477 22804 5513 23074
rect 5793 22804 5829 23074
rect 6031 22804 6067 23074
rect 6347 22804 6383 23074
rect 6585 22804 6621 23074
rect 6901 22804 6937 23074
rect 7139 22804 7175 23074
rect 7455 22804 7491 23074
rect 7693 22804 7729 23074
rect 5239 21099 5275 21340
rect 5477 21099 5513 21340
rect 5793 21099 5829 21340
rect 6031 21099 6067 21340
rect 6347 21099 6383 21340
rect 6585 21099 6621 21340
rect 6901 21099 6937 21340
rect 7139 21099 7175 21340
rect 7455 21099 7491 21340
rect 7693 21099 7729 21340
rect 5239 21083 7729 21099
rect 5239 21049 5255 21083
rect 5289 21049 5325 21083
rect 5359 21049 5395 21083
rect 5429 21049 5465 21083
rect 5499 21049 5535 21083
rect 5569 21049 5605 21083
rect 5639 21049 5675 21083
rect 5709 21049 5745 21083
rect 5779 21049 5815 21083
rect 5849 21049 5885 21083
rect 5919 21049 5954 21083
rect 5988 21049 6023 21083
rect 6057 21049 6092 21083
rect 6126 21049 6161 21083
rect 6195 21049 6230 21083
rect 6264 21049 6299 21083
rect 6333 21049 6368 21083
rect 6402 21049 6437 21083
rect 6471 21049 6506 21083
rect 6540 21049 6575 21083
rect 6609 21049 6644 21083
rect 6678 21049 6713 21083
rect 6747 21049 6782 21083
rect 6816 21049 6851 21083
rect 6885 21049 6920 21083
rect 6954 21049 6989 21083
rect 7023 21049 7058 21083
rect 7092 21049 7127 21083
rect 7161 21049 7196 21083
rect 7230 21049 7265 21083
rect 7299 21049 7334 21083
rect 7368 21049 7403 21083
rect 7437 21049 7472 21083
rect 7506 21049 7541 21083
rect 7575 21049 7610 21083
rect 7644 21049 7679 21083
rect 7713 21049 7729 21083
rect 5239 21033 7729 21049
rect 5239 20804 5275 21033
rect 5477 20804 5513 21033
rect 5793 20804 5829 21033
rect 6031 20804 6067 21033
rect 6347 20804 6383 21033
rect 6585 20804 6621 21033
rect 6901 20804 6937 21033
rect 7139 20804 7175 21033
rect 7455 20804 7491 21033
rect 7693 20804 7729 21033
rect 5239 19135 5275 19340
rect 5477 19135 5513 19340
rect 5793 19135 5829 19340
rect 6031 19135 6067 19340
rect 6347 19135 6383 19340
rect 6585 19135 6621 19340
rect 6901 19135 6937 19340
rect 7139 19135 7175 19340
rect 7455 19135 7491 19340
rect 7693 19135 7729 19340
rect 5239 19119 7729 19135
rect 5239 19085 5255 19119
rect 5289 19085 5325 19119
rect 5359 19085 5395 19119
rect 5429 19085 5465 19119
rect 5499 19085 5535 19119
rect 5569 19085 5605 19119
rect 5639 19085 5675 19119
rect 5709 19085 5745 19119
rect 5779 19085 5815 19119
rect 5849 19085 5885 19119
rect 5919 19085 5954 19119
rect 5988 19085 6023 19119
rect 6057 19085 6092 19119
rect 6126 19085 6161 19119
rect 6195 19085 6230 19119
rect 6264 19085 6299 19119
rect 6333 19085 6368 19119
rect 6402 19085 6437 19119
rect 6471 19085 6506 19119
rect 6540 19085 6575 19119
rect 6609 19085 6644 19119
rect 6678 19085 6713 19119
rect 6747 19085 6782 19119
rect 6816 19085 6851 19119
rect 6885 19085 6920 19119
rect 6954 19085 6989 19119
rect 7023 19085 7058 19119
rect 7092 19085 7127 19119
rect 7161 19085 7196 19119
rect 7230 19085 7265 19119
rect 7299 19085 7334 19119
rect 7368 19085 7403 19119
rect 7437 19085 7472 19119
rect 7506 19085 7541 19119
rect 7575 19085 7610 19119
rect 7644 19085 7679 19119
rect 7713 19085 7729 19119
rect 5239 19069 7729 19085
rect 5239 18804 5275 19069
rect 5477 18804 5513 19069
rect 5793 18804 5829 19069
rect 6031 18804 6067 19069
rect 6347 18804 6383 19069
rect 6585 18804 6621 19069
rect 6901 18804 6937 19069
rect 7139 18804 7175 19069
rect 7455 18804 7491 19069
rect 7693 18804 7729 19069
rect 5239 17261 5275 17340
rect 5477 17261 5513 17340
rect 5793 17261 5829 17340
rect 6031 17261 6067 17340
rect 6347 17261 6383 17340
rect 6585 17261 6621 17340
rect 6901 17261 6937 17340
rect 7139 17261 7175 17340
rect 7455 17261 7491 17340
rect 7693 17261 7729 17340
rect 5239 17245 7729 17261
rect 5239 17211 5255 17245
rect 5289 17211 5325 17245
rect 5359 17211 5395 17245
rect 5429 17211 5465 17245
rect 5499 17211 5535 17245
rect 5569 17211 5605 17245
rect 5639 17211 5675 17245
rect 5709 17211 5745 17245
rect 5779 17211 5815 17245
rect 5849 17211 5885 17245
rect 5919 17211 5954 17245
rect 5988 17211 6023 17245
rect 6057 17211 6092 17245
rect 6126 17211 6161 17245
rect 6195 17211 6230 17245
rect 6264 17211 6299 17245
rect 6333 17211 6368 17245
rect 6402 17211 6437 17245
rect 6471 17211 6506 17245
rect 6540 17211 6575 17245
rect 6609 17211 6644 17245
rect 6678 17211 6713 17245
rect 6747 17211 6782 17245
rect 6816 17211 6851 17245
rect 6885 17211 6920 17245
rect 6954 17211 6989 17245
rect 7023 17211 7058 17245
rect 7092 17211 7127 17245
rect 7161 17211 7196 17245
rect 7230 17211 7265 17245
rect 7299 17211 7334 17245
rect 7368 17211 7403 17245
rect 7437 17211 7472 17245
rect 7506 17211 7541 17245
rect 7575 17211 7610 17245
rect 7644 17211 7679 17245
rect 7713 17211 7729 17245
rect 5239 17195 7729 17211
rect 3023 15586 7729 15602
rect 3023 15552 3039 15586
rect 3073 15552 3108 15586
rect 3142 15552 3177 15586
rect 3211 15552 3246 15586
rect 3280 15552 3315 15586
rect 3349 15552 3384 15586
rect 3418 15552 3453 15586
rect 3487 15552 3522 15586
rect 3556 15552 3591 15586
rect 3625 15552 3660 15586
rect 3694 15552 3729 15586
rect 3763 15552 3798 15586
rect 3832 15552 3867 15586
rect 3901 15552 3936 15586
rect 3970 15552 4005 15586
rect 4039 15552 4074 15586
rect 4108 15552 4143 15586
rect 4177 15552 4211 15586
rect 4245 15552 4279 15586
rect 4313 15552 4347 15586
rect 4381 15552 4415 15586
rect 4449 15552 4483 15586
rect 4517 15552 4551 15586
rect 4585 15552 4619 15586
rect 4653 15552 4687 15586
rect 4721 15552 4755 15586
rect 4789 15552 4823 15586
rect 4857 15552 4891 15586
rect 4925 15552 4959 15586
rect 4993 15552 5027 15586
rect 5061 15552 5095 15586
rect 5129 15552 5163 15586
rect 5197 15552 5231 15586
rect 5265 15552 5299 15586
rect 5333 15552 5367 15586
rect 5401 15552 5435 15586
rect 5469 15552 5503 15586
rect 5537 15552 5571 15586
rect 5605 15552 5639 15586
rect 5673 15552 5707 15586
rect 5741 15552 5775 15586
rect 5809 15552 5843 15586
rect 5877 15552 5911 15586
rect 5945 15552 5979 15586
rect 6013 15552 6047 15586
rect 6081 15552 6115 15586
rect 6149 15552 6183 15586
rect 6217 15552 6251 15586
rect 6285 15552 6319 15586
rect 6353 15552 6387 15586
rect 6421 15552 6455 15586
rect 6489 15552 6523 15586
rect 6557 15552 6591 15586
rect 6625 15552 6659 15586
rect 6693 15552 6727 15586
rect 6761 15552 6795 15586
rect 6829 15552 6863 15586
rect 6897 15552 6931 15586
rect 6965 15552 6999 15586
rect 7033 15552 7067 15586
rect 7101 15552 7135 15586
rect 7169 15552 7203 15586
rect 7237 15552 7271 15586
rect 7305 15552 7339 15586
rect 7373 15552 7407 15586
rect 7441 15552 7475 15586
rect 7509 15552 7543 15586
rect 7577 15552 7611 15586
rect 7645 15552 7679 15586
rect 7713 15552 7729 15586
rect 3023 15536 7729 15552
rect 3023 13872 3059 14072
rect 3261 13872 3297 14072
rect 3577 13872 3613 14072
rect 3815 13872 3851 14072
rect 4131 13872 4167 14072
rect 4369 13872 4405 14072
rect 4685 13872 4721 14072
rect 4923 13872 4959 14072
rect 5239 13872 5275 14072
rect 5477 13872 5513 14072
rect 5793 13872 5829 14072
rect 6031 13872 6067 14072
rect 6347 13872 6383 14072
rect 6585 13872 6621 14072
rect 6901 13872 6937 14072
rect 7139 13872 7175 14072
rect 7455 13872 7491 14072
rect 7693 13872 7729 14072
rect 3023 13856 7729 13872
rect 3023 13822 3039 13856
rect 3073 13822 3108 13856
rect 3142 13822 3177 13856
rect 3211 13822 3246 13856
rect 3280 13822 3315 13856
rect 3349 13822 3384 13856
rect 3418 13822 3453 13856
rect 3487 13822 3522 13856
rect 3556 13822 3591 13856
rect 3625 13822 3660 13856
rect 3694 13822 3729 13856
rect 3763 13822 3798 13856
rect 3832 13822 3867 13856
rect 3901 13822 3936 13856
rect 3970 13822 4005 13856
rect 4039 13822 4073 13856
rect 4107 13822 4141 13856
rect 4175 13822 4209 13856
rect 4243 13822 4277 13856
rect 4311 13822 4345 13856
rect 4379 13822 4413 13856
rect 4447 13822 4481 13856
rect 4515 13822 4549 13856
rect 4583 13822 4617 13856
rect 4651 13822 4685 13856
rect 4719 13822 4753 13856
rect 4787 13822 4821 13856
rect 4855 13822 4889 13856
rect 4923 13822 4957 13856
rect 4991 13822 5025 13856
rect 5059 13822 5093 13856
rect 5127 13822 5161 13856
rect 5195 13822 5229 13856
rect 5263 13822 5297 13856
rect 5331 13822 5365 13856
rect 5399 13822 5433 13856
rect 5467 13822 5501 13856
rect 5535 13822 5569 13856
rect 5603 13822 5637 13856
rect 5671 13822 5705 13856
rect 5739 13822 5773 13856
rect 5807 13822 5841 13856
rect 5875 13822 5909 13856
rect 5943 13822 5977 13856
rect 6011 13822 6045 13856
rect 6079 13822 6113 13856
rect 6147 13822 6181 13856
rect 6215 13822 6249 13856
rect 6283 13822 6317 13856
rect 6351 13822 6385 13856
rect 6419 13822 6453 13856
rect 6487 13822 6521 13856
rect 6555 13822 6589 13856
rect 6623 13822 6657 13856
rect 6691 13822 6725 13856
rect 6759 13822 6793 13856
rect 6827 13822 6861 13856
rect 6895 13822 6929 13856
rect 6963 13822 6997 13856
rect 7031 13822 7065 13856
rect 7099 13822 7133 13856
rect 7167 13822 7201 13856
rect 7235 13822 7269 13856
rect 7303 13822 7337 13856
rect 7371 13822 7405 13856
rect 7439 13822 7473 13856
rect 7507 13822 7541 13856
rect 7575 13822 7609 13856
rect 7643 13822 7677 13856
rect 7711 13822 7729 13856
rect 3023 13806 7729 13822
rect 3023 13536 3059 13806
rect 3261 13536 3297 13806
rect 3577 13536 3613 13806
rect 3815 13536 3851 13806
rect 4131 13536 4167 13806
rect 4369 13536 4405 13806
rect 4685 13536 4721 13806
rect 4923 13536 4959 13806
rect 5239 13536 5275 13806
rect 5477 13536 5513 13806
rect 5793 13536 5829 13806
rect 6031 13536 6067 13806
rect 6347 13536 6383 13806
rect 6585 13536 6621 13806
rect 6901 13536 6937 13806
rect 7139 13536 7175 13806
rect 7455 13536 7491 13806
rect 7693 13536 7729 13806
rect 3023 11834 3059 12072
rect 3261 11834 3297 12072
rect 3577 11834 3613 12072
rect 3815 11834 3851 12072
rect 4131 11834 4167 12072
rect 4369 11834 4405 12072
rect 4685 11834 4721 12072
rect 4923 11834 4959 12072
rect 5239 11834 5275 12072
rect 5477 11834 5513 12072
rect 5793 11834 5829 12072
rect 6031 11834 6067 12072
rect 6347 11834 6383 12072
rect 6585 11834 6621 12072
rect 6901 11834 6937 12072
rect 7139 11834 7175 12072
rect 7455 11834 7491 12072
rect 7693 11834 7729 12072
rect 3023 11818 7729 11834
rect 3023 11784 3039 11818
rect 3073 11784 3108 11818
rect 3142 11784 3177 11818
rect 3211 11784 3246 11818
rect 3280 11784 3315 11818
rect 3349 11784 3384 11818
rect 3418 11784 3453 11818
rect 3487 11784 3522 11818
rect 3556 11784 3591 11818
rect 3625 11784 3660 11818
rect 3694 11784 3729 11818
rect 3763 11784 3798 11818
rect 3832 11784 3867 11818
rect 3901 11784 3936 11818
rect 3970 11784 4005 11818
rect 4039 11784 4073 11818
rect 4107 11784 4141 11818
rect 4175 11784 4209 11818
rect 4243 11784 4277 11818
rect 4311 11784 4345 11818
rect 4379 11784 4413 11818
rect 4447 11784 4481 11818
rect 4515 11784 4549 11818
rect 4583 11784 4617 11818
rect 4651 11784 4685 11818
rect 4719 11784 4753 11818
rect 4787 11784 4821 11818
rect 4855 11784 4889 11818
rect 4923 11784 4957 11818
rect 4991 11784 5025 11818
rect 5059 11784 5093 11818
rect 5127 11784 5161 11818
rect 5195 11784 5229 11818
rect 5263 11784 5297 11818
rect 5331 11784 5365 11818
rect 5399 11784 5433 11818
rect 5467 11784 5501 11818
rect 5535 11784 5569 11818
rect 5603 11784 5637 11818
rect 5671 11784 5705 11818
rect 5739 11784 5773 11818
rect 5807 11784 5841 11818
rect 5875 11784 5909 11818
rect 5943 11784 5977 11818
rect 6011 11784 6045 11818
rect 6079 11784 6113 11818
rect 6147 11784 6181 11818
rect 6215 11784 6249 11818
rect 6283 11784 6317 11818
rect 6351 11784 6385 11818
rect 6419 11784 6453 11818
rect 6487 11784 6521 11818
rect 6555 11784 6589 11818
rect 6623 11784 6657 11818
rect 6691 11784 6725 11818
rect 6759 11784 6793 11818
rect 6827 11784 6861 11818
rect 6895 11784 6929 11818
rect 6963 11784 6997 11818
rect 7031 11784 7065 11818
rect 7099 11784 7133 11818
rect 7167 11784 7201 11818
rect 7235 11784 7269 11818
rect 7303 11784 7337 11818
rect 7371 11784 7405 11818
rect 7439 11784 7473 11818
rect 7507 11784 7541 11818
rect 7575 11784 7609 11818
rect 7643 11784 7677 11818
rect 7711 11784 7729 11818
rect 3023 11768 7729 11784
rect 3023 11536 3059 11768
rect 3261 11536 3297 11768
rect 3577 11536 3613 11768
rect 3815 11536 3851 11768
rect 4131 11536 4167 11768
rect 4369 11536 4405 11768
rect 4685 11536 4721 11768
rect 4923 11536 4959 11768
rect 5239 11536 5275 11768
rect 5477 11536 5513 11768
rect 5793 11536 5829 11768
rect 6031 11536 6067 11768
rect 6347 11536 6383 11768
rect 6585 11536 6621 11768
rect 6901 11536 6937 11768
rect 7139 11536 7175 11768
rect 7455 11536 7491 11768
rect 7693 11536 7729 11768
rect 3023 10056 7729 10072
rect 3023 10022 3039 10056
rect 3073 10022 3108 10056
rect 3142 10022 3177 10056
rect 3211 10022 3246 10056
rect 3280 10022 3315 10056
rect 3349 10022 3384 10056
rect 3418 10022 3453 10056
rect 3487 10022 3522 10056
rect 3556 10022 3591 10056
rect 3625 10022 3660 10056
rect 3694 10022 3729 10056
rect 3763 10022 3798 10056
rect 3832 10022 3867 10056
rect 3901 10022 3936 10056
rect 3970 10022 4005 10056
rect 4039 10022 4074 10056
rect 4108 10022 4143 10056
rect 4177 10022 4211 10056
rect 4245 10022 4279 10056
rect 4313 10022 4347 10056
rect 4381 10022 4415 10056
rect 4449 10022 4483 10056
rect 4517 10022 4551 10056
rect 4585 10022 4619 10056
rect 4653 10022 4687 10056
rect 4721 10022 4755 10056
rect 4789 10022 4823 10056
rect 4857 10022 4891 10056
rect 4925 10022 4959 10056
rect 4993 10022 5027 10056
rect 5061 10022 5095 10056
rect 5129 10022 5163 10056
rect 5197 10022 5231 10056
rect 5265 10022 5299 10056
rect 5333 10022 5367 10056
rect 5401 10022 5435 10056
rect 5469 10022 5503 10056
rect 5537 10022 5571 10056
rect 5605 10022 5639 10056
rect 5673 10022 5707 10056
rect 5741 10022 5775 10056
rect 5809 10022 5843 10056
rect 5877 10022 5911 10056
rect 5945 10022 5979 10056
rect 6013 10022 6047 10056
rect 6081 10022 6115 10056
rect 6149 10022 6183 10056
rect 6217 10022 6251 10056
rect 6285 10022 6319 10056
rect 6353 10022 6387 10056
rect 6421 10022 6455 10056
rect 6489 10022 6523 10056
rect 6557 10022 6591 10056
rect 6625 10022 6659 10056
rect 6693 10022 6727 10056
rect 6761 10022 6795 10056
rect 6829 10022 6863 10056
rect 6897 10022 6931 10056
rect 6965 10022 6999 10056
rect 7033 10022 7067 10056
rect 7101 10022 7135 10056
rect 7169 10022 7203 10056
rect 7237 10022 7271 10056
rect 7305 10022 7339 10056
rect 7373 10022 7407 10056
rect 7441 10022 7475 10056
rect 7509 10022 7543 10056
rect 7577 10022 7611 10056
rect 7645 10022 7679 10056
rect 7713 10022 7729 10056
rect 3023 10006 7729 10022
rect 2468 9340 7380 9356
rect 2468 9306 2488 9340
rect 2522 9306 2556 9340
rect 2590 9306 2624 9340
rect 2658 9306 2692 9340
rect 2726 9306 2760 9340
rect 2794 9306 2828 9340
rect 2862 9306 2896 9340
rect 2930 9306 2964 9340
rect 2998 9306 3032 9340
rect 3066 9306 3100 9340
rect 3134 9306 3168 9340
rect 3202 9306 3236 9340
rect 3270 9306 3304 9340
rect 3338 9306 3372 9340
rect 3406 9306 3440 9340
rect 3474 9306 3508 9340
rect 3542 9306 3576 9340
rect 3610 9306 3644 9340
rect 3678 9306 3712 9340
rect 3746 9306 3780 9340
rect 3814 9306 3848 9340
rect 3882 9306 3916 9340
rect 3950 9306 3984 9340
rect 4018 9306 4052 9340
rect 4086 9306 4120 9340
rect 4154 9306 4188 9340
rect 4222 9306 4256 9340
rect 4290 9306 4324 9340
rect 4358 9306 4392 9340
rect 4426 9306 4460 9340
rect 4494 9306 4528 9340
rect 4562 9306 4596 9340
rect 4630 9306 4664 9340
rect 4698 9306 4732 9340
rect 4766 9306 4800 9340
rect 4834 9306 4868 9340
rect 4902 9306 4936 9340
rect 4970 9306 5004 9340
rect 5038 9306 5072 9340
rect 5106 9306 5140 9340
rect 5174 9306 5208 9340
rect 5242 9306 5276 9340
rect 5310 9306 5344 9340
rect 5378 9306 5412 9340
rect 5446 9306 5480 9340
rect 5514 9306 5548 9340
rect 5582 9306 5616 9340
rect 5650 9306 5684 9340
rect 5718 9306 5752 9340
rect 5786 9306 5820 9340
rect 5854 9306 5888 9340
rect 5922 9306 5956 9340
rect 5990 9306 6024 9340
rect 6058 9306 6092 9340
rect 6126 9306 6160 9340
rect 6194 9306 6228 9340
rect 6262 9306 6296 9340
rect 6330 9306 6364 9340
rect 6398 9306 6432 9340
rect 6466 9306 6500 9340
rect 6534 9306 6568 9340
rect 6602 9306 6636 9340
rect 6670 9306 6704 9340
rect 6738 9306 6772 9340
rect 6806 9306 6840 9340
rect 6874 9306 6908 9340
rect 6942 9306 6976 9340
rect 7010 9306 7044 9340
rect 7078 9306 7112 9340
rect 7146 9306 7180 9340
rect 7214 9306 7248 9340
rect 7282 9306 7316 9340
rect 7350 9306 7380 9340
rect 2468 9290 7380 9306
rect 2468 7540 7380 7556
rect 2468 7506 2488 7540
rect 2522 7506 2556 7540
rect 2590 7506 2624 7540
rect 2658 7506 2692 7540
rect 2726 7506 2760 7540
rect 2794 7506 2828 7540
rect 2862 7506 2896 7540
rect 2930 7506 2964 7540
rect 2998 7506 3032 7540
rect 3066 7506 3100 7540
rect 3134 7506 3168 7540
rect 3202 7506 3236 7540
rect 3270 7506 3304 7540
rect 3338 7506 3372 7540
rect 3406 7506 3440 7540
rect 3474 7506 3508 7540
rect 3542 7506 3576 7540
rect 3610 7506 3644 7540
rect 3678 7506 3712 7540
rect 3746 7506 3780 7540
rect 3814 7506 3848 7540
rect 3882 7506 3916 7540
rect 3950 7506 3984 7540
rect 4018 7506 4052 7540
rect 4086 7506 4120 7540
rect 4154 7506 4188 7540
rect 4222 7506 4256 7540
rect 4290 7506 4324 7540
rect 4358 7506 4392 7540
rect 4426 7506 4460 7540
rect 4494 7506 4528 7540
rect 4562 7506 4596 7540
rect 4630 7506 4664 7540
rect 4698 7506 4732 7540
rect 4766 7506 4800 7540
rect 4834 7506 4868 7540
rect 4902 7506 4936 7540
rect 4970 7506 5004 7540
rect 5038 7506 5072 7540
rect 5106 7506 5140 7540
rect 5174 7506 5208 7540
rect 5242 7506 5276 7540
rect 5310 7506 5344 7540
rect 5378 7506 5412 7540
rect 5446 7506 5480 7540
rect 5514 7506 5548 7540
rect 5582 7506 5616 7540
rect 5650 7506 5684 7540
rect 5718 7506 5752 7540
rect 5786 7506 5820 7540
rect 5854 7506 5888 7540
rect 5922 7506 5956 7540
rect 5990 7506 6024 7540
rect 6058 7506 6092 7540
rect 6126 7506 6160 7540
rect 6194 7506 6228 7540
rect 6262 7506 6296 7540
rect 6330 7506 6364 7540
rect 6398 7506 6432 7540
rect 6466 7506 6500 7540
rect 6534 7506 6568 7540
rect 6602 7506 6636 7540
rect 6670 7506 6704 7540
rect 6738 7506 6772 7540
rect 6806 7506 6840 7540
rect 6874 7506 6908 7540
rect 6942 7506 6976 7540
rect 7010 7506 7044 7540
rect 7078 7506 7112 7540
rect 7146 7506 7180 7540
rect 7214 7506 7248 7540
rect 7282 7506 7316 7540
rect 7350 7506 7380 7540
rect 2468 7490 7380 7506
rect 2640 5645 7048 5661
rect 2640 5611 2660 5645
rect 2694 5611 2728 5645
rect 2762 5611 2796 5645
rect 2830 5611 2864 5645
rect 2898 5611 2932 5645
rect 2966 5611 3000 5645
rect 3034 5611 3068 5645
rect 3102 5611 3136 5645
rect 3170 5611 3204 5645
rect 3238 5611 3272 5645
rect 3306 5611 3340 5645
rect 3374 5611 3408 5645
rect 3442 5611 3476 5645
rect 3510 5611 3544 5645
rect 3578 5611 3612 5645
rect 3646 5611 3680 5645
rect 3714 5611 3748 5645
rect 3782 5611 3816 5645
rect 3850 5611 3884 5645
rect 3918 5611 3952 5645
rect 3986 5611 4020 5645
rect 4054 5611 4088 5645
rect 4122 5611 4156 5645
rect 4190 5611 4224 5645
rect 4258 5611 4292 5645
rect 4326 5611 4360 5645
rect 4394 5611 4428 5645
rect 4462 5611 4496 5645
rect 4530 5611 4564 5645
rect 4598 5611 4632 5645
rect 4666 5611 4700 5645
rect 4734 5611 4768 5645
rect 4802 5611 4836 5645
rect 4870 5611 4904 5645
rect 4938 5611 4972 5645
rect 5006 5611 5040 5645
rect 5074 5611 5108 5645
rect 5142 5611 5176 5645
rect 5210 5611 5244 5645
rect 5278 5611 5312 5645
rect 5346 5611 5380 5645
rect 5414 5611 5448 5645
rect 5482 5611 5516 5645
rect 5550 5611 5584 5645
rect 5618 5611 5652 5645
rect 5686 5611 5720 5645
rect 5754 5611 5788 5645
rect 5822 5611 5856 5645
rect 5890 5611 5924 5645
rect 5958 5611 5992 5645
rect 6026 5611 6060 5645
rect 6094 5611 6128 5645
rect 6162 5611 6196 5645
rect 6230 5611 6264 5645
rect 6298 5611 6332 5645
rect 6366 5611 6400 5645
rect 6434 5611 6468 5645
rect 6502 5611 6536 5645
rect 6570 5611 6604 5645
rect 6638 5611 6672 5645
rect 6706 5611 6740 5645
rect 6774 5611 6808 5645
rect 6842 5611 6876 5645
rect 6910 5611 6944 5645
rect 6978 5611 7048 5645
rect 2640 5595 7048 5611
rect 1903 1856 1969 1872
rect 1903 1822 1919 1856
rect 1953 1822 1969 1856
rect 1903 1784 1969 1822
rect 1903 1750 1919 1784
rect 1953 1750 1969 1784
rect 1903 1712 1969 1750
rect 1903 1678 1919 1712
rect 1953 1678 1969 1712
rect 1903 1640 1969 1678
rect 1903 1606 1919 1640
rect 1953 1606 1969 1640
rect 1903 1568 1969 1606
rect 1903 1534 1919 1568
rect 1953 1534 1969 1568
rect 1903 1496 1969 1534
rect 1903 1462 1919 1496
rect 1953 1462 1969 1496
rect 1903 1423 1969 1462
rect 1903 1389 1919 1423
rect 1953 1389 1969 1423
rect 1903 1350 1969 1389
rect 1903 1316 1919 1350
rect 1953 1316 1969 1350
rect 1903 1277 1969 1316
rect 1903 1243 1919 1277
rect 1953 1243 1969 1277
rect 1903 1204 1969 1243
rect 1903 1170 1919 1204
rect 1953 1170 1969 1204
rect 1903 1131 1969 1170
rect 1903 1097 1919 1131
rect 1953 1097 1969 1131
rect 1903 1058 1969 1097
rect 1903 1024 1919 1058
rect 1953 1024 1969 1058
rect 1903 1008 1969 1024
rect 3433 1856 3499 1872
rect 3433 1822 3449 1856
rect 3483 1822 3499 1856
rect 3433 1784 3499 1822
rect 3433 1750 3449 1784
rect 3483 1750 3499 1784
rect 3433 1712 3499 1750
rect 3433 1678 3449 1712
rect 3483 1678 3499 1712
rect 3433 1640 3499 1678
rect 3433 1606 3449 1640
rect 3483 1606 3499 1640
rect 3433 1568 3499 1606
rect 3433 1534 3449 1568
rect 3483 1534 3499 1568
rect 3433 1496 3499 1534
rect 3433 1462 3449 1496
rect 3483 1462 3499 1496
rect 3433 1423 3499 1462
rect 3433 1389 3449 1423
rect 3483 1389 3499 1423
rect 3433 1350 3499 1389
rect 3433 1316 3449 1350
rect 3483 1316 3499 1350
rect 3433 1277 3499 1316
rect 3433 1243 3449 1277
rect 3483 1243 3499 1277
rect 3433 1204 3499 1243
rect 3433 1170 3449 1204
rect 3483 1170 3499 1204
rect 3433 1131 3499 1170
rect 3433 1097 3449 1131
rect 3483 1097 3499 1131
rect 3433 1058 3499 1097
rect 3433 1024 3449 1058
rect 3483 1024 3499 1058
rect 3433 1008 3499 1024
rect 154 221 220 244
rect 154 187 170 221
rect 204 187 220 221
rect 154 153 220 187
rect 154 119 170 153
rect 204 119 220 153
rect 154 103 220 119
rect 1612 221 1678 244
rect 1612 187 1628 221
rect 1662 187 1678 221
rect 1612 153 1678 187
rect 1612 119 1628 153
rect 1662 119 1678 153
rect 1612 103 1678 119
<< polycont >>
rect 3039 38820 3073 38854
rect 3108 38820 3142 38854
rect 3177 38820 3211 38854
rect 3246 38820 3280 38854
rect 3315 38820 3349 38854
rect 3384 38820 3418 38854
rect 3453 38820 3487 38854
rect 3522 38820 3556 38854
rect 3591 38820 3625 38854
rect 3660 38820 3694 38854
rect 3729 38820 3763 38854
rect 3798 38820 3832 38854
rect 3867 38820 3901 38854
rect 3936 38820 3970 38854
rect 4005 38820 4039 38854
rect 4074 38820 4108 38854
rect 4143 38820 4177 38854
rect 4211 38820 4245 38854
rect 4279 38820 4313 38854
rect 4347 38820 4381 38854
rect 4415 38820 4449 38854
rect 4483 38820 4517 38854
rect 4551 38820 4585 38854
rect 4619 38820 4653 38854
rect 4687 38820 4721 38854
rect 4755 38820 4789 38854
rect 4823 38820 4857 38854
rect 4891 38820 4925 38854
rect 4959 38820 4993 38854
rect 5027 38820 5061 38854
rect 5095 38820 5129 38854
rect 5163 38820 5197 38854
rect 5231 38820 5265 38854
rect 5299 38820 5333 38854
rect 5367 38820 5401 38854
rect 5435 38820 5469 38854
rect 5503 38820 5537 38854
rect 5571 38820 5605 38854
rect 5639 38820 5673 38854
rect 5707 38820 5741 38854
rect 5775 38820 5809 38854
rect 5843 38820 5877 38854
rect 5911 38820 5945 38854
rect 5979 38820 6013 38854
rect 6047 38820 6081 38854
rect 6115 38820 6149 38854
rect 6183 38820 6217 38854
rect 6251 38820 6285 38854
rect 6319 38820 6353 38854
rect 6387 38820 6421 38854
rect 6455 38820 6489 38854
rect 6523 38820 6557 38854
rect 6591 38820 6625 38854
rect 6659 38820 6693 38854
rect 6727 38820 6761 38854
rect 6795 38820 6829 38854
rect 6863 38820 6897 38854
rect 6931 38820 6965 38854
rect 6999 38820 7033 38854
rect 7067 38820 7101 38854
rect 7135 38820 7169 38854
rect 7203 38820 7237 38854
rect 7271 38820 7305 38854
rect 7339 38820 7373 38854
rect 7407 38820 7441 38854
rect 7475 38820 7509 38854
rect 7543 38820 7577 38854
rect 7611 38820 7645 38854
rect 7679 38820 7713 38854
rect 3039 37031 3073 37065
rect 3108 37031 3142 37065
rect 3177 37031 3211 37065
rect 3246 37031 3280 37065
rect 3315 37031 3349 37065
rect 3384 37031 3418 37065
rect 3453 37031 3487 37065
rect 3522 37031 3556 37065
rect 3591 37031 3625 37065
rect 3660 37031 3694 37065
rect 3729 37031 3763 37065
rect 3798 37031 3832 37065
rect 3867 37031 3901 37065
rect 3936 37031 3970 37065
rect 4005 37031 4039 37065
rect 4074 37031 4108 37065
rect 4143 37031 4177 37065
rect 4211 37031 4245 37065
rect 4279 37031 4313 37065
rect 4347 37031 4381 37065
rect 4415 37031 4449 37065
rect 4483 37031 4517 37065
rect 4551 37031 4585 37065
rect 4619 37031 4653 37065
rect 4687 37031 4721 37065
rect 4755 37031 4789 37065
rect 4823 37031 4857 37065
rect 4891 37031 4925 37065
rect 4959 37031 4993 37065
rect 5027 37031 5061 37065
rect 5095 37031 5129 37065
rect 5163 37031 5197 37065
rect 5231 37031 5265 37065
rect 5299 37031 5333 37065
rect 5367 37031 5401 37065
rect 5435 37031 5469 37065
rect 5503 37031 5537 37065
rect 5571 37031 5605 37065
rect 5639 37031 5673 37065
rect 5707 37031 5741 37065
rect 5775 37031 5809 37065
rect 5843 37031 5877 37065
rect 5911 37031 5945 37065
rect 5979 37031 6013 37065
rect 6047 37031 6081 37065
rect 6115 37031 6149 37065
rect 6183 37031 6217 37065
rect 6251 37031 6285 37065
rect 6319 37031 6353 37065
rect 6387 37031 6421 37065
rect 6455 37031 6489 37065
rect 6523 37031 6557 37065
rect 6591 37031 6625 37065
rect 6659 37031 6693 37065
rect 6727 37031 6761 37065
rect 6795 37031 6829 37065
rect 6863 37031 6897 37065
rect 6931 37031 6965 37065
rect 6999 37031 7033 37065
rect 7067 37031 7101 37065
rect 7135 37031 7169 37065
rect 7203 37031 7237 37065
rect 7271 37031 7305 37065
rect 7339 37031 7373 37065
rect 7407 37031 7441 37065
rect 7475 37031 7509 37065
rect 7543 37031 7577 37065
rect 7611 37031 7645 37065
rect 7679 37031 7713 37065
rect 3039 35065 3073 35099
rect 3108 35065 3142 35099
rect 3177 35065 3211 35099
rect 3246 35065 3280 35099
rect 3315 35065 3349 35099
rect 3384 35065 3418 35099
rect 3453 35065 3487 35099
rect 3522 35065 3556 35099
rect 3591 35065 3625 35099
rect 3660 35065 3694 35099
rect 3729 35065 3763 35099
rect 3798 35065 3832 35099
rect 3867 35065 3901 35099
rect 3936 35065 3970 35099
rect 4005 35065 4039 35099
rect 4074 35065 4108 35099
rect 4143 35065 4177 35099
rect 4211 35065 4245 35099
rect 4279 35065 4313 35099
rect 4347 35065 4381 35099
rect 4415 35065 4449 35099
rect 4483 35065 4517 35099
rect 4551 35065 4585 35099
rect 4619 35065 4653 35099
rect 4687 35065 4721 35099
rect 4755 35065 4789 35099
rect 4823 35065 4857 35099
rect 4891 35065 4925 35099
rect 4959 35065 4993 35099
rect 5027 35065 5061 35099
rect 5095 35065 5129 35099
rect 5163 35065 5197 35099
rect 5231 35065 5265 35099
rect 5299 35065 5333 35099
rect 5367 35065 5401 35099
rect 5435 35065 5469 35099
rect 5503 35065 5537 35099
rect 5571 35065 5605 35099
rect 5639 35065 5673 35099
rect 5707 35065 5741 35099
rect 5775 35065 5809 35099
rect 5843 35065 5877 35099
rect 5911 35065 5945 35099
rect 5979 35065 6013 35099
rect 6047 35065 6081 35099
rect 6115 35065 6149 35099
rect 6183 35065 6217 35099
rect 6251 35065 6285 35099
rect 6319 35065 6353 35099
rect 6387 35065 6421 35099
rect 6455 35065 6489 35099
rect 6523 35065 6557 35099
rect 6591 35065 6625 35099
rect 6659 35065 6693 35099
rect 6727 35065 6761 35099
rect 6795 35065 6829 35099
rect 6863 35065 6897 35099
rect 6931 35065 6965 35099
rect 6999 35065 7033 35099
rect 7067 35065 7101 35099
rect 7135 35065 7169 35099
rect 7203 35065 7237 35099
rect 7271 35065 7305 35099
rect 7339 35065 7373 35099
rect 7407 35065 7441 35099
rect 7475 35065 7509 35099
rect 7543 35065 7577 35099
rect 7611 35065 7645 35099
rect 7679 35065 7713 35099
rect 3039 33066 3073 33100
rect 3108 33066 3142 33100
rect 3177 33066 3211 33100
rect 3246 33066 3280 33100
rect 3315 33066 3349 33100
rect 3384 33066 3418 33100
rect 3453 33066 3487 33100
rect 3522 33066 3556 33100
rect 3591 33066 3625 33100
rect 3660 33066 3694 33100
rect 3729 33066 3763 33100
rect 3798 33066 3832 33100
rect 3867 33066 3901 33100
rect 3936 33066 3970 33100
rect 4005 33066 4039 33100
rect 4074 33066 4108 33100
rect 4143 33066 4177 33100
rect 4211 33066 4245 33100
rect 4279 33066 4313 33100
rect 4347 33066 4381 33100
rect 4415 33066 4449 33100
rect 4483 33066 4517 33100
rect 4551 33066 4585 33100
rect 4619 33066 4653 33100
rect 4687 33066 4721 33100
rect 4755 33066 4789 33100
rect 4823 33066 4857 33100
rect 4891 33066 4925 33100
rect 4959 33066 4993 33100
rect 5027 33066 5061 33100
rect 5095 33066 5129 33100
rect 5163 33066 5197 33100
rect 5231 33066 5265 33100
rect 5299 33066 5333 33100
rect 5367 33066 5401 33100
rect 5435 33066 5469 33100
rect 5503 33066 5537 33100
rect 5571 33066 5605 33100
rect 5639 33066 5673 33100
rect 5707 33066 5741 33100
rect 5775 33066 5809 33100
rect 5843 33066 5877 33100
rect 5911 33066 5945 33100
rect 5979 33066 6013 33100
rect 6047 33066 6081 33100
rect 6115 33066 6149 33100
rect 6183 33066 6217 33100
rect 6251 33066 6285 33100
rect 6319 33066 6353 33100
rect 6387 33066 6421 33100
rect 6455 33066 6489 33100
rect 6523 33066 6557 33100
rect 6591 33066 6625 33100
rect 6659 33066 6693 33100
rect 6727 33066 6761 33100
rect 6795 33066 6829 33100
rect 6863 33066 6897 33100
rect 6931 33066 6965 33100
rect 6999 33066 7033 33100
rect 7067 33066 7101 33100
rect 7135 33066 7169 33100
rect 7203 33066 7237 33100
rect 7271 33066 7305 33100
rect 7339 33066 7373 33100
rect 7407 33066 7441 33100
rect 7475 33066 7509 33100
rect 7543 33066 7577 33100
rect 7611 33066 7645 33100
rect 7679 33066 7713 33100
rect 3039 31043 3073 31077
rect 3108 31043 3142 31077
rect 3177 31043 3211 31077
rect 3246 31043 3280 31077
rect 3315 31043 3349 31077
rect 3384 31043 3418 31077
rect 3453 31043 3487 31077
rect 3522 31043 3556 31077
rect 3591 31043 3625 31077
rect 3660 31043 3694 31077
rect 3729 31043 3763 31077
rect 3798 31043 3832 31077
rect 3867 31043 3901 31077
rect 3936 31043 3970 31077
rect 4005 31043 4039 31077
rect 4074 31043 4108 31077
rect 4143 31043 4177 31077
rect 4211 31043 4245 31077
rect 4279 31043 4313 31077
rect 4347 31043 4381 31077
rect 4415 31043 4449 31077
rect 4483 31043 4517 31077
rect 4551 31043 4585 31077
rect 4619 31043 4653 31077
rect 4687 31043 4721 31077
rect 4755 31043 4789 31077
rect 4823 31043 4857 31077
rect 4891 31043 4925 31077
rect 4959 31043 4993 31077
rect 5027 31043 5061 31077
rect 5095 31043 5129 31077
rect 5163 31043 5197 31077
rect 5231 31043 5265 31077
rect 5299 31043 5333 31077
rect 5367 31043 5401 31077
rect 5435 31043 5469 31077
rect 5503 31043 5537 31077
rect 5571 31043 5605 31077
rect 5639 31043 5673 31077
rect 5707 31043 5741 31077
rect 5775 31043 5809 31077
rect 5843 31043 5877 31077
rect 5911 31043 5945 31077
rect 5979 31043 6013 31077
rect 6047 31043 6081 31077
rect 6115 31043 6149 31077
rect 6183 31043 6217 31077
rect 6251 31043 6285 31077
rect 6319 31043 6353 31077
rect 6387 31043 6421 31077
rect 6455 31043 6489 31077
rect 6523 31043 6557 31077
rect 6591 31043 6625 31077
rect 6659 31043 6693 31077
rect 6727 31043 6761 31077
rect 6795 31043 6829 31077
rect 6863 31043 6897 31077
rect 6931 31043 6965 31077
rect 6999 31043 7033 31077
rect 7067 31043 7101 31077
rect 7135 31043 7169 31077
rect 7203 31043 7237 31077
rect 7271 31043 7305 31077
rect 7339 31043 7373 31077
rect 7407 31043 7441 31077
rect 7475 31043 7509 31077
rect 7543 31043 7577 31077
rect 7611 31043 7645 31077
rect 7679 31043 7713 31077
rect 3039 29216 3073 29250
rect 3108 29216 3142 29250
rect 3177 29216 3211 29250
rect 3246 29216 3280 29250
rect 3315 29216 3349 29250
rect 3384 29216 3418 29250
rect 3453 29216 3487 29250
rect 3522 29216 3556 29250
rect 3591 29216 3625 29250
rect 3660 29216 3694 29250
rect 3729 29216 3763 29250
rect 3798 29216 3832 29250
rect 3867 29216 3901 29250
rect 3936 29216 3970 29250
rect 4005 29216 4039 29250
rect 4074 29216 4108 29250
rect 4143 29216 4177 29250
rect 4211 29216 4245 29250
rect 4279 29216 4313 29250
rect 4347 29216 4381 29250
rect 4415 29216 4449 29250
rect 4483 29216 4517 29250
rect 4551 29216 4585 29250
rect 4619 29216 4653 29250
rect 4687 29216 4721 29250
rect 4755 29216 4789 29250
rect 4823 29216 4857 29250
rect 4891 29216 4925 29250
rect 4959 29216 4993 29250
rect 5027 29216 5061 29250
rect 5095 29216 5129 29250
rect 5163 29216 5197 29250
rect 5231 29216 5265 29250
rect 5299 29216 5333 29250
rect 5367 29216 5401 29250
rect 5435 29216 5469 29250
rect 5503 29216 5537 29250
rect 5571 29216 5605 29250
rect 5639 29216 5673 29250
rect 5707 29216 5741 29250
rect 5775 29216 5809 29250
rect 5843 29216 5877 29250
rect 5911 29216 5945 29250
rect 5979 29216 6013 29250
rect 6047 29216 6081 29250
rect 6115 29216 6149 29250
rect 6183 29216 6217 29250
rect 6251 29216 6285 29250
rect 6319 29216 6353 29250
rect 6387 29216 6421 29250
rect 6455 29216 6489 29250
rect 6523 29216 6557 29250
rect 6591 29216 6625 29250
rect 6659 29216 6693 29250
rect 6727 29216 6761 29250
rect 6795 29216 6829 29250
rect 6863 29216 6897 29250
rect 6931 29216 6965 29250
rect 6999 29216 7033 29250
rect 7067 29216 7101 29250
rect 7135 29216 7169 29250
rect 7203 29216 7237 29250
rect 7271 29216 7305 29250
rect 7339 29216 7373 29250
rect 7407 29216 7441 29250
rect 7475 29216 7509 29250
rect 7543 29216 7577 29250
rect 7611 29216 7645 29250
rect 7679 29216 7713 29250
rect 5255 27071 5289 27105
rect 5325 27071 5359 27105
rect 5395 27071 5429 27105
rect 5465 27071 5499 27105
rect 5535 27071 5569 27105
rect 5605 27071 5639 27105
rect 5675 27071 5709 27105
rect 5745 27071 5779 27105
rect 5815 27071 5849 27105
rect 5885 27071 5919 27105
rect 5954 27071 5988 27105
rect 6023 27071 6057 27105
rect 6092 27071 6126 27105
rect 6161 27071 6195 27105
rect 6230 27071 6264 27105
rect 6299 27071 6333 27105
rect 6368 27071 6402 27105
rect 6437 27071 6471 27105
rect 6506 27071 6540 27105
rect 6575 27071 6609 27105
rect 6644 27071 6678 27105
rect 6713 27071 6747 27105
rect 6782 27071 6816 27105
rect 6851 27071 6885 27105
rect 6920 27071 6954 27105
rect 6989 27071 7023 27105
rect 7058 27071 7092 27105
rect 7127 27071 7161 27105
rect 7196 27071 7230 27105
rect 7265 27071 7299 27105
rect 7334 27071 7368 27105
rect 7403 27071 7437 27105
rect 7472 27071 7506 27105
rect 7541 27071 7575 27105
rect 7610 27071 7644 27105
rect 7679 27071 7713 27105
rect 5255 25078 5289 25112
rect 5325 25078 5359 25112
rect 5395 25078 5429 25112
rect 5465 25078 5499 25112
rect 5535 25078 5569 25112
rect 5605 25078 5639 25112
rect 5675 25078 5709 25112
rect 5745 25078 5779 25112
rect 5815 25078 5849 25112
rect 5885 25078 5919 25112
rect 5954 25078 5988 25112
rect 6023 25078 6057 25112
rect 6092 25078 6126 25112
rect 6161 25078 6195 25112
rect 6230 25078 6264 25112
rect 6299 25078 6333 25112
rect 6368 25078 6402 25112
rect 6437 25078 6471 25112
rect 6506 25078 6540 25112
rect 6575 25078 6609 25112
rect 6644 25078 6678 25112
rect 6713 25078 6747 25112
rect 6782 25078 6816 25112
rect 6851 25078 6885 25112
rect 6920 25078 6954 25112
rect 6989 25078 7023 25112
rect 7058 25078 7092 25112
rect 7127 25078 7161 25112
rect 7196 25078 7230 25112
rect 7265 25078 7299 25112
rect 7334 25078 7368 25112
rect 7403 25078 7437 25112
rect 7472 25078 7506 25112
rect 7541 25078 7575 25112
rect 7610 25078 7644 25112
rect 7679 25078 7713 25112
rect 5255 23090 5289 23124
rect 5325 23090 5359 23124
rect 5395 23090 5429 23124
rect 5465 23090 5499 23124
rect 5535 23090 5569 23124
rect 5605 23090 5639 23124
rect 5675 23090 5709 23124
rect 5745 23090 5779 23124
rect 5815 23090 5849 23124
rect 5885 23090 5919 23124
rect 5954 23090 5988 23124
rect 6023 23090 6057 23124
rect 6092 23090 6126 23124
rect 6161 23090 6195 23124
rect 6230 23090 6264 23124
rect 6299 23090 6333 23124
rect 6368 23090 6402 23124
rect 6437 23090 6471 23124
rect 6506 23090 6540 23124
rect 6575 23090 6609 23124
rect 6644 23090 6678 23124
rect 6713 23090 6747 23124
rect 6782 23090 6816 23124
rect 6851 23090 6885 23124
rect 6920 23090 6954 23124
rect 6989 23090 7023 23124
rect 7058 23090 7092 23124
rect 7127 23090 7161 23124
rect 7196 23090 7230 23124
rect 7265 23090 7299 23124
rect 7334 23090 7368 23124
rect 7403 23090 7437 23124
rect 7472 23090 7506 23124
rect 7541 23090 7575 23124
rect 7610 23090 7644 23124
rect 7679 23090 7713 23124
rect 5255 21049 5289 21083
rect 5325 21049 5359 21083
rect 5395 21049 5429 21083
rect 5465 21049 5499 21083
rect 5535 21049 5569 21083
rect 5605 21049 5639 21083
rect 5675 21049 5709 21083
rect 5745 21049 5779 21083
rect 5815 21049 5849 21083
rect 5885 21049 5919 21083
rect 5954 21049 5988 21083
rect 6023 21049 6057 21083
rect 6092 21049 6126 21083
rect 6161 21049 6195 21083
rect 6230 21049 6264 21083
rect 6299 21049 6333 21083
rect 6368 21049 6402 21083
rect 6437 21049 6471 21083
rect 6506 21049 6540 21083
rect 6575 21049 6609 21083
rect 6644 21049 6678 21083
rect 6713 21049 6747 21083
rect 6782 21049 6816 21083
rect 6851 21049 6885 21083
rect 6920 21049 6954 21083
rect 6989 21049 7023 21083
rect 7058 21049 7092 21083
rect 7127 21049 7161 21083
rect 7196 21049 7230 21083
rect 7265 21049 7299 21083
rect 7334 21049 7368 21083
rect 7403 21049 7437 21083
rect 7472 21049 7506 21083
rect 7541 21049 7575 21083
rect 7610 21049 7644 21083
rect 7679 21049 7713 21083
rect 5255 19085 5289 19119
rect 5325 19085 5359 19119
rect 5395 19085 5429 19119
rect 5465 19085 5499 19119
rect 5535 19085 5569 19119
rect 5605 19085 5639 19119
rect 5675 19085 5709 19119
rect 5745 19085 5779 19119
rect 5815 19085 5849 19119
rect 5885 19085 5919 19119
rect 5954 19085 5988 19119
rect 6023 19085 6057 19119
rect 6092 19085 6126 19119
rect 6161 19085 6195 19119
rect 6230 19085 6264 19119
rect 6299 19085 6333 19119
rect 6368 19085 6402 19119
rect 6437 19085 6471 19119
rect 6506 19085 6540 19119
rect 6575 19085 6609 19119
rect 6644 19085 6678 19119
rect 6713 19085 6747 19119
rect 6782 19085 6816 19119
rect 6851 19085 6885 19119
rect 6920 19085 6954 19119
rect 6989 19085 7023 19119
rect 7058 19085 7092 19119
rect 7127 19085 7161 19119
rect 7196 19085 7230 19119
rect 7265 19085 7299 19119
rect 7334 19085 7368 19119
rect 7403 19085 7437 19119
rect 7472 19085 7506 19119
rect 7541 19085 7575 19119
rect 7610 19085 7644 19119
rect 7679 19085 7713 19119
rect 5255 17211 5289 17245
rect 5325 17211 5359 17245
rect 5395 17211 5429 17245
rect 5465 17211 5499 17245
rect 5535 17211 5569 17245
rect 5605 17211 5639 17245
rect 5675 17211 5709 17245
rect 5745 17211 5779 17245
rect 5815 17211 5849 17245
rect 5885 17211 5919 17245
rect 5954 17211 5988 17245
rect 6023 17211 6057 17245
rect 6092 17211 6126 17245
rect 6161 17211 6195 17245
rect 6230 17211 6264 17245
rect 6299 17211 6333 17245
rect 6368 17211 6402 17245
rect 6437 17211 6471 17245
rect 6506 17211 6540 17245
rect 6575 17211 6609 17245
rect 6644 17211 6678 17245
rect 6713 17211 6747 17245
rect 6782 17211 6816 17245
rect 6851 17211 6885 17245
rect 6920 17211 6954 17245
rect 6989 17211 7023 17245
rect 7058 17211 7092 17245
rect 7127 17211 7161 17245
rect 7196 17211 7230 17245
rect 7265 17211 7299 17245
rect 7334 17211 7368 17245
rect 7403 17211 7437 17245
rect 7472 17211 7506 17245
rect 7541 17211 7575 17245
rect 7610 17211 7644 17245
rect 7679 17211 7713 17245
rect 3039 15552 3073 15586
rect 3108 15552 3142 15586
rect 3177 15552 3211 15586
rect 3246 15552 3280 15586
rect 3315 15552 3349 15586
rect 3384 15552 3418 15586
rect 3453 15552 3487 15586
rect 3522 15552 3556 15586
rect 3591 15552 3625 15586
rect 3660 15552 3694 15586
rect 3729 15552 3763 15586
rect 3798 15552 3832 15586
rect 3867 15552 3901 15586
rect 3936 15552 3970 15586
rect 4005 15552 4039 15586
rect 4074 15552 4108 15586
rect 4143 15552 4177 15586
rect 4211 15552 4245 15586
rect 4279 15552 4313 15586
rect 4347 15552 4381 15586
rect 4415 15552 4449 15586
rect 4483 15552 4517 15586
rect 4551 15552 4585 15586
rect 4619 15552 4653 15586
rect 4687 15552 4721 15586
rect 4755 15552 4789 15586
rect 4823 15552 4857 15586
rect 4891 15552 4925 15586
rect 4959 15552 4993 15586
rect 5027 15552 5061 15586
rect 5095 15552 5129 15586
rect 5163 15552 5197 15586
rect 5231 15552 5265 15586
rect 5299 15552 5333 15586
rect 5367 15552 5401 15586
rect 5435 15552 5469 15586
rect 5503 15552 5537 15586
rect 5571 15552 5605 15586
rect 5639 15552 5673 15586
rect 5707 15552 5741 15586
rect 5775 15552 5809 15586
rect 5843 15552 5877 15586
rect 5911 15552 5945 15586
rect 5979 15552 6013 15586
rect 6047 15552 6081 15586
rect 6115 15552 6149 15586
rect 6183 15552 6217 15586
rect 6251 15552 6285 15586
rect 6319 15552 6353 15586
rect 6387 15552 6421 15586
rect 6455 15552 6489 15586
rect 6523 15552 6557 15586
rect 6591 15552 6625 15586
rect 6659 15552 6693 15586
rect 6727 15552 6761 15586
rect 6795 15552 6829 15586
rect 6863 15552 6897 15586
rect 6931 15552 6965 15586
rect 6999 15552 7033 15586
rect 7067 15552 7101 15586
rect 7135 15552 7169 15586
rect 7203 15552 7237 15586
rect 7271 15552 7305 15586
rect 7339 15552 7373 15586
rect 7407 15552 7441 15586
rect 7475 15552 7509 15586
rect 7543 15552 7577 15586
rect 7611 15552 7645 15586
rect 7679 15552 7713 15586
rect 3039 13822 3073 13856
rect 3108 13822 3142 13856
rect 3177 13822 3211 13856
rect 3246 13822 3280 13856
rect 3315 13822 3349 13856
rect 3384 13822 3418 13856
rect 3453 13822 3487 13856
rect 3522 13822 3556 13856
rect 3591 13822 3625 13856
rect 3660 13822 3694 13856
rect 3729 13822 3763 13856
rect 3798 13822 3832 13856
rect 3867 13822 3901 13856
rect 3936 13822 3970 13856
rect 4005 13822 4039 13856
rect 4073 13822 4107 13856
rect 4141 13822 4175 13856
rect 4209 13822 4243 13856
rect 4277 13822 4311 13856
rect 4345 13822 4379 13856
rect 4413 13822 4447 13856
rect 4481 13822 4515 13856
rect 4549 13822 4583 13856
rect 4617 13822 4651 13856
rect 4685 13822 4719 13856
rect 4753 13822 4787 13856
rect 4821 13822 4855 13856
rect 4889 13822 4923 13856
rect 4957 13822 4991 13856
rect 5025 13822 5059 13856
rect 5093 13822 5127 13856
rect 5161 13822 5195 13856
rect 5229 13822 5263 13856
rect 5297 13822 5331 13856
rect 5365 13822 5399 13856
rect 5433 13822 5467 13856
rect 5501 13822 5535 13856
rect 5569 13822 5603 13856
rect 5637 13822 5671 13856
rect 5705 13822 5739 13856
rect 5773 13822 5807 13856
rect 5841 13822 5875 13856
rect 5909 13822 5943 13856
rect 5977 13822 6011 13856
rect 6045 13822 6079 13856
rect 6113 13822 6147 13856
rect 6181 13822 6215 13856
rect 6249 13822 6283 13856
rect 6317 13822 6351 13856
rect 6385 13822 6419 13856
rect 6453 13822 6487 13856
rect 6521 13822 6555 13856
rect 6589 13822 6623 13856
rect 6657 13822 6691 13856
rect 6725 13822 6759 13856
rect 6793 13822 6827 13856
rect 6861 13822 6895 13856
rect 6929 13822 6963 13856
rect 6997 13822 7031 13856
rect 7065 13822 7099 13856
rect 7133 13822 7167 13856
rect 7201 13822 7235 13856
rect 7269 13822 7303 13856
rect 7337 13822 7371 13856
rect 7405 13822 7439 13856
rect 7473 13822 7507 13856
rect 7541 13822 7575 13856
rect 7609 13822 7643 13856
rect 7677 13822 7711 13856
rect 3039 11784 3073 11818
rect 3108 11784 3142 11818
rect 3177 11784 3211 11818
rect 3246 11784 3280 11818
rect 3315 11784 3349 11818
rect 3384 11784 3418 11818
rect 3453 11784 3487 11818
rect 3522 11784 3556 11818
rect 3591 11784 3625 11818
rect 3660 11784 3694 11818
rect 3729 11784 3763 11818
rect 3798 11784 3832 11818
rect 3867 11784 3901 11818
rect 3936 11784 3970 11818
rect 4005 11784 4039 11818
rect 4073 11784 4107 11818
rect 4141 11784 4175 11818
rect 4209 11784 4243 11818
rect 4277 11784 4311 11818
rect 4345 11784 4379 11818
rect 4413 11784 4447 11818
rect 4481 11784 4515 11818
rect 4549 11784 4583 11818
rect 4617 11784 4651 11818
rect 4685 11784 4719 11818
rect 4753 11784 4787 11818
rect 4821 11784 4855 11818
rect 4889 11784 4923 11818
rect 4957 11784 4991 11818
rect 5025 11784 5059 11818
rect 5093 11784 5127 11818
rect 5161 11784 5195 11818
rect 5229 11784 5263 11818
rect 5297 11784 5331 11818
rect 5365 11784 5399 11818
rect 5433 11784 5467 11818
rect 5501 11784 5535 11818
rect 5569 11784 5603 11818
rect 5637 11784 5671 11818
rect 5705 11784 5739 11818
rect 5773 11784 5807 11818
rect 5841 11784 5875 11818
rect 5909 11784 5943 11818
rect 5977 11784 6011 11818
rect 6045 11784 6079 11818
rect 6113 11784 6147 11818
rect 6181 11784 6215 11818
rect 6249 11784 6283 11818
rect 6317 11784 6351 11818
rect 6385 11784 6419 11818
rect 6453 11784 6487 11818
rect 6521 11784 6555 11818
rect 6589 11784 6623 11818
rect 6657 11784 6691 11818
rect 6725 11784 6759 11818
rect 6793 11784 6827 11818
rect 6861 11784 6895 11818
rect 6929 11784 6963 11818
rect 6997 11784 7031 11818
rect 7065 11784 7099 11818
rect 7133 11784 7167 11818
rect 7201 11784 7235 11818
rect 7269 11784 7303 11818
rect 7337 11784 7371 11818
rect 7405 11784 7439 11818
rect 7473 11784 7507 11818
rect 7541 11784 7575 11818
rect 7609 11784 7643 11818
rect 7677 11784 7711 11818
rect 3039 10022 3073 10056
rect 3108 10022 3142 10056
rect 3177 10022 3211 10056
rect 3246 10022 3280 10056
rect 3315 10022 3349 10056
rect 3384 10022 3418 10056
rect 3453 10022 3487 10056
rect 3522 10022 3556 10056
rect 3591 10022 3625 10056
rect 3660 10022 3694 10056
rect 3729 10022 3763 10056
rect 3798 10022 3832 10056
rect 3867 10022 3901 10056
rect 3936 10022 3970 10056
rect 4005 10022 4039 10056
rect 4074 10022 4108 10056
rect 4143 10022 4177 10056
rect 4211 10022 4245 10056
rect 4279 10022 4313 10056
rect 4347 10022 4381 10056
rect 4415 10022 4449 10056
rect 4483 10022 4517 10056
rect 4551 10022 4585 10056
rect 4619 10022 4653 10056
rect 4687 10022 4721 10056
rect 4755 10022 4789 10056
rect 4823 10022 4857 10056
rect 4891 10022 4925 10056
rect 4959 10022 4993 10056
rect 5027 10022 5061 10056
rect 5095 10022 5129 10056
rect 5163 10022 5197 10056
rect 5231 10022 5265 10056
rect 5299 10022 5333 10056
rect 5367 10022 5401 10056
rect 5435 10022 5469 10056
rect 5503 10022 5537 10056
rect 5571 10022 5605 10056
rect 5639 10022 5673 10056
rect 5707 10022 5741 10056
rect 5775 10022 5809 10056
rect 5843 10022 5877 10056
rect 5911 10022 5945 10056
rect 5979 10022 6013 10056
rect 6047 10022 6081 10056
rect 6115 10022 6149 10056
rect 6183 10022 6217 10056
rect 6251 10022 6285 10056
rect 6319 10022 6353 10056
rect 6387 10022 6421 10056
rect 6455 10022 6489 10056
rect 6523 10022 6557 10056
rect 6591 10022 6625 10056
rect 6659 10022 6693 10056
rect 6727 10022 6761 10056
rect 6795 10022 6829 10056
rect 6863 10022 6897 10056
rect 6931 10022 6965 10056
rect 6999 10022 7033 10056
rect 7067 10022 7101 10056
rect 7135 10022 7169 10056
rect 7203 10022 7237 10056
rect 7271 10022 7305 10056
rect 7339 10022 7373 10056
rect 7407 10022 7441 10056
rect 7475 10022 7509 10056
rect 7543 10022 7577 10056
rect 7611 10022 7645 10056
rect 7679 10022 7713 10056
rect 2488 9306 2522 9340
rect 2556 9306 2590 9340
rect 2624 9306 2658 9340
rect 2692 9306 2726 9340
rect 2760 9306 2794 9340
rect 2828 9306 2862 9340
rect 2896 9306 2930 9340
rect 2964 9306 2998 9340
rect 3032 9306 3066 9340
rect 3100 9306 3134 9340
rect 3168 9306 3202 9340
rect 3236 9306 3270 9340
rect 3304 9306 3338 9340
rect 3372 9306 3406 9340
rect 3440 9306 3474 9340
rect 3508 9306 3542 9340
rect 3576 9306 3610 9340
rect 3644 9306 3678 9340
rect 3712 9306 3746 9340
rect 3780 9306 3814 9340
rect 3848 9306 3882 9340
rect 3916 9306 3950 9340
rect 3984 9306 4018 9340
rect 4052 9306 4086 9340
rect 4120 9306 4154 9340
rect 4188 9306 4222 9340
rect 4256 9306 4290 9340
rect 4324 9306 4358 9340
rect 4392 9306 4426 9340
rect 4460 9306 4494 9340
rect 4528 9306 4562 9340
rect 4596 9306 4630 9340
rect 4664 9306 4698 9340
rect 4732 9306 4766 9340
rect 4800 9306 4834 9340
rect 4868 9306 4902 9340
rect 4936 9306 4970 9340
rect 5004 9306 5038 9340
rect 5072 9306 5106 9340
rect 5140 9306 5174 9340
rect 5208 9306 5242 9340
rect 5276 9306 5310 9340
rect 5344 9306 5378 9340
rect 5412 9306 5446 9340
rect 5480 9306 5514 9340
rect 5548 9306 5582 9340
rect 5616 9306 5650 9340
rect 5684 9306 5718 9340
rect 5752 9306 5786 9340
rect 5820 9306 5854 9340
rect 5888 9306 5922 9340
rect 5956 9306 5990 9340
rect 6024 9306 6058 9340
rect 6092 9306 6126 9340
rect 6160 9306 6194 9340
rect 6228 9306 6262 9340
rect 6296 9306 6330 9340
rect 6364 9306 6398 9340
rect 6432 9306 6466 9340
rect 6500 9306 6534 9340
rect 6568 9306 6602 9340
rect 6636 9306 6670 9340
rect 6704 9306 6738 9340
rect 6772 9306 6806 9340
rect 6840 9306 6874 9340
rect 6908 9306 6942 9340
rect 6976 9306 7010 9340
rect 7044 9306 7078 9340
rect 7112 9306 7146 9340
rect 7180 9306 7214 9340
rect 7248 9306 7282 9340
rect 7316 9306 7350 9340
rect 2488 7506 2522 7540
rect 2556 7506 2590 7540
rect 2624 7506 2658 7540
rect 2692 7506 2726 7540
rect 2760 7506 2794 7540
rect 2828 7506 2862 7540
rect 2896 7506 2930 7540
rect 2964 7506 2998 7540
rect 3032 7506 3066 7540
rect 3100 7506 3134 7540
rect 3168 7506 3202 7540
rect 3236 7506 3270 7540
rect 3304 7506 3338 7540
rect 3372 7506 3406 7540
rect 3440 7506 3474 7540
rect 3508 7506 3542 7540
rect 3576 7506 3610 7540
rect 3644 7506 3678 7540
rect 3712 7506 3746 7540
rect 3780 7506 3814 7540
rect 3848 7506 3882 7540
rect 3916 7506 3950 7540
rect 3984 7506 4018 7540
rect 4052 7506 4086 7540
rect 4120 7506 4154 7540
rect 4188 7506 4222 7540
rect 4256 7506 4290 7540
rect 4324 7506 4358 7540
rect 4392 7506 4426 7540
rect 4460 7506 4494 7540
rect 4528 7506 4562 7540
rect 4596 7506 4630 7540
rect 4664 7506 4698 7540
rect 4732 7506 4766 7540
rect 4800 7506 4834 7540
rect 4868 7506 4902 7540
rect 4936 7506 4970 7540
rect 5004 7506 5038 7540
rect 5072 7506 5106 7540
rect 5140 7506 5174 7540
rect 5208 7506 5242 7540
rect 5276 7506 5310 7540
rect 5344 7506 5378 7540
rect 5412 7506 5446 7540
rect 5480 7506 5514 7540
rect 5548 7506 5582 7540
rect 5616 7506 5650 7540
rect 5684 7506 5718 7540
rect 5752 7506 5786 7540
rect 5820 7506 5854 7540
rect 5888 7506 5922 7540
rect 5956 7506 5990 7540
rect 6024 7506 6058 7540
rect 6092 7506 6126 7540
rect 6160 7506 6194 7540
rect 6228 7506 6262 7540
rect 6296 7506 6330 7540
rect 6364 7506 6398 7540
rect 6432 7506 6466 7540
rect 6500 7506 6534 7540
rect 6568 7506 6602 7540
rect 6636 7506 6670 7540
rect 6704 7506 6738 7540
rect 6772 7506 6806 7540
rect 6840 7506 6874 7540
rect 6908 7506 6942 7540
rect 6976 7506 7010 7540
rect 7044 7506 7078 7540
rect 7112 7506 7146 7540
rect 7180 7506 7214 7540
rect 7248 7506 7282 7540
rect 7316 7506 7350 7540
rect 2660 5611 2694 5645
rect 2728 5611 2762 5645
rect 2796 5611 2830 5645
rect 2864 5611 2898 5645
rect 2932 5611 2966 5645
rect 3000 5611 3034 5645
rect 3068 5611 3102 5645
rect 3136 5611 3170 5645
rect 3204 5611 3238 5645
rect 3272 5611 3306 5645
rect 3340 5611 3374 5645
rect 3408 5611 3442 5645
rect 3476 5611 3510 5645
rect 3544 5611 3578 5645
rect 3612 5611 3646 5645
rect 3680 5611 3714 5645
rect 3748 5611 3782 5645
rect 3816 5611 3850 5645
rect 3884 5611 3918 5645
rect 3952 5611 3986 5645
rect 4020 5611 4054 5645
rect 4088 5611 4122 5645
rect 4156 5611 4190 5645
rect 4224 5611 4258 5645
rect 4292 5611 4326 5645
rect 4360 5611 4394 5645
rect 4428 5611 4462 5645
rect 4496 5611 4530 5645
rect 4564 5611 4598 5645
rect 4632 5611 4666 5645
rect 4700 5611 4734 5645
rect 4768 5611 4802 5645
rect 4836 5611 4870 5645
rect 4904 5611 4938 5645
rect 4972 5611 5006 5645
rect 5040 5611 5074 5645
rect 5108 5611 5142 5645
rect 5176 5611 5210 5645
rect 5244 5611 5278 5645
rect 5312 5611 5346 5645
rect 5380 5611 5414 5645
rect 5448 5611 5482 5645
rect 5516 5611 5550 5645
rect 5584 5611 5618 5645
rect 5652 5611 5686 5645
rect 5720 5611 5754 5645
rect 5788 5611 5822 5645
rect 5856 5611 5890 5645
rect 5924 5611 5958 5645
rect 5992 5611 6026 5645
rect 6060 5611 6094 5645
rect 6128 5611 6162 5645
rect 6196 5611 6230 5645
rect 6264 5611 6298 5645
rect 6332 5611 6366 5645
rect 6400 5611 6434 5645
rect 6468 5611 6502 5645
rect 6536 5611 6570 5645
rect 6604 5611 6638 5645
rect 6672 5611 6706 5645
rect 6740 5611 6774 5645
rect 6808 5611 6842 5645
rect 6876 5611 6910 5645
rect 6944 5611 6978 5645
rect 1919 1822 1953 1856
rect 1919 1750 1953 1784
rect 1919 1678 1953 1712
rect 1919 1606 1953 1640
rect 1919 1534 1953 1568
rect 1919 1462 1953 1496
rect 1919 1389 1953 1423
rect 1919 1316 1953 1350
rect 1919 1243 1953 1277
rect 1919 1170 1953 1204
rect 1919 1097 1953 1131
rect 1919 1024 1953 1058
rect 3449 1822 3483 1856
rect 3449 1750 3483 1784
rect 3449 1678 3483 1712
rect 3449 1606 3483 1640
rect 3449 1534 3483 1568
rect 3449 1462 3483 1496
rect 3449 1389 3483 1423
rect 3449 1316 3483 1350
rect 3449 1243 3483 1277
rect 3449 1170 3483 1204
rect 3449 1097 3483 1131
rect 3449 1024 3483 1058
rect 170 187 204 221
rect 170 119 204 153
rect 1628 187 1662 221
rect 1628 119 1662 153
<< locali >>
rect 1938 39474 2163 39476
rect 2989 39474 3028 39476
rect 3062 39474 3101 39476
rect 3135 39474 3174 39476
rect 3208 39474 3247 39476
rect 3281 39474 3320 39476
rect 3354 39474 3393 39476
rect 3427 39474 3466 39476
rect 3500 39474 3539 39476
rect 3573 39474 3612 39476
rect 3646 39474 3685 39476
rect 3719 39474 3758 39476
rect 3792 39474 3831 39476
rect 3865 39474 3904 39476
rect 3938 39474 3977 39476
rect 4011 39474 4050 39476
rect 4084 39474 4123 39476
rect 4157 39474 4196 39476
rect 4230 39474 4269 39476
rect 4303 39474 4342 39476
rect 4376 39474 4415 39476
rect 4449 39474 4488 39476
rect 4522 39474 4561 39476
rect 4595 39474 4634 39476
rect 4668 39474 4707 39476
rect 4741 39474 4780 39476
rect 4814 39474 4853 39476
rect 4887 39474 4926 39476
rect 4960 39474 4999 39476
rect 5033 39474 5072 39476
rect 5106 39474 5145 39476
rect 5179 39474 5218 39476
rect 5252 39474 5291 39476
rect 5325 39474 5364 39476
rect 5398 39474 5437 39476
rect 5471 39474 5510 39476
rect 5544 39474 5583 39476
rect 5617 39474 5656 39476
rect 5690 39474 5729 39476
rect 5763 39474 5802 39476
rect 5836 39474 5875 39476
rect 5909 39474 5948 39476
rect 5982 39474 6021 39476
rect 6055 39474 6094 39476
rect 6128 39474 6167 39476
rect 6201 39474 6240 39476
rect 6274 39474 6313 39476
rect 6347 39474 6386 39476
rect 6420 39474 6459 39476
rect 6493 39474 6532 39476
rect 6566 39474 6605 39476
rect 6639 39474 6678 39476
rect 6712 39474 6751 39476
rect 6785 39474 6824 39476
rect 6858 39474 6897 39476
rect 6931 39474 6970 39476
rect 7004 39474 7043 39476
rect 7077 39474 7116 39476
rect 7150 39474 7189 39476
rect 7223 39474 7262 39476
rect 7296 39474 7335 39476
rect 7369 39474 7408 39476
rect 7442 39474 7481 39476
rect 7515 39474 7554 39476
rect 7588 39474 7627 39476
rect 7661 39474 7786 39476
rect 7820 39474 7866 39476
rect 7900 39474 7946 39476
rect 7980 39474 8026 39476
rect 8060 39474 8106 39476
rect 8140 39474 8186 39476
rect 8220 39474 8267 39476
rect 8301 39474 8348 39476
rect 8382 39474 8429 39476
rect 8463 39474 8535 39476
rect 1938 39470 2039 39474
rect 1938 34108 1944 39470
rect 2073 39440 2107 39474
rect 2050 39372 2107 39440
rect 8465 39404 8535 39474
rect 2050 39370 2163 39372
rect 2989 39370 3028 39372
rect 3062 39370 3101 39372
rect 3135 39370 3174 39372
rect 3208 39370 3247 39372
rect 3281 39370 3320 39372
rect 3354 39370 3393 39372
rect 3427 39370 3466 39372
rect 3500 39370 3539 39372
rect 3573 39370 3612 39372
rect 3646 39370 3685 39372
rect 3719 39370 3758 39372
rect 3792 39370 3831 39372
rect 3865 39370 3904 39372
rect 3938 39370 3977 39372
rect 4011 39370 4050 39372
rect 4084 39370 4123 39372
rect 4157 39370 4196 39372
rect 4230 39370 4269 39372
rect 4303 39370 4342 39372
rect 4376 39370 4415 39372
rect 4449 39370 4488 39372
rect 4522 39370 4561 39372
rect 4595 39370 4634 39372
rect 4668 39370 4707 39372
rect 4741 39370 4780 39372
rect 4814 39370 4853 39372
rect 4887 39370 4926 39372
rect 4960 39370 4999 39372
rect 5033 39370 5072 39372
rect 5106 39370 5145 39372
rect 5179 39370 5218 39372
rect 5252 39370 5291 39372
rect 5325 39370 5364 39372
rect 5398 39370 5437 39372
rect 5471 39370 5510 39372
rect 5544 39370 5583 39372
rect 5617 39370 5656 39372
rect 5690 39370 5729 39372
rect 5763 39370 5802 39372
rect 5836 39370 5875 39372
rect 5909 39370 5948 39372
rect 5982 39370 6021 39372
rect 6055 39370 6094 39372
rect 6128 39370 6167 39372
rect 6201 39370 6240 39372
rect 6274 39370 6313 39372
rect 6347 39370 6386 39372
rect 6420 39370 6459 39372
rect 6493 39370 6532 39372
rect 6566 39370 6605 39372
rect 6639 39370 6678 39372
rect 6712 39370 6751 39372
rect 6785 39370 6824 39372
rect 6858 39370 6897 39372
rect 6931 39370 6970 39372
rect 7004 39370 7043 39372
rect 7077 39370 7116 39372
rect 7150 39370 7189 39372
rect 7223 39370 7262 39372
rect 7296 39370 7335 39372
rect 7369 39370 7408 39372
rect 7442 39370 7481 39372
rect 7515 39370 7554 39372
rect 7588 39370 7627 39372
rect 7661 39370 7786 39372
rect 7820 39370 7866 39372
rect 7900 39370 7946 39372
rect 7980 39370 8026 39372
rect 8060 39370 8106 39372
rect 8140 39370 8186 39372
rect 8220 39370 8267 39372
rect 8301 39370 8348 39372
rect 8382 39370 8429 39372
rect 2050 34108 2056 39370
rect 1938 34069 1946 34108
rect 2048 34069 2056 34108
rect 1938 34035 1944 34069
rect 2050 34035 2056 34069
rect 1938 33996 1946 34035
rect 2048 33996 2056 34035
rect 1938 33962 1944 33996
rect 2050 33962 2056 33996
rect 1938 33923 1946 33962
rect 2048 33923 2056 33962
rect 1938 33889 1944 33923
rect 2050 33889 2056 33923
rect 1938 33850 1946 33889
rect 2048 33850 2056 33889
rect 1938 33816 1944 33850
rect 2050 33816 2056 33850
rect 1938 33777 1946 33816
rect 2048 33777 2056 33816
rect 1938 33743 1944 33777
rect 2050 33743 2056 33777
rect 1938 33704 1946 33743
rect 2048 33704 2056 33743
rect 1938 33670 1944 33704
rect 2050 33670 2056 33704
rect 1938 33607 1946 33670
rect 2048 33607 2056 33670
rect 1938 11037 1944 33607
rect 2050 11037 2056 33607
rect 1938 10998 1946 11037
rect 2048 10998 2056 11037
rect 1938 10964 1944 10998
rect 2050 10964 2056 10998
rect 1938 10925 1946 10964
rect 2048 10925 2056 10964
rect 1938 10891 1944 10925
rect 2050 10891 2056 10925
rect 1938 10847 1946 10891
rect 2048 10847 2056 10891
rect 1938 10813 1944 10847
rect 2050 10813 2056 10847
rect 1938 10774 1946 10813
rect 2048 10774 2056 10813
rect 1938 10740 1944 10774
rect 2050 10740 2056 10774
rect 1938 10701 1946 10740
rect 2048 10701 2056 10740
rect 1938 10667 1944 10701
rect 2050 10667 2056 10701
rect 1938 10628 1946 10667
rect 2048 10628 2056 10667
rect 1938 8938 1944 10628
rect 2050 9705 2056 10628
rect 2274 39141 2405 39142
rect 2439 39141 2473 39142
rect 2274 39107 2348 39141
rect 2382 39108 2405 39141
rect 2382 39107 2420 39108
rect 2454 39107 2473 39141
rect 2274 39074 2473 39107
rect 2376 39040 2473 39074
rect 8151 39069 8219 39142
rect 8151 39040 8184 39069
rect 2376 39007 2541 39040
rect 8083 39035 8184 39040
rect 8218 39035 8219 39069
rect 8083 39023 8219 39035
rect 8083 39007 8185 39023
rect 2376 39006 2410 39007
rect 2444 38973 2482 39007
rect 2516 38973 2541 39007
rect 8084 38997 8185 39007
rect 8084 38973 8184 38997
rect 2444 38972 2541 38973
rect 8083 38972 8184 38973
rect 8049 38963 8184 38972
rect 8218 38963 8219 38989
rect 8049 38955 8219 38963
rect 8049 38935 8117 38955
rect 8049 38901 8050 38935
rect 8084 38901 8117 38935
rect 8049 38887 8117 38901
rect 3023 38820 3035 38854
rect 3073 38820 3108 38854
rect 3142 38820 3177 38854
rect 3215 38820 3246 38854
rect 3288 38820 3315 38854
rect 3361 38820 3384 38854
rect 3434 38820 3453 38854
rect 3507 38820 3522 38854
rect 3580 38820 3591 38854
rect 3653 38820 3660 38854
rect 3726 38820 3729 38854
rect 3763 38820 3765 38854
rect 3832 38820 3838 38854
rect 3901 38820 3911 38854
rect 3970 38820 3984 38854
rect 4039 38820 4057 38854
rect 4108 38820 4130 38854
rect 4177 38820 4203 38854
rect 4245 38820 4276 38854
rect 4313 38820 4347 38854
rect 4383 38820 4415 38854
rect 4456 38820 4483 38854
rect 4529 38820 4551 38854
rect 4602 38820 4619 38854
rect 4675 38820 4687 38854
rect 4748 38820 4755 38854
rect 4821 38820 4823 38854
rect 4857 38820 4860 38854
rect 4925 38820 4933 38854
rect 4993 38820 5006 38854
rect 5061 38820 5079 38854
rect 5129 38820 5152 38854
rect 5197 38820 5225 38854
rect 5265 38820 5298 38854
rect 5333 38820 5367 38854
rect 5405 38820 5435 38854
rect 5478 38820 5503 38854
rect 5551 38820 5571 38854
rect 5624 38820 5639 38854
rect 5697 38820 5707 38854
rect 5770 38820 5775 38854
rect 5877 38820 5882 38854
rect 5945 38820 5955 38854
rect 6013 38820 6027 38854
rect 6081 38820 6099 38854
rect 6149 38820 6171 38854
rect 6217 38820 6243 38854
rect 6285 38820 6315 38854
rect 6353 38820 6387 38854
rect 6421 38820 6455 38854
rect 6493 38820 6523 38854
rect 6565 38820 6591 38854
rect 6637 38820 6659 38854
rect 6709 38820 6727 38854
rect 6781 38820 6795 38854
rect 6853 38820 6863 38854
rect 6925 38820 6931 38854
rect 6997 38820 6999 38854
rect 7033 38820 7035 38854
rect 7101 38820 7107 38854
rect 7169 38820 7179 38854
rect 7237 38820 7251 38854
rect 7305 38820 7323 38854
rect 7373 38820 7395 38854
rect 7441 38820 7467 38854
rect 7509 38820 7539 38854
rect 7577 38820 7611 38854
rect 7645 38820 7679 38854
rect 7717 38820 7729 38854
rect 3109 38714 3211 38726
rect 3663 38714 3765 38726
rect 4217 38714 4319 38726
rect 4771 38714 4873 38726
rect 5325 38714 5427 38726
rect 5879 38714 5981 38726
rect 6987 38714 7089 38726
rect 7539 38714 7645 38726
rect 2864 38680 2902 38714
rect 2830 38641 2936 38680
rect 2864 38607 2902 38641
rect 2830 38568 2936 38607
rect 2864 38534 2902 38568
rect 2830 38495 2936 38534
rect 2864 38461 2902 38495
rect 2830 38422 2936 38461
rect 3141 38680 3179 38714
rect 3107 38641 3213 38680
rect 3141 38607 3179 38641
rect 3107 38568 3213 38607
rect 3141 38534 3179 38568
rect 3107 38495 3213 38534
rect 3141 38461 3179 38495
rect 3107 38422 3213 38461
rect 3418 38680 3456 38714
rect 3384 38641 3490 38680
rect 3418 38607 3456 38641
rect 3384 38568 3490 38607
rect 3418 38534 3456 38568
rect 3384 38495 3490 38534
rect 3418 38461 3456 38495
rect 3384 38422 3490 38461
rect 3695 38680 3733 38714
rect 3661 38641 3767 38680
rect 3695 38607 3733 38641
rect 3661 38568 3767 38607
rect 3695 38534 3733 38568
rect 3661 38495 3767 38534
rect 3695 38461 3733 38495
rect 3661 38422 3767 38461
rect 3972 38680 4010 38714
rect 3938 38641 4044 38680
rect 3972 38607 4010 38641
rect 3938 38568 4044 38607
rect 3972 38534 4010 38568
rect 3938 38495 4044 38534
rect 3972 38461 4010 38495
rect 3938 38422 4044 38461
rect 4249 38680 4287 38714
rect 4215 38641 4321 38680
rect 4249 38607 4287 38641
rect 4215 38568 4321 38607
rect 4249 38534 4287 38568
rect 4215 38495 4321 38534
rect 4249 38461 4287 38495
rect 4215 38422 4321 38461
rect 4526 38680 4564 38714
rect 4492 38641 4598 38680
rect 4526 38607 4564 38641
rect 4492 38568 4598 38607
rect 4526 38534 4564 38568
rect 4492 38495 4598 38534
rect 4526 38461 4564 38495
rect 4492 38422 4598 38461
rect 4803 38680 4841 38714
rect 4769 38641 4875 38680
rect 4803 38607 4841 38641
rect 4769 38568 4875 38607
rect 4803 38534 4841 38568
rect 4769 38495 4875 38534
rect 4803 38461 4841 38495
rect 4769 38422 4875 38461
rect 5080 38680 5118 38714
rect 5046 38641 5152 38680
rect 5080 38607 5118 38641
rect 5046 38568 5152 38607
rect 5080 38534 5118 38568
rect 5046 38495 5152 38534
rect 5080 38461 5118 38495
rect 5046 38422 5152 38461
rect 5357 38680 5395 38714
rect 5323 38641 5429 38680
rect 5357 38607 5395 38641
rect 5323 38568 5429 38607
rect 5357 38534 5395 38568
rect 5323 38495 5429 38534
rect 5357 38461 5395 38495
rect 5323 38422 5429 38461
rect 5634 38680 5672 38714
rect 5600 38641 5706 38680
rect 5634 38607 5672 38641
rect 5600 38568 5706 38607
rect 5634 38534 5672 38568
rect 5600 38495 5706 38534
rect 5634 38461 5672 38495
rect 5600 38422 5706 38461
rect 5911 38680 5949 38714
rect 5877 38641 5983 38680
rect 5911 38607 5949 38641
rect 5877 38568 5983 38607
rect 5911 38534 5949 38568
rect 5877 38495 5983 38534
rect 5911 38461 5949 38495
rect 5877 38422 5983 38461
rect 6188 38680 6226 38714
rect 6154 38641 6260 38680
rect 6188 38607 6226 38641
rect 6154 38568 6260 38607
rect 6188 38534 6226 38568
rect 6154 38495 6260 38534
rect 6188 38461 6226 38495
rect 6154 38422 6260 38461
rect 6465 38680 6503 38714
rect 6431 38641 6537 38680
rect 6465 38607 6503 38641
rect 6431 38568 6537 38607
rect 6465 38534 6503 38568
rect 6431 38495 6537 38534
rect 6465 38461 6503 38495
rect 6431 38422 6537 38461
rect 6742 38680 6780 38714
rect 6708 38641 6814 38680
rect 6742 38607 6780 38641
rect 6708 38568 6814 38607
rect 6742 38534 6780 38568
rect 6708 38495 6814 38534
rect 6742 38461 6780 38495
rect 6708 38422 6814 38461
rect 7019 38680 7057 38714
rect 6985 38641 7091 38680
rect 7019 38607 7057 38641
rect 6985 38568 7091 38607
rect 7019 38534 7057 38568
rect 6985 38495 7091 38534
rect 7019 38461 7057 38495
rect 6985 38422 7091 38461
rect 7296 38680 7334 38714
rect 7262 38641 7368 38680
rect 7296 38607 7334 38641
rect 7262 38568 7368 38607
rect 7296 38534 7334 38568
rect 7262 38495 7368 38534
rect 7296 38461 7334 38495
rect 7262 38422 7368 38461
rect 7573 38680 7611 38714
rect 7539 38641 7645 38680
rect 7573 38607 7611 38641
rect 7539 38568 7645 38607
rect 7573 38534 7611 38568
rect 7539 38495 7645 38534
rect 7573 38461 7611 38495
rect 7539 38422 7645 38461
rect 7850 38680 7888 38714
rect 7816 38641 7922 38680
rect 7850 38607 7888 38641
rect 7816 38568 7922 38607
rect 7850 38534 7888 38568
rect 7816 38495 7922 38534
rect 7850 38461 7888 38495
rect 7816 38422 7922 38461
rect 3109 37368 3211 37380
rect 3663 37368 3765 37380
rect 4217 37368 4319 37380
rect 4771 37368 4873 37380
rect 5325 37368 5427 37380
rect 5879 37368 5981 37380
rect 6987 37368 7089 37380
rect 7539 37368 7645 37380
rect 3023 37031 3035 37065
rect 3073 37031 3108 37065
rect 3142 37031 3177 37065
rect 3215 37031 3246 37065
rect 3288 37031 3315 37065
rect 3361 37031 3384 37065
rect 3434 37031 3453 37065
rect 3507 37031 3522 37065
rect 3580 37031 3591 37065
rect 3653 37031 3660 37065
rect 3726 37031 3729 37065
rect 3763 37031 3765 37065
rect 3832 37031 3838 37065
rect 3901 37031 3911 37065
rect 3970 37031 3984 37065
rect 4039 37031 4057 37065
rect 4108 37031 4130 37065
rect 4177 37031 4203 37065
rect 4245 37031 4276 37065
rect 4313 37031 4347 37065
rect 4383 37031 4415 37065
rect 4456 37031 4483 37065
rect 4529 37031 4551 37065
rect 4602 37031 4619 37065
rect 4675 37031 4687 37065
rect 4748 37031 4755 37065
rect 4821 37031 4823 37065
rect 4857 37031 4860 37065
rect 4925 37031 4933 37065
rect 4993 37031 5006 37065
rect 5061 37031 5079 37065
rect 5129 37031 5152 37065
rect 5197 37031 5225 37065
rect 5265 37031 5298 37065
rect 5333 37031 5367 37065
rect 5405 37031 5435 37065
rect 5478 37031 5503 37065
rect 5551 37031 5571 37065
rect 5624 37031 5639 37065
rect 5697 37031 5707 37065
rect 5770 37031 5775 37065
rect 5877 37031 5882 37065
rect 5945 37031 5955 37065
rect 6013 37031 6027 37065
rect 6081 37031 6099 37065
rect 6149 37031 6171 37065
rect 6217 37031 6243 37065
rect 6285 37031 6315 37065
rect 6353 37031 6387 37065
rect 6421 37031 6455 37065
rect 6493 37031 6523 37065
rect 6565 37031 6591 37065
rect 6637 37031 6659 37065
rect 6709 37031 6727 37065
rect 6781 37031 6795 37065
rect 6853 37031 6863 37065
rect 6925 37031 6931 37065
rect 6997 37031 6999 37065
rect 7033 37031 7035 37065
rect 7101 37031 7107 37065
rect 7169 37031 7179 37065
rect 7237 37031 7251 37065
rect 7305 37031 7323 37065
rect 7373 37031 7395 37065
rect 7441 37031 7467 37065
rect 7509 37031 7539 37065
rect 7577 37031 7611 37065
rect 7645 37031 7679 37065
rect 7717 37031 7729 37065
rect 3109 36714 3211 36726
rect 3663 36714 3765 36726
rect 4217 36714 4319 36726
rect 4771 36714 4873 36726
rect 5325 36714 5427 36726
rect 5879 36714 5981 36726
rect 6987 36714 7089 36726
rect 7539 36714 7645 36726
rect 2864 36680 2902 36714
rect 2830 36641 2936 36680
rect 2864 36607 2902 36641
rect 2830 36568 2936 36607
rect 2864 36534 2902 36568
rect 2830 36495 2936 36534
rect 2864 36461 2902 36495
rect 2830 36422 2936 36461
rect 3141 36680 3179 36714
rect 3107 36641 3213 36680
rect 3141 36607 3179 36641
rect 3107 36568 3213 36607
rect 3141 36534 3179 36568
rect 3107 36495 3213 36534
rect 3141 36461 3179 36495
rect 3107 36422 3213 36461
rect 3418 36680 3456 36714
rect 3384 36641 3490 36680
rect 3418 36607 3456 36641
rect 3384 36568 3490 36607
rect 3418 36534 3456 36568
rect 3384 36495 3490 36534
rect 3418 36461 3456 36495
rect 3384 36422 3490 36461
rect 3695 36680 3733 36714
rect 3661 36641 3767 36680
rect 3695 36607 3733 36641
rect 3661 36568 3767 36607
rect 3695 36534 3733 36568
rect 3661 36495 3767 36534
rect 3695 36461 3733 36495
rect 3661 36422 3767 36461
rect 3972 36680 4010 36714
rect 3938 36641 4044 36680
rect 3972 36607 4010 36641
rect 3938 36568 4044 36607
rect 3972 36534 4010 36568
rect 3938 36495 4044 36534
rect 3972 36461 4010 36495
rect 3938 36422 4044 36461
rect 4249 36680 4287 36714
rect 4215 36641 4321 36680
rect 4249 36607 4287 36641
rect 4215 36568 4321 36607
rect 4249 36534 4287 36568
rect 4215 36495 4321 36534
rect 4249 36461 4287 36495
rect 4215 36422 4321 36461
rect 4526 36680 4564 36714
rect 4492 36641 4598 36680
rect 4526 36607 4564 36641
rect 4492 36568 4598 36607
rect 4526 36534 4564 36568
rect 4492 36495 4598 36534
rect 4526 36461 4564 36495
rect 4492 36422 4598 36461
rect 4803 36680 4841 36714
rect 4769 36641 4875 36680
rect 4803 36607 4841 36641
rect 4769 36568 4875 36607
rect 4803 36534 4841 36568
rect 4769 36495 4875 36534
rect 4803 36461 4841 36495
rect 4769 36422 4875 36461
rect 5080 36680 5118 36714
rect 5046 36641 5152 36680
rect 5080 36607 5118 36641
rect 5046 36568 5152 36607
rect 5080 36534 5118 36568
rect 5046 36495 5152 36534
rect 5080 36461 5118 36495
rect 5046 36422 5152 36461
rect 5357 36680 5395 36714
rect 5323 36641 5429 36680
rect 5357 36607 5395 36641
rect 5323 36568 5429 36607
rect 5357 36534 5395 36568
rect 5323 36495 5429 36534
rect 5357 36461 5395 36495
rect 5323 36422 5429 36461
rect 5634 36680 5672 36714
rect 5600 36641 5706 36680
rect 5634 36607 5672 36641
rect 5600 36568 5706 36607
rect 5634 36534 5672 36568
rect 5600 36495 5706 36534
rect 5634 36461 5672 36495
rect 5600 36422 5706 36461
rect 5911 36680 5949 36714
rect 5877 36641 5983 36680
rect 5911 36607 5949 36641
rect 5877 36568 5983 36607
rect 5911 36534 5949 36568
rect 5877 36495 5983 36534
rect 5911 36461 5949 36495
rect 5877 36422 5983 36461
rect 6188 36680 6226 36714
rect 6154 36641 6260 36680
rect 6188 36607 6226 36641
rect 6154 36568 6260 36607
rect 6188 36534 6226 36568
rect 6154 36495 6260 36534
rect 6188 36461 6226 36495
rect 6154 36422 6260 36461
rect 6465 36680 6503 36714
rect 6431 36641 6537 36680
rect 6465 36607 6503 36641
rect 6431 36568 6537 36607
rect 6465 36534 6503 36568
rect 6431 36495 6537 36534
rect 6465 36461 6503 36495
rect 6431 36422 6537 36461
rect 6742 36680 6780 36714
rect 6708 36641 6814 36680
rect 6742 36607 6780 36641
rect 6708 36568 6814 36607
rect 6742 36534 6780 36568
rect 6708 36495 6814 36534
rect 6742 36461 6780 36495
rect 6708 36422 6814 36461
rect 7019 36680 7057 36714
rect 6985 36641 7091 36680
rect 7019 36607 7057 36641
rect 6985 36568 7091 36607
rect 7019 36534 7057 36568
rect 6985 36495 7091 36534
rect 7019 36461 7057 36495
rect 6985 36422 7091 36461
rect 7296 36680 7334 36714
rect 7262 36641 7368 36680
rect 7296 36607 7334 36641
rect 7262 36568 7368 36607
rect 7296 36534 7334 36568
rect 7262 36495 7368 36534
rect 7296 36461 7334 36495
rect 7262 36422 7368 36461
rect 7573 36680 7611 36714
rect 7539 36641 7645 36680
rect 7573 36607 7611 36641
rect 7539 36568 7645 36607
rect 7573 36534 7611 36568
rect 7539 36495 7645 36534
rect 7573 36461 7611 36495
rect 7539 36422 7645 36461
rect 7850 36680 7888 36714
rect 7816 36641 7922 36680
rect 7850 36607 7888 36641
rect 7816 36568 7922 36607
rect 7850 36534 7888 36568
rect 7816 36495 7922 36534
rect 7850 36461 7888 36495
rect 7816 36422 7922 36461
rect 3109 35368 3211 35380
rect 3663 35368 3765 35380
rect 4217 35368 4319 35380
rect 4771 35368 4873 35380
rect 5325 35368 5427 35380
rect 5879 35368 5981 35380
rect 6987 35368 7089 35380
rect 7539 35368 7645 35380
rect 3023 35065 3035 35099
rect 3073 35065 3108 35099
rect 3142 35065 3177 35099
rect 3215 35065 3246 35099
rect 3288 35065 3315 35099
rect 3361 35065 3384 35099
rect 3434 35065 3453 35099
rect 3507 35065 3522 35099
rect 3580 35065 3591 35099
rect 3653 35065 3660 35099
rect 3726 35065 3729 35099
rect 3763 35065 3765 35099
rect 3832 35065 3838 35099
rect 3901 35065 3911 35099
rect 3970 35065 3984 35099
rect 4039 35065 4057 35099
rect 4108 35065 4130 35099
rect 4177 35065 4203 35099
rect 4245 35065 4276 35099
rect 4313 35065 4347 35099
rect 4383 35065 4415 35099
rect 4456 35065 4483 35099
rect 4529 35065 4551 35099
rect 4602 35065 4619 35099
rect 4675 35065 4687 35099
rect 4748 35065 4755 35099
rect 4821 35065 4823 35099
rect 4857 35065 4860 35099
rect 4925 35065 4933 35099
rect 4993 35065 5006 35099
rect 5061 35065 5079 35099
rect 5129 35065 5152 35099
rect 5197 35065 5225 35099
rect 5265 35065 5298 35099
rect 5333 35065 5367 35099
rect 5405 35065 5435 35099
rect 5478 35065 5503 35099
rect 5551 35065 5571 35099
rect 5624 35065 5639 35099
rect 5697 35065 5707 35099
rect 5770 35065 5775 35099
rect 5877 35065 5882 35099
rect 5945 35065 5955 35099
rect 6013 35065 6027 35099
rect 6081 35065 6099 35099
rect 6149 35065 6171 35099
rect 6217 35065 6243 35099
rect 6285 35065 6315 35099
rect 6353 35065 6387 35099
rect 6421 35065 6455 35099
rect 6493 35065 6523 35099
rect 6565 35065 6591 35099
rect 6637 35065 6659 35099
rect 6709 35065 6727 35099
rect 6781 35065 6795 35099
rect 6853 35065 6863 35099
rect 6925 35065 6931 35099
rect 6997 35065 6999 35099
rect 7033 35065 7035 35099
rect 7101 35065 7107 35099
rect 7169 35065 7179 35099
rect 7237 35065 7251 35099
rect 7305 35065 7323 35099
rect 7373 35065 7395 35099
rect 7441 35065 7467 35099
rect 7509 35065 7539 35099
rect 7577 35065 7611 35099
rect 7645 35065 7679 35099
rect 7717 35065 7729 35099
rect 3109 34714 3211 34726
rect 3663 34714 3765 34726
rect 4217 34714 4319 34726
rect 4771 34714 4873 34726
rect 5325 34714 5427 34726
rect 5879 34714 5981 34726
rect 6433 34714 6535 34726
rect 6987 34714 7089 34726
rect 7539 34714 7645 34726
rect 2864 34680 2902 34714
rect 2830 34641 2936 34680
rect 2864 34607 2902 34641
rect 2830 34568 2936 34607
rect 2864 34534 2902 34568
rect 2830 34495 2936 34534
rect 2864 34461 2902 34495
rect 2830 34422 2936 34461
rect 3141 34680 3179 34714
rect 3107 34641 3213 34680
rect 3141 34607 3179 34641
rect 3107 34568 3213 34607
rect 3141 34534 3179 34568
rect 3107 34495 3213 34534
rect 3141 34461 3179 34495
rect 3107 34422 3213 34461
rect 3418 34680 3456 34714
rect 3384 34641 3490 34680
rect 3418 34607 3456 34641
rect 3384 34568 3490 34607
rect 3418 34534 3456 34568
rect 3384 34495 3490 34534
rect 3418 34461 3456 34495
rect 3384 34422 3490 34461
rect 3695 34680 3733 34714
rect 3661 34641 3767 34680
rect 3695 34607 3733 34641
rect 3661 34568 3767 34607
rect 3695 34534 3733 34568
rect 3661 34495 3767 34534
rect 3695 34461 3733 34495
rect 3661 34422 3767 34461
rect 3972 34680 4010 34714
rect 3938 34641 4044 34680
rect 3972 34607 4010 34641
rect 3938 34568 4044 34607
rect 3972 34534 4010 34568
rect 3938 34495 4044 34534
rect 3972 34461 4010 34495
rect 3938 34422 4044 34461
rect 4249 34680 4287 34714
rect 4215 34641 4321 34680
rect 4249 34607 4287 34641
rect 4215 34568 4321 34607
rect 4249 34534 4287 34568
rect 4215 34495 4321 34534
rect 4249 34461 4287 34495
rect 4215 34422 4321 34461
rect 4526 34680 4564 34714
rect 4492 34641 4598 34680
rect 4526 34607 4564 34641
rect 4492 34568 4598 34607
rect 4526 34534 4564 34568
rect 4492 34495 4598 34534
rect 4526 34461 4564 34495
rect 4492 34422 4598 34461
rect 4803 34680 4841 34714
rect 4769 34641 4875 34680
rect 4803 34607 4841 34641
rect 4769 34568 4875 34607
rect 4803 34534 4841 34568
rect 4769 34495 4875 34534
rect 4803 34461 4841 34495
rect 4769 34422 4875 34461
rect 5080 34680 5118 34714
rect 5046 34641 5152 34680
rect 5080 34607 5118 34641
rect 5046 34568 5152 34607
rect 5080 34534 5118 34568
rect 5046 34495 5152 34534
rect 5080 34461 5118 34495
rect 5046 34422 5152 34461
rect 5357 34680 5395 34714
rect 5323 34641 5429 34680
rect 5357 34607 5395 34641
rect 5323 34568 5429 34607
rect 5357 34534 5395 34568
rect 5323 34495 5429 34534
rect 5357 34461 5395 34495
rect 5323 34422 5429 34461
rect 5634 34680 5672 34714
rect 5600 34641 5706 34680
rect 5634 34607 5672 34641
rect 5600 34568 5706 34607
rect 5634 34534 5672 34568
rect 5600 34495 5706 34534
rect 5634 34461 5672 34495
rect 5600 34422 5706 34461
rect 5911 34680 5949 34714
rect 5877 34641 5983 34680
rect 5911 34607 5949 34641
rect 5877 34568 5983 34607
rect 5911 34534 5949 34568
rect 5877 34495 5983 34534
rect 5911 34461 5949 34495
rect 5877 34422 5983 34461
rect 6188 34680 6226 34714
rect 6154 34641 6260 34680
rect 6188 34607 6226 34641
rect 6154 34568 6260 34607
rect 6188 34534 6226 34568
rect 6154 34495 6260 34534
rect 6188 34461 6226 34495
rect 6154 34422 6260 34461
rect 6465 34680 6503 34714
rect 6431 34641 6537 34680
rect 6465 34607 6503 34641
rect 6431 34568 6537 34607
rect 6465 34534 6503 34568
rect 6431 34495 6537 34534
rect 6465 34461 6503 34495
rect 6431 34422 6537 34461
rect 6742 34680 6780 34714
rect 6708 34641 6814 34680
rect 6742 34607 6780 34641
rect 6708 34568 6814 34607
rect 6742 34534 6780 34568
rect 6708 34495 6814 34534
rect 6742 34461 6780 34495
rect 6708 34422 6814 34461
rect 7019 34680 7057 34714
rect 6985 34641 7091 34680
rect 7019 34607 7057 34641
rect 6985 34568 7091 34607
rect 7019 34534 7057 34568
rect 6985 34495 7091 34534
rect 7019 34461 7057 34495
rect 6985 34422 7091 34461
rect 7296 34680 7334 34714
rect 7262 34641 7368 34680
rect 7296 34607 7334 34641
rect 7262 34568 7368 34607
rect 7296 34534 7334 34568
rect 7262 34495 7368 34534
rect 7296 34461 7334 34495
rect 7262 34422 7368 34461
rect 7573 34680 7611 34714
rect 7539 34641 7645 34680
rect 7573 34607 7611 34641
rect 7539 34568 7645 34607
rect 7573 34534 7611 34568
rect 7539 34495 7645 34534
rect 7573 34461 7611 34495
rect 7539 34422 7645 34461
rect 7850 34680 7888 34714
rect 7816 34641 7922 34680
rect 7850 34607 7888 34641
rect 7816 34568 7922 34607
rect 7850 34534 7888 34568
rect 7816 34495 7922 34534
rect 7850 34461 7888 34495
rect 7816 34422 7922 34461
rect 3109 33368 3211 33380
rect 3663 33368 3765 33380
rect 4217 33368 4319 33380
rect 4771 33368 4873 33380
rect 5325 33368 5427 33380
rect 5879 33368 5981 33380
rect 6433 33368 6535 33380
rect 6987 33368 7089 33380
rect 7539 33368 7645 33380
rect 3023 33066 3035 33100
rect 3073 33066 3108 33100
rect 3142 33066 3177 33100
rect 3215 33066 3246 33100
rect 3288 33066 3315 33100
rect 3361 33066 3384 33100
rect 3434 33066 3453 33100
rect 3507 33066 3522 33100
rect 3580 33066 3591 33100
rect 3653 33066 3660 33100
rect 3726 33066 3729 33100
rect 3763 33066 3765 33100
rect 3832 33066 3838 33100
rect 3901 33066 3911 33100
rect 3970 33066 3984 33100
rect 4039 33066 4057 33100
rect 4108 33066 4130 33100
rect 4177 33066 4203 33100
rect 4245 33066 4276 33100
rect 4313 33066 4347 33100
rect 4383 33066 4415 33100
rect 4456 33066 4483 33100
rect 4529 33066 4551 33100
rect 4602 33066 4619 33100
rect 4675 33066 4687 33100
rect 4748 33066 4755 33100
rect 4821 33066 4823 33100
rect 4857 33066 4860 33100
rect 4925 33066 4933 33100
rect 4993 33066 5006 33100
rect 5061 33066 5079 33100
rect 5129 33066 5152 33100
rect 5197 33066 5225 33100
rect 5265 33066 5298 33100
rect 5333 33066 5367 33100
rect 5405 33066 5435 33100
rect 5478 33066 5503 33100
rect 5551 33066 5571 33100
rect 5624 33066 5639 33100
rect 5697 33066 5707 33100
rect 5770 33066 5775 33100
rect 5877 33066 5882 33100
rect 5945 33066 5955 33100
rect 6013 33066 6027 33100
rect 6081 33066 6099 33100
rect 6149 33066 6171 33100
rect 6217 33066 6243 33100
rect 6285 33066 6315 33100
rect 6353 33066 6387 33100
rect 6421 33066 6455 33100
rect 6493 33066 6523 33100
rect 6565 33066 6591 33100
rect 6637 33066 6659 33100
rect 6709 33066 6727 33100
rect 6781 33066 6795 33100
rect 6853 33066 6863 33100
rect 6925 33066 6931 33100
rect 6997 33066 6999 33100
rect 7033 33066 7035 33100
rect 7101 33066 7107 33100
rect 7169 33066 7179 33100
rect 7237 33066 7251 33100
rect 7305 33066 7323 33100
rect 7373 33066 7395 33100
rect 7441 33066 7467 33100
rect 7509 33066 7539 33100
rect 7577 33066 7611 33100
rect 7645 33066 7679 33100
rect 7717 33066 7729 33100
rect 3109 32714 3211 32726
rect 3663 32714 3765 32726
rect 4217 32714 4319 32726
rect 4771 32714 4873 32726
rect 5325 32714 5427 32726
rect 5879 32714 5981 32726
rect 6433 32714 6535 32726
rect 6987 32714 7089 32726
rect 7539 32714 7645 32726
rect 2864 32680 2902 32714
rect 2830 32641 2936 32680
rect 2864 32607 2902 32641
rect 2830 32568 2936 32607
rect 2864 32534 2902 32568
rect 2830 32495 2936 32534
rect 2864 32461 2902 32495
rect 2830 32422 2936 32461
rect 3141 32680 3179 32714
rect 3107 32641 3213 32680
rect 3141 32607 3179 32641
rect 3107 32568 3213 32607
rect 3141 32534 3179 32568
rect 3107 32495 3213 32534
rect 3141 32461 3179 32495
rect 3107 32422 3213 32461
rect 3418 32680 3456 32714
rect 3384 32641 3490 32680
rect 3418 32607 3456 32641
rect 3384 32568 3490 32607
rect 3418 32534 3456 32568
rect 3384 32495 3490 32534
rect 3418 32461 3456 32495
rect 3384 32422 3490 32461
rect 3695 32680 3733 32714
rect 3661 32641 3767 32680
rect 3695 32607 3733 32641
rect 3661 32568 3767 32607
rect 3695 32534 3733 32568
rect 3661 32495 3767 32534
rect 3695 32461 3733 32495
rect 3661 32422 3767 32461
rect 3972 32680 4010 32714
rect 3938 32641 4044 32680
rect 3972 32607 4010 32641
rect 3938 32568 4044 32607
rect 3972 32534 4010 32568
rect 3938 32495 4044 32534
rect 3972 32461 4010 32495
rect 3938 32422 4044 32461
rect 4249 32680 4287 32714
rect 4215 32641 4321 32680
rect 4249 32607 4287 32641
rect 4215 32568 4321 32607
rect 4249 32534 4287 32568
rect 4215 32495 4321 32534
rect 4249 32461 4287 32495
rect 4215 32422 4321 32461
rect 4526 32680 4564 32714
rect 4492 32641 4598 32680
rect 4526 32607 4564 32641
rect 4492 32568 4598 32607
rect 4526 32534 4564 32568
rect 4492 32495 4598 32534
rect 4526 32461 4564 32495
rect 4492 32422 4598 32461
rect 4803 32680 4841 32714
rect 4769 32641 4875 32680
rect 4803 32607 4841 32641
rect 4769 32568 4875 32607
rect 4803 32534 4841 32568
rect 4769 32495 4875 32534
rect 4803 32461 4841 32495
rect 4769 32422 4875 32461
rect 5080 32680 5118 32714
rect 5046 32641 5152 32680
rect 5080 32607 5118 32641
rect 5046 32568 5152 32607
rect 5080 32534 5118 32568
rect 5046 32495 5152 32534
rect 5080 32461 5118 32495
rect 5046 32422 5152 32461
rect 5357 32680 5395 32714
rect 5323 32641 5429 32680
rect 5357 32607 5395 32641
rect 5323 32568 5429 32607
rect 5357 32534 5395 32568
rect 5323 32495 5429 32534
rect 5357 32461 5395 32495
rect 5323 32422 5429 32461
rect 5634 32680 5672 32714
rect 5600 32641 5706 32680
rect 5634 32607 5672 32641
rect 5600 32568 5706 32607
rect 5634 32534 5672 32568
rect 5600 32495 5706 32534
rect 5634 32461 5672 32495
rect 5600 32422 5706 32461
rect 5911 32680 5949 32714
rect 5877 32641 5983 32680
rect 5911 32607 5949 32641
rect 5877 32568 5983 32607
rect 5911 32534 5949 32568
rect 5877 32495 5983 32534
rect 5911 32461 5949 32495
rect 5877 32422 5983 32461
rect 6188 32680 6226 32714
rect 6154 32641 6260 32680
rect 6188 32607 6226 32641
rect 6154 32568 6260 32607
rect 6188 32534 6226 32568
rect 6154 32495 6260 32534
rect 6188 32461 6226 32495
rect 6154 32422 6260 32461
rect 6465 32680 6503 32714
rect 6431 32641 6537 32680
rect 6465 32607 6503 32641
rect 6431 32568 6537 32607
rect 6465 32534 6503 32568
rect 6431 32495 6537 32534
rect 6465 32461 6503 32495
rect 6431 32422 6537 32461
rect 6742 32680 6780 32714
rect 6708 32641 6814 32680
rect 6742 32607 6780 32641
rect 6708 32568 6814 32607
rect 6742 32534 6780 32568
rect 6708 32495 6814 32534
rect 6742 32461 6780 32495
rect 6708 32422 6814 32461
rect 7019 32680 7057 32714
rect 6985 32641 7091 32680
rect 7019 32607 7057 32641
rect 6985 32568 7091 32607
rect 7019 32534 7057 32568
rect 6985 32495 7091 32534
rect 7019 32461 7057 32495
rect 6985 32422 7091 32461
rect 7296 32680 7334 32714
rect 7262 32641 7368 32680
rect 7296 32607 7334 32641
rect 7262 32568 7368 32607
rect 7296 32534 7334 32568
rect 7262 32495 7368 32534
rect 7296 32461 7334 32495
rect 7262 32422 7368 32461
rect 7573 32680 7611 32714
rect 7539 32641 7645 32680
rect 7573 32607 7611 32641
rect 7539 32568 7645 32607
rect 7573 32534 7611 32568
rect 7539 32495 7645 32534
rect 7573 32461 7611 32495
rect 7539 32422 7645 32461
rect 7850 32680 7888 32714
rect 7816 32641 7922 32680
rect 7850 32607 7888 32641
rect 7816 32568 7922 32607
rect 7850 32534 7888 32568
rect 7816 32495 7922 32534
rect 7850 32461 7888 32495
rect 7816 32422 7922 32461
rect 3109 31368 3211 31380
rect 3663 31368 3765 31380
rect 4217 31368 4319 31380
rect 4771 31368 4873 31380
rect 5325 31368 5427 31380
rect 5879 31368 5981 31380
rect 6433 31368 6535 31380
rect 6987 31368 7089 31380
rect 7539 31368 7645 31380
rect 3023 31043 3035 31077
rect 3073 31043 3108 31077
rect 3142 31043 3177 31077
rect 3215 31043 3246 31077
rect 3288 31043 3315 31077
rect 3361 31043 3384 31077
rect 3434 31043 3453 31077
rect 3507 31043 3522 31077
rect 3580 31043 3591 31077
rect 3653 31043 3660 31077
rect 3726 31043 3729 31077
rect 3763 31043 3765 31077
rect 3832 31043 3838 31077
rect 3901 31043 3911 31077
rect 3970 31043 3984 31077
rect 4039 31043 4057 31077
rect 4108 31043 4130 31077
rect 4177 31043 4203 31077
rect 4245 31043 4276 31077
rect 4313 31043 4347 31077
rect 4383 31043 4415 31077
rect 4456 31043 4483 31077
rect 4529 31043 4551 31077
rect 4602 31043 4619 31077
rect 4675 31043 4687 31077
rect 4748 31043 4755 31077
rect 4821 31043 4823 31077
rect 4857 31043 4860 31077
rect 4925 31043 4933 31077
rect 4993 31043 5006 31077
rect 5061 31043 5079 31077
rect 5129 31043 5152 31077
rect 5197 31043 5225 31077
rect 5265 31043 5298 31077
rect 5333 31043 5367 31077
rect 5405 31043 5435 31077
rect 5478 31043 5503 31077
rect 5551 31043 5571 31077
rect 5624 31043 5639 31077
rect 5697 31043 5707 31077
rect 5770 31043 5775 31077
rect 5877 31043 5882 31077
rect 5945 31043 5955 31077
rect 6013 31043 6027 31077
rect 6081 31043 6099 31077
rect 6149 31043 6171 31077
rect 6217 31043 6243 31077
rect 6285 31043 6315 31077
rect 6353 31043 6387 31077
rect 6421 31043 6455 31077
rect 6493 31043 6523 31077
rect 6565 31043 6591 31077
rect 6637 31043 6659 31077
rect 6709 31043 6727 31077
rect 6781 31043 6795 31077
rect 6853 31043 6863 31077
rect 6925 31043 6931 31077
rect 6997 31043 6999 31077
rect 7033 31043 7035 31077
rect 7101 31043 7107 31077
rect 7169 31043 7179 31077
rect 7237 31043 7251 31077
rect 7305 31043 7323 31077
rect 7373 31043 7395 31077
rect 7441 31043 7467 31077
rect 7509 31043 7539 31077
rect 7577 31043 7611 31077
rect 7645 31043 7679 31077
rect 7717 31043 7729 31077
rect 3109 30714 3211 30726
rect 3663 30714 3765 30726
rect 4217 30714 4319 30726
rect 4771 30714 4873 30726
rect 5325 30714 5427 30726
rect 5879 30714 5981 30726
rect 6433 30714 6535 30726
rect 6987 30714 7089 30726
rect 7539 30714 7645 30726
rect 2864 30680 2902 30714
rect 2830 30641 2936 30680
rect 2864 30607 2902 30641
rect 2830 30568 2936 30607
rect 2864 30534 2902 30568
rect 2830 30495 2936 30534
rect 2864 30461 2902 30495
rect 2830 30422 2936 30461
rect 3141 30680 3179 30714
rect 3107 30641 3213 30680
rect 3141 30607 3179 30641
rect 3107 30568 3213 30607
rect 3141 30534 3179 30568
rect 3107 30495 3213 30534
rect 3141 30461 3179 30495
rect 3107 30422 3213 30461
rect 3418 30680 3456 30714
rect 3384 30641 3490 30680
rect 3418 30607 3456 30641
rect 3384 30568 3490 30607
rect 3418 30534 3456 30568
rect 3384 30495 3490 30534
rect 3418 30461 3456 30495
rect 3384 30422 3490 30461
rect 3695 30680 3733 30714
rect 3661 30641 3767 30680
rect 3695 30607 3733 30641
rect 3661 30568 3767 30607
rect 3695 30534 3733 30568
rect 3661 30495 3767 30534
rect 3695 30461 3733 30495
rect 3661 30422 3767 30461
rect 3972 30680 4010 30714
rect 3938 30641 4044 30680
rect 3972 30607 4010 30641
rect 3938 30568 4044 30607
rect 3972 30534 4010 30568
rect 3938 30495 4044 30534
rect 3972 30461 4010 30495
rect 3938 30422 4044 30461
rect 4249 30680 4287 30714
rect 4215 30641 4321 30680
rect 4249 30607 4287 30641
rect 4215 30568 4321 30607
rect 4249 30534 4287 30568
rect 4215 30495 4321 30534
rect 4249 30461 4287 30495
rect 4215 30422 4321 30461
rect 4526 30680 4564 30714
rect 4492 30641 4598 30680
rect 4526 30607 4564 30641
rect 4492 30568 4598 30607
rect 4526 30534 4564 30568
rect 4492 30495 4598 30534
rect 4526 30461 4564 30495
rect 4492 30422 4598 30461
rect 4803 30680 4841 30714
rect 4769 30641 4875 30680
rect 4803 30607 4841 30641
rect 4769 30568 4875 30607
rect 4803 30534 4841 30568
rect 4769 30495 4875 30534
rect 4803 30461 4841 30495
rect 4769 30422 4875 30461
rect 5080 30680 5118 30714
rect 5046 30641 5152 30680
rect 5080 30607 5118 30641
rect 5046 30568 5152 30607
rect 5080 30534 5118 30568
rect 5046 30495 5152 30534
rect 5080 30461 5118 30495
rect 5046 30422 5152 30461
rect 5357 30680 5395 30714
rect 5323 30641 5429 30680
rect 5357 30607 5395 30641
rect 5323 30568 5429 30607
rect 5357 30534 5395 30568
rect 5323 30495 5429 30534
rect 5357 30461 5395 30495
rect 5323 30422 5429 30461
rect 5634 30680 5672 30714
rect 5600 30641 5706 30680
rect 5634 30607 5672 30641
rect 5600 30568 5706 30607
rect 5634 30534 5672 30568
rect 5600 30495 5706 30534
rect 5634 30461 5672 30495
rect 5600 30422 5706 30461
rect 5911 30680 5949 30714
rect 5877 30641 5983 30680
rect 5911 30607 5949 30641
rect 5877 30568 5983 30607
rect 5911 30534 5949 30568
rect 5877 30495 5983 30534
rect 5911 30461 5949 30495
rect 5877 30422 5983 30461
rect 6188 30680 6226 30714
rect 6154 30641 6260 30680
rect 6188 30607 6226 30641
rect 6154 30568 6260 30607
rect 6188 30534 6226 30568
rect 6154 30495 6260 30534
rect 6188 30461 6226 30495
rect 6154 30422 6260 30461
rect 6465 30680 6503 30714
rect 6431 30641 6537 30680
rect 6465 30607 6503 30641
rect 6431 30568 6537 30607
rect 6465 30534 6503 30568
rect 6431 30495 6537 30534
rect 6465 30461 6503 30495
rect 6431 30422 6537 30461
rect 6742 30680 6780 30714
rect 6708 30641 6814 30680
rect 6742 30607 6780 30641
rect 6708 30568 6814 30607
rect 6742 30534 6780 30568
rect 6708 30495 6814 30534
rect 6742 30461 6780 30495
rect 6708 30422 6814 30461
rect 7019 30680 7057 30714
rect 6985 30641 7091 30680
rect 7019 30607 7057 30641
rect 6985 30568 7091 30607
rect 7019 30534 7057 30568
rect 6985 30495 7091 30534
rect 7019 30461 7057 30495
rect 6985 30422 7091 30461
rect 7296 30680 7334 30714
rect 7262 30641 7368 30680
rect 7296 30607 7334 30641
rect 7262 30568 7368 30607
rect 7296 30534 7334 30568
rect 7262 30495 7368 30534
rect 7296 30461 7334 30495
rect 7262 30422 7368 30461
rect 7573 30680 7611 30714
rect 7539 30641 7645 30680
rect 7573 30607 7611 30641
rect 7539 30568 7645 30607
rect 7573 30534 7611 30568
rect 7539 30495 7645 30534
rect 7573 30461 7611 30495
rect 7539 30422 7645 30461
rect 7850 30680 7888 30714
rect 7816 30641 7922 30680
rect 7850 30607 7888 30641
rect 7816 30568 7922 30607
rect 7850 30534 7888 30568
rect 7816 30495 7922 30534
rect 7850 30461 7888 30495
rect 7816 30422 7922 30461
rect 3109 29368 3211 29380
rect 3663 29368 3765 29380
rect 4217 29368 4319 29380
rect 4771 29368 4873 29380
rect 5325 29368 5427 29380
rect 5879 29368 5981 29380
rect 6433 29368 6535 29380
rect 6987 29368 7089 29380
rect 7539 29368 7645 29380
rect 3023 29216 3035 29250
rect 3073 29216 3108 29250
rect 3142 29216 3177 29250
rect 3215 29216 3246 29250
rect 3288 29216 3315 29250
rect 3361 29216 3384 29250
rect 3434 29216 3453 29250
rect 3507 29216 3522 29250
rect 3580 29216 3591 29250
rect 3653 29216 3660 29250
rect 3726 29216 3729 29250
rect 3763 29216 3765 29250
rect 3832 29216 3838 29250
rect 3901 29216 3911 29250
rect 3970 29216 3984 29250
rect 4039 29216 4057 29250
rect 4108 29216 4130 29250
rect 4177 29216 4203 29250
rect 4245 29216 4276 29250
rect 4313 29216 4347 29250
rect 4383 29216 4415 29250
rect 4456 29216 4483 29250
rect 4529 29216 4551 29250
rect 4602 29216 4619 29250
rect 4675 29216 4687 29250
rect 4748 29216 4755 29250
rect 4821 29216 4823 29250
rect 4857 29216 4860 29250
rect 4925 29216 4933 29250
rect 4993 29216 5006 29250
rect 5061 29216 5079 29250
rect 5129 29216 5152 29250
rect 5197 29216 5225 29250
rect 5265 29216 5298 29250
rect 5333 29216 5367 29250
rect 5405 29216 5435 29250
rect 5478 29216 5503 29250
rect 5551 29216 5571 29250
rect 5624 29216 5639 29250
rect 5697 29216 5707 29250
rect 5770 29216 5775 29250
rect 5877 29216 5882 29250
rect 5945 29216 5955 29250
rect 6013 29216 6027 29250
rect 6081 29216 6099 29250
rect 6149 29216 6171 29250
rect 6217 29216 6243 29250
rect 6285 29216 6315 29250
rect 6353 29216 6387 29250
rect 6421 29216 6455 29250
rect 6493 29216 6523 29250
rect 6565 29216 6591 29250
rect 6637 29216 6659 29250
rect 6709 29216 6727 29250
rect 6781 29216 6795 29250
rect 6853 29216 6863 29250
rect 6925 29216 6931 29250
rect 6997 29216 6999 29250
rect 7033 29216 7035 29250
rect 7101 29216 7107 29250
rect 7169 29216 7179 29250
rect 7237 29216 7251 29250
rect 7305 29216 7323 29250
rect 7373 29216 7395 29250
rect 7441 29216 7467 29250
rect 7509 29216 7539 29250
rect 7577 29216 7611 29250
rect 7645 29216 7679 29250
rect 7717 29216 7729 29250
rect 2704 28965 4692 28982
rect 2648 18563 2663 28965
rect 4569 28958 4692 28965
rect 4569 28924 4647 28958
rect 4681 28924 4692 28958
rect 4569 28822 4692 28924
rect 4569 28788 4647 28822
rect 4681 28788 4692 28822
rect 4569 28686 4692 28788
rect 5325 28714 5427 28726
rect 5879 28714 5981 28726
rect 6433 28714 6535 28726
rect 6987 28714 7089 28726
rect 7539 28714 7645 28726
rect 4569 28652 4647 28686
rect 4681 28652 4692 28686
rect 4569 28550 4692 28652
rect 4569 28516 4647 28550
rect 4681 28516 4692 28550
rect 4569 28414 4692 28516
rect 4569 28380 4647 28414
rect 4681 28380 4692 28414
rect 4569 28278 4692 28380
rect 4569 28244 4647 28278
rect 4681 28244 4692 28278
rect 4569 28142 4692 28244
rect 4569 28108 4647 28142
rect 4681 28108 4692 28142
rect 4569 28006 4692 28108
rect 4569 27972 4647 28006
rect 4681 27972 4692 28006
rect 4569 27870 4692 27972
rect 4569 27836 4647 27870
rect 4681 27836 4692 27870
rect 4569 27734 4692 27836
rect 4569 27700 4647 27734
rect 4681 27700 4692 27734
rect 4569 27598 4692 27700
rect 4569 27564 4647 27598
rect 4681 27564 4692 27598
rect 4569 27462 4692 27564
rect 4569 27428 4647 27462
rect 4681 27428 4692 27462
rect 4569 27326 4692 27428
rect 5080 28680 5118 28714
rect 5046 28641 5152 28680
rect 5080 28607 5118 28641
rect 5046 28568 5152 28607
rect 5080 28534 5118 28568
rect 5046 28495 5152 28534
rect 5080 28461 5118 28495
rect 5046 28422 5152 28461
rect 5357 28680 5395 28714
rect 5323 28641 5429 28680
rect 5357 28607 5395 28641
rect 5323 28568 5429 28607
rect 5357 28534 5395 28568
rect 5323 28495 5429 28534
rect 5357 28461 5395 28495
rect 5323 28422 5429 28461
rect 5634 28680 5672 28714
rect 5600 28641 5706 28680
rect 5634 28607 5672 28641
rect 5600 28568 5706 28607
rect 5634 28534 5672 28568
rect 5600 28495 5706 28534
rect 5634 28461 5672 28495
rect 5600 28422 5706 28461
rect 5911 28680 5949 28714
rect 5877 28641 5983 28680
rect 5911 28607 5949 28641
rect 5877 28568 5983 28607
rect 5911 28534 5949 28568
rect 5877 28495 5983 28534
rect 5911 28461 5949 28495
rect 5877 28422 5983 28461
rect 6188 28680 6226 28714
rect 6154 28641 6260 28680
rect 6188 28607 6226 28641
rect 6154 28568 6260 28607
rect 6188 28534 6226 28568
rect 6154 28495 6260 28534
rect 6188 28461 6226 28495
rect 6154 28422 6260 28461
rect 6465 28680 6503 28714
rect 6431 28641 6537 28680
rect 6465 28607 6503 28641
rect 6431 28568 6537 28607
rect 6465 28534 6503 28568
rect 6431 28495 6537 28534
rect 6465 28461 6503 28495
rect 6431 28422 6537 28461
rect 6742 28680 6780 28714
rect 6708 28641 6814 28680
rect 6742 28607 6780 28641
rect 6708 28568 6814 28607
rect 6742 28534 6780 28568
rect 6708 28495 6814 28534
rect 6742 28461 6780 28495
rect 6708 28422 6814 28461
rect 7019 28680 7057 28714
rect 6985 28641 7091 28680
rect 7019 28607 7057 28641
rect 6985 28568 7091 28607
rect 7019 28534 7057 28568
rect 6985 28495 7091 28534
rect 7019 28461 7057 28495
rect 6985 28422 7091 28461
rect 7296 28680 7334 28714
rect 7262 28641 7368 28680
rect 7296 28607 7334 28641
rect 7262 28568 7368 28607
rect 7296 28534 7334 28568
rect 7262 28495 7368 28534
rect 7296 28461 7334 28495
rect 7262 28422 7368 28461
rect 7573 28680 7611 28714
rect 7539 28641 7645 28680
rect 7573 28607 7611 28641
rect 7539 28568 7645 28607
rect 7573 28534 7611 28568
rect 7539 28495 7645 28534
rect 7573 28461 7611 28495
rect 7539 28422 7645 28461
rect 7850 28680 7888 28714
rect 7816 28641 7922 28680
rect 7850 28607 7888 28641
rect 7816 28568 7922 28607
rect 7850 28534 7888 28568
rect 7816 28495 7922 28534
rect 7850 28461 7888 28495
rect 7816 28422 7922 28461
rect 5325 27368 5427 27380
rect 5879 27368 5981 27380
rect 6433 27368 6535 27380
rect 6987 27368 7089 27380
rect 7539 27368 7645 27380
rect 4569 27292 4647 27326
rect 4681 27292 4692 27326
rect 4569 27190 4692 27292
rect 4569 27156 4647 27190
rect 4681 27156 4692 27190
rect 4569 27054 4692 27156
rect 5239 27071 5251 27105
rect 5289 27071 5325 27105
rect 5360 27071 5395 27105
rect 5435 27071 5465 27105
rect 5510 27071 5535 27105
rect 5585 27071 5605 27105
rect 5660 27071 5675 27105
rect 5735 27071 5745 27105
rect 5810 27071 5815 27105
rect 5849 27071 5851 27105
rect 5919 27071 5926 27105
rect 5988 27071 6001 27105
rect 6057 27071 6076 27105
rect 6126 27071 6151 27105
rect 6195 27071 6225 27105
rect 6264 27071 6299 27105
rect 6333 27071 6368 27105
rect 6407 27071 6437 27105
rect 6481 27071 6506 27105
rect 6555 27071 6575 27105
rect 6629 27071 6644 27105
rect 6703 27071 6713 27105
rect 6777 27071 6782 27105
rect 6816 27071 6817 27105
rect 6885 27071 6891 27105
rect 6954 27071 6989 27105
rect 7023 27071 7058 27105
rect 7092 27071 7127 27105
rect 7161 27071 7196 27105
rect 7230 27071 7265 27105
rect 7299 27071 7334 27105
rect 7368 27071 7403 27105
rect 7437 27071 7472 27105
rect 7506 27071 7541 27105
rect 7575 27071 7610 27105
rect 7644 27071 7679 27105
rect 7713 27071 7729 27105
rect 4569 27020 4647 27054
rect 4681 27020 4692 27054
rect 4569 26918 4692 27020
rect 4569 26884 4647 26918
rect 4681 26884 4692 26918
rect 4569 26782 4692 26884
rect 4569 26748 4647 26782
rect 4681 26748 4692 26782
rect 4569 26646 4692 26748
rect 5325 26714 5427 26726
rect 5879 26714 5981 26726
rect 6433 26714 6535 26726
rect 6987 26714 7089 26726
rect 7539 26714 7645 26726
rect 4569 26612 4647 26646
rect 4681 26612 4692 26646
rect 4569 26510 4692 26612
rect 4569 26476 4647 26510
rect 4681 26476 4692 26510
rect 4569 26374 4692 26476
rect 4569 26340 4647 26374
rect 4681 26340 4692 26374
rect 4569 26238 4692 26340
rect 4569 26204 4647 26238
rect 4681 26204 4692 26238
rect 4569 26102 4692 26204
rect 4569 26068 4647 26102
rect 4681 26068 4692 26102
rect 4569 25966 4692 26068
rect 4569 25932 4647 25966
rect 4681 25932 4692 25966
rect 4569 25830 4692 25932
rect 4569 25796 4647 25830
rect 4681 25796 4692 25830
rect 4569 25694 4692 25796
rect 4569 25660 4647 25694
rect 4681 25660 4692 25694
rect 4569 25558 4692 25660
rect 4569 25524 4647 25558
rect 4681 25524 4692 25558
rect 4569 25422 4692 25524
rect 4569 25388 4647 25422
rect 4681 25388 4692 25422
rect 4569 25286 4692 25388
rect 5080 26680 5118 26714
rect 5046 26641 5152 26680
rect 5080 26607 5118 26641
rect 5046 26568 5152 26607
rect 5080 26534 5118 26568
rect 5046 26495 5152 26534
rect 5080 26461 5118 26495
rect 5046 26422 5152 26461
rect 5357 26680 5395 26714
rect 5323 26641 5429 26680
rect 5357 26607 5395 26641
rect 5323 26568 5429 26607
rect 5357 26534 5395 26568
rect 5323 26495 5429 26534
rect 5357 26461 5395 26495
rect 5323 26422 5429 26461
rect 5634 26680 5672 26714
rect 5600 26641 5706 26680
rect 5634 26607 5672 26641
rect 5600 26568 5706 26607
rect 5634 26534 5672 26568
rect 5600 26495 5706 26534
rect 5634 26461 5672 26495
rect 5600 26422 5706 26461
rect 5911 26680 5949 26714
rect 5877 26641 5983 26680
rect 5911 26607 5949 26641
rect 5877 26568 5983 26607
rect 5911 26534 5949 26568
rect 5877 26495 5983 26534
rect 5911 26461 5949 26495
rect 5877 26422 5983 26461
rect 6188 26680 6226 26714
rect 6154 26641 6260 26680
rect 6188 26607 6226 26641
rect 6154 26568 6260 26607
rect 6188 26534 6226 26568
rect 6154 26495 6260 26534
rect 6188 26461 6226 26495
rect 6154 26422 6260 26461
rect 6465 26680 6503 26714
rect 6431 26641 6537 26680
rect 6465 26607 6503 26641
rect 6431 26568 6537 26607
rect 6465 26534 6503 26568
rect 6431 26495 6537 26534
rect 6465 26461 6503 26495
rect 6431 26422 6537 26461
rect 6742 26680 6780 26714
rect 6708 26641 6814 26680
rect 6742 26607 6780 26641
rect 6708 26568 6814 26607
rect 6742 26534 6780 26568
rect 6708 26495 6814 26534
rect 6742 26461 6780 26495
rect 6708 26422 6814 26461
rect 7019 26680 7057 26714
rect 6985 26641 7091 26680
rect 7019 26607 7057 26641
rect 6985 26568 7091 26607
rect 7019 26534 7057 26568
rect 6985 26495 7091 26534
rect 7019 26461 7057 26495
rect 6985 26422 7091 26461
rect 7296 26680 7334 26714
rect 7262 26641 7368 26680
rect 7296 26607 7334 26641
rect 7262 26568 7368 26607
rect 7296 26534 7334 26568
rect 7262 26495 7368 26534
rect 7296 26461 7334 26495
rect 7262 26422 7368 26461
rect 7573 26680 7611 26714
rect 7539 26641 7645 26680
rect 7573 26607 7611 26641
rect 7539 26568 7645 26607
rect 7573 26534 7611 26568
rect 7539 26495 7645 26534
rect 7573 26461 7611 26495
rect 7539 26422 7645 26461
rect 7850 26680 7888 26714
rect 7816 26641 7922 26680
rect 7850 26607 7888 26641
rect 7816 26568 7922 26607
rect 7850 26534 7888 26568
rect 7816 26495 7922 26534
rect 7850 26461 7888 26495
rect 7816 26422 7922 26461
rect 5325 25368 5427 25380
rect 5879 25368 5981 25380
rect 6433 25368 6535 25380
rect 6987 25368 7089 25380
rect 7539 25368 7645 25380
rect 4569 25252 4647 25286
rect 4681 25252 4692 25286
rect 4569 25149 4692 25252
rect 4569 25115 4647 25149
rect 4681 25115 4692 25149
rect 4569 25012 4692 25115
rect 5239 25078 5251 25112
rect 5289 25078 5325 25112
rect 5359 25078 5395 25112
rect 5433 25078 5465 25112
rect 5507 25078 5535 25112
rect 5581 25078 5605 25112
rect 5655 25078 5675 25112
rect 5729 25078 5745 25112
rect 5803 25078 5815 25112
rect 5877 25078 5885 25112
rect 5951 25078 5954 25112
rect 5988 25078 5991 25112
rect 6057 25078 6065 25112
rect 6126 25078 6139 25112
rect 6195 25078 6213 25112
rect 6264 25078 6287 25112
rect 6333 25078 6361 25112
rect 6402 25078 6435 25112
rect 6471 25078 6506 25112
rect 6543 25078 6575 25112
rect 6617 25078 6644 25112
rect 6691 25078 6713 25112
rect 6765 25078 6782 25112
rect 6839 25078 6851 25112
rect 6913 25078 6920 25112
rect 6987 25078 6989 25112
rect 7023 25078 7026 25112
rect 7092 25078 7099 25112
rect 7161 25078 7172 25112
rect 7230 25078 7245 25112
rect 7299 25078 7318 25112
rect 7368 25078 7391 25112
rect 7437 25078 7464 25112
rect 7506 25078 7537 25112
rect 7575 25078 7610 25112
rect 7644 25078 7679 25112
rect 7717 25078 7729 25112
rect 4569 24978 4647 25012
rect 4681 24978 4692 25012
rect 4569 24875 4692 24978
rect 4569 24841 4647 24875
rect 4681 24841 4692 24875
rect 4569 24738 4692 24841
rect 4569 24704 4647 24738
rect 4681 24704 4692 24738
rect 5325 24714 5427 24726
rect 5879 24714 5981 24726
rect 6433 24714 6535 24726
rect 6987 24714 7089 24726
rect 7539 24714 7645 24726
rect 4569 24601 4692 24704
rect 4569 24567 4647 24601
rect 4681 24567 4692 24601
rect 4569 24464 4692 24567
rect 4569 24430 4647 24464
rect 4681 24430 4692 24464
rect 4569 24327 4692 24430
rect 4569 24293 4647 24327
rect 4681 24293 4692 24327
rect 4569 24190 4692 24293
rect 4569 24156 4647 24190
rect 4681 24156 4692 24190
rect 4569 24053 4692 24156
rect 4569 24019 4647 24053
rect 4681 24019 4692 24053
rect 4569 23916 4692 24019
rect 4569 23882 4647 23916
rect 4681 23882 4692 23916
rect 4569 23779 4692 23882
rect 4569 23745 4647 23779
rect 4681 23745 4692 23779
rect 4569 23642 4692 23745
rect 4569 23608 4647 23642
rect 4681 23608 4692 23642
rect 4569 23505 4692 23608
rect 4569 23471 4647 23505
rect 4681 23471 4692 23505
rect 4569 23368 4692 23471
rect 5080 24680 5118 24714
rect 5046 24641 5152 24680
rect 5080 24607 5118 24641
rect 5046 24568 5152 24607
rect 5080 24534 5118 24568
rect 5046 24495 5152 24534
rect 5080 24461 5118 24495
rect 5046 24422 5152 24461
rect 5357 24680 5395 24714
rect 5323 24641 5429 24680
rect 5357 24607 5395 24641
rect 5323 24568 5429 24607
rect 5357 24534 5395 24568
rect 5323 24495 5429 24534
rect 5357 24461 5395 24495
rect 5323 24422 5429 24461
rect 5634 24680 5672 24714
rect 5600 24641 5706 24680
rect 5634 24607 5672 24641
rect 5600 24568 5706 24607
rect 5634 24534 5672 24568
rect 5600 24495 5706 24534
rect 5634 24461 5672 24495
rect 5600 24422 5706 24461
rect 5911 24680 5949 24714
rect 5877 24641 5983 24680
rect 5911 24607 5949 24641
rect 5877 24568 5983 24607
rect 5911 24534 5949 24568
rect 5877 24495 5983 24534
rect 5911 24461 5949 24495
rect 5877 24422 5983 24461
rect 6188 24680 6226 24714
rect 6154 24641 6260 24680
rect 6188 24607 6226 24641
rect 6154 24568 6260 24607
rect 6188 24534 6226 24568
rect 6154 24495 6260 24534
rect 6188 24461 6226 24495
rect 6154 24422 6260 24461
rect 6465 24680 6503 24714
rect 6431 24641 6537 24680
rect 6465 24607 6503 24641
rect 6431 24568 6537 24607
rect 6465 24534 6503 24568
rect 6431 24495 6537 24534
rect 6465 24461 6503 24495
rect 6431 24422 6537 24461
rect 6742 24680 6780 24714
rect 6708 24641 6814 24680
rect 6742 24607 6780 24641
rect 6708 24568 6814 24607
rect 6742 24534 6780 24568
rect 6708 24495 6814 24534
rect 6742 24461 6780 24495
rect 6708 24422 6814 24461
rect 7019 24680 7057 24714
rect 6985 24641 7091 24680
rect 7019 24607 7057 24641
rect 6985 24568 7091 24607
rect 7019 24534 7057 24568
rect 6985 24495 7091 24534
rect 7019 24461 7057 24495
rect 6985 24422 7091 24461
rect 7296 24680 7334 24714
rect 7262 24641 7368 24680
rect 7296 24607 7334 24641
rect 7262 24568 7368 24607
rect 7296 24534 7334 24568
rect 7262 24495 7368 24534
rect 7296 24461 7334 24495
rect 7262 24422 7368 24461
rect 7573 24680 7611 24714
rect 7539 24641 7645 24680
rect 7573 24607 7611 24641
rect 7539 24568 7645 24607
rect 7573 24534 7611 24568
rect 7539 24495 7645 24534
rect 7573 24461 7611 24495
rect 7539 24422 7645 24461
rect 7850 24680 7888 24714
rect 7816 24641 7922 24680
rect 7850 24607 7888 24641
rect 7816 24568 7922 24607
rect 7850 24534 7888 24568
rect 7816 24495 7922 24534
rect 7850 24461 7888 24495
rect 7816 24422 7922 24461
rect 5325 23368 5427 23380
rect 5879 23368 5981 23380
rect 6433 23368 6535 23380
rect 6987 23368 7089 23380
rect 7539 23368 7645 23380
rect 4569 23334 4647 23368
rect 4681 23334 4692 23368
rect 4569 23231 4692 23334
rect 4569 23197 4647 23231
rect 4681 23197 4692 23231
rect 4569 23094 4692 23197
rect 4569 23060 4647 23094
rect 4681 23060 4692 23094
rect 5239 23090 5251 23124
rect 5289 23090 5325 23124
rect 5359 23090 5395 23124
rect 5433 23090 5465 23124
rect 5507 23090 5535 23124
rect 5581 23090 5605 23124
rect 5655 23090 5675 23124
rect 5729 23090 5745 23124
rect 5803 23090 5815 23124
rect 5877 23090 5885 23124
rect 5951 23090 5954 23124
rect 5988 23090 5991 23124
rect 6057 23090 6065 23124
rect 6126 23090 6139 23124
rect 6195 23090 6213 23124
rect 6264 23090 6287 23124
rect 6333 23090 6361 23124
rect 6402 23090 6435 23124
rect 6471 23090 6506 23124
rect 6543 23090 6575 23124
rect 6617 23090 6644 23124
rect 6691 23090 6713 23124
rect 6765 23090 6782 23124
rect 6839 23090 6851 23124
rect 6913 23090 6920 23124
rect 6987 23090 6989 23124
rect 7023 23090 7026 23124
rect 7092 23090 7099 23124
rect 7161 23090 7172 23124
rect 7230 23090 7245 23124
rect 7299 23090 7318 23124
rect 7368 23090 7391 23124
rect 7437 23090 7464 23124
rect 7506 23090 7537 23124
rect 7575 23090 7610 23124
rect 7644 23090 7679 23124
rect 7717 23090 7729 23124
rect 4569 22957 4692 23060
rect 4569 22923 4647 22957
rect 4681 22923 4692 22957
rect 4569 22820 4692 22923
rect 4569 22786 4647 22820
rect 4681 22786 4692 22820
rect 4569 22683 4692 22786
rect 5325 22714 5427 22726
rect 5879 22714 5981 22726
rect 6433 22714 6535 22726
rect 6987 22714 7089 22726
rect 7539 22714 7645 22726
rect 4569 22649 4647 22683
rect 4681 22649 4692 22683
rect 4569 22546 4692 22649
rect 4569 22512 4647 22546
rect 4681 22512 4692 22546
rect 4569 22409 4692 22512
rect 4569 22375 4647 22409
rect 4681 22375 4692 22409
rect 4569 22272 4692 22375
rect 4569 22238 4647 22272
rect 4681 22238 4692 22272
rect 4569 22135 4692 22238
rect 4569 22101 4647 22135
rect 4681 22101 4692 22135
rect 4569 21998 4692 22101
rect 4569 21964 4647 21998
rect 4681 21964 4692 21998
rect 4569 21861 4692 21964
rect 4569 21827 4647 21861
rect 4681 21827 4692 21861
rect 4569 21724 4692 21827
rect 4569 21690 4647 21724
rect 4681 21690 4692 21724
rect 4569 21587 4692 21690
rect 4569 21553 4647 21587
rect 4681 21553 4692 21587
rect 4569 21450 4692 21553
rect 4569 21416 4647 21450
rect 4681 21416 4692 21450
rect 4569 21313 4692 21416
rect 5080 22680 5118 22714
rect 5046 22641 5152 22680
rect 5080 22607 5118 22641
rect 5046 22568 5152 22607
rect 5080 22534 5118 22568
rect 5046 22495 5152 22534
rect 5080 22461 5118 22495
rect 5046 22422 5152 22461
rect 5357 22680 5395 22714
rect 5323 22641 5429 22680
rect 5357 22607 5395 22641
rect 5323 22568 5429 22607
rect 5357 22534 5395 22568
rect 5323 22495 5429 22534
rect 5357 22461 5395 22495
rect 5323 22422 5429 22461
rect 5634 22680 5672 22714
rect 5600 22641 5706 22680
rect 5634 22607 5672 22641
rect 5600 22568 5706 22607
rect 5634 22534 5672 22568
rect 5600 22495 5706 22534
rect 5634 22461 5672 22495
rect 5600 22422 5706 22461
rect 5911 22680 5949 22714
rect 5877 22641 5983 22680
rect 5911 22607 5949 22641
rect 5877 22568 5983 22607
rect 5911 22534 5949 22568
rect 5877 22495 5983 22534
rect 5911 22461 5949 22495
rect 5877 22422 5983 22461
rect 6188 22680 6226 22714
rect 6154 22641 6260 22680
rect 6188 22607 6226 22641
rect 6154 22568 6260 22607
rect 6188 22534 6226 22568
rect 6154 22495 6260 22534
rect 6188 22461 6226 22495
rect 6154 22422 6260 22461
rect 6465 22680 6503 22714
rect 6431 22641 6537 22680
rect 6465 22607 6503 22641
rect 6431 22568 6537 22607
rect 6465 22534 6503 22568
rect 6431 22495 6537 22534
rect 6465 22461 6503 22495
rect 6431 22422 6537 22461
rect 6742 22680 6780 22714
rect 6708 22641 6814 22680
rect 6742 22607 6780 22641
rect 6708 22568 6814 22607
rect 6742 22534 6780 22568
rect 6708 22495 6814 22534
rect 6742 22461 6780 22495
rect 6708 22422 6814 22461
rect 7019 22680 7057 22714
rect 6985 22641 7091 22680
rect 7019 22607 7057 22641
rect 6985 22568 7091 22607
rect 7019 22534 7057 22568
rect 6985 22495 7091 22534
rect 7019 22461 7057 22495
rect 6985 22422 7091 22461
rect 7296 22680 7334 22714
rect 7262 22641 7368 22680
rect 7296 22607 7334 22641
rect 7262 22568 7368 22607
rect 7296 22534 7334 22568
rect 7262 22495 7368 22534
rect 7296 22461 7334 22495
rect 7262 22422 7368 22461
rect 7573 22680 7611 22714
rect 7539 22641 7645 22680
rect 7573 22607 7611 22641
rect 7539 22568 7645 22607
rect 7573 22534 7611 22568
rect 7539 22495 7645 22534
rect 7573 22461 7611 22495
rect 7539 22422 7645 22461
rect 7850 22680 7888 22714
rect 7816 22641 7922 22680
rect 7850 22607 7888 22641
rect 7816 22568 7922 22607
rect 7850 22534 7888 22568
rect 7816 22495 7922 22534
rect 7850 22461 7888 22495
rect 7816 22422 7922 22461
rect 5325 21368 5427 21380
rect 5879 21368 5981 21380
rect 6433 21368 6535 21380
rect 6987 21368 7089 21380
rect 7539 21368 7645 21380
rect 4569 21279 4647 21313
rect 4681 21279 4692 21313
rect 4569 21176 4692 21279
rect 4569 21142 4647 21176
rect 4681 21142 4692 21176
rect 4569 21039 4692 21142
rect 5239 21049 5251 21083
rect 5289 21049 5325 21083
rect 5360 21049 5395 21083
rect 5435 21049 5465 21083
rect 5510 21049 5535 21083
rect 5585 21049 5605 21083
rect 5660 21049 5675 21083
rect 5735 21049 5745 21083
rect 5810 21049 5815 21083
rect 5849 21049 5851 21083
rect 5919 21049 5926 21083
rect 5988 21049 6001 21083
rect 6057 21049 6076 21083
rect 6126 21049 6151 21083
rect 6195 21049 6225 21083
rect 6264 21049 6299 21083
rect 6333 21049 6368 21083
rect 6407 21049 6437 21083
rect 6481 21049 6506 21083
rect 6555 21049 6575 21083
rect 6629 21049 6644 21083
rect 6703 21049 6713 21083
rect 6777 21049 6782 21083
rect 6816 21049 6817 21083
rect 6885 21049 6891 21083
rect 6954 21049 6989 21083
rect 7023 21049 7058 21083
rect 7092 21049 7127 21083
rect 7161 21049 7196 21083
rect 7230 21049 7265 21083
rect 7299 21049 7334 21083
rect 7368 21049 7403 21083
rect 7437 21049 7472 21083
rect 7506 21049 7541 21083
rect 7575 21049 7610 21083
rect 7644 21049 7679 21083
rect 7713 21049 7729 21083
rect 4569 21005 4647 21039
rect 4681 21005 4692 21039
rect 4569 20902 4692 21005
rect 4569 20868 4647 20902
rect 4681 20868 4692 20902
rect 4569 20765 4692 20868
rect 4569 20731 4647 20765
rect 4681 20731 4692 20765
rect 4569 20628 4692 20731
rect 5325 20714 5427 20726
rect 5879 20714 5981 20726
rect 6433 20714 6535 20726
rect 6987 20714 7089 20726
rect 7539 20714 7645 20726
rect 4569 20594 4647 20628
rect 4681 20594 4692 20628
rect 4569 20491 4692 20594
rect 4569 20457 4647 20491
rect 4681 20457 4692 20491
rect 4569 20354 4692 20457
rect 4569 20320 4647 20354
rect 4681 20320 4692 20354
rect 4569 20217 4692 20320
rect 4569 20183 4647 20217
rect 4681 20183 4692 20217
rect 4569 20080 4692 20183
rect 4569 20046 4647 20080
rect 4681 20046 4692 20080
rect 4569 19943 4692 20046
rect 4569 19909 4647 19943
rect 4681 19909 4692 19943
rect 4569 19806 4692 19909
rect 4569 19772 4647 19806
rect 4681 19772 4692 19806
rect 4569 19669 4692 19772
rect 4569 19635 4647 19669
rect 4681 19635 4692 19669
rect 4569 19532 4692 19635
rect 4569 19498 4647 19532
rect 4681 19498 4692 19532
rect 4569 19395 4692 19498
rect 4569 19361 4647 19395
rect 4681 19361 4692 19395
rect 5080 20680 5118 20714
rect 5046 20641 5152 20680
rect 5080 20607 5118 20641
rect 5046 20568 5152 20607
rect 5080 20534 5118 20568
rect 5046 20495 5152 20534
rect 5080 20461 5118 20495
rect 5046 20422 5152 20461
rect 5357 20680 5395 20714
rect 5323 20641 5429 20680
rect 5357 20607 5395 20641
rect 5323 20568 5429 20607
rect 5357 20534 5395 20568
rect 5323 20495 5429 20534
rect 5357 20461 5395 20495
rect 5323 20422 5429 20461
rect 5634 20680 5672 20714
rect 5600 20641 5706 20680
rect 5634 20607 5672 20641
rect 5600 20568 5706 20607
rect 5634 20534 5672 20568
rect 5600 20495 5706 20534
rect 5634 20461 5672 20495
rect 5600 20422 5706 20461
rect 5911 20680 5949 20714
rect 5877 20641 5983 20680
rect 5911 20607 5949 20641
rect 5877 20568 5983 20607
rect 5911 20534 5949 20568
rect 5877 20495 5983 20534
rect 5911 20461 5949 20495
rect 5877 20422 5983 20461
rect 6188 20680 6226 20714
rect 6154 20641 6260 20680
rect 6188 20607 6226 20641
rect 6154 20568 6260 20607
rect 6188 20534 6226 20568
rect 6154 20495 6260 20534
rect 6188 20461 6226 20495
rect 6154 20422 6260 20461
rect 6465 20680 6503 20714
rect 6431 20641 6537 20680
rect 6465 20607 6503 20641
rect 6431 20568 6537 20607
rect 6465 20534 6503 20568
rect 6431 20495 6537 20534
rect 6465 20461 6503 20495
rect 6431 20422 6537 20461
rect 6742 20680 6780 20714
rect 6708 20641 6814 20680
rect 6742 20607 6780 20641
rect 6708 20568 6814 20607
rect 6742 20534 6780 20568
rect 6708 20495 6814 20534
rect 6742 20461 6780 20495
rect 6708 20422 6814 20461
rect 7019 20680 7057 20714
rect 6985 20641 7091 20680
rect 7019 20607 7057 20641
rect 6985 20568 7091 20607
rect 7019 20534 7057 20568
rect 6985 20495 7091 20534
rect 7019 20461 7057 20495
rect 6985 20422 7091 20461
rect 7296 20680 7334 20714
rect 7262 20641 7368 20680
rect 7296 20607 7334 20641
rect 7262 20568 7368 20607
rect 7296 20534 7334 20568
rect 7262 20495 7368 20534
rect 7296 20461 7334 20495
rect 7262 20422 7368 20461
rect 7573 20680 7611 20714
rect 7539 20641 7645 20680
rect 7573 20607 7611 20641
rect 7539 20568 7645 20607
rect 7573 20534 7611 20568
rect 7539 20495 7645 20534
rect 7573 20461 7611 20495
rect 7539 20422 7645 20461
rect 7850 20680 7888 20714
rect 7816 20641 7922 20680
rect 7850 20607 7888 20641
rect 7816 20568 7922 20607
rect 7850 20534 7888 20568
rect 7816 20495 7922 20534
rect 7850 20461 7888 20495
rect 7816 20422 7922 20461
rect 5325 19368 5427 19380
rect 5879 19368 5981 19380
rect 6433 19368 6535 19380
rect 6987 19368 7089 19380
rect 7539 19368 7645 19380
rect 4569 19258 4692 19361
rect 4569 19224 4647 19258
rect 4681 19224 4692 19258
rect 4569 19121 4692 19224
rect 4569 19087 4647 19121
rect 4681 19087 4692 19121
rect 4569 18984 4692 19087
rect 5239 19085 5251 19119
rect 5289 19085 5325 19119
rect 5359 19085 5395 19119
rect 5433 19085 5465 19119
rect 5507 19085 5535 19119
rect 5581 19085 5605 19119
rect 5655 19085 5675 19119
rect 5729 19085 5745 19119
rect 5803 19085 5815 19119
rect 5877 19085 5885 19119
rect 5951 19085 5954 19119
rect 5988 19085 5991 19119
rect 6057 19085 6065 19119
rect 6126 19085 6139 19119
rect 6195 19085 6213 19119
rect 6264 19085 6287 19119
rect 6333 19085 6361 19119
rect 6402 19085 6435 19119
rect 6471 19085 6506 19119
rect 6543 19085 6575 19119
rect 6617 19085 6644 19119
rect 6691 19085 6713 19119
rect 6765 19085 6782 19119
rect 6839 19085 6851 19119
rect 6913 19085 6920 19119
rect 6987 19085 6989 19119
rect 7023 19085 7026 19119
rect 7092 19085 7099 19119
rect 7161 19085 7172 19119
rect 7230 19085 7245 19119
rect 7299 19085 7318 19119
rect 7368 19085 7391 19119
rect 7437 19085 7464 19119
rect 7506 19085 7537 19119
rect 7575 19085 7610 19119
rect 7644 19085 7679 19119
rect 7717 19085 7729 19119
rect 4569 18950 4647 18984
rect 4681 18950 4692 18984
rect 4569 18847 4692 18950
rect 4569 18813 4647 18847
rect 4681 18813 4692 18847
rect 4569 18710 4692 18813
rect 5325 18714 5427 18726
rect 5879 18714 5981 18726
rect 6433 18714 6535 18726
rect 6987 18714 7089 18726
rect 7539 18714 7645 18726
rect 4569 18676 4647 18710
rect 4681 18676 4692 18710
rect 4569 18573 4692 18676
rect 4569 18563 4647 18573
rect 2648 18539 2715 18563
rect 2749 18539 2853 18563
rect 2887 18539 2991 18563
rect 3025 18539 3129 18563
rect 3163 18539 3267 18563
rect 3301 18539 3405 18563
rect 3439 18539 3543 18563
rect 3577 18539 3681 18563
rect 3715 18539 3819 18563
rect 3853 18539 3957 18563
rect 3991 18539 4095 18563
rect 4129 18539 4233 18563
rect 4267 18539 4371 18563
rect 4405 18539 4509 18563
rect 4543 18539 4647 18563
rect 4681 18539 4692 18573
rect 2648 18524 4692 18539
rect 2648 18490 2663 18524
rect 2697 18490 2735 18524
rect 2769 18490 2807 18524
rect 2841 18490 2879 18524
rect 2913 18490 2951 18524
rect 2985 18490 3023 18524
rect 3057 18490 3095 18524
rect 3129 18490 3167 18524
rect 3201 18490 3239 18524
rect 3273 18490 3311 18524
rect 3345 18490 3383 18524
rect 3417 18490 3455 18524
rect 3489 18490 3527 18524
rect 3561 18490 3599 18524
rect 3633 18490 3671 18524
rect 3705 18490 3743 18524
rect 3777 18490 3815 18524
rect 3849 18490 3887 18524
rect 3921 18490 3959 18524
rect 3993 18490 4031 18524
rect 4065 18490 4103 18524
rect 4137 18490 4175 18524
rect 4209 18490 4247 18524
rect 4281 18490 4319 18524
rect 4353 18490 4391 18524
rect 4425 18490 4463 18524
rect 4497 18490 4535 18524
rect 4569 18490 4692 18524
rect 2648 18451 4692 18490
rect 2648 18417 2663 18451
rect 2697 18436 2735 18451
rect 2697 18417 2715 18436
rect 2769 18417 2807 18451
rect 2841 18436 2879 18451
rect 2841 18417 2853 18436
rect 2913 18417 2951 18451
rect 2985 18436 3023 18451
rect 2985 18417 2991 18436
rect 3057 18417 3095 18451
rect 3129 18436 3167 18451
rect 2648 18402 2715 18417
rect 2749 18402 2853 18417
rect 2887 18402 2991 18417
rect 3025 18402 3129 18417
rect 3163 18417 3167 18436
rect 3201 18417 3239 18451
rect 3273 18436 3311 18451
rect 3301 18417 3311 18436
rect 3345 18417 3383 18451
rect 3417 18436 3455 18451
rect 3439 18417 3455 18436
rect 3489 18417 3527 18451
rect 3561 18436 3599 18451
rect 3577 18417 3599 18436
rect 3633 18417 3671 18451
rect 3705 18436 3743 18451
rect 3715 18417 3743 18436
rect 3777 18417 3815 18451
rect 3849 18436 3887 18451
rect 3853 18417 3887 18436
rect 3921 18436 3959 18451
rect 3921 18417 3957 18436
rect 3993 18417 4031 18451
rect 4065 18436 4103 18451
rect 4065 18417 4095 18436
rect 4137 18417 4175 18451
rect 4209 18436 4247 18451
rect 4209 18417 4233 18436
rect 4281 18417 4319 18451
rect 4353 18436 4391 18451
rect 4353 18417 4371 18436
rect 4425 18417 4463 18451
rect 4497 18436 4535 18451
rect 4569 18436 4692 18451
rect 4497 18417 4509 18436
rect 4569 18417 4647 18436
rect 3163 18402 3267 18417
rect 3301 18402 3405 18417
rect 3439 18402 3543 18417
rect 3577 18402 3681 18417
rect 3715 18402 3819 18417
rect 3853 18402 3957 18417
rect 3991 18402 4095 18417
rect 4129 18402 4233 18417
rect 4267 18402 4371 18417
rect 4405 18402 4509 18417
rect 4543 18402 4647 18417
rect 4681 18402 4692 18436
rect 2648 18378 4692 18402
rect 2648 18344 2663 18378
rect 2697 18344 2735 18378
rect 2769 18344 2807 18378
rect 2841 18344 2879 18378
rect 2913 18344 2951 18378
rect 2985 18344 3023 18378
rect 3057 18344 3095 18378
rect 3129 18344 3167 18378
rect 3201 18344 3239 18378
rect 3273 18344 3311 18378
rect 3345 18344 3383 18378
rect 3417 18344 3455 18378
rect 3489 18344 3527 18378
rect 3561 18344 3599 18378
rect 3633 18344 3671 18378
rect 3705 18344 3743 18378
rect 3777 18344 3815 18378
rect 3849 18344 3887 18378
rect 3921 18344 3959 18378
rect 3993 18344 4031 18378
rect 4065 18344 4103 18378
rect 4137 18344 4175 18378
rect 4209 18344 4247 18378
rect 4281 18344 4319 18378
rect 4353 18344 4391 18378
rect 4425 18344 4463 18378
rect 4497 18344 4535 18378
rect 4569 18344 4692 18378
rect 2648 18305 4692 18344
rect 2648 18271 2663 18305
rect 2697 18299 2735 18305
rect 2697 18271 2715 18299
rect 2769 18271 2807 18305
rect 2841 18299 2879 18305
rect 2841 18271 2853 18299
rect 2913 18271 2951 18305
rect 2985 18299 3023 18305
rect 2985 18271 2991 18299
rect 3057 18271 3095 18305
rect 3129 18299 3167 18305
rect 2648 18265 2715 18271
rect 2749 18265 2853 18271
rect 2887 18265 2991 18271
rect 3025 18265 3129 18271
rect 3163 18271 3167 18299
rect 3201 18271 3239 18305
rect 3273 18299 3311 18305
rect 3301 18271 3311 18299
rect 3345 18271 3383 18305
rect 3417 18299 3455 18305
rect 3439 18271 3455 18299
rect 3489 18271 3527 18305
rect 3561 18299 3599 18305
rect 3577 18271 3599 18299
rect 3633 18271 3671 18305
rect 3705 18299 3743 18305
rect 3715 18271 3743 18299
rect 3777 18271 3815 18305
rect 3849 18299 3887 18305
rect 3853 18271 3887 18299
rect 3921 18299 3959 18305
rect 3921 18271 3957 18299
rect 3993 18271 4031 18305
rect 4065 18299 4103 18305
rect 4065 18271 4095 18299
rect 4137 18271 4175 18305
rect 4209 18299 4247 18305
rect 4209 18271 4233 18299
rect 4281 18271 4319 18305
rect 4353 18299 4391 18305
rect 4353 18271 4371 18299
rect 4425 18271 4463 18305
rect 4497 18299 4535 18305
rect 4569 18299 4692 18305
rect 4497 18271 4509 18299
rect 4569 18271 4647 18299
rect 3163 18265 3267 18271
rect 3301 18265 3405 18271
rect 3439 18265 3543 18271
rect 3577 18265 3681 18271
rect 3715 18265 3819 18271
rect 3853 18265 3957 18271
rect 3991 18265 4095 18271
rect 4129 18265 4233 18271
rect 4267 18265 4371 18271
rect 4405 18265 4509 18271
rect 4543 18265 4647 18271
rect 4681 18265 4692 18299
rect 2648 18232 4692 18265
rect 2648 18198 2663 18232
rect 2697 18198 2735 18232
rect 2769 18198 2807 18232
rect 2841 18198 2879 18232
rect 2913 18198 2951 18232
rect 2985 18198 3023 18232
rect 3057 18198 3095 18232
rect 3129 18198 3167 18232
rect 3201 18198 3239 18232
rect 3273 18198 3311 18232
rect 3345 18198 3383 18232
rect 3417 18198 3455 18232
rect 3489 18198 3527 18232
rect 3561 18198 3599 18232
rect 3633 18198 3671 18232
rect 3705 18198 3743 18232
rect 3777 18198 3815 18232
rect 3849 18198 3887 18232
rect 3921 18198 3959 18232
rect 3993 18198 4031 18232
rect 4065 18198 4103 18232
rect 4137 18198 4175 18232
rect 4209 18198 4247 18232
rect 4281 18198 4319 18232
rect 4353 18198 4391 18232
rect 4425 18198 4463 18232
rect 4497 18198 4535 18232
rect 4569 18198 4692 18232
rect 2648 18162 4692 18198
rect 2648 18159 2715 18162
rect 2749 18159 2853 18162
rect 2887 18159 2991 18162
rect 3025 18159 3129 18162
rect 2648 18125 2663 18159
rect 2697 18128 2715 18159
rect 2697 18125 2735 18128
rect 2769 18125 2807 18159
rect 2841 18128 2853 18159
rect 2841 18125 2879 18128
rect 2913 18125 2951 18159
rect 2985 18128 2991 18159
rect 2985 18125 3023 18128
rect 3057 18125 3095 18159
rect 3163 18159 3267 18162
rect 3301 18159 3405 18162
rect 3439 18159 3543 18162
rect 3577 18159 3681 18162
rect 3715 18159 3819 18162
rect 3853 18159 3957 18162
rect 3991 18159 4095 18162
rect 4129 18159 4233 18162
rect 4267 18159 4371 18162
rect 4405 18159 4509 18162
rect 4543 18159 4647 18162
rect 3163 18128 3167 18159
rect 3129 18125 3167 18128
rect 3201 18125 3239 18159
rect 3301 18128 3311 18159
rect 3273 18125 3311 18128
rect 3345 18125 3383 18159
rect 3439 18128 3455 18159
rect 3417 18125 3455 18128
rect 3489 18125 3527 18159
rect 3577 18128 3599 18159
rect 3561 18125 3599 18128
rect 3633 18125 3671 18159
rect 3715 18128 3743 18159
rect 3705 18125 3743 18128
rect 3777 18125 3815 18159
rect 3853 18128 3887 18159
rect 3849 18125 3887 18128
rect 3921 18128 3957 18159
rect 3921 18125 3959 18128
rect 3993 18125 4031 18159
rect 4065 18128 4095 18159
rect 4065 18125 4103 18128
rect 4137 18125 4175 18159
rect 4209 18128 4233 18159
rect 4209 18125 4247 18128
rect 4281 18125 4319 18159
rect 4353 18128 4371 18159
rect 4353 18125 4391 18128
rect 4425 18125 4463 18159
rect 4497 18128 4509 18159
rect 4569 18128 4647 18159
rect 4681 18128 4692 18162
rect 4497 18125 4535 18128
rect 4569 18125 4692 18128
rect 2648 18086 4692 18125
rect 2648 18052 2663 18086
rect 2697 18052 2735 18086
rect 2769 18052 2807 18086
rect 2841 18052 2879 18086
rect 2913 18052 2951 18086
rect 2985 18052 3023 18086
rect 3057 18052 3095 18086
rect 3129 18052 3167 18086
rect 3201 18052 3239 18086
rect 3273 18052 3311 18086
rect 3345 18052 3383 18086
rect 3417 18052 3455 18086
rect 3489 18052 3527 18086
rect 3561 18052 3599 18086
rect 3633 18052 3671 18086
rect 3705 18052 3743 18086
rect 3777 18052 3815 18086
rect 3849 18052 3887 18086
rect 3921 18052 3959 18086
rect 3993 18052 4031 18086
rect 4065 18052 4103 18086
rect 4137 18052 4175 18086
rect 4209 18052 4247 18086
rect 4281 18052 4319 18086
rect 4353 18052 4391 18086
rect 4425 18052 4463 18086
rect 4497 18052 4535 18086
rect 4569 18052 4692 18086
rect 2648 18025 4692 18052
rect 2648 18013 2715 18025
rect 2749 18013 2853 18025
rect 2887 18013 2991 18025
rect 3025 18013 3129 18025
rect 2648 17979 2663 18013
rect 2697 17991 2715 18013
rect 2697 17979 2735 17991
rect 2769 17979 2807 18013
rect 2841 17991 2853 18013
rect 2841 17979 2879 17991
rect 2913 17979 2951 18013
rect 2985 17991 2991 18013
rect 2985 17979 3023 17991
rect 3057 17979 3095 18013
rect 3163 18013 3267 18025
rect 3301 18013 3405 18025
rect 3439 18013 3543 18025
rect 3577 18013 3681 18025
rect 3715 18013 3819 18025
rect 3853 18013 3957 18025
rect 3991 18013 4095 18025
rect 4129 18013 4233 18025
rect 4267 18013 4371 18025
rect 4405 18013 4509 18025
rect 4543 18013 4647 18025
rect 3163 17991 3167 18013
rect 3129 17979 3167 17991
rect 3201 17979 3239 18013
rect 3301 17991 3311 18013
rect 3273 17979 3311 17991
rect 3345 17979 3383 18013
rect 3439 17991 3455 18013
rect 3417 17979 3455 17991
rect 3489 17979 3527 18013
rect 3577 17991 3599 18013
rect 3561 17979 3599 17991
rect 3633 17979 3671 18013
rect 3715 17991 3743 18013
rect 3705 17979 3743 17991
rect 3777 17979 3815 18013
rect 3853 17991 3887 18013
rect 3849 17979 3887 17991
rect 3921 17991 3957 18013
rect 3921 17979 3959 17991
rect 3993 17979 4031 18013
rect 4065 17991 4095 18013
rect 4065 17979 4103 17991
rect 4137 17979 4175 18013
rect 4209 17991 4233 18013
rect 4209 17979 4247 17991
rect 4281 17979 4319 18013
rect 4353 17991 4371 18013
rect 4353 17979 4391 17991
rect 4425 17979 4463 18013
rect 4497 17991 4509 18013
rect 4569 17991 4647 18013
rect 4681 17991 4692 18025
rect 4497 17979 4535 17991
rect 4569 17979 4692 17991
rect 2648 17940 4692 17979
rect 2648 17906 2663 17940
rect 2697 17906 2735 17940
rect 2769 17906 2807 17940
rect 2841 17906 2879 17940
rect 2913 17906 2951 17940
rect 2985 17906 3023 17940
rect 3057 17906 3095 17940
rect 3129 17906 3167 17940
rect 3201 17906 3239 17940
rect 3273 17906 3311 17940
rect 3345 17906 3383 17940
rect 3417 17906 3455 17940
rect 3489 17906 3527 17940
rect 3561 17906 3599 17940
rect 3633 17906 3671 17940
rect 3705 17906 3743 17940
rect 3777 17906 3815 17940
rect 3849 17906 3887 17940
rect 3921 17906 3959 17940
rect 3993 17906 4031 17940
rect 4065 17906 4103 17940
rect 4137 17906 4175 17940
rect 4209 17906 4247 17940
rect 4281 17906 4319 17940
rect 4353 17906 4391 17940
rect 4425 17906 4463 17940
rect 4497 17906 4535 17940
rect 4569 17906 4692 17940
rect 2648 17888 4692 17906
rect 2648 17867 2715 17888
rect 2749 17867 2853 17888
rect 2887 17867 2991 17888
rect 3025 17867 3129 17888
rect 2648 17833 2663 17867
rect 2697 17854 2715 17867
rect 2697 17833 2735 17854
rect 2769 17833 2807 17867
rect 2841 17854 2853 17867
rect 2841 17833 2879 17854
rect 2913 17833 2951 17867
rect 2985 17854 2991 17867
rect 2985 17833 3023 17854
rect 3057 17833 3095 17867
rect 3163 17867 3267 17888
rect 3301 17867 3405 17888
rect 3439 17867 3543 17888
rect 3577 17867 3681 17888
rect 3715 17867 3819 17888
rect 3853 17867 3957 17888
rect 3991 17867 4095 17888
rect 4129 17867 4233 17888
rect 4267 17867 4371 17888
rect 4405 17867 4509 17888
rect 4543 17867 4647 17888
rect 3163 17854 3167 17867
rect 3129 17833 3167 17854
rect 3201 17833 3239 17867
rect 3301 17854 3311 17867
rect 3273 17833 3311 17854
rect 3345 17833 3383 17867
rect 3439 17854 3455 17867
rect 3417 17833 3455 17854
rect 3489 17833 3527 17867
rect 3577 17854 3599 17867
rect 3561 17833 3599 17854
rect 3633 17833 3671 17867
rect 3715 17854 3743 17867
rect 3705 17833 3743 17854
rect 3777 17833 3815 17867
rect 3853 17854 3887 17867
rect 3849 17833 3887 17854
rect 3921 17854 3957 17867
rect 3921 17833 3959 17854
rect 3993 17833 4031 17867
rect 4065 17854 4095 17867
rect 4065 17833 4103 17854
rect 4137 17833 4175 17867
rect 4209 17854 4233 17867
rect 4209 17833 4247 17854
rect 4281 17833 4319 17867
rect 4353 17854 4371 17867
rect 4353 17833 4391 17854
rect 4425 17833 4463 17867
rect 4497 17854 4509 17867
rect 4569 17854 4647 17867
rect 4681 17854 4692 17888
rect 4497 17833 4535 17854
rect 4569 17833 4692 17854
rect 2648 17794 4692 17833
rect 2648 17760 2663 17794
rect 2697 17760 2735 17794
rect 2769 17760 2807 17794
rect 2841 17760 2879 17794
rect 2913 17760 2951 17794
rect 2985 17760 3023 17794
rect 3057 17760 3095 17794
rect 3129 17760 3167 17794
rect 3201 17760 3239 17794
rect 3273 17760 3311 17794
rect 3345 17760 3383 17794
rect 3417 17760 3455 17794
rect 3489 17760 3527 17794
rect 3561 17760 3599 17794
rect 3633 17760 3671 17794
rect 3705 17760 3743 17794
rect 3777 17760 3815 17794
rect 3849 17760 3887 17794
rect 3921 17760 3959 17794
rect 3993 17760 4031 17794
rect 4065 17760 4103 17794
rect 4137 17760 4175 17794
rect 4209 17760 4247 17794
rect 4281 17760 4319 17794
rect 4353 17760 4391 17794
rect 4425 17760 4463 17794
rect 4497 17760 4535 17794
rect 4569 17760 4692 17794
rect 2648 17751 4692 17760
rect 2648 17721 2715 17751
rect 2749 17721 2853 17751
rect 2887 17721 2991 17751
rect 3025 17721 3129 17751
rect 2648 17687 2663 17721
rect 2697 17717 2715 17721
rect 2697 17687 2735 17717
rect 2769 17687 2807 17721
rect 2841 17717 2853 17721
rect 2841 17687 2879 17717
rect 2913 17687 2951 17721
rect 2985 17717 2991 17721
rect 2985 17687 3023 17717
rect 3057 17687 3095 17721
rect 3163 17721 3267 17751
rect 3301 17721 3405 17751
rect 3439 17721 3543 17751
rect 3577 17721 3681 17751
rect 3715 17721 3819 17751
rect 3853 17721 3957 17751
rect 3991 17721 4095 17751
rect 4129 17721 4233 17751
rect 4267 17721 4371 17751
rect 4405 17721 4509 17751
rect 4543 17721 4647 17751
rect 3163 17717 3167 17721
rect 3129 17687 3167 17717
rect 3201 17687 3239 17721
rect 3301 17717 3311 17721
rect 3273 17687 3311 17717
rect 3345 17687 3383 17721
rect 3439 17717 3455 17721
rect 3417 17687 3455 17717
rect 3489 17687 3527 17721
rect 3577 17717 3599 17721
rect 3561 17687 3599 17717
rect 3633 17687 3671 17721
rect 3715 17717 3743 17721
rect 3705 17687 3743 17717
rect 3777 17687 3815 17721
rect 3853 17717 3887 17721
rect 3849 17687 3887 17717
rect 3921 17717 3957 17721
rect 3921 17687 3959 17717
rect 3993 17687 4031 17721
rect 4065 17717 4095 17721
rect 4065 17687 4103 17717
rect 4137 17687 4175 17721
rect 4209 17717 4233 17721
rect 4209 17687 4247 17717
rect 4281 17687 4319 17721
rect 4353 17717 4371 17721
rect 4353 17687 4391 17717
rect 4425 17687 4463 17721
rect 4497 17717 4509 17721
rect 4569 17717 4647 17721
rect 4681 17717 4692 17751
rect 4497 17687 4535 17717
rect 4569 17687 4692 17717
rect 2648 17648 4692 17687
rect 2648 17614 2663 17648
rect 2697 17614 2735 17648
rect 2769 17614 2807 17648
rect 2841 17614 2879 17648
rect 2913 17614 2951 17648
rect 2985 17614 3023 17648
rect 3057 17614 3095 17648
rect 3129 17614 3167 17648
rect 3201 17614 3239 17648
rect 3273 17614 3311 17648
rect 3345 17614 3383 17648
rect 3417 17614 3455 17648
rect 3489 17614 3527 17648
rect 3561 17614 3599 17648
rect 3633 17614 3671 17648
rect 3705 17614 3743 17648
rect 3777 17614 3815 17648
rect 3849 17614 3887 17648
rect 3921 17614 3959 17648
rect 3993 17614 4031 17648
rect 4065 17614 4103 17648
rect 4137 17614 4175 17648
rect 4209 17614 4247 17648
rect 4281 17614 4319 17648
rect 4353 17614 4391 17648
rect 4425 17614 4463 17648
rect 4497 17614 4535 17648
rect 4569 17614 4692 17648
rect 2648 17580 2715 17614
rect 2749 17580 2853 17614
rect 2887 17580 2991 17614
rect 3025 17580 3129 17614
rect 3163 17580 3267 17614
rect 3301 17580 3405 17614
rect 3439 17580 3543 17614
rect 3577 17580 3681 17614
rect 3715 17580 3819 17614
rect 3853 17580 3957 17614
rect 3991 17580 4095 17614
rect 4129 17580 4233 17614
rect 4267 17580 4371 17614
rect 4405 17580 4509 17614
rect 4543 17580 4647 17614
rect 4681 17580 4692 17614
rect 2648 17575 4692 17580
rect 2648 17541 2663 17575
rect 2697 17541 2735 17575
rect 2769 17541 2807 17575
rect 2841 17541 2879 17575
rect 2913 17541 2951 17575
rect 2985 17541 3023 17575
rect 3057 17541 3095 17575
rect 3129 17541 3167 17575
rect 3201 17541 3239 17575
rect 3273 17541 3311 17575
rect 3345 17541 3383 17575
rect 3417 17541 3455 17575
rect 3489 17541 3527 17575
rect 3561 17541 3599 17575
rect 3633 17541 3671 17575
rect 3705 17541 3743 17575
rect 3777 17541 3815 17575
rect 3849 17541 3887 17575
rect 3921 17541 3959 17575
rect 3993 17541 4031 17575
rect 4065 17541 4103 17575
rect 4137 17541 4175 17575
rect 4209 17541 4247 17575
rect 4281 17541 4319 17575
rect 4353 17541 4391 17575
rect 4425 17541 4463 17575
rect 4497 17541 4535 17575
rect 4569 17541 4692 17575
rect 2648 17502 4692 17541
rect 2648 17468 2663 17502
rect 2697 17477 2735 17502
rect 2697 17468 2715 17477
rect 2769 17468 2807 17502
rect 2841 17477 2879 17502
rect 2841 17468 2853 17477
rect 2913 17468 2951 17502
rect 2985 17477 3023 17502
rect 2985 17468 2991 17477
rect 3057 17468 3095 17502
rect 3129 17477 3167 17502
rect 2648 17443 2715 17468
rect 2749 17443 2853 17468
rect 2887 17443 2991 17468
rect 3025 17443 3129 17468
rect 3163 17468 3167 17477
rect 3201 17468 3239 17502
rect 3273 17477 3311 17502
rect 3301 17468 3311 17477
rect 3345 17468 3383 17502
rect 3417 17477 3455 17502
rect 3439 17468 3455 17477
rect 3489 17468 3527 17502
rect 3561 17477 3599 17502
rect 3577 17468 3599 17477
rect 3633 17468 3671 17502
rect 3705 17477 3743 17502
rect 3715 17468 3743 17477
rect 3777 17468 3815 17502
rect 3849 17477 3887 17502
rect 3853 17468 3887 17477
rect 3921 17477 3959 17502
rect 3921 17468 3957 17477
rect 3993 17468 4031 17502
rect 4065 17477 4103 17502
rect 4065 17468 4095 17477
rect 4137 17468 4175 17502
rect 4209 17477 4247 17502
rect 4209 17468 4233 17477
rect 4281 17468 4319 17502
rect 4353 17477 4391 17502
rect 4353 17468 4371 17477
rect 4425 17468 4463 17502
rect 4497 17477 4535 17502
rect 4569 17477 4692 17502
rect 4497 17468 4509 17477
rect 4569 17468 4647 17477
rect 3163 17443 3267 17468
rect 3301 17443 3405 17468
rect 3439 17443 3543 17468
rect 3577 17443 3681 17468
rect 3715 17443 3819 17468
rect 3853 17443 3957 17468
rect 3991 17443 4095 17468
rect 4129 17443 4233 17468
rect 4267 17443 4371 17468
rect 4405 17443 4509 17468
rect 4543 17443 4647 17468
rect 4681 17443 4692 17477
rect 2648 17429 4692 17443
rect 2648 17395 2663 17429
rect 2697 17395 2735 17429
rect 2769 17395 2807 17429
rect 2841 17395 2879 17429
rect 2913 17395 2951 17429
rect 2985 17395 3023 17429
rect 3057 17395 3095 17429
rect 3129 17395 3167 17429
rect 3201 17395 3239 17429
rect 3273 17395 3311 17429
rect 3345 17395 3383 17429
rect 3417 17395 3455 17429
rect 3489 17395 3527 17429
rect 3561 17395 3599 17429
rect 3633 17395 3671 17429
rect 3705 17395 3743 17429
rect 3777 17395 3815 17429
rect 3849 17395 3887 17429
rect 3921 17395 3959 17429
rect 3993 17395 4031 17429
rect 4065 17395 4103 17429
rect 4137 17395 4175 17429
rect 4209 17395 4247 17429
rect 4281 17395 4319 17429
rect 4353 17395 4391 17429
rect 4425 17395 4463 17429
rect 4497 17395 4535 17429
rect 4569 17395 4692 17429
rect 2648 17356 4692 17395
rect 5080 18680 5118 18714
rect 5046 18641 5152 18680
rect 5080 18607 5118 18641
rect 5046 18568 5152 18607
rect 5080 18534 5118 18568
rect 5046 18495 5152 18534
rect 5080 18461 5118 18495
rect 5046 18422 5152 18461
rect 5357 18680 5395 18714
rect 5323 18641 5429 18680
rect 5357 18607 5395 18641
rect 5323 18568 5429 18607
rect 5357 18534 5395 18568
rect 5323 18495 5429 18534
rect 5357 18461 5395 18495
rect 5323 18422 5429 18461
rect 5634 18680 5672 18714
rect 5600 18641 5706 18680
rect 5634 18607 5672 18641
rect 5600 18568 5706 18607
rect 5634 18534 5672 18568
rect 5600 18495 5706 18534
rect 5634 18461 5672 18495
rect 5600 18422 5706 18461
rect 5911 18680 5949 18714
rect 5877 18641 5983 18680
rect 5911 18607 5949 18641
rect 5877 18568 5983 18607
rect 5911 18534 5949 18568
rect 5877 18495 5983 18534
rect 5911 18461 5949 18495
rect 5877 18422 5983 18461
rect 6188 18680 6226 18714
rect 6154 18641 6260 18680
rect 6188 18607 6226 18641
rect 6154 18568 6260 18607
rect 6188 18534 6226 18568
rect 6154 18495 6260 18534
rect 6188 18461 6226 18495
rect 6154 18422 6260 18461
rect 6465 18680 6503 18714
rect 6431 18641 6537 18680
rect 6465 18607 6503 18641
rect 6431 18568 6537 18607
rect 6465 18534 6503 18568
rect 6431 18495 6537 18534
rect 6465 18461 6503 18495
rect 6431 18422 6537 18461
rect 6742 18680 6780 18714
rect 6708 18641 6814 18680
rect 6742 18607 6780 18641
rect 6708 18568 6814 18607
rect 6742 18534 6780 18568
rect 6708 18495 6814 18534
rect 6742 18461 6780 18495
rect 6708 18422 6814 18461
rect 7019 18680 7057 18714
rect 6985 18641 7091 18680
rect 7019 18607 7057 18641
rect 6985 18568 7091 18607
rect 7019 18534 7057 18568
rect 6985 18495 7091 18534
rect 7019 18461 7057 18495
rect 6985 18422 7091 18461
rect 7296 18680 7334 18714
rect 7262 18641 7368 18680
rect 7296 18607 7334 18641
rect 7262 18568 7368 18607
rect 7296 18534 7334 18568
rect 7262 18495 7368 18534
rect 7296 18461 7334 18495
rect 7262 18422 7368 18461
rect 7573 18680 7611 18714
rect 7539 18641 7645 18680
rect 7573 18607 7611 18641
rect 7539 18568 7645 18607
rect 7573 18534 7611 18568
rect 7539 18495 7645 18534
rect 7573 18461 7611 18495
rect 7539 18422 7645 18461
rect 7850 18680 7888 18714
rect 7816 18641 7922 18680
rect 7850 18607 7888 18641
rect 7816 18568 7922 18607
rect 7850 18534 7888 18568
rect 7816 18495 7922 18534
rect 7850 18461 7888 18495
rect 7816 18422 7922 18461
rect 5325 17368 5427 17380
rect 5879 17368 5981 17380
rect 6433 17368 6535 17380
rect 6987 17368 7089 17380
rect 7539 17368 7645 17380
rect 2648 17322 2663 17356
rect 2697 17340 2735 17356
rect 2697 17322 2715 17340
rect 2769 17322 2807 17356
rect 2841 17340 2879 17356
rect 2841 17322 2853 17340
rect 2913 17322 2951 17356
rect 2985 17340 3023 17356
rect 2985 17322 2991 17340
rect 3057 17322 3095 17356
rect 3129 17340 3167 17356
rect 2648 17306 2715 17322
rect 2749 17306 2853 17322
rect 2887 17306 2991 17322
rect 3025 17306 3129 17322
rect 3163 17322 3167 17340
rect 3201 17322 3239 17356
rect 3273 17340 3311 17356
rect 3301 17322 3311 17340
rect 3345 17322 3383 17356
rect 3417 17340 3455 17356
rect 3439 17322 3455 17340
rect 3489 17322 3527 17356
rect 3561 17340 3599 17356
rect 3577 17322 3599 17340
rect 3633 17322 3671 17356
rect 3705 17340 3743 17356
rect 3715 17322 3743 17340
rect 3777 17322 3815 17356
rect 3849 17340 3887 17356
rect 3853 17322 3887 17340
rect 3921 17340 3959 17356
rect 3921 17322 3957 17340
rect 3993 17322 4031 17356
rect 4065 17340 4103 17356
rect 4065 17322 4095 17340
rect 4137 17322 4175 17356
rect 4209 17340 4247 17356
rect 4209 17322 4233 17340
rect 4281 17322 4319 17356
rect 4353 17340 4391 17356
rect 4353 17322 4371 17340
rect 4425 17322 4463 17356
rect 4497 17340 4535 17356
rect 4569 17340 4692 17356
rect 4497 17322 4509 17340
rect 4569 17322 4647 17340
rect 3163 17306 3267 17322
rect 3301 17306 3405 17322
rect 3439 17306 3543 17322
rect 3577 17306 3681 17322
rect 3715 17306 3819 17322
rect 3853 17306 3957 17322
rect 3991 17306 4095 17322
rect 4129 17306 4233 17322
rect 4267 17306 4371 17322
rect 4405 17306 4509 17322
rect 4543 17306 4647 17322
rect 4681 17306 4692 17340
rect 2648 17283 4692 17306
rect 2648 17249 2663 17283
rect 2697 17249 2735 17283
rect 2769 17249 2807 17283
rect 2841 17249 2879 17283
rect 2913 17249 2951 17283
rect 2985 17249 3023 17283
rect 3057 17249 3095 17283
rect 3129 17249 3167 17283
rect 3201 17249 3239 17283
rect 3273 17249 3311 17283
rect 3345 17249 3383 17283
rect 3417 17249 3455 17283
rect 3489 17249 3527 17283
rect 3561 17249 3599 17283
rect 3633 17249 3671 17283
rect 3705 17249 3743 17283
rect 3777 17249 3815 17283
rect 3849 17249 3887 17283
rect 3921 17249 3959 17283
rect 3993 17249 4031 17283
rect 4065 17249 4103 17283
rect 4137 17249 4175 17283
rect 4209 17249 4247 17283
rect 4281 17249 4319 17283
rect 4353 17249 4391 17283
rect 4425 17249 4463 17283
rect 4497 17249 4535 17283
rect 4569 17249 4692 17283
rect 2648 17210 4692 17249
rect 5239 17211 5251 17245
rect 5289 17211 5325 17245
rect 5359 17211 5395 17245
rect 5433 17211 5465 17245
rect 5507 17211 5535 17245
rect 5581 17211 5605 17245
rect 5655 17211 5675 17245
rect 5729 17211 5745 17245
rect 5803 17211 5815 17245
rect 5877 17211 5885 17245
rect 5951 17211 5954 17245
rect 5988 17211 5991 17245
rect 6057 17211 6065 17245
rect 6126 17211 6139 17245
rect 6195 17211 6213 17245
rect 6264 17211 6287 17245
rect 6333 17211 6361 17245
rect 6402 17211 6435 17245
rect 6471 17211 6506 17245
rect 6543 17211 6575 17245
rect 6617 17211 6644 17245
rect 6691 17211 6713 17245
rect 6765 17211 6782 17245
rect 6839 17211 6851 17245
rect 6913 17211 6920 17245
rect 6987 17211 6989 17245
rect 7023 17211 7026 17245
rect 7092 17211 7099 17245
rect 7161 17211 7172 17245
rect 7230 17211 7245 17245
rect 7299 17211 7318 17245
rect 7368 17211 7391 17245
rect 7437 17211 7464 17245
rect 7506 17211 7537 17245
rect 7575 17211 7610 17245
rect 7644 17211 7679 17245
rect 7717 17211 7729 17245
rect 2648 17176 2663 17210
rect 2697 17203 2735 17210
rect 2697 17176 2715 17203
rect 2769 17176 2807 17210
rect 2841 17203 2879 17210
rect 2841 17176 2853 17203
rect 2913 17176 2951 17210
rect 2985 17203 3023 17210
rect 2985 17176 2991 17203
rect 3057 17176 3095 17210
rect 3129 17203 3167 17210
rect 2648 17169 2715 17176
rect 2749 17169 2853 17176
rect 2887 17169 2991 17176
rect 3025 17169 3129 17176
rect 3163 17176 3167 17203
rect 3201 17176 3239 17210
rect 3273 17203 3311 17210
rect 3301 17176 3311 17203
rect 3345 17176 3383 17210
rect 3417 17203 3455 17210
rect 3439 17176 3455 17203
rect 3489 17176 3527 17210
rect 3561 17203 3599 17210
rect 3577 17176 3599 17203
rect 3633 17176 3671 17210
rect 3705 17203 3743 17210
rect 3715 17176 3743 17203
rect 3777 17176 3815 17210
rect 3849 17203 3887 17210
rect 3853 17176 3887 17203
rect 3921 17203 3959 17210
rect 3921 17176 3957 17203
rect 3993 17176 4031 17210
rect 4065 17203 4103 17210
rect 4065 17176 4095 17203
rect 4137 17176 4175 17210
rect 4209 17203 4247 17210
rect 4209 17176 4233 17203
rect 4281 17176 4319 17210
rect 4353 17203 4391 17210
rect 4353 17176 4371 17203
rect 4425 17176 4463 17210
rect 4497 17203 4535 17210
rect 4569 17203 4692 17210
rect 4497 17176 4509 17203
rect 4569 17176 4647 17203
rect 3163 17169 3267 17176
rect 3301 17169 3405 17176
rect 3439 17169 3543 17176
rect 3577 17169 3681 17176
rect 3715 17169 3819 17176
rect 3853 17169 3957 17176
rect 3991 17169 4095 17176
rect 4129 17169 4233 17176
rect 4267 17169 4371 17176
rect 4405 17169 4509 17176
rect 4543 17169 4647 17176
rect 4681 17169 4692 17203
rect 2648 17137 4692 17169
rect 2648 17103 2663 17137
rect 2697 17103 2735 17137
rect 2769 17103 2807 17137
rect 2841 17103 2879 17137
rect 2913 17103 2951 17137
rect 2985 17103 3023 17137
rect 3057 17103 3095 17137
rect 3129 17103 3167 17137
rect 3201 17103 3239 17137
rect 3273 17103 3311 17137
rect 3345 17103 3383 17137
rect 3417 17103 3455 17137
rect 3489 17103 3527 17137
rect 3561 17103 3599 17137
rect 3633 17103 3671 17137
rect 3705 17103 3743 17137
rect 3777 17103 3815 17137
rect 3849 17103 3887 17137
rect 3921 17103 3959 17137
rect 3993 17103 4031 17137
rect 4065 17103 4103 17137
rect 4137 17103 4175 17137
rect 4209 17103 4247 17137
rect 4281 17103 4319 17137
rect 4353 17103 4391 17137
rect 4425 17103 4463 17137
rect 4497 17103 4535 17137
rect 4569 17103 4692 17137
rect 2648 17072 4692 17103
rect 2648 17066 7908 17072
rect 2648 17064 2715 17066
rect 2749 17064 2853 17066
rect 2887 17064 2991 17066
rect 3025 17064 3129 17066
rect 2648 17030 2663 17064
rect 2697 17032 2715 17064
rect 2697 17030 2735 17032
rect 2769 17030 2807 17064
rect 2841 17032 2853 17064
rect 2841 17030 2879 17032
rect 2913 17030 2951 17064
rect 2985 17032 2991 17064
rect 2985 17030 3023 17032
rect 3057 17030 3095 17064
rect 3163 17064 3267 17066
rect 3301 17064 3405 17066
rect 3439 17064 3543 17066
rect 3577 17064 3681 17066
rect 3715 17064 3819 17066
rect 3853 17064 3957 17066
rect 3991 17064 4095 17066
rect 4129 17064 4233 17066
rect 4267 17064 4371 17066
rect 4405 17064 4509 17066
rect 4543 17064 4647 17066
rect 3163 17032 3167 17064
rect 3129 17030 3167 17032
rect 3201 17030 3239 17064
rect 3301 17032 3311 17064
rect 3273 17030 3311 17032
rect 3345 17030 3383 17064
rect 3439 17032 3455 17064
rect 3417 17030 3455 17032
rect 3489 17030 3527 17064
rect 3577 17032 3599 17064
rect 3561 17030 3599 17032
rect 3633 17030 3671 17064
rect 3715 17032 3743 17064
rect 3705 17030 3743 17032
rect 3777 17030 3815 17064
rect 3853 17032 3887 17064
rect 3849 17030 3887 17032
rect 3921 17032 3957 17064
rect 3921 17030 3959 17032
rect 3993 17030 4031 17064
rect 4065 17032 4095 17064
rect 4065 17030 4103 17032
rect 4137 17030 4175 17064
rect 4209 17032 4233 17064
rect 4209 17030 4247 17032
rect 4281 17030 4319 17064
rect 4353 17032 4371 17064
rect 4353 17030 4391 17032
rect 4425 17030 4463 17064
rect 4497 17032 4509 17064
rect 4569 17032 4647 17064
rect 4681 17034 7908 17066
rect 4681 17032 4740 17034
rect 4497 17030 4535 17032
rect 4569 17030 4740 17032
rect 2648 17000 4740 17030
rect 4774 17000 4809 17034
rect 4843 17000 4878 17034
rect 4912 17000 4947 17034
rect 4981 17000 5016 17034
rect 5050 17000 5085 17034
rect 5119 17000 5154 17034
rect 5188 17000 5223 17034
rect 5257 17000 5292 17034
rect 5326 17000 5361 17034
rect 5395 17000 5430 17034
rect 5464 17000 5499 17034
rect 5533 17000 5568 17034
rect 5602 17000 5637 17034
rect 5671 17000 5706 17034
rect 5740 17000 5775 17034
rect 5809 17000 5844 17034
rect 5878 17000 5913 17034
rect 5947 17000 5982 17034
rect 6016 17000 6051 17034
rect 6085 17000 6120 17034
rect 6154 17000 6189 17034
rect 6223 17000 6258 17034
rect 6292 17000 6327 17034
rect 6361 17000 6396 17034
rect 6430 17000 6465 17034
rect 6499 17000 6534 17034
rect 6568 17000 6603 17034
rect 6637 17000 6672 17034
rect 6706 17000 6741 17034
rect 6775 17000 6810 17034
rect 6844 17000 6879 17034
rect 6913 17000 6948 17034
rect 6982 17000 7017 17034
rect 7051 17000 7086 17034
rect 7120 17000 7155 17034
rect 7189 17000 7224 17034
rect 7258 17000 7293 17034
rect 7327 17000 7362 17034
rect 7396 17000 7431 17034
rect 7465 17000 7500 17034
rect 7534 17000 7568 17034
rect 7602 17000 7636 17034
rect 7670 17000 7704 17034
rect 7738 17000 7772 17034
rect 7806 17000 7840 17034
rect 7874 17000 7908 17034
rect 2648 16991 7908 17000
rect 2648 16957 2663 16991
rect 2697 16957 2735 16991
rect 2769 16957 2807 16991
rect 2841 16957 2879 16991
rect 2913 16957 2951 16991
rect 2985 16957 3023 16991
rect 3057 16957 3095 16991
rect 3129 16957 3167 16991
rect 3201 16957 3239 16991
rect 3273 16957 3311 16991
rect 3345 16957 3383 16991
rect 3417 16957 3455 16991
rect 3489 16957 3527 16991
rect 3561 16957 3599 16991
rect 3633 16957 3671 16991
rect 3705 16957 3743 16991
rect 3777 16957 3815 16991
rect 3849 16957 3887 16991
rect 3921 16957 3959 16991
rect 3993 16957 4031 16991
rect 4065 16957 4103 16991
rect 4137 16957 4175 16991
rect 4209 16957 4247 16991
rect 4281 16957 4319 16991
rect 4353 16957 4391 16991
rect 4425 16957 4463 16991
rect 4497 16957 4535 16991
rect 4569 16989 7908 16991
rect 4569 16964 5089 16989
rect 5123 16964 5162 16989
rect 5196 16964 5235 16989
rect 5269 16964 5308 16989
rect 5342 16964 5381 16989
rect 5415 16964 5454 16989
rect 5488 16964 5527 16989
rect 5561 16964 5600 16989
rect 5634 16964 5673 16989
rect 5707 16964 5746 16989
rect 5780 16964 5819 16989
rect 5853 16964 5892 16989
rect 5926 16964 5965 16989
rect 5999 16964 6038 16989
rect 6072 16964 6110 16989
rect 6144 16964 6182 16989
rect 6216 16964 6254 16989
rect 6288 16964 6326 16989
rect 6360 16964 6398 16989
rect 6432 16964 6470 16989
rect 6504 16964 6542 16989
rect 6576 16964 6614 16989
rect 6648 16964 6686 16989
rect 6720 16964 6758 16989
rect 6792 16964 6830 16989
rect 6864 16964 6902 16989
rect 6936 16964 6974 16989
rect 7008 16964 7046 16989
rect 7080 16964 7118 16989
rect 7152 16964 7190 16989
rect 4569 16957 4740 16964
rect 2648 16930 4740 16957
rect 4774 16930 4809 16964
rect 4843 16930 4878 16964
rect 4912 16930 4947 16964
rect 4981 16930 5016 16964
rect 5050 16930 5085 16964
rect 5123 16955 5154 16964
rect 5196 16955 5223 16964
rect 5269 16955 5292 16964
rect 5342 16955 5361 16964
rect 5415 16955 5430 16964
rect 5488 16955 5499 16964
rect 5561 16955 5568 16964
rect 5634 16955 5637 16964
rect 5119 16930 5154 16955
rect 5188 16930 5223 16955
rect 5257 16930 5292 16955
rect 5326 16930 5361 16955
rect 5395 16930 5430 16955
rect 5464 16930 5499 16955
rect 5533 16930 5568 16955
rect 5602 16930 5637 16955
rect 5671 16955 5673 16964
rect 5740 16955 5746 16964
rect 5809 16955 5819 16964
rect 5878 16955 5892 16964
rect 5947 16955 5965 16964
rect 6016 16955 6038 16964
rect 6085 16955 6110 16964
rect 6154 16955 6182 16964
rect 6223 16955 6254 16964
rect 6292 16955 6326 16964
rect 5671 16930 5706 16955
rect 5740 16930 5775 16955
rect 5809 16930 5844 16955
rect 5878 16930 5913 16955
rect 5947 16930 5982 16955
rect 6016 16930 6051 16955
rect 6085 16930 6120 16955
rect 6154 16930 6189 16955
rect 6223 16930 6258 16955
rect 6292 16930 6327 16955
rect 6361 16930 6396 16964
rect 6432 16955 6465 16964
rect 6504 16955 6534 16964
rect 6576 16955 6603 16964
rect 6648 16955 6672 16964
rect 6720 16955 6741 16964
rect 6792 16955 6810 16964
rect 6864 16955 6879 16964
rect 6936 16955 6948 16964
rect 7008 16955 7017 16964
rect 7080 16955 7086 16964
rect 7152 16955 7155 16964
rect 6430 16930 6465 16955
rect 6499 16930 6534 16955
rect 6568 16930 6603 16955
rect 6637 16930 6672 16955
rect 6706 16930 6741 16955
rect 6775 16930 6810 16955
rect 6844 16930 6879 16955
rect 6913 16930 6948 16955
rect 6982 16930 7017 16955
rect 7051 16930 7086 16955
rect 7120 16930 7155 16955
rect 7189 16955 7190 16964
rect 7224 16964 7262 16989
rect 7296 16964 7334 16989
rect 7368 16964 7406 16989
rect 7440 16964 7478 16989
rect 7512 16964 7550 16989
rect 7584 16964 7622 16989
rect 7656 16964 7694 16989
rect 7728 16964 7766 16989
rect 7800 16964 7838 16989
rect 7872 16964 7908 16989
rect 7189 16930 7224 16955
rect 7258 16955 7262 16964
rect 7327 16955 7334 16964
rect 7396 16955 7406 16964
rect 7465 16955 7478 16964
rect 7534 16955 7550 16964
rect 7602 16955 7622 16964
rect 7670 16955 7694 16964
rect 7738 16955 7766 16964
rect 7806 16955 7838 16964
rect 7258 16930 7293 16955
rect 7327 16930 7362 16955
rect 7396 16930 7431 16955
rect 7465 16930 7500 16955
rect 7534 16930 7568 16955
rect 7602 16930 7636 16955
rect 7670 16930 7704 16955
rect 7738 16930 7772 16955
rect 7806 16930 7840 16955
rect 7874 16930 7908 16964
rect 2648 16929 7908 16930
rect 2648 16918 2715 16929
rect 2749 16918 2853 16929
rect 2887 16918 2991 16929
rect 3025 16918 3129 16929
rect 2648 16884 2663 16918
rect 2697 16895 2715 16918
rect 2697 16884 2735 16895
rect 2769 16884 2807 16918
rect 2841 16895 2853 16918
rect 2841 16884 2879 16895
rect 2913 16884 2951 16918
rect 2985 16895 2991 16918
rect 2985 16884 3023 16895
rect 3057 16884 3095 16918
rect 3163 16918 3267 16929
rect 3301 16918 3405 16929
rect 3439 16918 3543 16929
rect 3577 16918 3681 16929
rect 3715 16918 3819 16929
rect 3853 16918 3957 16929
rect 3991 16918 4095 16929
rect 4129 16918 4233 16929
rect 4267 16918 4371 16929
rect 4405 16918 4509 16929
rect 4543 16918 4647 16929
rect 3163 16895 3167 16918
rect 3129 16884 3167 16895
rect 3201 16884 3239 16918
rect 3301 16895 3311 16918
rect 3273 16884 3311 16895
rect 3345 16884 3383 16918
rect 3439 16895 3455 16918
rect 3417 16884 3455 16895
rect 3489 16884 3527 16918
rect 3577 16895 3599 16918
rect 3561 16884 3599 16895
rect 3633 16884 3671 16918
rect 3715 16895 3743 16918
rect 3705 16884 3743 16895
rect 3777 16884 3815 16918
rect 3853 16895 3887 16918
rect 3849 16884 3887 16895
rect 3921 16895 3957 16918
rect 3921 16884 3959 16895
rect 3993 16884 4031 16918
rect 4065 16895 4095 16918
rect 4065 16884 4103 16895
rect 4137 16884 4175 16918
rect 4209 16895 4233 16918
rect 4209 16884 4247 16895
rect 4281 16884 4319 16918
rect 4353 16895 4371 16918
rect 4353 16884 4391 16895
rect 4425 16884 4463 16918
rect 4497 16895 4509 16918
rect 4569 16895 4647 16918
rect 4681 16913 7908 16929
rect 4681 16895 5089 16913
rect 4497 16884 4535 16895
rect 4569 16894 5089 16895
rect 5123 16894 5162 16913
rect 5196 16894 5235 16913
rect 5269 16894 5308 16913
rect 5342 16894 5381 16913
rect 5415 16894 5454 16913
rect 5488 16894 5527 16913
rect 5561 16894 5600 16913
rect 5634 16894 5673 16913
rect 5707 16894 5746 16913
rect 5780 16894 5819 16913
rect 5853 16894 5892 16913
rect 5926 16894 5965 16913
rect 5999 16894 6038 16913
rect 6072 16894 6110 16913
rect 6144 16894 6182 16913
rect 6216 16894 6254 16913
rect 6288 16894 6326 16913
rect 6360 16894 6398 16913
rect 6432 16894 6470 16913
rect 6504 16894 6542 16913
rect 6576 16894 6614 16913
rect 6648 16894 6686 16913
rect 6720 16894 6758 16913
rect 6792 16894 6830 16913
rect 6864 16894 6902 16913
rect 6936 16894 6974 16913
rect 7008 16894 7046 16913
rect 7080 16894 7118 16913
rect 7152 16894 7190 16913
rect 4569 16884 4740 16894
rect 2648 16860 4740 16884
rect 4774 16860 4809 16894
rect 4843 16860 4878 16894
rect 4912 16860 4947 16894
rect 4981 16860 5016 16894
rect 5050 16860 5085 16894
rect 5123 16879 5154 16894
rect 5196 16879 5223 16894
rect 5269 16879 5292 16894
rect 5342 16879 5361 16894
rect 5415 16879 5430 16894
rect 5488 16879 5499 16894
rect 5561 16879 5568 16894
rect 5634 16879 5637 16894
rect 5119 16860 5154 16879
rect 5188 16860 5223 16879
rect 5257 16860 5292 16879
rect 5326 16860 5361 16879
rect 5395 16860 5430 16879
rect 5464 16860 5499 16879
rect 5533 16860 5568 16879
rect 5602 16860 5637 16879
rect 5671 16879 5673 16894
rect 5740 16879 5746 16894
rect 5809 16879 5819 16894
rect 5878 16879 5892 16894
rect 5947 16879 5965 16894
rect 6016 16879 6038 16894
rect 6085 16879 6110 16894
rect 6154 16879 6182 16894
rect 6223 16879 6254 16894
rect 6292 16879 6326 16894
rect 5671 16860 5706 16879
rect 5740 16860 5775 16879
rect 5809 16860 5844 16879
rect 5878 16860 5913 16879
rect 5947 16860 5982 16879
rect 6016 16860 6051 16879
rect 6085 16860 6120 16879
rect 6154 16860 6189 16879
rect 6223 16860 6258 16879
rect 6292 16860 6327 16879
rect 6361 16860 6396 16894
rect 6432 16879 6465 16894
rect 6504 16879 6534 16894
rect 6576 16879 6603 16894
rect 6648 16879 6672 16894
rect 6720 16879 6741 16894
rect 6792 16879 6810 16894
rect 6864 16879 6879 16894
rect 6936 16879 6948 16894
rect 7008 16879 7017 16894
rect 7080 16879 7086 16894
rect 7152 16879 7155 16894
rect 6430 16860 6465 16879
rect 6499 16860 6534 16879
rect 6568 16860 6603 16879
rect 6637 16860 6672 16879
rect 6706 16860 6741 16879
rect 6775 16860 6810 16879
rect 6844 16860 6879 16879
rect 6913 16860 6948 16879
rect 6982 16860 7017 16879
rect 7051 16860 7086 16879
rect 7120 16860 7155 16879
rect 7189 16879 7190 16894
rect 7224 16894 7262 16913
rect 7296 16894 7334 16913
rect 7368 16894 7406 16913
rect 7440 16894 7478 16913
rect 7512 16894 7550 16913
rect 7584 16894 7622 16913
rect 7656 16894 7694 16913
rect 7728 16894 7766 16913
rect 7800 16894 7838 16913
rect 7872 16894 7908 16913
rect 7189 16860 7224 16879
rect 7258 16879 7262 16894
rect 7327 16879 7334 16894
rect 7396 16879 7406 16894
rect 7465 16879 7478 16894
rect 7534 16879 7550 16894
rect 7602 16879 7622 16894
rect 7670 16879 7694 16894
rect 7738 16879 7766 16894
rect 7806 16879 7838 16894
rect 7258 16860 7293 16879
rect 7327 16860 7362 16879
rect 7396 16860 7431 16879
rect 7465 16860 7500 16879
rect 7534 16860 7568 16879
rect 7602 16860 7636 16879
rect 7670 16860 7704 16879
rect 7738 16860 7772 16879
rect 7806 16860 7840 16879
rect 7874 16860 7908 16894
rect 2648 16845 7908 16860
rect 2648 16811 2663 16845
rect 2697 16811 2735 16845
rect 2769 16811 2807 16845
rect 2841 16811 2879 16845
rect 2913 16811 2951 16845
rect 2985 16811 3023 16845
rect 3057 16811 3095 16845
rect 3129 16811 3167 16845
rect 3201 16811 3239 16845
rect 3273 16811 3311 16845
rect 3345 16811 3383 16845
rect 3417 16811 3455 16845
rect 3489 16811 3527 16845
rect 3561 16811 3599 16845
rect 3633 16811 3671 16845
rect 3705 16811 3743 16845
rect 3777 16811 3815 16845
rect 3849 16811 3887 16845
rect 3921 16811 3959 16845
rect 3993 16811 4031 16845
rect 4065 16811 4103 16845
rect 4137 16811 4175 16845
rect 4209 16811 4247 16845
rect 4281 16811 4319 16845
rect 4353 16811 4391 16845
rect 4425 16811 4463 16845
rect 4497 16811 4535 16845
rect 4569 16837 7908 16845
rect 4569 16824 5089 16837
rect 5123 16824 5162 16837
rect 5196 16824 5235 16837
rect 5269 16824 5308 16837
rect 5342 16824 5381 16837
rect 5415 16824 5454 16837
rect 5488 16824 5527 16837
rect 5561 16824 5600 16837
rect 5634 16824 5673 16837
rect 5707 16824 5746 16837
rect 5780 16824 5819 16837
rect 5853 16824 5892 16837
rect 5926 16824 5965 16837
rect 5999 16824 6038 16837
rect 6072 16824 6110 16837
rect 6144 16824 6182 16837
rect 6216 16824 6254 16837
rect 6288 16824 6326 16837
rect 6360 16824 6398 16837
rect 6432 16824 6470 16837
rect 6504 16824 6542 16837
rect 6576 16824 6614 16837
rect 6648 16824 6686 16837
rect 6720 16824 6758 16837
rect 6792 16824 6830 16837
rect 6864 16824 6902 16837
rect 6936 16824 6974 16837
rect 7008 16824 7046 16837
rect 7080 16824 7118 16837
rect 7152 16824 7190 16837
rect 4569 16811 4740 16824
rect 2648 16792 4740 16811
rect 2648 16772 2715 16792
rect 2749 16772 2853 16792
rect 2887 16772 2991 16792
rect 3025 16772 3129 16792
rect 2648 16738 2663 16772
rect 2697 16758 2715 16772
rect 2697 16738 2735 16758
rect 2769 16738 2807 16772
rect 2841 16758 2853 16772
rect 2841 16738 2879 16758
rect 2913 16738 2951 16772
rect 2985 16758 2991 16772
rect 2985 16738 3023 16758
rect 3057 16738 3095 16772
rect 3163 16772 3267 16792
rect 3301 16772 3405 16792
rect 3439 16772 3543 16792
rect 3577 16772 3681 16792
rect 3715 16772 3819 16792
rect 3853 16772 3957 16792
rect 3991 16772 4095 16792
rect 4129 16772 4233 16792
rect 4267 16772 4371 16792
rect 4405 16772 4509 16792
rect 4543 16772 4647 16792
rect 3163 16758 3167 16772
rect 3129 16738 3167 16758
rect 3201 16738 3239 16772
rect 3301 16758 3311 16772
rect 3273 16738 3311 16758
rect 3345 16738 3383 16772
rect 3439 16758 3455 16772
rect 3417 16738 3455 16758
rect 3489 16738 3527 16772
rect 3577 16758 3599 16772
rect 3561 16738 3599 16758
rect 3633 16738 3671 16772
rect 3715 16758 3743 16772
rect 3705 16738 3743 16758
rect 3777 16738 3815 16772
rect 3853 16758 3887 16772
rect 3849 16738 3887 16758
rect 3921 16758 3957 16772
rect 3921 16738 3959 16758
rect 3993 16738 4031 16772
rect 4065 16758 4095 16772
rect 4065 16738 4103 16758
rect 4137 16738 4175 16772
rect 4209 16758 4233 16772
rect 4209 16738 4247 16758
rect 4281 16738 4319 16772
rect 4353 16758 4371 16772
rect 4353 16738 4391 16758
rect 4425 16738 4463 16772
rect 4497 16758 4509 16772
rect 4569 16758 4647 16772
rect 4681 16790 4740 16792
rect 4774 16790 4809 16824
rect 4843 16790 4878 16824
rect 4912 16790 4947 16824
rect 4981 16790 5016 16824
rect 5050 16790 5085 16824
rect 5123 16803 5154 16824
rect 5196 16803 5223 16824
rect 5269 16803 5292 16824
rect 5342 16803 5361 16824
rect 5415 16803 5430 16824
rect 5488 16803 5499 16824
rect 5561 16803 5568 16824
rect 5634 16803 5637 16824
rect 5119 16790 5154 16803
rect 5188 16790 5223 16803
rect 5257 16790 5292 16803
rect 5326 16790 5361 16803
rect 5395 16790 5430 16803
rect 5464 16790 5499 16803
rect 5533 16790 5568 16803
rect 5602 16790 5637 16803
rect 5671 16803 5673 16824
rect 5740 16803 5746 16824
rect 5809 16803 5819 16824
rect 5878 16803 5892 16824
rect 5947 16803 5965 16824
rect 6016 16803 6038 16824
rect 6085 16803 6110 16824
rect 6154 16803 6182 16824
rect 6223 16803 6254 16824
rect 6292 16803 6326 16824
rect 5671 16790 5706 16803
rect 5740 16790 5775 16803
rect 5809 16790 5844 16803
rect 5878 16790 5913 16803
rect 5947 16790 5982 16803
rect 6016 16790 6051 16803
rect 6085 16790 6120 16803
rect 6154 16790 6189 16803
rect 6223 16790 6258 16803
rect 6292 16790 6327 16803
rect 6361 16790 6396 16824
rect 6432 16803 6465 16824
rect 6504 16803 6534 16824
rect 6576 16803 6603 16824
rect 6648 16803 6672 16824
rect 6720 16803 6741 16824
rect 6792 16803 6810 16824
rect 6864 16803 6879 16824
rect 6936 16803 6948 16824
rect 7008 16803 7017 16824
rect 7080 16803 7086 16824
rect 7152 16803 7155 16824
rect 6430 16790 6465 16803
rect 6499 16790 6534 16803
rect 6568 16790 6603 16803
rect 6637 16790 6672 16803
rect 6706 16790 6741 16803
rect 6775 16790 6810 16803
rect 6844 16790 6879 16803
rect 6913 16790 6948 16803
rect 6982 16790 7017 16803
rect 7051 16790 7086 16803
rect 7120 16790 7155 16803
rect 7189 16803 7190 16824
rect 7224 16824 7262 16837
rect 7296 16824 7334 16837
rect 7368 16824 7406 16837
rect 7440 16824 7478 16837
rect 7512 16824 7550 16837
rect 7584 16824 7622 16837
rect 7656 16824 7694 16837
rect 7728 16824 7766 16837
rect 7800 16824 7838 16837
rect 7872 16824 7908 16837
rect 7189 16790 7224 16803
rect 7258 16803 7262 16824
rect 7327 16803 7334 16824
rect 7396 16803 7406 16824
rect 7465 16803 7478 16824
rect 7534 16803 7550 16824
rect 7602 16803 7622 16824
rect 7670 16803 7694 16824
rect 7738 16803 7766 16824
rect 7806 16803 7838 16824
rect 7258 16790 7293 16803
rect 7327 16790 7362 16803
rect 7396 16790 7431 16803
rect 7465 16790 7500 16803
rect 7534 16790 7568 16803
rect 7602 16790 7636 16803
rect 7670 16790 7704 16803
rect 7738 16790 7772 16803
rect 7806 16790 7840 16803
rect 7874 16790 7908 16824
rect 4681 16761 7908 16790
rect 4681 16758 5089 16761
rect 4497 16738 4535 16758
rect 4569 16754 5089 16758
rect 5123 16754 5162 16761
rect 5196 16754 5235 16761
rect 5269 16754 5308 16761
rect 5342 16754 5381 16761
rect 5415 16754 5454 16761
rect 5488 16754 5527 16761
rect 5561 16754 5600 16761
rect 5634 16754 5673 16761
rect 5707 16754 5746 16761
rect 5780 16754 5819 16761
rect 5853 16754 5892 16761
rect 5926 16754 5965 16761
rect 5999 16754 6038 16761
rect 6072 16754 6110 16761
rect 6144 16754 6182 16761
rect 6216 16754 6254 16761
rect 6288 16754 6326 16761
rect 6360 16754 6398 16761
rect 6432 16754 6470 16761
rect 6504 16754 6542 16761
rect 6576 16754 6614 16761
rect 6648 16754 6686 16761
rect 6720 16754 6758 16761
rect 6792 16754 6830 16761
rect 6864 16754 6902 16761
rect 6936 16754 6974 16761
rect 7008 16754 7046 16761
rect 7080 16754 7118 16761
rect 7152 16754 7190 16761
rect 4569 16738 4740 16754
rect 2648 16720 4740 16738
rect 4774 16720 4809 16754
rect 4843 16720 4878 16754
rect 4912 16720 4947 16754
rect 4981 16720 5016 16754
rect 5050 16720 5085 16754
rect 5123 16727 5154 16754
rect 5196 16727 5223 16754
rect 5269 16727 5292 16754
rect 5342 16727 5361 16754
rect 5415 16727 5430 16754
rect 5488 16727 5499 16754
rect 5561 16727 5568 16754
rect 5634 16727 5637 16754
rect 5119 16720 5154 16727
rect 5188 16720 5223 16727
rect 5257 16720 5292 16727
rect 5326 16720 5361 16727
rect 5395 16720 5430 16727
rect 5464 16720 5499 16727
rect 5533 16720 5568 16727
rect 5602 16720 5637 16727
rect 5671 16727 5673 16754
rect 5740 16727 5746 16754
rect 5809 16727 5819 16754
rect 5878 16727 5892 16754
rect 5947 16727 5965 16754
rect 6016 16727 6038 16754
rect 6085 16727 6110 16754
rect 6154 16727 6182 16754
rect 6223 16727 6254 16754
rect 6292 16727 6326 16754
rect 5671 16720 5706 16727
rect 5740 16720 5775 16727
rect 5809 16720 5844 16727
rect 5878 16720 5913 16727
rect 5947 16720 5982 16727
rect 6016 16720 6051 16727
rect 6085 16720 6120 16727
rect 6154 16720 6189 16727
rect 6223 16720 6258 16727
rect 6292 16720 6327 16727
rect 6361 16720 6396 16754
rect 6432 16727 6465 16754
rect 6504 16727 6534 16754
rect 6576 16727 6603 16754
rect 6648 16727 6672 16754
rect 6720 16727 6741 16754
rect 6792 16727 6810 16754
rect 6864 16727 6879 16754
rect 6936 16727 6948 16754
rect 7008 16727 7017 16754
rect 7080 16727 7086 16754
rect 7152 16727 7155 16754
rect 6430 16720 6465 16727
rect 6499 16720 6534 16727
rect 6568 16720 6603 16727
rect 6637 16720 6672 16727
rect 6706 16720 6741 16727
rect 6775 16720 6810 16727
rect 6844 16720 6879 16727
rect 6913 16720 6948 16727
rect 6982 16720 7017 16727
rect 7051 16720 7086 16727
rect 7120 16720 7155 16727
rect 7189 16727 7190 16754
rect 7224 16754 7262 16761
rect 7296 16754 7334 16761
rect 7368 16754 7406 16761
rect 7440 16754 7478 16761
rect 7512 16754 7550 16761
rect 7584 16754 7622 16761
rect 7656 16754 7694 16761
rect 7728 16754 7766 16761
rect 7800 16754 7838 16761
rect 7872 16754 7908 16761
rect 7189 16720 7224 16727
rect 7258 16727 7262 16754
rect 7327 16727 7334 16754
rect 7396 16727 7406 16754
rect 7465 16727 7478 16754
rect 7534 16727 7550 16754
rect 7602 16727 7622 16754
rect 7670 16727 7694 16754
rect 7738 16727 7766 16754
rect 7806 16727 7838 16754
rect 7258 16720 7293 16727
rect 7327 16720 7362 16727
rect 7396 16720 7431 16727
rect 7465 16720 7500 16727
rect 7534 16720 7568 16727
rect 7602 16720 7636 16727
rect 7670 16720 7704 16727
rect 7738 16720 7772 16727
rect 7806 16720 7840 16727
rect 7874 16720 7908 16754
rect 2648 16699 7908 16720
rect 2648 16665 2663 16699
rect 2697 16665 2735 16699
rect 2769 16665 2807 16699
rect 2841 16665 2879 16699
rect 2913 16665 2951 16699
rect 2985 16665 3023 16699
rect 3057 16665 3095 16699
rect 3129 16665 3167 16699
rect 3201 16665 3239 16699
rect 3273 16665 3311 16699
rect 3345 16665 3383 16699
rect 3417 16665 3455 16699
rect 3489 16665 3527 16699
rect 3561 16665 3599 16699
rect 3633 16665 3671 16699
rect 3705 16665 3743 16699
rect 3777 16665 3815 16699
rect 3849 16665 3887 16699
rect 3921 16665 3959 16699
rect 3993 16665 4031 16699
rect 4065 16665 4103 16699
rect 4137 16665 4175 16699
rect 4209 16665 4247 16699
rect 4281 16665 4319 16699
rect 4353 16665 4391 16699
rect 4425 16665 4463 16699
rect 4497 16665 4535 16699
rect 4569 16685 7908 16699
rect 4569 16684 5089 16685
rect 5123 16684 5162 16685
rect 5196 16684 5235 16685
rect 5269 16684 5308 16685
rect 5342 16684 5381 16685
rect 5415 16684 5454 16685
rect 5488 16684 5527 16685
rect 5561 16684 5600 16685
rect 5634 16684 5673 16685
rect 5707 16684 5746 16685
rect 5780 16684 5819 16685
rect 5853 16684 5892 16685
rect 5926 16684 5965 16685
rect 5999 16684 6038 16685
rect 6072 16684 6110 16685
rect 6144 16684 6182 16685
rect 6216 16684 6254 16685
rect 6288 16684 6326 16685
rect 6360 16684 6398 16685
rect 6432 16684 6470 16685
rect 6504 16684 6542 16685
rect 6576 16684 6614 16685
rect 6648 16684 6686 16685
rect 6720 16684 6758 16685
rect 6792 16684 6830 16685
rect 6864 16684 6902 16685
rect 6936 16684 6974 16685
rect 7008 16684 7046 16685
rect 7080 16684 7118 16685
rect 7152 16684 7190 16685
rect 4569 16665 4740 16684
rect 2648 16655 4740 16665
rect 2648 16626 2715 16655
rect 2749 16626 2853 16655
rect 2887 16626 2991 16655
rect 3025 16626 3129 16655
rect 2648 16592 2663 16626
rect 2697 16621 2715 16626
rect 2697 16592 2735 16621
rect 2769 16592 2807 16626
rect 2841 16621 2853 16626
rect 2841 16592 2879 16621
rect 2913 16592 2951 16626
rect 2985 16621 2991 16626
rect 2985 16592 3023 16621
rect 3057 16592 3095 16626
rect 3163 16626 3267 16655
rect 3301 16626 3405 16655
rect 3439 16626 3543 16655
rect 3577 16626 3681 16655
rect 3715 16626 3819 16655
rect 3853 16626 3957 16655
rect 3991 16626 4095 16655
rect 4129 16626 4233 16655
rect 4267 16626 4371 16655
rect 4405 16626 4509 16655
rect 4543 16626 4647 16655
rect 3163 16621 3167 16626
rect 3129 16592 3167 16621
rect 3201 16592 3239 16626
rect 3301 16621 3311 16626
rect 3273 16592 3311 16621
rect 3345 16592 3383 16626
rect 3439 16621 3455 16626
rect 3417 16592 3455 16621
rect 3489 16592 3527 16626
rect 3577 16621 3599 16626
rect 3561 16592 3599 16621
rect 3633 16592 3671 16626
rect 3715 16621 3743 16626
rect 3705 16592 3743 16621
rect 3777 16592 3815 16626
rect 3853 16621 3887 16626
rect 3849 16592 3887 16621
rect 3921 16621 3957 16626
rect 3921 16592 3959 16621
rect 3993 16592 4031 16626
rect 4065 16621 4095 16626
rect 4065 16592 4103 16621
rect 4137 16592 4175 16626
rect 4209 16621 4233 16626
rect 4209 16592 4247 16621
rect 4281 16592 4319 16626
rect 4353 16621 4371 16626
rect 4353 16592 4391 16621
rect 4425 16592 4463 16626
rect 4497 16621 4509 16626
rect 4569 16621 4647 16626
rect 4681 16650 4740 16655
rect 4774 16650 4809 16684
rect 4843 16650 4878 16684
rect 4912 16650 4947 16684
rect 4981 16650 5016 16684
rect 5050 16650 5085 16684
rect 5123 16651 5154 16684
rect 5196 16651 5223 16684
rect 5269 16651 5292 16684
rect 5342 16651 5361 16684
rect 5415 16651 5430 16684
rect 5488 16651 5499 16684
rect 5561 16651 5568 16684
rect 5634 16651 5637 16684
rect 5119 16650 5154 16651
rect 5188 16650 5223 16651
rect 5257 16650 5292 16651
rect 5326 16650 5361 16651
rect 5395 16650 5430 16651
rect 5464 16650 5499 16651
rect 5533 16650 5568 16651
rect 5602 16650 5637 16651
rect 5671 16651 5673 16684
rect 5740 16651 5746 16684
rect 5809 16651 5819 16684
rect 5878 16651 5892 16684
rect 5947 16651 5965 16684
rect 6016 16651 6038 16684
rect 6085 16651 6110 16684
rect 6154 16651 6182 16684
rect 6223 16651 6254 16684
rect 6292 16651 6326 16684
rect 5671 16650 5706 16651
rect 5740 16650 5775 16651
rect 5809 16650 5844 16651
rect 5878 16650 5913 16651
rect 5947 16650 5982 16651
rect 6016 16650 6051 16651
rect 6085 16650 6120 16651
rect 6154 16650 6189 16651
rect 6223 16650 6258 16651
rect 6292 16650 6327 16651
rect 6361 16650 6396 16684
rect 6432 16651 6465 16684
rect 6504 16651 6534 16684
rect 6576 16651 6603 16684
rect 6648 16651 6672 16684
rect 6720 16651 6741 16684
rect 6792 16651 6810 16684
rect 6864 16651 6879 16684
rect 6936 16651 6948 16684
rect 7008 16651 7017 16684
rect 7080 16651 7086 16684
rect 7152 16651 7155 16684
rect 6430 16650 6465 16651
rect 6499 16650 6534 16651
rect 6568 16650 6603 16651
rect 6637 16650 6672 16651
rect 6706 16650 6741 16651
rect 6775 16650 6810 16651
rect 6844 16650 6879 16651
rect 6913 16650 6948 16651
rect 6982 16650 7017 16651
rect 7051 16650 7086 16651
rect 7120 16650 7155 16651
rect 7189 16651 7190 16684
rect 7224 16684 7262 16685
rect 7296 16684 7334 16685
rect 7368 16684 7406 16685
rect 7440 16684 7478 16685
rect 7512 16684 7550 16685
rect 7584 16684 7622 16685
rect 7656 16684 7694 16685
rect 7728 16684 7766 16685
rect 7800 16684 7838 16685
rect 7872 16684 7908 16685
rect 7189 16650 7224 16651
rect 7258 16651 7262 16684
rect 7327 16651 7334 16684
rect 7396 16651 7406 16684
rect 7465 16651 7478 16684
rect 7534 16651 7550 16684
rect 7602 16651 7622 16684
rect 7670 16651 7694 16684
rect 7738 16651 7766 16684
rect 7806 16651 7838 16684
rect 7258 16650 7293 16651
rect 7327 16650 7362 16651
rect 7396 16650 7431 16651
rect 7465 16650 7500 16651
rect 7534 16650 7568 16651
rect 7602 16650 7636 16651
rect 7670 16650 7704 16651
rect 7738 16650 7772 16651
rect 7806 16650 7840 16651
rect 7874 16650 7908 16684
rect 4681 16621 7908 16650
rect 4497 16592 4535 16621
rect 4569 16614 7908 16621
rect 4569 16592 4740 16614
rect 2648 16580 4740 16592
rect 4774 16580 4809 16614
rect 4843 16580 4878 16614
rect 4912 16580 4947 16614
rect 4981 16580 5016 16614
rect 5050 16580 5085 16614
rect 5119 16609 5154 16614
rect 5188 16609 5223 16614
rect 5257 16609 5292 16614
rect 5326 16609 5361 16614
rect 5395 16609 5430 16614
rect 5464 16609 5499 16614
rect 5533 16609 5568 16614
rect 5602 16609 5637 16614
rect 5123 16580 5154 16609
rect 5196 16580 5223 16609
rect 5269 16580 5292 16609
rect 5342 16580 5361 16609
rect 5415 16580 5430 16609
rect 5488 16580 5499 16609
rect 5561 16580 5568 16609
rect 5634 16580 5637 16609
rect 5671 16609 5706 16614
rect 5740 16609 5775 16614
rect 5809 16609 5844 16614
rect 5878 16609 5913 16614
rect 5947 16609 5982 16614
rect 6016 16609 6051 16614
rect 6085 16609 6120 16614
rect 6154 16609 6189 16614
rect 6223 16609 6258 16614
rect 6292 16609 6327 16614
rect 5671 16580 5673 16609
rect 5740 16580 5746 16609
rect 5809 16580 5819 16609
rect 5878 16580 5892 16609
rect 5947 16580 5965 16609
rect 6016 16580 6038 16609
rect 6085 16580 6110 16609
rect 6154 16580 6182 16609
rect 6223 16580 6254 16609
rect 6292 16580 6326 16609
rect 6361 16580 6396 16614
rect 6430 16609 6465 16614
rect 6499 16609 6534 16614
rect 6568 16609 6603 16614
rect 6637 16609 6672 16614
rect 6706 16609 6741 16614
rect 6775 16609 6810 16614
rect 6844 16609 6879 16614
rect 6913 16609 6948 16614
rect 6982 16609 7017 16614
rect 7051 16609 7086 16614
rect 7120 16609 7155 16614
rect 6432 16580 6465 16609
rect 6504 16580 6534 16609
rect 6576 16580 6603 16609
rect 6648 16580 6672 16609
rect 6720 16580 6741 16609
rect 6792 16580 6810 16609
rect 6864 16580 6879 16609
rect 6936 16580 6948 16609
rect 7008 16580 7017 16609
rect 7080 16580 7086 16609
rect 7152 16580 7155 16609
rect 7189 16609 7224 16614
rect 7189 16580 7190 16609
rect 2648 16575 5089 16580
rect 5123 16575 5162 16580
rect 5196 16575 5235 16580
rect 5269 16575 5308 16580
rect 5342 16575 5381 16580
rect 5415 16575 5454 16580
rect 5488 16575 5527 16580
rect 5561 16575 5600 16580
rect 5634 16575 5673 16580
rect 5707 16575 5746 16580
rect 5780 16575 5819 16580
rect 5853 16575 5892 16580
rect 5926 16575 5965 16580
rect 5999 16575 6038 16580
rect 6072 16575 6110 16580
rect 6144 16575 6182 16580
rect 6216 16575 6254 16580
rect 6288 16575 6326 16580
rect 6360 16575 6398 16580
rect 6432 16575 6470 16580
rect 6504 16575 6542 16580
rect 6576 16575 6614 16580
rect 6648 16575 6686 16580
rect 6720 16575 6758 16580
rect 6792 16575 6830 16580
rect 6864 16575 6902 16580
rect 6936 16575 6974 16580
rect 7008 16575 7046 16580
rect 7080 16575 7118 16580
rect 7152 16575 7190 16580
rect 7258 16609 7293 16614
rect 7327 16609 7362 16614
rect 7396 16609 7431 16614
rect 7465 16609 7500 16614
rect 7534 16609 7568 16614
rect 7602 16609 7636 16614
rect 7670 16609 7704 16614
rect 7738 16609 7772 16614
rect 7806 16609 7840 16614
rect 7258 16580 7262 16609
rect 7327 16580 7334 16609
rect 7396 16580 7406 16609
rect 7465 16580 7478 16609
rect 7534 16580 7550 16609
rect 7602 16580 7622 16609
rect 7670 16580 7694 16609
rect 7738 16580 7766 16609
rect 7806 16580 7838 16609
rect 7874 16580 7908 16614
rect 7224 16575 7262 16580
rect 7296 16575 7334 16580
rect 7368 16575 7406 16580
rect 7440 16575 7478 16580
rect 7512 16575 7550 16580
rect 7584 16575 7622 16580
rect 7656 16575 7694 16580
rect 7728 16575 7766 16580
rect 7800 16575 7838 16580
rect 7872 16575 7908 16580
rect 2648 16553 7908 16575
rect 2648 16519 2663 16553
rect 2697 16519 2735 16553
rect 2769 16519 2807 16553
rect 2841 16519 2879 16553
rect 2913 16519 2951 16553
rect 2985 16519 3023 16553
rect 3057 16519 3095 16553
rect 3129 16519 3167 16553
rect 3201 16519 3239 16553
rect 3273 16519 3311 16553
rect 3345 16519 3383 16553
rect 3417 16519 3455 16553
rect 3489 16519 3527 16553
rect 3561 16519 3599 16553
rect 3633 16519 3671 16553
rect 3705 16519 3743 16553
rect 3777 16519 3815 16553
rect 3849 16519 3887 16553
rect 3921 16519 3959 16553
rect 3993 16519 4031 16553
rect 4065 16519 4103 16553
rect 4137 16519 4175 16553
rect 4209 16519 4247 16553
rect 4281 16519 4319 16553
rect 4353 16519 4391 16553
rect 4425 16519 4463 16553
rect 4497 16519 4535 16553
rect 4569 16544 7908 16553
rect 4569 16519 4740 16544
rect 2648 16518 4740 16519
rect 2648 16484 2715 16518
rect 2749 16484 2853 16518
rect 2887 16484 2991 16518
rect 3025 16484 3129 16518
rect 3163 16484 3267 16518
rect 3301 16484 3405 16518
rect 3439 16484 3543 16518
rect 3577 16484 3681 16518
rect 3715 16484 3819 16518
rect 3853 16484 3957 16518
rect 3991 16484 4095 16518
rect 4129 16484 4233 16518
rect 4267 16484 4371 16518
rect 4405 16484 4509 16518
rect 4543 16484 4647 16518
rect 4681 16510 4740 16518
rect 4774 16510 4809 16544
rect 4843 16510 4878 16544
rect 4912 16510 4947 16544
rect 4981 16510 5016 16544
rect 5050 16510 5085 16544
rect 5119 16533 5154 16544
rect 5188 16533 5223 16544
rect 5257 16533 5292 16544
rect 5326 16533 5361 16544
rect 5395 16533 5430 16544
rect 5464 16533 5499 16544
rect 5533 16533 5568 16544
rect 5602 16533 5637 16544
rect 5123 16510 5154 16533
rect 5196 16510 5223 16533
rect 5269 16510 5292 16533
rect 5342 16510 5361 16533
rect 5415 16510 5430 16533
rect 5488 16510 5499 16533
rect 5561 16510 5568 16533
rect 5634 16510 5637 16533
rect 5671 16533 5706 16544
rect 5740 16533 5775 16544
rect 5809 16533 5844 16544
rect 5878 16533 5913 16544
rect 5947 16533 5982 16544
rect 6016 16533 6051 16544
rect 6085 16533 6120 16544
rect 6154 16533 6189 16544
rect 6223 16533 6258 16544
rect 6292 16533 6327 16544
rect 5671 16510 5673 16533
rect 5740 16510 5746 16533
rect 5809 16510 5819 16533
rect 5878 16510 5892 16533
rect 5947 16510 5965 16533
rect 6016 16510 6038 16533
rect 6085 16510 6110 16533
rect 6154 16510 6182 16533
rect 6223 16510 6254 16533
rect 6292 16510 6326 16533
rect 6361 16510 6396 16544
rect 6430 16533 6465 16544
rect 6499 16533 6534 16544
rect 6568 16533 6603 16544
rect 6637 16533 6672 16544
rect 6706 16533 6741 16544
rect 6775 16533 6810 16544
rect 6844 16533 6879 16544
rect 6913 16533 6948 16544
rect 6982 16533 7017 16544
rect 7051 16533 7086 16544
rect 7120 16533 7155 16544
rect 6432 16510 6465 16533
rect 6504 16510 6534 16533
rect 6576 16510 6603 16533
rect 6648 16510 6672 16533
rect 6720 16510 6741 16533
rect 6792 16510 6810 16533
rect 6864 16510 6879 16533
rect 6936 16510 6948 16533
rect 7008 16510 7017 16533
rect 7080 16510 7086 16533
rect 7152 16510 7155 16533
rect 7189 16533 7224 16544
rect 7189 16510 7190 16533
rect 4681 16499 5089 16510
rect 5123 16499 5162 16510
rect 5196 16499 5235 16510
rect 5269 16499 5308 16510
rect 5342 16499 5381 16510
rect 5415 16499 5454 16510
rect 5488 16499 5527 16510
rect 5561 16499 5600 16510
rect 5634 16499 5673 16510
rect 5707 16499 5746 16510
rect 5780 16499 5819 16510
rect 5853 16499 5892 16510
rect 5926 16499 5965 16510
rect 5999 16499 6038 16510
rect 6072 16499 6110 16510
rect 6144 16499 6182 16510
rect 6216 16499 6254 16510
rect 6288 16499 6326 16510
rect 6360 16499 6398 16510
rect 6432 16499 6470 16510
rect 6504 16499 6542 16510
rect 6576 16499 6614 16510
rect 6648 16499 6686 16510
rect 6720 16499 6758 16510
rect 6792 16499 6830 16510
rect 6864 16499 6902 16510
rect 6936 16499 6974 16510
rect 7008 16499 7046 16510
rect 7080 16499 7118 16510
rect 7152 16499 7190 16510
rect 7258 16533 7293 16544
rect 7327 16533 7362 16544
rect 7396 16533 7431 16544
rect 7465 16533 7500 16544
rect 7534 16533 7568 16544
rect 7602 16533 7636 16544
rect 7670 16533 7704 16544
rect 7738 16533 7772 16544
rect 7806 16533 7840 16544
rect 7258 16510 7262 16533
rect 7327 16510 7334 16533
rect 7396 16510 7406 16533
rect 7465 16510 7478 16533
rect 7534 16510 7550 16533
rect 7602 16510 7622 16533
rect 7670 16510 7694 16533
rect 7738 16510 7766 16533
rect 7806 16510 7838 16533
rect 7874 16510 7908 16544
rect 7224 16499 7262 16510
rect 7296 16499 7334 16510
rect 7368 16499 7406 16510
rect 7440 16499 7478 16510
rect 7512 16499 7550 16510
rect 7584 16499 7622 16510
rect 7656 16499 7694 16510
rect 7728 16499 7766 16510
rect 7800 16499 7838 16510
rect 7872 16499 7908 16510
rect 4681 16484 7908 16499
rect 2648 16480 7908 16484
rect 2648 16446 2663 16480
rect 2697 16446 2735 16480
rect 2769 16446 2807 16480
rect 2841 16446 2879 16480
rect 2913 16446 2951 16480
rect 2985 16446 3023 16480
rect 3057 16446 3095 16480
rect 3129 16446 3167 16480
rect 3201 16446 3239 16480
rect 3273 16446 3311 16480
rect 3345 16446 3383 16480
rect 3417 16446 3455 16480
rect 3489 16446 3527 16480
rect 3561 16446 3599 16480
rect 3633 16446 3671 16480
rect 3705 16446 3743 16480
rect 3777 16446 3815 16480
rect 3849 16446 3887 16480
rect 3921 16446 3959 16480
rect 3993 16446 4031 16480
rect 4065 16446 4103 16480
rect 4137 16446 4175 16480
rect 4209 16446 4247 16480
rect 4281 16446 4319 16480
rect 4353 16446 4391 16480
rect 4425 16446 4463 16480
rect 4497 16446 4535 16480
rect 4569 16474 7908 16480
rect 4569 16446 4740 16474
rect 2648 16440 4740 16446
rect 4774 16440 4809 16474
rect 4843 16440 4878 16474
rect 4912 16440 4947 16474
rect 4981 16440 5016 16474
rect 5050 16440 5085 16474
rect 5119 16457 5154 16474
rect 5188 16457 5223 16474
rect 5257 16457 5292 16474
rect 5326 16457 5361 16474
rect 5395 16457 5430 16474
rect 5464 16457 5499 16474
rect 5533 16457 5568 16474
rect 5602 16457 5637 16474
rect 5123 16440 5154 16457
rect 5196 16440 5223 16457
rect 5269 16440 5292 16457
rect 5342 16440 5361 16457
rect 5415 16440 5430 16457
rect 5488 16440 5499 16457
rect 5561 16440 5568 16457
rect 5634 16440 5637 16457
rect 5671 16457 5706 16474
rect 5740 16457 5775 16474
rect 5809 16457 5844 16474
rect 5878 16457 5913 16474
rect 5947 16457 5982 16474
rect 6016 16457 6051 16474
rect 6085 16457 6120 16474
rect 6154 16457 6189 16474
rect 6223 16457 6258 16474
rect 6292 16457 6327 16474
rect 5671 16440 5673 16457
rect 5740 16440 5746 16457
rect 5809 16440 5819 16457
rect 5878 16440 5892 16457
rect 5947 16440 5965 16457
rect 6016 16440 6038 16457
rect 6085 16440 6110 16457
rect 6154 16440 6182 16457
rect 6223 16440 6254 16457
rect 6292 16440 6326 16457
rect 6361 16440 6396 16474
rect 6430 16457 6465 16474
rect 6499 16457 6534 16474
rect 6568 16457 6603 16474
rect 6637 16457 6672 16474
rect 6706 16457 6741 16474
rect 6775 16457 6810 16474
rect 6844 16457 6879 16474
rect 6913 16457 6948 16474
rect 6982 16457 7017 16474
rect 7051 16457 7086 16474
rect 7120 16457 7155 16474
rect 6432 16440 6465 16457
rect 6504 16440 6534 16457
rect 6576 16440 6603 16457
rect 6648 16440 6672 16457
rect 6720 16440 6741 16457
rect 6792 16440 6810 16457
rect 6864 16440 6879 16457
rect 6936 16440 6948 16457
rect 7008 16440 7017 16457
rect 7080 16440 7086 16457
rect 7152 16440 7155 16457
rect 7189 16457 7224 16474
rect 7189 16440 7190 16457
rect 2648 16423 5089 16440
rect 5123 16423 5162 16440
rect 5196 16423 5235 16440
rect 5269 16423 5308 16440
rect 5342 16423 5381 16440
rect 5415 16423 5454 16440
rect 5488 16423 5527 16440
rect 5561 16423 5600 16440
rect 5634 16423 5673 16440
rect 5707 16423 5746 16440
rect 5780 16423 5819 16440
rect 5853 16423 5892 16440
rect 5926 16423 5965 16440
rect 5999 16423 6038 16440
rect 6072 16423 6110 16440
rect 6144 16423 6182 16440
rect 6216 16423 6254 16440
rect 6288 16423 6326 16440
rect 6360 16423 6398 16440
rect 6432 16423 6470 16440
rect 6504 16423 6542 16440
rect 6576 16423 6614 16440
rect 6648 16423 6686 16440
rect 6720 16423 6758 16440
rect 6792 16423 6830 16440
rect 6864 16423 6902 16440
rect 6936 16423 6974 16440
rect 7008 16423 7046 16440
rect 7080 16423 7118 16440
rect 7152 16423 7190 16440
rect 7258 16457 7293 16474
rect 7327 16457 7362 16474
rect 7396 16457 7431 16474
rect 7465 16457 7500 16474
rect 7534 16457 7568 16474
rect 7602 16457 7636 16474
rect 7670 16457 7704 16474
rect 7738 16457 7772 16474
rect 7806 16457 7840 16474
rect 7258 16440 7262 16457
rect 7327 16440 7334 16457
rect 7396 16440 7406 16457
rect 7465 16440 7478 16457
rect 7534 16440 7550 16457
rect 7602 16440 7622 16457
rect 7670 16440 7694 16457
rect 7738 16440 7766 16457
rect 7806 16440 7838 16457
rect 7874 16440 7908 16474
rect 7224 16423 7262 16440
rect 7296 16423 7334 16440
rect 7368 16423 7406 16440
rect 7440 16423 7478 16440
rect 7512 16423 7550 16440
rect 7584 16423 7622 16440
rect 7656 16423 7694 16440
rect 7728 16423 7766 16440
rect 7800 16423 7838 16440
rect 7872 16423 7908 16440
rect 2648 16407 7908 16423
rect 2648 16373 2663 16407
rect 2697 16381 2735 16407
rect 2697 16373 2715 16381
rect 2769 16373 2807 16407
rect 2841 16381 2879 16407
rect 2841 16373 2853 16381
rect 2913 16373 2951 16407
rect 2985 16381 3023 16407
rect 2985 16373 2991 16381
rect 3057 16373 3095 16407
rect 3129 16381 3167 16407
rect 2648 16347 2715 16373
rect 2749 16347 2853 16373
rect 2887 16347 2991 16373
rect 3025 16347 3129 16373
rect 3163 16373 3167 16381
rect 3201 16373 3239 16407
rect 3273 16381 3311 16407
rect 3301 16373 3311 16381
rect 3345 16373 3383 16407
rect 3417 16381 3455 16407
rect 3439 16373 3455 16381
rect 3489 16373 3527 16407
rect 3561 16381 3599 16407
rect 3577 16373 3599 16381
rect 3633 16373 3671 16407
rect 3705 16381 3743 16407
rect 3715 16373 3743 16381
rect 3777 16373 3815 16407
rect 3849 16381 3887 16407
rect 3853 16373 3887 16381
rect 3921 16381 3959 16407
rect 3921 16373 3957 16381
rect 3993 16373 4031 16407
rect 4065 16381 4103 16407
rect 4065 16373 4095 16381
rect 4137 16373 4175 16407
rect 4209 16381 4247 16407
rect 4209 16373 4233 16381
rect 4281 16373 4319 16407
rect 4353 16381 4391 16407
rect 4353 16373 4371 16381
rect 4425 16373 4463 16407
rect 4497 16381 4535 16407
rect 4569 16404 7908 16407
rect 4569 16381 4740 16404
rect 4497 16373 4509 16381
rect 4569 16373 4647 16381
rect 3163 16347 3267 16373
rect 3301 16347 3405 16373
rect 3439 16347 3543 16373
rect 3577 16347 3681 16373
rect 3715 16347 3819 16373
rect 3853 16347 3957 16373
rect 3991 16347 4095 16373
rect 4129 16347 4233 16373
rect 4267 16347 4371 16373
rect 4405 16347 4509 16373
rect 4543 16347 4647 16373
rect 4681 16370 4740 16381
rect 4774 16370 4809 16404
rect 4843 16370 4878 16404
rect 4912 16370 4947 16404
rect 4981 16370 5016 16404
rect 5050 16370 5085 16404
rect 5119 16381 5154 16404
rect 5188 16381 5223 16404
rect 5257 16381 5292 16404
rect 5326 16381 5361 16404
rect 5395 16381 5430 16404
rect 5464 16381 5499 16404
rect 5533 16381 5568 16404
rect 5602 16381 5637 16404
rect 5123 16370 5154 16381
rect 5196 16370 5223 16381
rect 5269 16370 5292 16381
rect 5342 16370 5361 16381
rect 5415 16370 5430 16381
rect 5488 16370 5499 16381
rect 5561 16370 5568 16381
rect 5634 16370 5637 16381
rect 5671 16381 5706 16404
rect 5740 16381 5775 16404
rect 5809 16381 5844 16404
rect 5878 16381 5913 16404
rect 5947 16381 5982 16404
rect 6016 16381 6051 16404
rect 6085 16381 6120 16404
rect 6154 16381 6189 16404
rect 6223 16381 6258 16404
rect 6292 16381 6327 16404
rect 5671 16370 5673 16381
rect 5740 16370 5746 16381
rect 5809 16370 5819 16381
rect 5878 16370 5892 16381
rect 5947 16370 5965 16381
rect 6016 16370 6038 16381
rect 6085 16370 6110 16381
rect 6154 16370 6182 16381
rect 6223 16370 6254 16381
rect 6292 16370 6326 16381
rect 6361 16370 6396 16404
rect 6430 16381 6465 16404
rect 6499 16381 6534 16404
rect 6568 16381 6603 16404
rect 6637 16381 6672 16404
rect 6706 16381 6741 16404
rect 6775 16381 6810 16404
rect 6844 16381 6879 16404
rect 6913 16381 6948 16404
rect 6982 16381 7017 16404
rect 7051 16381 7086 16404
rect 7120 16381 7155 16404
rect 6432 16370 6465 16381
rect 6504 16370 6534 16381
rect 6576 16370 6603 16381
rect 6648 16370 6672 16381
rect 6720 16370 6741 16381
rect 6792 16370 6810 16381
rect 6864 16370 6879 16381
rect 6936 16370 6948 16381
rect 7008 16370 7017 16381
rect 7080 16370 7086 16381
rect 7152 16370 7155 16381
rect 7189 16381 7224 16404
rect 7189 16370 7190 16381
rect 4681 16347 5089 16370
rect 5123 16347 5162 16370
rect 5196 16347 5235 16370
rect 5269 16347 5308 16370
rect 5342 16347 5381 16370
rect 5415 16347 5454 16370
rect 5488 16347 5527 16370
rect 5561 16347 5600 16370
rect 5634 16347 5673 16370
rect 5707 16347 5746 16370
rect 5780 16347 5819 16370
rect 5853 16347 5892 16370
rect 5926 16347 5965 16370
rect 5999 16347 6038 16370
rect 6072 16347 6110 16370
rect 6144 16347 6182 16370
rect 6216 16347 6254 16370
rect 6288 16347 6326 16370
rect 6360 16347 6398 16370
rect 6432 16347 6470 16370
rect 6504 16347 6542 16370
rect 6576 16347 6614 16370
rect 6648 16347 6686 16370
rect 6720 16347 6758 16370
rect 6792 16347 6830 16370
rect 6864 16347 6902 16370
rect 6936 16347 6974 16370
rect 7008 16347 7046 16370
rect 7080 16347 7118 16370
rect 7152 16347 7190 16370
rect 7258 16381 7293 16404
rect 7327 16381 7362 16404
rect 7396 16381 7431 16404
rect 7465 16381 7500 16404
rect 7534 16381 7568 16404
rect 7602 16381 7636 16404
rect 7670 16381 7704 16404
rect 7738 16381 7772 16404
rect 7806 16381 7840 16404
rect 7258 16370 7262 16381
rect 7327 16370 7334 16381
rect 7396 16370 7406 16381
rect 7465 16370 7478 16381
rect 7534 16370 7550 16381
rect 7602 16370 7622 16381
rect 7670 16370 7694 16381
rect 7738 16370 7766 16381
rect 7806 16370 7838 16381
rect 7874 16370 7908 16404
rect 7224 16347 7262 16370
rect 7296 16347 7334 16370
rect 7368 16347 7406 16370
rect 7440 16347 7478 16370
rect 7512 16347 7550 16370
rect 7584 16347 7622 16370
rect 7656 16347 7694 16370
rect 7728 16347 7766 16370
rect 7800 16347 7838 16370
rect 7872 16347 7908 16370
rect 2648 16334 7908 16347
rect 2648 16300 2663 16334
rect 2697 16300 2735 16334
rect 2769 16300 2807 16334
rect 2841 16300 2879 16334
rect 2913 16300 2951 16334
rect 2985 16300 3023 16334
rect 3057 16300 3095 16334
rect 3129 16300 3167 16334
rect 3201 16300 3239 16334
rect 3273 16300 3311 16334
rect 3345 16300 3383 16334
rect 3417 16300 3455 16334
rect 3489 16300 3527 16334
rect 3561 16300 3599 16334
rect 3633 16300 3671 16334
rect 3705 16300 3743 16334
rect 3777 16300 3815 16334
rect 3849 16300 3887 16334
rect 3921 16300 3959 16334
rect 3993 16300 4031 16334
rect 4065 16300 4103 16334
rect 4137 16300 4175 16334
rect 4209 16300 4247 16334
rect 4281 16300 4319 16334
rect 4353 16300 4391 16334
rect 4425 16300 4463 16334
rect 4497 16300 4535 16334
rect 4569 16300 4740 16334
rect 4774 16300 4809 16334
rect 4843 16300 4878 16334
rect 4912 16300 4947 16334
rect 4981 16300 5016 16334
rect 5050 16300 5085 16334
rect 5119 16305 5154 16334
rect 5188 16305 5223 16334
rect 5257 16305 5292 16334
rect 5326 16305 5361 16334
rect 5395 16305 5430 16334
rect 5464 16305 5499 16334
rect 5533 16305 5568 16334
rect 5602 16305 5637 16334
rect 5123 16300 5154 16305
rect 5196 16300 5223 16305
rect 5269 16300 5292 16305
rect 5342 16300 5361 16305
rect 5415 16300 5430 16305
rect 5488 16300 5499 16305
rect 5561 16300 5568 16305
rect 5634 16300 5637 16305
rect 5671 16305 5706 16334
rect 5740 16305 5775 16334
rect 5809 16305 5844 16334
rect 5878 16305 5913 16334
rect 5947 16305 5982 16334
rect 6016 16305 6051 16334
rect 6085 16305 6120 16334
rect 6154 16305 6189 16334
rect 6223 16305 6258 16334
rect 6292 16305 6327 16334
rect 5671 16300 5673 16305
rect 5740 16300 5746 16305
rect 5809 16300 5819 16305
rect 5878 16300 5892 16305
rect 5947 16300 5965 16305
rect 6016 16300 6038 16305
rect 6085 16300 6110 16305
rect 6154 16300 6182 16305
rect 6223 16300 6254 16305
rect 6292 16300 6326 16305
rect 6361 16300 6396 16334
rect 6430 16305 6465 16334
rect 6499 16305 6534 16334
rect 6568 16305 6603 16334
rect 6637 16305 6672 16334
rect 6706 16305 6741 16334
rect 6775 16305 6810 16334
rect 6844 16305 6879 16334
rect 6913 16305 6948 16334
rect 6982 16305 7017 16334
rect 7051 16305 7086 16334
rect 7120 16305 7155 16334
rect 6432 16300 6465 16305
rect 6504 16300 6534 16305
rect 6576 16300 6603 16305
rect 6648 16300 6672 16305
rect 6720 16300 6741 16305
rect 6792 16300 6810 16305
rect 6864 16300 6879 16305
rect 6936 16300 6948 16305
rect 7008 16300 7017 16305
rect 7080 16300 7086 16305
rect 7152 16300 7155 16305
rect 7189 16305 7224 16334
rect 7189 16300 7190 16305
rect 2648 16271 5089 16300
rect 5123 16271 5162 16300
rect 5196 16271 5235 16300
rect 5269 16271 5308 16300
rect 5342 16271 5381 16300
rect 5415 16271 5454 16300
rect 5488 16271 5527 16300
rect 5561 16271 5600 16300
rect 5634 16271 5673 16300
rect 5707 16271 5746 16300
rect 5780 16271 5819 16300
rect 5853 16271 5892 16300
rect 5926 16271 5965 16300
rect 5999 16271 6038 16300
rect 6072 16271 6110 16300
rect 6144 16271 6182 16300
rect 6216 16271 6254 16300
rect 6288 16271 6326 16300
rect 6360 16271 6398 16300
rect 6432 16271 6470 16300
rect 6504 16271 6542 16300
rect 6576 16271 6614 16300
rect 6648 16271 6686 16300
rect 6720 16271 6758 16300
rect 6792 16271 6830 16300
rect 6864 16271 6902 16300
rect 6936 16271 6974 16300
rect 7008 16271 7046 16300
rect 7080 16271 7118 16300
rect 7152 16271 7190 16300
rect 7258 16305 7293 16334
rect 7327 16305 7362 16334
rect 7396 16305 7431 16334
rect 7465 16305 7500 16334
rect 7534 16305 7568 16334
rect 7602 16305 7636 16334
rect 7670 16305 7704 16334
rect 7738 16305 7772 16334
rect 7806 16305 7840 16334
rect 7258 16300 7262 16305
rect 7327 16300 7334 16305
rect 7396 16300 7406 16305
rect 7465 16300 7478 16305
rect 7534 16300 7550 16305
rect 7602 16300 7622 16305
rect 7670 16300 7694 16305
rect 7738 16300 7766 16305
rect 7806 16300 7838 16305
rect 7874 16300 7908 16334
rect 7224 16271 7262 16300
rect 7296 16271 7334 16300
rect 7368 16271 7406 16300
rect 7440 16271 7478 16300
rect 7512 16271 7550 16300
rect 7584 16271 7622 16300
rect 7656 16271 7694 16300
rect 7728 16271 7766 16300
rect 7800 16271 7838 16300
rect 7872 16271 7908 16300
rect 2648 16264 7908 16271
rect 2648 16261 4740 16264
rect 2648 16227 2663 16261
rect 2697 16244 2735 16261
rect 2697 16227 2715 16244
rect 2769 16227 2807 16261
rect 2841 16244 2879 16261
rect 2841 16227 2853 16244
rect 2913 16227 2951 16261
rect 2985 16244 3023 16261
rect 2985 16227 2991 16244
rect 3057 16227 3095 16261
rect 3129 16244 3167 16261
rect 2648 16210 2715 16227
rect 2749 16210 2853 16227
rect 2887 16210 2991 16227
rect 3025 16210 3129 16227
rect 3163 16227 3167 16244
rect 3201 16227 3239 16261
rect 3273 16244 3311 16261
rect 3301 16227 3311 16244
rect 3345 16227 3383 16261
rect 3417 16244 3455 16261
rect 3439 16227 3455 16244
rect 3489 16227 3527 16261
rect 3561 16244 3599 16261
rect 3577 16227 3599 16244
rect 3633 16227 3671 16261
rect 3705 16244 3743 16261
rect 3715 16227 3743 16244
rect 3777 16227 3815 16261
rect 3849 16244 3887 16261
rect 3853 16227 3887 16244
rect 3921 16244 3959 16261
rect 3921 16227 3957 16244
rect 3993 16227 4031 16261
rect 4065 16244 4103 16261
rect 4065 16227 4095 16244
rect 4137 16227 4175 16261
rect 4209 16244 4247 16261
rect 4209 16227 4233 16244
rect 4281 16227 4319 16261
rect 4353 16244 4391 16261
rect 4353 16227 4371 16244
rect 4425 16227 4463 16261
rect 4497 16244 4535 16261
rect 4569 16244 4740 16261
rect 4497 16227 4509 16244
rect 4569 16227 4647 16244
rect 3163 16210 3267 16227
rect 3301 16210 3405 16227
rect 3439 16210 3543 16227
rect 3577 16210 3681 16227
rect 3715 16210 3819 16227
rect 3853 16210 3957 16227
rect 3991 16210 4095 16227
rect 4129 16210 4233 16227
rect 4267 16210 4371 16227
rect 4405 16210 4509 16227
rect 4543 16210 4647 16227
rect 4681 16230 4740 16244
rect 4774 16230 4809 16264
rect 4843 16230 4878 16264
rect 4912 16230 4947 16264
rect 4981 16230 5016 16264
rect 5050 16230 5085 16264
rect 5119 16230 5154 16264
rect 5188 16230 5223 16264
rect 5257 16230 5292 16264
rect 5326 16230 5361 16264
rect 5395 16230 5430 16264
rect 5464 16230 5499 16264
rect 5533 16230 5568 16264
rect 5602 16230 5637 16264
rect 5671 16230 5706 16264
rect 5740 16230 5775 16264
rect 5809 16230 5844 16264
rect 5878 16230 5913 16264
rect 5947 16230 5982 16264
rect 6016 16230 6051 16264
rect 6085 16230 6120 16264
rect 6154 16230 6189 16264
rect 6223 16230 6258 16264
rect 6292 16230 6327 16264
rect 6361 16230 6396 16264
rect 6430 16230 6465 16264
rect 6499 16230 6534 16264
rect 6568 16230 6603 16264
rect 6637 16230 6672 16264
rect 6706 16230 6741 16264
rect 6775 16230 6810 16264
rect 6844 16230 6879 16264
rect 6913 16230 6948 16264
rect 6982 16230 7017 16264
rect 7051 16230 7086 16264
rect 7120 16230 7155 16264
rect 7189 16230 7224 16264
rect 7258 16230 7293 16264
rect 7327 16230 7362 16264
rect 7396 16230 7431 16264
rect 7465 16230 7500 16264
rect 7534 16230 7568 16264
rect 7602 16230 7636 16264
rect 7670 16230 7704 16264
rect 7738 16230 7772 16264
rect 7806 16230 7840 16264
rect 7874 16230 7908 16264
rect 4681 16229 7908 16230
rect 4681 16210 5089 16229
rect 2648 16195 5089 16210
rect 5123 16195 5162 16229
rect 5196 16195 5235 16229
rect 5269 16195 5308 16229
rect 5342 16195 5381 16229
rect 5415 16195 5454 16229
rect 5488 16195 5527 16229
rect 5561 16195 5600 16229
rect 5634 16195 5673 16229
rect 5707 16195 5746 16229
rect 5780 16195 5819 16229
rect 5853 16195 5892 16229
rect 5926 16195 5965 16229
rect 5999 16195 6038 16229
rect 6072 16195 6110 16229
rect 6144 16195 6182 16229
rect 6216 16195 6254 16229
rect 6288 16195 6326 16229
rect 6360 16195 6398 16229
rect 6432 16195 6470 16229
rect 6504 16195 6542 16229
rect 6576 16195 6614 16229
rect 6648 16195 6686 16229
rect 6720 16195 6758 16229
rect 6792 16195 6830 16229
rect 6864 16195 6902 16229
rect 6936 16195 6974 16229
rect 7008 16195 7046 16229
rect 7080 16195 7118 16229
rect 7152 16195 7190 16229
rect 7224 16195 7262 16229
rect 7296 16195 7334 16229
rect 7368 16195 7406 16229
rect 7440 16195 7478 16229
rect 7512 16195 7550 16229
rect 7584 16195 7622 16229
rect 7656 16195 7694 16229
rect 7728 16195 7766 16229
rect 7800 16195 7838 16229
rect 7872 16195 7908 16229
rect 2648 16194 7908 16195
rect 2648 16188 4740 16194
rect 2648 16154 2663 16188
rect 2697 16154 2735 16188
rect 2769 16154 2807 16188
rect 2841 16154 2879 16188
rect 2913 16154 2951 16188
rect 2985 16154 3023 16188
rect 3057 16154 3095 16188
rect 3129 16154 3167 16188
rect 3201 16154 3239 16188
rect 3273 16154 3311 16188
rect 3345 16154 3383 16188
rect 3417 16154 3455 16188
rect 3489 16154 3527 16188
rect 3561 16154 3599 16188
rect 3633 16154 3671 16188
rect 3705 16154 3743 16188
rect 3777 16154 3815 16188
rect 3849 16154 3887 16188
rect 3921 16154 3959 16188
rect 3993 16154 4031 16188
rect 4065 16154 4103 16188
rect 4137 16154 4175 16188
rect 4209 16154 4247 16188
rect 4281 16154 4319 16188
rect 4353 16154 4391 16188
rect 4425 16154 4463 16188
rect 4497 16154 4535 16188
rect 4569 16160 4740 16188
rect 4774 16160 4809 16194
rect 4843 16160 4878 16194
rect 4912 16160 4947 16194
rect 4981 16160 5016 16194
rect 5050 16160 5085 16194
rect 5119 16160 5154 16194
rect 5188 16160 5223 16194
rect 5257 16160 5292 16194
rect 5326 16160 5361 16194
rect 5395 16160 5430 16194
rect 5464 16160 5499 16194
rect 5533 16160 5568 16194
rect 5602 16160 5637 16194
rect 5671 16160 5706 16194
rect 5740 16160 5775 16194
rect 5809 16160 5844 16194
rect 5878 16160 5913 16194
rect 5947 16160 5982 16194
rect 6016 16160 6051 16194
rect 6085 16160 6120 16194
rect 6154 16160 6189 16194
rect 6223 16160 6258 16194
rect 6292 16160 6327 16194
rect 6361 16160 6396 16194
rect 6430 16160 6465 16194
rect 6499 16160 6534 16194
rect 6568 16160 6603 16194
rect 6637 16160 6672 16194
rect 6706 16160 6741 16194
rect 6775 16160 6810 16194
rect 6844 16160 6879 16194
rect 6913 16160 6948 16194
rect 6982 16160 7017 16194
rect 7051 16160 7086 16194
rect 7120 16160 7155 16194
rect 7189 16160 7224 16194
rect 7258 16160 7293 16194
rect 7327 16160 7362 16194
rect 7396 16160 7431 16194
rect 7465 16160 7500 16194
rect 7534 16160 7568 16194
rect 7602 16160 7636 16194
rect 7670 16160 7704 16194
rect 7738 16160 7772 16194
rect 7806 16160 7840 16194
rect 7874 16160 7908 16194
rect 4569 16154 7908 16160
rect 2648 16153 7908 16154
rect 2648 16124 5089 16153
rect 5123 16124 5162 16153
rect 5196 16124 5235 16153
rect 5269 16124 5308 16153
rect 5342 16124 5381 16153
rect 5415 16124 5454 16153
rect 5488 16124 5527 16153
rect 5561 16124 5600 16153
rect 5634 16124 5673 16153
rect 5707 16124 5746 16153
rect 5780 16124 5819 16153
rect 5853 16124 5892 16153
rect 5926 16124 5965 16153
rect 5999 16124 6038 16153
rect 6072 16124 6110 16153
rect 6144 16124 6182 16153
rect 6216 16124 6254 16153
rect 6288 16124 6326 16153
rect 6360 16124 6398 16153
rect 6432 16124 6470 16153
rect 6504 16124 6542 16153
rect 6576 16124 6614 16153
rect 6648 16124 6686 16153
rect 6720 16124 6758 16153
rect 6792 16124 6830 16153
rect 6864 16124 6902 16153
rect 6936 16124 6974 16153
rect 7008 16124 7046 16153
rect 7080 16124 7118 16153
rect 7152 16124 7190 16153
rect 2648 16115 4740 16124
rect 2648 16081 2663 16115
rect 2697 16107 2735 16115
rect 2697 16081 2715 16107
rect 2769 16081 2807 16115
rect 2841 16107 2879 16115
rect 2841 16081 2853 16107
rect 2913 16081 2951 16115
rect 2985 16107 3023 16115
rect 2985 16081 2991 16107
rect 3057 16081 3095 16115
rect 3129 16107 3167 16115
rect 2648 16073 2715 16081
rect 2749 16073 2853 16081
rect 2887 16073 2991 16081
rect 3025 16073 3129 16081
rect 3163 16081 3167 16107
rect 3201 16081 3239 16115
rect 3273 16107 3311 16115
rect 3301 16081 3311 16107
rect 3345 16081 3383 16115
rect 3417 16107 3455 16115
rect 3439 16081 3455 16107
rect 3489 16081 3527 16115
rect 3561 16107 3599 16115
rect 3577 16081 3599 16107
rect 3633 16081 3671 16115
rect 3705 16107 3743 16115
rect 3715 16081 3743 16107
rect 3777 16081 3815 16115
rect 3849 16107 3887 16115
rect 3853 16081 3887 16107
rect 3921 16107 3959 16115
rect 3921 16081 3957 16107
rect 3993 16081 4031 16115
rect 4065 16107 4103 16115
rect 4065 16081 4095 16107
rect 4137 16081 4175 16115
rect 4209 16107 4247 16115
rect 4209 16081 4233 16107
rect 4281 16081 4319 16115
rect 4353 16107 4391 16115
rect 4353 16081 4371 16107
rect 4425 16081 4463 16115
rect 4497 16107 4535 16115
rect 4569 16107 4740 16115
rect 4497 16081 4509 16107
rect 4569 16081 4647 16107
rect 3163 16073 3267 16081
rect 3301 16073 3405 16081
rect 3439 16073 3543 16081
rect 3577 16073 3681 16081
rect 3715 16073 3819 16081
rect 3853 16073 3957 16081
rect 3991 16073 4095 16081
rect 4129 16073 4233 16081
rect 4267 16073 4371 16081
rect 4405 16073 4509 16081
rect 4543 16073 4647 16081
rect 4681 16090 4740 16107
rect 4774 16090 4809 16124
rect 4843 16090 4878 16124
rect 4912 16090 4947 16124
rect 4981 16090 5016 16124
rect 5050 16090 5085 16124
rect 5123 16119 5154 16124
rect 5196 16119 5223 16124
rect 5269 16119 5292 16124
rect 5342 16119 5361 16124
rect 5415 16119 5430 16124
rect 5488 16119 5499 16124
rect 5561 16119 5568 16124
rect 5634 16119 5637 16124
rect 5119 16090 5154 16119
rect 5188 16090 5223 16119
rect 5257 16090 5292 16119
rect 5326 16090 5361 16119
rect 5395 16090 5430 16119
rect 5464 16090 5499 16119
rect 5533 16090 5568 16119
rect 5602 16090 5637 16119
rect 5671 16119 5673 16124
rect 5740 16119 5746 16124
rect 5809 16119 5819 16124
rect 5878 16119 5892 16124
rect 5947 16119 5965 16124
rect 6016 16119 6038 16124
rect 6085 16119 6110 16124
rect 6154 16119 6182 16124
rect 6223 16119 6254 16124
rect 6292 16119 6326 16124
rect 5671 16090 5706 16119
rect 5740 16090 5775 16119
rect 5809 16090 5844 16119
rect 5878 16090 5913 16119
rect 5947 16090 5982 16119
rect 6016 16090 6051 16119
rect 6085 16090 6120 16119
rect 6154 16090 6189 16119
rect 6223 16090 6258 16119
rect 6292 16090 6327 16119
rect 6361 16090 6396 16124
rect 6432 16119 6465 16124
rect 6504 16119 6534 16124
rect 6576 16119 6603 16124
rect 6648 16119 6672 16124
rect 6720 16119 6741 16124
rect 6792 16119 6810 16124
rect 6864 16119 6879 16124
rect 6936 16119 6948 16124
rect 7008 16119 7017 16124
rect 7080 16119 7086 16124
rect 7152 16119 7155 16124
rect 6430 16090 6465 16119
rect 6499 16090 6534 16119
rect 6568 16090 6603 16119
rect 6637 16090 6672 16119
rect 6706 16090 6741 16119
rect 6775 16090 6810 16119
rect 6844 16090 6879 16119
rect 6913 16090 6948 16119
rect 6982 16090 7017 16119
rect 7051 16090 7086 16119
rect 7120 16090 7155 16119
rect 7189 16119 7190 16124
rect 7224 16124 7262 16153
rect 7296 16124 7334 16153
rect 7368 16124 7406 16153
rect 7440 16124 7478 16153
rect 7512 16124 7550 16153
rect 7584 16124 7622 16153
rect 7656 16124 7694 16153
rect 7728 16124 7766 16153
rect 7800 16124 7838 16153
rect 7872 16124 7908 16153
rect 7189 16090 7224 16119
rect 7258 16119 7262 16124
rect 7327 16119 7334 16124
rect 7396 16119 7406 16124
rect 7465 16119 7478 16124
rect 7534 16119 7550 16124
rect 7602 16119 7622 16124
rect 7670 16119 7694 16124
rect 7738 16119 7766 16124
rect 7806 16119 7838 16124
rect 7258 16090 7293 16119
rect 7327 16090 7362 16119
rect 7396 16090 7431 16119
rect 7465 16090 7500 16119
rect 7534 16090 7568 16119
rect 7602 16090 7636 16119
rect 7670 16090 7704 16119
rect 7738 16090 7772 16119
rect 7806 16090 7840 16119
rect 7874 16090 7908 16124
rect 4681 16077 7908 16090
rect 4681 16073 5089 16077
rect 2648 16054 5089 16073
rect 5123 16054 5162 16077
rect 5196 16054 5235 16077
rect 5269 16054 5308 16077
rect 5342 16054 5381 16077
rect 5415 16054 5454 16077
rect 5488 16054 5527 16077
rect 5561 16054 5600 16077
rect 5634 16054 5673 16077
rect 5707 16054 5746 16077
rect 5780 16054 5819 16077
rect 5853 16054 5892 16077
rect 5926 16054 5965 16077
rect 5999 16054 6038 16077
rect 6072 16054 6110 16077
rect 6144 16054 6182 16077
rect 6216 16054 6254 16077
rect 6288 16054 6326 16077
rect 6360 16054 6398 16077
rect 6432 16054 6470 16077
rect 6504 16054 6542 16077
rect 6576 16054 6614 16077
rect 6648 16054 6686 16077
rect 6720 16054 6758 16077
rect 6792 16054 6830 16077
rect 6864 16054 6902 16077
rect 6936 16054 6974 16077
rect 7008 16054 7046 16077
rect 7080 16054 7118 16077
rect 7152 16054 7190 16077
rect 2648 16042 4740 16054
rect 2648 16008 2663 16042
rect 2697 16008 2735 16042
rect 2769 16008 2807 16042
rect 2841 16008 2879 16042
rect 2913 16008 2951 16042
rect 2985 16008 3023 16042
rect 3057 16008 3095 16042
rect 3129 16008 3167 16042
rect 3201 16008 3239 16042
rect 3273 16008 3311 16042
rect 3345 16008 3383 16042
rect 3417 16008 3455 16042
rect 3489 16008 3527 16042
rect 3561 16008 3599 16042
rect 3633 16008 3671 16042
rect 3705 16008 3743 16042
rect 3777 16008 3815 16042
rect 3849 16008 3887 16042
rect 3921 16008 3959 16042
rect 3993 16008 4031 16042
rect 4065 16008 4103 16042
rect 4137 16008 4175 16042
rect 4209 16008 4247 16042
rect 4281 16008 4319 16042
rect 4353 16008 4391 16042
rect 4425 16008 4463 16042
rect 4497 16008 4535 16042
rect 4569 16020 4740 16042
rect 4774 16020 4809 16054
rect 4843 16020 4878 16054
rect 4912 16020 4947 16054
rect 4981 16020 5016 16054
rect 5050 16020 5085 16054
rect 5123 16043 5154 16054
rect 5196 16043 5223 16054
rect 5269 16043 5292 16054
rect 5342 16043 5361 16054
rect 5415 16043 5430 16054
rect 5488 16043 5499 16054
rect 5561 16043 5568 16054
rect 5634 16043 5637 16054
rect 5119 16020 5154 16043
rect 5188 16020 5223 16043
rect 5257 16020 5292 16043
rect 5326 16020 5361 16043
rect 5395 16020 5430 16043
rect 5464 16020 5499 16043
rect 5533 16020 5568 16043
rect 5602 16020 5637 16043
rect 5671 16043 5673 16054
rect 5740 16043 5746 16054
rect 5809 16043 5819 16054
rect 5878 16043 5892 16054
rect 5947 16043 5965 16054
rect 6016 16043 6038 16054
rect 6085 16043 6110 16054
rect 6154 16043 6182 16054
rect 6223 16043 6254 16054
rect 6292 16043 6326 16054
rect 5671 16020 5706 16043
rect 5740 16020 5775 16043
rect 5809 16020 5844 16043
rect 5878 16020 5913 16043
rect 5947 16020 5982 16043
rect 6016 16020 6051 16043
rect 6085 16020 6120 16043
rect 6154 16020 6189 16043
rect 6223 16020 6258 16043
rect 6292 16020 6327 16043
rect 6361 16020 6396 16054
rect 6432 16043 6465 16054
rect 6504 16043 6534 16054
rect 6576 16043 6603 16054
rect 6648 16043 6672 16054
rect 6720 16043 6741 16054
rect 6792 16043 6810 16054
rect 6864 16043 6879 16054
rect 6936 16043 6948 16054
rect 7008 16043 7017 16054
rect 7080 16043 7086 16054
rect 7152 16043 7155 16054
rect 6430 16020 6465 16043
rect 6499 16020 6534 16043
rect 6568 16020 6603 16043
rect 6637 16020 6672 16043
rect 6706 16020 6741 16043
rect 6775 16020 6810 16043
rect 6844 16020 6879 16043
rect 6913 16020 6948 16043
rect 6982 16020 7017 16043
rect 7051 16020 7086 16043
rect 7120 16020 7155 16043
rect 7189 16043 7190 16054
rect 7224 16054 7262 16077
rect 7296 16054 7334 16077
rect 7368 16054 7406 16077
rect 7440 16054 7478 16077
rect 7512 16054 7550 16077
rect 7584 16054 7622 16077
rect 7656 16054 7694 16077
rect 7728 16054 7766 16077
rect 7800 16054 7838 16077
rect 7872 16054 7908 16077
rect 7189 16020 7224 16043
rect 7258 16043 7262 16054
rect 7327 16043 7334 16054
rect 7396 16043 7406 16054
rect 7465 16043 7478 16054
rect 7534 16043 7550 16054
rect 7602 16043 7622 16054
rect 7670 16043 7694 16054
rect 7738 16043 7766 16054
rect 7806 16043 7838 16054
rect 7258 16020 7293 16043
rect 7327 16020 7362 16043
rect 7396 16020 7431 16043
rect 7465 16020 7500 16043
rect 7534 16020 7568 16043
rect 7602 16020 7636 16043
rect 7670 16020 7704 16043
rect 7738 16020 7772 16043
rect 7806 16020 7840 16043
rect 7874 16020 7908 16054
rect 4569 16008 7908 16020
rect 2648 16001 7908 16008
rect 2648 15984 5089 16001
rect 5123 15984 5162 16001
rect 5196 15984 5235 16001
rect 5269 15984 5308 16001
rect 5342 15984 5381 16001
rect 5415 15984 5454 16001
rect 5488 15984 5527 16001
rect 5561 15984 5600 16001
rect 5634 15984 5673 16001
rect 5707 15984 5746 16001
rect 5780 15984 5819 16001
rect 5853 15984 5892 16001
rect 5926 15984 5965 16001
rect 5999 15984 6038 16001
rect 6072 15984 6110 16001
rect 6144 15984 6182 16001
rect 6216 15984 6254 16001
rect 6288 15984 6326 16001
rect 6360 15984 6398 16001
rect 6432 15984 6470 16001
rect 6504 15984 6542 16001
rect 6576 15984 6614 16001
rect 6648 15984 6686 16001
rect 6720 15984 6758 16001
rect 6792 15984 6830 16001
rect 6864 15984 6902 16001
rect 6936 15984 6974 16001
rect 7008 15984 7046 16001
rect 7080 15984 7118 16001
rect 7152 15984 7190 16001
rect 2648 15970 4740 15984
rect 2648 15969 2715 15970
rect 2749 15969 2853 15970
rect 2887 15969 2991 15970
rect 3025 15969 3129 15970
rect 2648 15935 2663 15969
rect 2697 15936 2715 15969
rect 2697 15935 2735 15936
rect 2769 15935 2807 15969
rect 2841 15936 2853 15969
rect 2841 15935 2879 15936
rect 2913 15935 2951 15969
rect 2985 15936 2991 15969
rect 2985 15935 3023 15936
rect 3057 15935 3095 15969
rect 3163 15969 3267 15970
rect 3301 15969 3405 15970
rect 3439 15969 3543 15970
rect 3577 15969 3681 15970
rect 3715 15969 3819 15970
rect 3853 15969 3957 15970
rect 3991 15969 4095 15970
rect 4129 15969 4233 15970
rect 4267 15969 4371 15970
rect 4405 15969 4509 15970
rect 4543 15969 4647 15970
rect 3163 15936 3167 15969
rect 3129 15935 3167 15936
rect 3201 15935 3239 15969
rect 3301 15936 3311 15969
rect 3273 15935 3311 15936
rect 3345 15935 3383 15969
rect 3439 15936 3455 15969
rect 3417 15935 3455 15936
rect 3489 15935 3527 15969
rect 3577 15936 3599 15969
rect 3561 15935 3599 15936
rect 3633 15935 3671 15969
rect 3715 15936 3743 15969
rect 3705 15935 3743 15936
rect 3777 15935 3815 15969
rect 3853 15936 3887 15969
rect 3849 15935 3887 15936
rect 3921 15936 3957 15969
rect 3921 15935 3959 15936
rect 3993 15935 4031 15969
rect 4065 15936 4095 15969
rect 4065 15935 4103 15936
rect 4137 15935 4175 15969
rect 4209 15936 4233 15969
rect 4209 15935 4247 15936
rect 4281 15935 4319 15969
rect 4353 15936 4371 15969
rect 4353 15935 4391 15936
rect 4425 15935 4463 15969
rect 4497 15936 4509 15969
rect 4569 15936 4647 15969
rect 4681 15950 4740 15970
rect 4774 15950 4809 15984
rect 4843 15950 4878 15984
rect 4912 15950 4947 15984
rect 4981 15950 5016 15984
rect 5050 15950 5085 15984
rect 5123 15967 5154 15984
rect 5196 15967 5223 15984
rect 5269 15967 5292 15984
rect 5342 15967 5361 15984
rect 5415 15967 5430 15984
rect 5488 15967 5499 15984
rect 5561 15967 5568 15984
rect 5634 15967 5637 15984
rect 5119 15950 5154 15967
rect 5188 15950 5223 15967
rect 5257 15950 5292 15967
rect 5326 15950 5361 15967
rect 5395 15950 5430 15967
rect 5464 15950 5499 15967
rect 5533 15950 5568 15967
rect 5602 15950 5637 15967
rect 5671 15967 5673 15984
rect 5740 15967 5746 15984
rect 5809 15967 5819 15984
rect 5878 15967 5892 15984
rect 5947 15967 5965 15984
rect 6016 15967 6038 15984
rect 6085 15967 6110 15984
rect 6154 15967 6182 15984
rect 6223 15967 6254 15984
rect 6292 15967 6326 15984
rect 5671 15950 5706 15967
rect 5740 15950 5775 15967
rect 5809 15950 5844 15967
rect 5878 15950 5913 15967
rect 5947 15950 5982 15967
rect 6016 15950 6051 15967
rect 6085 15950 6120 15967
rect 6154 15950 6189 15967
rect 6223 15950 6258 15967
rect 6292 15950 6327 15967
rect 6361 15950 6396 15984
rect 6432 15967 6465 15984
rect 6504 15967 6534 15984
rect 6576 15967 6603 15984
rect 6648 15967 6672 15984
rect 6720 15967 6741 15984
rect 6792 15967 6810 15984
rect 6864 15967 6879 15984
rect 6936 15967 6948 15984
rect 7008 15967 7017 15984
rect 7080 15967 7086 15984
rect 7152 15967 7155 15984
rect 6430 15950 6465 15967
rect 6499 15950 6534 15967
rect 6568 15950 6603 15967
rect 6637 15950 6672 15967
rect 6706 15950 6741 15967
rect 6775 15950 6810 15967
rect 6844 15950 6879 15967
rect 6913 15950 6948 15967
rect 6982 15950 7017 15967
rect 7051 15950 7086 15967
rect 7120 15950 7155 15967
rect 7189 15967 7190 15984
rect 7224 15984 7262 16001
rect 7296 15984 7334 16001
rect 7368 15984 7406 16001
rect 7440 15984 7478 16001
rect 7512 15984 7550 16001
rect 7584 15984 7622 16001
rect 7656 15984 7694 16001
rect 7728 15984 7766 16001
rect 7800 15984 7838 16001
rect 7872 15984 7908 16001
rect 7189 15950 7224 15967
rect 7258 15967 7262 15984
rect 7327 15967 7334 15984
rect 7396 15967 7406 15984
rect 7465 15967 7478 15984
rect 7534 15967 7550 15984
rect 7602 15967 7622 15984
rect 7670 15967 7694 15984
rect 7738 15967 7766 15984
rect 7806 15967 7838 15984
rect 7258 15950 7293 15967
rect 7327 15950 7362 15967
rect 7396 15950 7431 15967
rect 7465 15950 7500 15967
rect 7534 15950 7568 15967
rect 7602 15950 7636 15967
rect 7670 15950 7704 15967
rect 7738 15950 7772 15967
rect 7806 15950 7840 15967
rect 7874 15950 7908 15984
rect 4681 15936 7908 15950
rect 4497 15935 4535 15936
rect 4569 15935 7908 15936
rect 2704 15912 7908 15935
rect 3023 15552 3035 15586
rect 3073 15552 3108 15586
rect 3142 15552 3177 15586
rect 3215 15552 3246 15586
rect 3288 15552 3315 15586
rect 3361 15552 3384 15586
rect 3434 15552 3453 15586
rect 3507 15552 3522 15586
rect 3580 15552 3591 15586
rect 3653 15552 3660 15586
rect 3726 15552 3729 15586
rect 3763 15552 3765 15586
rect 3832 15552 3838 15586
rect 3901 15552 3911 15586
rect 3970 15552 3984 15586
rect 4039 15552 4057 15586
rect 4108 15552 4130 15586
rect 4177 15552 4203 15586
rect 4245 15552 4276 15586
rect 4313 15552 4347 15586
rect 4383 15552 4415 15586
rect 4456 15552 4483 15586
rect 4529 15552 4551 15586
rect 4602 15552 4619 15586
rect 4675 15552 4687 15586
rect 4748 15552 4755 15586
rect 4821 15552 4823 15586
rect 4857 15552 4860 15586
rect 4925 15552 4933 15586
rect 4993 15552 5006 15586
rect 5061 15552 5079 15586
rect 5129 15552 5152 15586
rect 5197 15552 5225 15586
rect 5265 15552 5298 15586
rect 5333 15552 5367 15586
rect 5405 15552 5435 15586
rect 5478 15552 5503 15586
rect 5551 15552 5571 15586
rect 5624 15552 5639 15586
rect 5697 15552 5707 15586
rect 5770 15552 5775 15586
rect 5877 15552 5881 15586
rect 5945 15552 5953 15586
rect 6013 15552 6025 15586
rect 6081 15552 6097 15586
rect 6149 15552 6169 15586
rect 6217 15552 6241 15586
rect 6285 15552 6313 15586
rect 6353 15552 6385 15586
rect 6421 15552 6455 15586
rect 6491 15552 6523 15586
rect 6563 15552 6591 15586
rect 6635 15552 6659 15586
rect 6707 15552 6727 15586
rect 6779 15552 6795 15586
rect 6851 15552 6863 15586
rect 6923 15552 6931 15586
rect 6995 15552 6999 15586
rect 7101 15552 7105 15586
rect 7169 15552 7177 15586
rect 7237 15552 7249 15586
rect 7305 15552 7321 15586
rect 7373 15552 7393 15586
rect 7441 15552 7465 15586
rect 7509 15552 7537 15586
rect 7577 15552 7609 15586
rect 7645 15552 7679 15586
rect 7715 15552 7729 15586
rect 3109 15446 3211 15458
rect 3663 15446 3765 15458
rect 4217 15446 4319 15458
rect 4771 15446 4873 15458
rect 5325 15446 5427 15458
rect 5879 15446 5981 15458
rect 6433 15446 6535 15458
rect 6987 15446 7089 15458
rect 7539 15446 7645 15458
rect 2864 15412 2902 15446
rect 2830 15373 2936 15412
rect 2864 15339 2902 15373
rect 2830 15300 2936 15339
rect 2864 15266 2902 15300
rect 2830 15227 2936 15266
rect 2864 15193 2902 15227
rect 2830 15154 2936 15193
rect 3141 15412 3179 15446
rect 3107 15373 3213 15412
rect 3141 15339 3179 15373
rect 3107 15300 3213 15339
rect 3141 15266 3179 15300
rect 3107 15227 3213 15266
rect 3141 15193 3179 15227
rect 3107 15154 3213 15193
rect 3418 15412 3456 15446
rect 3384 15373 3490 15412
rect 3418 15339 3456 15373
rect 3384 15300 3490 15339
rect 3418 15266 3456 15300
rect 3384 15227 3490 15266
rect 3418 15193 3456 15227
rect 3384 15154 3490 15193
rect 3695 15412 3733 15446
rect 3661 15373 3767 15412
rect 3695 15339 3733 15373
rect 3661 15300 3767 15339
rect 3695 15266 3733 15300
rect 3661 15227 3767 15266
rect 3695 15193 3733 15227
rect 3661 15154 3767 15193
rect 3972 15412 4010 15446
rect 3938 15373 4044 15412
rect 3972 15339 4010 15373
rect 3938 15300 4044 15339
rect 3972 15266 4010 15300
rect 3938 15227 4044 15266
rect 3972 15193 4010 15227
rect 3938 15154 4044 15193
rect 4249 15412 4287 15446
rect 4215 15373 4321 15412
rect 4249 15339 4287 15373
rect 4215 15300 4321 15339
rect 4249 15266 4287 15300
rect 4215 15227 4321 15266
rect 4249 15193 4287 15227
rect 4215 15154 4321 15193
rect 4526 15412 4564 15446
rect 4492 15373 4598 15412
rect 4526 15339 4564 15373
rect 4492 15300 4598 15339
rect 4526 15266 4564 15300
rect 4492 15227 4598 15266
rect 4526 15193 4564 15227
rect 4492 15154 4598 15193
rect 4803 15412 4841 15446
rect 4769 15373 4875 15412
rect 4803 15339 4841 15373
rect 4769 15300 4875 15339
rect 4803 15266 4841 15300
rect 4769 15227 4875 15266
rect 4803 15193 4841 15227
rect 4769 15154 4875 15193
rect 5080 15412 5118 15446
rect 5046 15373 5152 15412
rect 5080 15339 5118 15373
rect 5046 15300 5152 15339
rect 5080 15266 5118 15300
rect 5046 15227 5152 15266
rect 5080 15193 5118 15227
rect 5046 15154 5152 15193
rect 5357 15412 5395 15446
rect 5323 15373 5429 15412
rect 5357 15339 5395 15373
rect 5323 15300 5429 15339
rect 5357 15266 5395 15300
rect 5323 15227 5429 15266
rect 5357 15193 5395 15227
rect 5323 15154 5429 15193
rect 5634 15412 5672 15446
rect 5600 15373 5706 15412
rect 5634 15339 5672 15373
rect 5600 15300 5706 15339
rect 5634 15266 5672 15300
rect 5600 15227 5706 15266
rect 5634 15193 5672 15227
rect 5600 15154 5706 15193
rect 5911 15412 5949 15446
rect 5877 15373 5983 15412
rect 5911 15339 5949 15373
rect 5877 15300 5983 15339
rect 5911 15266 5949 15300
rect 5877 15227 5983 15266
rect 5911 15193 5949 15227
rect 5877 15154 5983 15193
rect 6188 15412 6226 15446
rect 6154 15373 6260 15412
rect 6188 15339 6226 15373
rect 6154 15300 6260 15339
rect 6188 15266 6226 15300
rect 6154 15227 6260 15266
rect 6188 15193 6226 15227
rect 6154 15154 6260 15193
rect 6465 15412 6503 15446
rect 6431 15373 6537 15412
rect 6465 15339 6503 15373
rect 6431 15300 6537 15339
rect 6465 15266 6503 15300
rect 6431 15227 6537 15266
rect 6465 15193 6503 15227
rect 6431 15154 6537 15193
rect 6742 15412 6780 15446
rect 6708 15373 6814 15412
rect 6742 15339 6780 15373
rect 6708 15300 6814 15339
rect 6742 15266 6780 15300
rect 6708 15227 6814 15266
rect 6742 15193 6780 15227
rect 6708 15154 6814 15193
rect 7019 15412 7057 15446
rect 6985 15373 7091 15412
rect 7019 15339 7057 15373
rect 6985 15300 7091 15339
rect 7019 15266 7057 15300
rect 6985 15227 7091 15266
rect 7019 15193 7057 15227
rect 6985 15154 7091 15193
rect 7296 15412 7334 15446
rect 7262 15373 7368 15412
rect 7296 15339 7334 15373
rect 7262 15300 7368 15339
rect 7296 15266 7334 15300
rect 7262 15227 7368 15266
rect 7296 15193 7334 15227
rect 7262 15154 7368 15193
rect 7573 15412 7611 15446
rect 7539 15373 7645 15412
rect 7573 15339 7611 15373
rect 7539 15300 7645 15339
rect 7573 15266 7611 15300
rect 7539 15227 7645 15266
rect 7573 15193 7611 15227
rect 7539 15154 7645 15193
rect 7850 15412 7888 15446
rect 7816 15373 7922 15412
rect 7850 15339 7888 15373
rect 7816 15300 7922 15339
rect 7850 15266 7888 15300
rect 7816 15227 7922 15266
rect 7850 15193 7888 15227
rect 7816 15154 7922 15193
rect 3109 14100 3211 14112
rect 3663 14100 3765 14112
rect 4217 14100 4319 14112
rect 4771 14100 4873 14112
rect 5325 14100 5427 14112
rect 5879 14100 5981 14112
rect 6433 14100 6535 14112
rect 6987 14100 7089 14112
rect 7539 14100 7645 14112
rect 3023 13822 3035 13856
rect 3073 13822 3108 13856
rect 3142 13822 3177 13856
rect 3215 13822 3246 13856
rect 3288 13822 3315 13856
rect 3361 13822 3384 13856
rect 3434 13822 3453 13856
rect 3507 13822 3522 13856
rect 3580 13822 3591 13856
rect 3653 13822 3660 13856
rect 3726 13822 3729 13856
rect 3763 13822 3765 13856
rect 3832 13822 3838 13856
rect 3901 13822 3911 13856
rect 3970 13822 3984 13856
rect 4039 13822 4057 13856
rect 4107 13822 4130 13856
rect 4175 13822 4203 13856
rect 4243 13822 4276 13856
rect 4311 13822 4345 13856
rect 4383 13822 4413 13856
rect 4456 13822 4481 13856
rect 4529 13822 4549 13856
rect 4602 13822 4617 13856
rect 4675 13822 4685 13856
rect 4748 13822 4753 13856
rect 4855 13822 4860 13856
rect 4923 13822 4933 13856
rect 4991 13822 5006 13856
rect 5059 13822 5079 13856
rect 5127 13822 5152 13856
rect 5195 13822 5225 13856
rect 5263 13822 5297 13856
rect 5332 13822 5365 13856
rect 5405 13822 5433 13856
rect 5478 13822 5501 13856
rect 5551 13822 5569 13856
rect 5624 13822 5637 13856
rect 5697 13822 5705 13856
rect 5770 13822 5773 13856
rect 5807 13822 5809 13856
rect 5875 13822 5881 13856
rect 5943 13822 5953 13856
rect 6011 13822 6025 13856
rect 6079 13822 6097 13856
rect 6147 13822 6169 13856
rect 6215 13822 6241 13856
rect 6283 13822 6313 13856
rect 6351 13822 6385 13856
rect 6419 13822 6453 13856
rect 6491 13822 6521 13856
rect 6563 13822 6589 13856
rect 6635 13822 6657 13856
rect 6707 13822 6725 13856
rect 6779 13822 6793 13856
rect 6851 13822 6861 13856
rect 6923 13822 6929 13856
rect 6995 13822 6997 13856
rect 7031 13822 7033 13856
rect 7099 13822 7105 13856
rect 7167 13822 7177 13856
rect 7235 13822 7249 13856
rect 7303 13822 7321 13856
rect 7371 13822 7393 13856
rect 7439 13822 7465 13856
rect 7507 13822 7537 13856
rect 7575 13822 7609 13856
rect 7643 13822 7677 13856
rect 7715 13822 7727 13856
rect 3109 13446 3211 13458
rect 3663 13446 3765 13458
rect 4217 13446 4319 13458
rect 4771 13446 4873 13458
rect 5325 13446 5427 13458
rect 5879 13446 5981 13458
rect 6433 13446 6535 13458
rect 6987 13446 7089 13458
rect 7539 13446 7645 13458
rect 2864 13412 2902 13446
rect 2830 13373 2936 13412
rect 2864 13339 2902 13373
rect 2830 13300 2936 13339
rect 2864 13266 2902 13300
rect 2830 13227 2936 13266
rect 2864 13193 2902 13227
rect 2830 13154 2936 13193
rect 3141 13412 3179 13446
rect 3107 13373 3213 13412
rect 3141 13339 3179 13373
rect 3107 13300 3213 13339
rect 3141 13266 3179 13300
rect 3107 13227 3213 13266
rect 3141 13193 3179 13227
rect 3107 13154 3213 13193
rect 3418 13412 3456 13446
rect 3384 13373 3490 13412
rect 3418 13339 3456 13373
rect 3384 13300 3490 13339
rect 3418 13266 3456 13300
rect 3384 13227 3490 13266
rect 3418 13193 3456 13227
rect 3384 13154 3490 13193
rect 3695 13412 3733 13446
rect 3661 13373 3767 13412
rect 3695 13339 3733 13373
rect 3661 13300 3767 13339
rect 3695 13266 3733 13300
rect 3661 13227 3767 13266
rect 3695 13193 3733 13227
rect 3661 13154 3767 13193
rect 3972 13412 4010 13446
rect 3938 13373 4044 13412
rect 3972 13339 4010 13373
rect 3938 13300 4044 13339
rect 3972 13266 4010 13300
rect 3938 13227 4044 13266
rect 3972 13193 4010 13227
rect 3938 13154 4044 13193
rect 4249 13412 4287 13446
rect 4215 13373 4321 13412
rect 4249 13339 4287 13373
rect 4215 13300 4321 13339
rect 4249 13266 4287 13300
rect 4215 13227 4321 13266
rect 4249 13193 4287 13227
rect 4215 13154 4321 13193
rect 4526 13412 4564 13446
rect 4492 13373 4598 13412
rect 4526 13339 4564 13373
rect 4492 13300 4598 13339
rect 4526 13266 4564 13300
rect 4492 13227 4598 13266
rect 4526 13193 4564 13227
rect 4492 13154 4598 13193
rect 4803 13412 4841 13446
rect 4769 13373 4875 13412
rect 4803 13339 4841 13373
rect 4769 13300 4875 13339
rect 4803 13266 4841 13300
rect 4769 13227 4875 13266
rect 4803 13193 4841 13227
rect 4769 13154 4875 13193
rect 5080 13412 5118 13446
rect 5046 13373 5152 13412
rect 5080 13339 5118 13373
rect 5046 13300 5152 13339
rect 5080 13266 5118 13300
rect 5046 13227 5152 13266
rect 5080 13193 5118 13227
rect 5046 13154 5152 13193
rect 5357 13412 5395 13446
rect 5323 13373 5429 13412
rect 5357 13339 5395 13373
rect 5323 13300 5429 13339
rect 5357 13266 5395 13300
rect 5323 13227 5429 13266
rect 5357 13193 5395 13227
rect 5323 13154 5429 13193
rect 5634 13412 5672 13446
rect 5600 13373 5706 13412
rect 5634 13339 5672 13373
rect 5600 13300 5706 13339
rect 5634 13266 5672 13300
rect 5600 13227 5706 13266
rect 5634 13193 5672 13227
rect 5600 13154 5706 13193
rect 5911 13412 5949 13446
rect 5877 13373 5983 13412
rect 5911 13339 5949 13373
rect 5877 13300 5983 13339
rect 5911 13266 5949 13300
rect 5877 13227 5983 13266
rect 5911 13193 5949 13227
rect 5877 13154 5983 13193
rect 6188 13412 6226 13446
rect 6154 13373 6260 13412
rect 6188 13339 6226 13373
rect 6154 13300 6260 13339
rect 6188 13266 6226 13300
rect 6154 13227 6260 13266
rect 6188 13193 6226 13227
rect 6154 13154 6260 13193
rect 6465 13412 6503 13446
rect 6431 13373 6537 13412
rect 6465 13339 6503 13373
rect 6431 13300 6537 13339
rect 6465 13266 6503 13300
rect 6431 13227 6537 13266
rect 6465 13193 6503 13227
rect 6431 13154 6537 13193
rect 6742 13412 6780 13446
rect 6708 13373 6814 13412
rect 6742 13339 6780 13373
rect 6708 13300 6814 13339
rect 6742 13266 6780 13300
rect 6708 13227 6814 13266
rect 6742 13193 6780 13227
rect 6708 13154 6814 13193
rect 7019 13412 7057 13446
rect 6985 13373 7091 13412
rect 7019 13339 7057 13373
rect 6985 13300 7091 13339
rect 7019 13266 7057 13300
rect 6985 13227 7091 13266
rect 7019 13193 7057 13227
rect 6985 13154 7091 13193
rect 7296 13412 7334 13446
rect 7262 13373 7368 13412
rect 7296 13339 7334 13373
rect 7262 13300 7368 13339
rect 7296 13266 7334 13300
rect 7262 13227 7368 13266
rect 7296 13193 7334 13227
rect 7262 13154 7368 13193
rect 7573 13412 7611 13446
rect 7539 13373 7645 13412
rect 7573 13339 7611 13373
rect 7539 13300 7645 13339
rect 7573 13266 7611 13300
rect 7539 13227 7645 13266
rect 7573 13193 7611 13227
rect 7539 13154 7645 13193
rect 7850 13412 7888 13446
rect 7816 13373 7922 13412
rect 7850 13339 7888 13373
rect 7816 13300 7922 13339
rect 7850 13266 7888 13300
rect 7816 13227 7922 13266
rect 7850 13193 7888 13227
rect 7816 13154 7922 13193
rect 3109 12100 3211 12112
rect 3663 12100 3765 12112
rect 4217 12100 4319 12112
rect 4771 12100 4873 12112
rect 5325 12100 5427 12112
rect 5879 12100 5981 12112
rect 6433 12100 6535 12112
rect 6987 12100 7089 12112
rect 7539 12100 7645 12112
rect 3023 11784 3035 11818
rect 3073 11784 3108 11818
rect 3142 11784 3177 11818
rect 3215 11784 3246 11818
rect 3288 11784 3315 11818
rect 3361 11784 3384 11818
rect 3434 11784 3453 11818
rect 3507 11784 3522 11818
rect 3580 11784 3591 11818
rect 3653 11784 3660 11818
rect 3726 11784 3729 11818
rect 3763 11784 3765 11818
rect 3832 11784 3838 11818
rect 3901 11784 3911 11818
rect 3970 11784 3984 11818
rect 4039 11784 4057 11818
rect 4107 11784 4130 11818
rect 4175 11784 4203 11818
rect 4243 11784 4276 11818
rect 4311 11784 4345 11818
rect 4383 11784 4413 11818
rect 4456 11784 4481 11818
rect 4529 11784 4549 11818
rect 4602 11784 4617 11818
rect 4675 11784 4685 11818
rect 4748 11784 4753 11818
rect 4855 11784 4860 11818
rect 4923 11784 4933 11818
rect 4991 11784 5006 11818
rect 5059 11784 5079 11818
rect 5127 11784 5152 11818
rect 5195 11784 5225 11818
rect 5263 11784 5297 11818
rect 5332 11784 5365 11818
rect 5405 11784 5433 11818
rect 5478 11784 5501 11818
rect 5551 11784 5569 11818
rect 5624 11784 5637 11818
rect 5697 11784 5705 11818
rect 5770 11784 5773 11818
rect 5807 11784 5809 11818
rect 5875 11784 5881 11818
rect 5943 11784 5953 11818
rect 6011 11784 6025 11818
rect 6079 11784 6097 11818
rect 6147 11784 6169 11818
rect 6215 11784 6241 11818
rect 6283 11784 6313 11818
rect 6351 11784 6385 11818
rect 6419 11784 6453 11818
rect 6491 11784 6521 11818
rect 6563 11784 6589 11818
rect 6635 11784 6657 11818
rect 6707 11784 6725 11818
rect 6779 11784 6793 11818
rect 6851 11784 6861 11818
rect 6923 11784 6929 11818
rect 6995 11784 6997 11818
rect 7031 11784 7033 11818
rect 7099 11784 7105 11818
rect 7167 11784 7177 11818
rect 7235 11784 7249 11818
rect 7303 11784 7321 11818
rect 7371 11784 7393 11818
rect 7439 11784 7465 11818
rect 7507 11784 7537 11818
rect 7575 11784 7609 11818
rect 7643 11784 7677 11818
rect 7715 11784 7727 11818
rect 3109 11446 3211 11458
rect 3663 11446 3765 11458
rect 4217 11446 4319 11458
rect 4771 11446 4873 11458
rect 5325 11446 5427 11458
rect 5879 11446 5981 11458
rect 6433 11446 6535 11458
rect 6987 11446 7089 11458
rect 7539 11446 7645 11458
rect 2864 11412 2902 11446
rect 2830 11373 2936 11412
rect 2864 11339 2902 11373
rect 2830 11300 2936 11339
rect 2864 11266 2902 11300
rect 2830 11227 2936 11266
rect 2864 11193 2902 11227
rect 2830 11154 2936 11193
rect 3141 11412 3179 11446
rect 3107 11373 3213 11412
rect 3141 11339 3179 11373
rect 3107 11300 3213 11339
rect 3141 11266 3179 11300
rect 3107 11227 3213 11266
rect 3141 11193 3179 11227
rect 3107 11154 3213 11193
rect 3418 11412 3456 11446
rect 3384 11373 3490 11412
rect 3418 11339 3456 11373
rect 3384 11300 3490 11339
rect 3418 11266 3456 11300
rect 3384 11227 3490 11266
rect 3418 11193 3456 11227
rect 3384 11154 3490 11193
rect 3695 11412 3733 11446
rect 3661 11373 3767 11412
rect 3695 11339 3733 11373
rect 3661 11300 3767 11339
rect 3695 11266 3733 11300
rect 3661 11227 3767 11266
rect 3695 11193 3733 11227
rect 3661 11154 3767 11193
rect 3972 11412 4010 11446
rect 3938 11373 4044 11412
rect 3972 11339 4010 11373
rect 3938 11300 4044 11339
rect 3972 11266 4010 11300
rect 3938 11227 4044 11266
rect 3972 11193 4010 11227
rect 3938 11154 4044 11193
rect 4249 11412 4287 11446
rect 4215 11373 4321 11412
rect 4249 11339 4287 11373
rect 4215 11300 4321 11339
rect 4249 11266 4287 11300
rect 4215 11227 4321 11266
rect 4249 11193 4287 11227
rect 4215 11154 4321 11193
rect 4526 11412 4564 11446
rect 4492 11373 4598 11412
rect 4526 11339 4564 11373
rect 4492 11300 4598 11339
rect 4526 11266 4564 11300
rect 4492 11227 4598 11266
rect 4526 11193 4564 11227
rect 4492 11154 4598 11193
rect 4803 11412 4841 11446
rect 4769 11373 4875 11412
rect 4803 11339 4841 11373
rect 4769 11300 4875 11339
rect 4803 11266 4841 11300
rect 4769 11227 4875 11266
rect 4803 11193 4841 11227
rect 4769 11154 4875 11193
rect 5080 11412 5118 11446
rect 5046 11373 5152 11412
rect 5080 11339 5118 11373
rect 5046 11300 5152 11339
rect 5080 11266 5118 11300
rect 5046 11227 5152 11266
rect 5080 11193 5118 11227
rect 5046 11154 5152 11193
rect 5357 11412 5395 11446
rect 5323 11373 5429 11412
rect 5357 11339 5395 11373
rect 5323 11300 5429 11339
rect 5357 11266 5395 11300
rect 5323 11227 5429 11266
rect 5357 11193 5395 11227
rect 5323 11154 5429 11193
rect 5634 11412 5672 11446
rect 5600 11373 5706 11412
rect 5634 11339 5672 11373
rect 5600 11300 5706 11339
rect 5634 11266 5672 11300
rect 5600 11227 5706 11266
rect 5634 11193 5672 11227
rect 5600 11154 5706 11193
rect 5911 11412 5949 11446
rect 5877 11373 5983 11412
rect 5911 11339 5949 11373
rect 5877 11300 5983 11339
rect 5911 11266 5949 11300
rect 5877 11227 5983 11266
rect 5911 11193 5949 11227
rect 5877 11154 5983 11193
rect 6188 11412 6226 11446
rect 6154 11373 6260 11412
rect 6188 11339 6226 11373
rect 6154 11300 6260 11339
rect 6188 11266 6226 11300
rect 6154 11227 6260 11266
rect 6188 11193 6226 11227
rect 6154 11154 6260 11193
rect 6465 11412 6503 11446
rect 6431 11373 6537 11412
rect 6465 11339 6503 11373
rect 6431 11300 6537 11339
rect 6465 11266 6503 11300
rect 6431 11227 6537 11266
rect 6465 11193 6503 11227
rect 6431 11154 6537 11193
rect 6742 11412 6780 11446
rect 6708 11373 6814 11412
rect 6742 11339 6780 11373
rect 6708 11300 6814 11339
rect 6742 11266 6780 11300
rect 6708 11227 6814 11266
rect 6742 11193 6780 11227
rect 6708 11154 6814 11193
rect 7019 11412 7057 11446
rect 6985 11373 7091 11412
rect 7019 11339 7057 11373
rect 6985 11300 7091 11339
rect 7019 11266 7057 11300
rect 6985 11227 7091 11266
rect 7019 11193 7057 11227
rect 6985 11154 7091 11193
rect 7296 11412 7334 11446
rect 7262 11373 7368 11412
rect 7296 11339 7334 11373
rect 7262 11300 7368 11339
rect 7296 11266 7334 11300
rect 7262 11227 7368 11266
rect 7296 11193 7334 11227
rect 7262 11154 7368 11193
rect 7573 11412 7611 11446
rect 7539 11373 7645 11412
rect 7573 11339 7611 11373
rect 7539 11300 7645 11339
rect 7573 11266 7611 11300
rect 7539 11227 7645 11266
rect 7573 11193 7611 11227
rect 7539 11154 7645 11193
rect 7850 11412 7888 11446
rect 7816 11373 7922 11412
rect 7850 11339 7888 11373
rect 7816 11300 7922 11339
rect 7850 11266 7888 11300
rect 7816 11227 7922 11266
rect 7850 11193 7888 11227
rect 7816 11154 7922 11193
rect 3109 10100 3211 10112
rect 3663 10100 3765 10112
rect 4217 10100 4319 10112
rect 4771 10100 4873 10112
rect 5325 10100 5427 10112
rect 5879 10100 5981 10112
rect 6433 10100 6535 10112
rect 6987 10100 7089 10112
rect 7539 10100 7645 10112
rect 3023 10050 3039 10056
rect 3023 10022 3035 10050
rect 3073 10022 3108 10056
rect 3142 10022 3177 10056
rect 3211 10050 3246 10056
rect 3280 10050 3315 10056
rect 3349 10050 3384 10056
rect 3418 10050 3453 10056
rect 3487 10050 3522 10056
rect 3556 10050 3591 10056
rect 3625 10050 3660 10056
rect 3694 10050 3729 10056
rect 3215 10022 3246 10050
rect 3288 10022 3315 10050
rect 3361 10022 3384 10050
rect 3434 10022 3453 10050
rect 3507 10022 3522 10050
rect 3580 10022 3591 10050
rect 3653 10022 3660 10050
rect 3726 10022 3729 10050
rect 3763 10050 3798 10056
rect 3832 10050 3867 10056
rect 3901 10050 3936 10056
rect 3970 10050 4005 10056
rect 4039 10050 4074 10056
rect 4108 10050 4143 10056
rect 4177 10050 4211 10056
rect 4245 10050 4279 10056
rect 3763 10022 3765 10050
rect 3832 10022 3838 10050
rect 3901 10022 3911 10050
rect 3970 10022 3984 10050
rect 4039 10022 4057 10050
rect 4108 10022 4130 10050
rect 4177 10022 4203 10050
rect 4245 10022 4276 10050
rect 4313 10022 4347 10056
rect 4381 10050 4415 10056
rect 4449 10050 4483 10056
rect 4517 10050 4551 10056
rect 4585 10050 4619 10056
rect 4653 10050 4687 10056
rect 4721 10050 4755 10056
rect 4789 10050 4823 10056
rect 4383 10022 4415 10050
rect 4456 10022 4483 10050
rect 4529 10022 4551 10050
rect 4602 10022 4619 10050
rect 4675 10022 4687 10050
rect 4748 10022 4755 10050
rect 4821 10022 4823 10050
rect 4857 10050 4891 10056
rect 4925 10050 4959 10056
rect 4993 10050 5027 10056
rect 5061 10050 5095 10056
rect 5129 10050 5163 10056
rect 5197 10050 5231 10056
rect 5265 10050 5299 10056
rect 4857 10022 4860 10050
rect 4925 10022 4933 10050
rect 4993 10022 5006 10050
rect 5061 10022 5079 10050
rect 5129 10022 5152 10050
rect 5197 10022 5225 10050
rect 5265 10022 5298 10050
rect 5333 10022 5367 10056
rect 5401 10050 5435 10056
rect 5469 10050 5503 10056
rect 5537 10050 5571 10056
rect 5605 10050 5639 10056
rect 5673 10050 5707 10056
rect 5741 10050 5775 10056
rect 5405 10022 5435 10050
rect 5478 10022 5503 10050
rect 5551 10022 5571 10050
rect 5624 10022 5639 10050
rect 5697 10022 5707 10050
rect 5770 10022 5775 10050
rect 5809 10050 5843 10056
rect 3069 10016 3108 10022
rect 3142 10016 3181 10022
rect 3215 10016 3254 10022
rect 3288 10016 3327 10022
rect 3361 10016 3400 10022
rect 3434 10016 3473 10022
rect 3507 10016 3546 10022
rect 3580 10016 3619 10022
rect 3653 10016 3692 10022
rect 3726 10016 3765 10022
rect 3799 10016 3838 10022
rect 3872 10016 3911 10022
rect 3945 10016 3984 10022
rect 4018 10016 4057 10022
rect 4091 10016 4130 10022
rect 4164 10016 4203 10022
rect 4237 10016 4276 10022
rect 4310 10016 4349 10022
rect 4383 10016 4422 10022
rect 4456 10016 4495 10022
rect 4529 10016 4568 10022
rect 4602 10016 4641 10022
rect 4675 10016 4714 10022
rect 4748 10016 4787 10022
rect 4821 10016 4860 10022
rect 4894 10016 4933 10022
rect 4967 10016 5006 10022
rect 5040 10016 5079 10022
rect 5113 10016 5152 10022
rect 5186 10016 5225 10022
rect 5259 10016 5298 10022
rect 5332 10016 5371 10022
rect 5405 10016 5444 10022
rect 5478 10016 5517 10022
rect 5551 10016 5590 10022
rect 5624 10016 5663 10022
rect 5697 10016 5736 10022
rect 5770 10016 5809 10022
rect 5877 10050 5911 10056
rect 5945 10050 5979 10056
rect 6013 10050 6047 10056
rect 6081 10050 6115 10056
rect 6149 10050 6183 10056
rect 6217 10050 6251 10056
rect 6285 10050 6319 10056
rect 5877 10022 5882 10050
rect 5945 10022 5955 10050
rect 6013 10022 6027 10050
rect 6081 10022 6099 10050
rect 6149 10022 6171 10050
rect 6217 10022 6243 10050
rect 6285 10022 6315 10050
rect 6353 10022 6387 10056
rect 6421 10022 6455 10056
rect 6489 10050 6523 10056
rect 6557 10050 6591 10056
rect 6625 10050 6659 10056
rect 6693 10050 6727 10056
rect 6761 10050 6795 10056
rect 6829 10050 6863 10056
rect 6897 10050 6931 10056
rect 6965 10050 6999 10056
rect 6493 10022 6523 10050
rect 6565 10022 6591 10050
rect 6637 10022 6659 10050
rect 6709 10022 6727 10050
rect 6781 10022 6795 10050
rect 6853 10022 6863 10050
rect 6925 10022 6931 10050
rect 6997 10022 6999 10050
rect 7033 10050 7067 10056
rect 7101 10050 7135 10056
rect 7169 10050 7203 10056
rect 7237 10050 7271 10056
rect 7305 10050 7339 10056
rect 7373 10050 7407 10056
rect 7441 10050 7475 10056
rect 7509 10050 7543 10056
rect 7033 10022 7035 10050
rect 7101 10022 7107 10050
rect 7169 10022 7179 10050
rect 7237 10022 7251 10050
rect 7305 10022 7323 10050
rect 7373 10022 7395 10050
rect 7441 10022 7467 10050
rect 7509 10022 7539 10050
rect 7577 10022 7611 10056
rect 7645 10022 7679 10056
rect 7713 10050 7729 10056
rect 7717 10022 7729 10050
rect 5843 10016 5882 10022
rect 5916 10016 5955 10022
rect 5989 10016 6027 10022
rect 6061 10016 6099 10022
rect 6133 10016 6171 10022
rect 6205 10016 6243 10022
rect 6277 10016 6315 10022
rect 6349 10016 6387 10022
rect 6421 10016 6459 10022
rect 6493 10016 6531 10022
rect 6565 10016 6603 10022
rect 6637 10016 6675 10022
rect 6709 10016 6747 10022
rect 6781 10016 6819 10022
rect 6853 10016 6891 10022
rect 6925 10016 6963 10022
rect 6997 10016 7035 10022
rect 7069 10016 7107 10022
rect 7141 10016 7179 10022
rect 7213 10016 7251 10022
rect 7285 10016 7323 10022
rect 7357 10016 7395 10022
rect 7429 10016 7467 10022
rect 7501 10016 7539 10022
rect 7573 10016 7611 10022
rect 7645 10016 7683 10022
rect 2274 9986 2276 10004
rect 2310 9986 2410 10004
rect 2274 9948 2444 9986
rect 2274 9914 2276 9948
rect 2310 9919 2410 9948
rect 8195 9949 8219 9953
rect 2274 9885 2298 9914
rect 2332 9885 2367 9919
rect 2401 9914 2410 9919
rect 2401 9885 2436 9914
rect 2470 9885 2505 9919
rect 2539 9885 2574 9919
rect 2608 9885 2643 9919
rect 2677 9885 2712 9919
rect 2746 9885 2781 9919
rect 2815 9885 2850 9919
rect 2884 9885 2919 9919
rect 2953 9885 2988 9919
rect 3022 9885 3057 9919
rect 3091 9885 3126 9919
rect 3160 9885 3195 9919
rect 3229 9885 3264 9919
rect 3298 9885 3333 9919
rect 3367 9885 3401 9919
rect 3435 9885 3469 9919
rect 3503 9885 3537 9919
rect 3571 9885 3605 9919
rect 3639 9885 3673 9919
rect 3707 9885 3741 9919
rect 3775 9885 3809 9919
rect 3843 9885 3877 9919
rect 3911 9885 3945 9919
rect 3979 9885 4013 9919
rect 4047 9885 4081 9919
rect 4115 9885 4149 9919
rect 4183 9885 4217 9919
rect 4251 9885 4285 9919
rect 4319 9885 4353 9919
rect 4387 9885 4421 9919
rect 4455 9885 4489 9919
rect 4523 9885 4557 9919
rect 4591 9885 4625 9919
rect 4659 9885 4693 9919
rect 4727 9885 4761 9919
rect 4795 9885 4829 9919
rect 4863 9885 4897 9919
rect 4931 9885 4965 9919
rect 4999 9885 5033 9919
rect 5067 9885 5101 9919
rect 5135 9885 5169 9919
rect 5203 9885 5237 9919
rect 5271 9885 5305 9919
rect 5339 9885 5373 9919
rect 5407 9885 5441 9919
rect 5475 9885 5509 9919
rect 5543 9885 5577 9919
rect 5611 9885 5645 9919
rect 5679 9885 5713 9919
rect 5747 9885 5781 9919
rect 5815 9885 5849 9919
rect 5883 9885 5917 9919
rect 5951 9885 5985 9919
rect 6019 9885 6053 9919
rect 6087 9885 6121 9919
rect 6155 9885 6189 9919
rect 6223 9885 6257 9919
rect 6291 9885 6325 9919
rect 6359 9885 6393 9919
rect 6427 9885 6461 9919
rect 6495 9885 6529 9919
rect 6563 9885 6597 9919
rect 6631 9885 6665 9919
rect 6699 9885 6733 9919
rect 6767 9885 6801 9919
rect 6835 9885 6869 9919
rect 6903 9885 6937 9919
rect 6971 9885 7005 9919
rect 7039 9885 7073 9919
rect 7107 9885 7141 9919
rect 7175 9885 7209 9919
rect 7243 9885 7277 9919
rect 7311 9885 7345 9919
rect 7379 9885 7413 9919
rect 7447 9885 7481 9919
rect 7515 9885 7549 9919
rect 7583 9885 7617 9919
rect 7651 9885 7685 9919
rect 7719 9885 7753 9919
rect 7787 9885 7821 9919
rect 7855 9885 7889 9919
rect 7923 9885 7957 9919
rect 7991 9885 8025 9919
rect 8218 9915 8219 9949
rect 8195 9885 8219 9915
rect 2274 9876 8219 9885
rect 2274 9842 2276 9876
rect 2310 9842 2410 9876
rect 2444 9870 8050 9876
rect 2444 9842 2482 9870
rect 2274 9836 2482 9842
rect 2516 9836 2555 9870
rect 2589 9836 2628 9870
rect 2662 9836 2701 9870
rect 2735 9836 2774 9870
rect 2808 9836 2847 9870
rect 2881 9836 2920 9870
rect 2954 9836 2993 9870
rect 3027 9836 3066 9870
rect 3100 9836 3139 9870
rect 3173 9836 3212 9870
rect 3246 9836 3285 9870
rect 3319 9836 3358 9870
rect 3392 9836 3431 9870
rect 3465 9836 3504 9870
rect 3538 9836 3577 9870
rect 3611 9836 3650 9870
rect 3684 9836 3723 9870
rect 3757 9836 3796 9870
rect 3830 9836 3869 9870
rect 3903 9836 3942 9870
rect 3976 9836 4015 9870
rect 4049 9836 4088 9870
rect 4122 9836 4161 9870
rect 4195 9836 4234 9870
rect 4268 9836 4306 9870
rect 4340 9836 4378 9870
rect 4412 9836 4450 9870
rect 4484 9836 4522 9870
rect 4556 9836 4594 9870
rect 4628 9836 4666 9870
rect 4700 9836 4738 9870
rect 4772 9836 4810 9870
rect 4844 9836 4882 9870
rect 4916 9836 4954 9870
rect 4988 9836 5026 9870
rect 5060 9836 5098 9870
rect 5132 9836 5170 9870
rect 5204 9836 5242 9870
rect 5276 9836 5314 9870
rect 5348 9836 5386 9870
rect 5420 9836 5458 9870
rect 5492 9836 5530 9870
rect 5564 9836 5602 9870
rect 5636 9836 5674 9870
rect 5708 9836 5746 9870
rect 5780 9836 5818 9870
rect 5852 9836 5890 9870
rect 5924 9836 5962 9870
rect 5996 9836 6034 9870
rect 6068 9836 6106 9870
rect 6140 9836 6178 9870
rect 6212 9836 6250 9870
rect 6284 9836 6322 9870
rect 6356 9836 6394 9870
rect 6428 9836 6466 9870
rect 6500 9836 6538 9870
rect 6572 9836 6610 9870
rect 6644 9836 6682 9870
rect 6716 9836 6754 9870
rect 6788 9836 6826 9870
rect 6860 9836 6898 9870
rect 6932 9836 6970 9870
rect 7004 9836 7042 9870
rect 7076 9836 7114 9870
rect 7148 9836 7186 9870
rect 7220 9836 7258 9870
rect 7292 9836 7330 9870
rect 7364 9836 7402 9870
rect 7436 9836 7474 9870
rect 7508 9836 7546 9870
rect 7580 9836 7618 9870
rect 7652 9836 7690 9870
rect 7724 9836 7762 9870
rect 7796 9836 7834 9870
rect 7868 9836 7906 9870
rect 7940 9836 7978 9870
rect 8012 9842 8050 9870
rect 8084 9842 8184 9876
rect 8218 9842 8219 9876
rect 8012 9836 8219 9842
rect 2274 9830 8219 9836
rect 8429 14491 8431 14530
rect 8533 14491 8535 14530
rect 8429 14418 8431 14457
rect 8533 14418 8535 14457
rect 8429 14345 8431 14384
rect 8533 14345 8535 14384
rect 8429 14272 8431 14311
rect 8533 14272 8535 14311
rect 8429 14199 8431 14238
rect 8533 14199 8535 14238
rect 8429 14126 8431 14165
rect 8533 14126 8535 14165
rect 8429 14053 8431 14092
rect 8533 14053 8535 14092
rect 8429 13980 8431 14019
rect 8533 13980 8535 14019
rect 8429 13907 8431 13946
rect 8533 13907 8535 13946
rect 8429 13834 8431 13873
rect 8533 13834 8535 13873
rect 8429 13761 8431 13800
rect 8533 13761 8535 13800
rect 8429 13688 8431 13727
rect 8533 13688 8535 13727
rect 8429 13615 8431 13654
rect 8533 13615 8535 13654
rect 8429 13542 8431 13581
rect 8533 13542 8535 13581
rect 8429 13469 8431 13508
rect 8533 13469 8535 13508
rect 8429 13396 8431 13435
rect 8533 13396 8535 13435
rect 8429 13323 8431 13362
rect 8533 13323 8535 13362
rect 8429 13250 8431 13289
rect 8533 13250 8535 13289
rect 8429 13177 8431 13216
rect 8533 13177 8535 13216
rect 8429 13104 8431 13143
rect 8533 13104 8535 13143
rect 8429 13031 8431 13070
rect 8533 13031 8535 13070
rect 8429 12958 8431 12997
rect 8533 12958 8535 12997
rect 8429 12885 8431 12924
rect 8533 12885 8535 12924
rect 8429 12812 8431 12851
rect 8533 12812 8535 12851
rect 8429 12739 8431 12778
rect 8533 12739 8535 12778
rect 8429 12666 8431 12705
rect 8533 12666 8535 12705
rect 8429 12593 8431 12632
rect 8533 12593 8535 12632
rect 8429 12520 8431 12559
rect 8533 12520 8535 12559
rect 8429 12447 8431 12486
rect 8533 12447 8535 12486
rect 8429 12374 8431 12413
rect 8533 12374 8535 12413
rect 8429 12301 8431 12340
rect 8533 12301 8535 12340
rect 8429 12228 8431 12267
rect 8533 12228 8535 12267
rect 8429 12155 8431 12194
rect 8533 12155 8535 12194
rect 8429 12082 8431 12121
rect 8533 12082 8535 12121
rect 8429 12009 8431 12048
rect 8533 12009 8535 12048
rect 8429 11936 8431 11975
rect 8533 11936 8535 11975
rect 8429 11863 8431 11902
rect 8533 11863 8535 11902
rect 8429 11790 8431 11829
rect 8533 11790 8535 11829
rect 8429 11717 8431 11756
rect 8533 11717 8535 11756
rect 8429 11644 8431 11683
rect 8533 11644 8535 11683
rect 8429 11571 8431 11610
rect 8533 11571 8535 11610
rect 8429 11498 8431 11537
rect 8533 11498 8535 11537
rect 8429 11425 8431 11464
rect 8533 11425 8535 11464
rect 8429 11352 8431 11391
rect 8533 11352 8535 11391
rect 8429 11279 8431 11318
rect 8533 11279 8535 11318
rect 8429 11206 8431 11245
rect 8533 11206 8535 11245
rect 8429 11133 8431 11172
rect 8533 11133 8535 11172
rect 8429 11060 8431 11099
rect 8533 11060 8535 11099
rect 8429 10987 8431 11026
rect 8533 10987 8535 11026
rect 8429 10914 8431 10953
rect 8533 10914 8535 10953
rect 8429 10841 8431 10880
rect 8533 10841 8535 10880
rect 8429 10768 8431 10807
rect 8533 10768 8535 10807
rect 8429 10695 8431 10734
rect 8533 10695 8535 10734
rect 8429 10622 8431 10661
rect 8533 10622 8535 10661
rect 8429 10549 8431 10588
rect 8533 10549 8535 10588
rect 8429 10476 8431 10515
rect 8533 10476 8535 10515
rect 8429 10403 8431 10442
rect 8533 10403 8535 10442
rect 8429 10330 8431 10369
rect 8533 10330 8535 10369
rect 8429 10257 8431 10296
rect 8533 10257 8535 10296
rect 8429 10184 8431 10223
rect 8533 10184 8535 10223
rect 8429 10111 8431 10150
rect 8533 10111 8535 10150
rect 8429 10038 8431 10077
rect 8533 10038 8535 10077
rect 8429 9965 8431 10004
rect 8533 9965 8535 10004
rect 8429 9892 8431 9931
rect 8533 9892 8535 9931
rect 8429 9819 8431 9858
rect 8533 9819 8535 9858
rect 8429 9746 8431 9785
rect 8533 9746 8535 9785
rect 7733 9712 7805 9746
rect 7839 9712 7883 9746
rect 7917 9712 7961 9746
rect 7995 9712 8039 9746
rect 8073 9712 8116 9746
rect 8150 9712 8193 9746
rect 8227 9712 8270 9746
rect 8304 9712 8347 9746
rect 8381 9712 8429 9746
rect 7733 9705 8431 9712
rect 2050 9699 8431 9705
rect 2122 9665 2161 9699
rect 2195 9697 2234 9699
rect 2268 9697 2307 9699
rect 2341 9697 2380 9699
rect 2414 9697 2453 9699
rect 2487 9697 2526 9699
rect 2560 9697 2599 9699
rect 2633 9697 2672 9699
rect 2706 9697 2745 9699
rect 2779 9697 2818 9699
rect 2852 9697 2891 9699
rect 2925 9697 2964 9699
rect 2998 9697 3037 9699
rect 3071 9697 3110 9699
rect 3144 9697 3183 9699
rect 3217 9697 3256 9699
rect 3290 9697 3329 9699
rect 3363 9697 3402 9699
rect 3436 9697 3475 9699
rect 3509 9697 3548 9699
rect 3582 9697 3621 9699
rect 3655 9697 3694 9699
rect 3728 9697 3767 9699
rect 3801 9697 3840 9699
rect 3874 9697 3913 9699
rect 3947 9697 3986 9699
rect 4020 9697 4059 9699
rect 4093 9697 4132 9699
rect 4166 9697 4205 9699
rect 2195 9665 2208 9697
rect 2122 9627 2208 9665
rect 2122 9593 2161 9627
rect 2195 9595 2208 9627
rect 7695 9674 8431 9699
rect 7839 9640 7883 9674
rect 7917 9640 7961 9674
rect 7995 9640 8039 9674
rect 8073 9640 8116 9674
rect 8150 9640 8193 9674
rect 8227 9640 8270 9674
rect 8304 9640 8347 9674
rect 8381 9640 8424 9674
rect 7839 9638 8431 9640
rect 2195 9593 2234 9595
rect 2268 9593 2307 9595
rect 2341 9593 2380 9595
rect 2414 9593 2453 9595
rect 2487 9593 2526 9595
rect 2560 9593 2599 9595
rect 2633 9593 2672 9595
rect 2706 9593 2745 9595
rect 2779 9593 2818 9595
rect 2852 9593 2891 9595
rect 2925 9593 2964 9595
rect 2998 9593 3037 9595
rect 3071 9593 3110 9595
rect 3144 9593 3183 9595
rect 3217 9593 3256 9595
rect 3290 9593 3329 9595
rect 3363 9593 3402 9595
rect 3436 9593 3475 9595
rect 3509 9593 3548 9595
rect 3582 9593 3621 9595
rect 3655 9593 3694 9595
rect 3728 9593 3767 9595
rect 3801 9593 3840 9595
rect 3874 9593 3913 9595
rect 3947 9593 3986 9595
rect 4020 9593 4059 9595
rect 4093 9593 4132 9595
rect 4166 9593 4205 9595
rect 2050 9587 7733 9593
rect 2050 8938 2056 9587
rect 8381 9604 8431 9638
rect 8533 9604 8535 9712
rect 8381 9570 8535 9604
rect 8381 9536 8415 9570
rect 8449 9536 8535 9570
rect 1938 8874 1946 8938
rect 2048 8874 2056 8938
rect 1938 8840 1944 8874
rect 2050 8840 2056 8874
rect 1938 8801 1946 8840
rect 2048 8801 2056 8840
rect 1938 8767 1944 8801
rect 2050 8767 2056 8801
rect 1938 8728 1946 8767
rect 2048 8728 2056 8767
rect 1938 8694 1944 8728
rect 2050 8694 2056 8728
rect 1938 8655 1946 8694
rect 2048 8655 2056 8694
rect 1938 8621 1944 8655
rect 2050 8621 2056 8655
rect 1938 8582 1946 8621
rect 2048 8582 2056 8621
rect 1938 8548 1944 8582
rect 2050 8548 2056 8582
rect 1938 8509 1946 8548
rect 2048 8509 2056 8548
rect 1938 8475 1944 8509
rect 2050 8475 2056 8509
rect 1938 8436 1946 8475
rect 2048 8436 2056 8475
rect 1938 8402 1944 8436
rect 2050 8402 2056 8436
rect 1938 8363 1946 8402
rect 2048 8363 2056 8402
rect 1938 8329 1944 8363
rect 2050 8329 2056 8363
rect 1938 8290 1946 8329
rect 2048 8290 2056 8329
rect 1938 8256 1944 8290
rect 2050 8256 2056 8290
rect 1938 8217 1946 8256
rect 2048 8217 2056 8256
rect 1938 8183 1944 8217
rect 2050 8183 2056 8217
rect 1938 8144 1946 8183
rect 2048 8144 2056 8183
rect 1938 8110 1944 8144
rect 2050 8110 2056 8144
rect 1938 8071 1946 8110
rect 2048 8071 2056 8110
rect 1938 8037 1944 8071
rect 2050 8037 2056 8071
rect 1938 7998 1946 8037
rect 2048 7998 2056 8037
rect 1938 7964 1944 7998
rect 2050 7964 2056 7998
rect 1938 7925 1946 7964
rect 2048 7925 2056 7964
rect 1938 7891 1944 7925
rect 2050 7891 2056 7925
rect 1938 7852 1946 7891
rect 2048 7852 2056 7891
rect 1938 7818 1944 7852
rect 2050 7818 2056 7852
rect 1938 7779 1946 7818
rect 2048 7779 2056 7818
rect 1938 7745 1944 7779
rect 2050 7745 2056 7779
rect 1938 7706 1946 7745
rect 2048 7706 2056 7745
rect 1938 7672 1944 7706
rect 2050 7672 2056 7706
rect 1938 7633 1946 7672
rect 2048 7633 2056 7672
rect 1938 7599 1944 7633
rect 2050 7599 2056 7633
rect 1938 7560 1946 7599
rect 2048 7560 2056 7599
rect 1938 7526 1944 7560
rect 2050 7526 2056 7560
rect 1938 7487 1946 7526
rect 2048 7487 2056 7526
rect 1938 7453 1944 7487
rect 2050 7453 2056 7487
rect 1938 7414 1946 7453
rect 2048 7414 2056 7453
rect 1938 7380 1944 7414
rect 2050 7380 2056 7414
rect 1938 7341 1946 7380
rect 2048 7341 2056 7380
rect 1938 3491 1944 7341
rect 2050 3491 2056 7341
rect 2141 9449 7613 9455
rect 2141 9443 2359 9449
rect 2319 9430 2359 9443
rect 2393 9430 2432 9449
rect 2466 9430 2505 9449
rect 2539 9430 2578 9449
rect 2612 9430 2651 9449
rect 2685 9430 2724 9449
rect 2758 9430 2797 9449
rect 2831 9430 2870 9449
rect 2904 9430 2943 9449
rect 2977 9430 3016 9449
rect 3050 9430 3089 9449
rect 3123 9430 3162 9449
rect 3196 9430 3235 9449
rect 3269 9430 3308 9449
rect 3342 9430 3381 9449
rect 3415 9430 3454 9449
rect 3488 9430 3527 9449
rect 3561 9430 3600 9449
rect 3634 9430 3673 9449
rect 3707 9430 3746 9449
rect 3780 9430 3819 9449
rect 3853 9430 3892 9449
rect 3926 9430 3965 9449
rect 3999 9430 4038 9449
rect 4072 9430 4111 9449
rect 4145 9430 4184 9449
rect 2338 9415 2359 9430
rect 2407 9415 2432 9430
rect 2476 9415 2505 9430
rect 2545 9415 2578 9430
rect 2338 9396 2373 9415
rect 2407 9396 2442 9415
rect 2476 9396 2511 9415
rect 2545 9396 2580 9415
rect 2614 9396 2649 9430
rect 2685 9415 2718 9430
rect 2758 9415 2787 9430
rect 2831 9415 2856 9430
rect 2904 9415 2925 9430
rect 2977 9415 2994 9430
rect 3050 9415 3062 9430
rect 3123 9415 3130 9430
rect 3196 9415 3198 9430
rect 2683 9396 2718 9415
rect 2752 9396 2787 9415
rect 2821 9396 2856 9415
rect 2890 9396 2925 9415
rect 2959 9396 2994 9415
rect 3028 9396 3062 9415
rect 3096 9396 3130 9415
rect 3164 9396 3198 9415
rect 3232 9415 3235 9430
rect 3300 9415 3308 9430
rect 3368 9415 3381 9430
rect 3436 9415 3454 9430
rect 3504 9415 3527 9430
rect 3572 9415 3600 9430
rect 3640 9415 3673 9430
rect 3232 9396 3266 9415
rect 3300 9396 3334 9415
rect 3368 9396 3402 9415
rect 3436 9396 3470 9415
rect 3504 9396 3538 9415
rect 3572 9396 3606 9415
rect 3640 9396 3674 9415
rect 3708 9396 3742 9430
rect 3780 9415 3810 9430
rect 3853 9415 3878 9430
rect 3926 9415 3946 9430
rect 3999 9415 4014 9430
rect 4072 9415 4082 9430
rect 4145 9415 4150 9430
rect 3776 9396 3810 9415
rect 3844 9396 3878 9415
rect 3912 9396 3946 9415
rect 3980 9396 4014 9415
rect 4048 9396 4082 9415
rect 4116 9396 4150 9415
rect 4218 9430 4257 9449
rect 4291 9430 4330 9449
rect 4364 9430 4403 9449
rect 4437 9430 4476 9449
rect 4510 9430 4549 9449
rect 4583 9430 4622 9449
rect 4656 9430 4694 9449
rect 4728 9430 4766 9449
rect 4800 9430 4838 9449
rect 4872 9430 4910 9449
rect 4944 9430 4982 9449
rect 5016 9430 5054 9449
rect 5088 9430 5126 9449
rect 5160 9430 5198 9449
rect 5232 9430 5270 9449
rect 5304 9430 5342 9449
rect 5376 9430 5414 9449
rect 5448 9430 5486 9449
rect 5520 9430 5558 9449
rect 5592 9430 5630 9449
rect 5664 9430 5702 9449
rect 5736 9430 5774 9449
rect 5808 9430 5846 9449
rect 5880 9430 5918 9449
rect 5952 9430 5990 9449
rect 6024 9430 6062 9449
rect 6096 9430 6134 9449
rect 6168 9430 6206 9449
rect 6240 9430 6278 9449
rect 6312 9430 6350 9449
rect 6384 9430 6422 9449
rect 6456 9430 6494 9449
rect 6528 9430 6566 9449
rect 6600 9430 6638 9449
rect 6672 9430 6710 9449
rect 6744 9430 6782 9449
rect 6816 9430 6854 9449
rect 6888 9430 6926 9449
rect 6960 9430 6998 9449
rect 7032 9430 7070 9449
rect 7104 9430 7142 9449
rect 7176 9430 7214 9449
rect 7248 9430 7286 9449
rect 7320 9430 7358 9449
rect 7392 9437 7613 9449
rect 7392 9430 7493 9437
rect 4184 9396 4218 9415
rect 4252 9415 4257 9430
rect 4320 9415 4330 9430
rect 4388 9415 4403 9430
rect 4456 9415 4476 9430
rect 4524 9415 4549 9430
rect 4592 9415 4622 9430
rect 4252 9396 4286 9415
rect 4320 9396 4354 9415
rect 4388 9396 4422 9415
rect 4456 9396 4490 9415
rect 4524 9396 4558 9415
rect 4592 9396 4626 9415
rect 4660 9396 4694 9430
rect 4728 9396 4762 9430
rect 4800 9415 4830 9430
rect 4872 9415 4898 9430
rect 4944 9415 4966 9430
rect 5016 9415 5034 9430
rect 5088 9415 5102 9430
rect 5160 9415 5170 9430
rect 5232 9415 5238 9430
rect 5304 9415 5306 9430
rect 4796 9396 4830 9415
rect 4864 9396 4898 9415
rect 4932 9396 4966 9415
rect 5000 9396 5034 9415
rect 5068 9396 5102 9415
rect 5136 9396 5170 9415
rect 5204 9396 5238 9415
rect 5272 9396 5306 9415
rect 5340 9415 5342 9430
rect 5408 9415 5414 9430
rect 5476 9415 5486 9430
rect 5544 9415 5558 9430
rect 5612 9415 5630 9430
rect 5680 9415 5702 9430
rect 5748 9415 5774 9430
rect 5816 9415 5846 9430
rect 5340 9396 5374 9415
rect 5408 9396 5442 9415
rect 5476 9396 5510 9415
rect 5544 9396 5578 9415
rect 5612 9396 5646 9415
rect 5680 9396 5714 9415
rect 5748 9396 5782 9415
rect 5816 9396 5850 9415
rect 5884 9396 5918 9430
rect 5952 9396 5986 9430
rect 6024 9415 6054 9430
rect 6096 9415 6122 9430
rect 6168 9415 6190 9430
rect 6240 9415 6258 9430
rect 6312 9415 6326 9430
rect 6384 9415 6394 9430
rect 6456 9415 6462 9430
rect 6528 9415 6530 9430
rect 6020 9396 6054 9415
rect 6088 9396 6122 9415
rect 6156 9396 6190 9415
rect 6224 9396 6258 9415
rect 6292 9396 6326 9415
rect 6360 9396 6394 9415
rect 6428 9396 6462 9415
rect 6496 9396 6530 9415
rect 6564 9415 6566 9430
rect 6632 9415 6638 9430
rect 6700 9415 6710 9430
rect 6768 9415 6782 9430
rect 6836 9415 6854 9430
rect 6904 9415 6926 9430
rect 6972 9415 6998 9430
rect 7040 9415 7070 9430
rect 6564 9396 6598 9415
rect 6632 9396 6666 9415
rect 6700 9396 6734 9415
rect 6768 9396 6802 9415
rect 6836 9396 6870 9415
rect 6904 9396 6938 9415
rect 6972 9396 7006 9415
rect 7040 9396 7074 9415
rect 7108 9396 7142 9430
rect 7176 9396 7210 9430
rect 7248 9415 7278 9430
rect 7320 9415 7346 9430
rect 7392 9415 7414 9430
rect 7244 9396 7278 9415
rect 7312 9396 7346 9415
rect 7380 9396 7414 9415
rect 7448 9403 7493 9430
rect 7527 9403 7579 9437
rect 7448 9396 7613 9403
rect 2319 9362 2334 9396
rect 2324 9328 2334 9362
rect 7487 9370 7613 9396
rect 7521 9365 7613 9370
rect 2514 9340 2553 9341
rect 2587 9340 2626 9341
rect 2660 9340 2699 9341
rect 2733 9340 2772 9341
rect 2806 9340 2845 9341
rect 2879 9340 2918 9341
rect 2952 9340 2991 9341
rect 3025 9340 3064 9341
rect 3098 9340 3137 9341
rect 3171 9340 3210 9341
rect 3244 9340 3283 9341
rect 3317 9340 3356 9341
rect 3390 9340 3429 9341
rect 3463 9340 3502 9341
rect 3536 9340 3575 9341
rect 3609 9340 3648 9341
rect 3682 9340 3721 9341
rect 3755 9340 3794 9341
rect 3828 9340 3867 9341
rect 3901 9340 3940 9341
rect 3974 9340 4013 9341
rect 4047 9340 4086 9341
rect 2319 9294 2334 9328
rect 2468 9307 2480 9340
rect 2522 9307 2553 9340
rect 2468 9306 2488 9307
rect 2522 9306 2556 9307
rect 2590 9306 2624 9340
rect 2660 9307 2692 9340
rect 2733 9307 2760 9340
rect 2806 9307 2828 9340
rect 2879 9307 2896 9340
rect 2952 9307 2964 9340
rect 3025 9307 3032 9340
rect 3098 9307 3100 9340
rect 2658 9306 2692 9307
rect 2726 9306 2760 9307
rect 2794 9306 2828 9307
rect 2862 9306 2896 9307
rect 2930 9306 2964 9307
rect 2998 9306 3032 9307
rect 3066 9306 3100 9307
rect 3134 9307 3137 9340
rect 3202 9307 3210 9340
rect 3270 9307 3283 9340
rect 3338 9307 3356 9340
rect 3406 9307 3429 9340
rect 3474 9307 3502 9340
rect 3542 9307 3575 9340
rect 3134 9306 3168 9307
rect 3202 9306 3236 9307
rect 3270 9306 3304 9307
rect 3338 9306 3372 9307
rect 3406 9306 3440 9307
rect 3474 9306 3508 9307
rect 3542 9306 3576 9307
rect 3610 9306 3644 9340
rect 3682 9307 3712 9340
rect 3755 9307 3780 9340
rect 3828 9307 3848 9340
rect 3901 9307 3916 9340
rect 3974 9307 3984 9340
rect 4047 9307 4052 9340
rect 3678 9306 3712 9307
rect 3746 9306 3780 9307
rect 3814 9306 3848 9307
rect 3882 9306 3916 9307
rect 3950 9306 3984 9307
rect 4018 9306 4052 9307
rect 4120 9340 4159 9341
rect 4193 9340 4232 9341
rect 4266 9340 4305 9341
rect 4339 9340 4378 9341
rect 4412 9340 4451 9341
rect 4485 9340 4524 9341
rect 4558 9340 4597 9341
rect 4631 9340 4670 9341
rect 4704 9340 4742 9341
rect 4776 9340 4814 9341
rect 4848 9340 4886 9341
rect 4920 9340 4958 9341
rect 4992 9340 5030 9341
rect 5064 9340 5102 9341
rect 5136 9340 5174 9341
rect 4086 9306 4120 9307
rect 4154 9307 4159 9340
rect 4222 9307 4232 9340
rect 4290 9307 4305 9340
rect 4358 9307 4378 9340
rect 4426 9307 4451 9340
rect 4494 9307 4524 9340
rect 4154 9306 4188 9307
rect 4222 9306 4256 9307
rect 4290 9306 4324 9307
rect 4358 9306 4392 9307
rect 4426 9306 4460 9307
rect 4494 9306 4528 9307
rect 4562 9306 4596 9340
rect 4631 9307 4664 9340
rect 4704 9307 4732 9340
rect 4776 9307 4800 9340
rect 4848 9307 4868 9340
rect 4920 9307 4936 9340
rect 4992 9307 5004 9340
rect 5064 9307 5072 9340
rect 5136 9307 5140 9340
rect 4630 9306 4664 9307
rect 4698 9306 4732 9307
rect 4766 9306 4800 9307
rect 4834 9306 4868 9307
rect 4902 9306 4936 9307
rect 4970 9306 5004 9307
rect 5038 9306 5072 9307
rect 5106 9306 5140 9307
rect 5208 9340 5246 9341
rect 5280 9340 5318 9341
rect 5352 9340 5390 9341
rect 5424 9340 5462 9341
rect 5496 9340 5534 9341
rect 5568 9340 5606 9341
rect 5640 9340 5678 9341
rect 5712 9340 5750 9341
rect 5784 9340 5822 9341
rect 5856 9340 5894 9341
rect 5928 9340 5966 9341
rect 6000 9340 6038 9341
rect 6072 9340 6110 9341
rect 6144 9340 6182 9341
rect 6216 9340 6254 9341
rect 6288 9340 6326 9341
rect 6360 9340 6398 9341
rect 5174 9306 5208 9307
rect 5242 9307 5246 9340
rect 5310 9307 5318 9340
rect 5378 9307 5390 9340
rect 5446 9307 5462 9340
rect 5514 9307 5534 9340
rect 5582 9307 5606 9340
rect 5650 9307 5678 9340
rect 5718 9307 5750 9340
rect 5242 9306 5276 9307
rect 5310 9306 5344 9307
rect 5378 9306 5412 9307
rect 5446 9306 5480 9307
rect 5514 9306 5548 9307
rect 5582 9306 5616 9307
rect 5650 9306 5684 9307
rect 5718 9306 5752 9307
rect 5786 9306 5820 9340
rect 5856 9307 5888 9340
rect 5928 9307 5956 9340
rect 6000 9307 6024 9340
rect 6072 9307 6092 9340
rect 6144 9307 6160 9340
rect 6216 9307 6228 9340
rect 6288 9307 6296 9340
rect 6360 9307 6364 9340
rect 5854 9306 5888 9307
rect 5922 9306 5956 9307
rect 5990 9306 6024 9307
rect 6058 9306 6092 9307
rect 6126 9306 6160 9307
rect 6194 9306 6228 9307
rect 6262 9306 6296 9307
rect 6330 9306 6364 9307
rect 6432 9340 6470 9341
rect 6504 9340 6542 9341
rect 6576 9340 6614 9341
rect 6648 9340 6686 9341
rect 6720 9340 6758 9341
rect 6792 9340 6830 9341
rect 6864 9340 6902 9341
rect 6936 9340 6974 9341
rect 7008 9340 7046 9341
rect 7080 9340 7118 9341
rect 7152 9340 7190 9341
rect 7224 9340 7262 9341
rect 7296 9340 7334 9341
rect 6398 9306 6432 9307
rect 6466 9307 6470 9340
rect 6534 9307 6542 9340
rect 6602 9307 6614 9340
rect 6670 9307 6686 9340
rect 6738 9307 6758 9340
rect 6806 9307 6830 9340
rect 6874 9307 6902 9340
rect 6942 9307 6974 9340
rect 6466 9306 6500 9307
rect 6534 9306 6568 9307
rect 6602 9306 6636 9307
rect 6670 9306 6704 9307
rect 6738 9306 6772 9307
rect 6806 9306 6840 9307
rect 6874 9306 6908 9307
rect 6942 9306 6976 9307
rect 7010 9306 7044 9340
rect 7080 9307 7112 9340
rect 7152 9307 7180 9340
rect 7224 9307 7248 9340
rect 7296 9307 7316 9340
rect 7368 9307 7380 9340
rect 7078 9306 7112 9307
rect 7146 9306 7180 9307
rect 7214 9306 7248 9307
rect 7282 9306 7316 9307
rect 7350 9306 7380 9307
rect 7487 9331 7493 9336
rect 7527 9331 7579 9365
rect 2324 9260 2334 9294
rect 2319 9226 2334 9260
rect 2324 9192 2334 9226
rect 7487 9302 7613 9331
rect 7521 9293 7613 9302
rect 7487 9259 7493 9268
rect 7527 9259 7579 9293
rect 7487 9234 7613 9259
rect 7521 9221 7613 9234
rect 2319 9158 2334 9192
rect 2324 9124 2334 9158
rect 2319 9090 2334 9124
rect 2324 9056 2334 9090
rect 2319 9022 2334 9056
rect 2324 8988 2334 9022
rect 2319 8954 2334 8988
rect 2324 8920 2334 8954
rect 2319 8886 2334 8920
rect 2324 8852 2334 8886
rect 2319 8818 2334 8852
rect 2324 8784 2334 8818
rect 2319 8750 2334 8784
rect 2324 8716 2334 8750
rect 2319 8682 2334 8716
rect 2324 8648 2334 8682
rect 2319 8614 2334 8648
rect 2324 8580 2334 8614
rect 2319 8546 2334 8580
rect 2324 8512 2334 8546
rect 2319 8478 2334 8512
rect 2324 8444 2334 8478
rect 2319 8410 2334 8444
rect 2324 8376 2334 8410
rect 2319 8342 2334 8376
rect 2324 8308 2334 8342
rect 2319 8274 2334 8308
rect 2324 8240 2334 8274
rect 2319 8206 2334 8240
rect 2324 8172 2334 8206
rect 2319 8138 2334 8172
rect 2324 8104 2334 8138
rect 2319 8070 2334 8104
rect 2324 8036 2334 8070
rect 2319 8002 2334 8036
rect 2324 7968 2334 8002
rect 2319 7934 2334 7968
rect 2324 7900 2334 7934
rect 2319 7866 2334 7900
rect 2324 7832 2334 7866
rect 2417 9178 2422 9212
rect 2456 9178 2461 9212
rect 2417 9139 2461 9178
rect 2417 9105 2422 9139
rect 2456 9105 2461 9139
rect 2417 9066 2461 9105
rect 2417 9032 2422 9066
rect 2456 9032 2461 9066
rect 2417 8993 2461 9032
rect 2417 8959 2422 8993
rect 2456 8959 2461 8993
rect 2417 8920 2461 8959
rect 2417 8886 2422 8920
rect 2456 8886 2461 8920
rect 2417 8847 2461 8886
rect 2417 8813 2422 8847
rect 2456 8813 2461 8847
rect 2417 8774 2461 8813
rect 2417 8740 2422 8774
rect 2456 8740 2461 8774
rect 2417 8701 2461 8740
rect 2417 8667 2422 8701
rect 2456 8667 2461 8701
rect 2417 8628 2461 8667
rect 2417 8594 2422 8628
rect 2456 8594 2461 8628
rect 2417 8554 2461 8594
rect 2417 8520 2422 8554
rect 2456 8520 2461 8554
rect 2417 8480 2461 8520
rect 2417 8446 2422 8480
rect 2456 8446 2461 8480
rect 2417 8406 2461 8446
rect 2417 8372 2422 8406
rect 2456 8372 2461 8406
rect 2417 8332 2461 8372
rect 2417 8298 2422 8332
rect 2456 8298 2461 8332
rect 2417 8258 2461 8298
rect 2417 8224 2422 8258
rect 2456 8224 2461 8258
rect 2417 8184 2461 8224
rect 2417 8150 2422 8184
rect 2456 8150 2461 8184
rect 2417 8110 2461 8150
rect 2417 8076 2422 8110
rect 2456 8076 2461 8110
rect 2417 8036 2461 8076
rect 2417 8002 2422 8036
rect 2456 8002 2461 8036
rect 2417 7962 2461 8002
rect 2417 7928 2422 7962
rect 2456 7928 2461 7962
rect 2417 7888 2461 7928
rect 2417 7854 2422 7888
rect 2456 7854 2461 7888
rect 4074 9178 4079 9212
rect 4113 9178 4118 9212
rect 4074 9139 4118 9178
rect 4074 9105 4079 9139
rect 4113 9105 4118 9139
rect 4074 9066 4118 9105
rect 4074 9032 4079 9066
rect 4113 9032 4118 9066
rect 4074 8993 4118 9032
rect 4074 8959 4079 8993
rect 4113 8959 4118 8993
rect 4074 8920 4118 8959
rect 4074 8886 4079 8920
rect 4113 8886 4118 8920
rect 4074 8847 4118 8886
rect 4074 8813 4079 8847
rect 4113 8813 4118 8847
rect 4074 8774 4118 8813
rect 4074 8740 4079 8774
rect 4113 8740 4118 8774
rect 4074 8701 4118 8740
rect 4074 8667 4079 8701
rect 4113 8667 4118 8701
rect 4074 8628 4118 8667
rect 4074 8594 4079 8628
rect 4113 8594 4118 8628
rect 4074 8554 4118 8594
rect 4074 8520 4079 8554
rect 4113 8520 4118 8554
rect 4074 8480 4118 8520
rect 4074 8446 4079 8480
rect 4113 8446 4118 8480
rect 4074 8406 4118 8446
rect 4074 8372 4079 8406
rect 4113 8372 4118 8406
rect 4074 8332 4118 8372
rect 4074 8298 4079 8332
rect 4113 8298 4118 8332
rect 4074 8258 4118 8298
rect 4074 8224 4079 8258
rect 4113 8224 4118 8258
rect 4074 8184 4118 8224
rect 4074 8150 4079 8184
rect 4113 8150 4118 8184
rect 4074 8110 4118 8150
rect 4074 8076 4079 8110
rect 4113 8076 4118 8110
rect 4074 8036 4118 8076
rect 4074 8002 4079 8036
rect 4113 8002 4118 8036
rect 4074 7962 4118 8002
rect 4074 7928 4079 7962
rect 4113 7928 4118 7962
rect 4074 7888 4118 7928
rect 4074 7854 4079 7888
rect 4113 7854 4118 7888
rect 5732 9178 5737 9212
rect 5771 9178 5776 9212
rect 5732 9139 5776 9178
rect 5732 9105 5737 9139
rect 5771 9105 5776 9139
rect 5732 9066 5776 9105
rect 5732 9032 5737 9066
rect 5771 9032 5776 9066
rect 5732 8993 5776 9032
rect 5732 8959 5737 8993
rect 5771 8959 5776 8993
rect 5732 8920 5776 8959
rect 5732 8886 5737 8920
rect 5771 8886 5776 8920
rect 5732 8847 5776 8886
rect 5732 8813 5737 8847
rect 5771 8813 5776 8847
rect 5732 8774 5776 8813
rect 5732 8740 5737 8774
rect 5771 8740 5776 8774
rect 5732 8701 5776 8740
rect 5732 8667 5737 8701
rect 5771 8667 5776 8701
rect 5732 8628 5776 8667
rect 5732 8594 5737 8628
rect 5771 8594 5776 8628
rect 5732 8554 5776 8594
rect 5732 8520 5737 8554
rect 5771 8520 5776 8554
rect 5732 8480 5776 8520
rect 5732 8446 5737 8480
rect 5771 8446 5776 8480
rect 5732 8406 5776 8446
rect 5732 8372 5737 8406
rect 5771 8372 5776 8406
rect 5732 8332 5776 8372
rect 5732 8298 5737 8332
rect 5771 8298 5776 8332
rect 5732 8258 5776 8298
rect 5732 8224 5737 8258
rect 5771 8224 5776 8258
rect 5732 8184 5776 8224
rect 5732 8150 5737 8184
rect 5771 8150 5776 8184
rect 5732 8110 5776 8150
rect 5732 8076 5737 8110
rect 5771 8076 5776 8110
rect 5732 8036 5776 8076
rect 5732 8002 5737 8036
rect 5771 8002 5776 8036
rect 5732 7962 5776 8002
rect 5732 7928 5737 7962
rect 5771 7928 5776 7962
rect 5732 7888 5776 7928
rect 5732 7854 5737 7888
rect 5771 7854 5776 7888
rect 7381 9178 7386 9212
rect 7420 9178 7425 9212
rect 7381 9139 7425 9178
rect 7381 9105 7386 9139
rect 7420 9105 7425 9139
rect 7381 9066 7425 9105
rect 7381 9032 7386 9066
rect 7420 9032 7425 9066
rect 7381 8993 7425 9032
rect 7381 8959 7386 8993
rect 7420 8959 7425 8993
rect 7381 8920 7425 8959
rect 7381 8886 7386 8920
rect 7420 8886 7425 8920
rect 7381 8847 7425 8886
rect 7381 8813 7386 8847
rect 7420 8813 7425 8847
rect 7381 8774 7425 8813
rect 7381 8740 7386 8774
rect 7420 8740 7425 8774
rect 7381 8701 7425 8740
rect 7381 8667 7386 8701
rect 7420 8667 7425 8701
rect 7381 8628 7425 8667
rect 7381 8594 7386 8628
rect 7420 8594 7425 8628
rect 7381 8554 7425 8594
rect 7381 8520 7386 8554
rect 7420 8520 7425 8554
rect 7381 8480 7425 8520
rect 7381 8446 7386 8480
rect 7420 8446 7425 8480
rect 7381 8406 7425 8446
rect 7381 8372 7386 8406
rect 7420 8372 7425 8406
rect 7381 8332 7425 8372
rect 7381 8298 7386 8332
rect 7420 8298 7425 8332
rect 7381 8258 7425 8298
rect 7381 8224 7386 8258
rect 7420 8224 7425 8258
rect 7381 8184 7425 8224
rect 7381 8150 7386 8184
rect 7420 8150 7425 8184
rect 7381 8110 7425 8150
rect 7381 8076 7386 8110
rect 7420 8076 7425 8110
rect 7381 8036 7425 8076
rect 7381 8002 7386 8036
rect 7420 8002 7425 8036
rect 7381 7962 7425 8002
rect 7381 7928 7386 7962
rect 7420 7928 7425 7962
rect 7381 7888 7425 7928
rect 7381 7854 7386 7888
rect 7420 7854 7425 7888
rect 7487 9187 7493 9200
rect 7527 9187 7579 9221
rect 7487 9166 7613 9187
rect 7521 9149 7613 9166
rect 7487 9115 7493 9132
rect 7527 9115 7579 9149
rect 7487 9098 7613 9115
rect 7521 9077 7613 9098
rect 7487 9043 7493 9064
rect 7527 9043 7579 9077
rect 7487 9030 7613 9043
rect 7521 9005 7613 9030
rect 7487 8971 7493 8996
rect 7527 8971 7579 9005
rect 7487 8962 7613 8971
rect 7521 8933 7613 8962
rect 7487 8899 7493 8928
rect 7527 8899 7579 8933
rect 7487 8894 7613 8899
rect 7521 8861 7613 8894
rect 7487 8827 7493 8860
rect 7527 8827 7579 8861
rect 7487 8826 7613 8827
rect 7521 8792 7613 8826
rect 7487 8789 7613 8792
rect 7487 8758 7493 8789
rect 7527 8755 7579 8789
rect 7521 8724 7613 8755
rect 7487 8717 7613 8724
rect 7487 8690 7493 8717
rect 7527 8683 7579 8717
rect 7521 8656 7613 8683
rect 7487 8645 7613 8656
rect 7487 8622 7493 8645
rect 7527 8611 7579 8645
rect 7521 8588 7613 8611
rect 7487 8573 7613 8588
rect 7487 8554 7493 8573
rect 7527 8539 7579 8573
rect 7521 8520 7613 8539
rect 7487 8501 7613 8520
rect 7487 8486 7493 8501
rect 7527 8467 7579 8501
rect 7521 8452 7613 8467
rect 7487 8429 7613 8452
rect 7487 8418 7493 8429
rect 7527 8395 7579 8429
rect 7521 8384 7613 8395
rect 7487 8357 7613 8384
rect 7487 8350 7493 8357
rect 7527 8323 7579 8357
rect 7521 8316 7613 8323
rect 7487 8285 7613 8316
rect 7487 8282 7493 8285
rect 7527 8251 7579 8285
rect 7521 8248 7613 8251
rect 7487 8214 7613 8248
rect 7521 8213 7613 8214
rect 7487 8179 7493 8180
rect 7527 8179 7579 8213
rect 7487 8146 7613 8179
rect 7521 8141 7613 8146
rect 7487 8107 7493 8112
rect 7527 8107 7579 8141
rect 7487 8078 7613 8107
rect 7521 8069 7613 8078
rect 7487 8035 7493 8044
rect 7527 8035 7579 8069
rect 7487 8010 7613 8035
rect 7521 7997 7613 8010
rect 7487 7963 7493 7976
rect 7527 7963 7579 7997
rect 7487 7942 7613 7963
rect 7521 7925 7613 7942
rect 7487 7891 7493 7908
rect 7527 7891 7579 7925
rect 7487 7874 7613 7891
rect 2319 7798 2334 7832
rect 2324 7764 2334 7798
rect 2319 7730 2334 7764
rect 2324 7696 2334 7730
rect 2319 7687 2334 7696
rect 7521 7853 7613 7874
rect 7487 7819 7493 7840
rect 7527 7819 7579 7853
rect 7487 7806 7613 7819
rect 7521 7781 7613 7806
rect 7487 7747 7493 7772
rect 7527 7747 7579 7781
rect 7487 7738 7613 7747
rect 7521 7709 7613 7738
rect 7487 7687 7493 7704
rect 2319 7681 7493 7687
rect 2319 7662 2357 7681
rect 2324 7647 2357 7662
rect 2392 7647 2427 7681
rect 2463 7647 2496 7681
rect 2535 7647 2565 7681
rect 2607 7647 2634 7681
rect 2679 7647 2703 7681
rect 2751 7647 2772 7681
rect 2823 7647 2841 7681
rect 2895 7647 2910 7681
rect 2967 7647 2979 7681
rect 3039 7647 3048 7681
rect 3111 7647 3117 7681
rect 3183 7647 3186 7681
rect 3220 7647 3221 7681
rect 3289 7647 3293 7681
rect 3358 7647 3365 7681
rect 3427 7647 3437 7681
rect 3496 7647 3509 7681
rect 3565 7647 3581 7681
rect 3634 7647 3653 7681
rect 3703 7647 3725 7681
rect 3772 7647 3797 7681
rect 3841 7647 3869 7681
rect 3909 7647 3941 7681
rect 3977 7647 4011 7681
rect 4047 7647 4079 7681
rect 4119 7647 4147 7681
rect 4191 7647 4215 7681
rect 4263 7647 4283 7681
rect 4335 7647 4351 7681
rect 4407 7647 4419 7681
rect 4479 7647 4487 7681
rect 4551 7647 4555 7681
rect 4657 7647 4661 7681
rect 4725 7647 4733 7681
rect 4793 7647 4805 7681
rect 4861 7647 4877 7681
rect 4929 7647 4949 7681
rect 4997 7647 5021 7681
rect 5065 7647 5093 7681
rect 5133 7647 5165 7681
rect 5201 7647 5235 7681
rect 5271 7647 5303 7681
rect 5343 7647 5371 7681
rect 5415 7647 5439 7681
rect 5487 7647 5507 7681
rect 5559 7647 5575 7681
rect 5631 7647 5643 7681
rect 5703 7647 5711 7681
rect 5775 7647 5779 7681
rect 5881 7647 5885 7681
rect 5949 7647 5957 7681
rect 6017 7647 6029 7681
rect 6085 7647 6101 7681
rect 6153 7647 6173 7681
rect 6221 7647 6245 7681
rect 6289 7647 6317 7681
rect 6357 7647 6389 7681
rect 6425 7647 6459 7681
rect 6495 7647 6527 7681
rect 6567 7647 6595 7681
rect 6639 7647 6663 7681
rect 6711 7647 6731 7681
rect 6783 7647 6799 7681
rect 6855 7647 6867 7681
rect 6927 7647 6935 7681
rect 6999 7647 7003 7681
rect 7105 7647 7109 7681
rect 7173 7647 7181 7681
rect 7241 7647 7253 7681
rect 7309 7647 7325 7681
rect 7377 7647 7397 7681
rect 7445 7675 7493 7681
rect 7527 7675 7579 7709
rect 7445 7670 7613 7675
rect 7445 7647 7487 7670
rect 2324 7641 7487 7647
rect 2324 7628 2334 7641
rect 2319 7594 2334 7628
rect 2324 7560 2334 7594
rect 2319 7526 2334 7560
rect 7521 7637 7613 7670
rect 7487 7603 7493 7636
rect 7527 7603 7579 7637
rect 7487 7602 7613 7603
rect 7521 7568 7613 7602
rect 7487 7565 7613 7568
rect 2324 7492 2334 7526
rect 2468 7506 2480 7540
rect 2522 7506 2553 7540
rect 2590 7506 2624 7540
rect 2660 7506 2692 7540
rect 2733 7506 2760 7540
rect 2806 7506 2828 7540
rect 2879 7506 2896 7540
rect 2952 7506 2964 7540
rect 3025 7506 3032 7540
rect 3098 7506 3100 7540
rect 3134 7506 3137 7540
rect 3202 7506 3210 7540
rect 3270 7506 3283 7540
rect 3338 7506 3356 7540
rect 3406 7506 3429 7540
rect 3474 7506 3502 7540
rect 3542 7506 3575 7540
rect 3610 7506 3644 7540
rect 3682 7506 3712 7540
rect 3755 7506 3780 7540
rect 3828 7506 3848 7540
rect 3901 7506 3916 7540
rect 3974 7506 3984 7540
rect 4047 7506 4052 7540
rect 4154 7506 4159 7540
rect 4222 7506 4232 7540
rect 4290 7506 4305 7540
rect 4358 7506 4378 7540
rect 4426 7506 4451 7540
rect 4494 7506 4524 7540
rect 4562 7506 4596 7540
rect 4631 7506 4664 7540
rect 4704 7506 4732 7540
rect 4776 7506 4800 7540
rect 4848 7506 4868 7540
rect 4920 7506 4936 7540
rect 4992 7506 5004 7540
rect 5064 7506 5072 7540
rect 5136 7506 5140 7540
rect 5242 7506 5246 7540
rect 5310 7506 5318 7540
rect 5378 7506 5390 7540
rect 5446 7506 5462 7540
rect 5514 7506 5534 7540
rect 5582 7506 5606 7540
rect 5650 7506 5678 7540
rect 5718 7506 5750 7540
rect 5786 7506 5820 7540
rect 5856 7506 5888 7540
rect 5928 7506 5956 7540
rect 6000 7506 6024 7540
rect 6072 7506 6092 7540
rect 6144 7506 6160 7540
rect 6216 7506 6228 7540
rect 6288 7506 6296 7540
rect 6360 7506 6364 7540
rect 6466 7506 6470 7540
rect 6534 7506 6542 7540
rect 6602 7506 6614 7540
rect 6670 7506 6686 7540
rect 6738 7506 6758 7540
rect 6806 7506 6830 7540
rect 6874 7506 6902 7540
rect 6942 7506 6974 7540
rect 7010 7506 7044 7540
rect 7080 7506 7112 7540
rect 7152 7506 7180 7540
rect 7224 7506 7248 7540
rect 7296 7506 7316 7540
rect 7368 7506 7380 7540
rect 7487 7534 7493 7565
rect 7527 7531 7579 7565
rect 2319 7458 2334 7492
rect 2324 7424 2334 7458
rect 2319 7390 2334 7424
rect 7521 7500 7613 7531
rect 7487 7493 7613 7500
rect 7487 7466 7493 7493
rect 7527 7459 7579 7493
rect 7521 7432 7613 7459
rect 7487 7421 7613 7432
rect 2324 7356 2334 7390
rect 2319 7322 2334 7356
rect 2324 7288 2334 7322
rect 2319 7254 2334 7288
rect 2324 7220 2334 7254
rect 2319 7186 2334 7220
rect 2324 7152 2334 7186
rect 2319 7118 2334 7152
rect 2324 7084 2334 7118
rect 2319 7050 2334 7084
rect 2324 7016 2334 7050
rect 2319 6982 2334 7016
rect 2324 6948 2334 6982
rect 2319 6914 2334 6948
rect 2324 6880 2334 6914
rect 2319 6846 2334 6880
rect 2324 6812 2334 6846
rect 2319 6778 2334 6812
rect 2324 6744 2334 6778
rect 2319 6710 2334 6744
rect 2324 6676 2334 6710
rect 2319 6642 2334 6676
rect 2324 6608 2334 6642
rect 2319 6574 2334 6608
rect 2324 6540 2334 6574
rect 2319 6506 2334 6540
rect 2324 6472 2334 6506
rect 2319 6438 2334 6472
rect 2324 6404 2334 6438
rect 2319 6370 2334 6404
rect 2324 6336 2334 6370
rect 2319 6302 2334 6336
rect 2324 6268 2334 6302
rect 2319 6234 2334 6268
rect 2324 6200 2334 6234
rect 2319 6166 2334 6200
rect 2324 6132 2334 6166
rect 2319 6098 2334 6132
rect 2324 6064 2334 6098
rect 2319 6030 2334 6064
rect 2417 7378 2422 7412
rect 2456 7378 2461 7412
rect 2417 7339 2461 7378
rect 2417 7305 2422 7339
rect 2456 7305 2461 7339
rect 2417 7266 2461 7305
rect 2417 7232 2422 7266
rect 2456 7232 2461 7266
rect 2417 7193 2461 7232
rect 2417 7159 2422 7193
rect 2456 7159 2461 7193
rect 2417 7120 2461 7159
rect 2417 7086 2422 7120
rect 2456 7086 2461 7120
rect 2417 7047 2461 7086
rect 2417 7013 2422 7047
rect 2456 7013 2461 7047
rect 2417 6974 2461 7013
rect 2417 6940 2422 6974
rect 2456 6940 2461 6974
rect 2417 6901 2461 6940
rect 2417 6867 2422 6901
rect 2456 6867 2461 6901
rect 2417 6828 2461 6867
rect 2417 6794 2422 6828
rect 2456 6794 2461 6828
rect 2417 6754 2461 6794
rect 2417 6720 2422 6754
rect 2456 6720 2461 6754
rect 2417 6680 2461 6720
rect 2417 6646 2422 6680
rect 2456 6646 2461 6680
rect 2417 6606 2461 6646
rect 2417 6572 2422 6606
rect 2456 6572 2461 6606
rect 2417 6532 2461 6572
rect 2417 6498 2422 6532
rect 2456 6498 2461 6532
rect 2417 6458 2461 6498
rect 2417 6424 2422 6458
rect 2456 6424 2461 6458
rect 2417 6384 2461 6424
rect 2417 6350 2422 6384
rect 2456 6350 2461 6384
rect 2417 6310 2461 6350
rect 2417 6276 2422 6310
rect 2456 6276 2461 6310
rect 2417 6236 2461 6276
rect 2417 6202 2422 6236
rect 2456 6202 2461 6236
rect 2417 6162 2461 6202
rect 2417 6128 2422 6162
rect 2456 6128 2461 6162
rect 2417 6088 2461 6128
rect 2417 6054 2422 6088
rect 2456 6054 2461 6088
rect 4074 7378 4079 7412
rect 4113 7378 4118 7412
rect 4074 7339 4118 7378
rect 4074 7305 4079 7339
rect 4113 7305 4118 7339
rect 4074 7266 4118 7305
rect 4074 7232 4079 7266
rect 4113 7232 4118 7266
rect 4074 7193 4118 7232
rect 4074 7159 4079 7193
rect 4113 7159 4118 7193
rect 4074 7120 4118 7159
rect 4074 7086 4079 7120
rect 4113 7086 4118 7120
rect 4074 7047 4118 7086
rect 4074 7013 4079 7047
rect 4113 7013 4118 7047
rect 4074 6974 4118 7013
rect 4074 6940 4079 6974
rect 4113 6940 4118 6974
rect 4074 6901 4118 6940
rect 4074 6867 4079 6901
rect 4113 6867 4118 6901
rect 4074 6828 4118 6867
rect 4074 6794 4079 6828
rect 4113 6794 4118 6828
rect 4074 6754 4118 6794
rect 4074 6720 4079 6754
rect 4113 6720 4118 6754
rect 4074 6680 4118 6720
rect 4074 6646 4079 6680
rect 4113 6646 4118 6680
rect 4074 6606 4118 6646
rect 4074 6572 4079 6606
rect 4113 6572 4118 6606
rect 4074 6532 4118 6572
rect 4074 6498 4079 6532
rect 4113 6498 4118 6532
rect 4074 6458 4118 6498
rect 4074 6424 4079 6458
rect 4113 6424 4118 6458
rect 4074 6384 4118 6424
rect 4074 6350 4079 6384
rect 4113 6350 4118 6384
rect 4074 6310 4118 6350
rect 4074 6276 4079 6310
rect 4113 6276 4118 6310
rect 4074 6236 4118 6276
rect 4074 6202 4079 6236
rect 4113 6202 4118 6236
rect 4074 6162 4118 6202
rect 4074 6128 4079 6162
rect 4113 6128 4118 6162
rect 4074 6088 4118 6128
rect 4074 6054 4079 6088
rect 4113 6054 4118 6088
rect 5732 7378 5737 7412
rect 5771 7378 5776 7412
rect 5732 7339 5776 7378
rect 5732 7305 5737 7339
rect 5771 7305 5776 7339
rect 5732 7266 5776 7305
rect 5732 7232 5737 7266
rect 5771 7232 5776 7266
rect 5732 7193 5776 7232
rect 5732 7159 5737 7193
rect 5771 7159 5776 7193
rect 5732 7120 5776 7159
rect 5732 7086 5737 7120
rect 5771 7086 5776 7120
rect 5732 7047 5776 7086
rect 5732 7013 5737 7047
rect 5771 7013 5776 7047
rect 5732 6974 5776 7013
rect 5732 6940 5737 6974
rect 5771 6940 5776 6974
rect 5732 6901 5776 6940
rect 5732 6867 5737 6901
rect 5771 6867 5776 6901
rect 5732 6828 5776 6867
rect 5732 6794 5737 6828
rect 5771 6794 5776 6828
rect 5732 6754 5776 6794
rect 5732 6720 5737 6754
rect 5771 6720 5776 6754
rect 5732 6680 5776 6720
rect 5732 6646 5737 6680
rect 5771 6646 5776 6680
rect 5732 6606 5776 6646
rect 5732 6572 5737 6606
rect 5771 6572 5776 6606
rect 5732 6532 5776 6572
rect 5732 6498 5737 6532
rect 5771 6498 5776 6532
rect 5732 6458 5776 6498
rect 5732 6424 5737 6458
rect 5771 6424 5776 6458
rect 5732 6384 5776 6424
rect 5732 6350 5737 6384
rect 5771 6350 5776 6384
rect 5732 6310 5776 6350
rect 5732 6276 5737 6310
rect 5771 6276 5776 6310
rect 5732 6236 5776 6276
rect 5732 6202 5737 6236
rect 5771 6202 5776 6236
rect 5732 6162 5776 6202
rect 5732 6128 5737 6162
rect 5771 6128 5776 6162
rect 5732 6088 5776 6128
rect 5732 6054 5737 6088
rect 5771 6054 5776 6088
rect 7381 7378 7386 7412
rect 7420 7378 7425 7412
rect 7381 7339 7425 7378
rect 7381 7305 7386 7339
rect 7420 7305 7425 7339
rect 7381 7266 7425 7305
rect 7381 7232 7386 7266
rect 7420 7232 7425 7266
rect 7381 7193 7425 7232
rect 7381 7159 7386 7193
rect 7420 7159 7425 7193
rect 7381 7120 7425 7159
rect 7381 7086 7386 7120
rect 7420 7086 7425 7120
rect 7381 7047 7425 7086
rect 7381 7013 7386 7047
rect 7420 7013 7425 7047
rect 7381 6974 7425 7013
rect 7381 6940 7386 6974
rect 7420 6940 7425 6974
rect 7381 6901 7425 6940
rect 7381 6867 7386 6901
rect 7420 6867 7425 6901
rect 7381 6828 7425 6867
rect 7381 6794 7386 6828
rect 7420 6794 7425 6828
rect 7381 6754 7425 6794
rect 7381 6720 7386 6754
rect 7420 6720 7425 6754
rect 7381 6680 7425 6720
rect 7381 6646 7386 6680
rect 7420 6646 7425 6680
rect 7381 6606 7425 6646
rect 7381 6572 7386 6606
rect 7420 6572 7425 6606
rect 7381 6532 7425 6572
rect 7381 6498 7386 6532
rect 7420 6498 7425 6532
rect 7381 6458 7425 6498
rect 7381 6424 7386 6458
rect 7420 6424 7425 6458
rect 7381 6384 7425 6424
rect 7381 6350 7386 6384
rect 7420 6350 7425 6384
rect 7381 6310 7425 6350
rect 7381 6276 7386 6310
rect 7420 6276 7425 6310
rect 7381 6236 7425 6276
rect 7381 6202 7386 6236
rect 7420 6202 7425 6236
rect 7381 6162 7425 6202
rect 7381 6128 7386 6162
rect 7420 6128 7425 6162
rect 7381 6088 7425 6128
rect 7381 6054 7386 6088
rect 7420 6054 7425 6088
rect 7487 7398 7493 7421
rect 7527 7387 7579 7421
rect 7521 7364 7613 7387
rect 7487 7349 7613 7364
rect 7487 7330 7493 7349
rect 7527 7315 7579 7349
rect 7521 7296 7613 7315
rect 7487 7277 7613 7296
rect 7487 7262 7493 7277
rect 7527 7243 7579 7277
rect 7521 7228 7613 7243
rect 7487 7205 7613 7228
rect 7487 7194 7493 7205
rect 7527 7171 7579 7205
rect 7521 7160 7613 7171
rect 7487 7133 7613 7160
rect 7487 7126 7493 7133
rect 7527 7099 7579 7133
rect 7521 7092 7613 7099
rect 7487 7061 7613 7092
rect 7487 7058 7493 7061
rect 7527 7027 7579 7061
rect 7521 7024 7613 7027
rect 7487 6990 7613 7024
rect 7521 6989 7613 6990
rect 7487 6955 7493 6956
rect 7527 6955 7579 6989
rect 7487 6922 7613 6955
rect 7521 6917 7613 6922
rect 7487 6883 7493 6888
rect 7527 6883 7579 6917
rect 7487 6854 7613 6883
rect 7521 6845 7613 6854
rect 7487 6811 7493 6820
rect 7527 6811 7579 6845
rect 7487 6786 7613 6811
rect 7521 6773 7613 6786
rect 7487 6739 7493 6752
rect 7527 6739 7579 6773
rect 7487 6718 7613 6739
rect 7521 6701 7613 6718
rect 7487 6667 7493 6684
rect 7527 6667 7579 6701
rect 7487 6650 7613 6667
rect 7521 6629 7613 6650
rect 7487 6595 7493 6616
rect 7527 6595 7579 6629
rect 7487 6582 7613 6595
rect 7521 6557 7613 6582
rect 7487 6523 7493 6548
rect 7527 6523 7579 6557
rect 7487 6514 7613 6523
rect 7521 6485 7613 6514
rect 7487 6451 7493 6480
rect 7527 6451 7579 6485
rect 7487 6446 7613 6451
rect 7521 6413 7613 6446
rect 7487 6379 7493 6412
rect 7527 6379 7579 6413
rect 7487 6378 7613 6379
rect 7521 6344 7613 6378
rect 7487 6341 7613 6344
rect 7487 6310 7493 6341
rect 7527 6307 7579 6341
rect 7521 6276 7613 6307
rect 7487 6269 7613 6276
rect 7487 6242 7493 6269
rect 7527 6235 7579 6269
rect 7521 6208 7613 6235
rect 7487 6197 7613 6208
rect 7487 6174 7493 6197
rect 7527 6163 7579 6197
rect 7521 6140 7613 6163
rect 7487 6125 7613 6140
rect 7487 6106 7493 6125
rect 7527 6091 7579 6125
rect 7521 6072 7613 6091
rect 2324 5996 2334 6030
rect 2319 5962 2334 5996
rect 2324 5928 2334 5962
rect 2319 5894 2334 5928
rect 2324 5860 2334 5894
rect 2319 5847 2334 5860
rect 7487 6053 7613 6072
rect 7487 6038 7493 6053
rect 7527 6019 7579 6053
rect 7521 6004 7613 6019
rect 7487 5981 7613 6004
rect 7487 5970 7493 5981
rect 7527 5947 7579 5981
rect 7521 5936 7613 5947
rect 7487 5909 7613 5936
rect 7487 5902 7493 5909
rect 7527 5875 7579 5909
rect 7521 5868 7613 5875
rect 7487 5847 7613 5868
rect 2319 5841 7613 5847
rect 2319 5826 2358 5841
rect 2324 5807 2358 5826
rect 2397 5807 2427 5841
rect 2470 5807 2496 5841
rect 2543 5807 2565 5841
rect 2616 5807 2634 5841
rect 2689 5807 2703 5841
rect 2762 5807 2772 5841
rect 2835 5807 2841 5841
rect 2908 5807 2910 5841
rect 2944 5807 2947 5841
rect 3013 5807 3020 5841
rect 3082 5807 3093 5841
rect 3151 5807 3166 5841
rect 3220 5807 3239 5841
rect 3289 5807 3312 5841
rect 3358 5807 3385 5841
rect 3427 5807 3458 5841
rect 3496 5807 3531 5841
rect 3565 5807 3600 5841
rect 3638 5807 3669 5841
rect 3711 5807 3737 5841
rect 3784 5807 3805 5841
rect 3857 5807 3873 5841
rect 3930 5807 3941 5841
rect 4003 5807 4009 5841
rect 4076 5807 4077 5841
rect 4111 5807 4115 5841
rect 4179 5807 4188 5841
rect 4247 5807 4261 5841
rect 4315 5807 4334 5841
rect 4383 5807 4407 5841
rect 4451 5807 4480 5841
rect 4519 5807 4553 5841
rect 4587 5807 4621 5841
rect 4660 5807 4689 5841
rect 4733 5807 4757 5841
rect 4806 5807 4825 5841
rect 4879 5807 4893 5841
rect 4952 5807 4961 5841
rect 5025 5807 5029 5841
rect 5063 5807 5064 5841
rect 5131 5807 5137 5841
rect 5199 5807 5210 5841
rect 5267 5807 5283 5841
rect 5335 5807 5356 5841
rect 5403 5807 5429 5841
rect 5471 5807 5502 5841
rect 5539 5807 5573 5841
rect 5609 5807 5641 5841
rect 5682 5807 5709 5841
rect 5755 5807 5777 5841
rect 5828 5807 5845 5841
rect 5901 5807 5913 5841
rect 5974 5807 5981 5841
rect 6047 5807 6049 5841
rect 6083 5807 6086 5841
rect 6151 5807 6159 5841
rect 6219 5807 6232 5841
rect 6287 5807 6305 5841
rect 6355 5807 6378 5841
rect 6423 5807 6451 5841
rect 6491 5807 6524 5841
rect 6559 5807 6593 5841
rect 6631 5807 6661 5841
rect 6704 5807 6729 5841
rect 6777 5807 6797 5841
rect 6850 5807 6865 5841
rect 6923 5807 6933 5841
rect 6996 5807 7001 5841
rect 7103 5807 7108 5841
rect 7171 5807 7181 5841
rect 7239 5807 7253 5841
rect 7307 5807 7325 5841
rect 7375 5807 7397 5841
rect 7443 5837 7613 5841
rect 7443 5834 7493 5837
rect 7443 5807 7487 5834
rect 2324 5801 7487 5807
rect 7527 5803 7579 5837
rect 2324 5792 2334 5801
rect 2319 5758 2334 5792
rect 2324 5724 2334 5758
rect 2319 5690 2334 5724
rect 2324 5656 2334 5690
rect 2319 5622 2334 5656
rect 7521 5800 7613 5803
rect 7487 5766 7613 5800
rect 7521 5765 7613 5766
rect 7487 5731 7493 5732
rect 7527 5731 7579 5765
rect 7487 5698 7613 5731
rect 7521 5693 7613 5698
rect 7487 5659 7493 5664
rect 7527 5659 7579 5693
rect 2324 5588 2334 5622
rect 2694 5611 2713 5645
rect 2762 5611 2786 5645
rect 2830 5611 2859 5645
rect 2898 5611 2932 5645
rect 2966 5611 3000 5645
rect 3039 5611 3068 5645
rect 3112 5611 3136 5645
rect 3185 5611 3204 5645
rect 3258 5611 3272 5645
rect 3331 5611 3340 5645
rect 3404 5611 3408 5645
rect 3442 5611 3443 5645
rect 3510 5611 3516 5645
rect 3578 5611 3589 5645
rect 3646 5611 3662 5645
rect 3714 5611 3735 5645
rect 3782 5611 3808 5645
rect 3850 5611 3881 5645
rect 3918 5611 3952 5645
rect 3988 5611 4020 5645
rect 4061 5611 4088 5645
rect 4134 5611 4156 5645
rect 4207 5611 4224 5645
rect 4280 5611 4292 5645
rect 4353 5611 4360 5645
rect 4426 5611 4428 5645
rect 4462 5611 4465 5645
rect 4530 5611 4538 5645
rect 4598 5611 4611 5645
rect 4666 5611 4684 5645
rect 4734 5611 4757 5645
rect 4802 5611 4830 5645
rect 4870 5611 4903 5645
rect 4938 5611 4972 5645
rect 5010 5611 5040 5645
rect 5083 5611 5108 5645
rect 5156 5611 5176 5645
rect 5229 5611 5244 5645
rect 5302 5611 5312 5645
rect 5375 5611 5380 5645
rect 5482 5611 5487 5645
rect 5550 5611 5560 5645
rect 5618 5611 5633 5645
rect 5686 5611 5706 5645
rect 5754 5611 5778 5645
rect 5822 5611 5850 5645
rect 5890 5611 5922 5645
rect 5958 5611 5992 5645
rect 6028 5611 6060 5645
rect 6100 5611 6128 5645
rect 6172 5611 6196 5645
rect 6244 5611 6264 5645
rect 6316 5611 6332 5645
rect 6388 5611 6400 5645
rect 6460 5611 6468 5645
rect 6532 5611 6536 5645
rect 6638 5611 6642 5645
rect 6706 5611 6714 5645
rect 6774 5611 6786 5645
rect 6842 5611 6858 5645
rect 6910 5611 6930 5645
rect 6978 5611 7002 5645
rect 7036 5611 7048 5645
rect 7487 5630 7613 5659
rect 7521 5621 7613 5630
rect 2319 5554 2334 5588
rect 2324 5520 2334 5554
rect 7487 5587 7493 5596
rect 7527 5587 7579 5621
rect 7487 5562 7613 5587
rect 7521 5549 7613 5562
rect 2319 5486 2334 5520
rect 2324 5452 2334 5486
rect 2319 5418 2334 5452
rect 2324 5384 2334 5418
rect 2319 5350 2334 5384
rect 2324 5316 2334 5350
rect 2687 5472 2721 5512
rect 2687 5398 2721 5438
rect 2687 5324 2721 5364
rect 2319 5305 2334 5316
rect 2141 5282 2334 5305
rect 2141 5266 2290 5282
rect 2175 5232 2213 5266
rect 2247 5232 2285 5266
rect 2324 5248 2334 5282
rect 2319 5232 2334 5248
rect 2141 5214 2334 5232
rect 2141 5193 2290 5214
rect 2175 5159 2213 5193
rect 2247 5159 2285 5193
rect 2324 5180 2334 5214
rect 2319 5159 2334 5180
rect 2141 5146 2334 5159
rect 2141 5120 2290 5146
rect 2175 5086 2213 5120
rect 2247 5086 2285 5120
rect 2324 5112 2334 5146
rect 2319 5086 2334 5112
rect 2141 5078 2334 5086
rect 2141 5047 2290 5078
rect 2175 5013 2213 5047
rect 2247 5013 2285 5047
rect 2324 5044 2334 5078
rect 2319 5013 2334 5044
rect 2141 5010 2334 5013
rect 2141 4976 2290 5010
rect 2324 4976 2334 5010
rect 2141 4974 2334 4976
rect 2175 4940 2213 4974
rect 2247 4940 2285 4974
rect 2319 4942 2334 4974
rect 2141 4908 2290 4940
rect 2324 4908 2334 4942
rect 2141 4901 2334 4908
rect 2175 4867 2213 4901
rect 2247 4867 2285 4901
rect 2319 4874 2334 4901
rect 2141 4840 2290 4867
rect 2324 4840 2334 4874
rect 2141 4828 2334 4840
rect 2175 4794 2213 4828
rect 2247 4794 2285 4828
rect 2319 4806 2334 4828
rect 2141 4772 2290 4794
rect 2324 4772 2334 4806
rect 2141 4755 2334 4772
rect 2175 4721 2213 4755
rect 2247 4721 2285 4755
rect 2319 4738 2334 4755
rect 2141 4704 2290 4721
rect 2324 4704 2334 4738
rect 2141 4682 2334 4704
rect 2175 4648 2213 4682
rect 2247 4648 2285 4682
rect 2319 4670 2334 4682
rect 2141 4636 2290 4648
rect 2324 4636 2334 4670
rect 2141 4609 2334 4636
rect 2175 4575 2213 4609
rect 2247 4575 2285 4609
rect 2319 4602 2334 4609
rect 2141 4568 2290 4575
rect 2324 4568 2334 4602
rect 2141 4536 2334 4568
rect 2175 4502 2213 4536
rect 2247 4502 2285 4536
rect 2319 4534 2334 4536
rect 2141 4500 2290 4502
rect 2324 4500 2334 4534
rect 2141 4466 2334 4500
rect 2141 4463 2290 4466
rect 2175 4429 2213 4463
rect 2247 4429 2285 4463
rect 2324 4432 2334 4466
rect 2319 4429 2334 4432
rect 2141 4398 2334 4429
rect 2141 4390 2290 4398
rect 2175 4356 2213 4390
rect 2247 4356 2285 4390
rect 2324 4364 2334 4398
rect 2319 4356 2334 4364
rect 2141 4330 2334 4356
rect 2141 4317 2290 4330
rect 2175 4283 2213 4317
rect 2247 4283 2285 4317
rect 2324 4296 2334 4330
rect 2319 4283 2334 4296
rect 2141 4262 2334 4283
rect 2141 4244 2290 4262
rect 2175 4210 2213 4244
rect 2247 4210 2285 4244
rect 2324 4228 2334 4262
rect 2319 4210 2334 4228
rect 2141 4194 2334 4210
rect 2141 4171 2290 4194
rect 2175 4137 2213 4171
rect 2247 4137 2285 4171
rect 2324 4160 2334 4194
rect 2595 5245 2629 5285
rect 2595 5171 2629 5211
rect 2595 5097 2629 5137
rect 2595 5023 2629 5063
rect 2595 4949 2629 4989
rect 2595 4875 2629 4915
rect 2595 4801 2629 4841
rect 2595 4727 2629 4767
rect 2595 4653 2629 4693
rect 2595 4579 2629 4619
rect 2595 4504 2629 4545
rect 2595 4429 2629 4470
rect 2595 4354 2629 4395
rect 2595 4279 2629 4320
rect 2595 4204 2629 4245
rect 7487 5515 7493 5528
rect 7527 5515 7579 5549
rect 7487 5494 7613 5515
rect 7521 5477 7613 5494
rect 7487 5443 7493 5460
rect 7527 5443 7579 5477
rect 7487 5426 7613 5443
rect 7521 5405 7613 5426
rect 7487 5371 7493 5392
rect 7527 5371 7579 5405
rect 7487 5358 7613 5371
rect 7521 5333 7613 5358
rect 2687 5250 2721 5290
rect 2687 5176 2721 5216
rect 2687 5102 2721 5142
rect 2687 5028 2721 5068
rect 2687 4954 2721 4994
rect 2687 4879 2721 4920
rect 2687 4804 2721 4845
rect 2687 4729 2721 4770
rect 2687 4654 2721 4695
rect 2687 4579 2721 4620
rect 2687 4504 2721 4545
rect 2687 4429 2721 4470
rect 2687 4354 2721 4395
rect 2687 4279 2721 4320
rect 2687 4204 2721 4245
rect 2779 5245 2813 5285
rect 2779 5171 2813 5211
rect 2779 5097 2813 5137
rect 2779 5023 2813 5063
rect 2779 4949 2813 4989
rect 2779 4875 2813 4915
rect 2779 4801 2813 4841
rect 2779 4727 2813 4767
rect 2779 4653 2813 4693
rect 2779 4579 2813 4619
rect 2779 4504 2813 4545
rect 2779 4429 2813 4470
rect 2779 4354 2813 4395
rect 2779 4279 2813 4320
rect 2779 4204 2813 4245
rect 3627 5285 3632 5319
rect 3666 5285 3671 5319
rect 3627 5244 3671 5285
rect 3627 5210 3632 5244
rect 3666 5210 3671 5244
rect 3627 5169 3671 5210
rect 3627 5135 3632 5169
rect 3666 5135 3671 5169
rect 3627 5094 3671 5135
rect 3627 5060 3632 5094
rect 3666 5060 3671 5094
rect 3627 5019 3671 5060
rect 3627 4985 3632 5019
rect 3666 4985 3671 5019
rect 3627 4944 3671 4985
rect 3627 4910 3632 4944
rect 3666 4910 3671 4944
rect 3627 4869 3671 4910
rect 3627 4835 3632 4869
rect 3666 4835 3671 4869
rect 3627 4794 3671 4835
rect 3627 4760 3632 4794
rect 3666 4760 3671 4794
rect 3627 4719 3671 4760
rect 3627 4685 3632 4719
rect 3666 4685 3671 4719
rect 3627 4644 3671 4685
rect 3627 4610 3632 4644
rect 3666 4610 3671 4644
rect 3627 4569 3671 4610
rect 3627 4535 3632 4569
rect 3666 4535 3671 4569
rect 3627 4494 3671 4535
rect 3627 4460 3632 4494
rect 3666 4460 3671 4494
rect 3627 4419 3671 4460
rect 3627 4385 3632 4419
rect 3666 4385 3671 4419
rect 3627 4344 3671 4385
rect 3627 4310 3632 4344
rect 3666 4310 3671 4344
rect 3627 4269 3671 4310
rect 3627 4235 3632 4269
rect 3666 4235 3671 4269
rect 3627 4193 3671 4235
rect 2319 4137 2334 4160
rect 3627 4159 3632 4193
rect 3666 4159 3671 4193
rect 4486 5285 4491 5319
rect 4525 5285 4530 5319
rect 4486 5244 4530 5285
rect 4486 5210 4491 5244
rect 4525 5210 4530 5244
rect 4486 5169 4530 5210
rect 4486 5135 4491 5169
rect 4525 5135 4530 5169
rect 4486 5094 4530 5135
rect 4486 5060 4491 5094
rect 4525 5060 4530 5094
rect 4486 5019 4530 5060
rect 4486 4985 4491 5019
rect 4525 4985 4530 5019
rect 4486 4944 4530 4985
rect 4486 4910 4491 4944
rect 4525 4910 4530 4944
rect 4486 4869 4530 4910
rect 4486 4835 4491 4869
rect 4525 4835 4530 4869
rect 4486 4794 4530 4835
rect 4486 4760 4491 4794
rect 4525 4760 4530 4794
rect 4486 4719 4530 4760
rect 4486 4685 4491 4719
rect 4525 4685 4530 4719
rect 4486 4644 4530 4685
rect 4486 4610 4491 4644
rect 4525 4610 4530 4644
rect 4486 4569 4530 4610
rect 4486 4535 4491 4569
rect 4525 4535 4530 4569
rect 4486 4494 4530 4535
rect 4486 4460 4491 4494
rect 4525 4460 4530 4494
rect 4486 4419 4530 4460
rect 4486 4385 4491 4419
rect 4525 4385 4530 4419
rect 4486 4344 4530 4385
rect 4486 4310 4491 4344
rect 4525 4310 4530 4344
rect 4486 4269 4530 4310
rect 4486 4235 4491 4269
rect 4525 4235 4530 4269
rect 4486 4193 4530 4235
rect 4486 4159 4491 4193
rect 4525 4159 4530 4193
rect 5342 5285 5347 5319
rect 5381 5285 5386 5319
rect 5342 5244 5386 5285
rect 5342 5210 5347 5244
rect 5381 5210 5386 5244
rect 5342 5169 5386 5210
rect 5342 5135 5347 5169
rect 5381 5135 5386 5169
rect 5342 5094 5386 5135
rect 5342 5060 5347 5094
rect 5381 5060 5386 5094
rect 5342 5019 5386 5060
rect 5342 4985 5347 5019
rect 5381 4985 5386 5019
rect 5342 4944 5386 4985
rect 5342 4910 5347 4944
rect 5381 4910 5386 4944
rect 5342 4869 5386 4910
rect 5342 4835 5347 4869
rect 5381 4835 5386 4869
rect 5342 4794 5386 4835
rect 5342 4760 5347 4794
rect 5381 4760 5386 4794
rect 5342 4719 5386 4760
rect 5342 4685 5347 4719
rect 5381 4685 5386 4719
rect 5342 4644 5386 4685
rect 5342 4610 5347 4644
rect 5381 4610 5386 4644
rect 5342 4569 5386 4610
rect 5342 4535 5347 4569
rect 5381 4535 5386 4569
rect 5342 4494 5386 4535
rect 5342 4460 5347 4494
rect 5381 4460 5386 4494
rect 5342 4419 5386 4460
rect 5342 4385 5347 4419
rect 5381 4385 5386 4419
rect 5342 4344 5386 4385
rect 5342 4310 5347 4344
rect 5381 4310 5386 4344
rect 5342 4269 5386 4310
rect 5342 4235 5347 4269
rect 5381 4235 5386 4269
rect 5342 4193 5386 4235
rect 5342 4159 5347 4193
rect 5381 4159 5386 4193
rect 6201 5285 6206 5319
rect 6240 5285 6245 5319
rect 6201 5244 6245 5285
rect 6201 5210 6206 5244
rect 6240 5210 6245 5244
rect 6201 5169 6245 5210
rect 6201 5135 6206 5169
rect 6240 5135 6245 5169
rect 6201 5094 6245 5135
rect 6201 5060 6206 5094
rect 6240 5060 6245 5094
rect 6201 5019 6245 5060
rect 6201 4985 6206 5019
rect 6240 4985 6245 5019
rect 6201 4944 6245 4985
rect 6201 4910 6206 4944
rect 6240 4910 6245 4944
rect 6201 4869 6245 4910
rect 6201 4835 6206 4869
rect 6240 4835 6245 4869
rect 6201 4794 6245 4835
rect 6201 4760 6206 4794
rect 6240 4760 6245 4794
rect 6201 4719 6245 4760
rect 6201 4685 6206 4719
rect 6240 4685 6245 4719
rect 6201 4644 6245 4685
rect 6201 4610 6206 4644
rect 6240 4610 6245 4644
rect 6201 4569 6245 4610
rect 6201 4535 6206 4569
rect 6240 4535 6245 4569
rect 6201 4494 6245 4535
rect 6201 4460 6206 4494
rect 6240 4460 6245 4494
rect 6201 4419 6245 4460
rect 6201 4385 6206 4419
rect 6240 4385 6245 4419
rect 6201 4344 6245 4385
rect 6201 4310 6206 4344
rect 6240 4310 6245 4344
rect 6201 4269 6245 4310
rect 6201 4235 6206 4269
rect 6240 4235 6245 4269
rect 6201 4193 6245 4235
rect 6201 4159 6206 4193
rect 6240 4159 6245 4193
rect 7054 5285 7059 5319
rect 7093 5285 7098 5319
rect 7054 5244 7098 5285
rect 7054 5210 7059 5244
rect 7093 5210 7098 5244
rect 7054 5169 7098 5210
rect 7054 5135 7059 5169
rect 7093 5135 7098 5169
rect 7054 5094 7098 5135
rect 7054 5060 7059 5094
rect 7093 5060 7098 5094
rect 7054 5019 7098 5060
rect 7054 4985 7059 5019
rect 7093 4985 7098 5019
rect 7054 4944 7098 4985
rect 7054 4910 7059 4944
rect 7093 4910 7098 4944
rect 7054 4869 7098 4910
rect 7054 4835 7059 4869
rect 7093 4835 7098 4869
rect 7054 4794 7098 4835
rect 7054 4760 7059 4794
rect 7093 4760 7098 4794
rect 7054 4719 7098 4760
rect 7054 4685 7059 4719
rect 7093 4685 7098 4719
rect 7054 4644 7098 4685
rect 7054 4610 7059 4644
rect 7093 4610 7098 4644
rect 7054 4569 7098 4610
rect 7054 4535 7059 4569
rect 7093 4535 7098 4569
rect 7054 4494 7098 4535
rect 7054 4460 7059 4494
rect 7093 4460 7098 4494
rect 7054 4419 7098 4460
rect 7054 4385 7059 4419
rect 7093 4385 7098 4419
rect 7054 4344 7098 4385
rect 7054 4310 7059 4344
rect 7093 4310 7098 4344
rect 7054 4269 7098 4310
rect 7054 4235 7059 4269
rect 7093 4235 7098 4269
rect 7054 4193 7098 4235
rect 7054 4159 7059 4193
rect 7093 4159 7098 4193
rect 7487 5299 7493 5324
rect 7527 5299 7579 5333
rect 7487 5290 7613 5299
rect 7521 5261 7613 5290
rect 7487 5227 7493 5256
rect 7527 5227 7579 5261
rect 7487 5222 7613 5227
rect 7521 5189 7613 5222
rect 7487 5155 7493 5188
rect 7527 5155 7579 5189
rect 7487 5154 7613 5155
rect 7521 5120 7613 5154
rect 7487 5117 7613 5120
rect 7487 5086 7493 5117
rect 7527 5083 7579 5117
rect 7521 5052 7613 5083
rect 7487 5045 7613 5052
rect 7487 5018 7493 5045
rect 7527 5011 7579 5045
rect 7521 4984 7613 5011
rect 7487 4973 7613 4984
rect 7487 4950 7493 4973
rect 7527 4939 7579 4973
rect 7521 4916 7613 4939
rect 7487 4901 7613 4916
rect 7487 4882 7493 4901
rect 7527 4867 7579 4901
rect 7521 4848 7613 4867
rect 7487 4829 7613 4848
rect 7487 4814 7493 4829
rect 7527 4795 7579 4829
rect 7521 4780 7613 4795
rect 7487 4757 7613 4780
rect 7487 4746 7493 4757
rect 7527 4723 7579 4757
rect 7521 4712 7613 4723
rect 7487 4685 7613 4712
rect 7487 4678 7493 4685
rect 7527 4651 7579 4685
rect 7521 4644 7613 4651
rect 7487 4613 7613 4644
rect 7487 4610 7493 4613
rect 7527 4579 7579 4613
rect 7521 4576 7613 4579
rect 7487 4542 7613 4576
rect 7521 4540 7613 4542
rect 7487 4506 7493 4508
rect 7527 4506 7579 4540
rect 7487 4474 7613 4506
rect 7521 4467 7613 4474
rect 7487 4433 7493 4440
rect 7527 4433 7579 4467
rect 7487 4406 7613 4433
rect 7521 4394 7613 4406
rect 7487 4360 7493 4372
rect 7527 4360 7579 4394
rect 7487 4338 7613 4360
rect 7521 4321 7613 4338
rect 7487 4287 7493 4304
rect 7527 4287 7579 4321
rect 7487 4270 7613 4287
rect 7521 4248 7613 4270
rect 7487 4214 7493 4236
rect 7527 4214 7579 4248
rect 7487 4202 7613 4214
rect 7521 4175 7613 4202
rect 2141 4126 2334 4137
rect 2141 4098 2290 4126
rect 2175 4064 2213 4098
rect 2247 4064 2285 4098
rect 2324 4092 2334 4126
rect 2319 4064 2334 4092
rect 2141 4058 2334 4064
rect 2141 4025 2290 4058
rect 2175 3991 2213 4025
rect 2247 3991 2285 4025
rect 2324 4024 2334 4058
rect 2319 3991 2334 4024
rect 2141 3943 2334 3991
rect 7487 4141 7493 4168
rect 7527 4141 7579 4175
rect 7487 4134 7613 4141
rect 7521 4102 7613 4134
rect 7487 4068 7493 4100
rect 7527 4068 7579 4102
rect 7487 4066 7613 4068
rect 7521 4032 7613 4066
rect 7487 4029 7613 4032
rect 7487 3998 7493 4029
rect 7527 3995 7579 4029
rect 7521 3964 7613 3995
rect 7487 3943 7613 3964
rect 2141 3909 2147 3943
rect 2181 3909 2220 3943
rect 2254 3909 2293 3943
rect 2327 3909 2366 3943
rect 2400 3909 2439 3943
rect 2473 3909 2512 3943
rect 2546 3909 2585 3943
rect 2619 3909 2658 3943
rect 2692 3909 2731 3943
rect 2765 3909 2804 3943
rect 2838 3909 2877 3943
rect 2911 3909 2950 3943
rect 2984 3909 3023 3943
rect 2141 3907 3023 3909
rect 2141 3873 2314 3907
rect 2348 3873 2382 3907
rect 2416 3873 2450 3907
rect 2484 3873 2518 3907
rect 2552 3873 2586 3907
rect 2620 3873 2654 3907
rect 2688 3873 2722 3907
rect 2756 3873 2790 3907
rect 2824 3873 2858 3907
rect 2892 3873 2926 3907
rect 2960 3873 2994 3907
rect 2141 3871 3023 3873
rect 2141 3837 2147 3871
rect 2181 3837 2220 3871
rect 2254 3837 2293 3871
rect 2327 3837 2366 3871
rect 2400 3837 2439 3871
rect 2473 3837 2512 3871
rect 2546 3837 2585 3871
rect 2619 3837 2658 3871
rect 2692 3837 2731 3871
rect 2765 3837 2804 3871
rect 2838 3837 2877 3871
rect 2911 3837 2950 3871
rect 2984 3837 3023 3871
rect 7593 3837 7613 3943
rect 7733 4489 7735 4528
rect 7837 4489 7839 4528
rect 7733 4416 7735 4455
rect 7837 4416 7839 4455
rect 7733 4343 7735 4382
rect 7837 4343 7839 4382
rect 7733 4270 7735 4309
rect 7837 4270 7839 4309
rect 7733 4197 7735 4236
rect 7837 4197 7839 4236
rect 7767 4163 7805 4175
rect 7733 4124 7839 4163
rect 7767 4090 7805 4124
rect 7733 4063 7839 4090
rect 7733 4051 7735 4063
rect 7837 4051 7839 4063
rect 7733 3978 7735 4017
rect 7837 3978 7839 4017
rect 7733 3905 7735 3944
rect 7837 3905 7839 3944
rect 1938 3459 1946 3491
rect 2048 3453 2056 3491
rect 7733 3832 7735 3871
rect 7837 3832 7839 3871
rect 7733 3759 7735 3798
rect 7837 3759 7839 3798
rect 7733 3686 7735 3725
rect 7837 3686 7839 3725
rect 7733 3613 7735 3652
rect 7837 3613 7839 3652
rect 7733 3540 7735 3579
rect 7837 3540 7839 3579
rect 7733 3467 7735 3506
rect 7837 3467 7839 3506
rect 2057 3451 2096 3453
rect 2130 3451 2169 3453
rect 2203 3451 2242 3453
rect 2276 3451 2315 3453
rect 2349 3451 2388 3453
rect 2422 3451 2461 3453
rect 2495 3451 2534 3453
rect 2568 3451 2607 3453
rect 2057 3419 2088 3451
rect 2598 3419 2607 3451
rect 2641 3451 2680 3453
rect 2714 3451 2753 3453
rect 2787 3451 2826 3453
rect 2860 3451 2899 3453
rect 2933 3451 2972 3453
rect 3006 3451 3045 3453
rect 3079 3451 3118 3453
rect 3152 3451 3191 3453
rect 3225 3451 3264 3453
rect 3298 3451 3337 3453
rect 3371 3451 3410 3453
rect 3444 3451 3483 3453
rect 3517 3451 3556 3453
rect 3590 3451 3629 3453
rect 3663 3451 3702 3453
rect 3736 3451 3775 3453
rect 3809 3451 3848 3453
rect 3882 3451 3921 3453
rect 3955 3451 3994 3453
rect 4028 3451 4067 3453
rect 4101 3451 4140 3453
rect 4174 3451 4213 3453
rect 4247 3451 4286 3453
rect 4320 3451 4359 3453
rect 4393 3451 4432 3453
rect 4466 3451 4505 3453
rect 4539 3451 4578 3453
rect 4612 3451 4651 3453
rect 4685 3451 4724 3453
rect 4758 3451 4797 3453
rect 4831 3451 4870 3453
rect 4904 3451 4943 3453
rect 4977 3451 5016 3453
rect 5050 3451 5089 3453
rect 5123 3451 5162 3453
rect 5196 3451 5235 3453
rect 5269 3451 5308 3453
rect 5342 3451 5381 3453
rect 5415 3451 5454 3453
rect 5488 3451 5527 3453
rect 5561 3451 5600 3453
rect 5634 3451 5673 3453
rect 5707 3451 5746 3453
rect 5780 3451 5819 3453
rect 5853 3451 5892 3453
rect 5926 3451 5965 3453
rect 5999 3451 6038 3453
rect 6072 3451 6111 3453
rect 6145 3451 6184 3453
rect 6218 3451 6257 3453
rect 6291 3451 6330 3453
rect 7660 3451 7733 3453
rect 2641 3419 2666 3451
rect 2048 3417 2088 3419
rect 1946 3383 2088 3417
rect 1946 3381 2020 3383
rect 2054 3381 2088 3383
rect 2598 3381 2666 3419
rect 1946 3347 1950 3381
rect 1984 3349 2020 3381
rect 2057 3349 2088 3381
rect 2598 3349 2607 3381
rect 1984 3347 2023 3349
rect 2057 3347 2096 3349
rect 2130 3347 2169 3349
rect 2203 3347 2242 3349
rect 2276 3347 2315 3349
rect 2349 3347 2388 3349
rect 2422 3347 2461 3349
rect 2495 3347 2534 3349
rect 2568 3347 2607 3349
rect 2641 3349 2666 3381
rect 7677 3433 7733 3451
rect 7677 3417 7735 3433
rect 7837 3417 7839 3433
rect 7677 3394 7839 3417
rect 7677 3383 7733 3394
rect 7677 3349 7711 3383
rect 7767 3360 7805 3394
rect 7745 3349 7839 3360
rect 2641 3347 2680 3349
rect 2714 3347 2753 3349
rect 2787 3347 2826 3349
rect 2860 3347 2899 3349
rect 2933 3347 2972 3349
rect 3006 3347 3045 3349
rect 3079 3347 3118 3349
rect 3152 3347 3191 3349
rect 3225 3347 3264 3349
rect 3298 3347 3337 3349
rect 3371 3347 3410 3349
rect 3444 3347 3483 3349
rect 3517 3347 3556 3349
rect 3590 3347 3629 3349
rect 3663 3347 3702 3349
rect 3736 3347 3775 3349
rect 3809 3347 3848 3349
rect 3882 3347 3921 3349
rect 3955 3347 3994 3349
rect 4028 3347 4067 3349
rect 4101 3347 4140 3349
rect 4174 3347 4213 3349
rect 4247 3347 4286 3349
rect 4320 3347 4359 3349
rect 4393 3347 4432 3349
rect 4466 3347 4505 3349
rect 4539 3347 4578 3349
rect 4612 3347 4651 3349
rect 4685 3347 4724 3349
rect 4758 3347 4797 3349
rect 4831 3347 4870 3349
rect 4904 3347 4943 3349
rect 4977 3347 5016 3349
rect 5050 3347 5089 3349
rect 5123 3347 5162 3349
rect 5196 3347 5235 3349
rect 5269 3347 5308 3349
rect 5342 3347 5381 3349
rect 5415 3347 5454 3349
rect 5488 3347 5527 3349
rect 5561 3347 5600 3349
rect 5634 3347 5673 3349
rect 5707 3347 5746 3349
rect 5780 3347 5819 3349
rect 5853 3347 5892 3349
rect 5926 3347 5965 3349
rect 5999 3347 6038 3349
rect 6072 3347 6111 3349
rect 6145 3347 6184 3349
rect 6218 3347 6257 3349
rect 6291 3347 6330 3349
rect 7660 3347 7839 3349
rect 1831 3126 7904 3127
rect 1831 3092 1855 3126
rect 1889 3092 1992 3126
rect 2026 3092 2129 3126
rect 2163 3092 2266 3126
rect 2300 3092 2403 3126
rect 2437 3092 2540 3126
rect 2574 3092 2677 3126
rect 2711 3092 2814 3126
rect 2848 3092 2950 3126
rect 2984 3092 3086 3126
rect 3120 3092 3222 3126
rect 3256 3092 3358 3126
rect 3392 3092 3494 3126
rect 3528 3092 3630 3126
rect 3664 3092 3766 3126
rect 3800 3092 3902 3126
rect 3936 3092 4038 3126
rect 4072 3092 4174 3126
rect 4208 3092 4310 3126
rect 4344 3092 4446 3126
rect 4480 3092 4582 3126
rect 4616 3092 4718 3126
rect 4752 3092 4854 3126
rect 4888 3092 4990 3126
rect 5024 3092 5126 3126
rect 5160 3092 5262 3126
rect 5296 3092 5398 3126
rect 5432 3092 5534 3126
rect 5568 3092 5670 3126
rect 5704 3092 5806 3126
rect 5840 3092 5942 3126
rect 5976 3092 6078 3126
rect 6112 3092 6214 3126
rect 6248 3092 6350 3126
rect 6384 3092 6486 3126
rect 6520 3092 6622 3126
rect 6656 3092 6758 3126
rect 6792 3092 6894 3126
rect 6928 3092 7030 3126
rect 7064 3092 7166 3126
rect 7200 3092 7302 3126
rect 7336 3092 7438 3126
rect 7472 3092 7574 3126
rect 7608 3092 7710 3126
rect 7744 3092 7846 3126
rect 7880 3092 7904 3126
rect 1831 3049 7904 3092
rect 1831 3015 1935 3049
rect 1969 3015 2008 3049
rect 2042 3015 2081 3049
rect 2115 3015 2154 3049
rect 2188 3015 2227 3049
rect 2261 3015 2300 3049
rect 2334 3015 2373 3049
rect 2407 3015 2446 3049
rect 2480 3015 2519 3049
rect 2553 3015 2592 3049
rect 2626 3015 2665 3049
rect 2699 3015 2738 3049
rect 2772 3015 2811 3049
rect 2845 3015 2884 3049
rect 2918 3015 2957 3049
rect 2991 3015 3030 3049
rect 3064 3015 3103 3049
rect 3137 3015 3176 3049
rect 3210 3015 3249 3049
rect 3283 3015 3322 3049
rect 3356 3015 3395 3049
rect 3429 3015 3468 3049
rect 3502 3015 3541 3049
rect 3575 3015 3614 3049
rect 3648 3015 3687 3049
rect 3721 3015 3760 3049
rect 3794 3015 3833 3049
rect 3867 3015 3906 3049
rect 3940 3015 3979 3049
rect 4013 3015 4052 3049
rect 4086 3015 4125 3049
rect 4159 3015 4198 3049
rect 4232 3015 4271 3049
rect 4305 3015 4344 3049
rect 4378 3015 4417 3049
rect 4451 3015 4490 3049
rect 4524 3015 4563 3049
rect 4597 3015 4636 3049
rect 4670 3015 4709 3049
rect 4743 3015 4782 3049
rect 4816 3015 4855 3049
rect 4889 3015 4928 3049
rect 4962 3015 5001 3049
rect 5035 3015 5074 3049
rect 5108 3015 5147 3049
rect 5181 3015 5220 3049
rect 5254 3015 5293 3049
rect 5327 3015 5366 3049
rect 5400 3015 5439 3049
rect 5473 3015 5511 3049
rect 5545 3015 5583 3049
rect 5617 3015 5655 3049
rect 5689 3015 5727 3049
rect 5761 3015 5799 3049
rect 5833 3015 5871 3049
rect 5905 3015 5943 3049
rect 5977 3015 6015 3049
rect 6049 3015 6087 3049
rect 6121 3015 6159 3049
rect 6193 3015 6231 3049
rect 6265 3015 6303 3049
rect 6337 3015 6375 3049
rect 6409 3015 6447 3049
rect 6481 3015 6519 3049
rect 6553 3015 6591 3049
rect 6625 3015 6663 3049
rect 6697 3015 6735 3049
rect 6769 3015 6807 3049
rect 6841 3015 6879 3049
rect 6913 3015 6951 3049
rect 6985 3015 7023 3049
rect 7057 3015 7095 3049
rect 7129 3015 7167 3049
rect 7201 3015 7239 3049
rect 7273 3015 7311 3049
rect 7345 3015 7383 3049
rect 7417 3015 7455 3049
rect 7489 3015 7527 3049
rect 7561 3015 7904 3049
rect 1831 3010 7904 3015
rect 1831 2976 1855 3010
rect 1889 2976 1992 3010
rect 2026 2976 2129 3010
rect 2163 2976 2266 3010
rect 2300 2976 2403 3010
rect 2437 2976 2540 3010
rect 2574 2976 2677 3010
rect 2711 2976 2814 3010
rect 2848 2976 2950 3010
rect 2984 2976 3086 3010
rect 3120 2976 3222 3010
rect 3256 2976 3358 3010
rect 3392 2976 3494 3010
rect 3528 2976 3630 3010
rect 3664 2976 3766 3010
rect 3800 2976 3902 3010
rect 3936 2976 4038 3010
rect 4072 2976 4174 3010
rect 4208 2976 4310 3010
rect 4344 2976 4446 3010
rect 4480 2976 4582 3010
rect 4616 2976 4718 3010
rect 4752 2976 4854 3010
rect 4888 2976 4990 3010
rect 5024 2976 5126 3010
rect 5160 2976 5262 3010
rect 5296 2976 5398 3010
rect 5432 2976 5534 3010
rect 5568 2976 5670 3010
rect 5704 2976 5806 3010
rect 5840 2976 5942 3010
rect 5976 2976 6078 3010
rect 6112 2976 6214 3010
rect 6248 2976 6350 3010
rect 6384 2976 6486 3010
rect 6520 2976 6622 3010
rect 6656 2976 6758 3010
rect 6792 2976 6894 3010
rect 6928 2976 7030 3010
rect 7064 2976 7166 3010
rect 7200 2976 7302 3010
rect 7336 2976 7438 3010
rect 7472 2976 7574 3010
rect 7608 2976 7710 3010
rect 7744 2976 7846 3010
rect 7880 2976 7904 3010
rect 1831 2971 7904 2976
rect 1831 2937 1935 2971
rect 1969 2937 2008 2971
rect 2042 2937 2081 2971
rect 2115 2937 2154 2971
rect 2188 2937 2227 2971
rect 2261 2937 2300 2971
rect 2334 2937 2373 2971
rect 2407 2937 2446 2971
rect 2480 2937 2519 2971
rect 2553 2937 2592 2971
rect 2626 2937 2665 2971
rect 2699 2937 2738 2971
rect 2772 2937 2811 2971
rect 2845 2937 2884 2971
rect 2918 2937 2957 2971
rect 2991 2937 3030 2971
rect 3064 2937 3103 2971
rect 3137 2937 3176 2971
rect 3210 2937 3249 2971
rect 3283 2937 3322 2971
rect 3356 2937 3395 2971
rect 3429 2937 3468 2971
rect 3502 2937 3541 2971
rect 3575 2937 3614 2971
rect 3648 2937 3687 2971
rect 3721 2937 3760 2971
rect 3794 2937 3833 2971
rect 3867 2937 3906 2971
rect 3940 2937 3979 2971
rect 4013 2937 4052 2971
rect 4086 2937 4125 2971
rect 4159 2937 4198 2971
rect 4232 2937 4271 2971
rect 4305 2937 4344 2971
rect 4378 2937 4417 2971
rect 4451 2937 4490 2971
rect 4524 2937 4563 2971
rect 4597 2937 4636 2971
rect 4670 2937 4709 2971
rect 4743 2937 4782 2971
rect 4816 2937 4855 2971
rect 4889 2937 4928 2971
rect 4962 2937 5001 2971
rect 5035 2937 5074 2971
rect 5108 2937 5147 2971
rect 5181 2937 5220 2971
rect 5254 2937 5293 2971
rect 5327 2937 5366 2971
rect 5400 2937 5439 2971
rect 5473 2937 5511 2971
rect 5545 2937 5583 2971
rect 5617 2937 5655 2971
rect 5689 2937 5727 2971
rect 5761 2937 5799 2971
rect 5833 2937 5871 2971
rect 5905 2937 5943 2971
rect 5977 2937 6015 2971
rect 6049 2937 6087 2971
rect 6121 2937 6159 2971
rect 6193 2937 6231 2971
rect 6265 2937 6303 2971
rect 6337 2937 6375 2971
rect 6409 2937 6447 2971
rect 6481 2937 6519 2971
rect 6553 2937 6591 2971
rect 6625 2937 6663 2971
rect 6697 2937 6735 2971
rect 6769 2937 6807 2971
rect 6841 2937 6879 2971
rect 6913 2937 6951 2971
rect 6985 2937 7023 2971
rect 7057 2937 7095 2971
rect 7129 2937 7167 2971
rect 7201 2937 7239 2971
rect 7273 2937 7311 2971
rect 7345 2937 7383 2971
rect 7417 2937 7455 2971
rect 7489 2937 7527 2971
rect 7561 2937 7904 2971
rect 1831 2894 7904 2937
rect 1831 2860 1855 2894
rect 1889 2893 1992 2894
rect 2026 2893 2129 2894
rect 2163 2893 2266 2894
rect 1889 2860 1935 2893
rect 1831 2859 1935 2860
rect 1969 2860 1992 2893
rect 1969 2859 2008 2860
rect 2042 2859 2081 2893
rect 2115 2860 2129 2893
rect 2115 2859 2154 2860
rect 2188 2859 2227 2893
rect 2261 2860 2266 2893
rect 2300 2893 2403 2894
rect 2437 2893 2540 2894
rect 2574 2893 2677 2894
rect 2711 2893 2814 2894
rect 2848 2893 2950 2894
rect 2984 2893 3086 2894
rect 3120 2893 3222 2894
rect 3256 2893 3358 2894
rect 2261 2859 2300 2860
rect 2334 2859 2373 2893
rect 2437 2860 2446 2893
rect 2407 2859 2446 2860
rect 2480 2859 2519 2893
rect 2574 2860 2592 2893
rect 2553 2859 2592 2860
rect 2626 2859 2665 2893
rect 2711 2860 2738 2893
rect 2699 2859 2738 2860
rect 2772 2859 2811 2893
rect 2848 2860 2884 2893
rect 2845 2859 2884 2860
rect 2918 2860 2950 2893
rect 2918 2859 2957 2860
rect 2991 2859 3030 2893
rect 3064 2860 3086 2893
rect 3064 2859 3103 2860
rect 3137 2859 3176 2893
rect 3210 2860 3222 2893
rect 3210 2859 3249 2860
rect 3283 2859 3322 2893
rect 3356 2860 3358 2893
rect 3392 2893 3494 2894
rect 3528 2893 3630 2894
rect 3664 2893 3766 2894
rect 3800 2893 3902 2894
rect 3936 2893 4038 2894
rect 4072 2893 4174 2894
rect 4208 2893 4310 2894
rect 3392 2860 3395 2893
rect 3356 2859 3395 2860
rect 3429 2859 3468 2893
rect 3528 2860 3541 2893
rect 3502 2859 3541 2860
rect 3575 2859 3614 2893
rect 3664 2860 3687 2893
rect 3648 2859 3687 2860
rect 3721 2859 3760 2893
rect 3800 2860 3833 2893
rect 3794 2859 3833 2860
rect 3867 2860 3902 2893
rect 3867 2859 3906 2860
rect 3940 2859 3979 2893
rect 4013 2860 4038 2893
rect 4013 2859 4052 2860
rect 4086 2859 4125 2893
rect 4159 2860 4174 2893
rect 4159 2859 4198 2860
rect 4232 2859 4271 2893
rect 4305 2860 4310 2893
rect 4344 2893 4446 2894
rect 4480 2893 4582 2894
rect 4616 2893 4718 2894
rect 4752 2893 4854 2894
rect 4888 2893 4990 2894
rect 5024 2893 5126 2894
rect 5160 2893 5262 2894
rect 5296 2893 5398 2894
rect 5432 2893 5534 2894
rect 5568 2893 5670 2894
rect 5704 2893 5806 2894
rect 5840 2893 5942 2894
rect 5976 2893 6078 2894
rect 6112 2893 6214 2894
rect 6248 2893 6350 2894
rect 6384 2893 6486 2894
rect 6520 2893 6622 2894
rect 6656 2893 6758 2894
rect 6792 2893 6894 2894
rect 6928 2893 7030 2894
rect 7064 2893 7166 2894
rect 7200 2893 7302 2894
rect 7336 2893 7438 2894
rect 7472 2893 7574 2894
rect 4305 2859 4344 2860
rect 4378 2859 4417 2893
rect 4480 2860 4490 2893
rect 4451 2859 4490 2860
rect 4524 2859 4563 2893
rect 4616 2860 4636 2893
rect 4597 2859 4636 2860
rect 4670 2859 4709 2893
rect 4752 2860 4782 2893
rect 4743 2859 4782 2860
rect 4816 2860 4854 2893
rect 4816 2859 4855 2860
rect 4889 2859 4928 2893
rect 4962 2860 4990 2893
rect 4962 2859 5001 2860
rect 5035 2859 5074 2893
rect 5108 2860 5126 2893
rect 5108 2859 5147 2860
rect 5181 2859 5220 2893
rect 5254 2860 5262 2893
rect 5254 2859 5293 2860
rect 5327 2859 5366 2893
rect 5432 2860 5439 2893
rect 5400 2859 5439 2860
rect 5473 2859 5511 2893
rect 5568 2860 5583 2893
rect 5545 2859 5583 2860
rect 5617 2859 5655 2893
rect 5704 2860 5727 2893
rect 5689 2859 5727 2860
rect 5761 2859 5799 2893
rect 5840 2860 5871 2893
rect 5833 2859 5871 2860
rect 5905 2860 5942 2893
rect 5905 2859 5943 2860
rect 5977 2859 6015 2893
rect 6049 2860 6078 2893
rect 6049 2859 6087 2860
rect 6121 2859 6159 2893
rect 6193 2860 6214 2893
rect 6193 2859 6231 2860
rect 6265 2859 6303 2893
rect 6337 2860 6350 2893
rect 6337 2859 6375 2860
rect 6409 2859 6447 2893
rect 6481 2860 6486 2893
rect 6481 2859 6519 2860
rect 6553 2859 6591 2893
rect 6656 2860 6663 2893
rect 6625 2859 6663 2860
rect 6697 2859 6735 2893
rect 6792 2860 6807 2893
rect 6769 2859 6807 2860
rect 6841 2859 6879 2893
rect 6928 2860 6951 2893
rect 6913 2859 6951 2860
rect 6985 2859 7023 2893
rect 7064 2860 7095 2893
rect 7057 2859 7095 2860
rect 7129 2860 7166 2893
rect 7129 2859 7167 2860
rect 7201 2859 7239 2893
rect 7273 2860 7302 2893
rect 7273 2859 7311 2860
rect 7345 2859 7383 2893
rect 7417 2860 7438 2893
rect 7417 2859 7455 2860
rect 7489 2859 7527 2893
rect 7561 2860 7574 2893
rect 7608 2860 7710 2894
rect 7744 2860 7846 2894
rect 7880 2860 7904 2894
rect 7561 2859 7904 2860
rect 1831 2815 7904 2859
rect 1831 2781 1935 2815
rect 1969 2781 2008 2815
rect 2042 2781 2081 2815
rect 2115 2781 2154 2815
rect 2188 2781 2227 2815
rect 2261 2781 2300 2815
rect 2334 2781 2373 2815
rect 2407 2781 2446 2815
rect 2480 2781 2519 2815
rect 2553 2781 2592 2815
rect 2626 2781 2665 2815
rect 2699 2781 2738 2815
rect 2772 2781 2811 2815
rect 2845 2781 2884 2815
rect 2918 2781 2957 2815
rect 2991 2781 3030 2815
rect 3064 2781 3103 2815
rect 3137 2781 3176 2815
rect 3210 2781 3249 2815
rect 3283 2781 3322 2815
rect 3356 2781 3395 2815
rect 3429 2781 3468 2815
rect 3502 2781 3541 2815
rect 3575 2781 3614 2815
rect 3648 2781 3687 2815
rect 3721 2781 3760 2815
rect 3794 2781 3833 2815
rect 3867 2781 3906 2815
rect 3940 2781 3979 2815
rect 4013 2781 4052 2815
rect 4086 2781 4125 2815
rect 4159 2781 4198 2815
rect 4232 2781 4271 2815
rect 4305 2781 4344 2815
rect 4378 2781 4417 2815
rect 4451 2781 4490 2815
rect 4524 2781 4563 2815
rect 4597 2781 4636 2815
rect 4670 2781 4709 2815
rect 4743 2781 4782 2815
rect 4816 2781 4855 2815
rect 4889 2781 4928 2815
rect 4962 2781 5001 2815
rect 5035 2781 5074 2815
rect 5108 2781 5147 2815
rect 5181 2781 5220 2815
rect 5254 2781 5293 2815
rect 5327 2781 5366 2815
rect 5400 2781 5439 2815
rect 5473 2781 5511 2815
rect 5545 2781 5583 2815
rect 5617 2781 5655 2815
rect 5689 2781 5727 2815
rect 5761 2781 5799 2815
rect 5833 2781 5871 2815
rect 5905 2781 5943 2815
rect 5977 2781 6015 2815
rect 6049 2781 6087 2815
rect 6121 2781 6159 2815
rect 6193 2781 6231 2815
rect 6265 2781 6303 2815
rect 6337 2781 6375 2815
rect 6409 2781 6447 2815
rect 6481 2781 6519 2815
rect 6553 2781 6591 2815
rect 6625 2781 6663 2815
rect 6697 2781 6735 2815
rect 6769 2781 6807 2815
rect 6841 2781 6879 2815
rect 6913 2781 6951 2815
rect 6985 2781 7023 2815
rect 7057 2781 7095 2815
rect 7129 2781 7167 2815
rect 7201 2781 7239 2815
rect 7273 2781 7311 2815
rect 7345 2781 7383 2815
rect 7417 2781 7455 2815
rect 7489 2781 7527 2815
rect 7561 2781 7904 2815
rect 1831 2778 7904 2781
rect 1831 2744 1855 2778
rect 1889 2744 1992 2778
rect 2026 2744 2129 2778
rect 2163 2744 2266 2778
rect 2300 2744 2403 2778
rect 2437 2744 2540 2778
rect 2574 2744 2677 2778
rect 2711 2744 2814 2778
rect 2848 2744 2950 2778
rect 2984 2744 3086 2778
rect 3120 2744 3222 2778
rect 3256 2744 3358 2778
rect 3392 2744 3494 2778
rect 3528 2744 3630 2778
rect 3664 2744 3766 2778
rect 3800 2744 3902 2778
rect 3936 2744 4038 2778
rect 4072 2744 4174 2778
rect 4208 2744 4310 2778
rect 4344 2744 4446 2778
rect 4480 2744 4582 2778
rect 4616 2744 4718 2778
rect 4752 2744 4854 2778
rect 4888 2744 4990 2778
rect 5024 2744 5126 2778
rect 5160 2744 5262 2778
rect 5296 2744 5398 2778
rect 5432 2744 5534 2778
rect 5568 2744 5670 2778
rect 5704 2744 5806 2778
rect 5840 2744 5942 2778
rect 5976 2744 6078 2778
rect 6112 2744 6214 2778
rect 6248 2744 6350 2778
rect 6384 2744 6486 2778
rect 6520 2744 6622 2778
rect 6656 2744 6758 2778
rect 6792 2744 6894 2778
rect 6928 2744 7030 2778
rect 7064 2744 7166 2778
rect 7200 2744 7302 2778
rect 7336 2744 7438 2778
rect 7472 2744 7574 2778
rect 7608 2744 7710 2778
rect 7744 2744 7846 2778
rect 7880 2744 7904 2778
rect 1831 2737 7904 2744
rect 1831 2703 1935 2737
rect 1969 2703 2008 2737
rect 2042 2703 2081 2737
rect 2115 2703 2154 2737
rect 2188 2703 2227 2737
rect 2261 2703 2300 2737
rect 2334 2703 2373 2737
rect 2407 2703 2446 2737
rect 2480 2703 2519 2737
rect 2553 2703 2592 2737
rect 2626 2703 2665 2737
rect 2699 2703 2738 2737
rect 2772 2703 2811 2737
rect 2845 2703 2884 2737
rect 2918 2703 2957 2737
rect 2991 2703 3030 2737
rect 3064 2703 3103 2737
rect 3137 2703 3176 2737
rect 3210 2703 3249 2737
rect 3283 2703 3322 2737
rect 3356 2703 3395 2737
rect 3429 2703 3468 2737
rect 3502 2703 3541 2737
rect 3575 2703 3614 2737
rect 3648 2703 3687 2737
rect 3721 2703 3760 2737
rect 3794 2703 3833 2737
rect 3867 2703 3906 2737
rect 3940 2703 3979 2737
rect 4013 2703 4052 2737
rect 4086 2703 4125 2737
rect 4159 2703 4198 2737
rect 4232 2703 4271 2737
rect 4305 2703 4344 2737
rect 4378 2703 4417 2737
rect 4451 2703 4490 2737
rect 4524 2703 4563 2737
rect 4597 2703 4636 2737
rect 4670 2703 4709 2737
rect 4743 2703 4782 2737
rect 4816 2703 4855 2737
rect 4889 2703 4928 2737
rect 4962 2703 5001 2737
rect 5035 2703 5074 2737
rect 5108 2703 5147 2737
rect 5181 2703 5220 2737
rect 5254 2703 5293 2737
rect 5327 2703 5366 2737
rect 5400 2703 5439 2737
rect 5473 2703 5511 2737
rect 5545 2703 5583 2737
rect 5617 2703 5655 2737
rect 5689 2703 5727 2737
rect 5761 2703 5799 2737
rect 5833 2703 5871 2737
rect 5905 2703 5943 2737
rect 5977 2703 6015 2737
rect 6049 2703 6087 2737
rect 6121 2703 6159 2737
rect 6193 2703 6231 2737
rect 6265 2703 6303 2737
rect 6337 2703 6375 2737
rect 6409 2703 6447 2737
rect 6481 2703 6519 2737
rect 6553 2703 6591 2737
rect 6625 2703 6663 2737
rect 6697 2703 6735 2737
rect 6769 2703 6807 2737
rect 6841 2703 6879 2737
rect 6913 2703 6951 2737
rect 6985 2703 7023 2737
rect 7057 2703 7095 2737
rect 7129 2703 7167 2737
rect 7201 2703 7239 2737
rect 7273 2703 7311 2737
rect 7345 2703 7383 2737
rect 7417 2703 7455 2737
rect 7489 2703 7527 2737
rect 7561 2703 7904 2737
rect 1831 2662 7904 2703
rect 1831 2628 1855 2662
rect 1889 2659 1992 2662
rect 2026 2659 2129 2662
rect 2163 2659 2266 2662
rect 1889 2628 1935 2659
rect 1831 2625 1935 2628
rect 1969 2628 1992 2659
rect 1969 2625 2008 2628
rect 2042 2625 2081 2659
rect 2115 2628 2129 2659
rect 2115 2625 2154 2628
rect 2188 2625 2227 2659
rect 2261 2628 2266 2659
rect 2300 2659 2403 2662
rect 2437 2659 2540 2662
rect 2574 2659 2677 2662
rect 2711 2659 2814 2662
rect 2848 2659 2950 2662
rect 2984 2659 3086 2662
rect 3120 2659 3222 2662
rect 3256 2659 3358 2662
rect 2261 2625 2300 2628
rect 2334 2625 2373 2659
rect 2437 2628 2446 2659
rect 2407 2625 2446 2628
rect 2480 2625 2519 2659
rect 2574 2628 2592 2659
rect 2553 2625 2592 2628
rect 2626 2625 2665 2659
rect 2711 2628 2738 2659
rect 2699 2625 2738 2628
rect 2772 2625 2811 2659
rect 2848 2628 2884 2659
rect 2845 2625 2884 2628
rect 2918 2628 2950 2659
rect 2918 2625 2957 2628
rect 2991 2625 3030 2659
rect 3064 2628 3086 2659
rect 3064 2625 3103 2628
rect 3137 2625 3176 2659
rect 3210 2628 3222 2659
rect 3210 2625 3249 2628
rect 3283 2625 3322 2659
rect 3356 2628 3358 2659
rect 3392 2659 3494 2662
rect 3528 2659 3630 2662
rect 3664 2659 3766 2662
rect 3800 2659 3902 2662
rect 3936 2659 4038 2662
rect 4072 2659 4174 2662
rect 4208 2659 4310 2662
rect 3392 2628 3395 2659
rect 3356 2625 3395 2628
rect 3429 2625 3468 2659
rect 3528 2628 3541 2659
rect 3502 2625 3541 2628
rect 3575 2625 3614 2659
rect 3664 2628 3687 2659
rect 3648 2625 3687 2628
rect 3721 2625 3760 2659
rect 3800 2628 3833 2659
rect 3794 2625 3833 2628
rect 3867 2628 3902 2659
rect 3867 2625 3906 2628
rect 3940 2625 3979 2659
rect 4013 2628 4038 2659
rect 4013 2625 4052 2628
rect 4086 2625 4125 2659
rect 4159 2628 4174 2659
rect 4159 2625 4198 2628
rect 4232 2625 4271 2659
rect 4305 2628 4310 2659
rect 4344 2659 4446 2662
rect 4480 2659 4582 2662
rect 4616 2659 4718 2662
rect 4752 2659 4854 2662
rect 4888 2659 4990 2662
rect 5024 2659 5126 2662
rect 5160 2659 5262 2662
rect 5296 2659 5398 2662
rect 5432 2659 5534 2662
rect 5568 2659 5670 2662
rect 5704 2659 5806 2662
rect 5840 2659 5942 2662
rect 5976 2659 6078 2662
rect 6112 2659 6214 2662
rect 6248 2659 6350 2662
rect 6384 2659 6486 2662
rect 6520 2659 6622 2662
rect 6656 2659 6758 2662
rect 6792 2659 6894 2662
rect 6928 2659 7030 2662
rect 7064 2659 7166 2662
rect 7200 2659 7302 2662
rect 7336 2659 7438 2662
rect 7472 2659 7574 2662
rect 4305 2625 4344 2628
rect 4378 2625 4417 2659
rect 4480 2628 4490 2659
rect 4451 2625 4490 2628
rect 4524 2625 4563 2659
rect 4616 2628 4636 2659
rect 4597 2625 4636 2628
rect 4670 2625 4709 2659
rect 4752 2628 4782 2659
rect 4743 2625 4782 2628
rect 4816 2628 4854 2659
rect 4816 2625 4855 2628
rect 4889 2625 4928 2659
rect 4962 2628 4990 2659
rect 4962 2625 5001 2628
rect 5035 2625 5074 2659
rect 5108 2628 5126 2659
rect 5108 2625 5147 2628
rect 5181 2625 5220 2659
rect 5254 2628 5262 2659
rect 5254 2625 5293 2628
rect 5327 2625 5366 2659
rect 5432 2628 5439 2659
rect 5400 2625 5439 2628
rect 5473 2625 5511 2659
rect 5568 2628 5583 2659
rect 5545 2625 5583 2628
rect 5617 2625 5655 2659
rect 5704 2628 5727 2659
rect 5689 2625 5727 2628
rect 5761 2625 5799 2659
rect 5840 2628 5871 2659
rect 5833 2625 5871 2628
rect 5905 2628 5942 2659
rect 5905 2625 5943 2628
rect 5977 2625 6015 2659
rect 6049 2628 6078 2659
rect 6049 2625 6087 2628
rect 6121 2625 6159 2659
rect 6193 2628 6214 2659
rect 6193 2625 6231 2628
rect 6265 2625 6303 2659
rect 6337 2628 6350 2659
rect 6337 2625 6375 2628
rect 6409 2625 6447 2659
rect 6481 2628 6486 2659
rect 6481 2625 6519 2628
rect 6553 2625 6591 2659
rect 6656 2628 6663 2659
rect 6625 2625 6663 2628
rect 6697 2625 6735 2659
rect 6792 2628 6807 2659
rect 6769 2625 6807 2628
rect 6841 2625 6879 2659
rect 6928 2628 6951 2659
rect 6913 2625 6951 2628
rect 6985 2625 7023 2659
rect 7064 2628 7095 2659
rect 7057 2625 7095 2628
rect 7129 2628 7166 2659
rect 7129 2625 7167 2628
rect 7201 2625 7239 2659
rect 7273 2628 7302 2659
rect 7273 2625 7311 2628
rect 7345 2625 7383 2659
rect 7417 2628 7438 2659
rect 7417 2625 7455 2628
rect 7489 2625 7527 2659
rect 7561 2628 7574 2659
rect 7608 2628 7710 2662
rect 7744 2628 7846 2662
rect 7880 2628 7904 2662
rect 7561 2625 7904 2628
rect 1831 2581 7904 2625
rect 1831 2547 1935 2581
rect 1969 2547 2008 2581
rect 2042 2547 2081 2581
rect 2115 2547 2154 2581
rect 2188 2547 2227 2581
rect 2261 2547 2300 2581
rect 2334 2547 2373 2581
rect 2407 2547 2446 2581
rect 2480 2547 2519 2581
rect 2553 2547 2592 2581
rect 2626 2547 2665 2581
rect 2699 2547 2738 2581
rect 2772 2547 2811 2581
rect 2845 2547 2884 2581
rect 2918 2547 2957 2581
rect 2991 2547 3030 2581
rect 3064 2547 3103 2581
rect 3137 2547 3176 2581
rect 3210 2547 3249 2581
rect 3283 2547 3322 2581
rect 3356 2547 3395 2581
rect 3429 2547 3468 2581
rect 3502 2547 3541 2581
rect 3575 2547 3614 2581
rect 3648 2547 3687 2581
rect 3721 2547 3760 2581
rect 3794 2547 3833 2581
rect 3867 2547 3906 2581
rect 3940 2547 3979 2581
rect 4013 2547 4052 2581
rect 4086 2547 4125 2581
rect 4159 2547 4198 2581
rect 4232 2547 4271 2581
rect 4305 2547 4344 2581
rect 4378 2547 4417 2581
rect 4451 2547 4490 2581
rect 4524 2547 4563 2581
rect 4597 2547 4636 2581
rect 4670 2547 4709 2581
rect 4743 2547 4782 2581
rect 4816 2547 4855 2581
rect 4889 2547 4928 2581
rect 4962 2547 5001 2581
rect 5035 2547 5074 2581
rect 5108 2547 5147 2581
rect 5181 2547 5220 2581
rect 5254 2547 5293 2581
rect 5327 2547 5366 2581
rect 5400 2547 5439 2581
rect 5473 2547 5511 2581
rect 5545 2547 5583 2581
rect 5617 2547 5655 2581
rect 5689 2547 5727 2581
rect 5761 2547 5799 2581
rect 5833 2547 5871 2581
rect 5905 2547 5943 2581
rect 5977 2547 6015 2581
rect 6049 2547 6087 2581
rect 6121 2547 6159 2581
rect 6193 2547 6231 2581
rect 6265 2547 6303 2581
rect 6337 2547 6375 2581
rect 6409 2547 6447 2581
rect 6481 2547 6519 2581
rect 6553 2547 6591 2581
rect 6625 2547 6663 2581
rect 6697 2547 6735 2581
rect 6769 2547 6807 2581
rect 6841 2547 6879 2581
rect 6913 2547 6951 2581
rect 6985 2547 7023 2581
rect 7057 2547 7095 2581
rect 7129 2547 7167 2581
rect 7201 2547 7239 2581
rect 7273 2547 7311 2581
rect 7345 2547 7383 2581
rect 7417 2547 7455 2581
rect 7489 2547 7527 2581
rect 7561 2547 7904 2581
rect 1831 2546 7904 2547
rect 1831 2512 1855 2546
rect 1889 2512 1992 2546
rect 2026 2512 2129 2546
rect 2163 2512 2266 2546
rect 2300 2512 2403 2546
rect 2437 2512 2540 2546
rect 2574 2512 2677 2546
rect 2711 2512 2814 2546
rect 2848 2512 2950 2546
rect 2984 2512 3086 2546
rect 3120 2512 3222 2546
rect 3256 2512 3358 2546
rect 3392 2512 3494 2546
rect 3528 2512 3630 2546
rect 3664 2512 3766 2546
rect 3800 2512 3902 2546
rect 3936 2512 4038 2546
rect 4072 2512 4174 2546
rect 4208 2512 4310 2546
rect 4344 2512 4446 2546
rect 4480 2512 4582 2546
rect 4616 2512 4718 2546
rect 4752 2512 4854 2546
rect 4888 2512 4990 2546
rect 5024 2512 5126 2546
rect 5160 2512 5262 2546
rect 5296 2512 5398 2546
rect 5432 2512 5534 2546
rect 5568 2512 5670 2546
rect 5704 2512 5806 2546
rect 5840 2512 5942 2546
rect 5976 2512 6078 2546
rect 6112 2512 6214 2546
rect 6248 2512 6350 2546
rect 6384 2512 6486 2546
rect 6520 2512 6622 2546
rect 6656 2512 6758 2546
rect 6792 2512 6894 2546
rect 6928 2512 7030 2546
rect 7064 2512 7166 2546
rect 7200 2512 7302 2546
rect 7336 2512 7438 2546
rect 7472 2512 7574 2546
rect 7608 2512 7710 2546
rect 7744 2512 7846 2546
rect 7880 2512 7904 2546
rect 1831 2503 7904 2512
rect 1831 2469 1935 2503
rect 1969 2469 2008 2503
rect 2042 2469 2081 2503
rect 2115 2469 2154 2503
rect 2188 2469 2227 2503
rect 2261 2469 2300 2503
rect 2334 2469 2373 2503
rect 2407 2469 2446 2503
rect 2480 2469 2519 2503
rect 2553 2469 2592 2503
rect 2626 2469 2665 2503
rect 2699 2469 2738 2503
rect 2772 2469 2811 2503
rect 2845 2469 2884 2503
rect 2918 2469 2957 2503
rect 2991 2469 3030 2503
rect 3064 2469 3103 2503
rect 3137 2469 3176 2503
rect 3210 2469 3249 2503
rect 3283 2469 3322 2503
rect 3356 2469 3395 2503
rect 3429 2469 3468 2503
rect 3502 2469 3541 2503
rect 3575 2469 3614 2503
rect 3648 2469 3687 2503
rect 3721 2469 3760 2503
rect 3794 2469 3833 2503
rect 3867 2469 3906 2503
rect 3940 2469 3979 2503
rect 4013 2469 4052 2503
rect 4086 2469 4125 2503
rect 4159 2469 4198 2503
rect 4232 2469 4271 2503
rect 4305 2469 4344 2503
rect 4378 2469 4417 2503
rect 4451 2469 4490 2503
rect 4524 2469 4563 2503
rect 4597 2469 4636 2503
rect 4670 2469 4709 2503
rect 4743 2469 4782 2503
rect 4816 2469 4855 2503
rect 4889 2469 4928 2503
rect 4962 2469 5001 2503
rect 5035 2469 5074 2503
rect 5108 2469 5147 2503
rect 5181 2469 5220 2503
rect 5254 2469 5293 2503
rect 5327 2469 5366 2503
rect 5400 2469 5439 2503
rect 5473 2469 5511 2503
rect 5545 2469 5583 2503
rect 5617 2469 5655 2503
rect 5689 2469 5727 2503
rect 5761 2469 5799 2503
rect 5833 2469 5871 2503
rect 5905 2469 5943 2503
rect 5977 2469 6015 2503
rect 6049 2469 6087 2503
rect 6121 2469 6159 2503
rect 6193 2469 6231 2503
rect 6265 2469 6303 2503
rect 6337 2469 6375 2503
rect 6409 2469 6447 2503
rect 6481 2469 6519 2503
rect 6553 2469 6591 2503
rect 6625 2469 6663 2503
rect 6697 2469 6735 2503
rect 6769 2469 6807 2503
rect 6841 2469 6879 2503
rect 6913 2469 6951 2503
rect 6985 2469 7023 2503
rect 7057 2469 7095 2503
rect 7129 2469 7167 2503
rect 7201 2469 7239 2503
rect 7273 2469 7311 2503
rect 7345 2469 7383 2503
rect 7417 2469 7455 2503
rect 7489 2469 7527 2503
rect 7561 2469 7904 2503
rect 1831 2430 7904 2469
rect 1831 2396 1855 2430
rect 1889 2396 1992 2430
rect 2026 2396 2129 2430
rect 2163 2396 2266 2430
rect 2300 2396 2403 2430
rect 2437 2396 2540 2430
rect 2574 2396 2677 2430
rect 2711 2396 2814 2430
rect 2848 2396 2950 2430
rect 2984 2396 3086 2430
rect 3120 2396 3222 2430
rect 3256 2396 3358 2430
rect 3392 2396 3494 2430
rect 3528 2396 3630 2430
rect 3664 2396 3766 2430
rect 3800 2396 3902 2430
rect 3936 2396 4038 2430
rect 4072 2396 4174 2430
rect 4208 2396 4310 2430
rect 4344 2396 4446 2430
rect 4480 2396 4582 2430
rect 4616 2396 4718 2430
rect 4752 2396 4854 2430
rect 4888 2396 4990 2430
rect 5024 2396 5126 2430
rect 5160 2396 5262 2430
rect 5296 2396 5398 2430
rect 5432 2396 5534 2430
rect 5568 2396 5670 2430
rect 5704 2396 5806 2430
rect 5840 2396 5942 2430
rect 5976 2396 6078 2430
rect 6112 2396 6214 2430
rect 6248 2396 6350 2430
rect 6384 2396 6486 2430
rect 6520 2396 6622 2430
rect 6656 2396 6758 2430
rect 6792 2396 6894 2430
rect 6928 2396 7030 2430
rect 7064 2396 7166 2430
rect 7200 2396 7302 2430
rect 7336 2396 7438 2430
rect 7472 2396 7574 2430
rect 7608 2396 7710 2430
rect 7744 2396 7846 2430
rect 7880 2396 7904 2430
rect 1831 2395 7904 2396
rect 5340 2361 7594 2395
rect 5340 2327 5346 2361
rect 5380 2327 5484 2361
rect 5518 2327 5622 2361
rect 5656 2327 5760 2361
rect 5794 2327 5898 2361
rect 5932 2327 6036 2361
rect 6070 2327 6174 2361
rect 6208 2327 6312 2361
rect 6346 2327 6450 2361
rect 6484 2327 6588 2361
rect 6622 2327 6726 2361
rect 6760 2327 6864 2361
rect 6898 2327 7002 2361
rect 7036 2327 7140 2361
rect 7174 2327 7278 2361
rect 7312 2327 7416 2361
rect 7450 2327 7554 2361
rect 7588 2327 7594 2361
rect 5340 2269 7594 2327
rect 5340 2235 5414 2269
rect 5448 2235 5486 2269
rect 5520 2235 5558 2269
rect 5592 2235 5630 2269
rect 5664 2235 5702 2269
rect 5736 2235 5774 2269
rect 5808 2235 5846 2269
rect 5880 2235 5918 2269
rect 5952 2235 5990 2269
rect 6024 2235 6062 2269
rect 6096 2235 6134 2269
rect 6168 2235 6206 2269
rect 6240 2235 6278 2269
rect 6312 2235 6350 2269
rect 6384 2235 6595 2269
rect 6629 2235 6667 2269
rect 6701 2235 6739 2269
rect 6773 2235 6811 2269
rect 6845 2235 6883 2269
rect 6917 2235 6955 2269
rect 6989 2235 7027 2269
rect 7061 2235 7099 2269
rect 7133 2235 7171 2269
rect 7205 2235 7243 2269
rect 7277 2235 7315 2269
rect 7349 2235 7387 2269
rect 7421 2235 7459 2269
rect 7493 2235 7531 2269
rect 7565 2235 7594 2269
rect 5340 2223 7594 2235
rect 5340 2189 5346 2223
rect 5380 2195 5484 2223
rect 5518 2195 5622 2223
rect 5656 2195 5760 2223
rect 5794 2195 5898 2223
rect 5932 2195 6036 2223
rect 6070 2195 6174 2223
rect 6208 2195 6312 2223
rect 5380 2189 5414 2195
rect 5340 2161 5414 2189
rect 5448 2189 5484 2195
rect 5448 2161 5486 2189
rect 5520 2161 5558 2195
rect 5592 2189 5622 2195
rect 5592 2161 5630 2189
rect 5664 2161 5702 2195
rect 5736 2189 5760 2195
rect 5736 2161 5774 2189
rect 5808 2161 5846 2195
rect 5880 2189 5898 2195
rect 5880 2161 5918 2189
rect 5952 2161 5990 2195
rect 6024 2189 6036 2195
rect 6024 2161 6062 2189
rect 6096 2161 6134 2195
rect 6168 2189 6174 2195
rect 6168 2161 6206 2189
rect 6240 2161 6278 2195
rect 6346 2195 6450 2223
rect 6346 2189 6350 2195
rect 6312 2161 6350 2189
rect 6384 2189 6450 2195
rect 6484 2189 6588 2223
rect 6622 2195 6726 2223
rect 6760 2195 6864 2223
rect 6898 2195 7002 2223
rect 7036 2195 7140 2223
rect 7174 2195 7278 2223
rect 6384 2161 6595 2189
rect 6629 2161 6667 2195
rect 6701 2189 6726 2195
rect 6701 2161 6739 2189
rect 6773 2161 6811 2195
rect 6845 2189 6864 2195
rect 6845 2161 6883 2189
rect 6917 2161 6955 2195
rect 6989 2189 7002 2195
rect 6989 2161 7027 2189
rect 7061 2161 7099 2195
rect 7133 2189 7140 2195
rect 7133 2161 7171 2189
rect 7205 2161 7243 2195
rect 7277 2189 7278 2195
rect 7312 2195 7416 2223
rect 7450 2195 7554 2223
rect 7312 2189 7315 2195
rect 7277 2161 7315 2189
rect 7349 2161 7387 2195
rect 7450 2189 7459 2195
rect 7421 2161 7459 2189
rect 7493 2161 7531 2195
rect 7588 2189 7594 2223
rect 7565 2161 7594 2189
rect 5340 2121 7594 2161
rect 5340 2087 5414 2121
rect 5448 2087 5486 2121
rect 5520 2087 5558 2121
rect 5592 2087 5630 2121
rect 5664 2087 5702 2121
rect 5736 2087 5774 2121
rect 5808 2087 5846 2121
rect 5880 2087 5918 2121
rect 5952 2087 5990 2121
rect 6024 2087 6062 2121
rect 6096 2087 6134 2121
rect 6168 2087 6206 2121
rect 6240 2087 6278 2121
rect 6312 2087 6350 2121
rect 6384 2087 6595 2121
rect 6629 2087 6667 2121
rect 6701 2087 6739 2121
rect 6773 2087 6811 2121
rect 6845 2087 6883 2121
rect 6917 2087 6955 2121
rect 6989 2087 7027 2121
rect 7061 2087 7099 2121
rect 7133 2087 7171 2121
rect 7205 2087 7243 2121
rect 7277 2087 7315 2121
rect 7349 2087 7387 2121
rect 7421 2087 7459 2121
rect 7493 2087 7531 2121
rect 7565 2087 7594 2121
rect 5340 2085 7594 2087
rect 5340 2051 5346 2085
rect 5380 2051 5484 2085
rect 5518 2051 5622 2085
rect 5656 2051 5760 2085
rect 5794 2051 5898 2085
rect 5932 2051 6036 2085
rect 6070 2051 6174 2085
rect 6208 2051 6312 2085
rect 6346 2051 6450 2085
rect 6484 2051 6588 2085
rect 6622 2051 6726 2085
rect 6760 2051 6864 2085
rect 6898 2051 7002 2085
rect 7036 2051 7140 2085
rect 7174 2051 7278 2085
rect 7312 2051 7416 2085
rect 7450 2051 7554 2085
rect 7588 2051 7594 2085
rect 5340 2047 7594 2051
rect 1801 1982 1869 2016
rect 1903 1982 1937 2016
rect 1971 1982 2005 2016
rect 2039 1982 2073 2016
rect 2107 1982 2141 2016
rect 2175 1982 2209 2016
rect 2243 1982 2253 2016
rect 2311 1982 2326 2016
rect 2379 1982 2399 2016
rect 2447 1982 2472 2016
rect 2515 1982 2545 2016
rect 2583 1982 2617 2016
rect 2652 1982 2685 2016
rect 2725 1982 2753 2016
rect 2798 1982 2821 2016
rect 2871 1982 2889 2016
rect 2944 1982 2957 2016
rect 3017 1982 3025 2016
rect 3090 1982 3093 2016
rect 3127 1982 3129 2016
rect 3195 1982 3202 2016
rect 3263 1982 3275 2016
rect 3331 1982 3348 2016
rect 3399 1982 3421 2016
rect 3467 1982 3493 2016
rect 3535 1982 3565 2016
rect 3603 1982 3637 2016
rect 3671 1982 3705 2016
rect 3743 1982 3773 2016
rect 3815 1982 3841 2016
rect 3887 1982 3909 2016
rect 3959 1982 3977 2016
rect 4031 1982 4045 2016
rect 4103 1982 4113 2016
rect 4175 1982 4181 2016
rect 4247 1982 4249 2016
rect 4283 1982 4285 2016
rect 4351 1982 4357 2016
rect 4419 1982 4429 2016
rect 4487 1982 4501 2016
rect 4555 1982 4573 2016
rect 4623 1982 4645 2016
rect 4691 1982 4717 2016
rect 4759 1982 4789 2016
rect 4827 1982 4861 2016
rect 4895 1982 4929 2016
rect 4967 1982 5039 2016
rect 1801 1918 1835 1982
rect 5005 1948 5039 1982
rect 1801 1850 1835 1884
rect 2043 1883 2084 1917
rect 2118 1883 2159 1917
rect 2193 1883 2234 1917
rect 2268 1883 2309 1917
rect 2343 1883 2384 1917
rect 2418 1883 2459 1917
rect 2493 1883 2534 1917
rect 2568 1883 2609 1917
rect 2643 1883 2684 1917
rect 2718 1883 2759 1917
rect 2793 1883 2834 1917
rect 2868 1883 2909 1917
rect 2943 1883 2984 1917
rect 3018 1883 3059 1917
rect 3093 1883 3133 1917
rect 3167 1883 3207 1917
rect 3241 1883 3281 1917
rect 3315 1883 3355 1917
rect 3573 1883 3614 1917
rect 3648 1883 3689 1917
rect 3723 1883 3764 1917
rect 3798 1883 3839 1917
rect 3873 1883 3914 1917
rect 3948 1883 3989 1917
rect 4023 1883 4064 1917
rect 4098 1883 4139 1917
rect 4173 1883 4214 1917
rect 4248 1883 4289 1917
rect 4323 1883 4364 1917
rect 4398 1883 4439 1917
rect 4473 1883 4514 1917
rect 4548 1883 4589 1917
rect 4623 1883 4663 1917
rect 4697 1883 4737 1917
rect 4771 1883 4811 1917
rect 4845 1883 4885 1917
rect 5005 1880 5039 1910
rect 1801 1782 1835 1816
rect 1801 1714 1835 1748
rect 1801 1646 1835 1680
rect 1801 1578 1835 1612
rect 1801 1510 1835 1544
rect 1801 1442 1835 1476
rect 1801 1374 1835 1408
rect 1801 1306 1835 1340
rect 1801 1238 1835 1272
rect 1801 1170 1835 1204
rect 1801 1102 1835 1136
rect 1801 1034 1835 1068
rect 1919 1860 1953 1872
rect 3449 1856 3483 1872
rect 1919 1787 1953 1822
rect 2129 1791 2170 1825
rect 2204 1791 2245 1825
rect 2279 1791 2319 1825
rect 2353 1791 2393 1825
rect 2427 1791 2467 1825
rect 2501 1791 2541 1825
rect 2575 1791 2615 1825
rect 2649 1791 2689 1825
rect 2723 1791 2763 1825
rect 2797 1791 2837 1825
rect 2871 1791 2911 1825
rect 2945 1791 2985 1825
rect 3019 1791 3059 1825
rect 3093 1791 3133 1825
rect 3167 1791 3207 1825
rect 3241 1791 3281 1825
rect 3315 1791 3355 1825
rect 1919 1714 1953 1750
rect 3449 1784 3483 1822
rect 3659 1791 3699 1825
rect 3733 1791 3773 1825
rect 3807 1791 3847 1825
rect 3881 1791 3921 1825
rect 3955 1791 3994 1825
rect 4028 1791 4067 1825
rect 4101 1791 4140 1825
rect 4174 1791 4213 1825
rect 4247 1791 4286 1825
rect 4320 1791 4359 1825
rect 4393 1791 4432 1825
rect 4466 1791 4505 1825
rect 4539 1791 4578 1825
rect 4612 1791 4651 1825
rect 5005 1812 5039 1835
rect 2275 1699 2316 1733
rect 2350 1699 2391 1733
rect 2425 1699 2466 1733
rect 2500 1699 2541 1733
rect 2575 1699 2615 1733
rect 2649 1699 2689 1733
rect 2723 1699 2763 1733
rect 2797 1699 2837 1733
rect 2871 1699 2911 1733
rect 2945 1699 2985 1733
rect 3019 1699 3059 1733
rect 3093 1699 3133 1733
rect 3167 1699 3207 1733
rect 3241 1699 3281 1733
rect 3315 1699 3355 1733
rect 3449 1712 3483 1750
rect 5005 1744 5039 1760
rect 1919 1641 1953 1678
rect 3573 1699 3614 1733
rect 3648 1699 3689 1733
rect 3723 1699 3764 1733
rect 3798 1699 3839 1733
rect 3873 1699 3914 1733
rect 3948 1699 3989 1733
rect 4023 1699 4064 1733
rect 4098 1699 4139 1733
rect 4173 1699 4214 1733
rect 4248 1699 4289 1733
rect 4323 1699 4364 1733
rect 4398 1699 4439 1733
rect 4473 1699 4514 1733
rect 4548 1699 4589 1733
rect 4623 1699 4663 1733
rect 4697 1699 4737 1733
rect 4771 1699 4811 1733
rect 4845 1699 4885 1733
rect 2129 1607 2170 1641
rect 2204 1607 2245 1641
rect 2279 1607 2319 1641
rect 2353 1607 2393 1641
rect 2427 1607 2467 1641
rect 2501 1607 2541 1641
rect 2575 1607 2615 1641
rect 2649 1607 2689 1641
rect 2723 1607 2763 1641
rect 2797 1607 2837 1641
rect 2871 1607 2911 1641
rect 2945 1607 2985 1641
rect 3019 1607 3059 1641
rect 3093 1607 3133 1641
rect 3167 1607 3207 1641
rect 3241 1607 3281 1641
rect 3315 1607 3355 1641
rect 3449 1640 3483 1678
rect 5005 1676 5039 1685
rect 1919 1568 1953 1606
rect 3659 1607 3699 1641
rect 3733 1607 3773 1641
rect 3807 1607 3847 1641
rect 3881 1607 3921 1641
rect 3955 1607 3994 1641
rect 4028 1607 4067 1641
rect 4101 1607 4140 1641
rect 4174 1607 4213 1641
rect 4247 1607 4286 1641
rect 4320 1607 4359 1641
rect 4393 1607 4432 1641
rect 4466 1607 4505 1641
rect 4539 1607 4578 1641
rect 4612 1607 4651 1641
rect 5005 1608 5039 1610
rect 3449 1568 3483 1606
rect 1919 1496 1953 1534
rect 2275 1515 2316 1549
rect 2350 1515 2391 1549
rect 2425 1515 2466 1549
rect 2500 1515 2541 1549
rect 2575 1515 2615 1549
rect 2649 1515 2689 1549
rect 2723 1515 2763 1549
rect 2797 1515 2837 1549
rect 2871 1515 2911 1549
rect 2945 1515 2985 1549
rect 3019 1515 3059 1549
rect 3093 1515 3133 1549
rect 3167 1515 3207 1549
rect 3241 1515 3281 1549
rect 3315 1515 3355 1549
rect 5005 1569 5039 1574
rect 1919 1423 1953 1461
rect 3449 1496 3483 1534
rect 3573 1515 3614 1549
rect 3648 1515 3689 1549
rect 3723 1515 3764 1549
rect 3798 1515 3839 1549
rect 3873 1515 3914 1549
rect 3948 1515 3989 1549
rect 4023 1515 4064 1549
rect 4098 1515 4139 1549
rect 4173 1515 4214 1549
rect 4248 1515 4289 1549
rect 4323 1515 4364 1549
rect 4398 1515 4439 1549
rect 4473 1515 4514 1549
rect 4548 1515 4589 1549
rect 4623 1515 4663 1549
rect 4697 1515 4737 1549
rect 4771 1515 4811 1549
rect 4845 1515 4885 1549
rect 2129 1423 2170 1457
rect 2204 1423 2245 1457
rect 2279 1423 2319 1457
rect 2353 1423 2393 1457
rect 2427 1423 2467 1457
rect 2501 1423 2541 1457
rect 2575 1423 2615 1457
rect 2649 1423 2689 1457
rect 2723 1423 2763 1457
rect 2797 1423 2837 1457
rect 2871 1423 2911 1457
rect 2945 1423 2985 1457
rect 3019 1423 3059 1457
rect 3093 1423 3133 1457
rect 3167 1423 3207 1457
rect 3241 1423 3281 1457
rect 3315 1423 3355 1457
rect 3449 1423 3483 1462
rect 5005 1494 5039 1506
rect 3659 1423 3699 1457
rect 3733 1423 3773 1457
rect 3807 1423 3847 1457
rect 3881 1423 3921 1457
rect 3955 1423 3994 1457
rect 4028 1423 4067 1457
rect 4101 1423 4140 1457
rect 4174 1423 4213 1457
rect 4247 1423 4286 1457
rect 4320 1423 4359 1457
rect 4393 1423 4432 1457
rect 4466 1423 4505 1457
rect 4539 1423 4578 1457
rect 4612 1423 4651 1457
rect 1919 1350 1953 1388
rect 2275 1331 2316 1365
rect 2350 1331 2391 1365
rect 2425 1331 2466 1365
rect 2500 1331 2541 1365
rect 2575 1331 2615 1365
rect 2649 1331 2689 1365
rect 2723 1331 2763 1365
rect 2797 1331 2837 1365
rect 2871 1331 2911 1365
rect 2945 1331 2985 1365
rect 3019 1331 3059 1365
rect 3093 1331 3133 1365
rect 3167 1331 3207 1365
rect 3241 1331 3281 1365
rect 3315 1331 3355 1365
rect 3449 1350 3483 1389
rect 5005 1419 5039 1438
rect 1919 1277 1953 1315
rect 3573 1331 3614 1365
rect 3648 1331 3689 1365
rect 3723 1331 3764 1365
rect 3798 1331 3839 1365
rect 3873 1331 3914 1365
rect 3948 1331 3989 1365
rect 4023 1331 4064 1365
rect 4098 1331 4139 1365
rect 4173 1331 4214 1365
rect 4248 1331 4289 1365
rect 4323 1331 4364 1365
rect 4398 1331 4439 1365
rect 4473 1331 4514 1365
rect 4548 1331 4589 1365
rect 4623 1331 4663 1365
rect 4697 1331 4737 1365
rect 4771 1331 4811 1365
rect 4845 1331 4885 1365
rect 5005 1344 5039 1370
rect 3449 1277 3483 1316
rect 1919 1204 1953 1242
rect 2129 1239 2170 1273
rect 2204 1239 2245 1273
rect 2279 1239 2319 1273
rect 2353 1239 2393 1273
rect 2427 1239 2467 1273
rect 2501 1239 2541 1273
rect 2575 1239 2615 1273
rect 2649 1239 2689 1273
rect 2723 1239 2763 1273
rect 2797 1239 2837 1273
rect 2871 1239 2911 1273
rect 2945 1239 2985 1273
rect 3019 1239 3059 1273
rect 3093 1239 3133 1273
rect 3167 1239 3207 1273
rect 3241 1239 3281 1273
rect 3315 1239 3355 1273
rect 3449 1204 3483 1243
rect 3659 1239 3699 1273
rect 3733 1239 3773 1273
rect 3807 1239 3847 1273
rect 3881 1239 3921 1273
rect 3955 1239 3994 1273
rect 4028 1239 4067 1273
rect 4101 1239 4140 1273
rect 4174 1239 4213 1273
rect 4247 1239 4286 1273
rect 4320 1239 4359 1273
rect 4393 1239 4432 1273
rect 4466 1239 4505 1273
rect 4539 1239 4578 1273
rect 4612 1239 4651 1273
rect 5005 1270 5039 1302
rect 1919 1131 1953 1168
rect 2275 1147 2316 1181
rect 2350 1147 2391 1181
rect 2425 1147 2466 1181
rect 2500 1147 2541 1181
rect 2575 1147 2615 1181
rect 2649 1147 2689 1181
rect 2723 1147 2763 1181
rect 2797 1147 2837 1181
rect 2871 1147 2911 1181
rect 2945 1147 2985 1181
rect 3019 1147 3059 1181
rect 3093 1147 3133 1181
rect 3167 1147 3207 1181
rect 3241 1147 3281 1181
rect 3315 1147 3355 1181
rect 5005 1200 5039 1234
rect 1919 1058 1953 1094
rect 3449 1131 3483 1170
rect 3573 1147 3614 1181
rect 3648 1147 3689 1181
rect 3723 1147 3764 1181
rect 3798 1147 3839 1181
rect 3873 1147 3914 1181
rect 3948 1147 3989 1181
rect 4023 1147 4064 1181
rect 4098 1147 4139 1181
rect 4173 1147 4214 1181
rect 4248 1147 4289 1181
rect 4323 1147 4364 1181
rect 4398 1147 4439 1181
rect 4473 1147 4514 1181
rect 4548 1147 4589 1181
rect 4623 1147 4663 1181
rect 4697 1147 4737 1181
rect 4771 1147 4811 1181
rect 4845 1147 4885 1181
rect 2129 1055 2170 1089
rect 2204 1055 2245 1089
rect 2279 1055 2319 1089
rect 2353 1055 2393 1089
rect 2427 1055 2467 1089
rect 2501 1055 2541 1089
rect 2575 1055 2615 1089
rect 2649 1055 2689 1089
rect 2723 1055 2763 1089
rect 2797 1055 2837 1089
rect 2871 1055 2911 1089
rect 2945 1055 2985 1089
rect 3019 1055 3059 1089
rect 3093 1055 3133 1089
rect 3167 1055 3207 1089
rect 3241 1055 3281 1089
rect 3315 1055 3355 1089
rect 3449 1058 3483 1097
rect 5005 1132 5039 1162
rect 1919 1008 1953 1020
rect 3659 1055 3699 1089
rect 3733 1055 3773 1089
rect 3807 1055 3847 1089
rect 3881 1055 3921 1089
rect 3955 1055 3994 1089
rect 4028 1055 4067 1089
rect 4101 1055 4140 1089
rect 4174 1055 4213 1089
rect 4247 1055 4286 1089
rect 4320 1055 4359 1089
rect 4393 1055 4432 1089
rect 4466 1055 4505 1089
rect 4539 1055 4578 1089
rect 4612 1055 4651 1089
rect 5005 1064 5039 1088
rect 3449 1008 3483 1024
rect 1801 966 1835 1000
rect 5005 998 5039 1030
rect 2275 963 2316 997
rect 2350 963 2391 997
rect 2425 963 2466 997
rect 2500 963 2541 997
rect 2575 963 2615 997
rect 2649 963 2689 997
rect 2723 963 2763 997
rect 2797 963 2837 997
rect 2871 963 2911 997
rect 2945 963 2985 997
rect 3019 963 3059 997
rect 3093 963 3133 997
rect 3167 963 3207 997
rect 3241 963 3281 997
rect 3315 963 3355 997
rect 3573 963 3614 997
rect 3648 963 3689 997
rect 3723 963 3764 997
rect 3798 963 3839 997
rect 3873 963 3914 997
rect 3948 963 3989 997
rect 4023 963 4064 997
rect 4098 963 4139 997
rect 4173 963 4214 997
rect 4248 963 4289 997
rect 4323 963 4364 997
rect 4398 963 4439 997
rect 4473 963 4514 997
rect 4548 963 4589 997
rect 4623 963 4663 997
rect 4697 963 4737 997
rect 4771 963 4811 997
rect 4845 963 4885 997
rect 1801 898 1835 932
rect 5005 898 5039 962
rect 1801 864 1945 898
rect 1979 864 2013 898
rect 2047 864 2081 898
rect 2115 864 2149 898
rect 2183 864 2217 898
rect 2251 864 2285 898
rect 2319 864 2353 898
rect 2387 864 2421 898
rect 2455 864 2471 898
rect 2523 864 2543 898
rect 2591 864 2615 898
rect 2659 864 2687 898
rect 2727 864 2759 898
rect 2795 864 2829 898
rect 2865 864 2897 898
rect 2937 864 2965 898
rect 3009 864 3033 898
rect 3081 864 3101 898
rect 3153 864 3169 898
rect 3225 864 3237 898
rect 3297 864 3305 898
rect 3369 864 3373 898
rect 3475 864 3479 898
rect 3543 864 3551 898
rect 3611 864 3623 898
rect 3679 864 3695 898
rect 3747 864 3767 898
rect 3815 864 3839 898
rect 3883 864 3911 898
rect 3951 864 3984 898
rect 4019 864 4053 898
rect 4091 864 4121 898
rect 4164 864 4189 898
rect 4237 864 4257 898
rect 4310 864 4325 898
rect 4383 864 4393 898
rect 4456 864 4461 898
rect 4563 864 4568 898
rect 4631 864 4641 898
rect 4699 864 4714 898
rect 4767 864 4787 898
rect 4835 864 4860 898
rect 4903 864 4933 898
rect 4971 864 5039 898
rect 5340 2013 5414 2047
rect 5448 2013 5486 2047
rect 5520 2013 5558 2047
rect 5592 2013 5630 2047
rect 5664 2013 5702 2047
rect 5736 2013 5774 2047
rect 5808 2013 5846 2047
rect 5880 2013 5918 2047
rect 5952 2013 5990 2047
rect 6024 2013 6062 2047
rect 6096 2013 6134 2047
rect 6168 2013 6206 2047
rect 6240 2013 6278 2047
rect 6312 2013 6350 2047
rect 6384 2013 6595 2047
rect 6629 2013 6667 2047
rect 6701 2013 6739 2047
rect 6773 2013 6811 2047
rect 6845 2013 6883 2047
rect 6917 2013 6955 2047
rect 6989 2013 7027 2047
rect 7061 2013 7099 2047
rect 7133 2013 7171 2047
rect 7205 2013 7243 2047
rect 7277 2013 7315 2047
rect 7349 2013 7387 2047
rect 7421 2013 7459 2047
rect 7493 2013 7531 2047
rect 7565 2013 7594 2047
rect 5340 1973 7594 2013
rect 5340 1947 5414 1973
rect 5340 1913 5346 1947
rect 5380 1939 5414 1947
rect 5448 1947 5486 1973
rect 5448 1939 5484 1947
rect 5520 1939 5558 1973
rect 5592 1947 5630 1973
rect 5592 1939 5622 1947
rect 5664 1939 5702 1973
rect 5736 1947 5774 1973
rect 5736 1939 5760 1947
rect 5808 1939 5846 1973
rect 5880 1947 5918 1973
rect 5880 1939 5898 1947
rect 5952 1939 5990 1973
rect 6024 1947 6062 1973
rect 6024 1939 6036 1947
rect 6096 1939 6134 1973
rect 6168 1947 6206 1973
rect 6168 1939 6174 1947
rect 6240 1939 6278 1973
rect 6312 1947 6350 1973
rect 5380 1913 5484 1939
rect 5518 1913 5622 1939
rect 5656 1913 5760 1939
rect 5794 1913 5898 1939
rect 5932 1913 6036 1939
rect 6070 1913 6174 1939
rect 6208 1913 6312 1939
rect 6346 1939 6350 1947
rect 6384 1947 6595 1973
rect 6384 1939 6450 1947
rect 6346 1913 6450 1939
rect 6484 1913 6588 1947
rect 6629 1939 6667 1973
rect 6701 1947 6739 1973
rect 6701 1939 6726 1947
rect 6773 1939 6811 1973
rect 6845 1947 6883 1973
rect 6845 1939 6864 1947
rect 6917 1939 6955 1973
rect 6989 1947 7027 1973
rect 6989 1939 7002 1947
rect 7061 1939 7099 1973
rect 7133 1947 7171 1973
rect 7133 1939 7140 1947
rect 7205 1939 7243 1973
rect 7277 1947 7315 1973
rect 7277 1939 7278 1947
rect 6622 1913 6726 1939
rect 6760 1913 6864 1939
rect 6898 1913 7002 1939
rect 7036 1913 7140 1939
rect 7174 1913 7278 1939
rect 7312 1939 7315 1947
rect 7349 1939 7387 1973
rect 7421 1947 7459 1973
rect 7450 1939 7459 1947
rect 7493 1939 7531 1973
rect 7565 1947 7594 1973
rect 7312 1913 7416 1939
rect 7450 1913 7554 1939
rect 7588 1913 7594 1947
rect 5340 1899 7594 1913
rect 5340 1865 5414 1899
rect 5448 1865 5486 1899
rect 5520 1865 5558 1899
rect 5592 1865 5630 1899
rect 5664 1865 5702 1899
rect 5736 1865 5774 1899
rect 5808 1865 5846 1899
rect 5880 1865 5918 1899
rect 5952 1865 5990 1899
rect 6024 1865 6062 1899
rect 6096 1865 6134 1899
rect 6168 1865 6206 1899
rect 6240 1865 6278 1899
rect 6312 1865 6350 1899
rect 6384 1865 6595 1899
rect 6629 1865 6667 1899
rect 6701 1865 6739 1899
rect 6773 1865 6811 1899
rect 6845 1865 6883 1899
rect 6917 1865 6955 1899
rect 6989 1865 7027 1899
rect 7061 1865 7099 1899
rect 7133 1865 7171 1899
rect 7205 1865 7243 1899
rect 7277 1865 7315 1899
rect 7349 1865 7387 1899
rect 7421 1865 7459 1899
rect 7493 1865 7531 1899
rect 7565 1865 7594 1899
rect 5340 1825 7594 1865
rect 5340 1809 5414 1825
rect 5340 1775 5346 1809
rect 5380 1791 5414 1809
rect 5448 1809 5486 1825
rect 5448 1791 5484 1809
rect 5520 1791 5558 1825
rect 5592 1809 5630 1825
rect 5592 1791 5622 1809
rect 5664 1791 5702 1825
rect 5736 1809 5774 1825
rect 5736 1791 5760 1809
rect 5808 1791 5846 1825
rect 5880 1809 5918 1825
rect 5880 1791 5898 1809
rect 5952 1791 5990 1825
rect 6024 1809 6062 1825
rect 6024 1791 6036 1809
rect 6096 1791 6134 1825
rect 6168 1809 6206 1825
rect 6168 1791 6174 1809
rect 6240 1791 6278 1825
rect 6312 1809 6350 1825
rect 5380 1775 5484 1791
rect 5518 1775 5622 1791
rect 5656 1775 5760 1791
rect 5794 1775 5898 1791
rect 5932 1775 6036 1791
rect 6070 1775 6174 1791
rect 6208 1775 6312 1791
rect 6346 1791 6350 1809
rect 6384 1809 6595 1825
rect 6384 1791 6450 1809
rect 6346 1775 6450 1791
rect 6484 1775 6588 1809
rect 6629 1791 6667 1825
rect 6701 1809 6739 1825
rect 6701 1791 6726 1809
rect 6773 1791 6811 1825
rect 6845 1809 6883 1825
rect 6845 1791 6864 1809
rect 6917 1791 6955 1825
rect 6989 1809 7027 1825
rect 6989 1791 7002 1809
rect 7061 1791 7099 1825
rect 7133 1809 7171 1825
rect 7133 1791 7140 1809
rect 7205 1791 7243 1825
rect 7277 1809 7315 1825
rect 7277 1791 7278 1809
rect 6622 1775 6726 1791
rect 6760 1775 6864 1791
rect 6898 1775 7002 1791
rect 7036 1775 7140 1791
rect 7174 1775 7278 1791
rect 7312 1791 7315 1809
rect 7349 1791 7387 1825
rect 7421 1809 7459 1825
rect 7450 1791 7459 1809
rect 7493 1791 7531 1825
rect 7565 1809 7594 1825
rect 7312 1775 7416 1791
rect 7450 1775 7554 1791
rect 7588 1775 7594 1809
rect 5340 1751 7594 1775
rect 5340 1717 5414 1751
rect 5448 1717 5486 1751
rect 5520 1717 5558 1751
rect 5592 1717 5630 1751
rect 5664 1717 5702 1751
rect 5736 1717 5774 1751
rect 5808 1717 5846 1751
rect 5880 1717 5918 1751
rect 5952 1717 5990 1751
rect 6024 1717 6062 1751
rect 6096 1717 6134 1751
rect 6168 1717 6206 1751
rect 6240 1717 6278 1751
rect 6312 1717 6350 1751
rect 6384 1717 6595 1751
rect 6629 1717 6667 1751
rect 6701 1717 6739 1751
rect 6773 1717 6811 1751
rect 6845 1717 6883 1751
rect 6917 1717 6955 1751
rect 6989 1717 7027 1751
rect 7061 1717 7099 1751
rect 7133 1717 7171 1751
rect 7205 1717 7243 1751
rect 7277 1717 7315 1751
rect 7349 1717 7387 1751
rect 7421 1717 7459 1751
rect 7493 1717 7531 1751
rect 7565 1717 7594 1751
rect 5340 1676 7594 1717
rect 5340 1671 5414 1676
rect 5340 1637 5346 1671
rect 5380 1642 5414 1671
rect 5448 1671 5486 1676
rect 5448 1642 5484 1671
rect 5520 1642 5558 1676
rect 5592 1671 5630 1676
rect 5592 1642 5622 1671
rect 5664 1642 5702 1676
rect 5736 1671 5774 1676
rect 5736 1642 5760 1671
rect 5808 1642 5846 1676
rect 5880 1671 5918 1676
rect 5880 1642 5898 1671
rect 5952 1642 5990 1676
rect 6024 1671 6062 1676
rect 6024 1642 6036 1671
rect 6096 1642 6134 1676
rect 6168 1671 6206 1676
rect 6168 1642 6174 1671
rect 6240 1642 6278 1676
rect 6312 1671 6350 1676
rect 5380 1637 5484 1642
rect 5518 1637 5622 1642
rect 5656 1637 5760 1642
rect 5794 1637 5898 1642
rect 5932 1637 6036 1642
rect 6070 1637 6174 1642
rect 6208 1637 6312 1642
rect 6346 1642 6350 1671
rect 6384 1671 6595 1676
rect 6384 1642 6450 1671
rect 6346 1637 6450 1642
rect 6484 1637 6588 1671
rect 6629 1642 6667 1676
rect 6701 1671 6739 1676
rect 6701 1642 6726 1671
rect 6773 1642 6811 1676
rect 6845 1671 6883 1676
rect 6845 1642 6864 1671
rect 6917 1642 6955 1676
rect 6989 1671 7027 1676
rect 6989 1642 7002 1671
rect 7061 1642 7099 1676
rect 7133 1671 7171 1676
rect 7133 1642 7140 1671
rect 7205 1642 7243 1676
rect 7277 1671 7315 1676
rect 7277 1642 7278 1671
rect 6622 1637 6726 1642
rect 6760 1637 6864 1642
rect 6898 1637 7002 1642
rect 7036 1637 7140 1642
rect 7174 1637 7278 1642
rect 7312 1642 7315 1671
rect 7349 1642 7387 1676
rect 7421 1671 7459 1676
rect 7450 1642 7459 1671
rect 7493 1642 7531 1676
rect 7565 1671 7594 1676
rect 7312 1637 7416 1642
rect 7450 1637 7554 1642
rect 7588 1637 7594 1671
rect 5340 1601 7594 1637
rect 5340 1567 5414 1601
rect 5448 1567 5486 1601
rect 5520 1567 5558 1601
rect 5592 1567 5630 1601
rect 5664 1567 5702 1601
rect 5736 1567 5774 1601
rect 5808 1567 5846 1601
rect 5880 1567 5918 1601
rect 5952 1567 5990 1601
rect 6024 1567 6062 1601
rect 6096 1567 6134 1601
rect 6168 1567 6206 1601
rect 6240 1567 6278 1601
rect 6312 1567 6350 1601
rect 6384 1567 6595 1601
rect 6629 1567 6667 1601
rect 6701 1567 6739 1601
rect 6773 1567 6811 1601
rect 6845 1567 6883 1601
rect 6917 1567 6955 1601
rect 6989 1567 7027 1601
rect 7061 1567 7099 1601
rect 7133 1567 7171 1601
rect 7205 1567 7243 1601
rect 7277 1567 7315 1601
rect 7349 1567 7387 1601
rect 7421 1567 7459 1601
rect 7493 1567 7531 1601
rect 7565 1567 7594 1601
rect 5340 1532 7594 1567
rect 5340 1498 5346 1532
rect 5380 1526 5484 1532
rect 5518 1526 5622 1532
rect 5656 1526 5760 1532
rect 5794 1526 5898 1532
rect 5932 1526 6036 1532
rect 6070 1526 6174 1532
rect 6208 1526 6312 1532
rect 5380 1498 5414 1526
rect 5340 1492 5414 1498
rect 5448 1498 5484 1526
rect 5448 1492 5486 1498
rect 5520 1492 5558 1526
rect 5592 1498 5622 1526
rect 5592 1492 5630 1498
rect 5664 1492 5702 1526
rect 5736 1498 5760 1526
rect 5736 1492 5774 1498
rect 5808 1492 5846 1526
rect 5880 1498 5898 1526
rect 5880 1492 5918 1498
rect 5952 1492 5990 1526
rect 6024 1498 6036 1526
rect 6024 1492 6062 1498
rect 6096 1492 6134 1526
rect 6168 1498 6174 1526
rect 6168 1492 6206 1498
rect 6240 1492 6278 1526
rect 6346 1526 6450 1532
rect 6346 1498 6350 1526
rect 6312 1492 6350 1498
rect 6384 1498 6450 1526
rect 6484 1498 6588 1532
rect 6622 1526 6726 1532
rect 6760 1526 6864 1532
rect 6898 1526 7002 1532
rect 7036 1526 7140 1532
rect 7174 1526 7278 1532
rect 6384 1492 6595 1498
rect 6629 1492 6667 1526
rect 6701 1498 6726 1526
rect 6701 1492 6739 1498
rect 6773 1492 6811 1526
rect 6845 1498 6864 1526
rect 6845 1492 6883 1498
rect 6917 1492 6955 1526
rect 6989 1498 7002 1526
rect 6989 1492 7027 1498
rect 7061 1492 7099 1526
rect 7133 1498 7140 1526
rect 7133 1492 7171 1498
rect 7205 1492 7243 1526
rect 7277 1498 7278 1526
rect 7312 1526 7416 1532
rect 7450 1526 7554 1532
rect 7312 1498 7315 1526
rect 7277 1492 7315 1498
rect 7349 1492 7387 1526
rect 7450 1498 7459 1526
rect 7421 1492 7459 1498
rect 7493 1492 7531 1526
rect 7588 1498 7594 1532
rect 7565 1492 7594 1498
rect 5340 1451 7594 1492
rect 5340 1417 5414 1451
rect 5448 1417 5486 1451
rect 5520 1417 5558 1451
rect 5592 1417 5630 1451
rect 5664 1417 5702 1451
rect 5736 1417 5774 1451
rect 5808 1417 5846 1451
rect 5880 1417 5918 1451
rect 5952 1417 5990 1451
rect 6024 1417 6062 1451
rect 6096 1417 6134 1451
rect 6168 1417 6206 1451
rect 6240 1417 6278 1451
rect 6312 1417 6350 1451
rect 6384 1417 6595 1451
rect 6629 1417 6667 1451
rect 6701 1417 6739 1451
rect 6773 1417 6811 1451
rect 6845 1417 6883 1451
rect 6917 1417 6955 1451
rect 6989 1417 7027 1451
rect 7061 1417 7099 1451
rect 7133 1417 7171 1451
rect 7205 1417 7243 1451
rect 7277 1417 7315 1451
rect 7349 1417 7387 1451
rect 7421 1417 7459 1451
rect 7493 1417 7531 1451
rect 7565 1417 7594 1451
rect 5340 1393 7594 1417
rect 5340 1359 5346 1393
rect 5380 1376 5484 1393
rect 5518 1376 5622 1393
rect 5656 1376 5760 1393
rect 5794 1376 5898 1393
rect 5932 1376 6036 1393
rect 6070 1376 6174 1393
rect 6208 1376 6312 1393
rect 5380 1359 5414 1376
rect 5340 1342 5414 1359
rect 5448 1359 5484 1376
rect 5448 1342 5486 1359
rect 5520 1342 5558 1376
rect 5592 1359 5622 1376
rect 5592 1342 5630 1359
rect 5664 1342 5702 1376
rect 5736 1359 5760 1376
rect 5736 1342 5774 1359
rect 5808 1342 5846 1376
rect 5880 1359 5898 1376
rect 5880 1342 5918 1359
rect 5952 1342 5990 1376
rect 6024 1359 6036 1376
rect 6024 1342 6062 1359
rect 6096 1342 6134 1376
rect 6168 1359 6174 1376
rect 6168 1342 6206 1359
rect 6240 1342 6278 1376
rect 6346 1376 6450 1393
rect 6346 1359 6350 1376
rect 6312 1342 6350 1359
rect 6384 1359 6450 1376
rect 6484 1359 6588 1393
rect 6622 1376 6726 1393
rect 6760 1376 6864 1393
rect 6898 1376 7002 1393
rect 7036 1376 7140 1393
rect 7174 1376 7278 1393
rect 6384 1342 6595 1359
rect 6629 1342 6667 1376
rect 6701 1359 6726 1376
rect 6701 1342 6739 1359
rect 6773 1342 6811 1376
rect 6845 1359 6864 1376
rect 6845 1342 6883 1359
rect 6917 1342 6955 1376
rect 6989 1359 7002 1376
rect 6989 1342 7027 1359
rect 7061 1342 7099 1376
rect 7133 1359 7140 1376
rect 7133 1342 7171 1359
rect 7205 1342 7243 1376
rect 7277 1359 7278 1376
rect 7312 1376 7416 1393
rect 7450 1376 7554 1393
rect 7312 1359 7315 1376
rect 7277 1342 7315 1359
rect 7349 1342 7387 1376
rect 7450 1359 7459 1376
rect 7421 1342 7459 1359
rect 7493 1342 7531 1376
rect 7588 1359 7594 1393
rect 7565 1342 7594 1359
rect 5340 1301 7594 1342
rect 5340 1267 5414 1301
rect 5448 1267 5486 1301
rect 5520 1267 5558 1301
rect 5592 1267 5630 1301
rect 5664 1267 5702 1301
rect 5736 1267 5774 1301
rect 5808 1267 5846 1301
rect 5880 1267 5918 1301
rect 5952 1267 5990 1301
rect 6024 1267 6062 1301
rect 6096 1267 6134 1301
rect 6168 1267 6206 1301
rect 6240 1267 6278 1301
rect 6312 1267 6350 1301
rect 6384 1267 6595 1301
rect 6629 1267 6667 1301
rect 6701 1267 6739 1301
rect 6773 1267 6811 1301
rect 6845 1267 6883 1301
rect 6917 1267 6955 1301
rect 6989 1267 7027 1301
rect 7061 1267 7099 1301
rect 7133 1267 7171 1301
rect 7205 1267 7243 1301
rect 7277 1267 7315 1301
rect 7349 1267 7387 1301
rect 7421 1267 7459 1301
rect 7493 1267 7531 1301
rect 7565 1267 7594 1301
rect 5340 1254 7594 1267
rect 5340 1220 5346 1254
rect 5380 1226 5484 1254
rect 5518 1226 5622 1254
rect 5656 1226 5760 1254
rect 5794 1226 5898 1254
rect 5932 1226 6036 1254
rect 6070 1226 6174 1254
rect 6208 1226 6312 1254
rect 5380 1220 5414 1226
rect 5340 1192 5414 1220
rect 5448 1220 5484 1226
rect 5448 1192 5486 1220
rect 5520 1192 5558 1226
rect 5592 1220 5622 1226
rect 5592 1192 5630 1220
rect 5664 1192 5702 1226
rect 5736 1220 5760 1226
rect 5736 1192 5774 1220
rect 5808 1192 5846 1226
rect 5880 1220 5898 1226
rect 5880 1192 5918 1220
rect 5952 1192 5990 1226
rect 6024 1220 6036 1226
rect 6024 1192 6062 1220
rect 6096 1192 6134 1226
rect 6168 1220 6174 1226
rect 6168 1192 6206 1220
rect 6240 1192 6278 1226
rect 6346 1226 6450 1254
rect 6346 1220 6350 1226
rect 6312 1192 6350 1220
rect 6384 1220 6450 1226
rect 6484 1220 6588 1254
rect 6622 1226 6726 1254
rect 6760 1226 6864 1254
rect 6898 1226 7002 1254
rect 7036 1226 7140 1254
rect 7174 1226 7278 1254
rect 6384 1192 6595 1220
rect 6629 1192 6667 1226
rect 6701 1220 6726 1226
rect 6701 1192 6739 1220
rect 6773 1192 6811 1226
rect 6845 1220 6864 1226
rect 6845 1192 6883 1220
rect 6917 1192 6955 1226
rect 6989 1220 7002 1226
rect 6989 1192 7027 1220
rect 7061 1192 7099 1226
rect 7133 1220 7140 1226
rect 7133 1192 7171 1220
rect 7205 1192 7243 1226
rect 7277 1220 7278 1226
rect 7312 1226 7416 1254
rect 7450 1226 7554 1254
rect 7312 1220 7315 1226
rect 7277 1192 7315 1220
rect 7349 1192 7387 1226
rect 7450 1220 7459 1226
rect 7421 1192 7459 1220
rect 7493 1192 7531 1226
rect 7588 1220 7594 1254
rect 7565 1192 7594 1220
rect 5340 1151 7594 1192
rect 5340 1117 5414 1151
rect 5448 1117 5486 1151
rect 5520 1117 5558 1151
rect 5592 1117 5630 1151
rect 5664 1117 5702 1151
rect 5736 1117 5774 1151
rect 5808 1117 5846 1151
rect 5880 1117 5918 1151
rect 5952 1117 5990 1151
rect 6024 1117 6062 1151
rect 6096 1117 6134 1151
rect 6168 1117 6206 1151
rect 6240 1117 6278 1151
rect 6312 1117 6350 1151
rect 6384 1117 6595 1151
rect 6629 1117 6667 1151
rect 6701 1117 6739 1151
rect 6773 1117 6811 1151
rect 6845 1117 6883 1151
rect 6917 1117 6955 1151
rect 6989 1117 7027 1151
rect 7061 1117 7099 1151
rect 7133 1117 7171 1151
rect 7205 1117 7243 1151
rect 7277 1117 7315 1151
rect 7349 1117 7387 1151
rect 7421 1117 7459 1151
rect 7493 1117 7531 1151
rect 7565 1117 7594 1151
rect 5340 1115 7594 1117
rect 5340 1081 5346 1115
rect 5380 1081 5484 1115
rect 5518 1081 5622 1115
rect 5656 1081 5760 1115
rect 5794 1081 5898 1115
rect 5932 1081 6036 1115
rect 6070 1081 6174 1115
rect 6208 1081 6312 1115
rect 6346 1081 6450 1115
rect 6484 1081 6588 1115
rect 6622 1081 6726 1115
rect 6760 1081 6864 1115
rect 6898 1081 7002 1115
rect 7036 1081 7140 1115
rect 7174 1081 7278 1115
rect 7312 1081 7416 1115
rect 7450 1081 7554 1115
rect 7588 1081 7594 1115
rect 5340 1076 7594 1081
rect 5340 1042 5414 1076
rect 5448 1042 5486 1076
rect 5520 1042 5558 1076
rect 5592 1042 5630 1076
rect 5664 1042 5702 1076
rect 5736 1042 5774 1076
rect 5808 1042 5846 1076
rect 5880 1042 5918 1076
rect 5952 1042 5990 1076
rect 6024 1042 6062 1076
rect 6096 1042 6134 1076
rect 6168 1042 6206 1076
rect 6240 1042 6278 1076
rect 6312 1042 6350 1076
rect 6384 1042 6595 1076
rect 6629 1042 6667 1076
rect 6701 1042 6739 1076
rect 6773 1042 6811 1076
rect 6845 1042 6883 1076
rect 6917 1042 6955 1076
rect 6989 1042 7027 1076
rect 7061 1042 7099 1076
rect 7133 1042 7171 1076
rect 7205 1042 7243 1076
rect 7277 1042 7315 1076
rect 7349 1042 7387 1076
rect 7421 1042 7459 1076
rect 7493 1042 7531 1076
rect 7565 1042 7594 1076
rect 5340 1001 7594 1042
rect 5340 976 5414 1001
rect 5340 942 5346 976
rect 5380 967 5414 976
rect 5448 976 5486 1001
rect 5448 967 5484 976
rect 5520 967 5558 1001
rect 5592 976 5630 1001
rect 5592 967 5622 976
rect 5664 967 5702 1001
rect 5736 976 5774 1001
rect 5736 967 5760 976
rect 5808 967 5846 1001
rect 5880 976 5918 1001
rect 5880 967 5898 976
rect 5952 967 5990 1001
rect 6024 976 6062 1001
rect 6024 967 6036 976
rect 6096 967 6134 1001
rect 6168 976 6206 1001
rect 6168 967 6174 976
rect 6240 967 6278 1001
rect 6312 976 6350 1001
rect 5380 942 5484 967
rect 5518 942 5622 967
rect 5656 942 5760 967
rect 5794 942 5898 967
rect 5932 942 6036 967
rect 6070 942 6174 967
rect 6208 942 6312 967
rect 6346 967 6350 976
rect 6384 976 6595 1001
rect 6384 967 6450 976
rect 6346 942 6450 967
rect 6484 942 6588 976
rect 6629 967 6667 1001
rect 6701 976 6739 1001
rect 6701 967 6726 976
rect 6773 967 6811 1001
rect 6845 976 6883 1001
rect 6845 967 6864 976
rect 6917 967 6955 1001
rect 6989 976 7027 1001
rect 6989 967 7002 976
rect 7061 967 7099 1001
rect 7133 976 7171 1001
rect 7133 967 7140 976
rect 7205 967 7243 1001
rect 7277 976 7315 1001
rect 7277 967 7278 976
rect 6622 942 6726 967
rect 6760 942 6864 967
rect 6898 942 7002 967
rect 7036 942 7140 967
rect 7174 942 7278 967
rect 7312 967 7315 976
rect 7349 967 7387 1001
rect 7421 976 7459 1001
rect 7450 967 7459 976
rect 7493 967 7531 1001
rect 7565 976 7594 1001
rect 7312 942 7416 967
rect 7450 942 7554 967
rect 7588 942 7594 976
rect 5340 926 7594 942
rect 5340 892 5414 926
rect 5448 892 5486 926
rect 5520 892 5558 926
rect 5592 892 5630 926
rect 5664 892 5702 926
rect 5736 892 5774 926
rect 5808 892 5846 926
rect 5880 892 5918 926
rect 5952 892 5990 926
rect 6024 892 6062 926
rect 6096 892 6134 926
rect 6168 892 6206 926
rect 6240 892 6278 926
rect 6312 892 6350 926
rect 6384 892 6595 926
rect 6629 892 6667 926
rect 6701 892 6739 926
rect 6773 892 6811 926
rect 6845 892 6883 926
rect 6917 892 6955 926
rect 6989 892 7027 926
rect 7061 892 7099 926
rect 7133 892 7171 926
rect 7205 892 7243 926
rect 7277 892 7315 926
rect 7349 892 7387 926
rect 7421 892 7459 926
rect 7493 892 7531 926
rect 7565 892 7594 926
rect 5340 851 7594 892
rect 5340 837 5414 851
rect 5340 803 5346 837
rect 5380 817 5414 837
rect 5448 837 5486 851
rect 5448 817 5484 837
rect 5520 817 5558 851
rect 5592 837 5630 851
rect 5592 817 5622 837
rect 5664 817 5702 851
rect 5736 837 5774 851
rect 5736 817 5760 837
rect 5808 817 5846 851
rect 5880 837 5918 851
rect 5880 817 5898 837
rect 5952 817 5990 851
rect 6024 837 6062 851
rect 6024 817 6036 837
rect 6096 817 6134 851
rect 6168 837 6206 851
rect 6168 817 6174 837
rect 6240 817 6278 851
rect 6312 837 6350 851
rect 5380 803 5484 817
rect 5518 803 5622 817
rect 5656 803 5760 817
rect 5794 803 5898 817
rect 5932 803 6036 817
rect 6070 803 6174 817
rect 6208 803 6312 817
rect 6346 817 6350 837
rect 6384 837 6595 851
rect 6384 817 6450 837
rect 6346 803 6450 817
rect 6484 803 6588 837
rect 6629 817 6667 851
rect 6701 837 6739 851
rect 6701 817 6726 837
rect 6773 817 6811 851
rect 6845 837 6883 851
rect 6845 817 6864 837
rect 6917 817 6955 851
rect 6989 837 7027 851
rect 6989 817 7002 837
rect 7061 817 7099 851
rect 7133 837 7171 851
rect 7133 817 7140 837
rect 7205 817 7243 851
rect 7277 837 7315 851
rect 7277 817 7278 837
rect 6622 803 6726 817
rect 6760 803 6864 817
rect 6898 803 7002 817
rect 7036 803 7140 817
rect 7174 803 7278 817
rect 7312 817 7315 837
rect 7349 817 7387 851
rect 7421 837 7459 851
rect 7450 817 7459 837
rect 7493 817 7531 851
rect 7565 837 7594 851
rect 7312 803 7416 817
rect 7450 803 7554 817
rect 7588 803 7594 837
rect 5340 776 7594 803
rect 5340 742 5414 776
rect 5448 742 5486 776
rect 5520 742 5558 776
rect 5592 742 5630 776
rect 5664 742 5702 776
rect 5736 742 5774 776
rect 5808 742 5846 776
rect 5880 742 5918 776
rect 5952 742 5990 776
rect 6024 742 6062 776
rect 6096 742 6134 776
rect 6168 742 6206 776
rect 6240 742 6278 776
rect 6312 742 6350 776
rect 6384 742 6595 776
rect 6629 742 6667 776
rect 6701 742 6739 776
rect 6773 742 6811 776
rect 6845 742 6883 776
rect 6917 742 6955 776
rect 6989 742 7027 776
rect 7061 742 7099 776
rect 7133 742 7171 776
rect 7205 742 7243 776
rect 7277 742 7315 776
rect 7349 742 7387 776
rect 7421 742 7459 776
rect 7493 742 7531 776
rect 7565 742 7594 776
rect 5340 701 7594 742
rect 5340 698 5414 701
rect 5340 664 5346 698
rect 5380 667 5414 698
rect 5448 698 5486 701
rect 5448 667 5484 698
rect 5520 667 5558 701
rect 5592 698 5630 701
rect 5592 667 5622 698
rect 5664 667 5702 701
rect 5736 698 5774 701
rect 5736 667 5760 698
rect 5808 667 5846 701
rect 5880 698 5918 701
rect 5880 667 5898 698
rect 5952 667 5990 701
rect 6024 698 6062 701
rect 6024 667 6036 698
rect 6096 667 6134 701
rect 6168 698 6206 701
rect 6168 667 6174 698
rect 6240 667 6278 701
rect 6312 698 6350 701
rect 5380 664 5484 667
rect 5518 664 5622 667
rect 5656 664 5760 667
rect 5794 664 5898 667
rect 5932 664 6036 667
rect 6070 664 6174 667
rect 6208 664 6312 667
rect 6346 667 6350 698
rect 6384 698 6595 701
rect 6384 667 6450 698
rect 6346 664 6450 667
rect 6484 664 6588 698
rect 6629 667 6667 701
rect 6701 698 6739 701
rect 6701 667 6726 698
rect 6773 667 6811 701
rect 6845 698 6883 701
rect 6845 667 6864 698
rect 6917 667 6955 701
rect 6989 698 7027 701
rect 6989 667 7002 698
rect 7061 667 7099 701
rect 7133 698 7171 701
rect 7133 667 7140 698
rect 7205 667 7243 701
rect 7277 698 7315 701
rect 7277 667 7278 698
rect 6622 664 6726 667
rect 6760 664 6864 667
rect 6898 664 7002 667
rect 7036 664 7140 667
rect 7174 664 7278 667
rect 7312 667 7315 698
rect 7349 667 7387 701
rect 7421 698 7459 701
rect 7450 667 7459 698
rect 7493 667 7531 701
rect 7565 698 7594 701
rect 7312 664 7416 667
rect 7450 664 7554 667
rect 7588 664 7594 698
rect 5340 626 7594 664
rect 5340 592 5414 626
rect 5448 592 5486 626
rect 5520 592 5558 626
rect 5592 592 5630 626
rect 5664 592 5702 626
rect 5736 592 5774 626
rect 5808 592 5846 626
rect 5880 592 5918 626
rect 5952 592 5990 626
rect 6024 592 6062 626
rect 6096 592 6134 626
rect 6168 592 6206 626
rect 6240 592 6278 626
rect 6312 592 6350 626
rect 6384 592 6595 626
rect 6629 592 6667 626
rect 6701 592 6739 626
rect 6773 592 6811 626
rect 6845 592 6883 626
rect 6917 592 6955 626
rect 6989 592 7027 626
rect 7061 592 7099 626
rect 7133 592 7171 626
rect 7205 592 7243 626
rect 7277 592 7315 626
rect 7349 592 7387 626
rect 7421 592 7459 626
rect 7493 592 7531 626
rect 7565 592 7594 626
rect 5340 559 7594 592
rect 5340 525 5346 559
rect 5380 551 5484 559
rect 5518 551 5622 559
rect 5656 551 5760 559
rect 5794 551 5898 559
rect 5932 551 6036 559
rect 6070 551 6174 559
rect 6208 551 6312 559
rect 5380 525 5414 551
rect 5340 517 5414 525
rect 5448 525 5484 551
rect 5448 517 5486 525
rect 5520 517 5558 551
rect 5592 525 5622 551
rect 5592 517 5630 525
rect 5664 517 5702 551
rect 5736 525 5760 551
rect 5736 517 5774 525
rect 5808 517 5846 551
rect 5880 525 5898 551
rect 5880 517 5918 525
rect 5952 517 5990 551
rect 6024 525 6036 551
rect 6024 517 6062 525
rect 6096 517 6134 551
rect 6168 525 6174 551
rect 6168 517 6206 525
rect 6240 517 6278 551
rect 6346 551 6450 559
rect 6346 525 6350 551
rect 6312 517 6350 525
rect 6384 525 6450 551
rect 6484 525 6588 559
rect 6622 551 6726 559
rect 6760 551 6864 559
rect 6898 551 7002 559
rect 7036 551 7140 559
rect 7174 551 7278 559
rect 6384 517 6595 525
rect 6629 517 6667 551
rect 6701 525 6726 551
rect 6701 517 6739 525
rect 6773 517 6811 551
rect 6845 525 6864 551
rect 6845 517 6883 525
rect 6917 517 6955 551
rect 6989 525 7002 551
rect 6989 517 7027 525
rect 7061 517 7099 551
rect 7133 525 7140 551
rect 7133 517 7171 525
rect 7205 517 7243 551
rect 7277 525 7278 551
rect 7312 551 7416 559
rect 7450 551 7554 559
rect 7312 525 7315 551
rect 7277 517 7315 525
rect 7349 517 7387 551
rect 7450 525 7459 551
rect 7421 517 7459 525
rect 7493 517 7531 551
rect 7588 525 7594 559
rect 7565 517 7594 525
rect 5340 476 7594 517
rect 5340 442 5414 476
rect 5448 442 5486 476
rect 5520 442 5558 476
rect 5592 442 5630 476
rect 5664 442 5702 476
rect 5736 442 5774 476
rect 5808 442 5846 476
rect 5880 442 5918 476
rect 5952 442 5990 476
rect 6024 442 6062 476
rect 6096 442 6134 476
rect 6168 442 6206 476
rect 6240 442 6278 476
rect 6312 442 6350 476
rect 6384 442 6595 476
rect 6629 442 6667 476
rect 6701 442 6739 476
rect 6773 442 6811 476
rect 6845 442 6883 476
rect 6917 442 6955 476
rect 6989 442 7027 476
rect 7061 442 7099 476
rect 7133 442 7171 476
rect 7205 442 7243 476
rect 7277 442 7315 476
rect 7349 442 7387 476
rect 7421 442 7459 476
rect 7493 442 7531 476
rect 7565 442 7594 476
rect 5340 420 7594 442
rect 5340 386 5346 420
rect 5380 386 5484 420
rect 5518 386 5622 420
rect 5656 386 5760 420
rect 5794 386 5898 420
rect 5932 386 6036 420
rect 6070 386 6174 420
rect 6208 386 6312 420
rect 6346 386 6450 420
rect 6484 386 6588 420
rect 6622 386 6726 420
rect 6760 386 6864 420
rect 6898 386 7002 420
rect 7036 386 7140 420
rect 7174 386 7278 420
rect 7312 386 7416 420
rect 7450 386 7554 420
rect 7588 386 7594 420
rect 5340 352 7594 386
rect 1392 307 1451 341
rect 1485 307 1543 341
rect 1577 307 1635 341
rect 1358 299 1669 307
rect 115 262 175 296
rect 209 262 219 296
rect 81 221 219 262
rect 81 213 170 221
rect 204 213 219 221
rect 115 187 170 213
rect 115 179 175 187
rect 209 179 219 213
rect 81 153 219 179
rect 81 130 170 153
rect 204 130 219 153
rect 115 119 170 130
rect 115 96 175 119
rect 209 96 219 130
rect 1358 269 1678 299
rect 1392 235 1451 269
rect 1485 235 1543 269
rect 1577 235 1635 269
rect 1669 235 1678 269
rect 1358 221 1678 235
rect 1358 187 1628 221
rect 1662 187 1678 221
rect 1358 153 1678 187
rect 1358 119 1628 153
rect 1662 119 1678 153
rect 1358 103 1678 119
<< viali >>
rect 2163 39474 2989 39476
rect 3028 39474 3062 39476
rect 3101 39474 3135 39476
rect 3174 39474 3208 39476
rect 3247 39474 3281 39476
rect 3320 39474 3354 39476
rect 3393 39474 3427 39476
rect 3466 39474 3500 39476
rect 3539 39474 3573 39476
rect 3612 39474 3646 39476
rect 3685 39474 3719 39476
rect 3758 39474 3792 39476
rect 3831 39474 3865 39476
rect 3904 39474 3938 39476
rect 3977 39474 4011 39476
rect 4050 39474 4084 39476
rect 4123 39474 4157 39476
rect 4196 39474 4230 39476
rect 4269 39474 4303 39476
rect 4342 39474 4376 39476
rect 4415 39474 4449 39476
rect 4488 39474 4522 39476
rect 4561 39474 4595 39476
rect 4634 39474 4668 39476
rect 4707 39474 4741 39476
rect 4780 39474 4814 39476
rect 4853 39474 4887 39476
rect 4926 39474 4960 39476
rect 4999 39474 5033 39476
rect 5072 39474 5106 39476
rect 5145 39474 5179 39476
rect 5218 39474 5252 39476
rect 5291 39474 5325 39476
rect 5364 39474 5398 39476
rect 5437 39474 5471 39476
rect 5510 39474 5544 39476
rect 5583 39474 5617 39476
rect 5656 39474 5690 39476
rect 5729 39474 5763 39476
rect 5802 39474 5836 39476
rect 5875 39474 5909 39476
rect 5948 39474 5982 39476
rect 6021 39474 6055 39476
rect 6094 39474 6128 39476
rect 6167 39474 6201 39476
rect 6240 39474 6274 39476
rect 6313 39474 6347 39476
rect 6386 39474 6420 39476
rect 6459 39474 6493 39476
rect 6532 39474 6566 39476
rect 6605 39474 6639 39476
rect 6678 39474 6712 39476
rect 6751 39474 6785 39476
rect 6824 39474 6858 39476
rect 6897 39474 6931 39476
rect 6970 39474 7004 39476
rect 7043 39474 7077 39476
rect 7116 39474 7150 39476
rect 7189 39474 7223 39476
rect 7262 39474 7296 39476
rect 7335 39474 7369 39476
rect 7408 39474 7442 39476
rect 7481 39474 7515 39476
rect 7554 39474 7588 39476
rect 7627 39474 7661 39476
rect 7786 39474 7820 39476
rect 7866 39474 7900 39476
rect 7946 39474 7980 39476
rect 8026 39474 8060 39476
rect 8106 39474 8140 39476
rect 8186 39474 8220 39476
rect 8267 39474 8301 39476
rect 8348 39474 8382 39476
rect 8429 39474 8463 39476
rect 1944 39440 2039 39470
rect 2039 39440 2050 39470
rect 1944 39406 2050 39440
rect 1944 34108 1946 39406
rect 1946 34108 2048 39406
rect 2048 34108 2050 39406
rect 2163 39372 2989 39474
rect 3028 39442 3062 39474
rect 3101 39442 3135 39474
rect 3174 39442 3208 39474
rect 3247 39442 3281 39474
rect 3320 39442 3354 39474
rect 3393 39442 3427 39474
rect 3466 39442 3500 39474
rect 3539 39442 3573 39474
rect 3612 39442 3646 39474
rect 3685 39442 3719 39474
rect 3758 39442 3792 39474
rect 3831 39442 3865 39474
rect 3904 39442 3938 39474
rect 3977 39442 4011 39474
rect 4050 39442 4084 39474
rect 4123 39442 4157 39474
rect 4196 39442 4230 39474
rect 4269 39442 4303 39474
rect 4342 39442 4376 39474
rect 4415 39442 4449 39474
rect 4488 39442 4522 39474
rect 4561 39442 4595 39474
rect 4634 39442 4668 39474
rect 4707 39442 4741 39474
rect 4780 39442 4814 39474
rect 4853 39442 4887 39474
rect 4926 39442 4960 39474
rect 4999 39442 5033 39474
rect 5072 39442 5106 39474
rect 5145 39442 5179 39474
rect 5218 39442 5252 39474
rect 5291 39442 5325 39474
rect 5364 39442 5398 39474
rect 5437 39442 5471 39474
rect 5510 39442 5544 39474
rect 5583 39442 5617 39474
rect 5656 39442 5690 39474
rect 5729 39442 5763 39474
rect 5802 39442 5836 39474
rect 5875 39442 5909 39474
rect 5948 39442 5982 39474
rect 6021 39442 6055 39474
rect 6094 39442 6128 39474
rect 6167 39442 6201 39474
rect 6240 39442 6274 39474
rect 6313 39442 6347 39474
rect 6386 39442 6420 39474
rect 6459 39442 6493 39474
rect 6532 39442 6566 39474
rect 6605 39442 6639 39474
rect 6678 39442 6712 39474
rect 6751 39442 6785 39474
rect 6824 39442 6858 39474
rect 6897 39442 6931 39474
rect 6970 39442 7004 39474
rect 7043 39442 7077 39474
rect 7116 39442 7150 39474
rect 7189 39442 7223 39474
rect 7262 39442 7296 39474
rect 7335 39442 7369 39474
rect 7408 39442 7442 39474
rect 7481 39442 7515 39474
rect 7554 39442 7588 39474
rect 7627 39442 7661 39474
rect 7786 39442 7820 39474
rect 7866 39442 7900 39474
rect 7946 39442 7980 39474
rect 8026 39442 8060 39474
rect 8106 39442 8140 39474
rect 8186 39442 8220 39474
rect 8267 39442 8301 39474
rect 8348 39442 8382 39474
rect 8429 39442 8463 39474
rect 3028 39372 3062 39404
rect 3101 39372 3135 39404
rect 3174 39372 3208 39404
rect 3247 39372 3281 39404
rect 3320 39372 3354 39404
rect 3393 39372 3427 39404
rect 3466 39372 3500 39404
rect 3539 39372 3573 39404
rect 3612 39372 3646 39404
rect 3685 39372 3719 39404
rect 3758 39372 3792 39404
rect 3831 39372 3865 39404
rect 3904 39372 3938 39404
rect 3977 39372 4011 39404
rect 4050 39372 4084 39404
rect 4123 39372 4157 39404
rect 4196 39372 4230 39404
rect 4269 39372 4303 39404
rect 4342 39372 4376 39404
rect 4415 39372 4449 39404
rect 4488 39372 4522 39404
rect 4561 39372 4595 39404
rect 4634 39372 4668 39404
rect 4707 39372 4741 39404
rect 4780 39372 4814 39404
rect 4853 39372 4887 39404
rect 4926 39372 4960 39404
rect 4999 39372 5033 39404
rect 5072 39372 5106 39404
rect 5145 39372 5179 39404
rect 5218 39372 5252 39404
rect 5291 39372 5325 39404
rect 5364 39372 5398 39404
rect 5437 39372 5471 39404
rect 5510 39372 5544 39404
rect 5583 39372 5617 39404
rect 5656 39372 5690 39404
rect 5729 39372 5763 39404
rect 5802 39372 5836 39404
rect 5875 39372 5909 39404
rect 5948 39372 5982 39404
rect 6021 39372 6055 39404
rect 6094 39372 6128 39404
rect 6167 39372 6201 39404
rect 6240 39372 6274 39404
rect 6313 39372 6347 39404
rect 6386 39372 6420 39404
rect 6459 39372 6493 39404
rect 6532 39372 6566 39404
rect 6605 39372 6639 39404
rect 6678 39372 6712 39404
rect 6751 39372 6785 39404
rect 6824 39372 6858 39404
rect 6897 39372 6931 39404
rect 6970 39372 7004 39404
rect 7043 39372 7077 39404
rect 7116 39372 7150 39404
rect 7189 39372 7223 39404
rect 7262 39372 7296 39404
rect 7335 39372 7369 39404
rect 7408 39372 7442 39404
rect 7481 39372 7515 39404
rect 7554 39372 7588 39404
rect 7627 39372 7661 39404
rect 7786 39372 7820 39404
rect 7866 39372 7900 39404
rect 7946 39372 7980 39404
rect 8026 39372 8060 39404
rect 8106 39372 8140 39404
rect 8186 39372 8220 39404
rect 8267 39372 8301 39404
rect 8348 39372 8382 39404
rect 8429 39372 8465 39404
rect 8465 39372 8535 39404
rect 2163 39370 2989 39372
rect 3028 39370 3062 39372
rect 3101 39370 3135 39372
rect 3174 39370 3208 39372
rect 3247 39370 3281 39372
rect 3320 39370 3354 39372
rect 3393 39370 3427 39372
rect 3466 39370 3500 39372
rect 3539 39370 3573 39372
rect 3612 39370 3646 39372
rect 3685 39370 3719 39372
rect 3758 39370 3792 39372
rect 3831 39370 3865 39372
rect 3904 39370 3938 39372
rect 3977 39370 4011 39372
rect 4050 39370 4084 39372
rect 4123 39370 4157 39372
rect 4196 39370 4230 39372
rect 4269 39370 4303 39372
rect 4342 39370 4376 39372
rect 4415 39370 4449 39372
rect 4488 39370 4522 39372
rect 4561 39370 4595 39372
rect 4634 39370 4668 39372
rect 4707 39370 4741 39372
rect 4780 39370 4814 39372
rect 4853 39370 4887 39372
rect 4926 39370 4960 39372
rect 4999 39370 5033 39372
rect 5072 39370 5106 39372
rect 5145 39370 5179 39372
rect 5218 39370 5252 39372
rect 5291 39370 5325 39372
rect 5364 39370 5398 39372
rect 5437 39370 5471 39372
rect 5510 39370 5544 39372
rect 5583 39370 5617 39372
rect 5656 39370 5690 39372
rect 5729 39370 5763 39372
rect 5802 39370 5836 39372
rect 5875 39370 5909 39372
rect 5948 39370 5982 39372
rect 6021 39370 6055 39372
rect 6094 39370 6128 39372
rect 6167 39370 6201 39372
rect 6240 39370 6274 39372
rect 6313 39370 6347 39372
rect 6386 39370 6420 39372
rect 6459 39370 6493 39372
rect 6532 39370 6566 39372
rect 6605 39370 6639 39372
rect 6678 39370 6712 39372
rect 6751 39370 6785 39372
rect 6824 39370 6858 39372
rect 6897 39370 6931 39372
rect 6970 39370 7004 39372
rect 7043 39370 7077 39372
rect 7116 39370 7150 39372
rect 7189 39370 7223 39372
rect 7262 39370 7296 39372
rect 7335 39370 7369 39372
rect 7408 39370 7442 39372
rect 7481 39370 7515 39372
rect 7554 39370 7588 39372
rect 7627 39370 7661 39372
rect 7786 39370 7820 39372
rect 7866 39370 7900 39372
rect 7946 39370 7980 39372
rect 8026 39370 8060 39372
rect 8106 39370 8140 39372
rect 8186 39370 8220 39372
rect 8267 39370 8301 39372
rect 8348 39370 8382 39372
rect 8429 39354 8535 39372
rect 8429 39320 8499 39354
rect 8499 39320 8533 39354
rect 8533 39320 8535 39354
rect 8429 39286 8535 39320
rect 1944 34035 1946 34069
rect 1946 34035 1978 34069
rect 2016 34035 2048 34069
rect 2048 34035 2050 34069
rect 1944 33962 1946 33996
rect 1946 33962 1978 33996
rect 2016 33962 2048 33996
rect 2048 33962 2050 33996
rect 1944 33889 1946 33923
rect 1946 33889 1978 33923
rect 2016 33889 2048 33923
rect 2048 33889 2050 33923
rect 1944 33816 1946 33850
rect 1946 33816 1978 33850
rect 2016 33816 2048 33850
rect 2048 33816 2050 33850
rect 1944 33743 1946 33777
rect 1946 33743 1978 33777
rect 2016 33743 2048 33777
rect 2048 33743 2050 33777
rect 1944 33670 1946 33704
rect 1946 33670 1978 33704
rect 2016 33670 2048 33704
rect 2048 33670 2050 33704
rect 1944 11037 1946 33607
rect 1946 11037 2048 33607
rect 2048 11037 2050 33607
rect 1944 10964 1946 10998
rect 1946 10964 1978 10998
rect 2016 10964 2048 10998
rect 2048 10964 2050 10998
rect 1944 10891 1946 10925
rect 1946 10891 1978 10925
rect 2016 10891 2048 10925
rect 2048 10891 2050 10925
rect 1944 10813 1946 10847
rect 1946 10813 1978 10847
rect 2016 10813 2048 10847
rect 2048 10813 2050 10847
rect 1944 10740 1946 10774
rect 1946 10740 1978 10774
rect 2016 10740 2048 10774
rect 2048 10740 2050 10774
rect 1944 10667 1946 10701
rect 1946 10667 1978 10701
rect 2016 10667 2048 10701
rect 2048 10667 2050 10701
rect 1944 8938 1946 10628
rect 1946 8938 2048 10628
rect 2048 9699 2050 10628
rect 2348 39107 2382 39141
rect 2420 39108 2439 39141
rect 2439 39108 2454 39141
rect 2420 39107 2454 39108
rect 2492 39107 2526 39141
rect 2564 39107 2598 39141
rect 2636 39107 2670 39141
rect 2708 39107 2742 39141
rect 2780 39107 2814 39141
rect 2852 39107 2886 39141
rect 2924 39107 2958 39141
rect 2996 39107 3030 39141
rect 3068 39107 3102 39141
rect 3140 39107 3174 39141
rect 3212 39107 3246 39141
rect 3284 39107 3318 39141
rect 3356 39107 3390 39141
rect 3428 39107 3462 39141
rect 3500 39107 3534 39141
rect 3572 39107 3606 39141
rect 3644 39107 3678 39141
rect 3716 39107 3750 39141
rect 3788 39107 3822 39141
rect 3860 39107 3894 39141
rect 3932 39107 3966 39141
rect 4004 39107 4038 39141
rect 4076 39107 4110 39141
rect 4148 39107 4182 39141
rect 4220 39107 4254 39141
rect 4292 39107 4326 39141
rect 4364 39107 4398 39141
rect 4436 39107 4470 39141
rect 4508 39107 4542 39141
rect 4580 39107 4614 39141
rect 4652 39107 4686 39141
rect 4724 39107 4758 39141
rect 4796 39107 4830 39141
rect 4868 39107 4902 39141
rect 4940 39107 4974 39141
rect 5012 39107 5046 39141
rect 5084 39107 5118 39141
rect 5156 39107 5190 39141
rect 5228 39107 5262 39141
rect 5300 39107 5334 39141
rect 5372 39107 5406 39141
rect 5444 39107 5478 39141
rect 5516 39107 5550 39141
rect 5588 39107 5622 39141
rect 5660 39107 5694 39141
rect 5732 39107 5766 39141
rect 5804 39107 5838 39141
rect 5877 39107 5911 39141
rect 5950 39107 5984 39141
rect 6023 39107 6057 39141
rect 6096 39107 6130 39141
rect 6169 39107 6203 39141
rect 6242 39107 6276 39141
rect 6315 39107 6349 39141
rect 6388 39107 6422 39141
rect 6461 39107 6495 39141
rect 6534 39107 6568 39141
rect 6607 39107 6641 39141
rect 6680 39107 6714 39141
rect 6753 39107 6787 39141
rect 6826 39107 6860 39141
rect 6963 39107 6997 39141
rect 7039 39107 7073 39141
rect 7115 39107 7149 39141
rect 7191 39107 7225 39141
rect 7267 39107 7301 39141
rect 7343 39107 7377 39141
rect 7419 39107 7453 39141
rect 7496 39107 7530 39141
rect 7573 39107 7607 39141
rect 7650 39107 7684 39141
rect 7727 39107 7761 39141
rect 7804 39107 7838 39141
rect 7881 39107 7915 39141
rect 7958 39107 7992 39141
rect 8035 39107 8069 39141
rect 8112 39107 8146 39141
rect 2276 39035 2310 39069
rect 8184 39035 8218 39069
rect 2410 39006 2444 39007
rect 2276 38962 2310 38996
rect 2410 38973 2444 39006
rect 2482 38973 2516 39007
rect 2554 38973 2588 39007
rect 2626 38973 2660 39007
rect 2698 38973 2732 39007
rect 2770 38973 2804 39007
rect 2842 38973 2876 39007
rect 2914 38973 2948 39007
rect 2986 38973 3020 39007
rect 3058 38973 3092 39007
rect 3130 38973 3164 39007
rect 3202 38973 3236 39007
rect 3274 38973 3308 39007
rect 3346 38973 3380 39007
rect 3418 38973 3452 39007
rect 3490 38973 3524 39007
rect 3562 38973 3596 39007
rect 3634 38973 3668 39007
rect 3706 38973 3740 39007
rect 3778 38973 3812 39007
rect 3850 38973 3884 39007
rect 3922 38973 3956 39007
rect 3994 38973 4028 39007
rect 4066 38973 4100 39007
rect 4138 38973 4172 39007
rect 4210 38973 4244 39007
rect 4282 38973 4316 39007
rect 4354 38973 4388 39007
rect 4426 38973 4460 39007
rect 4498 38973 4532 39007
rect 4570 38973 4604 39007
rect 4642 38973 4676 39007
rect 4714 38973 4748 39007
rect 4786 38973 4820 39007
rect 4858 38973 4892 39007
rect 4930 38973 4964 39007
rect 5002 38973 5036 39007
rect 5074 38973 5108 39007
rect 5147 38973 5181 39007
rect 5220 38973 5254 39007
rect 5293 38973 5327 39007
rect 5366 38973 5400 39007
rect 5439 38973 5473 39007
rect 5512 38973 5546 39007
rect 5585 38973 5619 39007
rect 5658 38973 5692 39007
rect 5731 38973 5765 39007
rect 5804 38973 5838 39007
rect 5877 38973 5911 39007
rect 5950 38973 5984 39007
rect 6023 38973 6057 39007
rect 6096 38973 6130 39007
rect 6169 38973 6203 39007
rect 6242 38973 6276 39007
rect 6315 38973 6349 39007
rect 6388 38973 6422 39007
rect 6461 38973 6495 39007
rect 6534 38973 6568 39007
rect 6607 38973 6641 39007
rect 6680 38973 6714 39007
rect 6753 38973 6787 39007
rect 6826 38973 6860 39007
rect 6963 38973 6997 39007
rect 7035 38973 7069 39007
rect 7107 38973 7141 39007
rect 7179 38973 7213 39007
rect 7251 38973 7285 39007
rect 7323 38973 7357 39007
rect 7395 38973 7429 39007
rect 7467 38973 7501 39007
rect 7539 38973 7573 39007
rect 7612 38973 7646 39007
rect 7685 38973 7719 39007
rect 7758 38973 7792 39007
rect 7831 38973 7865 39007
rect 7904 38973 7938 39007
rect 7977 38973 8011 39007
rect 8050 38973 8083 39007
rect 8083 38973 8084 39007
rect 8184 38989 8185 38997
rect 8185 38989 8218 38997
rect 2276 38889 2310 38923
rect 2410 38900 2444 38934
rect 2276 38816 2310 38850
rect 2410 38827 2444 38861
rect 8184 38963 8218 38989
rect 8050 38901 8084 38935
rect 8184 38891 8218 38925
rect 3035 38820 3039 38854
rect 3039 38820 3069 38854
rect 3108 38820 3142 38854
rect 3181 38820 3211 38854
rect 3211 38820 3215 38854
rect 3254 38820 3280 38854
rect 3280 38820 3288 38854
rect 3327 38820 3349 38854
rect 3349 38820 3361 38854
rect 3400 38820 3418 38854
rect 3418 38820 3434 38854
rect 3473 38820 3487 38854
rect 3487 38820 3507 38854
rect 3546 38820 3556 38854
rect 3556 38820 3580 38854
rect 3619 38820 3625 38854
rect 3625 38820 3653 38854
rect 3692 38820 3694 38854
rect 3694 38820 3726 38854
rect 3765 38820 3798 38854
rect 3798 38820 3799 38854
rect 3838 38820 3867 38854
rect 3867 38820 3872 38854
rect 3911 38820 3936 38854
rect 3936 38820 3945 38854
rect 3984 38820 4005 38854
rect 4005 38820 4018 38854
rect 4057 38820 4074 38854
rect 4074 38820 4091 38854
rect 4130 38820 4143 38854
rect 4143 38820 4164 38854
rect 4203 38820 4211 38854
rect 4211 38820 4237 38854
rect 4276 38820 4279 38854
rect 4279 38820 4310 38854
rect 4349 38820 4381 38854
rect 4381 38820 4383 38854
rect 4422 38820 4449 38854
rect 4449 38820 4456 38854
rect 4495 38820 4517 38854
rect 4517 38820 4529 38854
rect 4568 38820 4585 38854
rect 4585 38820 4602 38854
rect 4641 38820 4653 38854
rect 4653 38820 4675 38854
rect 4714 38820 4721 38854
rect 4721 38820 4748 38854
rect 4787 38820 4789 38854
rect 4789 38820 4821 38854
rect 4860 38820 4891 38854
rect 4891 38820 4894 38854
rect 4933 38820 4959 38854
rect 4959 38820 4967 38854
rect 5006 38820 5027 38854
rect 5027 38820 5040 38854
rect 5079 38820 5095 38854
rect 5095 38820 5113 38854
rect 5152 38820 5163 38854
rect 5163 38820 5186 38854
rect 5225 38820 5231 38854
rect 5231 38820 5259 38854
rect 5298 38820 5299 38854
rect 5299 38820 5332 38854
rect 5371 38820 5401 38854
rect 5401 38820 5405 38854
rect 5444 38820 5469 38854
rect 5469 38820 5478 38854
rect 5517 38820 5537 38854
rect 5537 38820 5551 38854
rect 5590 38820 5605 38854
rect 5605 38820 5624 38854
rect 5663 38820 5673 38854
rect 5673 38820 5697 38854
rect 5736 38820 5741 38854
rect 5741 38820 5770 38854
rect 5809 38820 5843 38854
rect 5882 38820 5911 38854
rect 5911 38820 5916 38854
rect 5955 38820 5979 38854
rect 5979 38820 5989 38854
rect 6027 38820 6047 38854
rect 6047 38820 6061 38854
rect 6099 38820 6115 38854
rect 6115 38820 6133 38854
rect 6171 38820 6183 38854
rect 6183 38820 6205 38854
rect 6243 38820 6251 38854
rect 6251 38820 6277 38854
rect 6315 38820 6319 38854
rect 6319 38820 6349 38854
rect 6387 38820 6421 38854
rect 6459 38820 6489 38854
rect 6489 38820 6493 38854
rect 6531 38820 6557 38854
rect 6557 38820 6565 38854
rect 6603 38820 6625 38854
rect 6625 38820 6637 38854
rect 6675 38820 6693 38854
rect 6693 38820 6709 38854
rect 6747 38820 6761 38854
rect 6761 38820 6781 38854
rect 6819 38820 6829 38854
rect 6829 38820 6853 38854
rect 6891 38820 6897 38854
rect 6897 38820 6925 38854
rect 6963 38820 6965 38854
rect 6965 38820 6997 38854
rect 7035 38820 7067 38854
rect 7067 38820 7069 38854
rect 7107 38820 7135 38854
rect 7135 38820 7141 38854
rect 7179 38820 7203 38854
rect 7203 38820 7213 38854
rect 7251 38820 7271 38854
rect 7271 38820 7285 38854
rect 7323 38820 7339 38854
rect 7339 38820 7357 38854
rect 7395 38820 7407 38854
rect 7407 38820 7429 38854
rect 7467 38820 7475 38854
rect 7475 38820 7501 38854
rect 7539 38820 7543 38854
rect 7543 38820 7573 38854
rect 7611 38820 7645 38854
rect 7683 38820 7713 38854
rect 7713 38820 7717 38854
rect 8050 38829 8084 38863
rect 2276 38743 2310 38777
rect 2410 38754 2444 38788
rect 8184 38819 8218 38853
rect 8050 38757 8084 38791
rect 8184 38747 8218 38781
rect 2276 38670 2310 38704
rect 2410 38681 2444 38715
rect 2276 38597 2310 38631
rect 2410 38608 2444 38642
rect 2276 38524 2310 38558
rect 2410 38535 2444 38569
rect 2276 38451 2310 38485
rect 2410 38462 2444 38496
rect 2276 38378 2310 38412
rect 2410 38389 2444 38423
rect 2276 38305 2310 38339
rect 2410 38316 2444 38350
rect 2276 38232 2310 38266
rect 2410 38243 2444 38277
rect 2276 38159 2310 38193
rect 2410 38170 2444 38204
rect 2276 38086 2310 38120
rect 2410 38097 2444 38131
rect 2276 38013 2310 38047
rect 2410 38024 2444 38058
rect 2276 37940 2310 37974
rect 2410 37951 2444 37985
rect 2276 37867 2310 37901
rect 2410 37878 2444 37912
rect 2276 37794 2310 37828
rect 2410 37805 2444 37839
rect 2276 37721 2310 37755
rect 2410 37732 2444 37766
rect 2276 37648 2310 37682
rect 2410 37659 2444 37693
rect 2276 37575 2310 37609
rect 2410 37586 2444 37620
rect 2276 37502 2310 37536
rect 2410 37513 2444 37547
rect 2276 37429 2310 37463
rect 2410 37440 2444 37474
rect 2276 37356 2310 37390
rect 2410 37367 2444 37401
rect 2830 38680 2864 38714
rect 2902 38680 2936 38714
rect 2830 38607 2864 38641
rect 2902 38607 2936 38641
rect 2830 38534 2864 38568
rect 2902 38534 2936 38568
rect 2830 38461 2864 38495
rect 2902 38461 2936 38495
rect 2830 37380 2936 38422
rect 3107 38680 3141 38714
rect 3179 38680 3213 38714
rect 3107 38607 3141 38641
rect 3179 38607 3213 38641
rect 3107 38534 3141 38568
rect 3179 38534 3213 38568
rect 3107 38461 3141 38495
rect 3179 38461 3213 38495
rect 3107 37380 3213 38422
rect 3384 38680 3418 38714
rect 3456 38680 3490 38714
rect 3384 38607 3418 38641
rect 3456 38607 3490 38641
rect 3384 38534 3418 38568
rect 3456 38534 3490 38568
rect 3384 38461 3418 38495
rect 3456 38461 3490 38495
rect 3384 37380 3490 38422
rect 3661 38680 3695 38714
rect 3733 38680 3767 38714
rect 3661 38607 3695 38641
rect 3733 38607 3767 38641
rect 3661 38534 3695 38568
rect 3733 38534 3767 38568
rect 3661 38461 3695 38495
rect 3733 38461 3767 38495
rect 3661 37380 3767 38422
rect 3938 38680 3972 38714
rect 4010 38680 4044 38714
rect 3938 38607 3972 38641
rect 4010 38607 4044 38641
rect 3938 38534 3972 38568
rect 4010 38534 4044 38568
rect 3938 38461 3972 38495
rect 4010 38461 4044 38495
rect 3938 37380 4044 38422
rect 4215 38680 4249 38714
rect 4287 38680 4321 38714
rect 4215 38607 4249 38641
rect 4287 38607 4321 38641
rect 4215 38534 4249 38568
rect 4287 38534 4321 38568
rect 4215 38461 4249 38495
rect 4287 38461 4321 38495
rect 4215 37380 4321 38422
rect 4492 38680 4526 38714
rect 4564 38680 4598 38714
rect 4492 38607 4526 38641
rect 4564 38607 4598 38641
rect 4492 38534 4526 38568
rect 4564 38534 4598 38568
rect 4492 38461 4526 38495
rect 4564 38461 4598 38495
rect 4492 37380 4598 38422
rect 4769 38680 4803 38714
rect 4841 38680 4875 38714
rect 4769 38607 4803 38641
rect 4841 38607 4875 38641
rect 4769 38534 4803 38568
rect 4841 38534 4875 38568
rect 4769 38461 4803 38495
rect 4841 38461 4875 38495
rect 4769 37380 4875 38422
rect 5046 38680 5080 38714
rect 5118 38680 5152 38714
rect 5046 38607 5080 38641
rect 5118 38607 5152 38641
rect 5046 38534 5080 38568
rect 5118 38534 5152 38568
rect 5046 38461 5080 38495
rect 5118 38461 5152 38495
rect 5046 37380 5152 38422
rect 5323 38680 5357 38714
rect 5395 38680 5429 38714
rect 5323 38607 5357 38641
rect 5395 38607 5429 38641
rect 5323 38534 5357 38568
rect 5395 38534 5429 38568
rect 5323 38461 5357 38495
rect 5395 38461 5429 38495
rect 5323 37380 5429 38422
rect 5600 38680 5634 38714
rect 5672 38680 5706 38714
rect 5600 38607 5634 38641
rect 5672 38607 5706 38641
rect 5600 38534 5634 38568
rect 5672 38534 5706 38568
rect 5600 38461 5634 38495
rect 5672 38461 5706 38495
rect 5600 37380 5706 38422
rect 5877 38680 5911 38714
rect 5949 38680 5983 38714
rect 5877 38607 5911 38641
rect 5949 38607 5983 38641
rect 5877 38534 5911 38568
rect 5949 38534 5983 38568
rect 5877 38461 5911 38495
rect 5949 38461 5983 38495
rect 5877 37380 5983 38422
rect 6154 38680 6188 38714
rect 6226 38680 6260 38714
rect 6154 38607 6188 38641
rect 6226 38607 6260 38641
rect 6154 38534 6188 38568
rect 6226 38534 6260 38568
rect 6154 38461 6188 38495
rect 6226 38461 6260 38495
rect 6154 37380 6260 38422
rect 6431 38680 6465 38714
rect 6503 38680 6537 38714
rect 6431 38607 6465 38641
rect 6503 38607 6537 38641
rect 6431 38534 6465 38568
rect 6503 38534 6537 38568
rect 6431 38461 6465 38495
rect 6503 38461 6537 38495
rect 6431 37380 6537 38422
rect 6708 38680 6742 38714
rect 6780 38680 6814 38714
rect 6708 38607 6742 38641
rect 6780 38607 6814 38641
rect 6708 38534 6742 38568
rect 6780 38534 6814 38568
rect 6708 38461 6742 38495
rect 6780 38461 6814 38495
rect 6708 37380 6814 38422
rect 6985 38680 7019 38714
rect 7057 38680 7091 38714
rect 6985 38607 7019 38641
rect 7057 38607 7091 38641
rect 6985 38534 7019 38568
rect 7057 38534 7091 38568
rect 6985 38461 7019 38495
rect 7057 38461 7091 38495
rect 6985 37380 7091 38422
rect 7262 38680 7296 38714
rect 7334 38680 7368 38714
rect 7262 38607 7296 38641
rect 7334 38607 7368 38641
rect 7262 38534 7296 38568
rect 7334 38534 7368 38568
rect 7262 38461 7296 38495
rect 7334 38461 7368 38495
rect 7262 37380 7368 38422
rect 7539 38680 7573 38714
rect 7611 38680 7645 38714
rect 7539 38607 7573 38641
rect 7611 38607 7645 38641
rect 7539 38534 7573 38568
rect 7611 38534 7645 38568
rect 7539 38461 7573 38495
rect 7611 38461 7645 38495
rect 7539 37380 7645 38422
rect 7816 38680 7850 38714
rect 7888 38680 7922 38714
rect 7816 38607 7850 38641
rect 7888 38607 7922 38641
rect 7816 38534 7850 38568
rect 7888 38534 7922 38568
rect 7816 38461 7850 38495
rect 7888 38461 7922 38495
rect 7816 37380 7922 38422
rect 8050 38685 8084 38719
rect 8184 38675 8218 38709
rect 8050 38613 8084 38647
rect 8184 38603 8218 38637
rect 8050 38541 8084 38575
rect 8184 38531 8218 38565
rect 8050 38469 8084 38503
rect 8184 38459 8218 38493
rect 8050 38397 8084 38431
rect 8184 38387 8218 38421
rect 8050 38325 8084 38359
rect 8184 38315 8218 38349
rect 8050 38253 8084 38287
rect 8184 38243 8218 38277
rect 8050 38181 8084 38215
rect 8184 38171 8218 38205
rect 8050 38109 8084 38143
rect 8184 38099 8218 38133
rect 8050 38037 8084 38071
rect 8184 38027 8218 38061
rect 8050 37965 8084 37999
rect 8184 37955 8218 37989
rect 8050 37893 8084 37927
rect 8184 37883 8218 37917
rect 8050 37821 8084 37855
rect 8184 37811 8218 37845
rect 8050 37749 8084 37783
rect 8184 37739 8218 37773
rect 8050 37677 8084 37711
rect 8184 37667 8218 37701
rect 8050 37605 8084 37639
rect 8184 37595 8218 37629
rect 8050 37533 8084 37567
rect 8184 37523 8218 37557
rect 8050 37461 8084 37495
rect 8184 37451 8218 37485
rect 8050 37389 8084 37423
rect 8184 37379 8218 37413
rect 2276 37283 2310 37317
rect 2410 37294 2444 37328
rect 2276 37210 2310 37244
rect 2410 37221 2444 37255
rect 2276 37137 2310 37171
rect 2410 37148 2444 37182
rect 2276 37064 2310 37098
rect 2410 37075 2444 37109
rect 8050 37317 8084 37351
rect 8184 37307 8218 37341
rect 8050 37245 8084 37279
rect 8184 37235 8218 37269
rect 8050 37173 8084 37207
rect 8184 37163 8218 37197
rect 8050 37101 8084 37135
rect 8184 37091 8218 37125
rect 2276 36991 2310 37025
rect 2410 37002 2444 37036
rect 3035 37031 3039 37065
rect 3039 37031 3069 37065
rect 3108 37031 3142 37065
rect 3181 37031 3211 37065
rect 3211 37031 3215 37065
rect 3254 37031 3280 37065
rect 3280 37031 3288 37065
rect 3327 37031 3349 37065
rect 3349 37031 3361 37065
rect 3400 37031 3418 37065
rect 3418 37031 3434 37065
rect 3473 37031 3487 37065
rect 3487 37031 3507 37065
rect 3546 37031 3556 37065
rect 3556 37031 3580 37065
rect 3619 37031 3625 37065
rect 3625 37031 3653 37065
rect 3692 37031 3694 37065
rect 3694 37031 3726 37065
rect 3765 37031 3798 37065
rect 3798 37031 3799 37065
rect 3838 37031 3867 37065
rect 3867 37031 3872 37065
rect 3911 37031 3936 37065
rect 3936 37031 3945 37065
rect 3984 37031 4005 37065
rect 4005 37031 4018 37065
rect 4057 37031 4074 37065
rect 4074 37031 4091 37065
rect 4130 37031 4143 37065
rect 4143 37031 4164 37065
rect 4203 37031 4211 37065
rect 4211 37031 4237 37065
rect 4276 37031 4279 37065
rect 4279 37031 4310 37065
rect 4349 37031 4381 37065
rect 4381 37031 4383 37065
rect 4422 37031 4449 37065
rect 4449 37031 4456 37065
rect 4495 37031 4517 37065
rect 4517 37031 4529 37065
rect 4568 37031 4585 37065
rect 4585 37031 4602 37065
rect 4641 37031 4653 37065
rect 4653 37031 4675 37065
rect 4714 37031 4721 37065
rect 4721 37031 4748 37065
rect 4787 37031 4789 37065
rect 4789 37031 4821 37065
rect 4860 37031 4891 37065
rect 4891 37031 4894 37065
rect 4933 37031 4959 37065
rect 4959 37031 4967 37065
rect 5006 37031 5027 37065
rect 5027 37031 5040 37065
rect 5079 37031 5095 37065
rect 5095 37031 5113 37065
rect 5152 37031 5163 37065
rect 5163 37031 5186 37065
rect 5225 37031 5231 37065
rect 5231 37031 5259 37065
rect 5298 37031 5299 37065
rect 5299 37031 5332 37065
rect 5371 37031 5401 37065
rect 5401 37031 5405 37065
rect 5444 37031 5469 37065
rect 5469 37031 5478 37065
rect 5517 37031 5537 37065
rect 5537 37031 5551 37065
rect 5590 37031 5605 37065
rect 5605 37031 5624 37065
rect 5663 37031 5673 37065
rect 5673 37031 5697 37065
rect 5736 37031 5741 37065
rect 5741 37031 5770 37065
rect 5809 37031 5843 37065
rect 5882 37031 5911 37065
rect 5911 37031 5916 37065
rect 5955 37031 5979 37065
rect 5979 37031 5989 37065
rect 6027 37031 6047 37065
rect 6047 37031 6061 37065
rect 6099 37031 6115 37065
rect 6115 37031 6133 37065
rect 6171 37031 6183 37065
rect 6183 37031 6205 37065
rect 6243 37031 6251 37065
rect 6251 37031 6277 37065
rect 6315 37031 6319 37065
rect 6319 37031 6349 37065
rect 6387 37031 6421 37065
rect 6459 37031 6489 37065
rect 6489 37031 6493 37065
rect 6531 37031 6557 37065
rect 6557 37031 6565 37065
rect 6603 37031 6625 37065
rect 6625 37031 6637 37065
rect 6675 37031 6693 37065
rect 6693 37031 6709 37065
rect 6747 37031 6761 37065
rect 6761 37031 6781 37065
rect 6819 37031 6829 37065
rect 6829 37031 6853 37065
rect 6891 37031 6897 37065
rect 6897 37031 6925 37065
rect 6963 37031 6965 37065
rect 6965 37031 6997 37065
rect 7035 37031 7067 37065
rect 7067 37031 7069 37065
rect 7107 37031 7135 37065
rect 7135 37031 7141 37065
rect 7179 37031 7203 37065
rect 7203 37031 7213 37065
rect 7251 37031 7271 37065
rect 7271 37031 7285 37065
rect 7323 37031 7339 37065
rect 7339 37031 7357 37065
rect 7395 37031 7407 37065
rect 7407 37031 7429 37065
rect 7467 37031 7475 37065
rect 7475 37031 7501 37065
rect 7539 37031 7543 37065
rect 7543 37031 7573 37065
rect 7611 37031 7645 37065
rect 7683 37031 7713 37065
rect 7713 37031 7717 37065
rect 2276 36918 2310 36952
rect 2410 36929 2444 36963
rect 2276 36845 2310 36879
rect 2410 36856 2444 36890
rect 2276 36772 2310 36806
rect 2410 36783 2444 36817
rect 2276 36699 2310 36733
rect 2410 36710 2444 36744
rect 8050 37029 8084 37063
rect 8184 37019 8218 37053
rect 8050 36957 8084 36991
rect 8184 36947 8218 36981
rect 8050 36885 8084 36919
rect 8184 36875 8218 36909
rect 8050 36813 8084 36847
rect 8184 36803 8218 36837
rect 8050 36741 8084 36775
rect 8184 36731 8218 36765
rect 2276 36626 2310 36660
rect 2410 36637 2444 36671
rect 2276 36554 2310 36588
rect 2410 36564 2444 36598
rect 2276 36482 2310 36516
rect 2410 36491 2444 36525
rect 2276 36410 2310 36444
rect 2410 36418 2444 36452
rect 2276 36338 2310 36372
rect 2410 36345 2444 36379
rect 2276 36266 2310 36300
rect 2410 36272 2444 36306
rect 2276 36194 2310 36228
rect 2410 36199 2444 36233
rect 2276 36122 2310 36156
rect 2410 36126 2444 36160
rect 2276 36050 2310 36084
rect 2410 36053 2444 36087
rect 2276 35978 2310 36012
rect 2410 35980 2444 36014
rect 2276 35906 2310 35940
rect 2410 35907 2444 35941
rect 2276 35834 2310 35868
rect 2410 35834 2444 35868
rect 2276 35762 2310 35796
rect 2410 35762 2444 35796
rect 2276 35690 2310 35724
rect 2410 35690 2444 35724
rect 2276 35618 2310 35652
rect 2410 35618 2444 35652
rect 2276 35546 2310 35580
rect 2410 35546 2444 35580
rect 2276 35474 2310 35508
rect 2410 35474 2444 35508
rect 2276 35402 2310 35436
rect 2410 35402 2444 35436
rect 2830 36680 2864 36714
rect 2902 36680 2936 36714
rect 2830 36607 2864 36641
rect 2902 36607 2936 36641
rect 2830 36534 2864 36568
rect 2902 36534 2936 36568
rect 2830 36461 2864 36495
rect 2902 36461 2936 36495
rect 2830 35380 2936 36422
rect 3107 36680 3141 36714
rect 3179 36680 3213 36714
rect 3107 36607 3141 36641
rect 3179 36607 3213 36641
rect 3107 36534 3141 36568
rect 3179 36534 3213 36568
rect 3107 36461 3141 36495
rect 3179 36461 3213 36495
rect 3107 35380 3213 36422
rect 3384 36680 3418 36714
rect 3456 36680 3490 36714
rect 3384 36607 3418 36641
rect 3456 36607 3490 36641
rect 3384 36534 3418 36568
rect 3456 36534 3490 36568
rect 3384 36461 3418 36495
rect 3456 36461 3490 36495
rect 3384 35380 3490 36422
rect 3661 36680 3695 36714
rect 3733 36680 3767 36714
rect 3661 36607 3695 36641
rect 3733 36607 3767 36641
rect 3661 36534 3695 36568
rect 3733 36534 3767 36568
rect 3661 36461 3695 36495
rect 3733 36461 3767 36495
rect 3661 35380 3767 36422
rect 3938 36680 3972 36714
rect 4010 36680 4044 36714
rect 3938 36607 3972 36641
rect 4010 36607 4044 36641
rect 3938 36534 3972 36568
rect 4010 36534 4044 36568
rect 3938 36461 3972 36495
rect 4010 36461 4044 36495
rect 3938 35380 4044 36422
rect 4215 36680 4249 36714
rect 4287 36680 4321 36714
rect 4215 36607 4249 36641
rect 4287 36607 4321 36641
rect 4215 36534 4249 36568
rect 4287 36534 4321 36568
rect 4215 36461 4249 36495
rect 4287 36461 4321 36495
rect 4215 35380 4321 36422
rect 4492 36680 4526 36714
rect 4564 36680 4598 36714
rect 4492 36607 4526 36641
rect 4564 36607 4598 36641
rect 4492 36534 4526 36568
rect 4564 36534 4598 36568
rect 4492 36461 4526 36495
rect 4564 36461 4598 36495
rect 4492 35380 4598 36422
rect 4769 36680 4803 36714
rect 4841 36680 4875 36714
rect 4769 36607 4803 36641
rect 4841 36607 4875 36641
rect 4769 36534 4803 36568
rect 4841 36534 4875 36568
rect 4769 36461 4803 36495
rect 4841 36461 4875 36495
rect 4769 35380 4875 36422
rect 5046 36680 5080 36714
rect 5118 36680 5152 36714
rect 5046 36607 5080 36641
rect 5118 36607 5152 36641
rect 5046 36534 5080 36568
rect 5118 36534 5152 36568
rect 5046 36461 5080 36495
rect 5118 36461 5152 36495
rect 5046 35380 5152 36422
rect 5323 36680 5357 36714
rect 5395 36680 5429 36714
rect 5323 36607 5357 36641
rect 5395 36607 5429 36641
rect 5323 36534 5357 36568
rect 5395 36534 5429 36568
rect 5323 36461 5357 36495
rect 5395 36461 5429 36495
rect 5323 35380 5429 36422
rect 5600 36680 5634 36714
rect 5672 36680 5706 36714
rect 5600 36607 5634 36641
rect 5672 36607 5706 36641
rect 5600 36534 5634 36568
rect 5672 36534 5706 36568
rect 5600 36461 5634 36495
rect 5672 36461 5706 36495
rect 5600 35380 5706 36422
rect 5877 36680 5911 36714
rect 5949 36680 5983 36714
rect 5877 36607 5911 36641
rect 5949 36607 5983 36641
rect 5877 36534 5911 36568
rect 5949 36534 5983 36568
rect 5877 36461 5911 36495
rect 5949 36461 5983 36495
rect 5877 35380 5983 36422
rect 6154 36680 6188 36714
rect 6226 36680 6260 36714
rect 6154 36607 6188 36641
rect 6226 36607 6260 36641
rect 6154 36534 6188 36568
rect 6226 36534 6260 36568
rect 6154 36461 6188 36495
rect 6226 36461 6260 36495
rect 6154 35380 6260 36422
rect 6431 36680 6465 36714
rect 6503 36680 6537 36714
rect 6431 36607 6465 36641
rect 6503 36607 6537 36641
rect 6431 36534 6465 36568
rect 6503 36534 6537 36568
rect 6431 36461 6465 36495
rect 6503 36461 6537 36495
rect 6431 35380 6537 36422
rect 6708 36680 6742 36714
rect 6780 36680 6814 36714
rect 6708 36607 6742 36641
rect 6780 36607 6814 36641
rect 6708 36534 6742 36568
rect 6780 36534 6814 36568
rect 6708 36461 6742 36495
rect 6780 36461 6814 36495
rect 6708 35380 6814 36422
rect 6985 36680 7019 36714
rect 7057 36680 7091 36714
rect 6985 36607 7019 36641
rect 7057 36607 7091 36641
rect 6985 36534 7019 36568
rect 7057 36534 7091 36568
rect 6985 36461 7019 36495
rect 7057 36461 7091 36495
rect 6985 35380 7091 36422
rect 7262 36680 7296 36714
rect 7334 36680 7368 36714
rect 7262 36607 7296 36641
rect 7334 36607 7368 36641
rect 7262 36534 7296 36568
rect 7334 36534 7368 36568
rect 7262 36461 7296 36495
rect 7334 36461 7368 36495
rect 7262 35380 7368 36422
rect 7539 36680 7573 36714
rect 7611 36680 7645 36714
rect 7539 36607 7573 36641
rect 7611 36607 7645 36641
rect 7539 36534 7573 36568
rect 7611 36534 7645 36568
rect 7539 36461 7573 36495
rect 7611 36461 7645 36495
rect 7539 35380 7645 36422
rect 7816 36680 7850 36714
rect 7888 36680 7922 36714
rect 7816 36607 7850 36641
rect 7888 36607 7922 36641
rect 7816 36534 7850 36568
rect 7888 36534 7922 36568
rect 7816 36461 7850 36495
rect 7888 36461 7922 36495
rect 7816 35380 7922 36422
rect 8050 36669 8084 36703
rect 8184 36659 8218 36693
rect 8050 36597 8084 36631
rect 8184 36587 8218 36621
rect 8050 36525 8084 36559
rect 8184 36515 8218 36549
rect 8050 36453 8084 36487
rect 8184 36443 8218 36477
rect 8050 36381 8084 36415
rect 8184 36371 8218 36405
rect 8050 36309 8084 36343
rect 8184 36299 8218 36333
rect 8050 36237 8084 36271
rect 8184 36227 8218 36261
rect 8050 36165 8084 36199
rect 8184 36155 8218 36189
rect 8050 36093 8084 36127
rect 8184 36083 8218 36117
rect 8050 36021 8084 36055
rect 8184 36011 8218 36045
rect 8050 35949 8084 35983
rect 8184 35939 8218 35973
rect 8050 35877 8084 35911
rect 8184 35867 8218 35901
rect 8050 35805 8084 35839
rect 8184 35795 8218 35829
rect 8050 35733 8084 35767
rect 8184 35723 8218 35757
rect 8050 35661 8084 35695
rect 8184 35651 8218 35685
rect 8050 35589 8084 35623
rect 8184 35579 8218 35613
rect 8050 35517 8084 35551
rect 8184 35507 8218 35541
rect 8050 35445 8084 35479
rect 8184 35435 8218 35469
rect 8050 35373 8084 35407
rect 2276 35330 2310 35364
rect 2410 35330 2444 35364
rect 2276 35258 2310 35292
rect 2410 35258 2444 35292
rect 2276 35186 2310 35220
rect 2410 35186 2444 35220
rect 2276 35114 2310 35148
rect 2410 35114 2444 35148
rect 8184 35363 8218 35397
rect 8050 35301 8084 35335
rect 8184 35291 8218 35325
rect 8050 35229 8084 35263
rect 8184 35219 8218 35253
rect 8050 35157 8084 35191
rect 8184 35147 8218 35181
rect 2276 35042 2310 35076
rect 2410 35042 2444 35076
rect 3035 35065 3039 35099
rect 3039 35065 3069 35099
rect 3108 35065 3142 35099
rect 3181 35065 3211 35099
rect 3211 35065 3215 35099
rect 3254 35065 3280 35099
rect 3280 35065 3288 35099
rect 3327 35065 3349 35099
rect 3349 35065 3361 35099
rect 3400 35065 3418 35099
rect 3418 35065 3434 35099
rect 3473 35065 3487 35099
rect 3487 35065 3507 35099
rect 3546 35065 3556 35099
rect 3556 35065 3580 35099
rect 3619 35065 3625 35099
rect 3625 35065 3653 35099
rect 3692 35065 3694 35099
rect 3694 35065 3726 35099
rect 3765 35065 3798 35099
rect 3798 35065 3799 35099
rect 3838 35065 3867 35099
rect 3867 35065 3872 35099
rect 3911 35065 3936 35099
rect 3936 35065 3945 35099
rect 3984 35065 4005 35099
rect 4005 35065 4018 35099
rect 4057 35065 4074 35099
rect 4074 35065 4091 35099
rect 4130 35065 4143 35099
rect 4143 35065 4164 35099
rect 4203 35065 4211 35099
rect 4211 35065 4237 35099
rect 4276 35065 4279 35099
rect 4279 35065 4310 35099
rect 4349 35065 4381 35099
rect 4381 35065 4383 35099
rect 4422 35065 4449 35099
rect 4449 35065 4456 35099
rect 4495 35065 4517 35099
rect 4517 35065 4529 35099
rect 4568 35065 4585 35099
rect 4585 35065 4602 35099
rect 4641 35065 4653 35099
rect 4653 35065 4675 35099
rect 4714 35065 4721 35099
rect 4721 35065 4748 35099
rect 4787 35065 4789 35099
rect 4789 35065 4821 35099
rect 4860 35065 4891 35099
rect 4891 35065 4894 35099
rect 4933 35065 4959 35099
rect 4959 35065 4967 35099
rect 5006 35065 5027 35099
rect 5027 35065 5040 35099
rect 5079 35065 5095 35099
rect 5095 35065 5113 35099
rect 5152 35065 5163 35099
rect 5163 35065 5186 35099
rect 5225 35065 5231 35099
rect 5231 35065 5259 35099
rect 5298 35065 5299 35099
rect 5299 35065 5332 35099
rect 5371 35065 5401 35099
rect 5401 35065 5405 35099
rect 5444 35065 5469 35099
rect 5469 35065 5478 35099
rect 5517 35065 5537 35099
rect 5537 35065 5551 35099
rect 5590 35065 5605 35099
rect 5605 35065 5624 35099
rect 5663 35065 5673 35099
rect 5673 35065 5697 35099
rect 5736 35065 5741 35099
rect 5741 35065 5770 35099
rect 5809 35065 5843 35099
rect 5882 35065 5911 35099
rect 5911 35065 5916 35099
rect 5955 35065 5979 35099
rect 5979 35065 5989 35099
rect 6027 35065 6047 35099
rect 6047 35065 6061 35099
rect 6099 35065 6115 35099
rect 6115 35065 6133 35099
rect 6171 35065 6183 35099
rect 6183 35065 6205 35099
rect 6243 35065 6251 35099
rect 6251 35065 6277 35099
rect 6315 35065 6319 35099
rect 6319 35065 6349 35099
rect 6387 35065 6421 35099
rect 6459 35065 6489 35099
rect 6489 35065 6493 35099
rect 6531 35065 6557 35099
rect 6557 35065 6565 35099
rect 6603 35065 6625 35099
rect 6625 35065 6637 35099
rect 6675 35065 6693 35099
rect 6693 35065 6709 35099
rect 6747 35065 6761 35099
rect 6761 35065 6781 35099
rect 6819 35065 6829 35099
rect 6829 35065 6853 35099
rect 6891 35065 6897 35099
rect 6897 35065 6925 35099
rect 6963 35065 6965 35099
rect 6965 35065 6997 35099
rect 7035 35065 7067 35099
rect 7067 35065 7069 35099
rect 7107 35065 7135 35099
rect 7135 35065 7141 35099
rect 7179 35065 7203 35099
rect 7203 35065 7213 35099
rect 7251 35065 7271 35099
rect 7271 35065 7285 35099
rect 7323 35065 7339 35099
rect 7339 35065 7357 35099
rect 7395 35065 7407 35099
rect 7407 35065 7429 35099
rect 7467 35065 7475 35099
rect 7475 35065 7501 35099
rect 7539 35065 7543 35099
rect 7543 35065 7573 35099
rect 7611 35065 7645 35099
rect 7683 35065 7713 35099
rect 7713 35065 7717 35099
rect 8050 35085 8084 35119
rect 8184 35075 8218 35109
rect 2276 34970 2310 35004
rect 2410 34970 2444 35004
rect 2276 34898 2310 34932
rect 2410 34898 2444 34932
rect 2276 34826 2310 34860
rect 2410 34826 2444 34860
rect 2276 34754 2310 34788
rect 2410 34754 2444 34788
rect 8050 35013 8084 35047
rect 8184 35003 8218 35037
rect 8050 34941 8084 34975
rect 8184 34931 8218 34965
rect 8050 34869 8084 34903
rect 8184 34859 8218 34893
rect 8050 34797 8084 34831
rect 8184 34787 8218 34821
rect 2276 34682 2310 34716
rect 2410 34682 2444 34716
rect 8050 34725 8084 34759
rect 8184 34715 8218 34749
rect 2276 34610 2310 34644
rect 2410 34610 2444 34644
rect 2276 34538 2310 34572
rect 2410 34538 2444 34572
rect 2276 34466 2310 34500
rect 2410 34466 2444 34500
rect 2276 34394 2310 34428
rect 2410 34394 2444 34428
rect 2276 34322 2310 34356
rect 2410 34322 2444 34356
rect 2276 34250 2310 34284
rect 2410 34250 2444 34284
rect 2276 34178 2310 34212
rect 2410 34178 2444 34212
rect 2276 34106 2310 34140
rect 2410 34106 2444 34140
rect 2276 34034 2310 34068
rect 2410 34034 2444 34068
rect 2276 33962 2310 33996
rect 2410 33962 2444 33996
rect 2276 33890 2310 33924
rect 2410 33890 2444 33924
rect 2276 33818 2310 33852
rect 2410 33818 2444 33852
rect 2276 33746 2310 33780
rect 2410 33746 2444 33780
rect 2276 33674 2310 33708
rect 2410 33674 2444 33708
rect 2276 33602 2310 33636
rect 2410 33602 2444 33636
rect 2276 33530 2310 33564
rect 2410 33530 2444 33564
rect 2276 33458 2310 33492
rect 2410 33458 2444 33492
rect 2276 33386 2310 33420
rect 2410 33386 2444 33420
rect 2830 34680 2864 34714
rect 2902 34680 2936 34714
rect 2830 34607 2864 34641
rect 2902 34607 2936 34641
rect 2830 34534 2864 34568
rect 2902 34534 2936 34568
rect 2830 34461 2864 34495
rect 2902 34461 2936 34495
rect 2830 33380 2936 34422
rect 3107 34680 3141 34714
rect 3179 34680 3213 34714
rect 3107 34607 3141 34641
rect 3179 34607 3213 34641
rect 3107 34534 3141 34568
rect 3179 34534 3213 34568
rect 3107 34461 3141 34495
rect 3179 34461 3213 34495
rect 3107 33380 3213 34422
rect 3384 34680 3418 34714
rect 3456 34680 3490 34714
rect 3384 34607 3418 34641
rect 3456 34607 3490 34641
rect 3384 34534 3418 34568
rect 3456 34534 3490 34568
rect 3384 34461 3418 34495
rect 3456 34461 3490 34495
rect 3384 33380 3490 34422
rect 3661 34680 3695 34714
rect 3733 34680 3767 34714
rect 3661 34607 3695 34641
rect 3733 34607 3767 34641
rect 3661 34534 3695 34568
rect 3733 34534 3767 34568
rect 3661 34461 3695 34495
rect 3733 34461 3767 34495
rect 3661 33380 3767 34422
rect 3938 34680 3972 34714
rect 4010 34680 4044 34714
rect 3938 34607 3972 34641
rect 4010 34607 4044 34641
rect 3938 34534 3972 34568
rect 4010 34534 4044 34568
rect 3938 34461 3972 34495
rect 4010 34461 4044 34495
rect 3938 33380 4044 34422
rect 4215 34680 4249 34714
rect 4287 34680 4321 34714
rect 4215 34607 4249 34641
rect 4287 34607 4321 34641
rect 4215 34534 4249 34568
rect 4287 34534 4321 34568
rect 4215 34461 4249 34495
rect 4287 34461 4321 34495
rect 4215 33380 4321 34422
rect 4492 34680 4526 34714
rect 4564 34680 4598 34714
rect 4492 34607 4526 34641
rect 4564 34607 4598 34641
rect 4492 34534 4526 34568
rect 4564 34534 4598 34568
rect 4492 34461 4526 34495
rect 4564 34461 4598 34495
rect 4492 33380 4598 34422
rect 4769 34680 4803 34714
rect 4841 34680 4875 34714
rect 4769 34607 4803 34641
rect 4841 34607 4875 34641
rect 4769 34534 4803 34568
rect 4841 34534 4875 34568
rect 4769 34461 4803 34495
rect 4841 34461 4875 34495
rect 4769 33380 4875 34422
rect 5046 34680 5080 34714
rect 5118 34680 5152 34714
rect 5046 34607 5080 34641
rect 5118 34607 5152 34641
rect 5046 34534 5080 34568
rect 5118 34534 5152 34568
rect 5046 34461 5080 34495
rect 5118 34461 5152 34495
rect 5046 33380 5152 34422
rect 5323 34680 5357 34714
rect 5395 34680 5429 34714
rect 5323 34607 5357 34641
rect 5395 34607 5429 34641
rect 5323 34534 5357 34568
rect 5395 34534 5429 34568
rect 5323 34461 5357 34495
rect 5395 34461 5429 34495
rect 5323 33380 5429 34422
rect 5600 34680 5634 34714
rect 5672 34680 5706 34714
rect 5600 34607 5634 34641
rect 5672 34607 5706 34641
rect 5600 34534 5634 34568
rect 5672 34534 5706 34568
rect 5600 34461 5634 34495
rect 5672 34461 5706 34495
rect 5600 33380 5706 34422
rect 5877 34680 5911 34714
rect 5949 34680 5983 34714
rect 5877 34607 5911 34641
rect 5949 34607 5983 34641
rect 5877 34534 5911 34568
rect 5949 34534 5983 34568
rect 5877 34461 5911 34495
rect 5949 34461 5983 34495
rect 5877 33380 5983 34422
rect 6154 34680 6188 34714
rect 6226 34680 6260 34714
rect 6154 34607 6188 34641
rect 6226 34607 6260 34641
rect 6154 34534 6188 34568
rect 6226 34534 6260 34568
rect 6154 34461 6188 34495
rect 6226 34461 6260 34495
rect 6154 33380 6260 34422
rect 6431 34680 6465 34714
rect 6503 34680 6537 34714
rect 6431 34607 6465 34641
rect 6503 34607 6537 34641
rect 6431 34534 6465 34568
rect 6503 34534 6537 34568
rect 6431 34461 6465 34495
rect 6503 34461 6537 34495
rect 6431 33380 6537 34422
rect 6708 34680 6742 34714
rect 6780 34680 6814 34714
rect 6708 34607 6742 34641
rect 6780 34607 6814 34641
rect 6708 34534 6742 34568
rect 6780 34534 6814 34568
rect 6708 34461 6742 34495
rect 6780 34461 6814 34495
rect 6708 33380 6814 34422
rect 6985 34680 7019 34714
rect 7057 34680 7091 34714
rect 6985 34607 7019 34641
rect 7057 34607 7091 34641
rect 6985 34534 7019 34568
rect 7057 34534 7091 34568
rect 6985 34461 7019 34495
rect 7057 34461 7091 34495
rect 6985 33380 7091 34422
rect 7262 34680 7296 34714
rect 7334 34680 7368 34714
rect 7262 34607 7296 34641
rect 7334 34607 7368 34641
rect 7262 34534 7296 34568
rect 7334 34534 7368 34568
rect 7262 34461 7296 34495
rect 7334 34461 7368 34495
rect 7262 33380 7368 34422
rect 7539 34680 7573 34714
rect 7611 34680 7645 34714
rect 7539 34607 7573 34641
rect 7611 34607 7645 34641
rect 7539 34534 7573 34568
rect 7611 34534 7645 34568
rect 7539 34461 7573 34495
rect 7611 34461 7645 34495
rect 7539 33380 7645 34422
rect 7816 34680 7850 34714
rect 7888 34680 7922 34714
rect 7816 34607 7850 34641
rect 7888 34607 7922 34641
rect 7816 34534 7850 34568
rect 7888 34534 7922 34568
rect 7816 34461 7850 34495
rect 7888 34461 7922 34495
rect 7816 33380 7922 34422
rect 8050 34653 8084 34687
rect 8184 34643 8218 34677
rect 8050 34581 8084 34615
rect 8184 34571 8218 34605
rect 8050 34509 8084 34543
rect 8184 34499 8218 34533
rect 8050 34437 8084 34471
rect 8184 34427 8218 34461
rect 8050 34365 8084 34399
rect 8184 34355 8218 34389
rect 8050 34293 8084 34327
rect 8184 34283 8218 34317
rect 8050 34221 8084 34255
rect 8184 34211 8218 34245
rect 8050 34149 8084 34183
rect 8184 34139 8218 34173
rect 8050 34077 8084 34111
rect 8184 34067 8218 34101
rect 8050 34005 8084 34039
rect 8184 33995 8218 34029
rect 8050 33933 8084 33967
rect 8184 33923 8218 33957
rect 8050 33861 8084 33895
rect 8184 33851 8218 33885
rect 8050 33789 8084 33823
rect 8184 33779 8218 33813
rect 8050 33717 8084 33751
rect 8184 33707 8218 33741
rect 8050 33645 8084 33679
rect 8184 33635 8218 33669
rect 8050 33573 8084 33607
rect 8184 33563 8218 33597
rect 8050 33501 8084 33535
rect 8184 33491 8218 33525
rect 8050 33429 8084 33463
rect 8184 33419 8218 33453
rect 2276 33314 2310 33348
rect 2410 33314 2444 33348
rect 2276 33242 2310 33276
rect 2410 33242 2444 33276
rect 2276 33170 2310 33204
rect 2410 33170 2444 33204
rect 2276 33098 2310 33132
rect 2410 33098 2444 33132
rect 8050 33357 8084 33391
rect 8184 33347 8218 33381
rect 8050 33285 8084 33319
rect 8184 33275 8218 33309
rect 8050 33213 8084 33247
rect 8184 33203 8218 33237
rect 8050 33141 8084 33175
rect 8184 33131 8218 33165
rect 3035 33066 3039 33100
rect 3039 33066 3069 33100
rect 3108 33066 3142 33100
rect 3181 33066 3211 33100
rect 3211 33066 3215 33100
rect 3254 33066 3280 33100
rect 3280 33066 3288 33100
rect 3327 33066 3349 33100
rect 3349 33066 3361 33100
rect 3400 33066 3418 33100
rect 3418 33066 3434 33100
rect 3473 33066 3487 33100
rect 3487 33066 3507 33100
rect 3546 33066 3556 33100
rect 3556 33066 3580 33100
rect 3619 33066 3625 33100
rect 3625 33066 3653 33100
rect 3692 33066 3694 33100
rect 3694 33066 3726 33100
rect 3765 33066 3798 33100
rect 3798 33066 3799 33100
rect 3838 33066 3867 33100
rect 3867 33066 3872 33100
rect 3911 33066 3936 33100
rect 3936 33066 3945 33100
rect 3984 33066 4005 33100
rect 4005 33066 4018 33100
rect 4057 33066 4074 33100
rect 4074 33066 4091 33100
rect 4130 33066 4143 33100
rect 4143 33066 4164 33100
rect 4203 33066 4211 33100
rect 4211 33066 4237 33100
rect 4276 33066 4279 33100
rect 4279 33066 4310 33100
rect 4349 33066 4381 33100
rect 4381 33066 4383 33100
rect 4422 33066 4449 33100
rect 4449 33066 4456 33100
rect 4495 33066 4517 33100
rect 4517 33066 4529 33100
rect 4568 33066 4585 33100
rect 4585 33066 4602 33100
rect 4641 33066 4653 33100
rect 4653 33066 4675 33100
rect 4714 33066 4721 33100
rect 4721 33066 4748 33100
rect 4787 33066 4789 33100
rect 4789 33066 4821 33100
rect 4860 33066 4891 33100
rect 4891 33066 4894 33100
rect 4933 33066 4959 33100
rect 4959 33066 4967 33100
rect 5006 33066 5027 33100
rect 5027 33066 5040 33100
rect 5079 33066 5095 33100
rect 5095 33066 5113 33100
rect 5152 33066 5163 33100
rect 5163 33066 5186 33100
rect 5225 33066 5231 33100
rect 5231 33066 5259 33100
rect 5298 33066 5299 33100
rect 5299 33066 5332 33100
rect 5371 33066 5401 33100
rect 5401 33066 5405 33100
rect 5444 33066 5469 33100
rect 5469 33066 5478 33100
rect 5517 33066 5537 33100
rect 5537 33066 5551 33100
rect 5590 33066 5605 33100
rect 5605 33066 5624 33100
rect 5663 33066 5673 33100
rect 5673 33066 5697 33100
rect 5736 33066 5741 33100
rect 5741 33066 5770 33100
rect 5809 33066 5843 33100
rect 5882 33066 5911 33100
rect 5911 33066 5916 33100
rect 5955 33066 5979 33100
rect 5979 33066 5989 33100
rect 6027 33066 6047 33100
rect 6047 33066 6061 33100
rect 6099 33066 6115 33100
rect 6115 33066 6133 33100
rect 6171 33066 6183 33100
rect 6183 33066 6205 33100
rect 6243 33066 6251 33100
rect 6251 33066 6277 33100
rect 6315 33066 6319 33100
rect 6319 33066 6349 33100
rect 6387 33066 6421 33100
rect 6459 33066 6489 33100
rect 6489 33066 6493 33100
rect 6531 33066 6557 33100
rect 6557 33066 6565 33100
rect 6603 33066 6625 33100
rect 6625 33066 6637 33100
rect 6675 33066 6693 33100
rect 6693 33066 6709 33100
rect 6747 33066 6761 33100
rect 6761 33066 6781 33100
rect 6819 33066 6829 33100
rect 6829 33066 6853 33100
rect 6891 33066 6897 33100
rect 6897 33066 6925 33100
rect 6963 33066 6965 33100
rect 6965 33066 6997 33100
rect 7035 33066 7067 33100
rect 7067 33066 7069 33100
rect 7107 33066 7135 33100
rect 7135 33066 7141 33100
rect 7179 33066 7203 33100
rect 7203 33066 7213 33100
rect 7251 33066 7271 33100
rect 7271 33066 7285 33100
rect 7323 33066 7339 33100
rect 7339 33066 7357 33100
rect 7395 33066 7407 33100
rect 7407 33066 7429 33100
rect 7467 33066 7475 33100
rect 7475 33066 7501 33100
rect 7539 33066 7543 33100
rect 7543 33066 7573 33100
rect 7611 33066 7645 33100
rect 7683 33066 7713 33100
rect 7713 33066 7717 33100
rect 8050 33069 8084 33103
rect 2276 33026 2310 33060
rect 2410 33026 2444 33060
rect 2276 32954 2310 32988
rect 2410 32954 2444 32988
rect 2276 32882 2310 32916
rect 2410 32882 2444 32916
rect 2276 32810 2310 32844
rect 2410 32810 2444 32844
rect 2276 32738 2310 32772
rect 2410 32738 2444 32772
rect 8184 33059 8218 33093
rect 8050 32997 8084 33031
rect 8184 32987 8218 33021
rect 8050 32925 8084 32959
rect 8184 32915 8218 32949
rect 8050 32853 8084 32887
rect 8184 32843 8218 32877
rect 8050 32781 8084 32815
rect 8184 32771 8218 32805
rect 2276 32666 2310 32700
rect 2410 32666 2444 32700
rect 2276 32594 2310 32628
rect 2410 32594 2444 32628
rect 2276 32522 2310 32556
rect 2410 32522 2444 32556
rect 2276 32450 2310 32484
rect 2410 32450 2444 32484
rect 2276 32378 2310 32412
rect 2410 32378 2444 32412
rect 2276 32306 2310 32340
rect 2410 32306 2444 32340
rect 2276 32234 2310 32268
rect 2410 32234 2444 32268
rect 2276 32162 2310 32196
rect 2410 32162 2444 32196
rect 2276 32090 2310 32124
rect 2410 32090 2444 32124
rect 2276 32018 2310 32052
rect 2410 32018 2444 32052
rect 2276 31946 2310 31980
rect 2410 31946 2444 31980
rect 2276 31874 2310 31908
rect 2410 31874 2444 31908
rect 2276 31802 2310 31836
rect 2410 31802 2444 31836
rect 2276 31730 2310 31764
rect 2410 31730 2444 31764
rect 2276 31658 2310 31692
rect 2410 31658 2444 31692
rect 2276 31586 2310 31620
rect 2410 31586 2444 31620
rect 2276 31514 2310 31548
rect 2410 31514 2444 31548
rect 2276 31442 2310 31476
rect 2410 31442 2444 31476
rect 2276 31370 2310 31404
rect 2410 31370 2444 31404
rect 2830 32680 2864 32714
rect 2902 32680 2936 32714
rect 2830 32607 2864 32641
rect 2902 32607 2936 32641
rect 2830 32534 2864 32568
rect 2902 32534 2936 32568
rect 2830 32461 2864 32495
rect 2902 32461 2936 32495
rect 2830 31380 2936 32422
rect 3107 32680 3141 32714
rect 3179 32680 3213 32714
rect 3107 32607 3141 32641
rect 3179 32607 3213 32641
rect 3107 32534 3141 32568
rect 3179 32534 3213 32568
rect 3107 32461 3141 32495
rect 3179 32461 3213 32495
rect 3107 31380 3213 32422
rect 3384 32680 3418 32714
rect 3456 32680 3490 32714
rect 3384 32607 3418 32641
rect 3456 32607 3490 32641
rect 3384 32534 3418 32568
rect 3456 32534 3490 32568
rect 3384 32461 3418 32495
rect 3456 32461 3490 32495
rect 3384 31380 3490 32422
rect 3661 32680 3695 32714
rect 3733 32680 3767 32714
rect 3661 32607 3695 32641
rect 3733 32607 3767 32641
rect 3661 32534 3695 32568
rect 3733 32534 3767 32568
rect 3661 32461 3695 32495
rect 3733 32461 3767 32495
rect 3661 31380 3767 32422
rect 3938 32680 3972 32714
rect 4010 32680 4044 32714
rect 3938 32607 3972 32641
rect 4010 32607 4044 32641
rect 3938 32534 3972 32568
rect 4010 32534 4044 32568
rect 3938 32461 3972 32495
rect 4010 32461 4044 32495
rect 3938 31380 4044 32422
rect 4215 32680 4249 32714
rect 4287 32680 4321 32714
rect 4215 32607 4249 32641
rect 4287 32607 4321 32641
rect 4215 32534 4249 32568
rect 4287 32534 4321 32568
rect 4215 32461 4249 32495
rect 4287 32461 4321 32495
rect 4215 31380 4321 32422
rect 4492 32680 4526 32714
rect 4564 32680 4598 32714
rect 4492 32607 4526 32641
rect 4564 32607 4598 32641
rect 4492 32534 4526 32568
rect 4564 32534 4598 32568
rect 4492 32461 4526 32495
rect 4564 32461 4598 32495
rect 4492 31380 4598 32422
rect 4769 32680 4803 32714
rect 4841 32680 4875 32714
rect 4769 32607 4803 32641
rect 4841 32607 4875 32641
rect 4769 32534 4803 32568
rect 4841 32534 4875 32568
rect 4769 32461 4803 32495
rect 4841 32461 4875 32495
rect 4769 31380 4875 32422
rect 5046 32680 5080 32714
rect 5118 32680 5152 32714
rect 5046 32607 5080 32641
rect 5118 32607 5152 32641
rect 5046 32534 5080 32568
rect 5118 32534 5152 32568
rect 5046 32461 5080 32495
rect 5118 32461 5152 32495
rect 5046 31380 5152 32422
rect 5323 32680 5357 32714
rect 5395 32680 5429 32714
rect 5323 32607 5357 32641
rect 5395 32607 5429 32641
rect 5323 32534 5357 32568
rect 5395 32534 5429 32568
rect 5323 32461 5357 32495
rect 5395 32461 5429 32495
rect 5323 31380 5429 32422
rect 5600 32680 5634 32714
rect 5672 32680 5706 32714
rect 5600 32607 5634 32641
rect 5672 32607 5706 32641
rect 5600 32534 5634 32568
rect 5672 32534 5706 32568
rect 5600 32461 5634 32495
rect 5672 32461 5706 32495
rect 5600 31380 5706 32422
rect 5877 32680 5911 32714
rect 5949 32680 5983 32714
rect 5877 32607 5911 32641
rect 5949 32607 5983 32641
rect 5877 32534 5911 32568
rect 5949 32534 5983 32568
rect 5877 32461 5911 32495
rect 5949 32461 5983 32495
rect 5877 31380 5983 32422
rect 6154 32680 6188 32714
rect 6226 32680 6260 32714
rect 6154 32607 6188 32641
rect 6226 32607 6260 32641
rect 6154 32534 6188 32568
rect 6226 32534 6260 32568
rect 6154 32461 6188 32495
rect 6226 32461 6260 32495
rect 6154 31380 6260 32422
rect 6431 32680 6465 32714
rect 6503 32680 6537 32714
rect 6431 32607 6465 32641
rect 6503 32607 6537 32641
rect 6431 32534 6465 32568
rect 6503 32534 6537 32568
rect 6431 32461 6465 32495
rect 6503 32461 6537 32495
rect 6431 31380 6537 32422
rect 6708 32680 6742 32714
rect 6780 32680 6814 32714
rect 6708 32607 6742 32641
rect 6780 32607 6814 32641
rect 6708 32534 6742 32568
rect 6780 32534 6814 32568
rect 6708 32461 6742 32495
rect 6780 32461 6814 32495
rect 6708 31380 6814 32422
rect 6985 32680 7019 32714
rect 7057 32680 7091 32714
rect 6985 32607 7019 32641
rect 7057 32607 7091 32641
rect 6985 32534 7019 32568
rect 7057 32534 7091 32568
rect 6985 32461 7019 32495
rect 7057 32461 7091 32495
rect 6985 31380 7091 32422
rect 7262 32680 7296 32714
rect 7334 32680 7368 32714
rect 7262 32607 7296 32641
rect 7334 32607 7368 32641
rect 7262 32534 7296 32568
rect 7334 32534 7368 32568
rect 7262 32461 7296 32495
rect 7334 32461 7368 32495
rect 7262 31380 7368 32422
rect 7539 32680 7573 32714
rect 7611 32680 7645 32714
rect 7539 32607 7573 32641
rect 7611 32607 7645 32641
rect 7539 32534 7573 32568
rect 7611 32534 7645 32568
rect 7539 32461 7573 32495
rect 7611 32461 7645 32495
rect 7539 31380 7645 32422
rect 7816 32680 7850 32714
rect 7888 32680 7922 32714
rect 7816 32607 7850 32641
rect 7888 32607 7922 32641
rect 7816 32534 7850 32568
rect 7888 32534 7922 32568
rect 7816 32461 7850 32495
rect 7888 32461 7922 32495
rect 7816 31380 7922 32422
rect 8050 32709 8084 32743
rect 8184 32699 8218 32733
rect 8050 32637 8084 32671
rect 8184 32627 8218 32661
rect 8050 32565 8084 32599
rect 8184 32555 8218 32589
rect 8050 32493 8084 32527
rect 8184 32483 8218 32517
rect 8050 32421 8084 32455
rect 8184 32411 8218 32445
rect 8050 32349 8084 32383
rect 8184 32339 8218 32373
rect 8050 32277 8084 32311
rect 8184 32267 8218 32301
rect 8050 32205 8084 32239
rect 8184 32195 8218 32229
rect 8050 32133 8084 32167
rect 8184 32123 8218 32157
rect 8050 32061 8084 32095
rect 8184 32051 8218 32085
rect 8050 31989 8084 32023
rect 8184 31979 8218 32013
rect 8050 31917 8084 31951
rect 8184 31907 8218 31941
rect 8050 31845 8084 31879
rect 8184 31835 8218 31869
rect 8050 31773 8084 31807
rect 8184 31763 8218 31797
rect 8050 31701 8084 31735
rect 8184 31691 8218 31725
rect 8050 31629 8084 31663
rect 8184 31619 8218 31653
rect 8050 31557 8084 31591
rect 8184 31547 8218 31581
rect 8050 31485 8084 31519
rect 8184 31475 8218 31509
rect 8050 31413 8084 31447
rect 8184 31403 8218 31437
rect 2276 31298 2310 31332
rect 2410 31298 2444 31332
rect 2276 31226 2310 31260
rect 2410 31226 2444 31260
rect 2276 31154 2310 31188
rect 2410 31154 2444 31188
rect 2276 31082 2310 31116
rect 2410 31082 2444 31116
rect 8050 31341 8084 31375
rect 8184 31331 8218 31365
rect 8050 31269 8084 31303
rect 8184 31259 8218 31293
rect 8050 31197 8084 31231
rect 8184 31187 8218 31221
rect 8050 31125 8084 31159
rect 8184 31115 8218 31149
rect 2276 31010 2310 31044
rect 2410 31010 2444 31044
rect 3035 31043 3039 31077
rect 3039 31043 3069 31077
rect 3108 31043 3142 31077
rect 3181 31043 3211 31077
rect 3211 31043 3215 31077
rect 3254 31043 3280 31077
rect 3280 31043 3288 31077
rect 3327 31043 3349 31077
rect 3349 31043 3361 31077
rect 3400 31043 3418 31077
rect 3418 31043 3434 31077
rect 3473 31043 3487 31077
rect 3487 31043 3507 31077
rect 3546 31043 3556 31077
rect 3556 31043 3580 31077
rect 3619 31043 3625 31077
rect 3625 31043 3653 31077
rect 3692 31043 3694 31077
rect 3694 31043 3726 31077
rect 3765 31043 3798 31077
rect 3798 31043 3799 31077
rect 3838 31043 3867 31077
rect 3867 31043 3872 31077
rect 3911 31043 3936 31077
rect 3936 31043 3945 31077
rect 3984 31043 4005 31077
rect 4005 31043 4018 31077
rect 4057 31043 4074 31077
rect 4074 31043 4091 31077
rect 4130 31043 4143 31077
rect 4143 31043 4164 31077
rect 4203 31043 4211 31077
rect 4211 31043 4237 31077
rect 4276 31043 4279 31077
rect 4279 31043 4310 31077
rect 4349 31043 4381 31077
rect 4381 31043 4383 31077
rect 4422 31043 4449 31077
rect 4449 31043 4456 31077
rect 4495 31043 4517 31077
rect 4517 31043 4529 31077
rect 4568 31043 4585 31077
rect 4585 31043 4602 31077
rect 4641 31043 4653 31077
rect 4653 31043 4675 31077
rect 4714 31043 4721 31077
rect 4721 31043 4748 31077
rect 4787 31043 4789 31077
rect 4789 31043 4821 31077
rect 4860 31043 4891 31077
rect 4891 31043 4894 31077
rect 4933 31043 4959 31077
rect 4959 31043 4967 31077
rect 5006 31043 5027 31077
rect 5027 31043 5040 31077
rect 5079 31043 5095 31077
rect 5095 31043 5113 31077
rect 5152 31043 5163 31077
rect 5163 31043 5186 31077
rect 5225 31043 5231 31077
rect 5231 31043 5259 31077
rect 5298 31043 5299 31077
rect 5299 31043 5332 31077
rect 5371 31043 5401 31077
rect 5401 31043 5405 31077
rect 5444 31043 5469 31077
rect 5469 31043 5478 31077
rect 5517 31043 5537 31077
rect 5537 31043 5551 31077
rect 5590 31043 5605 31077
rect 5605 31043 5624 31077
rect 5663 31043 5673 31077
rect 5673 31043 5697 31077
rect 5736 31043 5741 31077
rect 5741 31043 5770 31077
rect 5809 31043 5843 31077
rect 5882 31043 5911 31077
rect 5911 31043 5916 31077
rect 5955 31043 5979 31077
rect 5979 31043 5989 31077
rect 6027 31043 6047 31077
rect 6047 31043 6061 31077
rect 6099 31043 6115 31077
rect 6115 31043 6133 31077
rect 6171 31043 6183 31077
rect 6183 31043 6205 31077
rect 6243 31043 6251 31077
rect 6251 31043 6277 31077
rect 6315 31043 6319 31077
rect 6319 31043 6349 31077
rect 6387 31043 6421 31077
rect 6459 31043 6489 31077
rect 6489 31043 6493 31077
rect 6531 31043 6557 31077
rect 6557 31043 6565 31077
rect 6603 31043 6625 31077
rect 6625 31043 6637 31077
rect 6675 31043 6693 31077
rect 6693 31043 6709 31077
rect 6747 31043 6761 31077
rect 6761 31043 6781 31077
rect 6819 31043 6829 31077
rect 6829 31043 6853 31077
rect 6891 31043 6897 31077
rect 6897 31043 6925 31077
rect 6963 31043 6965 31077
rect 6965 31043 6997 31077
rect 7035 31043 7067 31077
rect 7067 31043 7069 31077
rect 7107 31043 7135 31077
rect 7135 31043 7141 31077
rect 7179 31043 7203 31077
rect 7203 31043 7213 31077
rect 7251 31043 7271 31077
rect 7271 31043 7285 31077
rect 7323 31043 7339 31077
rect 7339 31043 7357 31077
rect 7395 31043 7407 31077
rect 7407 31043 7429 31077
rect 7467 31043 7475 31077
rect 7475 31043 7501 31077
rect 7539 31043 7543 31077
rect 7543 31043 7573 31077
rect 7611 31043 7645 31077
rect 7683 31043 7713 31077
rect 7713 31043 7717 31077
rect 8050 31053 8084 31087
rect 8184 31043 8218 31077
rect 2276 30938 2310 30972
rect 2410 30938 2444 30972
rect 2276 30866 2310 30900
rect 2410 30866 2444 30900
rect 2276 30794 2310 30828
rect 2410 30794 2444 30828
rect 2276 30722 2310 30756
rect 2410 30722 2444 30756
rect 8050 30981 8084 31015
rect 8184 30971 8218 31005
rect 8050 30909 8084 30943
rect 8184 30899 8218 30933
rect 8050 30837 8084 30871
rect 8184 30827 8218 30861
rect 8050 30765 8084 30799
rect 8184 30755 8218 30789
rect 2276 30650 2310 30684
rect 2410 30650 2444 30684
rect 2276 30578 2310 30612
rect 2410 30578 2444 30612
rect 2276 30506 2310 30540
rect 2410 30506 2444 30540
rect 2276 30434 2310 30468
rect 2410 30434 2444 30468
rect 2276 30362 2310 30396
rect 2410 30362 2444 30396
rect 2276 30290 2310 30324
rect 2410 30290 2444 30324
rect 2276 30218 2310 30252
rect 2410 30218 2444 30252
rect 2276 30146 2310 30180
rect 2410 30146 2444 30180
rect 2276 30074 2310 30108
rect 2410 30074 2444 30108
rect 2276 30002 2310 30036
rect 2410 30002 2444 30036
rect 2276 29930 2310 29964
rect 2410 29930 2444 29964
rect 2276 29858 2310 29892
rect 2410 29858 2444 29892
rect 2276 29786 2310 29820
rect 2410 29786 2444 29820
rect 2276 29714 2310 29748
rect 2410 29714 2444 29748
rect 2276 29642 2310 29676
rect 2410 29642 2444 29676
rect 2276 29570 2310 29604
rect 2410 29570 2444 29604
rect 2276 29498 2310 29532
rect 2410 29498 2444 29532
rect 2276 29426 2310 29460
rect 2410 29426 2444 29460
rect 2276 29354 2310 29388
rect 2410 29354 2444 29388
rect 2830 30680 2864 30714
rect 2902 30680 2936 30714
rect 2830 30607 2864 30641
rect 2902 30607 2936 30641
rect 2830 30534 2864 30568
rect 2902 30534 2936 30568
rect 2830 30461 2864 30495
rect 2902 30461 2936 30495
rect 2830 29380 2936 30422
rect 3107 30680 3141 30714
rect 3179 30680 3213 30714
rect 3107 30607 3141 30641
rect 3179 30607 3213 30641
rect 3107 30534 3141 30568
rect 3179 30534 3213 30568
rect 3107 30461 3141 30495
rect 3179 30461 3213 30495
rect 3107 29380 3213 30422
rect 3384 30680 3418 30714
rect 3456 30680 3490 30714
rect 3384 30607 3418 30641
rect 3456 30607 3490 30641
rect 3384 30534 3418 30568
rect 3456 30534 3490 30568
rect 3384 30461 3418 30495
rect 3456 30461 3490 30495
rect 3384 29380 3490 30422
rect 3661 30680 3695 30714
rect 3733 30680 3767 30714
rect 3661 30607 3695 30641
rect 3733 30607 3767 30641
rect 3661 30534 3695 30568
rect 3733 30534 3767 30568
rect 3661 30461 3695 30495
rect 3733 30461 3767 30495
rect 3661 29380 3767 30422
rect 3938 30680 3972 30714
rect 4010 30680 4044 30714
rect 3938 30607 3972 30641
rect 4010 30607 4044 30641
rect 3938 30534 3972 30568
rect 4010 30534 4044 30568
rect 3938 30461 3972 30495
rect 4010 30461 4044 30495
rect 3938 29380 4044 30422
rect 4215 30680 4249 30714
rect 4287 30680 4321 30714
rect 4215 30607 4249 30641
rect 4287 30607 4321 30641
rect 4215 30534 4249 30568
rect 4287 30534 4321 30568
rect 4215 30461 4249 30495
rect 4287 30461 4321 30495
rect 4215 29380 4321 30422
rect 4492 30680 4526 30714
rect 4564 30680 4598 30714
rect 4492 30607 4526 30641
rect 4564 30607 4598 30641
rect 4492 30534 4526 30568
rect 4564 30534 4598 30568
rect 4492 30461 4526 30495
rect 4564 30461 4598 30495
rect 4492 29380 4598 30422
rect 4769 30680 4803 30714
rect 4841 30680 4875 30714
rect 4769 30607 4803 30641
rect 4841 30607 4875 30641
rect 4769 30534 4803 30568
rect 4841 30534 4875 30568
rect 4769 30461 4803 30495
rect 4841 30461 4875 30495
rect 4769 29380 4875 30422
rect 5046 30680 5080 30714
rect 5118 30680 5152 30714
rect 5046 30607 5080 30641
rect 5118 30607 5152 30641
rect 5046 30534 5080 30568
rect 5118 30534 5152 30568
rect 5046 30461 5080 30495
rect 5118 30461 5152 30495
rect 5046 29380 5152 30422
rect 5323 30680 5357 30714
rect 5395 30680 5429 30714
rect 5323 30607 5357 30641
rect 5395 30607 5429 30641
rect 5323 30534 5357 30568
rect 5395 30534 5429 30568
rect 5323 30461 5357 30495
rect 5395 30461 5429 30495
rect 5323 29380 5429 30422
rect 5600 30680 5634 30714
rect 5672 30680 5706 30714
rect 5600 30607 5634 30641
rect 5672 30607 5706 30641
rect 5600 30534 5634 30568
rect 5672 30534 5706 30568
rect 5600 30461 5634 30495
rect 5672 30461 5706 30495
rect 5600 29380 5706 30422
rect 5877 30680 5911 30714
rect 5949 30680 5983 30714
rect 5877 30607 5911 30641
rect 5949 30607 5983 30641
rect 5877 30534 5911 30568
rect 5949 30534 5983 30568
rect 5877 30461 5911 30495
rect 5949 30461 5983 30495
rect 5877 29380 5983 30422
rect 6154 30680 6188 30714
rect 6226 30680 6260 30714
rect 6154 30607 6188 30641
rect 6226 30607 6260 30641
rect 6154 30534 6188 30568
rect 6226 30534 6260 30568
rect 6154 30461 6188 30495
rect 6226 30461 6260 30495
rect 6154 29380 6260 30422
rect 6431 30680 6465 30714
rect 6503 30680 6537 30714
rect 6431 30607 6465 30641
rect 6503 30607 6537 30641
rect 6431 30534 6465 30568
rect 6503 30534 6537 30568
rect 6431 30461 6465 30495
rect 6503 30461 6537 30495
rect 6431 29380 6537 30422
rect 6708 30680 6742 30714
rect 6780 30680 6814 30714
rect 6708 30607 6742 30641
rect 6780 30607 6814 30641
rect 6708 30534 6742 30568
rect 6780 30534 6814 30568
rect 6708 30461 6742 30495
rect 6780 30461 6814 30495
rect 6708 29380 6814 30422
rect 6985 30680 7019 30714
rect 7057 30680 7091 30714
rect 6985 30607 7019 30641
rect 7057 30607 7091 30641
rect 6985 30534 7019 30568
rect 7057 30534 7091 30568
rect 6985 30461 7019 30495
rect 7057 30461 7091 30495
rect 6985 29380 7091 30422
rect 7262 30680 7296 30714
rect 7334 30680 7368 30714
rect 7262 30607 7296 30641
rect 7334 30607 7368 30641
rect 7262 30534 7296 30568
rect 7334 30534 7368 30568
rect 7262 30461 7296 30495
rect 7334 30461 7368 30495
rect 7262 29380 7368 30422
rect 7539 30680 7573 30714
rect 7611 30680 7645 30714
rect 7539 30607 7573 30641
rect 7611 30607 7645 30641
rect 7539 30534 7573 30568
rect 7611 30534 7645 30568
rect 7539 30461 7573 30495
rect 7611 30461 7645 30495
rect 7539 29380 7645 30422
rect 7816 30680 7850 30714
rect 7888 30680 7922 30714
rect 7816 30607 7850 30641
rect 7888 30607 7922 30641
rect 7816 30534 7850 30568
rect 7888 30534 7922 30568
rect 7816 30461 7850 30495
rect 7888 30461 7922 30495
rect 7816 29380 7922 30422
rect 8050 30693 8084 30727
rect 8184 30683 8218 30717
rect 8050 30621 8084 30655
rect 8184 30611 8218 30645
rect 8050 30549 8084 30583
rect 8184 30539 8218 30573
rect 8050 30477 8084 30511
rect 8184 30467 8218 30501
rect 8050 30405 8084 30439
rect 8184 30395 8218 30429
rect 8050 30333 8084 30367
rect 8184 30323 8218 30357
rect 8050 30261 8084 30295
rect 8184 30251 8218 30285
rect 8050 30189 8084 30223
rect 8184 30179 8218 30213
rect 8050 30117 8084 30151
rect 8184 30107 8218 30141
rect 8050 30045 8084 30079
rect 8184 30035 8218 30069
rect 8050 29973 8084 30007
rect 8184 29963 8218 29997
rect 8050 29901 8084 29935
rect 8184 29891 8218 29925
rect 8050 29829 8084 29863
rect 8184 29819 8218 29853
rect 8050 29757 8084 29791
rect 8184 29747 8218 29781
rect 8050 29685 8084 29719
rect 8184 29675 8218 29709
rect 8050 29613 8084 29647
rect 8184 29603 8218 29637
rect 8050 29541 8084 29575
rect 8184 29531 8218 29565
rect 8050 29469 8084 29503
rect 8184 29459 8218 29493
rect 8050 29397 8084 29431
rect 8184 29387 8218 29421
rect 2276 29282 2310 29316
rect 2410 29282 2444 29316
rect 8050 29325 8084 29359
rect 8184 29315 8218 29349
rect 8050 29253 8084 29287
rect 2276 29210 2310 29244
rect 2410 29210 2444 29244
rect 3035 29216 3039 29250
rect 3039 29216 3069 29250
rect 3108 29216 3142 29250
rect 3181 29216 3211 29250
rect 3211 29216 3215 29250
rect 3254 29216 3280 29250
rect 3280 29216 3288 29250
rect 3327 29216 3349 29250
rect 3349 29216 3361 29250
rect 3400 29216 3418 29250
rect 3418 29216 3434 29250
rect 3473 29216 3487 29250
rect 3487 29216 3507 29250
rect 3546 29216 3556 29250
rect 3556 29216 3580 29250
rect 3619 29216 3625 29250
rect 3625 29216 3653 29250
rect 3692 29216 3694 29250
rect 3694 29216 3726 29250
rect 3765 29216 3798 29250
rect 3798 29216 3799 29250
rect 3838 29216 3867 29250
rect 3867 29216 3872 29250
rect 3911 29216 3936 29250
rect 3936 29216 3945 29250
rect 3984 29216 4005 29250
rect 4005 29216 4018 29250
rect 4057 29216 4074 29250
rect 4074 29216 4091 29250
rect 4130 29216 4143 29250
rect 4143 29216 4164 29250
rect 4203 29216 4211 29250
rect 4211 29216 4237 29250
rect 4276 29216 4279 29250
rect 4279 29216 4310 29250
rect 4349 29216 4381 29250
rect 4381 29216 4383 29250
rect 4422 29216 4449 29250
rect 4449 29216 4456 29250
rect 4495 29216 4517 29250
rect 4517 29216 4529 29250
rect 4568 29216 4585 29250
rect 4585 29216 4602 29250
rect 4641 29216 4653 29250
rect 4653 29216 4675 29250
rect 4714 29216 4721 29250
rect 4721 29216 4748 29250
rect 4787 29216 4789 29250
rect 4789 29216 4821 29250
rect 4860 29216 4891 29250
rect 4891 29216 4894 29250
rect 4933 29216 4959 29250
rect 4959 29216 4967 29250
rect 5006 29216 5027 29250
rect 5027 29216 5040 29250
rect 5079 29216 5095 29250
rect 5095 29216 5113 29250
rect 5152 29216 5163 29250
rect 5163 29216 5186 29250
rect 5225 29216 5231 29250
rect 5231 29216 5259 29250
rect 5298 29216 5299 29250
rect 5299 29216 5332 29250
rect 5371 29216 5401 29250
rect 5401 29216 5405 29250
rect 5444 29216 5469 29250
rect 5469 29216 5478 29250
rect 5517 29216 5537 29250
rect 5537 29216 5551 29250
rect 5590 29216 5605 29250
rect 5605 29216 5624 29250
rect 5663 29216 5673 29250
rect 5673 29216 5697 29250
rect 5736 29216 5741 29250
rect 5741 29216 5770 29250
rect 5809 29216 5843 29250
rect 5882 29216 5911 29250
rect 5911 29216 5916 29250
rect 5955 29216 5979 29250
rect 5979 29216 5989 29250
rect 6027 29216 6047 29250
rect 6047 29216 6061 29250
rect 6099 29216 6115 29250
rect 6115 29216 6133 29250
rect 6171 29216 6183 29250
rect 6183 29216 6205 29250
rect 6243 29216 6251 29250
rect 6251 29216 6277 29250
rect 6315 29216 6319 29250
rect 6319 29216 6349 29250
rect 6387 29216 6421 29250
rect 6459 29216 6489 29250
rect 6489 29216 6493 29250
rect 6531 29216 6557 29250
rect 6557 29216 6565 29250
rect 6603 29216 6625 29250
rect 6625 29216 6637 29250
rect 6675 29216 6693 29250
rect 6693 29216 6709 29250
rect 6747 29216 6761 29250
rect 6761 29216 6781 29250
rect 6819 29216 6829 29250
rect 6829 29216 6853 29250
rect 6891 29216 6897 29250
rect 6897 29216 6925 29250
rect 6963 29216 6965 29250
rect 6965 29216 6997 29250
rect 7035 29216 7067 29250
rect 7067 29216 7069 29250
rect 7107 29216 7135 29250
rect 7135 29216 7141 29250
rect 7179 29216 7203 29250
rect 7203 29216 7213 29250
rect 7251 29216 7271 29250
rect 7271 29216 7285 29250
rect 7323 29216 7339 29250
rect 7339 29216 7357 29250
rect 7395 29216 7407 29250
rect 7407 29216 7429 29250
rect 7467 29216 7475 29250
rect 7475 29216 7501 29250
rect 7539 29216 7543 29250
rect 7543 29216 7573 29250
rect 7611 29216 7645 29250
rect 7683 29216 7713 29250
rect 7713 29216 7717 29250
rect 8184 29243 8218 29277
rect 2276 29138 2310 29172
rect 2410 29138 2444 29172
rect 2276 29066 2310 29100
rect 2410 29066 2444 29100
rect 2276 28994 2310 29028
rect 2410 28994 2444 29028
rect 8050 29181 8084 29215
rect 8184 29171 8218 29205
rect 8050 29109 8084 29143
rect 8184 29099 8218 29133
rect 8050 29037 8084 29071
rect 8184 29027 8218 29061
rect 2276 28922 2310 28956
rect 2410 28922 2444 28956
rect 2276 28850 2310 28884
rect 2410 28850 2444 28884
rect 2276 28778 2310 28812
rect 2410 28778 2444 28812
rect 2276 28706 2310 28740
rect 2410 28706 2444 28740
rect 2276 28634 2310 28668
rect 2410 28634 2444 28668
rect 2276 28562 2310 28596
rect 2410 28562 2444 28596
rect 2276 28490 2310 28524
rect 2410 28490 2444 28524
rect 2276 28418 2310 28452
rect 2410 28418 2444 28452
rect 2276 28346 2310 28380
rect 2410 28346 2444 28380
rect 2276 28274 2310 28308
rect 2410 28274 2444 28308
rect 2276 28202 2310 28236
rect 2410 28202 2444 28236
rect 2276 28130 2310 28164
rect 2410 28130 2444 28164
rect 2276 28058 2310 28092
rect 2410 28058 2444 28092
rect 2276 27986 2310 28020
rect 2410 27986 2444 28020
rect 2276 27914 2310 27948
rect 2410 27914 2444 27948
rect 2276 27842 2310 27876
rect 2410 27842 2444 27876
rect 2276 27770 2310 27804
rect 2410 27770 2444 27804
rect 2276 27698 2310 27732
rect 2410 27698 2444 27732
rect 2276 27626 2310 27660
rect 2410 27626 2444 27660
rect 2276 27554 2310 27588
rect 2410 27554 2444 27588
rect 2276 27482 2310 27516
rect 2410 27482 2444 27516
rect 2276 27410 2310 27444
rect 2410 27410 2444 27444
rect 2276 27338 2310 27372
rect 2410 27338 2444 27372
rect 2276 27266 2310 27300
rect 2410 27266 2444 27300
rect 2276 27194 2310 27228
rect 2410 27194 2444 27228
rect 2276 27122 2310 27156
rect 2410 27122 2444 27156
rect 2276 27050 2310 27084
rect 2410 27050 2444 27084
rect 2276 26978 2310 27012
rect 2410 26978 2444 27012
rect 2276 26906 2310 26940
rect 2410 26906 2444 26940
rect 2276 26834 2310 26868
rect 2410 26834 2444 26868
rect 2276 26762 2310 26796
rect 2410 26762 2444 26796
rect 2276 26690 2310 26724
rect 2410 26690 2444 26724
rect 2276 26618 2310 26652
rect 2410 26618 2444 26652
rect 2276 26546 2310 26580
rect 2410 26546 2444 26580
rect 2276 26474 2310 26508
rect 2410 26474 2444 26508
rect 2276 26402 2310 26436
rect 2410 26402 2444 26436
rect 2276 26330 2310 26364
rect 2410 26330 2444 26364
rect 2276 26258 2310 26292
rect 2410 26258 2444 26292
rect 2276 26186 2310 26220
rect 2410 26186 2444 26220
rect 2276 26114 2310 26148
rect 2410 26114 2444 26148
rect 2276 26042 2310 26076
rect 2410 26042 2444 26076
rect 2276 25970 2310 26004
rect 2410 25970 2444 26004
rect 2276 25898 2310 25932
rect 2410 25898 2444 25932
rect 2276 25826 2310 25860
rect 2410 25826 2444 25860
rect 2276 25754 2310 25788
rect 2410 25754 2444 25788
rect 2276 25682 2310 25716
rect 2410 25682 2444 25716
rect 2276 25610 2310 25644
rect 2410 25610 2444 25644
rect 2276 25538 2310 25572
rect 2410 25538 2444 25572
rect 2276 25466 2310 25500
rect 2410 25466 2444 25500
rect 2276 25394 2310 25428
rect 2410 25394 2444 25428
rect 2276 25322 2310 25356
rect 2410 25322 2444 25356
rect 2276 25250 2310 25284
rect 2410 25250 2444 25284
rect 2276 25178 2310 25212
rect 2410 25178 2444 25212
rect 2276 25106 2310 25140
rect 2410 25106 2444 25140
rect 2276 25034 2310 25068
rect 2410 25034 2444 25068
rect 2276 24962 2310 24996
rect 2410 24962 2444 24996
rect 2276 24890 2310 24924
rect 2410 24890 2444 24924
rect 2276 24818 2310 24852
rect 2410 24818 2444 24852
rect 2276 24746 2310 24780
rect 2410 24746 2444 24780
rect 2276 24674 2310 24708
rect 2410 24674 2444 24708
rect 2276 24602 2310 24636
rect 2410 24602 2444 24636
rect 2276 24530 2310 24564
rect 2410 24530 2444 24564
rect 2276 24458 2310 24492
rect 2410 24458 2444 24492
rect 2276 24386 2310 24420
rect 2410 24386 2444 24420
rect 2276 24314 2310 24348
rect 2410 24314 2444 24348
rect 2276 24242 2310 24276
rect 2410 24242 2444 24276
rect 2276 24170 2310 24204
rect 2410 24170 2444 24204
rect 2276 24098 2310 24132
rect 2410 24098 2444 24132
rect 2276 24026 2310 24060
rect 2410 24026 2444 24060
rect 2276 23954 2310 23988
rect 2410 23954 2444 23988
rect 2276 23882 2310 23916
rect 2410 23882 2444 23916
rect 2276 23810 2310 23844
rect 2410 23810 2444 23844
rect 2276 23738 2310 23772
rect 2410 23738 2444 23772
rect 2276 23666 2310 23700
rect 2410 23666 2444 23700
rect 2276 23594 2310 23628
rect 2410 23594 2444 23628
rect 2276 23522 2310 23556
rect 2410 23522 2444 23556
rect 2276 23450 2310 23484
rect 2410 23450 2444 23484
rect 2276 23378 2310 23412
rect 2410 23378 2444 23412
rect 2276 23306 2310 23340
rect 2410 23306 2444 23340
rect 2276 23234 2310 23268
rect 2410 23234 2444 23268
rect 2276 23162 2310 23196
rect 2410 23162 2444 23196
rect 2276 23090 2310 23124
rect 2410 23090 2444 23124
rect 2276 23018 2310 23052
rect 2410 23018 2444 23052
rect 2276 22946 2310 22980
rect 2410 22946 2444 22980
rect 2276 22874 2310 22908
rect 2410 22874 2444 22908
rect 2276 22802 2310 22836
rect 2410 22802 2444 22836
rect 2276 22730 2310 22764
rect 2410 22730 2444 22764
rect 2276 22658 2310 22692
rect 2410 22658 2444 22692
rect 2276 22586 2310 22620
rect 2410 22586 2444 22620
rect 2276 22514 2310 22548
rect 2410 22514 2444 22548
rect 2276 22442 2310 22476
rect 2410 22442 2444 22476
rect 2276 22370 2310 22404
rect 2410 22370 2444 22404
rect 2276 22298 2310 22332
rect 2410 22298 2444 22332
rect 2276 22226 2310 22260
rect 2410 22226 2444 22260
rect 2276 22154 2310 22188
rect 2410 22154 2444 22188
rect 2276 22082 2310 22116
rect 2410 22082 2444 22116
rect 2276 22010 2310 22044
rect 2410 22010 2444 22044
rect 2276 21938 2310 21972
rect 2410 21938 2444 21972
rect 2276 21866 2310 21900
rect 2410 21866 2444 21900
rect 2276 21794 2310 21828
rect 2410 21794 2444 21828
rect 2276 21722 2310 21756
rect 2410 21722 2444 21756
rect 2276 21650 2310 21684
rect 2410 21650 2444 21684
rect 2276 21578 2310 21612
rect 2410 21578 2444 21612
rect 2276 21506 2310 21540
rect 2410 21506 2444 21540
rect 2276 21434 2310 21468
rect 2410 21434 2444 21468
rect 2276 21362 2310 21396
rect 2410 21362 2444 21396
rect 2276 21290 2310 21324
rect 2410 21290 2444 21324
rect 2276 21218 2310 21252
rect 2410 21218 2444 21252
rect 2276 21146 2310 21180
rect 2410 21146 2444 21180
rect 2276 21074 2310 21108
rect 2410 21074 2444 21108
rect 2276 21002 2310 21036
rect 2410 21002 2444 21036
rect 2276 20930 2310 20964
rect 2410 20930 2444 20964
rect 2276 20858 2310 20892
rect 2410 20858 2444 20892
rect 2276 20786 2310 20820
rect 2410 20786 2444 20820
rect 2276 20714 2310 20748
rect 2410 20714 2444 20748
rect 2276 20642 2310 20676
rect 2410 20642 2444 20676
rect 2276 20570 2310 20604
rect 2410 20570 2444 20604
rect 2276 20498 2310 20532
rect 2410 20498 2444 20532
rect 2276 20426 2310 20460
rect 2410 20426 2444 20460
rect 2276 20354 2310 20388
rect 2410 20354 2444 20388
rect 2276 20282 2310 20316
rect 2410 20282 2444 20316
rect 2276 20210 2310 20244
rect 2410 20210 2444 20244
rect 2276 20138 2310 20172
rect 2410 20138 2444 20172
rect 2276 20066 2310 20100
rect 2410 20066 2444 20100
rect 2276 19994 2310 20028
rect 2410 19994 2444 20028
rect 2276 19922 2310 19956
rect 2410 19922 2444 19956
rect 2276 19850 2310 19884
rect 2410 19850 2444 19884
rect 2276 19778 2310 19812
rect 2410 19778 2444 19812
rect 2276 19706 2310 19740
rect 2410 19706 2444 19740
rect 2276 19634 2310 19668
rect 2410 19634 2444 19668
rect 2276 19562 2310 19596
rect 2410 19562 2444 19596
rect 2276 19490 2310 19524
rect 2410 19490 2444 19524
rect 2276 19418 2310 19452
rect 2410 19418 2444 19452
rect 2276 19346 2310 19380
rect 2410 19346 2444 19380
rect 2276 19274 2310 19308
rect 2410 19274 2444 19308
rect 2276 19202 2310 19236
rect 2410 19202 2444 19236
rect 2276 19130 2310 19164
rect 2410 19130 2444 19164
rect 2276 19058 2310 19092
rect 2410 19058 2444 19092
rect 2276 18986 2310 19020
rect 2410 18986 2444 19020
rect 2276 18914 2310 18948
rect 2410 18914 2444 18948
rect 2276 18842 2310 18876
rect 2410 18842 2444 18876
rect 2276 18770 2310 18804
rect 2410 18770 2444 18804
rect 2276 18698 2310 18732
rect 2410 18698 2444 18732
rect 2276 18626 2310 18660
rect 2410 18626 2444 18660
rect 2276 18554 2310 18588
rect 2410 18554 2444 18588
rect 2276 18482 2310 18516
rect 2410 18482 2444 18516
rect 2276 18410 2310 18444
rect 2410 18410 2444 18444
rect 2276 18338 2310 18372
rect 2410 18338 2444 18372
rect 2276 18266 2310 18300
rect 2410 18266 2444 18300
rect 2276 18194 2310 18228
rect 2410 18194 2444 18228
rect 2276 18122 2310 18156
rect 2410 18122 2444 18156
rect 2276 18050 2310 18084
rect 2410 18050 2444 18084
rect 2276 17978 2310 18012
rect 2410 17978 2444 18012
rect 2276 17906 2310 17940
rect 2410 17906 2444 17940
rect 2276 17834 2310 17868
rect 2410 17834 2444 17868
rect 2276 17762 2310 17796
rect 2410 17762 2444 17796
rect 2276 17690 2310 17724
rect 2410 17690 2444 17724
rect 2276 17618 2310 17652
rect 2410 17618 2444 17652
rect 2276 17546 2310 17580
rect 2410 17546 2444 17580
rect 2276 17474 2310 17508
rect 2410 17474 2444 17508
rect 2276 17402 2310 17436
rect 2410 17402 2444 17436
rect 2276 17330 2310 17364
rect 2410 17330 2444 17364
rect 2276 17258 2310 17292
rect 2410 17258 2444 17292
rect 2276 17186 2310 17220
rect 2410 17186 2444 17220
rect 2276 17114 2310 17148
rect 2410 17114 2444 17148
rect 2276 17042 2310 17076
rect 2410 17042 2444 17076
rect 2276 16970 2310 17004
rect 2410 16970 2444 17004
rect 2276 16898 2310 16932
rect 2410 16898 2444 16932
rect 2276 16826 2310 16860
rect 2410 16826 2444 16860
rect 2276 16754 2310 16788
rect 2410 16754 2444 16788
rect 2276 16682 2310 16716
rect 2410 16682 2444 16716
rect 2276 16610 2310 16644
rect 2410 16610 2444 16644
rect 2276 16538 2310 16572
rect 2410 16538 2444 16572
rect 2276 16466 2310 16500
rect 2410 16466 2444 16500
rect 2276 16394 2310 16428
rect 2410 16394 2444 16428
rect 2276 16322 2310 16356
rect 2410 16322 2444 16356
rect 2276 16250 2310 16284
rect 2410 16250 2444 16284
rect 2276 16178 2310 16212
rect 2410 16178 2444 16212
rect 2276 16106 2310 16140
rect 2410 16106 2444 16140
rect 2276 16034 2310 16068
rect 2410 16034 2444 16068
rect 2276 15962 2310 15996
rect 2410 15962 2444 15996
rect 2663 28958 4569 28965
rect 2663 28924 2715 28958
rect 2715 28924 2749 28958
rect 2749 28924 2853 28958
rect 2853 28924 2887 28958
rect 2887 28924 2991 28958
rect 2991 28924 3025 28958
rect 3025 28924 3129 28958
rect 3129 28924 3163 28958
rect 3163 28924 3267 28958
rect 3267 28924 3301 28958
rect 3301 28924 3405 28958
rect 3405 28924 3439 28958
rect 3439 28924 3543 28958
rect 3543 28924 3577 28958
rect 3577 28924 3681 28958
rect 3681 28924 3715 28958
rect 3715 28924 3819 28958
rect 3819 28924 3853 28958
rect 3853 28924 3957 28958
rect 3957 28924 3991 28958
rect 3991 28924 4095 28958
rect 4095 28924 4129 28958
rect 4129 28924 4233 28958
rect 4233 28924 4267 28958
rect 4267 28924 4371 28958
rect 4371 28924 4405 28958
rect 4405 28924 4509 28958
rect 4509 28924 4543 28958
rect 4543 28924 4569 28958
rect 2663 28822 4569 28924
rect 2663 28788 2715 28822
rect 2715 28788 2749 28822
rect 2749 28788 2853 28822
rect 2853 28788 2887 28822
rect 2887 28788 2991 28822
rect 2991 28788 3025 28822
rect 3025 28788 3129 28822
rect 3129 28788 3163 28822
rect 3163 28788 3267 28822
rect 3267 28788 3301 28822
rect 3301 28788 3405 28822
rect 3405 28788 3439 28822
rect 3439 28788 3543 28822
rect 3543 28788 3577 28822
rect 3577 28788 3681 28822
rect 3681 28788 3715 28822
rect 3715 28788 3819 28822
rect 3819 28788 3853 28822
rect 3853 28788 3957 28822
rect 3957 28788 3991 28822
rect 3991 28788 4095 28822
rect 4095 28788 4129 28822
rect 4129 28788 4233 28822
rect 4233 28788 4267 28822
rect 4267 28788 4371 28822
rect 4371 28788 4405 28822
rect 4405 28788 4509 28822
rect 4509 28788 4543 28822
rect 4543 28788 4569 28822
rect 2663 28686 4569 28788
rect 8050 28965 8084 28999
rect 8184 28955 8218 28989
rect 8050 28893 8084 28927
rect 8184 28883 8218 28917
rect 8050 28821 8084 28855
rect 8184 28811 8218 28845
rect 8050 28749 8084 28783
rect 8184 28739 8218 28773
rect 2663 28652 2715 28686
rect 2715 28652 2749 28686
rect 2749 28652 2853 28686
rect 2853 28652 2887 28686
rect 2887 28652 2991 28686
rect 2991 28652 3025 28686
rect 3025 28652 3129 28686
rect 3129 28652 3163 28686
rect 3163 28652 3267 28686
rect 3267 28652 3301 28686
rect 3301 28652 3405 28686
rect 3405 28652 3439 28686
rect 3439 28652 3543 28686
rect 3543 28652 3577 28686
rect 3577 28652 3681 28686
rect 3681 28652 3715 28686
rect 3715 28652 3819 28686
rect 3819 28652 3853 28686
rect 3853 28652 3957 28686
rect 3957 28652 3991 28686
rect 3991 28652 4095 28686
rect 4095 28652 4129 28686
rect 4129 28652 4233 28686
rect 4233 28652 4267 28686
rect 4267 28652 4371 28686
rect 4371 28652 4405 28686
rect 4405 28652 4509 28686
rect 4509 28652 4543 28686
rect 4543 28652 4569 28686
rect 2663 28550 4569 28652
rect 2663 28516 2715 28550
rect 2715 28516 2749 28550
rect 2749 28516 2853 28550
rect 2853 28516 2887 28550
rect 2887 28516 2991 28550
rect 2991 28516 3025 28550
rect 3025 28516 3129 28550
rect 3129 28516 3163 28550
rect 3163 28516 3267 28550
rect 3267 28516 3301 28550
rect 3301 28516 3405 28550
rect 3405 28516 3439 28550
rect 3439 28516 3543 28550
rect 3543 28516 3577 28550
rect 3577 28516 3681 28550
rect 3681 28516 3715 28550
rect 3715 28516 3819 28550
rect 3819 28516 3853 28550
rect 3853 28516 3957 28550
rect 3957 28516 3991 28550
rect 3991 28516 4095 28550
rect 4095 28516 4129 28550
rect 4129 28516 4233 28550
rect 4233 28516 4267 28550
rect 4267 28516 4371 28550
rect 4371 28516 4405 28550
rect 4405 28516 4509 28550
rect 4509 28516 4543 28550
rect 4543 28516 4569 28550
rect 2663 28414 4569 28516
rect 2663 28380 2715 28414
rect 2715 28380 2749 28414
rect 2749 28380 2853 28414
rect 2853 28380 2887 28414
rect 2887 28380 2991 28414
rect 2991 28380 3025 28414
rect 3025 28380 3129 28414
rect 3129 28380 3163 28414
rect 3163 28380 3267 28414
rect 3267 28380 3301 28414
rect 3301 28380 3405 28414
rect 3405 28380 3439 28414
rect 3439 28380 3543 28414
rect 3543 28380 3577 28414
rect 3577 28380 3681 28414
rect 3681 28380 3715 28414
rect 3715 28380 3819 28414
rect 3819 28380 3853 28414
rect 3853 28380 3957 28414
rect 3957 28380 3991 28414
rect 3991 28380 4095 28414
rect 4095 28380 4129 28414
rect 4129 28380 4233 28414
rect 4233 28380 4267 28414
rect 4267 28380 4371 28414
rect 4371 28380 4405 28414
rect 4405 28380 4509 28414
rect 4509 28380 4543 28414
rect 4543 28380 4569 28414
rect 2663 28278 4569 28380
rect 2663 28244 2715 28278
rect 2715 28244 2749 28278
rect 2749 28244 2853 28278
rect 2853 28244 2887 28278
rect 2887 28244 2991 28278
rect 2991 28244 3025 28278
rect 3025 28244 3129 28278
rect 3129 28244 3163 28278
rect 3163 28244 3267 28278
rect 3267 28244 3301 28278
rect 3301 28244 3405 28278
rect 3405 28244 3439 28278
rect 3439 28244 3543 28278
rect 3543 28244 3577 28278
rect 3577 28244 3681 28278
rect 3681 28244 3715 28278
rect 3715 28244 3819 28278
rect 3819 28244 3853 28278
rect 3853 28244 3957 28278
rect 3957 28244 3991 28278
rect 3991 28244 4095 28278
rect 4095 28244 4129 28278
rect 4129 28244 4233 28278
rect 4233 28244 4267 28278
rect 4267 28244 4371 28278
rect 4371 28244 4405 28278
rect 4405 28244 4509 28278
rect 4509 28244 4543 28278
rect 4543 28244 4569 28278
rect 2663 28142 4569 28244
rect 2663 28108 2715 28142
rect 2715 28108 2749 28142
rect 2749 28108 2853 28142
rect 2853 28108 2887 28142
rect 2887 28108 2991 28142
rect 2991 28108 3025 28142
rect 3025 28108 3129 28142
rect 3129 28108 3163 28142
rect 3163 28108 3267 28142
rect 3267 28108 3301 28142
rect 3301 28108 3405 28142
rect 3405 28108 3439 28142
rect 3439 28108 3543 28142
rect 3543 28108 3577 28142
rect 3577 28108 3681 28142
rect 3681 28108 3715 28142
rect 3715 28108 3819 28142
rect 3819 28108 3853 28142
rect 3853 28108 3957 28142
rect 3957 28108 3991 28142
rect 3991 28108 4095 28142
rect 4095 28108 4129 28142
rect 4129 28108 4233 28142
rect 4233 28108 4267 28142
rect 4267 28108 4371 28142
rect 4371 28108 4405 28142
rect 4405 28108 4509 28142
rect 4509 28108 4543 28142
rect 4543 28108 4569 28142
rect 2663 28006 4569 28108
rect 2663 27972 2715 28006
rect 2715 27972 2749 28006
rect 2749 27972 2853 28006
rect 2853 27972 2887 28006
rect 2887 27972 2991 28006
rect 2991 27972 3025 28006
rect 3025 27972 3129 28006
rect 3129 27972 3163 28006
rect 3163 27972 3267 28006
rect 3267 27972 3301 28006
rect 3301 27972 3405 28006
rect 3405 27972 3439 28006
rect 3439 27972 3543 28006
rect 3543 27972 3577 28006
rect 3577 27972 3681 28006
rect 3681 27972 3715 28006
rect 3715 27972 3819 28006
rect 3819 27972 3853 28006
rect 3853 27972 3957 28006
rect 3957 27972 3991 28006
rect 3991 27972 4095 28006
rect 4095 27972 4129 28006
rect 4129 27972 4233 28006
rect 4233 27972 4267 28006
rect 4267 27972 4371 28006
rect 4371 27972 4405 28006
rect 4405 27972 4509 28006
rect 4509 27972 4543 28006
rect 4543 27972 4569 28006
rect 2663 27870 4569 27972
rect 2663 27836 2715 27870
rect 2715 27836 2749 27870
rect 2749 27836 2853 27870
rect 2853 27836 2887 27870
rect 2887 27836 2991 27870
rect 2991 27836 3025 27870
rect 3025 27836 3129 27870
rect 3129 27836 3163 27870
rect 3163 27836 3267 27870
rect 3267 27836 3301 27870
rect 3301 27836 3405 27870
rect 3405 27836 3439 27870
rect 3439 27836 3543 27870
rect 3543 27836 3577 27870
rect 3577 27836 3681 27870
rect 3681 27836 3715 27870
rect 3715 27836 3819 27870
rect 3819 27836 3853 27870
rect 3853 27836 3957 27870
rect 3957 27836 3991 27870
rect 3991 27836 4095 27870
rect 4095 27836 4129 27870
rect 4129 27836 4233 27870
rect 4233 27836 4267 27870
rect 4267 27836 4371 27870
rect 4371 27836 4405 27870
rect 4405 27836 4509 27870
rect 4509 27836 4543 27870
rect 4543 27836 4569 27870
rect 2663 27734 4569 27836
rect 2663 27700 2715 27734
rect 2715 27700 2749 27734
rect 2749 27700 2853 27734
rect 2853 27700 2887 27734
rect 2887 27700 2991 27734
rect 2991 27700 3025 27734
rect 3025 27700 3129 27734
rect 3129 27700 3163 27734
rect 3163 27700 3267 27734
rect 3267 27700 3301 27734
rect 3301 27700 3405 27734
rect 3405 27700 3439 27734
rect 3439 27700 3543 27734
rect 3543 27700 3577 27734
rect 3577 27700 3681 27734
rect 3681 27700 3715 27734
rect 3715 27700 3819 27734
rect 3819 27700 3853 27734
rect 3853 27700 3957 27734
rect 3957 27700 3991 27734
rect 3991 27700 4095 27734
rect 4095 27700 4129 27734
rect 4129 27700 4233 27734
rect 4233 27700 4267 27734
rect 4267 27700 4371 27734
rect 4371 27700 4405 27734
rect 4405 27700 4509 27734
rect 4509 27700 4543 27734
rect 4543 27700 4569 27734
rect 2663 27598 4569 27700
rect 2663 27564 2715 27598
rect 2715 27564 2749 27598
rect 2749 27564 2853 27598
rect 2853 27564 2887 27598
rect 2887 27564 2991 27598
rect 2991 27564 3025 27598
rect 3025 27564 3129 27598
rect 3129 27564 3163 27598
rect 3163 27564 3267 27598
rect 3267 27564 3301 27598
rect 3301 27564 3405 27598
rect 3405 27564 3439 27598
rect 3439 27564 3543 27598
rect 3543 27564 3577 27598
rect 3577 27564 3681 27598
rect 3681 27564 3715 27598
rect 3715 27564 3819 27598
rect 3819 27564 3853 27598
rect 3853 27564 3957 27598
rect 3957 27564 3991 27598
rect 3991 27564 4095 27598
rect 4095 27564 4129 27598
rect 4129 27564 4233 27598
rect 4233 27564 4267 27598
rect 4267 27564 4371 27598
rect 4371 27564 4405 27598
rect 4405 27564 4509 27598
rect 4509 27564 4543 27598
rect 4543 27564 4569 27598
rect 2663 27462 4569 27564
rect 2663 27428 2715 27462
rect 2715 27428 2749 27462
rect 2749 27428 2853 27462
rect 2853 27428 2887 27462
rect 2887 27428 2991 27462
rect 2991 27428 3025 27462
rect 3025 27428 3129 27462
rect 3129 27428 3163 27462
rect 3163 27428 3267 27462
rect 3267 27428 3301 27462
rect 3301 27428 3405 27462
rect 3405 27428 3439 27462
rect 3439 27428 3543 27462
rect 3543 27428 3577 27462
rect 3577 27428 3681 27462
rect 3681 27428 3715 27462
rect 3715 27428 3819 27462
rect 3819 27428 3853 27462
rect 3853 27428 3957 27462
rect 3957 27428 3991 27462
rect 3991 27428 4095 27462
rect 4095 27428 4129 27462
rect 4129 27428 4233 27462
rect 4233 27428 4267 27462
rect 4267 27428 4371 27462
rect 4371 27428 4405 27462
rect 4405 27428 4509 27462
rect 4509 27428 4543 27462
rect 4543 27428 4569 27462
rect 2663 27326 4569 27428
rect 5046 28680 5080 28714
rect 5118 28680 5152 28714
rect 5046 28607 5080 28641
rect 5118 28607 5152 28641
rect 5046 28534 5080 28568
rect 5118 28534 5152 28568
rect 5046 28461 5080 28495
rect 5118 28461 5152 28495
rect 5046 27380 5152 28422
rect 5323 28680 5357 28714
rect 5395 28680 5429 28714
rect 5323 28607 5357 28641
rect 5395 28607 5429 28641
rect 5323 28534 5357 28568
rect 5395 28534 5429 28568
rect 5323 28461 5357 28495
rect 5395 28461 5429 28495
rect 5323 27380 5429 28422
rect 5600 28680 5634 28714
rect 5672 28680 5706 28714
rect 5600 28607 5634 28641
rect 5672 28607 5706 28641
rect 5600 28534 5634 28568
rect 5672 28534 5706 28568
rect 5600 28461 5634 28495
rect 5672 28461 5706 28495
rect 5600 27380 5706 28422
rect 5877 28680 5911 28714
rect 5949 28680 5983 28714
rect 5877 28607 5911 28641
rect 5949 28607 5983 28641
rect 5877 28534 5911 28568
rect 5949 28534 5983 28568
rect 5877 28461 5911 28495
rect 5949 28461 5983 28495
rect 5877 27380 5983 28422
rect 6154 28680 6188 28714
rect 6226 28680 6260 28714
rect 6154 28607 6188 28641
rect 6226 28607 6260 28641
rect 6154 28534 6188 28568
rect 6226 28534 6260 28568
rect 6154 28461 6188 28495
rect 6226 28461 6260 28495
rect 6154 27380 6260 28422
rect 6431 28680 6465 28714
rect 6503 28680 6537 28714
rect 6431 28607 6465 28641
rect 6503 28607 6537 28641
rect 6431 28534 6465 28568
rect 6503 28534 6537 28568
rect 6431 28461 6465 28495
rect 6503 28461 6537 28495
rect 6431 27380 6537 28422
rect 6708 28680 6742 28714
rect 6780 28680 6814 28714
rect 6708 28607 6742 28641
rect 6780 28607 6814 28641
rect 6708 28534 6742 28568
rect 6780 28534 6814 28568
rect 6708 28461 6742 28495
rect 6780 28461 6814 28495
rect 6708 27380 6814 28422
rect 6985 28680 7019 28714
rect 7057 28680 7091 28714
rect 6985 28607 7019 28641
rect 7057 28607 7091 28641
rect 6985 28534 7019 28568
rect 7057 28534 7091 28568
rect 6985 28461 7019 28495
rect 7057 28461 7091 28495
rect 6985 27380 7091 28422
rect 7262 28680 7296 28714
rect 7334 28680 7368 28714
rect 7262 28607 7296 28641
rect 7334 28607 7368 28641
rect 7262 28534 7296 28568
rect 7334 28534 7368 28568
rect 7262 28461 7296 28495
rect 7334 28461 7368 28495
rect 7262 27380 7368 28422
rect 7539 28680 7573 28714
rect 7611 28680 7645 28714
rect 7539 28607 7573 28641
rect 7611 28607 7645 28641
rect 7539 28534 7573 28568
rect 7611 28534 7645 28568
rect 7539 28461 7573 28495
rect 7611 28461 7645 28495
rect 7539 27380 7645 28422
rect 7816 28680 7850 28714
rect 7888 28680 7922 28714
rect 7816 28607 7850 28641
rect 7888 28607 7922 28641
rect 7816 28534 7850 28568
rect 7888 28534 7922 28568
rect 7816 28461 7850 28495
rect 7888 28461 7922 28495
rect 7816 27380 7922 28422
rect 8050 28677 8084 28711
rect 8184 28667 8218 28701
rect 8050 28605 8084 28639
rect 8184 28595 8218 28629
rect 8050 28533 8084 28567
rect 8184 28523 8218 28557
rect 8050 28461 8084 28495
rect 8184 28451 8218 28485
rect 8050 28389 8084 28423
rect 8184 28379 8218 28413
rect 8050 28317 8084 28351
rect 8184 28307 8218 28341
rect 8050 28245 8084 28279
rect 8184 28235 8218 28269
rect 8050 28173 8084 28207
rect 8184 28163 8218 28197
rect 8050 28101 8084 28135
rect 8184 28091 8218 28125
rect 8050 28029 8084 28063
rect 8184 28019 8218 28053
rect 8050 27957 8084 27991
rect 8184 27947 8218 27981
rect 8050 27885 8084 27919
rect 8184 27875 8218 27909
rect 8050 27813 8084 27847
rect 8184 27803 8218 27837
rect 8050 27741 8084 27775
rect 8184 27731 8218 27765
rect 8050 27669 8084 27703
rect 8184 27659 8218 27693
rect 8050 27597 8084 27631
rect 8184 27587 8218 27621
rect 8050 27525 8084 27559
rect 8184 27515 8218 27549
rect 8050 27453 8084 27487
rect 8184 27443 8218 27477
rect 8050 27381 8084 27415
rect 8184 27371 8218 27405
rect 2663 27292 2715 27326
rect 2715 27292 2749 27326
rect 2749 27292 2853 27326
rect 2853 27292 2887 27326
rect 2887 27292 2991 27326
rect 2991 27292 3025 27326
rect 3025 27292 3129 27326
rect 3129 27292 3163 27326
rect 3163 27292 3267 27326
rect 3267 27292 3301 27326
rect 3301 27292 3405 27326
rect 3405 27292 3439 27326
rect 3439 27292 3543 27326
rect 3543 27292 3577 27326
rect 3577 27292 3681 27326
rect 3681 27292 3715 27326
rect 3715 27292 3819 27326
rect 3819 27292 3853 27326
rect 3853 27292 3957 27326
rect 3957 27292 3991 27326
rect 3991 27292 4095 27326
rect 4095 27292 4129 27326
rect 4129 27292 4233 27326
rect 4233 27292 4267 27326
rect 4267 27292 4371 27326
rect 4371 27292 4405 27326
rect 4405 27292 4509 27326
rect 4509 27292 4543 27326
rect 4543 27292 4569 27326
rect 2663 27190 4569 27292
rect 2663 27156 2715 27190
rect 2715 27156 2749 27190
rect 2749 27156 2853 27190
rect 2853 27156 2887 27190
rect 2887 27156 2991 27190
rect 2991 27156 3025 27190
rect 3025 27156 3129 27190
rect 3129 27156 3163 27190
rect 3163 27156 3267 27190
rect 3267 27156 3301 27190
rect 3301 27156 3405 27190
rect 3405 27156 3439 27190
rect 3439 27156 3543 27190
rect 3543 27156 3577 27190
rect 3577 27156 3681 27190
rect 3681 27156 3715 27190
rect 3715 27156 3819 27190
rect 3819 27156 3853 27190
rect 3853 27156 3957 27190
rect 3957 27156 3991 27190
rect 3991 27156 4095 27190
rect 4095 27156 4129 27190
rect 4129 27156 4233 27190
rect 4233 27156 4267 27190
rect 4267 27156 4371 27190
rect 4371 27156 4405 27190
rect 4405 27156 4509 27190
rect 4509 27156 4543 27190
rect 4543 27156 4569 27190
rect 2663 27054 4569 27156
rect 8050 27309 8084 27343
rect 8184 27299 8218 27333
rect 8050 27237 8084 27271
rect 8184 27227 8218 27261
rect 8050 27165 8084 27199
rect 8184 27155 8218 27189
rect 5251 27071 5255 27105
rect 5255 27071 5285 27105
rect 5326 27071 5359 27105
rect 5359 27071 5360 27105
rect 5401 27071 5429 27105
rect 5429 27071 5435 27105
rect 5476 27071 5499 27105
rect 5499 27071 5510 27105
rect 5551 27071 5569 27105
rect 5569 27071 5585 27105
rect 5626 27071 5639 27105
rect 5639 27071 5660 27105
rect 5701 27071 5709 27105
rect 5709 27071 5735 27105
rect 5776 27071 5779 27105
rect 5779 27071 5810 27105
rect 5851 27071 5885 27105
rect 5926 27071 5954 27105
rect 5954 27071 5960 27105
rect 6001 27071 6023 27105
rect 6023 27071 6035 27105
rect 6076 27071 6092 27105
rect 6092 27071 6110 27105
rect 6151 27071 6161 27105
rect 6161 27071 6185 27105
rect 6225 27071 6230 27105
rect 6230 27071 6259 27105
rect 6299 27071 6333 27105
rect 6373 27071 6402 27105
rect 6402 27071 6407 27105
rect 6447 27071 6471 27105
rect 6471 27071 6481 27105
rect 6521 27071 6540 27105
rect 6540 27071 6555 27105
rect 6595 27071 6609 27105
rect 6609 27071 6629 27105
rect 6669 27071 6678 27105
rect 6678 27071 6703 27105
rect 6743 27071 6747 27105
rect 6747 27071 6777 27105
rect 6817 27071 6851 27105
rect 6891 27071 6920 27105
rect 6920 27071 6925 27105
rect 8050 27093 8084 27127
rect 8184 27083 8218 27117
rect 2663 27020 2715 27054
rect 2715 27020 2749 27054
rect 2749 27020 2853 27054
rect 2853 27020 2887 27054
rect 2887 27020 2991 27054
rect 2991 27020 3025 27054
rect 3025 27020 3129 27054
rect 3129 27020 3163 27054
rect 3163 27020 3267 27054
rect 3267 27020 3301 27054
rect 3301 27020 3405 27054
rect 3405 27020 3439 27054
rect 3439 27020 3543 27054
rect 3543 27020 3577 27054
rect 3577 27020 3681 27054
rect 3681 27020 3715 27054
rect 3715 27020 3819 27054
rect 3819 27020 3853 27054
rect 3853 27020 3957 27054
rect 3957 27020 3991 27054
rect 3991 27020 4095 27054
rect 4095 27020 4129 27054
rect 4129 27020 4233 27054
rect 4233 27020 4267 27054
rect 4267 27020 4371 27054
rect 4371 27020 4405 27054
rect 4405 27020 4509 27054
rect 4509 27020 4543 27054
rect 4543 27020 4569 27054
rect 2663 26918 4569 27020
rect 2663 26884 2715 26918
rect 2715 26884 2749 26918
rect 2749 26884 2853 26918
rect 2853 26884 2887 26918
rect 2887 26884 2991 26918
rect 2991 26884 3025 26918
rect 3025 26884 3129 26918
rect 3129 26884 3163 26918
rect 3163 26884 3267 26918
rect 3267 26884 3301 26918
rect 3301 26884 3405 26918
rect 3405 26884 3439 26918
rect 3439 26884 3543 26918
rect 3543 26884 3577 26918
rect 3577 26884 3681 26918
rect 3681 26884 3715 26918
rect 3715 26884 3819 26918
rect 3819 26884 3853 26918
rect 3853 26884 3957 26918
rect 3957 26884 3991 26918
rect 3991 26884 4095 26918
rect 4095 26884 4129 26918
rect 4129 26884 4233 26918
rect 4233 26884 4267 26918
rect 4267 26884 4371 26918
rect 4371 26884 4405 26918
rect 4405 26884 4509 26918
rect 4509 26884 4543 26918
rect 4543 26884 4569 26918
rect 2663 26782 4569 26884
rect 2663 26748 2715 26782
rect 2715 26748 2749 26782
rect 2749 26748 2853 26782
rect 2853 26748 2887 26782
rect 2887 26748 2991 26782
rect 2991 26748 3025 26782
rect 3025 26748 3129 26782
rect 3129 26748 3163 26782
rect 3163 26748 3267 26782
rect 3267 26748 3301 26782
rect 3301 26748 3405 26782
rect 3405 26748 3439 26782
rect 3439 26748 3543 26782
rect 3543 26748 3577 26782
rect 3577 26748 3681 26782
rect 3681 26748 3715 26782
rect 3715 26748 3819 26782
rect 3819 26748 3853 26782
rect 3853 26748 3957 26782
rect 3957 26748 3991 26782
rect 3991 26748 4095 26782
rect 4095 26748 4129 26782
rect 4129 26748 4233 26782
rect 4233 26748 4267 26782
rect 4267 26748 4371 26782
rect 4371 26748 4405 26782
rect 4405 26748 4509 26782
rect 4509 26748 4543 26782
rect 4543 26748 4569 26782
rect 2663 26646 4569 26748
rect 8050 27021 8084 27055
rect 8184 27011 8218 27045
rect 8050 26949 8084 26983
rect 8184 26939 8218 26973
rect 8050 26877 8084 26911
rect 8184 26867 8218 26901
rect 8050 26805 8084 26839
rect 8184 26795 8218 26829
rect 8050 26733 8084 26767
rect 8184 26723 8218 26757
rect 2663 26612 2715 26646
rect 2715 26612 2749 26646
rect 2749 26612 2853 26646
rect 2853 26612 2887 26646
rect 2887 26612 2991 26646
rect 2991 26612 3025 26646
rect 3025 26612 3129 26646
rect 3129 26612 3163 26646
rect 3163 26612 3267 26646
rect 3267 26612 3301 26646
rect 3301 26612 3405 26646
rect 3405 26612 3439 26646
rect 3439 26612 3543 26646
rect 3543 26612 3577 26646
rect 3577 26612 3681 26646
rect 3681 26612 3715 26646
rect 3715 26612 3819 26646
rect 3819 26612 3853 26646
rect 3853 26612 3957 26646
rect 3957 26612 3991 26646
rect 3991 26612 4095 26646
rect 4095 26612 4129 26646
rect 4129 26612 4233 26646
rect 4233 26612 4267 26646
rect 4267 26612 4371 26646
rect 4371 26612 4405 26646
rect 4405 26612 4509 26646
rect 4509 26612 4543 26646
rect 4543 26612 4569 26646
rect 2663 26510 4569 26612
rect 2663 26476 2715 26510
rect 2715 26476 2749 26510
rect 2749 26476 2853 26510
rect 2853 26476 2887 26510
rect 2887 26476 2991 26510
rect 2991 26476 3025 26510
rect 3025 26476 3129 26510
rect 3129 26476 3163 26510
rect 3163 26476 3267 26510
rect 3267 26476 3301 26510
rect 3301 26476 3405 26510
rect 3405 26476 3439 26510
rect 3439 26476 3543 26510
rect 3543 26476 3577 26510
rect 3577 26476 3681 26510
rect 3681 26476 3715 26510
rect 3715 26476 3819 26510
rect 3819 26476 3853 26510
rect 3853 26476 3957 26510
rect 3957 26476 3991 26510
rect 3991 26476 4095 26510
rect 4095 26476 4129 26510
rect 4129 26476 4233 26510
rect 4233 26476 4267 26510
rect 4267 26476 4371 26510
rect 4371 26476 4405 26510
rect 4405 26476 4509 26510
rect 4509 26476 4543 26510
rect 4543 26476 4569 26510
rect 2663 26374 4569 26476
rect 2663 26340 2715 26374
rect 2715 26340 2749 26374
rect 2749 26340 2853 26374
rect 2853 26340 2887 26374
rect 2887 26340 2991 26374
rect 2991 26340 3025 26374
rect 3025 26340 3129 26374
rect 3129 26340 3163 26374
rect 3163 26340 3267 26374
rect 3267 26340 3301 26374
rect 3301 26340 3405 26374
rect 3405 26340 3439 26374
rect 3439 26340 3543 26374
rect 3543 26340 3577 26374
rect 3577 26340 3681 26374
rect 3681 26340 3715 26374
rect 3715 26340 3819 26374
rect 3819 26340 3853 26374
rect 3853 26340 3957 26374
rect 3957 26340 3991 26374
rect 3991 26340 4095 26374
rect 4095 26340 4129 26374
rect 4129 26340 4233 26374
rect 4233 26340 4267 26374
rect 4267 26340 4371 26374
rect 4371 26340 4405 26374
rect 4405 26340 4509 26374
rect 4509 26340 4543 26374
rect 4543 26340 4569 26374
rect 2663 26238 4569 26340
rect 2663 26204 2715 26238
rect 2715 26204 2749 26238
rect 2749 26204 2853 26238
rect 2853 26204 2887 26238
rect 2887 26204 2991 26238
rect 2991 26204 3025 26238
rect 3025 26204 3129 26238
rect 3129 26204 3163 26238
rect 3163 26204 3267 26238
rect 3267 26204 3301 26238
rect 3301 26204 3405 26238
rect 3405 26204 3439 26238
rect 3439 26204 3543 26238
rect 3543 26204 3577 26238
rect 3577 26204 3681 26238
rect 3681 26204 3715 26238
rect 3715 26204 3819 26238
rect 3819 26204 3853 26238
rect 3853 26204 3957 26238
rect 3957 26204 3991 26238
rect 3991 26204 4095 26238
rect 4095 26204 4129 26238
rect 4129 26204 4233 26238
rect 4233 26204 4267 26238
rect 4267 26204 4371 26238
rect 4371 26204 4405 26238
rect 4405 26204 4509 26238
rect 4509 26204 4543 26238
rect 4543 26204 4569 26238
rect 2663 26102 4569 26204
rect 2663 26068 2715 26102
rect 2715 26068 2749 26102
rect 2749 26068 2853 26102
rect 2853 26068 2887 26102
rect 2887 26068 2991 26102
rect 2991 26068 3025 26102
rect 3025 26068 3129 26102
rect 3129 26068 3163 26102
rect 3163 26068 3267 26102
rect 3267 26068 3301 26102
rect 3301 26068 3405 26102
rect 3405 26068 3439 26102
rect 3439 26068 3543 26102
rect 3543 26068 3577 26102
rect 3577 26068 3681 26102
rect 3681 26068 3715 26102
rect 3715 26068 3819 26102
rect 3819 26068 3853 26102
rect 3853 26068 3957 26102
rect 3957 26068 3991 26102
rect 3991 26068 4095 26102
rect 4095 26068 4129 26102
rect 4129 26068 4233 26102
rect 4233 26068 4267 26102
rect 4267 26068 4371 26102
rect 4371 26068 4405 26102
rect 4405 26068 4509 26102
rect 4509 26068 4543 26102
rect 4543 26068 4569 26102
rect 2663 25966 4569 26068
rect 2663 25932 2715 25966
rect 2715 25932 2749 25966
rect 2749 25932 2853 25966
rect 2853 25932 2887 25966
rect 2887 25932 2991 25966
rect 2991 25932 3025 25966
rect 3025 25932 3129 25966
rect 3129 25932 3163 25966
rect 3163 25932 3267 25966
rect 3267 25932 3301 25966
rect 3301 25932 3405 25966
rect 3405 25932 3439 25966
rect 3439 25932 3543 25966
rect 3543 25932 3577 25966
rect 3577 25932 3681 25966
rect 3681 25932 3715 25966
rect 3715 25932 3819 25966
rect 3819 25932 3853 25966
rect 3853 25932 3957 25966
rect 3957 25932 3991 25966
rect 3991 25932 4095 25966
rect 4095 25932 4129 25966
rect 4129 25932 4233 25966
rect 4233 25932 4267 25966
rect 4267 25932 4371 25966
rect 4371 25932 4405 25966
rect 4405 25932 4509 25966
rect 4509 25932 4543 25966
rect 4543 25932 4569 25966
rect 2663 25830 4569 25932
rect 2663 25796 2715 25830
rect 2715 25796 2749 25830
rect 2749 25796 2853 25830
rect 2853 25796 2887 25830
rect 2887 25796 2991 25830
rect 2991 25796 3025 25830
rect 3025 25796 3129 25830
rect 3129 25796 3163 25830
rect 3163 25796 3267 25830
rect 3267 25796 3301 25830
rect 3301 25796 3405 25830
rect 3405 25796 3439 25830
rect 3439 25796 3543 25830
rect 3543 25796 3577 25830
rect 3577 25796 3681 25830
rect 3681 25796 3715 25830
rect 3715 25796 3819 25830
rect 3819 25796 3853 25830
rect 3853 25796 3957 25830
rect 3957 25796 3991 25830
rect 3991 25796 4095 25830
rect 4095 25796 4129 25830
rect 4129 25796 4233 25830
rect 4233 25796 4267 25830
rect 4267 25796 4371 25830
rect 4371 25796 4405 25830
rect 4405 25796 4509 25830
rect 4509 25796 4543 25830
rect 4543 25796 4569 25830
rect 2663 25694 4569 25796
rect 2663 25660 2715 25694
rect 2715 25660 2749 25694
rect 2749 25660 2853 25694
rect 2853 25660 2887 25694
rect 2887 25660 2991 25694
rect 2991 25660 3025 25694
rect 3025 25660 3129 25694
rect 3129 25660 3163 25694
rect 3163 25660 3267 25694
rect 3267 25660 3301 25694
rect 3301 25660 3405 25694
rect 3405 25660 3439 25694
rect 3439 25660 3543 25694
rect 3543 25660 3577 25694
rect 3577 25660 3681 25694
rect 3681 25660 3715 25694
rect 3715 25660 3819 25694
rect 3819 25660 3853 25694
rect 3853 25660 3957 25694
rect 3957 25660 3991 25694
rect 3991 25660 4095 25694
rect 4095 25660 4129 25694
rect 4129 25660 4233 25694
rect 4233 25660 4267 25694
rect 4267 25660 4371 25694
rect 4371 25660 4405 25694
rect 4405 25660 4509 25694
rect 4509 25660 4543 25694
rect 4543 25660 4569 25694
rect 2663 25558 4569 25660
rect 2663 25524 2715 25558
rect 2715 25524 2749 25558
rect 2749 25524 2853 25558
rect 2853 25524 2887 25558
rect 2887 25524 2991 25558
rect 2991 25524 3025 25558
rect 3025 25524 3129 25558
rect 3129 25524 3163 25558
rect 3163 25524 3267 25558
rect 3267 25524 3301 25558
rect 3301 25524 3405 25558
rect 3405 25524 3439 25558
rect 3439 25524 3543 25558
rect 3543 25524 3577 25558
rect 3577 25524 3681 25558
rect 3681 25524 3715 25558
rect 3715 25524 3819 25558
rect 3819 25524 3853 25558
rect 3853 25524 3957 25558
rect 3957 25524 3991 25558
rect 3991 25524 4095 25558
rect 4095 25524 4129 25558
rect 4129 25524 4233 25558
rect 4233 25524 4267 25558
rect 4267 25524 4371 25558
rect 4371 25524 4405 25558
rect 4405 25524 4509 25558
rect 4509 25524 4543 25558
rect 4543 25524 4569 25558
rect 2663 25422 4569 25524
rect 2663 25388 2715 25422
rect 2715 25388 2749 25422
rect 2749 25388 2853 25422
rect 2853 25388 2887 25422
rect 2887 25388 2991 25422
rect 2991 25388 3025 25422
rect 3025 25388 3129 25422
rect 3129 25388 3163 25422
rect 3163 25388 3267 25422
rect 3267 25388 3301 25422
rect 3301 25388 3405 25422
rect 3405 25388 3439 25422
rect 3439 25388 3543 25422
rect 3543 25388 3577 25422
rect 3577 25388 3681 25422
rect 3681 25388 3715 25422
rect 3715 25388 3819 25422
rect 3819 25388 3853 25422
rect 3853 25388 3957 25422
rect 3957 25388 3991 25422
rect 3991 25388 4095 25422
rect 4095 25388 4129 25422
rect 4129 25388 4233 25422
rect 4233 25388 4267 25422
rect 4267 25388 4371 25422
rect 4371 25388 4405 25422
rect 4405 25388 4509 25422
rect 4509 25388 4543 25422
rect 4543 25388 4569 25422
rect 2663 25286 4569 25388
rect 5046 26680 5080 26714
rect 5118 26680 5152 26714
rect 5046 26607 5080 26641
rect 5118 26607 5152 26641
rect 5046 26534 5080 26568
rect 5118 26534 5152 26568
rect 5046 26461 5080 26495
rect 5118 26461 5152 26495
rect 5046 25380 5152 26422
rect 5323 26680 5357 26714
rect 5395 26680 5429 26714
rect 5323 26607 5357 26641
rect 5395 26607 5429 26641
rect 5323 26534 5357 26568
rect 5395 26534 5429 26568
rect 5323 26461 5357 26495
rect 5395 26461 5429 26495
rect 5323 25380 5429 26422
rect 5600 26680 5634 26714
rect 5672 26680 5706 26714
rect 5600 26607 5634 26641
rect 5672 26607 5706 26641
rect 5600 26534 5634 26568
rect 5672 26534 5706 26568
rect 5600 26461 5634 26495
rect 5672 26461 5706 26495
rect 5600 25380 5706 26422
rect 5877 26680 5911 26714
rect 5949 26680 5983 26714
rect 5877 26607 5911 26641
rect 5949 26607 5983 26641
rect 5877 26534 5911 26568
rect 5949 26534 5983 26568
rect 5877 26461 5911 26495
rect 5949 26461 5983 26495
rect 5877 25380 5983 26422
rect 6154 26680 6188 26714
rect 6226 26680 6260 26714
rect 6154 26607 6188 26641
rect 6226 26607 6260 26641
rect 6154 26534 6188 26568
rect 6226 26534 6260 26568
rect 6154 26461 6188 26495
rect 6226 26461 6260 26495
rect 6154 25380 6260 26422
rect 6431 26680 6465 26714
rect 6503 26680 6537 26714
rect 6431 26607 6465 26641
rect 6503 26607 6537 26641
rect 6431 26534 6465 26568
rect 6503 26534 6537 26568
rect 6431 26461 6465 26495
rect 6503 26461 6537 26495
rect 6431 25380 6537 26422
rect 6708 26680 6742 26714
rect 6780 26680 6814 26714
rect 6708 26607 6742 26641
rect 6780 26607 6814 26641
rect 6708 26534 6742 26568
rect 6780 26534 6814 26568
rect 6708 26461 6742 26495
rect 6780 26461 6814 26495
rect 6708 25380 6814 26422
rect 6985 26680 7019 26714
rect 7057 26680 7091 26714
rect 6985 26607 7019 26641
rect 7057 26607 7091 26641
rect 6985 26534 7019 26568
rect 7057 26534 7091 26568
rect 6985 26461 7019 26495
rect 7057 26461 7091 26495
rect 6985 25380 7091 26422
rect 7262 26680 7296 26714
rect 7334 26680 7368 26714
rect 7262 26607 7296 26641
rect 7334 26607 7368 26641
rect 7262 26534 7296 26568
rect 7334 26534 7368 26568
rect 7262 26461 7296 26495
rect 7334 26461 7368 26495
rect 7262 25380 7368 26422
rect 7539 26680 7573 26714
rect 7611 26680 7645 26714
rect 7539 26607 7573 26641
rect 7611 26607 7645 26641
rect 7539 26534 7573 26568
rect 7611 26534 7645 26568
rect 7539 26461 7573 26495
rect 7611 26461 7645 26495
rect 7539 25380 7645 26422
rect 7816 26680 7850 26714
rect 7888 26680 7922 26714
rect 7816 26607 7850 26641
rect 7888 26607 7922 26641
rect 7816 26534 7850 26568
rect 7888 26534 7922 26568
rect 7816 26461 7850 26495
rect 7888 26461 7922 26495
rect 7816 25380 7922 26422
rect 8050 26661 8084 26695
rect 8184 26651 8218 26685
rect 8050 26589 8084 26623
rect 8184 26579 8218 26613
rect 8050 26517 8084 26551
rect 8184 26507 8218 26541
rect 8050 26445 8084 26479
rect 8184 26435 8218 26469
rect 8050 26373 8084 26407
rect 8184 26363 8218 26397
rect 8050 26301 8084 26335
rect 8184 26291 8218 26325
rect 8050 26229 8084 26263
rect 8184 26219 8218 26253
rect 8050 26157 8084 26191
rect 8184 26147 8218 26181
rect 8050 26085 8084 26119
rect 8184 26075 8218 26109
rect 8050 26013 8084 26047
rect 8184 26003 8218 26037
rect 8050 25941 8084 25975
rect 8184 25931 8218 25965
rect 8050 25869 8084 25903
rect 8184 25859 8218 25893
rect 8050 25797 8084 25831
rect 8184 25787 8218 25821
rect 8050 25725 8084 25759
rect 8184 25715 8218 25749
rect 8050 25653 8084 25687
rect 8184 25643 8218 25677
rect 8050 25581 8084 25615
rect 8184 25571 8218 25605
rect 8050 25509 8084 25543
rect 8184 25499 8218 25533
rect 8050 25437 8084 25471
rect 8184 25427 8218 25461
rect 2663 25252 2715 25286
rect 2715 25252 2749 25286
rect 2749 25252 2853 25286
rect 2853 25252 2887 25286
rect 2887 25252 2991 25286
rect 2991 25252 3025 25286
rect 3025 25252 3129 25286
rect 3129 25252 3163 25286
rect 3163 25252 3267 25286
rect 3267 25252 3301 25286
rect 3301 25252 3405 25286
rect 3405 25252 3439 25286
rect 3439 25252 3543 25286
rect 3543 25252 3577 25286
rect 3577 25252 3681 25286
rect 3681 25252 3715 25286
rect 3715 25252 3819 25286
rect 3819 25252 3853 25286
rect 3853 25252 3957 25286
rect 3957 25252 3991 25286
rect 3991 25252 4095 25286
rect 4095 25252 4129 25286
rect 4129 25252 4233 25286
rect 4233 25252 4267 25286
rect 4267 25252 4371 25286
rect 4371 25252 4405 25286
rect 4405 25252 4509 25286
rect 4509 25252 4543 25286
rect 4543 25252 4569 25286
rect 2663 25149 4569 25252
rect 2663 25115 2715 25149
rect 2715 25115 2749 25149
rect 2749 25115 2853 25149
rect 2853 25115 2887 25149
rect 2887 25115 2991 25149
rect 2991 25115 3025 25149
rect 3025 25115 3129 25149
rect 3129 25115 3163 25149
rect 3163 25115 3267 25149
rect 3267 25115 3301 25149
rect 3301 25115 3405 25149
rect 3405 25115 3439 25149
rect 3439 25115 3543 25149
rect 3543 25115 3577 25149
rect 3577 25115 3681 25149
rect 3681 25115 3715 25149
rect 3715 25115 3819 25149
rect 3819 25115 3853 25149
rect 3853 25115 3957 25149
rect 3957 25115 3991 25149
rect 3991 25115 4095 25149
rect 4095 25115 4129 25149
rect 4129 25115 4233 25149
rect 4233 25115 4267 25149
rect 4267 25115 4371 25149
rect 4371 25115 4405 25149
rect 4405 25115 4509 25149
rect 4509 25115 4543 25149
rect 4543 25115 4569 25149
rect 2663 25012 4569 25115
rect 8050 25365 8084 25399
rect 8184 25355 8218 25389
rect 8050 25293 8084 25327
rect 8184 25283 8218 25317
rect 8050 25221 8084 25255
rect 8184 25211 8218 25245
rect 8050 25149 8084 25183
rect 8184 25139 8218 25173
rect 5251 25078 5255 25112
rect 5255 25078 5285 25112
rect 5325 25078 5359 25112
rect 5399 25078 5429 25112
rect 5429 25078 5433 25112
rect 5473 25078 5499 25112
rect 5499 25078 5507 25112
rect 5547 25078 5569 25112
rect 5569 25078 5581 25112
rect 5621 25078 5639 25112
rect 5639 25078 5655 25112
rect 5695 25078 5709 25112
rect 5709 25078 5729 25112
rect 5769 25078 5779 25112
rect 5779 25078 5803 25112
rect 5843 25078 5849 25112
rect 5849 25078 5877 25112
rect 5917 25078 5919 25112
rect 5919 25078 5951 25112
rect 5991 25078 6023 25112
rect 6023 25078 6025 25112
rect 6065 25078 6092 25112
rect 6092 25078 6099 25112
rect 6139 25078 6161 25112
rect 6161 25078 6173 25112
rect 6213 25078 6230 25112
rect 6230 25078 6247 25112
rect 6287 25078 6299 25112
rect 6299 25078 6321 25112
rect 6361 25078 6368 25112
rect 6368 25078 6395 25112
rect 6435 25078 6437 25112
rect 6437 25078 6469 25112
rect 6509 25078 6540 25112
rect 6540 25078 6543 25112
rect 6583 25078 6609 25112
rect 6609 25078 6617 25112
rect 6657 25078 6678 25112
rect 6678 25078 6691 25112
rect 6731 25078 6747 25112
rect 6747 25078 6765 25112
rect 6805 25078 6816 25112
rect 6816 25078 6839 25112
rect 6879 25078 6885 25112
rect 6885 25078 6913 25112
rect 6953 25078 6954 25112
rect 6954 25078 6987 25112
rect 7026 25078 7058 25112
rect 7058 25078 7060 25112
rect 7099 25078 7127 25112
rect 7127 25078 7133 25112
rect 7172 25078 7196 25112
rect 7196 25078 7206 25112
rect 7245 25078 7265 25112
rect 7265 25078 7279 25112
rect 7318 25078 7334 25112
rect 7334 25078 7352 25112
rect 7391 25078 7403 25112
rect 7403 25078 7425 25112
rect 7464 25078 7472 25112
rect 7472 25078 7498 25112
rect 7537 25078 7541 25112
rect 7541 25078 7571 25112
rect 7610 25078 7644 25112
rect 7683 25078 7713 25112
rect 7713 25078 7717 25112
rect 2663 24978 2715 25012
rect 2715 24978 2749 25012
rect 2749 24978 2853 25012
rect 2853 24978 2887 25012
rect 2887 24978 2991 25012
rect 2991 24978 3025 25012
rect 3025 24978 3129 25012
rect 3129 24978 3163 25012
rect 3163 24978 3267 25012
rect 3267 24978 3301 25012
rect 3301 24978 3405 25012
rect 3405 24978 3439 25012
rect 3439 24978 3543 25012
rect 3543 24978 3577 25012
rect 3577 24978 3681 25012
rect 3681 24978 3715 25012
rect 3715 24978 3819 25012
rect 3819 24978 3853 25012
rect 3853 24978 3957 25012
rect 3957 24978 3991 25012
rect 3991 24978 4095 25012
rect 4095 24978 4129 25012
rect 4129 24978 4233 25012
rect 4233 24978 4267 25012
rect 4267 24978 4371 25012
rect 4371 24978 4405 25012
rect 4405 24978 4509 25012
rect 4509 24978 4543 25012
rect 4543 24978 4569 25012
rect 2663 24875 4569 24978
rect 2663 24841 2715 24875
rect 2715 24841 2749 24875
rect 2749 24841 2853 24875
rect 2853 24841 2887 24875
rect 2887 24841 2991 24875
rect 2991 24841 3025 24875
rect 3025 24841 3129 24875
rect 3129 24841 3163 24875
rect 3163 24841 3267 24875
rect 3267 24841 3301 24875
rect 3301 24841 3405 24875
rect 3405 24841 3439 24875
rect 3439 24841 3543 24875
rect 3543 24841 3577 24875
rect 3577 24841 3681 24875
rect 3681 24841 3715 24875
rect 3715 24841 3819 24875
rect 3819 24841 3853 24875
rect 3853 24841 3957 24875
rect 3957 24841 3991 24875
rect 3991 24841 4095 24875
rect 4095 24841 4129 24875
rect 4129 24841 4233 24875
rect 4233 24841 4267 24875
rect 4267 24841 4371 24875
rect 4371 24841 4405 24875
rect 4405 24841 4509 24875
rect 4509 24841 4543 24875
rect 4543 24841 4569 24875
rect 2663 24738 4569 24841
rect 2663 24704 2715 24738
rect 2715 24704 2749 24738
rect 2749 24704 2853 24738
rect 2853 24704 2887 24738
rect 2887 24704 2991 24738
rect 2991 24704 3025 24738
rect 3025 24704 3129 24738
rect 3129 24704 3163 24738
rect 3163 24704 3267 24738
rect 3267 24704 3301 24738
rect 3301 24704 3405 24738
rect 3405 24704 3439 24738
rect 3439 24704 3543 24738
rect 3543 24704 3577 24738
rect 3577 24704 3681 24738
rect 3681 24704 3715 24738
rect 3715 24704 3819 24738
rect 3819 24704 3853 24738
rect 3853 24704 3957 24738
rect 3957 24704 3991 24738
rect 3991 24704 4095 24738
rect 4095 24704 4129 24738
rect 4129 24704 4233 24738
rect 4233 24704 4267 24738
rect 4267 24704 4371 24738
rect 4371 24704 4405 24738
rect 4405 24704 4509 24738
rect 4509 24704 4543 24738
rect 4543 24704 4569 24738
rect 8050 25077 8084 25111
rect 8184 25067 8218 25101
rect 8050 25005 8084 25039
rect 8184 24995 8218 25029
rect 8050 24933 8084 24967
rect 8184 24923 8218 24957
rect 8050 24861 8084 24895
rect 8184 24851 8218 24885
rect 8050 24789 8084 24823
rect 8184 24779 8218 24813
rect 8050 24717 8084 24751
rect 2663 24601 4569 24704
rect 2663 24567 2715 24601
rect 2715 24567 2749 24601
rect 2749 24567 2853 24601
rect 2853 24567 2887 24601
rect 2887 24567 2991 24601
rect 2991 24567 3025 24601
rect 3025 24567 3129 24601
rect 3129 24567 3163 24601
rect 3163 24567 3267 24601
rect 3267 24567 3301 24601
rect 3301 24567 3405 24601
rect 3405 24567 3439 24601
rect 3439 24567 3543 24601
rect 3543 24567 3577 24601
rect 3577 24567 3681 24601
rect 3681 24567 3715 24601
rect 3715 24567 3819 24601
rect 3819 24567 3853 24601
rect 3853 24567 3957 24601
rect 3957 24567 3991 24601
rect 3991 24567 4095 24601
rect 4095 24567 4129 24601
rect 4129 24567 4233 24601
rect 4233 24567 4267 24601
rect 4267 24567 4371 24601
rect 4371 24567 4405 24601
rect 4405 24567 4509 24601
rect 4509 24567 4543 24601
rect 4543 24567 4569 24601
rect 2663 24464 4569 24567
rect 2663 24430 2715 24464
rect 2715 24430 2749 24464
rect 2749 24430 2853 24464
rect 2853 24430 2887 24464
rect 2887 24430 2991 24464
rect 2991 24430 3025 24464
rect 3025 24430 3129 24464
rect 3129 24430 3163 24464
rect 3163 24430 3267 24464
rect 3267 24430 3301 24464
rect 3301 24430 3405 24464
rect 3405 24430 3439 24464
rect 3439 24430 3543 24464
rect 3543 24430 3577 24464
rect 3577 24430 3681 24464
rect 3681 24430 3715 24464
rect 3715 24430 3819 24464
rect 3819 24430 3853 24464
rect 3853 24430 3957 24464
rect 3957 24430 3991 24464
rect 3991 24430 4095 24464
rect 4095 24430 4129 24464
rect 4129 24430 4233 24464
rect 4233 24430 4267 24464
rect 4267 24430 4371 24464
rect 4371 24430 4405 24464
rect 4405 24430 4509 24464
rect 4509 24430 4543 24464
rect 4543 24430 4569 24464
rect 2663 24327 4569 24430
rect 2663 24293 2715 24327
rect 2715 24293 2749 24327
rect 2749 24293 2853 24327
rect 2853 24293 2887 24327
rect 2887 24293 2991 24327
rect 2991 24293 3025 24327
rect 3025 24293 3129 24327
rect 3129 24293 3163 24327
rect 3163 24293 3267 24327
rect 3267 24293 3301 24327
rect 3301 24293 3405 24327
rect 3405 24293 3439 24327
rect 3439 24293 3543 24327
rect 3543 24293 3577 24327
rect 3577 24293 3681 24327
rect 3681 24293 3715 24327
rect 3715 24293 3819 24327
rect 3819 24293 3853 24327
rect 3853 24293 3957 24327
rect 3957 24293 3991 24327
rect 3991 24293 4095 24327
rect 4095 24293 4129 24327
rect 4129 24293 4233 24327
rect 4233 24293 4267 24327
rect 4267 24293 4371 24327
rect 4371 24293 4405 24327
rect 4405 24293 4509 24327
rect 4509 24293 4543 24327
rect 4543 24293 4569 24327
rect 2663 24190 4569 24293
rect 2663 24156 2715 24190
rect 2715 24156 2749 24190
rect 2749 24156 2853 24190
rect 2853 24156 2887 24190
rect 2887 24156 2991 24190
rect 2991 24156 3025 24190
rect 3025 24156 3129 24190
rect 3129 24156 3163 24190
rect 3163 24156 3267 24190
rect 3267 24156 3301 24190
rect 3301 24156 3405 24190
rect 3405 24156 3439 24190
rect 3439 24156 3543 24190
rect 3543 24156 3577 24190
rect 3577 24156 3681 24190
rect 3681 24156 3715 24190
rect 3715 24156 3819 24190
rect 3819 24156 3853 24190
rect 3853 24156 3957 24190
rect 3957 24156 3991 24190
rect 3991 24156 4095 24190
rect 4095 24156 4129 24190
rect 4129 24156 4233 24190
rect 4233 24156 4267 24190
rect 4267 24156 4371 24190
rect 4371 24156 4405 24190
rect 4405 24156 4509 24190
rect 4509 24156 4543 24190
rect 4543 24156 4569 24190
rect 2663 24053 4569 24156
rect 2663 24019 2715 24053
rect 2715 24019 2749 24053
rect 2749 24019 2853 24053
rect 2853 24019 2887 24053
rect 2887 24019 2991 24053
rect 2991 24019 3025 24053
rect 3025 24019 3129 24053
rect 3129 24019 3163 24053
rect 3163 24019 3267 24053
rect 3267 24019 3301 24053
rect 3301 24019 3405 24053
rect 3405 24019 3439 24053
rect 3439 24019 3543 24053
rect 3543 24019 3577 24053
rect 3577 24019 3681 24053
rect 3681 24019 3715 24053
rect 3715 24019 3819 24053
rect 3819 24019 3853 24053
rect 3853 24019 3957 24053
rect 3957 24019 3991 24053
rect 3991 24019 4095 24053
rect 4095 24019 4129 24053
rect 4129 24019 4233 24053
rect 4233 24019 4267 24053
rect 4267 24019 4371 24053
rect 4371 24019 4405 24053
rect 4405 24019 4509 24053
rect 4509 24019 4543 24053
rect 4543 24019 4569 24053
rect 2663 23916 4569 24019
rect 2663 23882 2715 23916
rect 2715 23882 2749 23916
rect 2749 23882 2853 23916
rect 2853 23882 2887 23916
rect 2887 23882 2991 23916
rect 2991 23882 3025 23916
rect 3025 23882 3129 23916
rect 3129 23882 3163 23916
rect 3163 23882 3267 23916
rect 3267 23882 3301 23916
rect 3301 23882 3405 23916
rect 3405 23882 3439 23916
rect 3439 23882 3543 23916
rect 3543 23882 3577 23916
rect 3577 23882 3681 23916
rect 3681 23882 3715 23916
rect 3715 23882 3819 23916
rect 3819 23882 3853 23916
rect 3853 23882 3957 23916
rect 3957 23882 3991 23916
rect 3991 23882 4095 23916
rect 4095 23882 4129 23916
rect 4129 23882 4233 23916
rect 4233 23882 4267 23916
rect 4267 23882 4371 23916
rect 4371 23882 4405 23916
rect 4405 23882 4509 23916
rect 4509 23882 4543 23916
rect 4543 23882 4569 23916
rect 2663 23779 4569 23882
rect 2663 23745 2715 23779
rect 2715 23745 2749 23779
rect 2749 23745 2853 23779
rect 2853 23745 2887 23779
rect 2887 23745 2991 23779
rect 2991 23745 3025 23779
rect 3025 23745 3129 23779
rect 3129 23745 3163 23779
rect 3163 23745 3267 23779
rect 3267 23745 3301 23779
rect 3301 23745 3405 23779
rect 3405 23745 3439 23779
rect 3439 23745 3543 23779
rect 3543 23745 3577 23779
rect 3577 23745 3681 23779
rect 3681 23745 3715 23779
rect 3715 23745 3819 23779
rect 3819 23745 3853 23779
rect 3853 23745 3957 23779
rect 3957 23745 3991 23779
rect 3991 23745 4095 23779
rect 4095 23745 4129 23779
rect 4129 23745 4233 23779
rect 4233 23745 4267 23779
rect 4267 23745 4371 23779
rect 4371 23745 4405 23779
rect 4405 23745 4509 23779
rect 4509 23745 4543 23779
rect 4543 23745 4569 23779
rect 2663 23642 4569 23745
rect 2663 23608 2715 23642
rect 2715 23608 2749 23642
rect 2749 23608 2853 23642
rect 2853 23608 2887 23642
rect 2887 23608 2991 23642
rect 2991 23608 3025 23642
rect 3025 23608 3129 23642
rect 3129 23608 3163 23642
rect 3163 23608 3267 23642
rect 3267 23608 3301 23642
rect 3301 23608 3405 23642
rect 3405 23608 3439 23642
rect 3439 23608 3543 23642
rect 3543 23608 3577 23642
rect 3577 23608 3681 23642
rect 3681 23608 3715 23642
rect 3715 23608 3819 23642
rect 3819 23608 3853 23642
rect 3853 23608 3957 23642
rect 3957 23608 3991 23642
rect 3991 23608 4095 23642
rect 4095 23608 4129 23642
rect 4129 23608 4233 23642
rect 4233 23608 4267 23642
rect 4267 23608 4371 23642
rect 4371 23608 4405 23642
rect 4405 23608 4509 23642
rect 4509 23608 4543 23642
rect 4543 23608 4569 23642
rect 2663 23505 4569 23608
rect 2663 23471 2715 23505
rect 2715 23471 2749 23505
rect 2749 23471 2853 23505
rect 2853 23471 2887 23505
rect 2887 23471 2991 23505
rect 2991 23471 3025 23505
rect 3025 23471 3129 23505
rect 3129 23471 3163 23505
rect 3163 23471 3267 23505
rect 3267 23471 3301 23505
rect 3301 23471 3405 23505
rect 3405 23471 3439 23505
rect 3439 23471 3543 23505
rect 3543 23471 3577 23505
rect 3577 23471 3681 23505
rect 3681 23471 3715 23505
rect 3715 23471 3819 23505
rect 3819 23471 3853 23505
rect 3853 23471 3957 23505
rect 3957 23471 3991 23505
rect 3991 23471 4095 23505
rect 4095 23471 4129 23505
rect 4129 23471 4233 23505
rect 4233 23471 4267 23505
rect 4267 23471 4371 23505
rect 4371 23471 4405 23505
rect 4405 23471 4509 23505
rect 4509 23471 4543 23505
rect 4543 23471 4569 23505
rect 2663 23368 4569 23471
rect 5046 24680 5080 24714
rect 5118 24680 5152 24714
rect 5046 24607 5080 24641
rect 5118 24607 5152 24641
rect 5046 24534 5080 24568
rect 5118 24534 5152 24568
rect 5046 24461 5080 24495
rect 5118 24461 5152 24495
rect 5046 23380 5152 24422
rect 5323 24680 5357 24714
rect 5395 24680 5429 24714
rect 5323 24607 5357 24641
rect 5395 24607 5429 24641
rect 5323 24534 5357 24568
rect 5395 24534 5429 24568
rect 5323 24461 5357 24495
rect 5395 24461 5429 24495
rect 5323 23380 5429 24422
rect 5600 24680 5634 24714
rect 5672 24680 5706 24714
rect 5600 24607 5634 24641
rect 5672 24607 5706 24641
rect 5600 24534 5634 24568
rect 5672 24534 5706 24568
rect 5600 24461 5634 24495
rect 5672 24461 5706 24495
rect 5600 23380 5706 24422
rect 5877 24680 5911 24714
rect 5949 24680 5983 24714
rect 5877 24607 5911 24641
rect 5949 24607 5983 24641
rect 5877 24534 5911 24568
rect 5949 24534 5983 24568
rect 5877 24461 5911 24495
rect 5949 24461 5983 24495
rect 5877 23380 5983 24422
rect 6154 24680 6188 24714
rect 6226 24680 6260 24714
rect 6154 24607 6188 24641
rect 6226 24607 6260 24641
rect 6154 24534 6188 24568
rect 6226 24534 6260 24568
rect 6154 24461 6188 24495
rect 6226 24461 6260 24495
rect 6154 23380 6260 24422
rect 6431 24680 6465 24714
rect 6503 24680 6537 24714
rect 6431 24607 6465 24641
rect 6503 24607 6537 24641
rect 6431 24534 6465 24568
rect 6503 24534 6537 24568
rect 6431 24461 6465 24495
rect 6503 24461 6537 24495
rect 6431 23380 6537 24422
rect 6708 24680 6742 24714
rect 6780 24680 6814 24714
rect 6708 24607 6742 24641
rect 6780 24607 6814 24641
rect 6708 24534 6742 24568
rect 6780 24534 6814 24568
rect 6708 24461 6742 24495
rect 6780 24461 6814 24495
rect 6708 23380 6814 24422
rect 6985 24680 7019 24714
rect 7057 24680 7091 24714
rect 6985 24607 7019 24641
rect 7057 24607 7091 24641
rect 6985 24534 7019 24568
rect 7057 24534 7091 24568
rect 6985 24461 7019 24495
rect 7057 24461 7091 24495
rect 6985 23380 7091 24422
rect 7262 24680 7296 24714
rect 7334 24680 7368 24714
rect 7262 24607 7296 24641
rect 7334 24607 7368 24641
rect 7262 24534 7296 24568
rect 7334 24534 7368 24568
rect 7262 24461 7296 24495
rect 7334 24461 7368 24495
rect 7262 23380 7368 24422
rect 7539 24680 7573 24714
rect 7611 24680 7645 24714
rect 7539 24607 7573 24641
rect 7611 24607 7645 24641
rect 7539 24534 7573 24568
rect 7611 24534 7645 24568
rect 7539 24461 7573 24495
rect 7611 24461 7645 24495
rect 7539 23380 7645 24422
rect 7816 24680 7850 24714
rect 7888 24680 7922 24714
rect 7816 24607 7850 24641
rect 7888 24607 7922 24641
rect 7816 24534 7850 24568
rect 7888 24534 7922 24568
rect 7816 24461 7850 24495
rect 7888 24461 7922 24495
rect 7816 23380 7922 24422
rect 8184 24707 8218 24741
rect 8050 24645 8084 24679
rect 8184 24635 8218 24669
rect 8050 24573 8084 24607
rect 8184 24563 8218 24597
rect 8050 24501 8084 24535
rect 8184 24491 8218 24525
rect 8050 24429 8084 24463
rect 8184 24419 8218 24453
rect 8050 24357 8084 24391
rect 8184 24347 8218 24381
rect 8050 24285 8084 24319
rect 8184 24275 8218 24309
rect 8050 24213 8084 24247
rect 8184 24203 8218 24237
rect 8050 24141 8084 24175
rect 8184 24131 8218 24165
rect 8050 24069 8084 24103
rect 8184 24059 8218 24093
rect 8050 23997 8084 24031
rect 8184 23987 8218 24021
rect 8050 23925 8084 23959
rect 8184 23915 8218 23949
rect 8050 23853 8084 23887
rect 8184 23843 8218 23877
rect 8050 23781 8084 23815
rect 8184 23771 8218 23805
rect 8050 23709 8084 23743
rect 8184 23699 8218 23733
rect 8050 23637 8084 23671
rect 8184 23627 8218 23661
rect 8050 23565 8084 23599
rect 8184 23555 8218 23589
rect 8050 23493 8084 23527
rect 8184 23483 8218 23517
rect 8050 23421 8084 23455
rect 8184 23411 8218 23445
rect 2663 23334 2715 23368
rect 2715 23334 2749 23368
rect 2749 23334 2853 23368
rect 2853 23334 2887 23368
rect 2887 23334 2991 23368
rect 2991 23334 3025 23368
rect 3025 23334 3129 23368
rect 3129 23334 3163 23368
rect 3163 23334 3267 23368
rect 3267 23334 3301 23368
rect 3301 23334 3405 23368
rect 3405 23334 3439 23368
rect 3439 23334 3543 23368
rect 3543 23334 3577 23368
rect 3577 23334 3681 23368
rect 3681 23334 3715 23368
rect 3715 23334 3819 23368
rect 3819 23334 3853 23368
rect 3853 23334 3957 23368
rect 3957 23334 3991 23368
rect 3991 23334 4095 23368
rect 4095 23334 4129 23368
rect 4129 23334 4233 23368
rect 4233 23334 4267 23368
rect 4267 23334 4371 23368
rect 4371 23334 4405 23368
rect 4405 23334 4509 23368
rect 4509 23334 4543 23368
rect 4543 23334 4569 23368
rect 2663 23231 4569 23334
rect 2663 23197 2715 23231
rect 2715 23197 2749 23231
rect 2749 23197 2853 23231
rect 2853 23197 2887 23231
rect 2887 23197 2991 23231
rect 2991 23197 3025 23231
rect 3025 23197 3129 23231
rect 3129 23197 3163 23231
rect 3163 23197 3267 23231
rect 3267 23197 3301 23231
rect 3301 23197 3405 23231
rect 3405 23197 3439 23231
rect 3439 23197 3543 23231
rect 3543 23197 3577 23231
rect 3577 23197 3681 23231
rect 3681 23197 3715 23231
rect 3715 23197 3819 23231
rect 3819 23197 3853 23231
rect 3853 23197 3957 23231
rect 3957 23197 3991 23231
rect 3991 23197 4095 23231
rect 4095 23197 4129 23231
rect 4129 23197 4233 23231
rect 4233 23197 4267 23231
rect 4267 23197 4371 23231
rect 4371 23197 4405 23231
rect 4405 23197 4509 23231
rect 4509 23197 4543 23231
rect 4543 23197 4569 23231
rect 2663 23094 4569 23197
rect 8050 23349 8084 23383
rect 8184 23339 8218 23373
rect 8050 23277 8084 23311
rect 8184 23267 8218 23301
rect 8050 23205 8084 23239
rect 8184 23195 8218 23229
rect 8050 23133 8084 23167
rect 2663 23060 2715 23094
rect 2715 23060 2749 23094
rect 2749 23060 2853 23094
rect 2853 23060 2887 23094
rect 2887 23060 2991 23094
rect 2991 23060 3025 23094
rect 3025 23060 3129 23094
rect 3129 23060 3163 23094
rect 3163 23060 3267 23094
rect 3267 23060 3301 23094
rect 3301 23060 3405 23094
rect 3405 23060 3439 23094
rect 3439 23060 3543 23094
rect 3543 23060 3577 23094
rect 3577 23060 3681 23094
rect 3681 23060 3715 23094
rect 3715 23060 3819 23094
rect 3819 23060 3853 23094
rect 3853 23060 3957 23094
rect 3957 23060 3991 23094
rect 3991 23060 4095 23094
rect 4095 23060 4129 23094
rect 4129 23060 4233 23094
rect 4233 23060 4267 23094
rect 4267 23060 4371 23094
rect 4371 23060 4405 23094
rect 4405 23060 4509 23094
rect 4509 23060 4543 23094
rect 4543 23060 4569 23094
rect 5251 23090 5255 23124
rect 5255 23090 5285 23124
rect 5325 23090 5359 23124
rect 5399 23090 5429 23124
rect 5429 23090 5433 23124
rect 5473 23090 5499 23124
rect 5499 23090 5507 23124
rect 5547 23090 5569 23124
rect 5569 23090 5581 23124
rect 5621 23090 5639 23124
rect 5639 23090 5655 23124
rect 5695 23090 5709 23124
rect 5709 23090 5729 23124
rect 5769 23090 5779 23124
rect 5779 23090 5803 23124
rect 5843 23090 5849 23124
rect 5849 23090 5877 23124
rect 5917 23090 5919 23124
rect 5919 23090 5951 23124
rect 5991 23090 6023 23124
rect 6023 23090 6025 23124
rect 6065 23090 6092 23124
rect 6092 23090 6099 23124
rect 6139 23090 6161 23124
rect 6161 23090 6173 23124
rect 6213 23090 6230 23124
rect 6230 23090 6247 23124
rect 6287 23090 6299 23124
rect 6299 23090 6321 23124
rect 6361 23090 6368 23124
rect 6368 23090 6395 23124
rect 6435 23090 6437 23124
rect 6437 23090 6469 23124
rect 6509 23090 6540 23124
rect 6540 23090 6543 23124
rect 6583 23090 6609 23124
rect 6609 23090 6617 23124
rect 6657 23090 6678 23124
rect 6678 23090 6691 23124
rect 6731 23090 6747 23124
rect 6747 23090 6765 23124
rect 6805 23090 6816 23124
rect 6816 23090 6839 23124
rect 6879 23090 6885 23124
rect 6885 23090 6913 23124
rect 6953 23090 6954 23124
rect 6954 23090 6987 23124
rect 7026 23090 7058 23124
rect 7058 23090 7060 23124
rect 7099 23090 7127 23124
rect 7127 23090 7133 23124
rect 7172 23090 7196 23124
rect 7196 23090 7206 23124
rect 7245 23090 7265 23124
rect 7265 23090 7279 23124
rect 7318 23090 7334 23124
rect 7334 23090 7352 23124
rect 7391 23090 7403 23124
rect 7403 23090 7425 23124
rect 7464 23090 7472 23124
rect 7472 23090 7498 23124
rect 7537 23090 7541 23124
rect 7541 23090 7571 23124
rect 7610 23090 7644 23124
rect 7683 23090 7713 23124
rect 7713 23090 7717 23124
rect 8184 23123 8218 23157
rect 2663 22957 4569 23060
rect 2663 22923 2715 22957
rect 2715 22923 2749 22957
rect 2749 22923 2853 22957
rect 2853 22923 2887 22957
rect 2887 22923 2991 22957
rect 2991 22923 3025 22957
rect 3025 22923 3129 22957
rect 3129 22923 3163 22957
rect 3163 22923 3267 22957
rect 3267 22923 3301 22957
rect 3301 22923 3405 22957
rect 3405 22923 3439 22957
rect 3439 22923 3543 22957
rect 3543 22923 3577 22957
rect 3577 22923 3681 22957
rect 3681 22923 3715 22957
rect 3715 22923 3819 22957
rect 3819 22923 3853 22957
rect 3853 22923 3957 22957
rect 3957 22923 3991 22957
rect 3991 22923 4095 22957
rect 4095 22923 4129 22957
rect 4129 22923 4233 22957
rect 4233 22923 4267 22957
rect 4267 22923 4371 22957
rect 4371 22923 4405 22957
rect 4405 22923 4509 22957
rect 4509 22923 4543 22957
rect 4543 22923 4569 22957
rect 2663 22820 4569 22923
rect 2663 22786 2715 22820
rect 2715 22786 2749 22820
rect 2749 22786 2853 22820
rect 2853 22786 2887 22820
rect 2887 22786 2991 22820
rect 2991 22786 3025 22820
rect 3025 22786 3129 22820
rect 3129 22786 3163 22820
rect 3163 22786 3267 22820
rect 3267 22786 3301 22820
rect 3301 22786 3405 22820
rect 3405 22786 3439 22820
rect 3439 22786 3543 22820
rect 3543 22786 3577 22820
rect 3577 22786 3681 22820
rect 3681 22786 3715 22820
rect 3715 22786 3819 22820
rect 3819 22786 3853 22820
rect 3853 22786 3957 22820
rect 3957 22786 3991 22820
rect 3991 22786 4095 22820
rect 4095 22786 4129 22820
rect 4129 22786 4233 22820
rect 4233 22786 4267 22820
rect 4267 22786 4371 22820
rect 4371 22786 4405 22820
rect 4405 22786 4509 22820
rect 4509 22786 4543 22820
rect 4543 22786 4569 22820
rect 2663 22683 4569 22786
rect 8050 23061 8084 23095
rect 8184 23051 8218 23085
rect 8050 22989 8084 23023
rect 8184 22979 8218 23013
rect 8050 22917 8084 22951
rect 8184 22907 8218 22941
rect 8050 22845 8084 22879
rect 8184 22835 8218 22869
rect 8050 22773 8084 22807
rect 8184 22763 8218 22797
rect 2663 22649 2715 22683
rect 2715 22649 2749 22683
rect 2749 22649 2853 22683
rect 2853 22649 2887 22683
rect 2887 22649 2991 22683
rect 2991 22649 3025 22683
rect 3025 22649 3129 22683
rect 3129 22649 3163 22683
rect 3163 22649 3267 22683
rect 3267 22649 3301 22683
rect 3301 22649 3405 22683
rect 3405 22649 3439 22683
rect 3439 22649 3543 22683
rect 3543 22649 3577 22683
rect 3577 22649 3681 22683
rect 3681 22649 3715 22683
rect 3715 22649 3819 22683
rect 3819 22649 3853 22683
rect 3853 22649 3957 22683
rect 3957 22649 3991 22683
rect 3991 22649 4095 22683
rect 4095 22649 4129 22683
rect 4129 22649 4233 22683
rect 4233 22649 4267 22683
rect 4267 22649 4371 22683
rect 4371 22649 4405 22683
rect 4405 22649 4509 22683
rect 4509 22649 4543 22683
rect 4543 22649 4569 22683
rect 2663 22546 4569 22649
rect 2663 22512 2715 22546
rect 2715 22512 2749 22546
rect 2749 22512 2853 22546
rect 2853 22512 2887 22546
rect 2887 22512 2991 22546
rect 2991 22512 3025 22546
rect 3025 22512 3129 22546
rect 3129 22512 3163 22546
rect 3163 22512 3267 22546
rect 3267 22512 3301 22546
rect 3301 22512 3405 22546
rect 3405 22512 3439 22546
rect 3439 22512 3543 22546
rect 3543 22512 3577 22546
rect 3577 22512 3681 22546
rect 3681 22512 3715 22546
rect 3715 22512 3819 22546
rect 3819 22512 3853 22546
rect 3853 22512 3957 22546
rect 3957 22512 3991 22546
rect 3991 22512 4095 22546
rect 4095 22512 4129 22546
rect 4129 22512 4233 22546
rect 4233 22512 4267 22546
rect 4267 22512 4371 22546
rect 4371 22512 4405 22546
rect 4405 22512 4509 22546
rect 4509 22512 4543 22546
rect 4543 22512 4569 22546
rect 2663 22409 4569 22512
rect 2663 22375 2715 22409
rect 2715 22375 2749 22409
rect 2749 22375 2853 22409
rect 2853 22375 2887 22409
rect 2887 22375 2991 22409
rect 2991 22375 3025 22409
rect 3025 22375 3129 22409
rect 3129 22375 3163 22409
rect 3163 22375 3267 22409
rect 3267 22375 3301 22409
rect 3301 22375 3405 22409
rect 3405 22375 3439 22409
rect 3439 22375 3543 22409
rect 3543 22375 3577 22409
rect 3577 22375 3681 22409
rect 3681 22375 3715 22409
rect 3715 22375 3819 22409
rect 3819 22375 3853 22409
rect 3853 22375 3957 22409
rect 3957 22375 3991 22409
rect 3991 22375 4095 22409
rect 4095 22375 4129 22409
rect 4129 22375 4233 22409
rect 4233 22375 4267 22409
rect 4267 22375 4371 22409
rect 4371 22375 4405 22409
rect 4405 22375 4509 22409
rect 4509 22375 4543 22409
rect 4543 22375 4569 22409
rect 2663 22272 4569 22375
rect 2663 22238 2715 22272
rect 2715 22238 2749 22272
rect 2749 22238 2853 22272
rect 2853 22238 2887 22272
rect 2887 22238 2991 22272
rect 2991 22238 3025 22272
rect 3025 22238 3129 22272
rect 3129 22238 3163 22272
rect 3163 22238 3267 22272
rect 3267 22238 3301 22272
rect 3301 22238 3405 22272
rect 3405 22238 3439 22272
rect 3439 22238 3543 22272
rect 3543 22238 3577 22272
rect 3577 22238 3681 22272
rect 3681 22238 3715 22272
rect 3715 22238 3819 22272
rect 3819 22238 3853 22272
rect 3853 22238 3957 22272
rect 3957 22238 3991 22272
rect 3991 22238 4095 22272
rect 4095 22238 4129 22272
rect 4129 22238 4233 22272
rect 4233 22238 4267 22272
rect 4267 22238 4371 22272
rect 4371 22238 4405 22272
rect 4405 22238 4509 22272
rect 4509 22238 4543 22272
rect 4543 22238 4569 22272
rect 2663 22135 4569 22238
rect 2663 22101 2715 22135
rect 2715 22101 2749 22135
rect 2749 22101 2853 22135
rect 2853 22101 2887 22135
rect 2887 22101 2991 22135
rect 2991 22101 3025 22135
rect 3025 22101 3129 22135
rect 3129 22101 3163 22135
rect 3163 22101 3267 22135
rect 3267 22101 3301 22135
rect 3301 22101 3405 22135
rect 3405 22101 3439 22135
rect 3439 22101 3543 22135
rect 3543 22101 3577 22135
rect 3577 22101 3681 22135
rect 3681 22101 3715 22135
rect 3715 22101 3819 22135
rect 3819 22101 3853 22135
rect 3853 22101 3957 22135
rect 3957 22101 3991 22135
rect 3991 22101 4095 22135
rect 4095 22101 4129 22135
rect 4129 22101 4233 22135
rect 4233 22101 4267 22135
rect 4267 22101 4371 22135
rect 4371 22101 4405 22135
rect 4405 22101 4509 22135
rect 4509 22101 4543 22135
rect 4543 22101 4569 22135
rect 2663 21998 4569 22101
rect 2663 21964 2715 21998
rect 2715 21964 2749 21998
rect 2749 21964 2853 21998
rect 2853 21964 2887 21998
rect 2887 21964 2991 21998
rect 2991 21964 3025 21998
rect 3025 21964 3129 21998
rect 3129 21964 3163 21998
rect 3163 21964 3267 21998
rect 3267 21964 3301 21998
rect 3301 21964 3405 21998
rect 3405 21964 3439 21998
rect 3439 21964 3543 21998
rect 3543 21964 3577 21998
rect 3577 21964 3681 21998
rect 3681 21964 3715 21998
rect 3715 21964 3819 21998
rect 3819 21964 3853 21998
rect 3853 21964 3957 21998
rect 3957 21964 3991 21998
rect 3991 21964 4095 21998
rect 4095 21964 4129 21998
rect 4129 21964 4233 21998
rect 4233 21964 4267 21998
rect 4267 21964 4371 21998
rect 4371 21964 4405 21998
rect 4405 21964 4509 21998
rect 4509 21964 4543 21998
rect 4543 21964 4569 21998
rect 2663 21861 4569 21964
rect 2663 21827 2715 21861
rect 2715 21827 2749 21861
rect 2749 21827 2853 21861
rect 2853 21827 2887 21861
rect 2887 21827 2991 21861
rect 2991 21827 3025 21861
rect 3025 21827 3129 21861
rect 3129 21827 3163 21861
rect 3163 21827 3267 21861
rect 3267 21827 3301 21861
rect 3301 21827 3405 21861
rect 3405 21827 3439 21861
rect 3439 21827 3543 21861
rect 3543 21827 3577 21861
rect 3577 21827 3681 21861
rect 3681 21827 3715 21861
rect 3715 21827 3819 21861
rect 3819 21827 3853 21861
rect 3853 21827 3957 21861
rect 3957 21827 3991 21861
rect 3991 21827 4095 21861
rect 4095 21827 4129 21861
rect 4129 21827 4233 21861
rect 4233 21827 4267 21861
rect 4267 21827 4371 21861
rect 4371 21827 4405 21861
rect 4405 21827 4509 21861
rect 4509 21827 4543 21861
rect 4543 21827 4569 21861
rect 2663 21724 4569 21827
rect 2663 21690 2715 21724
rect 2715 21690 2749 21724
rect 2749 21690 2853 21724
rect 2853 21690 2887 21724
rect 2887 21690 2991 21724
rect 2991 21690 3025 21724
rect 3025 21690 3129 21724
rect 3129 21690 3163 21724
rect 3163 21690 3267 21724
rect 3267 21690 3301 21724
rect 3301 21690 3405 21724
rect 3405 21690 3439 21724
rect 3439 21690 3543 21724
rect 3543 21690 3577 21724
rect 3577 21690 3681 21724
rect 3681 21690 3715 21724
rect 3715 21690 3819 21724
rect 3819 21690 3853 21724
rect 3853 21690 3957 21724
rect 3957 21690 3991 21724
rect 3991 21690 4095 21724
rect 4095 21690 4129 21724
rect 4129 21690 4233 21724
rect 4233 21690 4267 21724
rect 4267 21690 4371 21724
rect 4371 21690 4405 21724
rect 4405 21690 4509 21724
rect 4509 21690 4543 21724
rect 4543 21690 4569 21724
rect 2663 21587 4569 21690
rect 2663 21553 2715 21587
rect 2715 21553 2749 21587
rect 2749 21553 2853 21587
rect 2853 21553 2887 21587
rect 2887 21553 2991 21587
rect 2991 21553 3025 21587
rect 3025 21553 3129 21587
rect 3129 21553 3163 21587
rect 3163 21553 3267 21587
rect 3267 21553 3301 21587
rect 3301 21553 3405 21587
rect 3405 21553 3439 21587
rect 3439 21553 3543 21587
rect 3543 21553 3577 21587
rect 3577 21553 3681 21587
rect 3681 21553 3715 21587
rect 3715 21553 3819 21587
rect 3819 21553 3853 21587
rect 3853 21553 3957 21587
rect 3957 21553 3991 21587
rect 3991 21553 4095 21587
rect 4095 21553 4129 21587
rect 4129 21553 4233 21587
rect 4233 21553 4267 21587
rect 4267 21553 4371 21587
rect 4371 21553 4405 21587
rect 4405 21553 4509 21587
rect 4509 21553 4543 21587
rect 4543 21553 4569 21587
rect 2663 21450 4569 21553
rect 2663 21416 2715 21450
rect 2715 21416 2749 21450
rect 2749 21416 2853 21450
rect 2853 21416 2887 21450
rect 2887 21416 2991 21450
rect 2991 21416 3025 21450
rect 3025 21416 3129 21450
rect 3129 21416 3163 21450
rect 3163 21416 3267 21450
rect 3267 21416 3301 21450
rect 3301 21416 3405 21450
rect 3405 21416 3439 21450
rect 3439 21416 3543 21450
rect 3543 21416 3577 21450
rect 3577 21416 3681 21450
rect 3681 21416 3715 21450
rect 3715 21416 3819 21450
rect 3819 21416 3853 21450
rect 3853 21416 3957 21450
rect 3957 21416 3991 21450
rect 3991 21416 4095 21450
rect 4095 21416 4129 21450
rect 4129 21416 4233 21450
rect 4233 21416 4267 21450
rect 4267 21416 4371 21450
rect 4371 21416 4405 21450
rect 4405 21416 4509 21450
rect 4509 21416 4543 21450
rect 4543 21416 4569 21450
rect 2663 21313 4569 21416
rect 5046 22680 5080 22714
rect 5118 22680 5152 22714
rect 5046 22607 5080 22641
rect 5118 22607 5152 22641
rect 5046 22534 5080 22568
rect 5118 22534 5152 22568
rect 5046 22461 5080 22495
rect 5118 22461 5152 22495
rect 5046 21380 5152 22422
rect 5323 22680 5357 22714
rect 5395 22680 5429 22714
rect 5323 22607 5357 22641
rect 5395 22607 5429 22641
rect 5323 22534 5357 22568
rect 5395 22534 5429 22568
rect 5323 22461 5357 22495
rect 5395 22461 5429 22495
rect 5323 21380 5429 22422
rect 5600 22680 5634 22714
rect 5672 22680 5706 22714
rect 5600 22607 5634 22641
rect 5672 22607 5706 22641
rect 5600 22534 5634 22568
rect 5672 22534 5706 22568
rect 5600 22461 5634 22495
rect 5672 22461 5706 22495
rect 5600 21380 5706 22422
rect 5877 22680 5911 22714
rect 5949 22680 5983 22714
rect 5877 22607 5911 22641
rect 5949 22607 5983 22641
rect 5877 22534 5911 22568
rect 5949 22534 5983 22568
rect 5877 22461 5911 22495
rect 5949 22461 5983 22495
rect 5877 21380 5983 22422
rect 6154 22680 6188 22714
rect 6226 22680 6260 22714
rect 6154 22607 6188 22641
rect 6226 22607 6260 22641
rect 6154 22534 6188 22568
rect 6226 22534 6260 22568
rect 6154 22461 6188 22495
rect 6226 22461 6260 22495
rect 6154 21380 6260 22422
rect 6431 22680 6465 22714
rect 6503 22680 6537 22714
rect 6431 22607 6465 22641
rect 6503 22607 6537 22641
rect 6431 22534 6465 22568
rect 6503 22534 6537 22568
rect 6431 22461 6465 22495
rect 6503 22461 6537 22495
rect 6431 21380 6537 22422
rect 6708 22680 6742 22714
rect 6780 22680 6814 22714
rect 6708 22607 6742 22641
rect 6780 22607 6814 22641
rect 6708 22534 6742 22568
rect 6780 22534 6814 22568
rect 6708 22461 6742 22495
rect 6780 22461 6814 22495
rect 6708 21380 6814 22422
rect 6985 22680 7019 22714
rect 7057 22680 7091 22714
rect 6985 22607 7019 22641
rect 7057 22607 7091 22641
rect 6985 22534 7019 22568
rect 7057 22534 7091 22568
rect 6985 22461 7019 22495
rect 7057 22461 7091 22495
rect 6985 21380 7091 22422
rect 7262 22680 7296 22714
rect 7334 22680 7368 22714
rect 7262 22607 7296 22641
rect 7334 22607 7368 22641
rect 7262 22534 7296 22568
rect 7334 22534 7368 22568
rect 7262 22461 7296 22495
rect 7334 22461 7368 22495
rect 7262 21380 7368 22422
rect 7539 22680 7573 22714
rect 7611 22680 7645 22714
rect 7539 22607 7573 22641
rect 7611 22607 7645 22641
rect 7539 22534 7573 22568
rect 7611 22534 7645 22568
rect 7539 22461 7573 22495
rect 7611 22461 7645 22495
rect 7539 21380 7645 22422
rect 7816 22680 7850 22714
rect 7888 22680 7922 22714
rect 7816 22607 7850 22641
rect 7888 22607 7922 22641
rect 7816 22534 7850 22568
rect 7888 22534 7922 22568
rect 7816 22461 7850 22495
rect 7888 22461 7922 22495
rect 7816 21380 7922 22422
rect 8050 22701 8084 22735
rect 8184 22691 8218 22725
rect 8050 22629 8084 22663
rect 8184 22619 8218 22653
rect 8050 22557 8084 22591
rect 8184 22547 8218 22581
rect 8050 22485 8084 22519
rect 8184 22475 8218 22509
rect 8050 22413 8084 22447
rect 8184 22403 8218 22437
rect 8050 22341 8084 22375
rect 8184 22331 8218 22365
rect 8050 22269 8084 22303
rect 8184 22259 8218 22293
rect 8050 22197 8084 22231
rect 8184 22187 8218 22221
rect 8050 22125 8084 22159
rect 8184 22115 8218 22149
rect 8050 22053 8084 22087
rect 8184 22043 8218 22077
rect 8050 21981 8084 22015
rect 8184 21971 8218 22005
rect 8050 21909 8084 21943
rect 8184 21899 8218 21933
rect 8050 21837 8084 21871
rect 8184 21827 8218 21861
rect 8050 21765 8084 21799
rect 8184 21755 8218 21789
rect 8050 21693 8084 21727
rect 8184 21683 8218 21717
rect 8050 21621 8084 21655
rect 8184 21611 8218 21645
rect 8050 21549 8084 21583
rect 8184 21539 8218 21573
rect 8050 21477 8084 21511
rect 8184 21467 8218 21501
rect 8050 21405 8084 21439
rect 8184 21395 8218 21429
rect 2663 21279 2715 21313
rect 2715 21279 2749 21313
rect 2749 21279 2853 21313
rect 2853 21279 2887 21313
rect 2887 21279 2991 21313
rect 2991 21279 3025 21313
rect 3025 21279 3129 21313
rect 3129 21279 3163 21313
rect 3163 21279 3267 21313
rect 3267 21279 3301 21313
rect 3301 21279 3405 21313
rect 3405 21279 3439 21313
rect 3439 21279 3543 21313
rect 3543 21279 3577 21313
rect 3577 21279 3681 21313
rect 3681 21279 3715 21313
rect 3715 21279 3819 21313
rect 3819 21279 3853 21313
rect 3853 21279 3957 21313
rect 3957 21279 3991 21313
rect 3991 21279 4095 21313
rect 4095 21279 4129 21313
rect 4129 21279 4233 21313
rect 4233 21279 4267 21313
rect 4267 21279 4371 21313
rect 4371 21279 4405 21313
rect 4405 21279 4509 21313
rect 4509 21279 4543 21313
rect 4543 21279 4569 21313
rect 2663 21176 4569 21279
rect 2663 21142 2715 21176
rect 2715 21142 2749 21176
rect 2749 21142 2853 21176
rect 2853 21142 2887 21176
rect 2887 21142 2991 21176
rect 2991 21142 3025 21176
rect 3025 21142 3129 21176
rect 3129 21142 3163 21176
rect 3163 21142 3267 21176
rect 3267 21142 3301 21176
rect 3301 21142 3405 21176
rect 3405 21142 3439 21176
rect 3439 21142 3543 21176
rect 3543 21142 3577 21176
rect 3577 21142 3681 21176
rect 3681 21142 3715 21176
rect 3715 21142 3819 21176
rect 3819 21142 3853 21176
rect 3853 21142 3957 21176
rect 3957 21142 3991 21176
rect 3991 21142 4095 21176
rect 4095 21142 4129 21176
rect 4129 21142 4233 21176
rect 4233 21142 4267 21176
rect 4267 21142 4371 21176
rect 4371 21142 4405 21176
rect 4405 21142 4509 21176
rect 4509 21142 4543 21176
rect 4543 21142 4569 21176
rect 2663 21039 4569 21142
rect 8050 21333 8084 21367
rect 8184 21323 8218 21357
rect 8050 21261 8084 21295
rect 8184 21251 8218 21285
rect 8050 21189 8084 21223
rect 8184 21179 8218 21213
rect 8050 21117 8084 21151
rect 8184 21107 8218 21141
rect 5251 21049 5255 21083
rect 5255 21049 5285 21083
rect 5326 21049 5359 21083
rect 5359 21049 5360 21083
rect 5401 21049 5429 21083
rect 5429 21049 5435 21083
rect 5476 21049 5499 21083
rect 5499 21049 5510 21083
rect 5551 21049 5569 21083
rect 5569 21049 5585 21083
rect 5626 21049 5639 21083
rect 5639 21049 5660 21083
rect 5701 21049 5709 21083
rect 5709 21049 5735 21083
rect 5776 21049 5779 21083
rect 5779 21049 5810 21083
rect 5851 21049 5885 21083
rect 5926 21049 5954 21083
rect 5954 21049 5960 21083
rect 6001 21049 6023 21083
rect 6023 21049 6035 21083
rect 6076 21049 6092 21083
rect 6092 21049 6110 21083
rect 6151 21049 6161 21083
rect 6161 21049 6185 21083
rect 6225 21049 6230 21083
rect 6230 21049 6259 21083
rect 6299 21049 6333 21083
rect 6373 21049 6402 21083
rect 6402 21049 6407 21083
rect 6447 21049 6471 21083
rect 6471 21049 6481 21083
rect 6521 21049 6540 21083
rect 6540 21049 6555 21083
rect 6595 21049 6609 21083
rect 6609 21049 6629 21083
rect 6669 21049 6678 21083
rect 6678 21049 6703 21083
rect 6743 21049 6747 21083
rect 6747 21049 6777 21083
rect 6817 21049 6851 21083
rect 6891 21049 6920 21083
rect 6920 21049 6925 21083
rect 2663 21005 2715 21039
rect 2715 21005 2749 21039
rect 2749 21005 2853 21039
rect 2853 21005 2887 21039
rect 2887 21005 2991 21039
rect 2991 21005 3025 21039
rect 3025 21005 3129 21039
rect 3129 21005 3163 21039
rect 3163 21005 3267 21039
rect 3267 21005 3301 21039
rect 3301 21005 3405 21039
rect 3405 21005 3439 21039
rect 3439 21005 3543 21039
rect 3543 21005 3577 21039
rect 3577 21005 3681 21039
rect 3681 21005 3715 21039
rect 3715 21005 3819 21039
rect 3819 21005 3853 21039
rect 3853 21005 3957 21039
rect 3957 21005 3991 21039
rect 3991 21005 4095 21039
rect 4095 21005 4129 21039
rect 4129 21005 4233 21039
rect 4233 21005 4267 21039
rect 4267 21005 4371 21039
rect 4371 21005 4405 21039
rect 4405 21005 4509 21039
rect 4509 21005 4543 21039
rect 4543 21005 4569 21039
rect 2663 20902 4569 21005
rect 2663 20868 2715 20902
rect 2715 20868 2749 20902
rect 2749 20868 2853 20902
rect 2853 20868 2887 20902
rect 2887 20868 2991 20902
rect 2991 20868 3025 20902
rect 3025 20868 3129 20902
rect 3129 20868 3163 20902
rect 3163 20868 3267 20902
rect 3267 20868 3301 20902
rect 3301 20868 3405 20902
rect 3405 20868 3439 20902
rect 3439 20868 3543 20902
rect 3543 20868 3577 20902
rect 3577 20868 3681 20902
rect 3681 20868 3715 20902
rect 3715 20868 3819 20902
rect 3819 20868 3853 20902
rect 3853 20868 3957 20902
rect 3957 20868 3991 20902
rect 3991 20868 4095 20902
rect 4095 20868 4129 20902
rect 4129 20868 4233 20902
rect 4233 20868 4267 20902
rect 4267 20868 4371 20902
rect 4371 20868 4405 20902
rect 4405 20868 4509 20902
rect 4509 20868 4543 20902
rect 4543 20868 4569 20902
rect 2663 20765 4569 20868
rect 2663 20731 2715 20765
rect 2715 20731 2749 20765
rect 2749 20731 2853 20765
rect 2853 20731 2887 20765
rect 2887 20731 2991 20765
rect 2991 20731 3025 20765
rect 3025 20731 3129 20765
rect 3129 20731 3163 20765
rect 3163 20731 3267 20765
rect 3267 20731 3301 20765
rect 3301 20731 3405 20765
rect 3405 20731 3439 20765
rect 3439 20731 3543 20765
rect 3543 20731 3577 20765
rect 3577 20731 3681 20765
rect 3681 20731 3715 20765
rect 3715 20731 3819 20765
rect 3819 20731 3853 20765
rect 3853 20731 3957 20765
rect 3957 20731 3991 20765
rect 3991 20731 4095 20765
rect 4095 20731 4129 20765
rect 4129 20731 4233 20765
rect 4233 20731 4267 20765
rect 4267 20731 4371 20765
rect 4371 20731 4405 20765
rect 4405 20731 4509 20765
rect 4509 20731 4543 20765
rect 4543 20731 4569 20765
rect 2663 20628 4569 20731
rect 8050 21045 8084 21079
rect 8184 21035 8218 21069
rect 8050 20973 8084 21007
rect 8184 20963 8218 20997
rect 8050 20901 8084 20935
rect 8184 20891 8218 20925
rect 8050 20829 8084 20863
rect 8184 20819 8218 20853
rect 8050 20757 8084 20791
rect 8184 20747 8218 20781
rect 2663 20594 2715 20628
rect 2715 20594 2749 20628
rect 2749 20594 2853 20628
rect 2853 20594 2887 20628
rect 2887 20594 2991 20628
rect 2991 20594 3025 20628
rect 3025 20594 3129 20628
rect 3129 20594 3163 20628
rect 3163 20594 3267 20628
rect 3267 20594 3301 20628
rect 3301 20594 3405 20628
rect 3405 20594 3439 20628
rect 3439 20594 3543 20628
rect 3543 20594 3577 20628
rect 3577 20594 3681 20628
rect 3681 20594 3715 20628
rect 3715 20594 3819 20628
rect 3819 20594 3853 20628
rect 3853 20594 3957 20628
rect 3957 20594 3991 20628
rect 3991 20594 4095 20628
rect 4095 20594 4129 20628
rect 4129 20594 4233 20628
rect 4233 20594 4267 20628
rect 4267 20594 4371 20628
rect 4371 20594 4405 20628
rect 4405 20594 4509 20628
rect 4509 20594 4543 20628
rect 4543 20594 4569 20628
rect 2663 20491 4569 20594
rect 2663 20457 2715 20491
rect 2715 20457 2749 20491
rect 2749 20457 2853 20491
rect 2853 20457 2887 20491
rect 2887 20457 2991 20491
rect 2991 20457 3025 20491
rect 3025 20457 3129 20491
rect 3129 20457 3163 20491
rect 3163 20457 3267 20491
rect 3267 20457 3301 20491
rect 3301 20457 3405 20491
rect 3405 20457 3439 20491
rect 3439 20457 3543 20491
rect 3543 20457 3577 20491
rect 3577 20457 3681 20491
rect 3681 20457 3715 20491
rect 3715 20457 3819 20491
rect 3819 20457 3853 20491
rect 3853 20457 3957 20491
rect 3957 20457 3991 20491
rect 3991 20457 4095 20491
rect 4095 20457 4129 20491
rect 4129 20457 4233 20491
rect 4233 20457 4267 20491
rect 4267 20457 4371 20491
rect 4371 20457 4405 20491
rect 4405 20457 4509 20491
rect 4509 20457 4543 20491
rect 4543 20457 4569 20491
rect 2663 20354 4569 20457
rect 2663 20320 2715 20354
rect 2715 20320 2749 20354
rect 2749 20320 2853 20354
rect 2853 20320 2887 20354
rect 2887 20320 2991 20354
rect 2991 20320 3025 20354
rect 3025 20320 3129 20354
rect 3129 20320 3163 20354
rect 3163 20320 3267 20354
rect 3267 20320 3301 20354
rect 3301 20320 3405 20354
rect 3405 20320 3439 20354
rect 3439 20320 3543 20354
rect 3543 20320 3577 20354
rect 3577 20320 3681 20354
rect 3681 20320 3715 20354
rect 3715 20320 3819 20354
rect 3819 20320 3853 20354
rect 3853 20320 3957 20354
rect 3957 20320 3991 20354
rect 3991 20320 4095 20354
rect 4095 20320 4129 20354
rect 4129 20320 4233 20354
rect 4233 20320 4267 20354
rect 4267 20320 4371 20354
rect 4371 20320 4405 20354
rect 4405 20320 4509 20354
rect 4509 20320 4543 20354
rect 4543 20320 4569 20354
rect 2663 20217 4569 20320
rect 2663 20183 2715 20217
rect 2715 20183 2749 20217
rect 2749 20183 2853 20217
rect 2853 20183 2887 20217
rect 2887 20183 2991 20217
rect 2991 20183 3025 20217
rect 3025 20183 3129 20217
rect 3129 20183 3163 20217
rect 3163 20183 3267 20217
rect 3267 20183 3301 20217
rect 3301 20183 3405 20217
rect 3405 20183 3439 20217
rect 3439 20183 3543 20217
rect 3543 20183 3577 20217
rect 3577 20183 3681 20217
rect 3681 20183 3715 20217
rect 3715 20183 3819 20217
rect 3819 20183 3853 20217
rect 3853 20183 3957 20217
rect 3957 20183 3991 20217
rect 3991 20183 4095 20217
rect 4095 20183 4129 20217
rect 4129 20183 4233 20217
rect 4233 20183 4267 20217
rect 4267 20183 4371 20217
rect 4371 20183 4405 20217
rect 4405 20183 4509 20217
rect 4509 20183 4543 20217
rect 4543 20183 4569 20217
rect 2663 20080 4569 20183
rect 2663 20046 2715 20080
rect 2715 20046 2749 20080
rect 2749 20046 2853 20080
rect 2853 20046 2887 20080
rect 2887 20046 2991 20080
rect 2991 20046 3025 20080
rect 3025 20046 3129 20080
rect 3129 20046 3163 20080
rect 3163 20046 3267 20080
rect 3267 20046 3301 20080
rect 3301 20046 3405 20080
rect 3405 20046 3439 20080
rect 3439 20046 3543 20080
rect 3543 20046 3577 20080
rect 3577 20046 3681 20080
rect 3681 20046 3715 20080
rect 3715 20046 3819 20080
rect 3819 20046 3853 20080
rect 3853 20046 3957 20080
rect 3957 20046 3991 20080
rect 3991 20046 4095 20080
rect 4095 20046 4129 20080
rect 4129 20046 4233 20080
rect 4233 20046 4267 20080
rect 4267 20046 4371 20080
rect 4371 20046 4405 20080
rect 4405 20046 4509 20080
rect 4509 20046 4543 20080
rect 4543 20046 4569 20080
rect 2663 19943 4569 20046
rect 2663 19909 2715 19943
rect 2715 19909 2749 19943
rect 2749 19909 2853 19943
rect 2853 19909 2887 19943
rect 2887 19909 2991 19943
rect 2991 19909 3025 19943
rect 3025 19909 3129 19943
rect 3129 19909 3163 19943
rect 3163 19909 3267 19943
rect 3267 19909 3301 19943
rect 3301 19909 3405 19943
rect 3405 19909 3439 19943
rect 3439 19909 3543 19943
rect 3543 19909 3577 19943
rect 3577 19909 3681 19943
rect 3681 19909 3715 19943
rect 3715 19909 3819 19943
rect 3819 19909 3853 19943
rect 3853 19909 3957 19943
rect 3957 19909 3991 19943
rect 3991 19909 4095 19943
rect 4095 19909 4129 19943
rect 4129 19909 4233 19943
rect 4233 19909 4267 19943
rect 4267 19909 4371 19943
rect 4371 19909 4405 19943
rect 4405 19909 4509 19943
rect 4509 19909 4543 19943
rect 4543 19909 4569 19943
rect 2663 19806 4569 19909
rect 2663 19772 2715 19806
rect 2715 19772 2749 19806
rect 2749 19772 2853 19806
rect 2853 19772 2887 19806
rect 2887 19772 2991 19806
rect 2991 19772 3025 19806
rect 3025 19772 3129 19806
rect 3129 19772 3163 19806
rect 3163 19772 3267 19806
rect 3267 19772 3301 19806
rect 3301 19772 3405 19806
rect 3405 19772 3439 19806
rect 3439 19772 3543 19806
rect 3543 19772 3577 19806
rect 3577 19772 3681 19806
rect 3681 19772 3715 19806
rect 3715 19772 3819 19806
rect 3819 19772 3853 19806
rect 3853 19772 3957 19806
rect 3957 19772 3991 19806
rect 3991 19772 4095 19806
rect 4095 19772 4129 19806
rect 4129 19772 4233 19806
rect 4233 19772 4267 19806
rect 4267 19772 4371 19806
rect 4371 19772 4405 19806
rect 4405 19772 4509 19806
rect 4509 19772 4543 19806
rect 4543 19772 4569 19806
rect 2663 19669 4569 19772
rect 2663 19635 2715 19669
rect 2715 19635 2749 19669
rect 2749 19635 2853 19669
rect 2853 19635 2887 19669
rect 2887 19635 2991 19669
rect 2991 19635 3025 19669
rect 3025 19635 3129 19669
rect 3129 19635 3163 19669
rect 3163 19635 3267 19669
rect 3267 19635 3301 19669
rect 3301 19635 3405 19669
rect 3405 19635 3439 19669
rect 3439 19635 3543 19669
rect 3543 19635 3577 19669
rect 3577 19635 3681 19669
rect 3681 19635 3715 19669
rect 3715 19635 3819 19669
rect 3819 19635 3853 19669
rect 3853 19635 3957 19669
rect 3957 19635 3991 19669
rect 3991 19635 4095 19669
rect 4095 19635 4129 19669
rect 4129 19635 4233 19669
rect 4233 19635 4267 19669
rect 4267 19635 4371 19669
rect 4371 19635 4405 19669
rect 4405 19635 4509 19669
rect 4509 19635 4543 19669
rect 4543 19635 4569 19669
rect 2663 19532 4569 19635
rect 2663 19498 2715 19532
rect 2715 19498 2749 19532
rect 2749 19498 2853 19532
rect 2853 19498 2887 19532
rect 2887 19498 2991 19532
rect 2991 19498 3025 19532
rect 3025 19498 3129 19532
rect 3129 19498 3163 19532
rect 3163 19498 3267 19532
rect 3267 19498 3301 19532
rect 3301 19498 3405 19532
rect 3405 19498 3439 19532
rect 3439 19498 3543 19532
rect 3543 19498 3577 19532
rect 3577 19498 3681 19532
rect 3681 19498 3715 19532
rect 3715 19498 3819 19532
rect 3819 19498 3853 19532
rect 3853 19498 3957 19532
rect 3957 19498 3991 19532
rect 3991 19498 4095 19532
rect 4095 19498 4129 19532
rect 4129 19498 4233 19532
rect 4233 19498 4267 19532
rect 4267 19498 4371 19532
rect 4371 19498 4405 19532
rect 4405 19498 4509 19532
rect 4509 19498 4543 19532
rect 4543 19498 4569 19532
rect 2663 19395 4569 19498
rect 2663 19361 2715 19395
rect 2715 19361 2749 19395
rect 2749 19361 2853 19395
rect 2853 19361 2887 19395
rect 2887 19361 2991 19395
rect 2991 19361 3025 19395
rect 3025 19361 3129 19395
rect 3129 19361 3163 19395
rect 3163 19361 3267 19395
rect 3267 19361 3301 19395
rect 3301 19361 3405 19395
rect 3405 19361 3439 19395
rect 3439 19361 3543 19395
rect 3543 19361 3577 19395
rect 3577 19361 3681 19395
rect 3681 19361 3715 19395
rect 3715 19361 3819 19395
rect 3819 19361 3853 19395
rect 3853 19361 3957 19395
rect 3957 19361 3991 19395
rect 3991 19361 4095 19395
rect 4095 19361 4129 19395
rect 4129 19361 4233 19395
rect 4233 19361 4267 19395
rect 4267 19361 4371 19395
rect 4371 19361 4405 19395
rect 4405 19361 4509 19395
rect 4509 19361 4543 19395
rect 4543 19361 4569 19395
rect 5046 20680 5080 20714
rect 5118 20680 5152 20714
rect 5046 20607 5080 20641
rect 5118 20607 5152 20641
rect 5046 20534 5080 20568
rect 5118 20534 5152 20568
rect 5046 20461 5080 20495
rect 5118 20461 5152 20495
rect 5046 19380 5152 20422
rect 5323 20680 5357 20714
rect 5395 20680 5429 20714
rect 5323 20607 5357 20641
rect 5395 20607 5429 20641
rect 5323 20534 5357 20568
rect 5395 20534 5429 20568
rect 5323 20461 5357 20495
rect 5395 20461 5429 20495
rect 5323 19380 5429 20422
rect 5600 20680 5634 20714
rect 5672 20680 5706 20714
rect 5600 20607 5634 20641
rect 5672 20607 5706 20641
rect 5600 20534 5634 20568
rect 5672 20534 5706 20568
rect 5600 20461 5634 20495
rect 5672 20461 5706 20495
rect 5600 19380 5706 20422
rect 5877 20680 5911 20714
rect 5949 20680 5983 20714
rect 5877 20607 5911 20641
rect 5949 20607 5983 20641
rect 5877 20534 5911 20568
rect 5949 20534 5983 20568
rect 5877 20461 5911 20495
rect 5949 20461 5983 20495
rect 5877 19380 5983 20422
rect 6154 20680 6188 20714
rect 6226 20680 6260 20714
rect 6154 20607 6188 20641
rect 6226 20607 6260 20641
rect 6154 20534 6188 20568
rect 6226 20534 6260 20568
rect 6154 20461 6188 20495
rect 6226 20461 6260 20495
rect 6154 19380 6260 20422
rect 6431 20680 6465 20714
rect 6503 20680 6537 20714
rect 6431 20607 6465 20641
rect 6503 20607 6537 20641
rect 6431 20534 6465 20568
rect 6503 20534 6537 20568
rect 6431 20461 6465 20495
rect 6503 20461 6537 20495
rect 6431 19380 6537 20422
rect 6708 20680 6742 20714
rect 6780 20680 6814 20714
rect 6708 20607 6742 20641
rect 6780 20607 6814 20641
rect 6708 20534 6742 20568
rect 6780 20534 6814 20568
rect 6708 20461 6742 20495
rect 6780 20461 6814 20495
rect 6708 19380 6814 20422
rect 6985 20680 7019 20714
rect 7057 20680 7091 20714
rect 6985 20607 7019 20641
rect 7057 20607 7091 20641
rect 6985 20534 7019 20568
rect 7057 20534 7091 20568
rect 6985 20461 7019 20495
rect 7057 20461 7091 20495
rect 6985 19380 7091 20422
rect 7262 20680 7296 20714
rect 7334 20680 7368 20714
rect 7262 20607 7296 20641
rect 7334 20607 7368 20641
rect 7262 20534 7296 20568
rect 7334 20534 7368 20568
rect 7262 20461 7296 20495
rect 7334 20461 7368 20495
rect 7262 19380 7368 20422
rect 7539 20680 7573 20714
rect 7611 20680 7645 20714
rect 7539 20607 7573 20641
rect 7611 20607 7645 20641
rect 7539 20534 7573 20568
rect 7611 20534 7645 20568
rect 7539 20461 7573 20495
rect 7611 20461 7645 20495
rect 7539 19380 7645 20422
rect 7816 20680 7850 20714
rect 7888 20680 7922 20714
rect 7816 20607 7850 20641
rect 7888 20607 7922 20641
rect 7816 20534 7850 20568
rect 7888 20534 7922 20568
rect 7816 20461 7850 20495
rect 7888 20461 7922 20495
rect 7816 19380 7922 20422
rect 8050 20685 8084 20719
rect 8184 20675 8218 20709
rect 8050 20613 8084 20647
rect 8184 20603 8218 20637
rect 8050 20541 8084 20575
rect 8184 20531 8218 20565
rect 8050 20469 8084 20503
rect 8184 20459 8218 20493
rect 8050 20397 8084 20431
rect 8184 20387 8218 20421
rect 8050 20325 8084 20359
rect 8184 20315 8218 20349
rect 8050 20253 8084 20287
rect 8184 20243 8218 20277
rect 8050 20181 8084 20215
rect 8184 20171 8218 20205
rect 8050 20109 8084 20143
rect 8184 20099 8218 20133
rect 8050 20037 8084 20071
rect 8184 20027 8218 20061
rect 8050 19965 8084 19999
rect 8184 19955 8218 19989
rect 8050 19893 8084 19927
rect 8184 19883 8218 19917
rect 8050 19821 8084 19855
rect 8184 19811 8218 19845
rect 8050 19749 8084 19783
rect 8184 19739 8218 19773
rect 8050 19677 8084 19711
rect 8184 19667 8218 19701
rect 8050 19605 8084 19639
rect 8184 19595 8218 19629
rect 8050 19533 8084 19567
rect 8184 19523 8218 19557
rect 8050 19461 8084 19495
rect 8184 19451 8218 19485
rect 8050 19389 8084 19423
rect 8184 19379 8218 19413
rect 2663 19258 4569 19361
rect 2663 19224 2715 19258
rect 2715 19224 2749 19258
rect 2749 19224 2853 19258
rect 2853 19224 2887 19258
rect 2887 19224 2991 19258
rect 2991 19224 3025 19258
rect 3025 19224 3129 19258
rect 3129 19224 3163 19258
rect 3163 19224 3267 19258
rect 3267 19224 3301 19258
rect 3301 19224 3405 19258
rect 3405 19224 3439 19258
rect 3439 19224 3543 19258
rect 3543 19224 3577 19258
rect 3577 19224 3681 19258
rect 3681 19224 3715 19258
rect 3715 19224 3819 19258
rect 3819 19224 3853 19258
rect 3853 19224 3957 19258
rect 3957 19224 3991 19258
rect 3991 19224 4095 19258
rect 4095 19224 4129 19258
rect 4129 19224 4233 19258
rect 4233 19224 4267 19258
rect 4267 19224 4371 19258
rect 4371 19224 4405 19258
rect 4405 19224 4509 19258
rect 4509 19224 4543 19258
rect 4543 19224 4569 19258
rect 2663 19121 4569 19224
rect 2663 19087 2715 19121
rect 2715 19087 2749 19121
rect 2749 19087 2853 19121
rect 2853 19087 2887 19121
rect 2887 19087 2991 19121
rect 2991 19087 3025 19121
rect 3025 19087 3129 19121
rect 3129 19087 3163 19121
rect 3163 19087 3267 19121
rect 3267 19087 3301 19121
rect 3301 19087 3405 19121
rect 3405 19087 3439 19121
rect 3439 19087 3543 19121
rect 3543 19087 3577 19121
rect 3577 19087 3681 19121
rect 3681 19087 3715 19121
rect 3715 19087 3819 19121
rect 3819 19087 3853 19121
rect 3853 19087 3957 19121
rect 3957 19087 3991 19121
rect 3991 19087 4095 19121
rect 4095 19087 4129 19121
rect 4129 19087 4233 19121
rect 4233 19087 4267 19121
rect 4267 19087 4371 19121
rect 4371 19087 4405 19121
rect 4405 19087 4509 19121
rect 4509 19087 4543 19121
rect 4543 19087 4569 19121
rect 8050 19317 8084 19351
rect 8184 19307 8218 19341
rect 8050 19245 8084 19279
rect 8184 19235 8218 19269
rect 8050 19173 8084 19207
rect 8184 19163 8218 19197
rect 2663 18984 4569 19087
rect 5251 19085 5255 19119
rect 5255 19085 5285 19119
rect 5325 19085 5359 19119
rect 5399 19085 5429 19119
rect 5429 19085 5433 19119
rect 5473 19085 5499 19119
rect 5499 19085 5507 19119
rect 5547 19085 5569 19119
rect 5569 19085 5581 19119
rect 5621 19085 5639 19119
rect 5639 19085 5655 19119
rect 5695 19085 5709 19119
rect 5709 19085 5729 19119
rect 5769 19085 5779 19119
rect 5779 19085 5803 19119
rect 5843 19085 5849 19119
rect 5849 19085 5877 19119
rect 5917 19085 5919 19119
rect 5919 19085 5951 19119
rect 5991 19085 6023 19119
rect 6023 19085 6025 19119
rect 6065 19085 6092 19119
rect 6092 19085 6099 19119
rect 6139 19085 6161 19119
rect 6161 19085 6173 19119
rect 6213 19085 6230 19119
rect 6230 19085 6247 19119
rect 6287 19085 6299 19119
rect 6299 19085 6321 19119
rect 6361 19085 6368 19119
rect 6368 19085 6395 19119
rect 6435 19085 6437 19119
rect 6437 19085 6469 19119
rect 6509 19085 6540 19119
rect 6540 19085 6543 19119
rect 6583 19085 6609 19119
rect 6609 19085 6617 19119
rect 6657 19085 6678 19119
rect 6678 19085 6691 19119
rect 6731 19085 6747 19119
rect 6747 19085 6765 19119
rect 6805 19085 6816 19119
rect 6816 19085 6839 19119
rect 6879 19085 6885 19119
rect 6885 19085 6913 19119
rect 6953 19085 6954 19119
rect 6954 19085 6987 19119
rect 7026 19085 7058 19119
rect 7058 19085 7060 19119
rect 7099 19085 7127 19119
rect 7127 19085 7133 19119
rect 7172 19085 7196 19119
rect 7196 19085 7206 19119
rect 7245 19085 7265 19119
rect 7265 19085 7279 19119
rect 7318 19085 7334 19119
rect 7334 19085 7352 19119
rect 7391 19085 7403 19119
rect 7403 19085 7425 19119
rect 7464 19085 7472 19119
rect 7472 19085 7498 19119
rect 7537 19085 7541 19119
rect 7541 19085 7571 19119
rect 7610 19085 7644 19119
rect 7683 19085 7713 19119
rect 7713 19085 7717 19119
rect 8050 19101 8084 19135
rect 8184 19091 8218 19125
rect 2663 18950 2715 18984
rect 2715 18950 2749 18984
rect 2749 18950 2853 18984
rect 2853 18950 2887 18984
rect 2887 18950 2991 18984
rect 2991 18950 3025 18984
rect 3025 18950 3129 18984
rect 3129 18950 3163 18984
rect 3163 18950 3267 18984
rect 3267 18950 3301 18984
rect 3301 18950 3405 18984
rect 3405 18950 3439 18984
rect 3439 18950 3543 18984
rect 3543 18950 3577 18984
rect 3577 18950 3681 18984
rect 3681 18950 3715 18984
rect 3715 18950 3819 18984
rect 3819 18950 3853 18984
rect 3853 18950 3957 18984
rect 3957 18950 3991 18984
rect 3991 18950 4095 18984
rect 4095 18950 4129 18984
rect 4129 18950 4233 18984
rect 4233 18950 4267 18984
rect 4267 18950 4371 18984
rect 4371 18950 4405 18984
rect 4405 18950 4509 18984
rect 4509 18950 4543 18984
rect 4543 18950 4569 18984
rect 2663 18847 4569 18950
rect 2663 18813 2715 18847
rect 2715 18813 2749 18847
rect 2749 18813 2853 18847
rect 2853 18813 2887 18847
rect 2887 18813 2991 18847
rect 2991 18813 3025 18847
rect 3025 18813 3129 18847
rect 3129 18813 3163 18847
rect 3163 18813 3267 18847
rect 3267 18813 3301 18847
rect 3301 18813 3405 18847
rect 3405 18813 3439 18847
rect 3439 18813 3543 18847
rect 3543 18813 3577 18847
rect 3577 18813 3681 18847
rect 3681 18813 3715 18847
rect 3715 18813 3819 18847
rect 3819 18813 3853 18847
rect 3853 18813 3957 18847
rect 3957 18813 3991 18847
rect 3991 18813 4095 18847
rect 4095 18813 4129 18847
rect 4129 18813 4233 18847
rect 4233 18813 4267 18847
rect 4267 18813 4371 18847
rect 4371 18813 4405 18847
rect 4405 18813 4509 18847
rect 4509 18813 4543 18847
rect 4543 18813 4569 18847
rect 2663 18710 4569 18813
rect 8050 19029 8084 19063
rect 8184 19019 8218 19053
rect 8050 18957 8084 18991
rect 8184 18947 8218 18981
rect 8050 18885 8084 18919
rect 8184 18875 8218 18909
rect 8050 18813 8084 18847
rect 8184 18803 8218 18837
rect 8050 18741 8084 18775
rect 8184 18731 8218 18765
rect 2663 18676 2715 18710
rect 2715 18676 2749 18710
rect 2749 18676 2853 18710
rect 2853 18676 2887 18710
rect 2887 18676 2991 18710
rect 2991 18676 3025 18710
rect 3025 18676 3129 18710
rect 3129 18676 3163 18710
rect 3163 18676 3267 18710
rect 3267 18676 3301 18710
rect 3301 18676 3405 18710
rect 3405 18676 3439 18710
rect 3439 18676 3543 18710
rect 3543 18676 3577 18710
rect 3577 18676 3681 18710
rect 3681 18676 3715 18710
rect 3715 18676 3819 18710
rect 3819 18676 3853 18710
rect 3853 18676 3957 18710
rect 3957 18676 3991 18710
rect 3991 18676 4095 18710
rect 4095 18676 4129 18710
rect 4129 18676 4233 18710
rect 4233 18676 4267 18710
rect 4267 18676 4371 18710
rect 4371 18676 4405 18710
rect 4405 18676 4509 18710
rect 4509 18676 4543 18710
rect 4543 18676 4569 18710
rect 2663 18573 4569 18676
rect 2663 18563 2715 18573
rect 2715 18563 2749 18573
rect 2749 18563 2853 18573
rect 2853 18563 2887 18573
rect 2887 18563 2991 18573
rect 2991 18563 3025 18573
rect 3025 18563 3129 18573
rect 3129 18563 3163 18573
rect 3163 18563 3267 18573
rect 3267 18563 3301 18573
rect 3301 18563 3405 18573
rect 3405 18563 3439 18573
rect 3439 18563 3543 18573
rect 3543 18563 3577 18573
rect 3577 18563 3681 18573
rect 3681 18563 3715 18573
rect 3715 18563 3819 18573
rect 3819 18563 3853 18573
rect 3853 18563 3957 18573
rect 3957 18563 3991 18573
rect 3991 18563 4095 18573
rect 4095 18563 4129 18573
rect 4129 18563 4233 18573
rect 4233 18563 4267 18573
rect 4267 18563 4371 18573
rect 4371 18563 4405 18573
rect 4405 18563 4509 18573
rect 4509 18563 4543 18573
rect 4543 18563 4569 18573
rect 2663 18490 2697 18524
rect 2735 18490 2769 18524
rect 2807 18490 2841 18524
rect 2879 18490 2913 18524
rect 2951 18490 2985 18524
rect 3023 18490 3057 18524
rect 3095 18490 3129 18524
rect 3167 18490 3201 18524
rect 3239 18490 3273 18524
rect 3311 18490 3345 18524
rect 3383 18490 3417 18524
rect 3455 18490 3489 18524
rect 3527 18490 3561 18524
rect 3599 18490 3633 18524
rect 3671 18490 3705 18524
rect 3743 18490 3777 18524
rect 3815 18490 3849 18524
rect 3887 18490 3921 18524
rect 3959 18490 3993 18524
rect 4031 18490 4065 18524
rect 4103 18490 4137 18524
rect 4175 18490 4209 18524
rect 4247 18490 4281 18524
rect 4319 18490 4353 18524
rect 4391 18490 4425 18524
rect 4463 18490 4497 18524
rect 4535 18490 4569 18524
rect 2663 18417 2697 18451
rect 2735 18436 2769 18451
rect 2735 18417 2749 18436
rect 2749 18417 2769 18436
rect 2807 18417 2841 18451
rect 2879 18436 2913 18451
rect 2879 18417 2887 18436
rect 2887 18417 2913 18436
rect 2951 18417 2985 18451
rect 3023 18436 3057 18451
rect 3023 18417 3025 18436
rect 3025 18417 3057 18436
rect 3095 18417 3129 18451
rect 3167 18417 3201 18451
rect 3239 18436 3273 18451
rect 3239 18417 3267 18436
rect 3267 18417 3273 18436
rect 3311 18417 3345 18451
rect 3383 18436 3417 18451
rect 3383 18417 3405 18436
rect 3405 18417 3417 18436
rect 3455 18417 3489 18451
rect 3527 18436 3561 18451
rect 3527 18417 3543 18436
rect 3543 18417 3561 18436
rect 3599 18417 3633 18451
rect 3671 18436 3705 18451
rect 3671 18417 3681 18436
rect 3681 18417 3705 18436
rect 3743 18417 3777 18451
rect 3815 18436 3849 18451
rect 3815 18417 3819 18436
rect 3819 18417 3849 18436
rect 3887 18417 3921 18451
rect 3959 18436 3993 18451
rect 3959 18417 3991 18436
rect 3991 18417 3993 18436
rect 4031 18417 4065 18451
rect 4103 18436 4137 18451
rect 4103 18417 4129 18436
rect 4129 18417 4137 18436
rect 4175 18417 4209 18451
rect 4247 18436 4281 18451
rect 4247 18417 4267 18436
rect 4267 18417 4281 18436
rect 4319 18417 4353 18451
rect 4391 18436 4425 18451
rect 4391 18417 4405 18436
rect 4405 18417 4425 18436
rect 4463 18417 4497 18451
rect 4535 18436 4569 18451
rect 4535 18417 4543 18436
rect 4543 18417 4569 18436
rect 2663 18344 2697 18378
rect 2735 18344 2769 18378
rect 2807 18344 2841 18378
rect 2879 18344 2913 18378
rect 2951 18344 2985 18378
rect 3023 18344 3057 18378
rect 3095 18344 3129 18378
rect 3167 18344 3201 18378
rect 3239 18344 3273 18378
rect 3311 18344 3345 18378
rect 3383 18344 3417 18378
rect 3455 18344 3489 18378
rect 3527 18344 3561 18378
rect 3599 18344 3633 18378
rect 3671 18344 3705 18378
rect 3743 18344 3777 18378
rect 3815 18344 3849 18378
rect 3887 18344 3921 18378
rect 3959 18344 3993 18378
rect 4031 18344 4065 18378
rect 4103 18344 4137 18378
rect 4175 18344 4209 18378
rect 4247 18344 4281 18378
rect 4319 18344 4353 18378
rect 4391 18344 4425 18378
rect 4463 18344 4497 18378
rect 4535 18344 4569 18378
rect 2663 18271 2697 18305
rect 2735 18299 2769 18305
rect 2735 18271 2749 18299
rect 2749 18271 2769 18299
rect 2807 18271 2841 18305
rect 2879 18299 2913 18305
rect 2879 18271 2887 18299
rect 2887 18271 2913 18299
rect 2951 18271 2985 18305
rect 3023 18299 3057 18305
rect 3023 18271 3025 18299
rect 3025 18271 3057 18299
rect 3095 18271 3129 18305
rect 3167 18271 3201 18305
rect 3239 18299 3273 18305
rect 3239 18271 3267 18299
rect 3267 18271 3273 18299
rect 3311 18271 3345 18305
rect 3383 18299 3417 18305
rect 3383 18271 3405 18299
rect 3405 18271 3417 18299
rect 3455 18271 3489 18305
rect 3527 18299 3561 18305
rect 3527 18271 3543 18299
rect 3543 18271 3561 18299
rect 3599 18271 3633 18305
rect 3671 18299 3705 18305
rect 3671 18271 3681 18299
rect 3681 18271 3705 18299
rect 3743 18271 3777 18305
rect 3815 18299 3849 18305
rect 3815 18271 3819 18299
rect 3819 18271 3849 18299
rect 3887 18271 3921 18305
rect 3959 18299 3993 18305
rect 3959 18271 3991 18299
rect 3991 18271 3993 18299
rect 4031 18271 4065 18305
rect 4103 18299 4137 18305
rect 4103 18271 4129 18299
rect 4129 18271 4137 18299
rect 4175 18271 4209 18305
rect 4247 18299 4281 18305
rect 4247 18271 4267 18299
rect 4267 18271 4281 18299
rect 4319 18271 4353 18305
rect 4391 18299 4425 18305
rect 4391 18271 4405 18299
rect 4405 18271 4425 18299
rect 4463 18271 4497 18305
rect 4535 18299 4569 18305
rect 4535 18271 4543 18299
rect 4543 18271 4569 18299
rect 2663 18198 2697 18232
rect 2735 18198 2769 18232
rect 2807 18198 2841 18232
rect 2879 18198 2913 18232
rect 2951 18198 2985 18232
rect 3023 18198 3057 18232
rect 3095 18198 3129 18232
rect 3167 18198 3201 18232
rect 3239 18198 3273 18232
rect 3311 18198 3345 18232
rect 3383 18198 3417 18232
rect 3455 18198 3489 18232
rect 3527 18198 3561 18232
rect 3599 18198 3633 18232
rect 3671 18198 3705 18232
rect 3743 18198 3777 18232
rect 3815 18198 3849 18232
rect 3887 18198 3921 18232
rect 3959 18198 3993 18232
rect 4031 18198 4065 18232
rect 4103 18198 4137 18232
rect 4175 18198 4209 18232
rect 4247 18198 4281 18232
rect 4319 18198 4353 18232
rect 4391 18198 4425 18232
rect 4463 18198 4497 18232
rect 4535 18198 4569 18232
rect 2663 18125 2697 18159
rect 2735 18128 2749 18159
rect 2749 18128 2769 18159
rect 2735 18125 2769 18128
rect 2807 18125 2841 18159
rect 2879 18128 2887 18159
rect 2887 18128 2913 18159
rect 2879 18125 2913 18128
rect 2951 18125 2985 18159
rect 3023 18128 3025 18159
rect 3025 18128 3057 18159
rect 3023 18125 3057 18128
rect 3095 18125 3129 18159
rect 3167 18125 3201 18159
rect 3239 18128 3267 18159
rect 3267 18128 3273 18159
rect 3239 18125 3273 18128
rect 3311 18125 3345 18159
rect 3383 18128 3405 18159
rect 3405 18128 3417 18159
rect 3383 18125 3417 18128
rect 3455 18125 3489 18159
rect 3527 18128 3543 18159
rect 3543 18128 3561 18159
rect 3527 18125 3561 18128
rect 3599 18125 3633 18159
rect 3671 18128 3681 18159
rect 3681 18128 3705 18159
rect 3671 18125 3705 18128
rect 3743 18125 3777 18159
rect 3815 18128 3819 18159
rect 3819 18128 3849 18159
rect 3815 18125 3849 18128
rect 3887 18125 3921 18159
rect 3959 18128 3991 18159
rect 3991 18128 3993 18159
rect 3959 18125 3993 18128
rect 4031 18125 4065 18159
rect 4103 18128 4129 18159
rect 4129 18128 4137 18159
rect 4103 18125 4137 18128
rect 4175 18125 4209 18159
rect 4247 18128 4267 18159
rect 4267 18128 4281 18159
rect 4247 18125 4281 18128
rect 4319 18125 4353 18159
rect 4391 18128 4405 18159
rect 4405 18128 4425 18159
rect 4391 18125 4425 18128
rect 4463 18125 4497 18159
rect 4535 18128 4543 18159
rect 4543 18128 4569 18159
rect 4535 18125 4569 18128
rect 2663 18052 2697 18086
rect 2735 18052 2769 18086
rect 2807 18052 2841 18086
rect 2879 18052 2913 18086
rect 2951 18052 2985 18086
rect 3023 18052 3057 18086
rect 3095 18052 3129 18086
rect 3167 18052 3201 18086
rect 3239 18052 3273 18086
rect 3311 18052 3345 18086
rect 3383 18052 3417 18086
rect 3455 18052 3489 18086
rect 3527 18052 3561 18086
rect 3599 18052 3633 18086
rect 3671 18052 3705 18086
rect 3743 18052 3777 18086
rect 3815 18052 3849 18086
rect 3887 18052 3921 18086
rect 3959 18052 3993 18086
rect 4031 18052 4065 18086
rect 4103 18052 4137 18086
rect 4175 18052 4209 18086
rect 4247 18052 4281 18086
rect 4319 18052 4353 18086
rect 4391 18052 4425 18086
rect 4463 18052 4497 18086
rect 4535 18052 4569 18086
rect 2663 17979 2697 18013
rect 2735 17991 2749 18013
rect 2749 17991 2769 18013
rect 2735 17979 2769 17991
rect 2807 17979 2841 18013
rect 2879 17991 2887 18013
rect 2887 17991 2913 18013
rect 2879 17979 2913 17991
rect 2951 17979 2985 18013
rect 3023 17991 3025 18013
rect 3025 17991 3057 18013
rect 3023 17979 3057 17991
rect 3095 17979 3129 18013
rect 3167 17979 3201 18013
rect 3239 17991 3267 18013
rect 3267 17991 3273 18013
rect 3239 17979 3273 17991
rect 3311 17979 3345 18013
rect 3383 17991 3405 18013
rect 3405 17991 3417 18013
rect 3383 17979 3417 17991
rect 3455 17979 3489 18013
rect 3527 17991 3543 18013
rect 3543 17991 3561 18013
rect 3527 17979 3561 17991
rect 3599 17979 3633 18013
rect 3671 17991 3681 18013
rect 3681 17991 3705 18013
rect 3671 17979 3705 17991
rect 3743 17979 3777 18013
rect 3815 17991 3819 18013
rect 3819 17991 3849 18013
rect 3815 17979 3849 17991
rect 3887 17979 3921 18013
rect 3959 17991 3991 18013
rect 3991 17991 3993 18013
rect 3959 17979 3993 17991
rect 4031 17979 4065 18013
rect 4103 17991 4129 18013
rect 4129 17991 4137 18013
rect 4103 17979 4137 17991
rect 4175 17979 4209 18013
rect 4247 17991 4267 18013
rect 4267 17991 4281 18013
rect 4247 17979 4281 17991
rect 4319 17979 4353 18013
rect 4391 17991 4405 18013
rect 4405 17991 4425 18013
rect 4391 17979 4425 17991
rect 4463 17979 4497 18013
rect 4535 17991 4543 18013
rect 4543 17991 4569 18013
rect 4535 17979 4569 17991
rect 2663 17906 2697 17940
rect 2735 17906 2769 17940
rect 2807 17906 2841 17940
rect 2879 17906 2913 17940
rect 2951 17906 2985 17940
rect 3023 17906 3057 17940
rect 3095 17906 3129 17940
rect 3167 17906 3201 17940
rect 3239 17906 3273 17940
rect 3311 17906 3345 17940
rect 3383 17906 3417 17940
rect 3455 17906 3489 17940
rect 3527 17906 3561 17940
rect 3599 17906 3633 17940
rect 3671 17906 3705 17940
rect 3743 17906 3777 17940
rect 3815 17906 3849 17940
rect 3887 17906 3921 17940
rect 3959 17906 3993 17940
rect 4031 17906 4065 17940
rect 4103 17906 4137 17940
rect 4175 17906 4209 17940
rect 4247 17906 4281 17940
rect 4319 17906 4353 17940
rect 4391 17906 4425 17940
rect 4463 17906 4497 17940
rect 4535 17906 4569 17940
rect 2663 17833 2697 17867
rect 2735 17854 2749 17867
rect 2749 17854 2769 17867
rect 2735 17833 2769 17854
rect 2807 17833 2841 17867
rect 2879 17854 2887 17867
rect 2887 17854 2913 17867
rect 2879 17833 2913 17854
rect 2951 17833 2985 17867
rect 3023 17854 3025 17867
rect 3025 17854 3057 17867
rect 3023 17833 3057 17854
rect 3095 17833 3129 17867
rect 3167 17833 3201 17867
rect 3239 17854 3267 17867
rect 3267 17854 3273 17867
rect 3239 17833 3273 17854
rect 3311 17833 3345 17867
rect 3383 17854 3405 17867
rect 3405 17854 3417 17867
rect 3383 17833 3417 17854
rect 3455 17833 3489 17867
rect 3527 17854 3543 17867
rect 3543 17854 3561 17867
rect 3527 17833 3561 17854
rect 3599 17833 3633 17867
rect 3671 17854 3681 17867
rect 3681 17854 3705 17867
rect 3671 17833 3705 17854
rect 3743 17833 3777 17867
rect 3815 17854 3819 17867
rect 3819 17854 3849 17867
rect 3815 17833 3849 17854
rect 3887 17833 3921 17867
rect 3959 17854 3991 17867
rect 3991 17854 3993 17867
rect 3959 17833 3993 17854
rect 4031 17833 4065 17867
rect 4103 17854 4129 17867
rect 4129 17854 4137 17867
rect 4103 17833 4137 17854
rect 4175 17833 4209 17867
rect 4247 17854 4267 17867
rect 4267 17854 4281 17867
rect 4247 17833 4281 17854
rect 4319 17833 4353 17867
rect 4391 17854 4405 17867
rect 4405 17854 4425 17867
rect 4391 17833 4425 17854
rect 4463 17833 4497 17867
rect 4535 17854 4543 17867
rect 4543 17854 4569 17867
rect 4535 17833 4569 17854
rect 2663 17760 2697 17794
rect 2735 17760 2769 17794
rect 2807 17760 2841 17794
rect 2879 17760 2913 17794
rect 2951 17760 2985 17794
rect 3023 17760 3057 17794
rect 3095 17760 3129 17794
rect 3167 17760 3201 17794
rect 3239 17760 3273 17794
rect 3311 17760 3345 17794
rect 3383 17760 3417 17794
rect 3455 17760 3489 17794
rect 3527 17760 3561 17794
rect 3599 17760 3633 17794
rect 3671 17760 3705 17794
rect 3743 17760 3777 17794
rect 3815 17760 3849 17794
rect 3887 17760 3921 17794
rect 3959 17760 3993 17794
rect 4031 17760 4065 17794
rect 4103 17760 4137 17794
rect 4175 17760 4209 17794
rect 4247 17760 4281 17794
rect 4319 17760 4353 17794
rect 4391 17760 4425 17794
rect 4463 17760 4497 17794
rect 4535 17760 4569 17794
rect 2663 17687 2697 17721
rect 2735 17717 2749 17721
rect 2749 17717 2769 17721
rect 2735 17687 2769 17717
rect 2807 17687 2841 17721
rect 2879 17717 2887 17721
rect 2887 17717 2913 17721
rect 2879 17687 2913 17717
rect 2951 17687 2985 17721
rect 3023 17717 3025 17721
rect 3025 17717 3057 17721
rect 3023 17687 3057 17717
rect 3095 17687 3129 17721
rect 3167 17687 3201 17721
rect 3239 17717 3267 17721
rect 3267 17717 3273 17721
rect 3239 17687 3273 17717
rect 3311 17687 3345 17721
rect 3383 17717 3405 17721
rect 3405 17717 3417 17721
rect 3383 17687 3417 17717
rect 3455 17687 3489 17721
rect 3527 17717 3543 17721
rect 3543 17717 3561 17721
rect 3527 17687 3561 17717
rect 3599 17687 3633 17721
rect 3671 17717 3681 17721
rect 3681 17717 3705 17721
rect 3671 17687 3705 17717
rect 3743 17687 3777 17721
rect 3815 17717 3819 17721
rect 3819 17717 3849 17721
rect 3815 17687 3849 17717
rect 3887 17687 3921 17721
rect 3959 17717 3991 17721
rect 3991 17717 3993 17721
rect 3959 17687 3993 17717
rect 4031 17687 4065 17721
rect 4103 17717 4129 17721
rect 4129 17717 4137 17721
rect 4103 17687 4137 17717
rect 4175 17687 4209 17721
rect 4247 17717 4267 17721
rect 4267 17717 4281 17721
rect 4247 17687 4281 17717
rect 4319 17687 4353 17721
rect 4391 17717 4405 17721
rect 4405 17717 4425 17721
rect 4391 17687 4425 17717
rect 4463 17687 4497 17721
rect 4535 17717 4543 17721
rect 4543 17717 4569 17721
rect 4535 17687 4569 17717
rect 2663 17614 2697 17648
rect 2735 17614 2769 17648
rect 2807 17614 2841 17648
rect 2879 17614 2913 17648
rect 2951 17614 2985 17648
rect 3023 17614 3057 17648
rect 3095 17614 3129 17648
rect 3167 17614 3201 17648
rect 3239 17614 3273 17648
rect 3311 17614 3345 17648
rect 3383 17614 3417 17648
rect 3455 17614 3489 17648
rect 3527 17614 3561 17648
rect 3599 17614 3633 17648
rect 3671 17614 3705 17648
rect 3743 17614 3777 17648
rect 3815 17614 3849 17648
rect 3887 17614 3921 17648
rect 3959 17614 3993 17648
rect 4031 17614 4065 17648
rect 4103 17614 4137 17648
rect 4175 17614 4209 17648
rect 4247 17614 4281 17648
rect 4319 17614 4353 17648
rect 4391 17614 4425 17648
rect 4463 17614 4497 17648
rect 4535 17614 4569 17648
rect 2663 17541 2697 17575
rect 2735 17541 2769 17575
rect 2807 17541 2841 17575
rect 2879 17541 2913 17575
rect 2951 17541 2985 17575
rect 3023 17541 3057 17575
rect 3095 17541 3129 17575
rect 3167 17541 3201 17575
rect 3239 17541 3273 17575
rect 3311 17541 3345 17575
rect 3383 17541 3417 17575
rect 3455 17541 3489 17575
rect 3527 17541 3561 17575
rect 3599 17541 3633 17575
rect 3671 17541 3705 17575
rect 3743 17541 3777 17575
rect 3815 17541 3849 17575
rect 3887 17541 3921 17575
rect 3959 17541 3993 17575
rect 4031 17541 4065 17575
rect 4103 17541 4137 17575
rect 4175 17541 4209 17575
rect 4247 17541 4281 17575
rect 4319 17541 4353 17575
rect 4391 17541 4425 17575
rect 4463 17541 4497 17575
rect 4535 17541 4569 17575
rect 2663 17468 2697 17502
rect 2735 17477 2769 17502
rect 2735 17468 2749 17477
rect 2749 17468 2769 17477
rect 2807 17468 2841 17502
rect 2879 17477 2913 17502
rect 2879 17468 2887 17477
rect 2887 17468 2913 17477
rect 2951 17468 2985 17502
rect 3023 17477 3057 17502
rect 3023 17468 3025 17477
rect 3025 17468 3057 17477
rect 3095 17468 3129 17502
rect 3167 17468 3201 17502
rect 3239 17477 3273 17502
rect 3239 17468 3267 17477
rect 3267 17468 3273 17477
rect 3311 17468 3345 17502
rect 3383 17477 3417 17502
rect 3383 17468 3405 17477
rect 3405 17468 3417 17477
rect 3455 17468 3489 17502
rect 3527 17477 3561 17502
rect 3527 17468 3543 17477
rect 3543 17468 3561 17477
rect 3599 17468 3633 17502
rect 3671 17477 3705 17502
rect 3671 17468 3681 17477
rect 3681 17468 3705 17477
rect 3743 17468 3777 17502
rect 3815 17477 3849 17502
rect 3815 17468 3819 17477
rect 3819 17468 3849 17477
rect 3887 17468 3921 17502
rect 3959 17477 3993 17502
rect 3959 17468 3991 17477
rect 3991 17468 3993 17477
rect 4031 17468 4065 17502
rect 4103 17477 4137 17502
rect 4103 17468 4129 17477
rect 4129 17468 4137 17477
rect 4175 17468 4209 17502
rect 4247 17477 4281 17502
rect 4247 17468 4267 17477
rect 4267 17468 4281 17477
rect 4319 17468 4353 17502
rect 4391 17477 4425 17502
rect 4391 17468 4405 17477
rect 4405 17468 4425 17477
rect 4463 17468 4497 17502
rect 4535 17477 4569 17502
rect 4535 17468 4543 17477
rect 4543 17468 4569 17477
rect 2663 17395 2697 17429
rect 2735 17395 2769 17429
rect 2807 17395 2841 17429
rect 2879 17395 2913 17429
rect 2951 17395 2985 17429
rect 3023 17395 3057 17429
rect 3095 17395 3129 17429
rect 3167 17395 3201 17429
rect 3239 17395 3273 17429
rect 3311 17395 3345 17429
rect 3383 17395 3417 17429
rect 3455 17395 3489 17429
rect 3527 17395 3561 17429
rect 3599 17395 3633 17429
rect 3671 17395 3705 17429
rect 3743 17395 3777 17429
rect 3815 17395 3849 17429
rect 3887 17395 3921 17429
rect 3959 17395 3993 17429
rect 4031 17395 4065 17429
rect 4103 17395 4137 17429
rect 4175 17395 4209 17429
rect 4247 17395 4281 17429
rect 4319 17395 4353 17429
rect 4391 17395 4425 17429
rect 4463 17395 4497 17429
rect 4535 17395 4569 17429
rect 5046 18680 5080 18714
rect 5118 18680 5152 18714
rect 5046 18607 5080 18641
rect 5118 18607 5152 18641
rect 5046 18534 5080 18568
rect 5118 18534 5152 18568
rect 5046 18461 5080 18495
rect 5118 18461 5152 18495
rect 5046 17380 5152 18422
rect 5323 18680 5357 18714
rect 5395 18680 5429 18714
rect 5323 18607 5357 18641
rect 5395 18607 5429 18641
rect 5323 18534 5357 18568
rect 5395 18534 5429 18568
rect 5323 18461 5357 18495
rect 5395 18461 5429 18495
rect 5323 17380 5429 18422
rect 5600 18680 5634 18714
rect 5672 18680 5706 18714
rect 5600 18607 5634 18641
rect 5672 18607 5706 18641
rect 5600 18534 5634 18568
rect 5672 18534 5706 18568
rect 5600 18461 5634 18495
rect 5672 18461 5706 18495
rect 5600 17380 5706 18422
rect 5877 18680 5911 18714
rect 5949 18680 5983 18714
rect 5877 18607 5911 18641
rect 5949 18607 5983 18641
rect 5877 18534 5911 18568
rect 5949 18534 5983 18568
rect 5877 18461 5911 18495
rect 5949 18461 5983 18495
rect 5877 17380 5983 18422
rect 6154 18680 6188 18714
rect 6226 18680 6260 18714
rect 6154 18607 6188 18641
rect 6226 18607 6260 18641
rect 6154 18534 6188 18568
rect 6226 18534 6260 18568
rect 6154 18461 6188 18495
rect 6226 18461 6260 18495
rect 6154 17380 6260 18422
rect 6431 18680 6465 18714
rect 6503 18680 6537 18714
rect 6431 18607 6465 18641
rect 6503 18607 6537 18641
rect 6431 18534 6465 18568
rect 6503 18534 6537 18568
rect 6431 18461 6465 18495
rect 6503 18461 6537 18495
rect 6431 17380 6537 18422
rect 6708 18680 6742 18714
rect 6780 18680 6814 18714
rect 6708 18607 6742 18641
rect 6780 18607 6814 18641
rect 6708 18534 6742 18568
rect 6780 18534 6814 18568
rect 6708 18461 6742 18495
rect 6780 18461 6814 18495
rect 6708 17380 6814 18422
rect 6985 18680 7019 18714
rect 7057 18680 7091 18714
rect 6985 18607 7019 18641
rect 7057 18607 7091 18641
rect 6985 18534 7019 18568
rect 7057 18534 7091 18568
rect 6985 18461 7019 18495
rect 7057 18461 7091 18495
rect 6985 17380 7091 18422
rect 7262 18680 7296 18714
rect 7334 18680 7368 18714
rect 7262 18607 7296 18641
rect 7334 18607 7368 18641
rect 7262 18534 7296 18568
rect 7334 18534 7368 18568
rect 7262 18461 7296 18495
rect 7334 18461 7368 18495
rect 7262 17380 7368 18422
rect 7539 18680 7573 18714
rect 7611 18680 7645 18714
rect 7539 18607 7573 18641
rect 7611 18607 7645 18641
rect 7539 18534 7573 18568
rect 7611 18534 7645 18568
rect 7539 18461 7573 18495
rect 7611 18461 7645 18495
rect 7539 17380 7645 18422
rect 7816 18680 7850 18714
rect 7888 18680 7922 18714
rect 7816 18607 7850 18641
rect 7888 18607 7922 18641
rect 7816 18534 7850 18568
rect 7888 18534 7922 18568
rect 7816 18461 7850 18495
rect 7888 18461 7922 18495
rect 7816 17380 7922 18422
rect 8050 18669 8084 18703
rect 8184 18659 8218 18693
rect 8050 18597 8084 18631
rect 8184 18587 8218 18621
rect 8050 18525 8084 18559
rect 8184 18515 8218 18549
rect 8050 18453 8084 18487
rect 8184 18443 8218 18477
rect 8050 18381 8084 18415
rect 8184 18371 8218 18405
rect 8050 18309 8084 18343
rect 8184 18299 8218 18333
rect 8050 18237 8084 18271
rect 8184 18227 8218 18261
rect 8050 18165 8084 18199
rect 8184 18155 8218 18189
rect 8050 18093 8084 18127
rect 8184 18083 8218 18117
rect 8050 18021 8084 18055
rect 8184 18011 8218 18045
rect 8050 17949 8084 17983
rect 8184 17939 8218 17973
rect 8050 17877 8084 17911
rect 8184 17867 8218 17901
rect 8050 17805 8084 17839
rect 8184 17795 8218 17829
rect 8050 17733 8084 17767
rect 8184 17723 8218 17757
rect 8050 17661 8084 17695
rect 8184 17651 8218 17685
rect 8050 17589 8084 17623
rect 8184 17579 8218 17613
rect 8050 17517 8084 17551
rect 8184 17507 8218 17541
rect 8050 17445 8084 17479
rect 8184 17435 8218 17469
rect 8050 17373 8084 17407
rect 2663 17322 2697 17356
rect 2735 17340 2769 17356
rect 2735 17322 2749 17340
rect 2749 17322 2769 17340
rect 2807 17322 2841 17356
rect 2879 17340 2913 17356
rect 2879 17322 2887 17340
rect 2887 17322 2913 17340
rect 2951 17322 2985 17356
rect 3023 17340 3057 17356
rect 3023 17322 3025 17340
rect 3025 17322 3057 17340
rect 3095 17322 3129 17356
rect 3167 17322 3201 17356
rect 3239 17340 3273 17356
rect 3239 17322 3267 17340
rect 3267 17322 3273 17340
rect 3311 17322 3345 17356
rect 3383 17340 3417 17356
rect 3383 17322 3405 17340
rect 3405 17322 3417 17340
rect 3455 17322 3489 17356
rect 3527 17340 3561 17356
rect 3527 17322 3543 17340
rect 3543 17322 3561 17340
rect 3599 17322 3633 17356
rect 3671 17340 3705 17356
rect 3671 17322 3681 17340
rect 3681 17322 3705 17340
rect 3743 17322 3777 17356
rect 3815 17340 3849 17356
rect 3815 17322 3819 17340
rect 3819 17322 3849 17340
rect 3887 17322 3921 17356
rect 3959 17340 3993 17356
rect 3959 17322 3991 17340
rect 3991 17322 3993 17340
rect 4031 17322 4065 17356
rect 4103 17340 4137 17356
rect 4103 17322 4129 17340
rect 4129 17322 4137 17340
rect 4175 17322 4209 17356
rect 4247 17340 4281 17356
rect 4247 17322 4267 17340
rect 4267 17322 4281 17340
rect 4319 17322 4353 17356
rect 4391 17340 4425 17356
rect 4391 17322 4405 17340
rect 4405 17322 4425 17340
rect 4463 17322 4497 17356
rect 4535 17340 4569 17356
rect 4535 17322 4543 17340
rect 4543 17322 4569 17340
rect 2663 17249 2697 17283
rect 2735 17249 2769 17283
rect 2807 17249 2841 17283
rect 2879 17249 2913 17283
rect 2951 17249 2985 17283
rect 3023 17249 3057 17283
rect 3095 17249 3129 17283
rect 3167 17249 3201 17283
rect 3239 17249 3273 17283
rect 3311 17249 3345 17283
rect 3383 17249 3417 17283
rect 3455 17249 3489 17283
rect 3527 17249 3561 17283
rect 3599 17249 3633 17283
rect 3671 17249 3705 17283
rect 3743 17249 3777 17283
rect 3815 17249 3849 17283
rect 3887 17249 3921 17283
rect 3959 17249 3993 17283
rect 4031 17249 4065 17283
rect 4103 17249 4137 17283
rect 4175 17249 4209 17283
rect 4247 17249 4281 17283
rect 4319 17249 4353 17283
rect 4391 17249 4425 17283
rect 4463 17249 4497 17283
rect 4535 17249 4569 17283
rect 8184 17363 8218 17397
rect 8050 17301 8084 17335
rect 8184 17291 8218 17325
rect 5251 17211 5255 17245
rect 5255 17211 5285 17245
rect 5325 17211 5359 17245
rect 5399 17211 5429 17245
rect 5429 17211 5433 17245
rect 5473 17211 5499 17245
rect 5499 17211 5507 17245
rect 5547 17211 5569 17245
rect 5569 17211 5581 17245
rect 5621 17211 5639 17245
rect 5639 17211 5655 17245
rect 5695 17211 5709 17245
rect 5709 17211 5729 17245
rect 5769 17211 5779 17245
rect 5779 17211 5803 17245
rect 5843 17211 5849 17245
rect 5849 17211 5877 17245
rect 5917 17211 5919 17245
rect 5919 17211 5951 17245
rect 5991 17211 6023 17245
rect 6023 17211 6025 17245
rect 6065 17211 6092 17245
rect 6092 17211 6099 17245
rect 6139 17211 6161 17245
rect 6161 17211 6173 17245
rect 6213 17211 6230 17245
rect 6230 17211 6247 17245
rect 6287 17211 6299 17245
rect 6299 17211 6321 17245
rect 6361 17211 6368 17245
rect 6368 17211 6395 17245
rect 6435 17211 6437 17245
rect 6437 17211 6469 17245
rect 6509 17211 6540 17245
rect 6540 17211 6543 17245
rect 6583 17211 6609 17245
rect 6609 17211 6617 17245
rect 6657 17211 6678 17245
rect 6678 17211 6691 17245
rect 6731 17211 6747 17245
rect 6747 17211 6765 17245
rect 6805 17211 6816 17245
rect 6816 17211 6839 17245
rect 6879 17211 6885 17245
rect 6885 17211 6913 17245
rect 6953 17211 6954 17245
rect 6954 17211 6987 17245
rect 7026 17211 7058 17245
rect 7058 17211 7060 17245
rect 7099 17211 7127 17245
rect 7127 17211 7133 17245
rect 7172 17211 7196 17245
rect 7196 17211 7206 17245
rect 7245 17211 7265 17245
rect 7265 17211 7279 17245
rect 7318 17211 7334 17245
rect 7334 17211 7352 17245
rect 7391 17211 7403 17245
rect 7403 17211 7425 17245
rect 7464 17211 7472 17245
rect 7472 17211 7498 17245
rect 7537 17211 7541 17245
rect 7541 17211 7571 17245
rect 7610 17211 7644 17245
rect 7683 17211 7713 17245
rect 7713 17211 7717 17245
rect 8050 17229 8084 17263
rect 8184 17219 8218 17253
rect 2663 17176 2697 17210
rect 2735 17203 2769 17210
rect 2735 17176 2749 17203
rect 2749 17176 2769 17203
rect 2807 17176 2841 17210
rect 2879 17203 2913 17210
rect 2879 17176 2887 17203
rect 2887 17176 2913 17203
rect 2951 17176 2985 17210
rect 3023 17203 3057 17210
rect 3023 17176 3025 17203
rect 3025 17176 3057 17203
rect 3095 17176 3129 17210
rect 3167 17176 3201 17210
rect 3239 17203 3273 17210
rect 3239 17176 3267 17203
rect 3267 17176 3273 17203
rect 3311 17176 3345 17210
rect 3383 17203 3417 17210
rect 3383 17176 3405 17203
rect 3405 17176 3417 17203
rect 3455 17176 3489 17210
rect 3527 17203 3561 17210
rect 3527 17176 3543 17203
rect 3543 17176 3561 17203
rect 3599 17176 3633 17210
rect 3671 17203 3705 17210
rect 3671 17176 3681 17203
rect 3681 17176 3705 17203
rect 3743 17176 3777 17210
rect 3815 17203 3849 17210
rect 3815 17176 3819 17203
rect 3819 17176 3849 17203
rect 3887 17176 3921 17210
rect 3959 17203 3993 17210
rect 3959 17176 3991 17203
rect 3991 17176 3993 17203
rect 4031 17176 4065 17210
rect 4103 17203 4137 17210
rect 4103 17176 4129 17203
rect 4129 17176 4137 17203
rect 4175 17176 4209 17210
rect 4247 17203 4281 17210
rect 4247 17176 4267 17203
rect 4267 17176 4281 17203
rect 4319 17176 4353 17210
rect 4391 17203 4425 17210
rect 4391 17176 4405 17203
rect 4405 17176 4425 17203
rect 4463 17176 4497 17210
rect 4535 17203 4569 17210
rect 4535 17176 4543 17203
rect 4543 17176 4569 17203
rect 2663 17103 2697 17137
rect 2735 17103 2769 17137
rect 2807 17103 2841 17137
rect 2879 17103 2913 17137
rect 2951 17103 2985 17137
rect 3023 17103 3057 17137
rect 3095 17103 3129 17137
rect 3167 17103 3201 17137
rect 3239 17103 3273 17137
rect 3311 17103 3345 17137
rect 3383 17103 3417 17137
rect 3455 17103 3489 17137
rect 3527 17103 3561 17137
rect 3599 17103 3633 17137
rect 3671 17103 3705 17137
rect 3743 17103 3777 17137
rect 3815 17103 3849 17137
rect 3887 17103 3921 17137
rect 3959 17103 3993 17137
rect 4031 17103 4065 17137
rect 4103 17103 4137 17137
rect 4175 17103 4209 17137
rect 4247 17103 4281 17137
rect 4319 17103 4353 17137
rect 4391 17103 4425 17137
rect 4463 17103 4497 17137
rect 4535 17103 4569 17137
rect 8050 17157 8084 17191
rect 8184 17147 8218 17181
rect 8050 17085 8084 17119
rect 8184 17075 8218 17109
rect 2663 17030 2697 17064
rect 2735 17032 2749 17064
rect 2749 17032 2769 17064
rect 2735 17030 2769 17032
rect 2807 17030 2841 17064
rect 2879 17032 2887 17064
rect 2887 17032 2913 17064
rect 2879 17030 2913 17032
rect 2951 17030 2985 17064
rect 3023 17032 3025 17064
rect 3025 17032 3057 17064
rect 3023 17030 3057 17032
rect 3095 17030 3129 17064
rect 3167 17030 3201 17064
rect 3239 17032 3267 17064
rect 3267 17032 3273 17064
rect 3239 17030 3273 17032
rect 3311 17030 3345 17064
rect 3383 17032 3405 17064
rect 3405 17032 3417 17064
rect 3383 17030 3417 17032
rect 3455 17030 3489 17064
rect 3527 17032 3543 17064
rect 3543 17032 3561 17064
rect 3527 17030 3561 17032
rect 3599 17030 3633 17064
rect 3671 17032 3681 17064
rect 3681 17032 3705 17064
rect 3671 17030 3705 17032
rect 3743 17030 3777 17064
rect 3815 17032 3819 17064
rect 3819 17032 3849 17064
rect 3815 17030 3849 17032
rect 3887 17030 3921 17064
rect 3959 17032 3991 17064
rect 3991 17032 3993 17064
rect 3959 17030 3993 17032
rect 4031 17030 4065 17064
rect 4103 17032 4129 17064
rect 4129 17032 4137 17064
rect 4103 17030 4137 17032
rect 4175 17030 4209 17064
rect 4247 17032 4267 17064
rect 4267 17032 4281 17064
rect 4247 17030 4281 17032
rect 4319 17030 4353 17064
rect 4391 17032 4405 17064
rect 4405 17032 4425 17064
rect 4391 17030 4425 17032
rect 4463 17030 4497 17064
rect 4535 17032 4543 17064
rect 4543 17032 4569 17064
rect 4535 17030 4569 17032
rect 2663 16957 2697 16991
rect 2735 16957 2769 16991
rect 2807 16957 2841 16991
rect 2879 16957 2913 16991
rect 2951 16957 2985 16991
rect 3023 16957 3057 16991
rect 3095 16957 3129 16991
rect 3167 16957 3201 16991
rect 3239 16957 3273 16991
rect 3311 16957 3345 16991
rect 3383 16957 3417 16991
rect 3455 16957 3489 16991
rect 3527 16957 3561 16991
rect 3599 16957 3633 16991
rect 3671 16957 3705 16991
rect 3743 16957 3777 16991
rect 3815 16957 3849 16991
rect 3887 16957 3921 16991
rect 3959 16957 3993 16991
rect 4031 16957 4065 16991
rect 4103 16957 4137 16991
rect 4175 16957 4209 16991
rect 4247 16957 4281 16991
rect 4319 16957 4353 16991
rect 4391 16957 4425 16991
rect 4463 16957 4497 16991
rect 4535 16957 4569 16991
rect 5089 16964 5123 16989
rect 5162 16964 5196 16989
rect 5235 16964 5269 16989
rect 5308 16964 5342 16989
rect 5381 16964 5415 16989
rect 5454 16964 5488 16989
rect 5527 16964 5561 16989
rect 5600 16964 5634 16989
rect 5673 16964 5707 16989
rect 5746 16964 5780 16989
rect 5819 16964 5853 16989
rect 5892 16964 5926 16989
rect 5965 16964 5999 16989
rect 6038 16964 6072 16989
rect 6110 16964 6144 16989
rect 6182 16964 6216 16989
rect 6254 16964 6288 16989
rect 6326 16964 6360 16989
rect 6398 16964 6432 16989
rect 6470 16964 6504 16989
rect 6542 16964 6576 16989
rect 6614 16964 6648 16989
rect 6686 16964 6720 16989
rect 6758 16964 6792 16989
rect 6830 16964 6864 16989
rect 6902 16964 6936 16989
rect 6974 16964 7008 16989
rect 7046 16964 7080 16989
rect 7118 16964 7152 16989
rect 5089 16955 5119 16964
rect 5119 16955 5123 16964
rect 5162 16955 5188 16964
rect 5188 16955 5196 16964
rect 5235 16955 5257 16964
rect 5257 16955 5269 16964
rect 5308 16955 5326 16964
rect 5326 16955 5342 16964
rect 5381 16955 5395 16964
rect 5395 16955 5415 16964
rect 5454 16955 5464 16964
rect 5464 16955 5488 16964
rect 5527 16955 5533 16964
rect 5533 16955 5561 16964
rect 5600 16955 5602 16964
rect 5602 16955 5634 16964
rect 5673 16955 5706 16964
rect 5706 16955 5707 16964
rect 5746 16955 5775 16964
rect 5775 16955 5780 16964
rect 5819 16955 5844 16964
rect 5844 16955 5853 16964
rect 5892 16955 5913 16964
rect 5913 16955 5926 16964
rect 5965 16955 5982 16964
rect 5982 16955 5999 16964
rect 6038 16955 6051 16964
rect 6051 16955 6072 16964
rect 6110 16955 6120 16964
rect 6120 16955 6144 16964
rect 6182 16955 6189 16964
rect 6189 16955 6216 16964
rect 6254 16955 6258 16964
rect 6258 16955 6288 16964
rect 6326 16955 6327 16964
rect 6327 16955 6360 16964
rect 6398 16955 6430 16964
rect 6430 16955 6432 16964
rect 6470 16955 6499 16964
rect 6499 16955 6504 16964
rect 6542 16955 6568 16964
rect 6568 16955 6576 16964
rect 6614 16955 6637 16964
rect 6637 16955 6648 16964
rect 6686 16955 6706 16964
rect 6706 16955 6720 16964
rect 6758 16955 6775 16964
rect 6775 16955 6792 16964
rect 6830 16955 6844 16964
rect 6844 16955 6864 16964
rect 6902 16955 6913 16964
rect 6913 16955 6936 16964
rect 6974 16955 6982 16964
rect 6982 16955 7008 16964
rect 7046 16955 7051 16964
rect 7051 16955 7080 16964
rect 7118 16955 7120 16964
rect 7120 16955 7152 16964
rect 7190 16955 7224 16989
rect 7262 16964 7296 16989
rect 7334 16964 7368 16989
rect 7406 16964 7440 16989
rect 7478 16964 7512 16989
rect 7550 16964 7584 16989
rect 7622 16964 7656 16989
rect 7694 16964 7728 16989
rect 7766 16964 7800 16989
rect 7838 16964 7872 16989
rect 7262 16955 7293 16964
rect 7293 16955 7296 16964
rect 7334 16955 7362 16964
rect 7362 16955 7368 16964
rect 7406 16955 7431 16964
rect 7431 16955 7440 16964
rect 7478 16955 7500 16964
rect 7500 16955 7512 16964
rect 7550 16955 7568 16964
rect 7568 16955 7584 16964
rect 7622 16955 7636 16964
rect 7636 16955 7656 16964
rect 7694 16955 7704 16964
rect 7704 16955 7728 16964
rect 7766 16955 7772 16964
rect 7772 16955 7800 16964
rect 7838 16955 7840 16964
rect 7840 16955 7872 16964
rect 2663 16884 2697 16918
rect 2735 16895 2749 16918
rect 2749 16895 2769 16918
rect 2735 16884 2769 16895
rect 2807 16884 2841 16918
rect 2879 16895 2887 16918
rect 2887 16895 2913 16918
rect 2879 16884 2913 16895
rect 2951 16884 2985 16918
rect 3023 16895 3025 16918
rect 3025 16895 3057 16918
rect 3023 16884 3057 16895
rect 3095 16884 3129 16918
rect 3167 16884 3201 16918
rect 3239 16895 3267 16918
rect 3267 16895 3273 16918
rect 3239 16884 3273 16895
rect 3311 16884 3345 16918
rect 3383 16895 3405 16918
rect 3405 16895 3417 16918
rect 3383 16884 3417 16895
rect 3455 16884 3489 16918
rect 3527 16895 3543 16918
rect 3543 16895 3561 16918
rect 3527 16884 3561 16895
rect 3599 16884 3633 16918
rect 3671 16895 3681 16918
rect 3681 16895 3705 16918
rect 3671 16884 3705 16895
rect 3743 16884 3777 16918
rect 3815 16895 3819 16918
rect 3819 16895 3849 16918
rect 3815 16884 3849 16895
rect 3887 16884 3921 16918
rect 3959 16895 3991 16918
rect 3991 16895 3993 16918
rect 3959 16884 3993 16895
rect 4031 16884 4065 16918
rect 4103 16895 4129 16918
rect 4129 16895 4137 16918
rect 4103 16884 4137 16895
rect 4175 16884 4209 16918
rect 4247 16895 4267 16918
rect 4267 16895 4281 16918
rect 4247 16884 4281 16895
rect 4319 16884 4353 16918
rect 4391 16895 4405 16918
rect 4405 16895 4425 16918
rect 4391 16884 4425 16895
rect 4463 16884 4497 16918
rect 4535 16895 4543 16918
rect 4543 16895 4569 16918
rect 4535 16884 4569 16895
rect 5089 16894 5123 16913
rect 5162 16894 5196 16913
rect 5235 16894 5269 16913
rect 5308 16894 5342 16913
rect 5381 16894 5415 16913
rect 5454 16894 5488 16913
rect 5527 16894 5561 16913
rect 5600 16894 5634 16913
rect 5673 16894 5707 16913
rect 5746 16894 5780 16913
rect 5819 16894 5853 16913
rect 5892 16894 5926 16913
rect 5965 16894 5999 16913
rect 6038 16894 6072 16913
rect 6110 16894 6144 16913
rect 6182 16894 6216 16913
rect 6254 16894 6288 16913
rect 6326 16894 6360 16913
rect 6398 16894 6432 16913
rect 6470 16894 6504 16913
rect 6542 16894 6576 16913
rect 6614 16894 6648 16913
rect 6686 16894 6720 16913
rect 6758 16894 6792 16913
rect 6830 16894 6864 16913
rect 6902 16894 6936 16913
rect 6974 16894 7008 16913
rect 7046 16894 7080 16913
rect 7118 16894 7152 16913
rect 5089 16879 5119 16894
rect 5119 16879 5123 16894
rect 5162 16879 5188 16894
rect 5188 16879 5196 16894
rect 5235 16879 5257 16894
rect 5257 16879 5269 16894
rect 5308 16879 5326 16894
rect 5326 16879 5342 16894
rect 5381 16879 5395 16894
rect 5395 16879 5415 16894
rect 5454 16879 5464 16894
rect 5464 16879 5488 16894
rect 5527 16879 5533 16894
rect 5533 16879 5561 16894
rect 5600 16879 5602 16894
rect 5602 16879 5634 16894
rect 5673 16879 5706 16894
rect 5706 16879 5707 16894
rect 5746 16879 5775 16894
rect 5775 16879 5780 16894
rect 5819 16879 5844 16894
rect 5844 16879 5853 16894
rect 5892 16879 5913 16894
rect 5913 16879 5926 16894
rect 5965 16879 5982 16894
rect 5982 16879 5999 16894
rect 6038 16879 6051 16894
rect 6051 16879 6072 16894
rect 6110 16879 6120 16894
rect 6120 16879 6144 16894
rect 6182 16879 6189 16894
rect 6189 16879 6216 16894
rect 6254 16879 6258 16894
rect 6258 16879 6288 16894
rect 6326 16879 6327 16894
rect 6327 16879 6360 16894
rect 6398 16879 6430 16894
rect 6430 16879 6432 16894
rect 6470 16879 6499 16894
rect 6499 16879 6504 16894
rect 6542 16879 6568 16894
rect 6568 16879 6576 16894
rect 6614 16879 6637 16894
rect 6637 16879 6648 16894
rect 6686 16879 6706 16894
rect 6706 16879 6720 16894
rect 6758 16879 6775 16894
rect 6775 16879 6792 16894
rect 6830 16879 6844 16894
rect 6844 16879 6864 16894
rect 6902 16879 6913 16894
rect 6913 16879 6936 16894
rect 6974 16879 6982 16894
rect 6982 16879 7008 16894
rect 7046 16879 7051 16894
rect 7051 16879 7080 16894
rect 7118 16879 7120 16894
rect 7120 16879 7152 16894
rect 7190 16879 7224 16913
rect 7262 16894 7296 16913
rect 7334 16894 7368 16913
rect 7406 16894 7440 16913
rect 7478 16894 7512 16913
rect 7550 16894 7584 16913
rect 7622 16894 7656 16913
rect 7694 16894 7728 16913
rect 7766 16894 7800 16913
rect 7838 16894 7872 16913
rect 7262 16879 7293 16894
rect 7293 16879 7296 16894
rect 7334 16879 7362 16894
rect 7362 16879 7368 16894
rect 7406 16879 7431 16894
rect 7431 16879 7440 16894
rect 7478 16879 7500 16894
rect 7500 16879 7512 16894
rect 7550 16879 7568 16894
rect 7568 16879 7584 16894
rect 7622 16879 7636 16894
rect 7636 16879 7656 16894
rect 7694 16879 7704 16894
rect 7704 16879 7728 16894
rect 7766 16879 7772 16894
rect 7772 16879 7800 16894
rect 7838 16879 7840 16894
rect 7840 16879 7872 16894
rect 2663 16811 2697 16845
rect 2735 16811 2769 16845
rect 2807 16811 2841 16845
rect 2879 16811 2913 16845
rect 2951 16811 2985 16845
rect 3023 16811 3057 16845
rect 3095 16811 3129 16845
rect 3167 16811 3201 16845
rect 3239 16811 3273 16845
rect 3311 16811 3345 16845
rect 3383 16811 3417 16845
rect 3455 16811 3489 16845
rect 3527 16811 3561 16845
rect 3599 16811 3633 16845
rect 3671 16811 3705 16845
rect 3743 16811 3777 16845
rect 3815 16811 3849 16845
rect 3887 16811 3921 16845
rect 3959 16811 3993 16845
rect 4031 16811 4065 16845
rect 4103 16811 4137 16845
rect 4175 16811 4209 16845
rect 4247 16811 4281 16845
rect 4319 16811 4353 16845
rect 4391 16811 4425 16845
rect 4463 16811 4497 16845
rect 4535 16811 4569 16845
rect 5089 16824 5123 16837
rect 5162 16824 5196 16837
rect 5235 16824 5269 16837
rect 5308 16824 5342 16837
rect 5381 16824 5415 16837
rect 5454 16824 5488 16837
rect 5527 16824 5561 16837
rect 5600 16824 5634 16837
rect 5673 16824 5707 16837
rect 5746 16824 5780 16837
rect 5819 16824 5853 16837
rect 5892 16824 5926 16837
rect 5965 16824 5999 16837
rect 6038 16824 6072 16837
rect 6110 16824 6144 16837
rect 6182 16824 6216 16837
rect 6254 16824 6288 16837
rect 6326 16824 6360 16837
rect 6398 16824 6432 16837
rect 6470 16824 6504 16837
rect 6542 16824 6576 16837
rect 6614 16824 6648 16837
rect 6686 16824 6720 16837
rect 6758 16824 6792 16837
rect 6830 16824 6864 16837
rect 6902 16824 6936 16837
rect 6974 16824 7008 16837
rect 7046 16824 7080 16837
rect 7118 16824 7152 16837
rect 2663 16738 2697 16772
rect 2735 16758 2749 16772
rect 2749 16758 2769 16772
rect 2735 16738 2769 16758
rect 2807 16738 2841 16772
rect 2879 16758 2887 16772
rect 2887 16758 2913 16772
rect 2879 16738 2913 16758
rect 2951 16738 2985 16772
rect 3023 16758 3025 16772
rect 3025 16758 3057 16772
rect 3023 16738 3057 16758
rect 3095 16738 3129 16772
rect 3167 16738 3201 16772
rect 3239 16758 3267 16772
rect 3267 16758 3273 16772
rect 3239 16738 3273 16758
rect 3311 16738 3345 16772
rect 3383 16758 3405 16772
rect 3405 16758 3417 16772
rect 3383 16738 3417 16758
rect 3455 16738 3489 16772
rect 3527 16758 3543 16772
rect 3543 16758 3561 16772
rect 3527 16738 3561 16758
rect 3599 16738 3633 16772
rect 3671 16758 3681 16772
rect 3681 16758 3705 16772
rect 3671 16738 3705 16758
rect 3743 16738 3777 16772
rect 3815 16758 3819 16772
rect 3819 16758 3849 16772
rect 3815 16738 3849 16758
rect 3887 16738 3921 16772
rect 3959 16758 3991 16772
rect 3991 16758 3993 16772
rect 3959 16738 3993 16758
rect 4031 16738 4065 16772
rect 4103 16758 4129 16772
rect 4129 16758 4137 16772
rect 4103 16738 4137 16758
rect 4175 16738 4209 16772
rect 4247 16758 4267 16772
rect 4267 16758 4281 16772
rect 4247 16738 4281 16758
rect 4319 16738 4353 16772
rect 4391 16758 4405 16772
rect 4405 16758 4425 16772
rect 4391 16738 4425 16758
rect 4463 16738 4497 16772
rect 4535 16758 4543 16772
rect 4543 16758 4569 16772
rect 5089 16803 5119 16824
rect 5119 16803 5123 16824
rect 5162 16803 5188 16824
rect 5188 16803 5196 16824
rect 5235 16803 5257 16824
rect 5257 16803 5269 16824
rect 5308 16803 5326 16824
rect 5326 16803 5342 16824
rect 5381 16803 5395 16824
rect 5395 16803 5415 16824
rect 5454 16803 5464 16824
rect 5464 16803 5488 16824
rect 5527 16803 5533 16824
rect 5533 16803 5561 16824
rect 5600 16803 5602 16824
rect 5602 16803 5634 16824
rect 5673 16803 5706 16824
rect 5706 16803 5707 16824
rect 5746 16803 5775 16824
rect 5775 16803 5780 16824
rect 5819 16803 5844 16824
rect 5844 16803 5853 16824
rect 5892 16803 5913 16824
rect 5913 16803 5926 16824
rect 5965 16803 5982 16824
rect 5982 16803 5999 16824
rect 6038 16803 6051 16824
rect 6051 16803 6072 16824
rect 6110 16803 6120 16824
rect 6120 16803 6144 16824
rect 6182 16803 6189 16824
rect 6189 16803 6216 16824
rect 6254 16803 6258 16824
rect 6258 16803 6288 16824
rect 6326 16803 6327 16824
rect 6327 16803 6360 16824
rect 6398 16803 6430 16824
rect 6430 16803 6432 16824
rect 6470 16803 6499 16824
rect 6499 16803 6504 16824
rect 6542 16803 6568 16824
rect 6568 16803 6576 16824
rect 6614 16803 6637 16824
rect 6637 16803 6648 16824
rect 6686 16803 6706 16824
rect 6706 16803 6720 16824
rect 6758 16803 6775 16824
rect 6775 16803 6792 16824
rect 6830 16803 6844 16824
rect 6844 16803 6864 16824
rect 6902 16803 6913 16824
rect 6913 16803 6936 16824
rect 6974 16803 6982 16824
rect 6982 16803 7008 16824
rect 7046 16803 7051 16824
rect 7051 16803 7080 16824
rect 7118 16803 7120 16824
rect 7120 16803 7152 16824
rect 7190 16803 7224 16837
rect 7262 16824 7296 16837
rect 7334 16824 7368 16837
rect 7406 16824 7440 16837
rect 7478 16824 7512 16837
rect 7550 16824 7584 16837
rect 7622 16824 7656 16837
rect 7694 16824 7728 16837
rect 7766 16824 7800 16837
rect 7838 16824 7872 16837
rect 7262 16803 7293 16824
rect 7293 16803 7296 16824
rect 7334 16803 7362 16824
rect 7362 16803 7368 16824
rect 7406 16803 7431 16824
rect 7431 16803 7440 16824
rect 7478 16803 7500 16824
rect 7500 16803 7512 16824
rect 7550 16803 7568 16824
rect 7568 16803 7584 16824
rect 7622 16803 7636 16824
rect 7636 16803 7656 16824
rect 7694 16803 7704 16824
rect 7704 16803 7728 16824
rect 7766 16803 7772 16824
rect 7772 16803 7800 16824
rect 7838 16803 7840 16824
rect 7840 16803 7872 16824
rect 4535 16738 4569 16758
rect 5089 16754 5123 16761
rect 5162 16754 5196 16761
rect 5235 16754 5269 16761
rect 5308 16754 5342 16761
rect 5381 16754 5415 16761
rect 5454 16754 5488 16761
rect 5527 16754 5561 16761
rect 5600 16754 5634 16761
rect 5673 16754 5707 16761
rect 5746 16754 5780 16761
rect 5819 16754 5853 16761
rect 5892 16754 5926 16761
rect 5965 16754 5999 16761
rect 6038 16754 6072 16761
rect 6110 16754 6144 16761
rect 6182 16754 6216 16761
rect 6254 16754 6288 16761
rect 6326 16754 6360 16761
rect 6398 16754 6432 16761
rect 6470 16754 6504 16761
rect 6542 16754 6576 16761
rect 6614 16754 6648 16761
rect 6686 16754 6720 16761
rect 6758 16754 6792 16761
rect 6830 16754 6864 16761
rect 6902 16754 6936 16761
rect 6974 16754 7008 16761
rect 7046 16754 7080 16761
rect 7118 16754 7152 16761
rect 5089 16727 5119 16754
rect 5119 16727 5123 16754
rect 5162 16727 5188 16754
rect 5188 16727 5196 16754
rect 5235 16727 5257 16754
rect 5257 16727 5269 16754
rect 5308 16727 5326 16754
rect 5326 16727 5342 16754
rect 5381 16727 5395 16754
rect 5395 16727 5415 16754
rect 5454 16727 5464 16754
rect 5464 16727 5488 16754
rect 5527 16727 5533 16754
rect 5533 16727 5561 16754
rect 5600 16727 5602 16754
rect 5602 16727 5634 16754
rect 5673 16727 5706 16754
rect 5706 16727 5707 16754
rect 5746 16727 5775 16754
rect 5775 16727 5780 16754
rect 5819 16727 5844 16754
rect 5844 16727 5853 16754
rect 5892 16727 5913 16754
rect 5913 16727 5926 16754
rect 5965 16727 5982 16754
rect 5982 16727 5999 16754
rect 6038 16727 6051 16754
rect 6051 16727 6072 16754
rect 6110 16727 6120 16754
rect 6120 16727 6144 16754
rect 6182 16727 6189 16754
rect 6189 16727 6216 16754
rect 6254 16727 6258 16754
rect 6258 16727 6288 16754
rect 6326 16727 6327 16754
rect 6327 16727 6360 16754
rect 6398 16727 6430 16754
rect 6430 16727 6432 16754
rect 6470 16727 6499 16754
rect 6499 16727 6504 16754
rect 6542 16727 6568 16754
rect 6568 16727 6576 16754
rect 6614 16727 6637 16754
rect 6637 16727 6648 16754
rect 6686 16727 6706 16754
rect 6706 16727 6720 16754
rect 6758 16727 6775 16754
rect 6775 16727 6792 16754
rect 6830 16727 6844 16754
rect 6844 16727 6864 16754
rect 6902 16727 6913 16754
rect 6913 16727 6936 16754
rect 6974 16727 6982 16754
rect 6982 16727 7008 16754
rect 7046 16727 7051 16754
rect 7051 16727 7080 16754
rect 7118 16727 7120 16754
rect 7120 16727 7152 16754
rect 7190 16727 7224 16761
rect 7262 16754 7296 16761
rect 7334 16754 7368 16761
rect 7406 16754 7440 16761
rect 7478 16754 7512 16761
rect 7550 16754 7584 16761
rect 7622 16754 7656 16761
rect 7694 16754 7728 16761
rect 7766 16754 7800 16761
rect 7838 16754 7872 16761
rect 7262 16727 7293 16754
rect 7293 16727 7296 16754
rect 7334 16727 7362 16754
rect 7362 16727 7368 16754
rect 7406 16727 7431 16754
rect 7431 16727 7440 16754
rect 7478 16727 7500 16754
rect 7500 16727 7512 16754
rect 7550 16727 7568 16754
rect 7568 16727 7584 16754
rect 7622 16727 7636 16754
rect 7636 16727 7656 16754
rect 7694 16727 7704 16754
rect 7704 16727 7728 16754
rect 7766 16727 7772 16754
rect 7772 16727 7800 16754
rect 7838 16727 7840 16754
rect 7840 16727 7872 16754
rect 2663 16665 2697 16699
rect 2735 16665 2769 16699
rect 2807 16665 2841 16699
rect 2879 16665 2913 16699
rect 2951 16665 2985 16699
rect 3023 16665 3057 16699
rect 3095 16665 3129 16699
rect 3167 16665 3201 16699
rect 3239 16665 3273 16699
rect 3311 16665 3345 16699
rect 3383 16665 3417 16699
rect 3455 16665 3489 16699
rect 3527 16665 3561 16699
rect 3599 16665 3633 16699
rect 3671 16665 3705 16699
rect 3743 16665 3777 16699
rect 3815 16665 3849 16699
rect 3887 16665 3921 16699
rect 3959 16665 3993 16699
rect 4031 16665 4065 16699
rect 4103 16665 4137 16699
rect 4175 16665 4209 16699
rect 4247 16665 4281 16699
rect 4319 16665 4353 16699
rect 4391 16665 4425 16699
rect 4463 16665 4497 16699
rect 4535 16665 4569 16699
rect 5089 16684 5123 16685
rect 5162 16684 5196 16685
rect 5235 16684 5269 16685
rect 5308 16684 5342 16685
rect 5381 16684 5415 16685
rect 5454 16684 5488 16685
rect 5527 16684 5561 16685
rect 5600 16684 5634 16685
rect 5673 16684 5707 16685
rect 5746 16684 5780 16685
rect 5819 16684 5853 16685
rect 5892 16684 5926 16685
rect 5965 16684 5999 16685
rect 6038 16684 6072 16685
rect 6110 16684 6144 16685
rect 6182 16684 6216 16685
rect 6254 16684 6288 16685
rect 6326 16684 6360 16685
rect 6398 16684 6432 16685
rect 6470 16684 6504 16685
rect 6542 16684 6576 16685
rect 6614 16684 6648 16685
rect 6686 16684 6720 16685
rect 6758 16684 6792 16685
rect 6830 16684 6864 16685
rect 6902 16684 6936 16685
rect 6974 16684 7008 16685
rect 7046 16684 7080 16685
rect 7118 16684 7152 16685
rect 2663 16592 2697 16626
rect 2735 16621 2749 16626
rect 2749 16621 2769 16626
rect 2735 16592 2769 16621
rect 2807 16592 2841 16626
rect 2879 16621 2887 16626
rect 2887 16621 2913 16626
rect 2879 16592 2913 16621
rect 2951 16592 2985 16626
rect 3023 16621 3025 16626
rect 3025 16621 3057 16626
rect 3023 16592 3057 16621
rect 3095 16592 3129 16626
rect 3167 16592 3201 16626
rect 3239 16621 3267 16626
rect 3267 16621 3273 16626
rect 3239 16592 3273 16621
rect 3311 16592 3345 16626
rect 3383 16621 3405 16626
rect 3405 16621 3417 16626
rect 3383 16592 3417 16621
rect 3455 16592 3489 16626
rect 3527 16621 3543 16626
rect 3543 16621 3561 16626
rect 3527 16592 3561 16621
rect 3599 16592 3633 16626
rect 3671 16621 3681 16626
rect 3681 16621 3705 16626
rect 3671 16592 3705 16621
rect 3743 16592 3777 16626
rect 3815 16621 3819 16626
rect 3819 16621 3849 16626
rect 3815 16592 3849 16621
rect 3887 16592 3921 16626
rect 3959 16621 3991 16626
rect 3991 16621 3993 16626
rect 3959 16592 3993 16621
rect 4031 16592 4065 16626
rect 4103 16621 4129 16626
rect 4129 16621 4137 16626
rect 4103 16592 4137 16621
rect 4175 16592 4209 16626
rect 4247 16621 4267 16626
rect 4267 16621 4281 16626
rect 4247 16592 4281 16621
rect 4319 16592 4353 16626
rect 4391 16621 4405 16626
rect 4405 16621 4425 16626
rect 4391 16592 4425 16621
rect 4463 16592 4497 16626
rect 4535 16621 4543 16626
rect 4543 16621 4569 16626
rect 5089 16651 5119 16684
rect 5119 16651 5123 16684
rect 5162 16651 5188 16684
rect 5188 16651 5196 16684
rect 5235 16651 5257 16684
rect 5257 16651 5269 16684
rect 5308 16651 5326 16684
rect 5326 16651 5342 16684
rect 5381 16651 5395 16684
rect 5395 16651 5415 16684
rect 5454 16651 5464 16684
rect 5464 16651 5488 16684
rect 5527 16651 5533 16684
rect 5533 16651 5561 16684
rect 5600 16651 5602 16684
rect 5602 16651 5634 16684
rect 5673 16651 5706 16684
rect 5706 16651 5707 16684
rect 5746 16651 5775 16684
rect 5775 16651 5780 16684
rect 5819 16651 5844 16684
rect 5844 16651 5853 16684
rect 5892 16651 5913 16684
rect 5913 16651 5926 16684
rect 5965 16651 5982 16684
rect 5982 16651 5999 16684
rect 6038 16651 6051 16684
rect 6051 16651 6072 16684
rect 6110 16651 6120 16684
rect 6120 16651 6144 16684
rect 6182 16651 6189 16684
rect 6189 16651 6216 16684
rect 6254 16651 6258 16684
rect 6258 16651 6288 16684
rect 6326 16651 6327 16684
rect 6327 16651 6360 16684
rect 6398 16651 6430 16684
rect 6430 16651 6432 16684
rect 6470 16651 6499 16684
rect 6499 16651 6504 16684
rect 6542 16651 6568 16684
rect 6568 16651 6576 16684
rect 6614 16651 6637 16684
rect 6637 16651 6648 16684
rect 6686 16651 6706 16684
rect 6706 16651 6720 16684
rect 6758 16651 6775 16684
rect 6775 16651 6792 16684
rect 6830 16651 6844 16684
rect 6844 16651 6864 16684
rect 6902 16651 6913 16684
rect 6913 16651 6936 16684
rect 6974 16651 6982 16684
rect 6982 16651 7008 16684
rect 7046 16651 7051 16684
rect 7051 16651 7080 16684
rect 7118 16651 7120 16684
rect 7120 16651 7152 16684
rect 7190 16651 7224 16685
rect 7262 16684 7296 16685
rect 7334 16684 7368 16685
rect 7406 16684 7440 16685
rect 7478 16684 7512 16685
rect 7550 16684 7584 16685
rect 7622 16684 7656 16685
rect 7694 16684 7728 16685
rect 7766 16684 7800 16685
rect 7838 16684 7872 16685
rect 7262 16651 7293 16684
rect 7293 16651 7296 16684
rect 7334 16651 7362 16684
rect 7362 16651 7368 16684
rect 7406 16651 7431 16684
rect 7431 16651 7440 16684
rect 7478 16651 7500 16684
rect 7500 16651 7512 16684
rect 7550 16651 7568 16684
rect 7568 16651 7584 16684
rect 7622 16651 7636 16684
rect 7636 16651 7656 16684
rect 7694 16651 7704 16684
rect 7704 16651 7728 16684
rect 7766 16651 7772 16684
rect 7772 16651 7800 16684
rect 7838 16651 7840 16684
rect 7840 16651 7872 16684
rect 4535 16592 4569 16621
rect 5089 16580 5119 16609
rect 5119 16580 5123 16609
rect 5162 16580 5188 16609
rect 5188 16580 5196 16609
rect 5235 16580 5257 16609
rect 5257 16580 5269 16609
rect 5308 16580 5326 16609
rect 5326 16580 5342 16609
rect 5381 16580 5395 16609
rect 5395 16580 5415 16609
rect 5454 16580 5464 16609
rect 5464 16580 5488 16609
rect 5527 16580 5533 16609
rect 5533 16580 5561 16609
rect 5600 16580 5602 16609
rect 5602 16580 5634 16609
rect 5673 16580 5706 16609
rect 5706 16580 5707 16609
rect 5746 16580 5775 16609
rect 5775 16580 5780 16609
rect 5819 16580 5844 16609
rect 5844 16580 5853 16609
rect 5892 16580 5913 16609
rect 5913 16580 5926 16609
rect 5965 16580 5982 16609
rect 5982 16580 5999 16609
rect 6038 16580 6051 16609
rect 6051 16580 6072 16609
rect 6110 16580 6120 16609
rect 6120 16580 6144 16609
rect 6182 16580 6189 16609
rect 6189 16580 6216 16609
rect 6254 16580 6258 16609
rect 6258 16580 6288 16609
rect 6326 16580 6327 16609
rect 6327 16580 6360 16609
rect 6398 16580 6430 16609
rect 6430 16580 6432 16609
rect 6470 16580 6499 16609
rect 6499 16580 6504 16609
rect 6542 16580 6568 16609
rect 6568 16580 6576 16609
rect 6614 16580 6637 16609
rect 6637 16580 6648 16609
rect 6686 16580 6706 16609
rect 6706 16580 6720 16609
rect 6758 16580 6775 16609
rect 6775 16580 6792 16609
rect 6830 16580 6844 16609
rect 6844 16580 6864 16609
rect 6902 16580 6913 16609
rect 6913 16580 6936 16609
rect 6974 16580 6982 16609
rect 6982 16580 7008 16609
rect 7046 16580 7051 16609
rect 7051 16580 7080 16609
rect 7118 16580 7120 16609
rect 7120 16580 7152 16609
rect 5089 16575 5123 16580
rect 5162 16575 5196 16580
rect 5235 16575 5269 16580
rect 5308 16575 5342 16580
rect 5381 16575 5415 16580
rect 5454 16575 5488 16580
rect 5527 16575 5561 16580
rect 5600 16575 5634 16580
rect 5673 16575 5707 16580
rect 5746 16575 5780 16580
rect 5819 16575 5853 16580
rect 5892 16575 5926 16580
rect 5965 16575 5999 16580
rect 6038 16575 6072 16580
rect 6110 16575 6144 16580
rect 6182 16575 6216 16580
rect 6254 16575 6288 16580
rect 6326 16575 6360 16580
rect 6398 16575 6432 16580
rect 6470 16575 6504 16580
rect 6542 16575 6576 16580
rect 6614 16575 6648 16580
rect 6686 16575 6720 16580
rect 6758 16575 6792 16580
rect 6830 16575 6864 16580
rect 6902 16575 6936 16580
rect 6974 16575 7008 16580
rect 7046 16575 7080 16580
rect 7118 16575 7152 16580
rect 7190 16575 7224 16609
rect 7262 16580 7293 16609
rect 7293 16580 7296 16609
rect 7334 16580 7362 16609
rect 7362 16580 7368 16609
rect 7406 16580 7431 16609
rect 7431 16580 7440 16609
rect 7478 16580 7500 16609
rect 7500 16580 7512 16609
rect 7550 16580 7568 16609
rect 7568 16580 7584 16609
rect 7622 16580 7636 16609
rect 7636 16580 7656 16609
rect 7694 16580 7704 16609
rect 7704 16580 7728 16609
rect 7766 16580 7772 16609
rect 7772 16580 7800 16609
rect 7838 16580 7840 16609
rect 7840 16580 7872 16609
rect 7262 16575 7296 16580
rect 7334 16575 7368 16580
rect 7406 16575 7440 16580
rect 7478 16575 7512 16580
rect 7550 16575 7584 16580
rect 7622 16575 7656 16580
rect 7694 16575 7728 16580
rect 7766 16575 7800 16580
rect 7838 16575 7872 16580
rect 2663 16519 2697 16553
rect 2735 16519 2769 16553
rect 2807 16519 2841 16553
rect 2879 16519 2913 16553
rect 2951 16519 2985 16553
rect 3023 16519 3057 16553
rect 3095 16519 3129 16553
rect 3167 16519 3201 16553
rect 3239 16519 3273 16553
rect 3311 16519 3345 16553
rect 3383 16519 3417 16553
rect 3455 16519 3489 16553
rect 3527 16519 3561 16553
rect 3599 16519 3633 16553
rect 3671 16519 3705 16553
rect 3743 16519 3777 16553
rect 3815 16519 3849 16553
rect 3887 16519 3921 16553
rect 3959 16519 3993 16553
rect 4031 16519 4065 16553
rect 4103 16519 4137 16553
rect 4175 16519 4209 16553
rect 4247 16519 4281 16553
rect 4319 16519 4353 16553
rect 4391 16519 4425 16553
rect 4463 16519 4497 16553
rect 4535 16519 4569 16553
rect 5089 16510 5119 16533
rect 5119 16510 5123 16533
rect 5162 16510 5188 16533
rect 5188 16510 5196 16533
rect 5235 16510 5257 16533
rect 5257 16510 5269 16533
rect 5308 16510 5326 16533
rect 5326 16510 5342 16533
rect 5381 16510 5395 16533
rect 5395 16510 5415 16533
rect 5454 16510 5464 16533
rect 5464 16510 5488 16533
rect 5527 16510 5533 16533
rect 5533 16510 5561 16533
rect 5600 16510 5602 16533
rect 5602 16510 5634 16533
rect 5673 16510 5706 16533
rect 5706 16510 5707 16533
rect 5746 16510 5775 16533
rect 5775 16510 5780 16533
rect 5819 16510 5844 16533
rect 5844 16510 5853 16533
rect 5892 16510 5913 16533
rect 5913 16510 5926 16533
rect 5965 16510 5982 16533
rect 5982 16510 5999 16533
rect 6038 16510 6051 16533
rect 6051 16510 6072 16533
rect 6110 16510 6120 16533
rect 6120 16510 6144 16533
rect 6182 16510 6189 16533
rect 6189 16510 6216 16533
rect 6254 16510 6258 16533
rect 6258 16510 6288 16533
rect 6326 16510 6327 16533
rect 6327 16510 6360 16533
rect 6398 16510 6430 16533
rect 6430 16510 6432 16533
rect 6470 16510 6499 16533
rect 6499 16510 6504 16533
rect 6542 16510 6568 16533
rect 6568 16510 6576 16533
rect 6614 16510 6637 16533
rect 6637 16510 6648 16533
rect 6686 16510 6706 16533
rect 6706 16510 6720 16533
rect 6758 16510 6775 16533
rect 6775 16510 6792 16533
rect 6830 16510 6844 16533
rect 6844 16510 6864 16533
rect 6902 16510 6913 16533
rect 6913 16510 6936 16533
rect 6974 16510 6982 16533
rect 6982 16510 7008 16533
rect 7046 16510 7051 16533
rect 7051 16510 7080 16533
rect 7118 16510 7120 16533
rect 7120 16510 7152 16533
rect 5089 16499 5123 16510
rect 5162 16499 5196 16510
rect 5235 16499 5269 16510
rect 5308 16499 5342 16510
rect 5381 16499 5415 16510
rect 5454 16499 5488 16510
rect 5527 16499 5561 16510
rect 5600 16499 5634 16510
rect 5673 16499 5707 16510
rect 5746 16499 5780 16510
rect 5819 16499 5853 16510
rect 5892 16499 5926 16510
rect 5965 16499 5999 16510
rect 6038 16499 6072 16510
rect 6110 16499 6144 16510
rect 6182 16499 6216 16510
rect 6254 16499 6288 16510
rect 6326 16499 6360 16510
rect 6398 16499 6432 16510
rect 6470 16499 6504 16510
rect 6542 16499 6576 16510
rect 6614 16499 6648 16510
rect 6686 16499 6720 16510
rect 6758 16499 6792 16510
rect 6830 16499 6864 16510
rect 6902 16499 6936 16510
rect 6974 16499 7008 16510
rect 7046 16499 7080 16510
rect 7118 16499 7152 16510
rect 7190 16499 7224 16533
rect 7262 16510 7293 16533
rect 7293 16510 7296 16533
rect 7334 16510 7362 16533
rect 7362 16510 7368 16533
rect 7406 16510 7431 16533
rect 7431 16510 7440 16533
rect 7478 16510 7500 16533
rect 7500 16510 7512 16533
rect 7550 16510 7568 16533
rect 7568 16510 7584 16533
rect 7622 16510 7636 16533
rect 7636 16510 7656 16533
rect 7694 16510 7704 16533
rect 7704 16510 7728 16533
rect 7766 16510 7772 16533
rect 7772 16510 7800 16533
rect 7838 16510 7840 16533
rect 7840 16510 7872 16533
rect 7262 16499 7296 16510
rect 7334 16499 7368 16510
rect 7406 16499 7440 16510
rect 7478 16499 7512 16510
rect 7550 16499 7584 16510
rect 7622 16499 7656 16510
rect 7694 16499 7728 16510
rect 7766 16499 7800 16510
rect 7838 16499 7872 16510
rect 2663 16446 2697 16480
rect 2735 16446 2769 16480
rect 2807 16446 2841 16480
rect 2879 16446 2913 16480
rect 2951 16446 2985 16480
rect 3023 16446 3057 16480
rect 3095 16446 3129 16480
rect 3167 16446 3201 16480
rect 3239 16446 3273 16480
rect 3311 16446 3345 16480
rect 3383 16446 3417 16480
rect 3455 16446 3489 16480
rect 3527 16446 3561 16480
rect 3599 16446 3633 16480
rect 3671 16446 3705 16480
rect 3743 16446 3777 16480
rect 3815 16446 3849 16480
rect 3887 16446 3921 16480
rect 3959 16446 3993 16480
rect 4031 16446 4065 16480
rect 4103 16446 4137 16480
rect 4175 16446 4209 16480
rect 4247 16446 4281 16480
rect 4319 16446 4353 16480
rect 4391 16446 4425 16480
rect 4463 16446 4497 16480
rect 4535 16446 4569 16480
rect 5089 16440 5119 16457
rect 5119 16440 5123 16457
rect 5162 16440 5188 16457
rect 5188 16440 5196 16457
rect 5235 16440 5257 16457
rect 5257 16440 5269 16457
rect 5308 16440 5326 16457
rect 5326 16440 5342 16457
rect 5381 16440 5395 16457
rect 5395 16440 5415 16457
rect 5454 16440 5464 16457
rect 5464 16440 5488 16457
rect 5527 16440 5533 16457
rect 5533 16440 5561 16457
rect 5600 16440 5602 16457
rect 5602 16440 5634 16457
rect 5673 16440 5706 16457
rect 5706 16440 5707 16457
rect 5746 16440 5775 16457
rect 5775 16440 5780 16457
rect 5819 16440 5844 16457
rect 5844 16440 5853 16457
rect 5892 16440 5913 16457
rect 5913 16440 5926 16457
rect 5965 16440 5982 16457
rect 5982 16440 5999 16457
rect 6038 16440 6051 16457
rect 6051 16440 6072 16457
rect 6110 16440 6120 16457
rect 6120 16440 6144 16457
rect 6182 16440 6189 16457
rect 6189 16440 6216 16457
rect 6254 16440 6258 16457
rect 6258 16440 6288 16457
rect 6326 16440 6327 16457
rect 6327 16440 6360 16457
rect 6398 16440 6430 16457
rect 6430 16440 6432 16457
rect 6470 16440 6499 16457
rect 6499 16440 6504 16457
rect 6542 16440 6568 16457
rect 6568 16440 6576 16457
rect 6614 16440 6637 16457
rect 6637 16440 6648 16457
rect 6686 16440 6706 16457
rect 6706 16440 6720 16457
rect 6758 16440 6775 16457
rect 6775 16440 6792 16457
rect 6830 16440 6844 16457
rect 6844 16440 6864 16457
rect 6902 16440 6913 16457
rect 6913 16440 6936 16457
rect 6974 16440 6982 16457
rect 6982 16440 7008 16457
rect 7046 16440 7051 16457
rect 7051 16440 7080 16457
rect 7118 16440 7120 16457
rect 7120 16440 7152 16457
rect 5089 16423 5123 16440
rect 5162 16423 5196 16440
rect 5235 16423 5269 16440
rect 5308 16423 5342 16440
rect 5381 16423 5415 16440
rect 5454 16423 5488 16440
rect 5527 16423 5561 16440
rect 5600 16423 5634 16440
rect 5673 16423 5707 16440
rect 5746 16423 5780 16440
rect 5819 16423 5853 16440
rect 5892 16423 5926 16440
rect 5965 16423 5999 16440
rect 6038 16423 6072 16440
rect 6110 16423 6144 16440
rect 6182 16423 6216 16440
rect 6254 16423 6288 16440
rect 6326 16423 6360 16440
rect 6398 16423 6432 16440
rect 6470 16423 6504 16440
rect 6542 16423 6576 16440
rect 6614 16423 6648 16440
rect 6686 16423 6720 16440
rect 6758 16423 6792 16440
rect 6830 16423 6864 16440
rect 6902 16423 6936 16440
rect 6974 16423 7008 16440
rect 7046 16423 7080 16440
rect 7118 16423 7152 16440
rect 7190 16423 7224 16457
rect 7262 16440 7293 16457
rect 7293 16440 7296 16457
rect 7334 16440 7362 16457
rect 7362 16440 7368 16457
rect 7406 16440 7431 16457
rect 7431 16440 7440 16457
rect 7478 16440 7500 16457
rect 7500 16440 7512 16457
rect 7550 16440 7568 16457
rect 7568 16440 7584 16457
rect 7622 16440 7636 16457
rect 7636 16440 7656 16457
rect 7694 16440 7704 16457
rect 7704 16440 7728 16457
rect 7766 16440 7772 16457
rect 7772 16440 7800 16457
rect 7838 16440 7840 16457
rect 7840 16440 7872 16457
rect 7262 16423 7296 16440
rect 7334 16423 7368 16440
rect 7406 16423 7440 16440
rect 7478 16423 7512 16440
rect 7550 16423 7584 16440
rect 7622 16423 7656 16440
rect 7694 16423 7728 16440
rect 7766 16423 7800 16440
rect 7838 16423 7872 16440
rect 2663 16373 2697 16407
rect 2735 16381 2769 16407
rect 2735 16373 2749 16381
rect 2749 16373 2769 16381
rect 2807 16373 2841 16407
rect 2879 16381 2913 16407
rect 2879 16373 2887 16381
rect 2887 16373 2913 16381
rect 2951 16373 2985 16407
rect 3023 16381 3057 16407
rect 3023 16373 3025 16381
rect 3025 16373 3057 16381
rect 3095 16373 3129 16407
rect 3167 16373 3201 16407
rect 3239 16381 3273 16407
rect 3239 16373 3267 16381
rect 3267 16373 3273 16381
rect 3311 16373 3345 16407
rect 3383 16381 3417 16407
rect 3383 16373 3405 16381
rect 3405 16373 3417 16381
rect 3455 16373 3489 16407
rect 3527 16381 3561 16407
rect 3527 16373 3543 16381
rect 3543 16373 3561 16381
rect 3599 16373 3633 16407
rect 3671 16381 3705 16407
rect 3671 16373 3681 16381
rect 3681 16373 3705 16381
rect 3743 16373 3777 16407
rect 3815 16381 3849 16407
rect 3815 16373 3819 16381
rect 3819 16373 3849 16381
rect 3887 16373 3921 16407
rect 3959 16381 3993 16407
rect 3959 16373 3991 16381
rect 3991 16373 3993 16381
rect 4031 16373 4065 16407
rect 4103 16381 4137 16407
rect 4103 16373 4129 16381
rect 4129 16373 4137 16381
rect 4175 16373 4209 16407
rect 4247 16381 4281 16407
rect 4247 16373 4267 16381
rect 4267 16373 4281 16381
rect 4319 16373 4353 16407
rect 4391 16381 4425 16407
rect 4391 16373 4405 16381
rect 4405 16373 4425 16381
rect 4463 16373 4497 16407
rect 4535 16381 4569 16407
rect 4535 16373 4543 16381
rect 4543 16373 4569 16381
rect 5089 16370 5119 16381
rect 5119 16370 5123 16381
rect 5162 16370 5188 16381
rect 5188 16370 5196 16381
rect 5235 16370 5257 16381
rect 5257 16370 5269 16381
rect 5308 16370 5326 16381
rect 5326 16370 5342 16381
rect 5381 16370 5395 16381
rect 5395 16370 5415 16381
rect 5454 16370 5464 16381
rect 5464 16370 5488 16381
rect 5527 16370 5533 16381
rect 5533 16370 5561 16381
rect 5600 16370 5602 16381
rect 5602 16370 5634 16381
rect 5673 16370 5706 16381
rect 5706 16370 5707 16381
rect 5746 16370 5775 16381
rect 5775 16370 5780 16381
rect 5819 16370 5844 16381
rect 5844 16370 5853 16381
rect 5892 16370 5913 16381
rect 5913 16370 5926 16381
rect 5965 16370 5982 16381
rect 5982 16370 5999 16381
rect 6038 16370 6051 16381
rect 6051 16370 6072 16381
rect 6110 16370 6120 16381
rect 6120 16370 6144 16381
rect 6182 16370 6189 16381
rect 6189 16370 6216 16381
rect 6254 16370 6258 16381
rect 6258 16370 6288 16381
rect 6326 16370 6327 16381
rect 6327 16370 6360 16381
rect 6398 16370 6430 16381
rect 6430 16370 6432 16381
rect 6470 16370 6499 16381
rect 6499 16370 6504 16381
rect 6542 16370 6568 16381
rect 6568 16370 6576 16381
rect 6614 16370 6637 16381
rect 6637 16370 6648 16381
rect 6686 16370 6706 16381
rect 6706 16370 6720 16381
rect 6758 16370 6775 16381
rect 6775 16370 6792 16381
rect 6830 16370 6844 16381
rect 6844 16370 6864 16381
rect 6902 16370 6913 16381
rect 6913 16370 6936 16381
rect 6974 16370 6982 16381
rect 6982 16370 7008 16381
rect 7046 16370 7051 16381
rect 7051 16370 7080 16381
rect 7118 16370 7120 16381
rect 7120 16370 7152 16381
rect 5089 16347 5123 16370
rect 5162 16347 5196 16370
rect 5235 16347 5269 16370
rect 5308 16347 5342 16370
rect 5381 16347 5415 16370
rect 5454 16347 5488 16370
rect 5527 16347 5561 16370
rect 5600 16347 5634 16370
rect 5673 16347 5707 16370
rect 5746 16347 5780 16370
rect 5819 16347 5853 16370
rect 5892 16347 5926 16370
rect 5965 16347 5999 16370
rect 6038 16347 6072 16370
rect 6110 16347 6144 16370
rect 6182 16347 6216 16370
rect 6254 16347 6288 16370
rect 6326 16347 6360 16370
rect 6398 16347 6432 16370
rect 6470 16347 6504 16370
rect 6542 16347 6576 16370
rect 6614 16347 6648 16370
rect 6686 16347 6720 16370
rect 6758 16347 6792 16370
rect 6830 16347 6864 16370
rect 6902 16347 6936 16370
rect 6974 16347 7008 16370
rect 7046 16347 7080 16370
rect 7118 16347 7152 16370
rect 7190 16347 7224 16381
rect 7262 16370 7293 16381
rect 7293 16370 7296 16381
rect 7334 16370 7362 16381
rect 7362 16370 7368 16381
rect 7406 16370 7431 16381
rect 7431 16370 7440 16381
rect 7478 16370 7500 16381
rect 7500 16370 7512 16381
rect 7550 16370 7568 16381
rect 7568 16370 7584 16381
rect 7622 16370 7636 16381
rect 7636 16370 7656 16381
rect 7694 16370 7704 16381
rect 7704 16370 7728 16381
rect 7766 16370 7772 16381
rect 7772 16370 7800 16381
rect 7838 16370 7840 16381
rect 7840 16370 7872 16381
rect 7262 16347 7296 16370
rect 7334 16347 7368 16370
rect 7406 16347 7440 16370
rect 7478 16347 7512 16370
rect 7550 16347 7584 16370
rect 7622 16347 7656 16370
rect 7694 16347 7728 16370
rect 7766 16347 7800 16370
rect 7838 16347 7872 16370
rect 2663 16300 2697 16334
rect 2735 16300 2769 16334
rect 2807 16300 2841 16334
rect 2879 16300 2913 16334
rect 2951 16300 2985 16334
rect 3023 16300 3057 16334
rect 3095 16300 3129 16334
rect 3167 16300 3201 16334
rect 3239 16300 3273 16334
rect 3311 16300 3345 16334
rect 3383 16300 3417 16334
rect 3455 16300 3489 16334
rect 3527 16300 3561 16334
rect 3599 16300 3633 16334
rect 3671 16300 3705 16334
rect 3743 16300 3777 16334
rect 3815 16300 3849 16334
rect 3887 16300 3921 16334
rect 3959 16300 3993 16334
rect 4031 16300 4065 16334
rect 4103 16300 4137 16334
rect 4175 16300 4209 16334
rect 4247 16300 4281 16334
rect 4319 16300 4353 16334
rect 4391 16300 4425 16334
rect 4463 16300 4497 16334
rect 4535 16300 4569 16334
rect 5089 16300 5119 16305
rect 5119 16300 5123 16305
rect 5162 16300 5188 16305
rect 5188 16300 5196 16305
rect 5235 16300 5257 16305
rect 5257 16300 5269 16305
rect 5308 16300 5326 16305
rect 5326 16300 5342 16305
rect 5381 16300 5395 16305
rect 5395 16300 5415 16305
rect 5454 16300 5464 16305
rect 5464 16300 5488 16305
rect 5527 16300 5533 16305
rect 5533 16300 5561 16305
rect 5600 16300 5602 16305
rect 5602 16300 5634 16305
rect 5673 16300 5706 16305
rect 5706 16300 5707 16305
rect 5746 16300 5775 16305
rect 5775 16300 5780 16305
rect 5819 16300 5844 16305
rect 5844 16300 5853 16305
rect 5892 16300 5913 16305
rect 5913 16300 5926 16305
rect 5965 16300 5982 16305
rect 5982 16300 5999 16305
rect 6038 16300 6051 16305
rect 6051 16300 6072 16305
rect 6110 16300 6120 16305
rect 6120 16300 6144 16305
rect 6182 16300 6189 16305
rect 6189 16300 6216 16305
rect 6254 16300 6258 16305
rect 6258 16300 6288 16305
rect 6326 16300 6327 16305
rect 6327 16300 6360 16305
rect 6398 16300 6430 16305
rect 6430 16300 6432 16305
rect 6470 16300 6499 16305
rect 6499 16300 6504 16305
rect 6542 16300 6568 16305
rect 6568 16300 6576 16305
rect 6614 16300 6637 16305
rect 6637 16300 6648 16305
rect 6686 16300 6706 16305
rect 6706 16300 6720 16305
rect 6758 16300 6775 16305
rect 6775 16300 6792 16305
rect 6830 16300 6844 16305
rect 6844 16300 6864 16305
rect 6902 16300 6913 16305
rect 6913 16300 6936 16305
rect 6974 16300 6982 16305
rect 6982 16300 7008 16305
rect 7046 16300 7051 16305
rect 7051 16300 7080 16305
rect 7118 16300 7120 16305
rect 7120 16300 7152 16305
rect 5089 16271 5123 16300
rect 5162 16271 5196 16300
rect 5235 16271 5269 16300
rect 5308 16271 5342 16300
rect 5381 16271 5415 16300
rect 5454 16271 5488 16300
rect 5527 16271 5561 16300
rect 5600 16271 5634 16300
rect 5673 16271 5707 16300
rect 5746 16271 5780 16300
rect 5819 16271 5853 16300
rect 5892 16271 5926 16300
rect 5965 16271 5999 16300
rect 6038 16271 6072 16300
rect 6110 16271 6144 16300
rect 6182 16271 6216 16300
rect 6254 16271 6288 16300
rect 6326 16271 6360 16300
rect 6398 16271 6432 16300
rect 6470 16271 6504 16300
rect 6542 16271 6576 16300
rect 6614 16271 6648 16300
rect 6686 16271 6720 16300
rect 6758 16271 6792 16300
rect 6830 16271 6864 16300
rect 6902 16271 6936 16300
rect 6974 16271 7008 16300
rect 7046 16271 7080 16300
rect 7118 16271 7152 16300
rect 7190 16271 7224 16305
rect 7262 16300 7293 16305
rect 7293 16300 7296 16305
rect 7334 16300 7362 16305
rect 7362 16300 7368 16305
rect 7406 16300 7431 16305
rect 7431 16300 7440 16305
rect 7478 16300 7500 16305
rect 7500 16300 7512 16305
rect 7550 16300 7568 16305
rect 7568 16300 7584 16305
rect 7622 16300 7636 16305
rect 7636 16300 7656 16305
rect 7694 16300 7704 16305
rect 7704 16300 7728 16305
rect 7766 16300 7772 16305
rect 7772 16300 7800 16305
rect 7838 16300 7840 16305
rect 7840 16300 7872 16305
rect 7262 16271 7296 16300
rect 7334 16271 7368 16300
rect 7406 16271 7440 16300
rect 7478 16271 7512 16300
rect 7550 16271 7584 16300
rect 7622 16271 7656 16300
rect 7694 16271 7728 16300
rect 7766 16271 7800 16300
rect 7838 16271 7872 16300
rect 2663 16227 2697 16261
rect 2735 16244 2769 16261
rect 2735 16227 2749 16244
rect 2749 16227 2769 16244
rect 2807 16227 2841 16261
rect 2879 16244 2913 16261
rect 2879 16227 2887 16244
rect 2887 16227 2913 16244
rect 2951 16227 2985 16261
rect 3023 16244 3057 16261
rect 3023 16227 3025 16244
rect 3025 16227 3057 16244
rect 3095 16227 3129 16261
rect 3167 16227 3201 16261
rect 3239 16244 3273 16261
rect 3239 16227 3267 16244
rect 3267 16227 3273 16244
rect 3311 16227 3345 16261
rect 3383 16244 3417 16261
rect 3383 16227 3405 16244
rect 3405 16227 3417 16244
rect 3455 16227 3489 16261
rect 3527 16244 3561 16261
rect 3527 16227 3543 16244
rect 3543 16227 3561 16244
rect 3599 16227 3633 16261
rect 3671 16244 3705 16261
rect 3671 16227 3681 16244
rect 3681 16227 3705 16244
rect 3743 16227 3777 16261
rect 3815 16244 3849 16261
rect 3815 16227 3819 16244
rect 3819 16227 3849 16244
rect 3887 16227 3921 16261
rect 3959 16244 3993 16261
rect 3959 16227 3991 16244
rect 3991 16227 3993 16244
rect 4031 16227 4065 16261
rect 4103 16244 4137 16261
rect 4103 16227 4129 16244
rect 4129 16227 4137 16244
rect 4175 16227 4209 16261
rect 4247 16244 4281 16261
rect 4247 16227 4267 16244
rect 4267 16227 4281 16244
rect 4319 16227 4353 16261
rect 4391 16244 4425 16261
rect 4391 16227 4405 16244
rect 4405 16227 4425 16244
rect 4463 16227 4497 16261
rect 4535 16244 4569 16261
rect 4535 16227 4543 16244
rect 4543 16227 4569 16244
rect 5089 16195 5123 16229
rect 5162 16195 5196 16229
rect 5235 16195 5269 16229
rect 5308 16195 5342 16229
rect 5381 16195 5415 16229
rect 5454 16195 5488 16229
rect 5527 16195 5561 16229
rect 5600 16195 5634 16229
rect 5673 16195 5707 16229
rect 5746 16195 5780 16229
rect 5819 16195 5853 16229
rect 5892 16195 5926 16229
rect 5965 16195 5999 16229
rect 6038 16195 6072 16229
rect 6110 16195 6144 16229
rect 6182 16195 6216 16229
rect 6254 16195 6288 16229
rect 6326 16195 6360 16229
rect 6398 16195 6432 16229
rect 6470 16195 6504 16229
rect 6542 16195 6576 16229
rect 6614 16195 6648 16229
rect 6686 16195 6720 16229
rect 6758 16195 6792 16229
rect 6830 16195 6864 16229
rect 6902 16195 6936 16229
rect 6974 16195 7008 16229
rect 7046 16195 7080 16229
rect 7118 16195 7152 16229
rect 7190 16195 7224 16229
rect 7262 16195 7296 16229
rect 7334 16195 7368 16229
rect 7406 16195 7440 16229
rect 7478 16195 7512 16229
rect 7550 16195 7584 16229
rect 7622 16195 7656 16229
rect 7694 16195 7728 16229
rect 7766 16195 7800 16229
rect 7838 16195 7872 16229
rect 2663 16154 2697 16188
rect 2735 16154 2769 16188
rect 2807 16154 2841 16188
rect 2879 16154 2913 16188
rect 2951 16154 2985 16188
rect 3023 16154 3057 16188
rect 3095 16154 3129 16188
rect 3167 16154 3201 16188
rect 3239 16154 3273 16188
rect 3311 16154 3345 16188
rect 3383 16154 3417 16188
rect 3455 16154 3489 16188
rect 3527 16154 3561 16188
rect 3599 16154 3633 16188
rect 3671 16154 3705 16188
rect 3743 16154 3777 16188
rect 3815 16154 3849 16188
rect 3887 16154 3921 16188
rect 3959 16154 3993 16188
rect 4031 16154 4065 16188
rect 4103 16154 4137 16188
rect 4175 16154 4209 16188
rect 4247 16154 4281 16188
rect 4319 16154 4353 16188
rect 4391 16154 4425 16188
rect 4463 16154 4497 16188
rect 4535 16154 4569 16188
rect 5089 16124 5123 16153
rect 5162 16124 5196 16153
rect 5235 16124 5269 16153
rect 5308 16124 5342 16153
rect 5381 16124 5415 16153
rect 5454 16124 5488 16153
rect 5527 16124 5561 16153
rect 5600 16124 5634 16153
rect 5673 16124 5707 16153
rect 5746 16124 5780 16153
rect 5819 16124 5853 16153
rect 5892 16124 5926 16153
rect 5965 16124 5999 16153
rect 6038 16124 6072 16153
rect 6110 16124 6144 16153
rect 6182 16124 6216 16153
rect 6254 16124 6288 16153
rect 6326 16124 6360 16153
rect 6398 16124 6432 16153
rect 6470 16124 6504 16153
rect 6542 16124 6576 16153
rect 6614 16124 6648 16153
rect 6686 16124 6720 16153
rect 6758 16124 6792 16153
rect 6830 16124 6864 16153
rect 6902 16124 6936 16153
rect 6974 16124 7008 16153
rect 7046 16124 7080 16153
rect 7118 16124 7152 16153
rect 2663 16081 2697 16115
rect 2735 16107 2769 16115
rect 2735 16081 2749 16107
rect 2749 16081 2769 16107
rect 2807 16081 2841 16115
rect 2879 16107 2913 16115
rect 2879 16081 2887 16107
rect 2887 16081 2913 16107
rect 2951 16081 2985 16115
rect 3023 16107 3057 16115
rect 3023 16081 3025 16107
rect 3025 16081 3057 16107
rect 3095 16081 3129 16115
rect 3167 16081 3201 16115
rect 3239 16107 3273 16115
rect 3239 16081 3267 16107
rect 3267 16081 3273 16107
rect 3311 16081 3345 16115
rect 3383 16107 3417 16115
rect 3383 16081 3405 16107
rect 3405 16081 3417 16107
rect 3455 16081 3489 16115
rect 3527 16107 3561 16115
rect 3527 16081 3543 16107
rect 3543 16081 3561 16107
rect 3599 16081 3633 16115
rect 3671 16107 3705 16115
rect 3671 16081 3681 16107
rect 3681 16081 3705 16107
rect 3743 16081 3777 16115
rect 3815 16107 3849 16115
rect 3815 16081 3819 16107
rect 3819 16081 3849 16107
rect 3887 16081 3921 16115
rect 3959 16107 3993 16115
rect 3959 16081 3991 16107
rect 3991 16081 3993 16107
rect 4031 16081 4065 16115
rect 4103 16107 4137 16115
rect 4103 16081 4129 16107
rect 4129 16081 4137 16107
rect 4175 16081 4209 16115
rect 4247 16107 4281 16115
rect 4247 16081 4267 16107
rect 4267 16081 4281 16107
rect 4319 16081 4353 16115
rect 4391 16107 4425 16115
rect 4391 16081 4405 16107
rect 4405 16081 4425 16107
rect 4463 16081 4497 16115
rect 4535 16107 4569 16115
rect 4535 16081 4543 16107
rect 4543 16081 4569 16107
rect 5089 16119 5119 16124
rect 5119 16119 5123 16124
rect 5162 16119 5188 16124
rect 5188 16119 5196 16124
rect 5235 16119 5257 16124
rect 5257 16119 5269 16124
rect 5308 16119 5326 16124
rect 5326 16119 5342 16124
rect 5381 16119 5395 16124
rect 5395 16119 5415 16124
rect 5454 16119 5464 16124
rect 5464 16119 5488 16124
rect 5527 16119 5533 16124
rect 5533 16119 5561 16124
rect 5600 16119 5602 16124
rect 5602 16119 5634 16124
rect 5673 16119 5706 16124
rect 5706 16119 5707 16124
rect 5746 16119 5775 16124
rect 5775 16119 5780 16124
rect 5819 16119 5844 16124
rect 5844 16119 5853 16124
rect 5892 16119 5913 16124
rect 5913 16119 5926 16124
rect 5965 16119 5982 16124
rect 5982 16119 5999 16124
rect 6038 16119 6051 16124
rect 6051 16119 6072 16124
rect 6110 16119 6120 16124
rect 6120 16119 6144 16124
rect 6182 16119 6189 16124
rect 6189 16119 6216 16124
rect 6254 16119 6258 16124
rect 6258 16119 6288 16124
rect 6326 16119 6327 16124
rect 6327 16119 6360 16124
rect 6398 16119 6430 16124
rect 6430 16119 6432 16124
rect 6470 16119 6499 16124
rect 6499 16119 6504 16124
rect 6542 16119 6568 16124
rect 6568 16119 6576 16124
rect 6614 16119 6637 16124
rect 6637 16119 6648 16124
rect 6686 16119 6706 16124
rect 6706 16119 6720 16124
rect 6758 16119 6775 16124
rect 6775 16119 6792 16124
rect 6830 16119 6844 16124
rect 6844 16119 6864 16124
rect 6902 16119 6913 16124
rect 6913 16119 6936 16124
rect 6974 16119 6982 16124
rect 6982 16119 7008 16124
rect 7046 16119 7051 16124
rect 7051 16119 7080 16124
rect 7118 16119 7120 16124
rect 7120 16119 7152 16124
rect 7190 16119 7224 16153
rect 7262 16124 7296 16153
rect 7334 16124 7368 16153
rect 7406 16124 7440 16153
rect 7478 16124 7512 16153
rect 7550 16124 7584 16153
rect 7622 16124 7656 16153
rect 7694 16124 7728 16153
rect 7766 16124 7800 16153
rect 7838 16124 7872 16153
rect 7262 16119 7293 16124
rect 7293 16119 7296 16124
rect 7334 16119 7362 16124
rect 7362 16119 7368 16124
rect 7406 16119 7431 16124
rect 7431 16119 7440 16124
rect 7478 16119 7500 16124
rect 7500 16119 7512 16124
rect 7550 16119 7568 16124
rect 7568 16119 7584 16124
rect 7622 16119 7636 16124
rect 7636 16119 7656 16124
rect 7694 16119 7704 16124
rect 7704 16119 7728 16124
rect 7766 16119 7772 16124
rect 7772 16119 7800 16124
rect 7838 16119 7840 16124
rect 7840 16119 7872 16124
rect 5089 16054 5123 16077
rect 5162 16054 5196 16077
rect 5235 16054 5269 16077
rect 5308 16054 5342 16077
rect 5381 16054 5415 16077
rect 5454 16054 5488 16077
rect 5527 16054 5561 16077
rect 5600 16054 5634 16077
rect 5673 16054 5707 16077
rect 5746 16054 5780 16077
rect 5819 16054 5853 16077
rect 5892 16054 5926 16077
rect 5965 16054 5999 16077
rect 6038 16054 6072 16077
rect 6110 16054 6144 16077
rect 6182 16054 6216 16077
rect 6254 16054 6288 16077
rect 6326 16054 6360 16077
rect 6398 16054 6432 16077
rect 6470 16054 6504 16077
rect 6542 16054 6576 16077
rect 6614 16054 6648 16077
rect 6686 16054 6720 16077
rect 6758 16054 6792 16077
rect 6830 16054 6864 16077
rect 6902 16054 6936 16077
rect 6974 16054 7008 16077
rect 7046 16054 7080 16077
rect 7118 16054 7152 16077
rect 2663 16008 2697 16042
rect 2735 16008 2769 16042
rect 2807 16008 2841 16042
rect 2879 16008 2913 16042
rect 2951 16008 2985 16042
rect 3023 16008 3057 16042
rect 3095 16008 3129 16042
rect 3167 16008 3201 16042
rect 3239 16008 3273 16042
rect 3311 16008 3345 16042
rect 3383 16008 3417 16042
rect 3455 16008 3489 16042
rect 3527 16008 3561 16042
rect 3599 16008 3633 16042
rect 3671 16008 3705 16042
rect 3743 16008 3777 16042
rect 3815 16008 3849 16042
rect 3887 16008 3921 16042
rect 3959 16008 3993 16042
rect 4031 16008 4065 16042
rect 4103 16008 4137 16042
rect 4175 16008 4209 16042
rect 4247 16008 4281 16042
rect 4319 16008 4353 16042
rect 4391 16008 4425 16042
rect 4463 16008 4497 16042
rect 4535 16008 4569 16042
rect 5089 16043 5119 16054
rect 5119 16043 5123 16054
rect 5162 16043 5188 16054
rect 5188 16043 5196 16054
rect 5235 16043 5257 16054
rect 5257 16043 5269 16054
rect 5308 16043 5326 16054
rect 5326 16043 5342 16054
rect 5381 16043 5395 16054
rect 5395 16043 5415 16054
rect 5454 16043 5464 16054
rect 5464 16043 5488 16054
rect 5527 16043 5533 16054
rect 5533 16043 5561 16054
rect 5600 16043 5602 16054
rect 5602 16043 5634 16054
rect 5673 16043 5706 16054
rect 5706 16043 5707 16054
rect 5746 16043 5775 16054
rect 5775 16043 5780 16054
rect 5819 16043 5844 16054
rect 5844 16043 5853 16054
rect 5892 16043 5913 16054
rect 5913 16043 5926 16054
rect 5965 16043 5982 16054
rect 5982 16043 5999 16054
rect 6038 16043 6051 16054
rect 6051 16043 6072 16054
rect 6110 16043 6120 16054
rect 6120 16043 6144 16054
rect 6182 16043 6189 16054
rect 6189 16043 6216 16054
rect 6254 16043 6258 16054
rect 6258 16043 6288 16054
rect 6326 16043 6327 16054
rect 6327 16043 6360 16054
rect 6398 16043 6430 16054
rect 6430 16043 6432 16054
rect 6470 16043 6499 16054
rect 6499 16043 6504 16054
rect 6542 16043 6568 16054
rect 6568 16043 6576 16054
rect 6614 16043 6637 16054
rect 6637 16043 6648 16054
rect 6686 16043 6706 16054
rect 6706 16043 6720 16054
rect 6758 16043 6775 16054
rect 6775 16043 6792 16054
rect 6830 16043 6844 16054
rect 6844 16043 6864 16054
rect 6902 16043 6913 16054
rect 6913 16043 6936 16054
rect 6974 16043 6982 16054
rect 6982 16043 7008 16054
rect 7046 16043 7051 16054
rect 7051 16043 7080 16054
rect 7118 16043 7120 16054
rect 7120 16043 7152 16054
rect 7190 16043 7224 16077
rect 7262 16054 7296 16077
rect 7334 16054 7368 16077
rect 7406 16054 7440 16077
rect 7478 16054 7512 16077
rect 7550 16054 7584 16077
rect 7622 16054 7656 16077
rect 7694 16054 7728 16077
rect 7766 16054 7800 16077
rect 7838 16054 7872 16077
rect 7262 16043 7293 16054
rect 7293 16043 7296 16054
rect 7334 16043 7362 16054
rect 7362 16043 7368 16054
rect 7406 16043 7431 16054
rect 7431 16043 7440 16054
rect 7478 16043 7500 16054
rect 7500 16043 7512 16054
rect 7550 16043 7568 16054
rect 7568 16043 7584 16054
rect 7622 16043 7636 16054
rect 7636 16043 7656 16054
rect 7694 16043 7704 16054
rect 7704 16043 7728 16054
rect 7766 16043 7772 16054
rect 7772 16043 7800 16054
rect 7838 16043 7840 16054
rect 7840 16043 7872 16054
rect 5089 15984 5123 16001
rect 5162 15984 5196 16001
rect 5235 15984 5269 16001
rect 5308 15984 5342 16001
rect 5381 15984 5415 16001
rect 5454 15984 5488 16001
rect 5527 15984 5561 16001
rect 5600 15984 5634 16001
rect 5673 15984 5707 16001
rect 5746 15984 5780 16001
rect 5819 15984 5853 16001
rect 5892 15984 5926 16001
rect 5965 15984 5999 16001
rect 6038 15984 6072 16001
rect 6110 15984 6144 16001
rect 6182 15984 6216 16001
rect 6254 15984 6288 16001
rect 6326 15984 6360 16001
rect 6398 15984 6432 16001
rect 6470 15984 6504 16001
rect 6542 15984 6576 16001
rect 6614 15984 6648 16001
rect 6686 15984 6720 16001
rect 6758 15984 6792 16001
rect 6830 15984 6864 16001
rect 6902 15984 6936 16001
rect 6974 15984 7008 16001
rect 7046 15984 7080 16001
rect 7118 15984 7152 16001
rect 2663 15935 2697 15969
rect 2735 15936 2749 15969
rect 2749 15936 2769 15969
rect 2735 15935 2769 15936
rect 2807 15935 2841 15969
rect 2879 15936 2887 15969
rect 2887 15936 2913 15969
rect 2879 15935 2913 15936
rect 2951 15935 2985 15969
rect 3023 15936 3025 15969
rect 3025 15936 3057 15969
rect 3023 15935 3057 15936
rect 3095 15935 3129 15969
rect 3167 15935 3201 15969
rect 3239 15936 3267 15969
rect 3267 15936 3273 15969
rect 3239 15935 3273 15936
rect 3311 15935 3345 15969
rect 3383 15936 3405 15969
rect 3405 15936 3417 15969
rect 3383 15935 3417 15936
rect 3455 15935 3489 15969
rect 3527 15936 3543 15969
rect 3543 15936 3561 15969
rect 3527 15935 3561 15936
rect 3599 15935 3633 15969
rect 3671 15936 3681 15969
rect 3681 15936 3705 15969
rect 3671 15935 3705 15936
rect 3743 15935 3777 15969
rect 3815 15936 3819 15969
rect 3819 15936 3849 15969
rect 3815 15935 3849 15936
rect 3887 15935 3921 15969
rect 3959 15936 3991 15969
rect 3991 15936 3993 15969
rect 3959 15935 3993 15936
rect 4031 15935 4065 15969
rect 4103 15936 4129 15969
rect 4129 15936 4137 15969
rect 4103 15935 4137 15936
rect 4175 15935 4209 15969
rect 4247 15936 4267 15969
rect 4267 15936 4281 15969
rect 4247 15935 4281 15936
rect 4319 15935 4353 15969
rect 4391 15936 4405 15969
rect 4405 15936 4425 15969
rect 4391 15935 4425 15936
rect 4463 15935 4497 15969
rect 4535 15936 4543 15969
rect 4543 15936 4569 15969
rect 5089 15967 5119 15984
rect 5119 15967 5123 15984
rect 5162 15967 5188 15984
rect 5188 15967 5196 15984
rect 5235 15967 5257 15984
rect 5257 15967 5269 15984
rect 5308 15967 5326 15984
rect 5326 15967 5342 15984
rect 5381 15967 5395 15984
rect 5395 15967 5415 15984
rect 5454 15967 5464 15984
rect 5464 15967 5488 15984
rect 5527 15967 5533 15984
rect 5533 15967 5561 15984
rect 5600 15967 5602 15984
rect 5602 15967 5634 15984
rect 5673 15967 5706 15984
rect 5706 15967 5707 15984
rect 5746 15967 5775 15984
rect 5775 15967 5780 15984
rect 5819 15967 5844 15984
rect 5844 15967 5853 15984
rect 5892 15967 5913 15984
rect 5913 15967 5926 15984
rect 5965 15967 5982 15984
rect 5982 15967 5999 15984
rect 6038 15967 6051 15984
rect 6051 15967 6072 15984
rect 6110 15967 6120 15984
rect 6120 15967 6144 15984
rect 6182 15967 6189 15984
rect 6189 15967 6216 15984
rect 6254 15967 6258 15984
rect 6258 15967 6288 15984
rect 6326 15967 6327 15984
rect 6327 15967 6360 15984
rect 6398 15967 6430 15984
rect 6430 15967 6432 15984
rect 6470 15967 6499 15984
rect 6499 15967 6504 15984
rect 6542 15967 6568 15984
rect 6568 15967 6576 15984
rect 6614 15967 6637 15984
rect 6637 15967 6648 15984
rect 6686 15967 6706 15984
rect 6706 15967 6720 15984
rect 6758 15967 6775 15984
rect 6775 15967 6792 15984
rect 6830 15967 6844 15984
rect 6844 15967 6864 15984
rect 6902 15967 6913 15984
rect 6913 15967 6936 15984
rect 6974 15967 6982 15984
rect 6982 15967 7008 15984
rect 7046 15967 7051 15984
rect 7051 15967 7080 15984
rect 7118 15967 7120 15984
rect 7120 15967 7152 15984
rect 7190 15967 7224 16001
rect 7262 15984 7296 16001
rect 7334 15984 7368 16001
rect 7406 15984 7440 16001
rect 7478 15984 7512 16001
rect 7550 15984 7584 16001
rect 7622 15984 7656 16001
rect 7694 15984 7728 16001
rect 7766 15984 7800 16001
rect 7838 15984 7872 16001
rect 7262 15967 7293 15984
rect 7293 15967 7296 15984
rect 7334 15967 7362 15984
rect 7362 15967 7368 15984
rect 7406 15967 7431 15984
rect 7431 15967 7440 15984
rect 7478 15967 7500 15984
rect 7500 15967 7512 15984
rect 7550 15967 7568 15984
rect 7568 15967 7584 15984
rect 7622 15967 7636 15984
rect 7636 15967 7656 15984
rect 7694 15967 7704 15984
rect 7704 15967 7728 15984
rect 7766 15967 7772 15984
rect 7772 15967 7800 15984
rect 7838 15967 7840 15984
rect 7840 15967 7872 15984
rect 4535 15935 4569 15936
rect 2276 15890 2310 15924
rect 2410 15890 2444 15924
rect 8050 17013 8084 17047
rect 8184 17003 8218 17037
rect 8050 16941 8084 16975
rect 8184 16931 8218 16965
rect 8050 16869 8084 16903
rect 8184 16859 8218 16893
rect 8050 16797 8084 16831
rect 8184 16787 8218 16821
rect 8050 16725 8084 16759
rect 8184 16715 8218 16749
rect 8050 16653 8084 16687
rect 8184 16643 8218 16677
rect 8050 16581 8084 16615
rect 8184 16571 8218 16605
rect 8050 16509 8084 16543
rect 8184 16499 8218 16533
rect 8050 16437 8084 16471
rect 8184 16427 8218 16461
rect 8050 16365 8084 16399
rect 8184 16355 8218 16389
rect 8050 16293 8084 16327
rect 8184 16283 8218 16317
rect 8050 16221 8084 16255
rect 8184 16211 8218 16245
rect 8050 16149 8084 16183
rect 8184 16139 8218 16173
rect 8050 16077 8084 16111
rect 8184 16067 8218 16101
rect 8050 16005 8084 16039
rect 8184 15995 8218 16029
rect 8050 15933 8084 15967
rect 8184 15923 8218 15957
rect 2276 15818 2310 15852
rect 2410 15818 2444 15852
rect 2276 15746 2310 15780
rect 2410 15746 2444 15780
rect 2276 15674 2310 15708
rect 2410 15674 2444 15708
rect 2276 15602 2310 15636
rect 2410 15602 2444 15636
rect 8050 15861 8084 15895
rect 8184 15851 8218 15885
rect 8050 15789 8084 15823
rect 8184 15779 8218 15813
rect 8050 15717 8084 15751
rect 8184 15707 8218 15741
rect 8050 15645 8084 15679
rect 8184 15635 8218 15669
rect 2276 15530 2310 15564
rect 2410 15530 2444 15564
rect 3035 15552 3039 15586
rect 3039 15552 3069 15586
rect 3108 15552 3142 15586
rect 3181 15552 3211 15586
rect 3211 15552 3215 15586
rect 3254 15552 3280 15586
rect 3280 15552 3288 15586
rect 3327 15552 3349 15586
rect 3349 15552 3361 15586
rect 3400 15552 3418 15586
rect 3418 15552 3434 15586
rect 3473 15552 3487 15586
rect 3487 15552 3507 15586
rect 3546 15552 3556 15586
rect 3556 15552 3580 15586
rect 3619 15552 3625 15586
rect 3625 15552 3653 15586
rect 3692 15552 3694 15586
rect 3694 15552 3726 15586
rect 3765 15552 3798 15586
rect 3798 15552 3799 15586
rect 3838 15552 3867 15586
rect 3867 15552 3872 15586
rect 3911 15552 3936 15586
rect 3936 15552 3945 15586
rect 3984 15552 4005 15586
rect 4005 15552 4018 15586
rect 4057 15552 4074 15586
rect 4074 15552 4091 15586
rect 4130 15552 4143 15586
rect 4143 15552 4164 15586
rect 4203 15552 4211 15586
rect 4211 15552 4237 15586
rect 4276 15552 4279 15586
rect 4279 15552 4310 15586
rect 4349 15552 4381 15586
rect 4381 15552 4383 15586
rect 4422 15552 4449 15586
rect 4449 15552 4456 15586
rect 4495 15552 4517 15586
rect 4517 15552 4529 15586
rect 4568 15552 4585 15586
rect 4585 15552 4602 15586
rect 4641 15552 4653 15586
rect 4653 15552 4675 15586
rect 4714 15552 4721 15586
rect 4721 15552 4748 15586
rect 4787 15552 4789 15586
rect 4789 15552 4821 15586
rect 4860 15552 4891 15586
rect 4891 15552 4894 15586
rect 4933 15552 4959 15586
rect 4959 15552 4967 15586
rect 5006 15552 5027 15586
rect 5027 15552 5040 15586
rect 5079 15552 5095 15586
rect 5095 15552 5113 15586
rect 5152 15552 5163 15586
rect 5163 15552 5186 15586
rect 5225 15552 5231 15586
rect 5231 15552 5259 15586
rect 5298 15552 5299 15586
rect 5299 15552 5332 15586
rect 5371 15552 5401 15586
rect 5401 15552 5405 15586
rect 5444 15552 5469 15586
rect 5469 15552 5478 15586
rect 5517 15552 5537 15586
rect 5537 15552 5551 15586
rect 5590 15552 5605 15586
rect 5605 15552 5624 15586
rect 5663 15552 5673 15586
rect 5673 15552 5697 15586
rect 5736 15552 5741 15586
rect 5741 15552 5770 15586
rect 5809 15552 5843 15586
rect 5881 15552 5911 15586
rect 5911 15552 5915 15586
rect 5953 15552 5979 15586
rect 5979 15552 5987 15586
rect 6025 15552 6047 15586
rect 6047 15552 6059 15586
rect 6097 15552 6115 15586
rect 6115 15552 6131 15586
rect 6169 15552 6183 15586
rect 6183 15552 6203 15586
rect 6241 15552 6251 15586
rect 6251 15552 6275 15586
rect 6313 15552 6319 15586
rect 6319 15552 6347 15586
rect 6385 15552 6387 15586
rect 6387 15552 6419 15586
rect 6457 15552 6489 15586
rect 6489 15552 6491 15586
rect 6529 15552 6557 15586
rect 6557 15552 6563 15586
rect 6601 15552 6625 15586
rect 6625 15552 6635 15586
rect 6673 15552 6693 15586
rect 6693 15552 6707 15586
rect 6745 15552 6761 15586
rect 6761 15552 6779 15586
rect 6817 15552 6829 15586
rect 6829 15552 6851 15586
rect 6889 15552 6897 15586
rect 6897 15552 6923 15586
rect 6961 15552 6965 15586
rect 6965 15552 6995 15586
rect 7033 15552 7067 15586
rect 7105 15552 7135 15586
rect 7135 15552 7139 15586
rect 7177 15552 7203 15586
rect 7203 15552 7211 15586
rect 7249 15552 7271 15586
rect 7271 15552 7283 15586
rect 7321 15552 7339 15586
rect 7339 15552 7355 15586
rect 7393 15552 7407 15586
rect 7407 15552 7427 15586
rect 7465 15552 7475 15586
rect 7475 15552 7499 15586
rect 7537 15552 7543 15586
rect 7543 15552 7571 15586
rect 7609 15552 7611 15586
rect 7611 15552 7643 15586
rect 7681 15552 7713 15586
rect 7713 15552 7715 15586
rect 8050 15573 8084 15607
rect 8184 15563 8218 15597
rect 2276 15458 2310 15492
rect 2410 15458 2444 15492
rect 8050 15501 8084 15535
rect 8184 15491 8218 15525
rect 2276 15386 2310 15420
rect 2410 15386 2444 15420
rect 2276 15314 2310 15348
rect 2410 15314 2444 15348
rect 2276 15242 2310 15276
rect 2410 15242 2444 15276
rect 2276 15170 2310 15204
rect 2410 15170 2444 15204
rect 2276 15098 2310 15132
rect 2410 15098 2444 15132
rect 2276 15026 2310 15060
rect 2410 15026 2444 15060
rect 2276 14954 2310 14988
rect 2410 14954 2444 14988
rect 2276 14882 2310 14916
rect 2410 14882 2444 14916
rect 2276 14810 2310 14844
rect 2410 14810 2444 14844
rect 2276 14738 2310 14772
rect 2410 14738 2444 14772
rect 2276 14666 2310 14700
rect 2410 14666 2444 14700
rect 2276 14594 2310 14628
rect 2410 14594 2444 14628
rect 2276 14522 2310 14556
rect 2410 14522 2444 14556
rect 2276 14450 2310 14484
rect 2410 14450 2444 14484
rect 2276 14378 2310 14412
rect 2410 14378 2444 14412
rect 2276 14306 2310 14340
rect 2410 14306 2444 14340
rect 2276 14234 2310 14268
rect 2410 14234 2444 14268
rect 2276 14162 2310 14196
rect 2410 14162 2444 14196
rect 2276 14090 2310 14124
rect 2410 14090 2444 14124
rect 2830 15412 2864 15446
rect 2902 15412 2936 15446
rect 2830 15339 2864 15373
rect 2902 15339 2936 15373
rect 2830 15266 2864 15300
rect 2902 15266 2936 15300
rect 2830 15193 2864 15227
rect 2902 15193 2936 15227
rect 2830 14112 2936 15154
rect 3107 15412 3141 15446
rect 3179 15412 3213 15446
rect 3107 15339 3141 15373
rect 3179 15339 3213 15373
rect 3107 15266 3141 15300
rect 3179 15266 3213 15300
rect 3107 15193 3141 15227
rect 3179 15193 3213 15227
rect 3107 14112 3213 15154
rect 3384 15412 3418 15446
rect 3456 15412 3490 15446
rect 3384 15339 3418 15373
rect 3456 15339 3490 15373
rect 3384 15266 3418 15300
rect 3456 15266 3490 15300
rect 3384 15193 3418 15227
rect 3456 15193 3490 15227
rect 3384 14112 3490 15154
rect 3661 15412 3695 15446
rect 3733 15412 3767 15446
rect 3661 15339 3695 15373
rect 3733 15339 3767 15373
rect 3661 15266 3695 15300
rect 3733 15266 3767 15300
rect 3661 15193 3695 15227
rect 3733 15193 3767 15227
rect 3661 14112 3767 15154
rect 3938 15412 3972 15446
rect 4010 15412 4044 15446
rect 3938 15339 3972 15373
rect 4010 15339 4044 15373
rect 3938 15266 3972 15300
rect 4010 15266 4044 15300
rect 3938 15193 3972 15227
rect 4010 15193 4044 15227
rect 3938 14112 4044 15154
rect 4215 15412 4249 15446
rect 4287 15412 4321 15446
rect 4215 15339 4249 15373
rect 4287 15339 4321 15373
rect 4215 15266 4249 15300
rect 4287 15266 4321 15300
rect 4215 15193 4249 15227
rect 4287 15193 4321 15227
rect 4215 14112 4321 15154
rect 4492 15412 4526 15446
rect 4564 15412 4598 15446
rect 4492 15339 4526 15373
rect 4564 15339 4598 15373
rect 4492 15266 4526 15300
rect 4564 15266 4598 15300
rect 4492 15193 4526 15227
rect 4564 15193 4598 15227
rect 4492 14112 4598 15154
rect 4769 15412 4803 15446
rect 4841 15412 4875 15446
rect 4769 15339 4803 15373
rect 4841 15339 4875 15373
rect 4769 15266 4803 15300
rect 4841 15266 4875 15300
rect 4769 15193 4803 15227
rect 4841 15193 4875 15227
rect 4769 14112 4875 15154
rect 5046 15412 5080 15446
rect 5118 15412 5152 15446
rect 5046 15339 5080 15373
rect 5118 15339 5152 15373
rect 5046 15266 5080 15300
rect 5118 15266 5152 15300
rect 5046 15193 5080 15227
rect 5118 15193 5152 15227
rect 5046 14112 5152 15154
rect 5323 15412 5357 15446
rect 5395 15412 5429 15446
rect 5323 15339 5357 15373
rect 5395 15339 5429 15373
rect 5323 15266 5357 15300
rect 5395 15266 5429 15300
rect 5323 15193 5357 15227
rect 5395 15193 5429 15227
rect 5323 14112 5429 15154
rect 5600 15412 5634 15446
rect 5672 15412 5706 15446
rect 5600 15339 5634 15373
rect 5672 15339 5706 15373
rect 5600 15266 5634 15300
rect 5672 15266 5706 15300
rect 5600 15193 5634 15227
rect 5672 15193 5706 15227
rect 5600 14112 5706 15154
rect 5877 15412 5911 15446
rect 5949 15412 5983 15446
rect 5877 15339 5911 15373
rect 5949 15339 5983 15373
rect 5877 15266 5911 15300
rect 5949 15266 5983 15300
rect 5877 15193 5911 15227
rect 5949 15193 5983 15227
rect 5877 14112 5983 15154
rect 6154 15412 6188 15446
rect 6226 15412 6260 15446
rect 6154 15339 6188 15373
rect 6226 15339 6260 15373
rect 6154 15266 6188 15300
rect 6226 15266 6260 15300
rect 6154 15193 6188 15227
rect 6226 15193 6260 15227
rect 6154 14112 6260 15154
rect 6431 15412 6465 15446
rect 6503 15412 6537 15446
rect 6431 15339 6465 15373
rect 6503 15339 6537 15373
rect 6431 15266 6465 15300
rect 6503 15266 6537 15300
rect 6431 15193 6465 15227
rect 6503 15193 6537 15227
rect 6431 14112 6537 15154
rect 6708 15412 6742 15446
rect 6780 15412 6814 15446
rect 6708 15339 6742 15373
rect 6780 15339 6814 15373
rect 6708 15266 6742 15300
rect 6780 15266 6814 15300
rect 6708 15193 6742 15227
rect 6780 15193 6814 15227
rect 6708 14112 6814 15154
rect 6985 15412 7019 15446
rect 7057 15412 7091 15446
rect 6985 15339 7019 15373
rect 7057 15339 7091 15373
rect 6985 15266 7019 15300
rect 7057 15266 7091 15300
rect 6985 15193 7019 15227
rect 7057 15193 7091 15227
rect 6985 14112 7091 15154
rect 7262 15412 7296 15446
rect 7334 15412 7368 15446
rect 7262 15339 7296 15373
rect 7334 15339 7368 15373
rect 7262 15266 7296 15300
rect 7334 15266 7368 15300
rect 7262 15193 7296 15227
rect 7334 15193 7368 15227
rect 7262 14112 7368 15154
rect 7539 15412 7573 15446
rect 7611 15412 7645 15446
rect 7539 15339 7573 15373
rect 7611 15339 7645 15373
rect 7539 15266 7573 15300
rect 7611 15266 7645 15300
rect 7539 15193 7573 15227
rect 7611 15193 7645 15227
rect 7539 14112 7645 15154
rect 7816 15412 7850 15446
rect 7888 15412 7922 15446
rect 7816 15339 7850 15373
rect 7888 15339 7922 15373
rect 7816 15266 7850 15300
rect 7888 15266 7922 15300
rect 7816 15193 7850 15227
rect 7888 15193 7922 15227
rect 7816 14112 7922 15154
rect 8050 15429 8084 15463
rect 8184 15419 8218 15453
rect 8050 15357 8084 15391
rect 8184 15347 8218 15381
rect 8050 15285 8084 15319
rect 8184 15275 8218 15309
rect 8050 15213 8084 15247
rect 8184 15203 8218 15237
rect 8050 15141 8084 15175
rect 8184 15131 8218 15165
rect 8050 15069 8084 15103
rect 8184 15059 8218 15093
rect 8050 14997 8084 15031
rect 8184 14987 8218 15021
rect 8050 14925 8084 14959
rect 8184 14915 8218 14949
rect 8050 14853 8084 14887
rect 8184 14843 8218 14877
rect 8050 14781 8084 14815
rect 8184 14771 8218 14805
rect 8050 14709 8084 14743
rect 8184 14699 8218 14733
rect 8050 14637 8084 14671
rect 8184 14627 8218 14661
rect 8050 14565 8084 14599
rect 8184 14555 8218 14589
rect 8050 14493 8084 14527
rect 8184 14483 8218 14517
rect 8050 14421 8084 14455
rect 8184 14411 8218 14445
rect 8050 14349 8084 14383
rect 8184 14339 8218 14373
rect 8050 14277 8084 14311
rect 8184 14267 8218 14301
rect 8050 14205 8084 14239
rect 8184 14195 8218 14229
rect 8050 14133 8084 14167
rect 8184 14123 8218 14157
rect 2276 14018 2310 14052
rect 2410 14018 2444 14052
rect 2276 13946 2310 13980
rect 2410 13946 2444 13980
rect 2276 13874 2310 13908
rect 2410 13874 2444 13908
rect 8050 14061 8084 14095
rect 8184 14051 8218 14085
rect 8050 13989 8084 14023
rect 8184 13979 8218 14013
rect 8050 13917 8084 13951
rect 8184 13907 8218 13941
rect 2276 13802 2310 13836
rect 2410 13802 2444 13836
rect 3035 13822 3039 13856
rect 3039 13822 3069 13856
rect 3108 13822 3142 13856
rect 3181 13822 3211 13856
rect 3211 13822 3215 13856
rect 3254 13822 3280 13856
rect 3280 13822 3288 13856
rect 3327 13822 3349 13856
rect 3349 13822 3361 13856
rect 3400 13822 3418 13856
rect 3418 13822 3434 13856
rect 3473 13822 3487 13856
rect 3487 13822 3507 13856
rect 3546 13822 3556 13856
rect 3556 13822 3580 13856
rect 3619 13822 3625 13856
rect 3625 13822 3653 13856
rect 3692 13822 3694 13856
rect 3694 13822 3726 13856
rect 3765 13822 3798 13856
rect 3798 13822 3799 13856
rect 3838 13822 3867 13856
rect 3867 13822 3872 13856
rect 3911 13822 3936 13856
rect 3936 13822 3945 13856
rect 3984 13822 4005 13856
rect 4005 13822 4018 13856
rect 4057 13822 4073 13856
rect 4073 13822 4091 13856
rect 4130 13822 4141 13856
rect 4141 13822 4164 13856
rect 4203 13822 4209 13856
rect 4209 13822 4237 13856
rect 4276 13822 4277 13856
rect 4277 13822 4310 13856
rect 4349 13822 4379 13856
rect 4379 13822 4383 13856
rect 4422 13822 4447 13856
rect 4447 13822 4456 13856
rect 4495 13822 4515 13856
rect 4515 13822 4529 13856
rect 4568 13822 4583 13856
rect 4583 13822 4602 13856
rect 4641 13822 4651 13856
rect 4651 13822 4675 13856
rect 4714 13822 4719 13856
rect 4719 13822 4748 13856
rect 4787 13822 4821 13856
rect 4860 13822 4889 13856
rect 4889 13822 4894 13856
rect 4933 13822 4957 13856
rect 4957 13822 4967 13856
rect 5006 13822 5025 13856
rect 5025 13822 5040 13856
rect 5079 13822 5093 13856
rect 5093 13822 5113 13856
rect 5152 13822 5161 13856
rect 5161 13822 5186 13856
rect 5225 13822 5229 13856
rect 5229 13822 5259 13856
rect 5298 13822 5331 13856
rect 5331 13822 5332 13856
rect 5371 13822 5399 13856
rect 5399 13822 5405 13856
rect 5444 13822 5467 13856
rect 5467 13822 5478 13856
rect 5517 13822 5535 13856
rect 5535 13822 5551 13856
rect 5590 13822 5603 13856
rect 5603 13822 5624 13856
rect 5663 13822 5671 13856
rect 5671 13822 5697 13856
rect 5736 13822 5739 13856
rect 5739 13822 5770 13856
rect 5809 13822 5841 13856
rect 5841 13822 5843 13856
rect 5881 13822 5909 13856
rect 5909 13822 5915 13856
rect 5953 13822 5977 13856
rect 5977 13822 5987 13856
rect 6025 13822 6045 13856
rect 6045 13822 6059 13856
rect 6097 13822 6113 13856
rect 6113 13822 6131 13856
rect 6169 13822 6181 13856
rect 6181 13822 6203 13856
rect 6241 13822 6249 13856
rect 6249 13822 6275 13856
rect 6313 13822 6317 13856
rect 6317 13822 6347 13856
rect 6385 13822 6419 13856
rect 6457 13822 6487 13856
rect 6487 13822 6491 13856
rect 6529 13822 6555 13856
rect 6555 13822 6563 13856
rect 6601 13822 6623 13856
rect 6623 13822 6635 13856
rect 6673 13822 6691 13856
rect 6691 13822 6707 13856
rect 6745 13822 6759 13856
rect 6759 13822 6779 13856
rect 6817 13822 6827 13856
rect 6827 13822 6851 13856
rect 6889 13822 6895 13856
rect 6895 13822 6923 13856
rect 6961 13822 6963 13856
rect 6963 13822 6995 13856
rect 7033 13822 7065 13856
rect 7065 13822 7067 13856
rect 7105 13822 7133 13856
rect 7133 13822 7139 13856
rect 7177 13822 7201 13856
rect 7201 13822 7211 13856
rect 7249 13822 7269 13856
rect 7269 13822 7283 13856
rect 7321 13822 7337 13856
rect 7337 13822 7355 13856
rect 7393 13822 7405 13856
rect 7405 13822 7427 13856
rect 7465 13822 7473 13856
rect 7473 13822 7499 13856
rect 7537 13822 7541 13856
rect 7541 13822 7571 13856
rect 7609 13822 7643 13856
rect 7681 13822 7711 13856
rect 7711 13822 7715 13856
rect 8050 13845 8084 13879
rect 8184 13835 8218 13869
rect 2276 13730 2310 13764
rect 2410 13730 2444 13764
rect 2276 13658 2310 13692
rect 2410 13658 2444 13692
rect 2276 13586 2310 13620
rect 2410 13586 2444 13620
rect 2276 13514 2310 13548
rect 2410 13514 2444 13548
rect 2276 13442 2310 13476
rect 2410 13442 2444 13476
rect 8050 13773 8084 13807
rect 8184 13763 8218 13797
rect 8050 13701 8084 13735
rect 8184 13691 8218 13725
rect 8050 13629 8084 13663
rect 8184 13619 8218 13653
rect 8050 13557 8084 13591
rect 8184 13547 8218 13581
rect 8050 13485 8084 13519
rect 8184 13475 8218 13509
rect 2276 13370 2310 13404
rect 2410 13370 2444 13404
rect 2276 13298 2310 13332
rect 2410 13298 2444 13332
rect 2276 13226 2310 13260
rect 2410 13226 2444 13260
rect 2276 13154 2310 13188
rect 2410 13154 2444 13188
rect 2276 13082 2310 13116
rect 2410 13082 2444 13116
rect 2276 13010 2310 13044
rect 2410 13010 2444 13044
rect 2276 12938 2310 12972
rect 2410 12938 2444 12972
rect 2276 12866 2310 12900
rect 2410 12866 2444 12900
rect 2276 12794 2310 12828
rect 2410 12794 2444 12828
rect 2276 12722 2310 12756
rect 2410 12722 2444 12756
rect 2276 12650 2310 12684
rect 2410 12650 2444 12684
rect 2276 12578 2310 12612
rect 2410 12578 2444 12612
rect 2276 12506 2310 12540
rect 2410 12506 2444 12540
rect 2276 12434 2310 12468
rect 2410 12434 2444 12468
rect 2276 12362 2310 12396
rect 2410 12362 2444 12396
rect 2276 12290 2310 12324
rect 2410 12290 2444 12324
rect 2276 12218 2310 12252
rect 2410 12218 2444 12252
rect 2276 12146 2310 12180
rect 2410 12146 2444 12180
rect 2830 13412 2864 13446
rect 2902 13412 2936 13446
rect 2830 13339 2864 13373
rect 2902 13339 2936 13373
rect 2830 13266 2864 13300
rect 2902 13266 2936 13300
rect 2830 13193 2864 13227
rect 2902 13193 2936 13227
rect 2830 12112 2936 13154
rect 3107 13412 3141 13446
rect 3179 13412 3213 13446
rect 3107 13339 3141 13373
rect 3179 13339 3213 13373
rect 3107 13266 3141 13300
rect 3179 13266 3213 13300
rect 3107 13193 3141 13227
rect 3179 13193 3213 13227
rect 3107 12112 3213 13154
rect 3384 13412 3418 13446
rect 3456 13412 3490 13446
rect 3384 13339 3418 13373
rect 3456 13339 3490 13373
rect 3384 13266 3418 13300
rect 3456 13266 3490 13300
rect 3384 13193 3418 13227
rect 3456 13193 3490 13227
rect 3384 12112 3490 13154
rect 3661 13412 3695 13446
rect 3733 13412 3767 13446
rect 3661 13339 3695 13373
rect 3733 13339 3767 13373
rect 3661 13266 3695 13300
rect 3733 13266 3767 13300
rect 3661 13193 3695 13227
rect 3733 13193 3767 13227
rect 3661 12112 3767 13154
rect 3938 13412 3972 13446
rect 4010 13412 4044 13446
rect 3938 13339 3972 13373
rect 4010 13339 4044 13373
rect 3938 13266 3972 13300
rect 4010 13266 4044 13300
rect 3938 13193 3972 13227
rect 4010 13193 4044 13227
rect 3938 12112 4044 13154
rect 4215 13412 4249 13446
rect 4287 13412 4321 13446
rect 4215 13339 4249 13373
rect 4287 13339 4321 13373
rect 4215 13266 4249 13300
rect 4287 13266 4321 13300
rect 4215 13193 4249 13227
rect 4287 13193 4321 13227
rect 4215 12112 4321 13154
rect 4492 13412 4526 13446
rect 4564 13412 4598 13446
rect 4492 13339 4526 13373
rect 4564 13339 4598 13373
rect 4492 13266 4526 13300
rect 4564 13266 4598 13300
rect 4492 13193 4526 13227
rect 4564 13193 4598 13227
rect 4492 12112 4598 13154
rect 4769 13412 4803 13446
rect 4841 13412 4875 13446
rect 4769 13339 4803 13373
rect 4841 13339 4875 13373
rect 4769 13266 4803 13300
rect 4841 13266 4875 13300
rect 4769 13193 4803 13227
rect 4841 13193 4875 13227
rect 4769 12112 4875 13154
rect 5046 13412 5080 13446
rect 5118 13412 5152 13446
rect 5046 13339 5080 13373
rect 5118 13339 5152 13373
rect 5046 13266 5080 13300
rect 5118 13266 5152 13300
rect 5046 13193 5080 13227
rect 5118 13193 5152 13227
rect 5046 12112 5152 13154
rect 5323 13412 5357 13446
rect 5395 13412 5429 13446
rect 5323 13339 5357 13373
rect 5395 13339 5429 13373
rect 5323 13266 5357 13300
rect 5395 13266 5429 13300
rect 5323 13193 5357 13227
rect 5395 13193 5429 13227
rect 5323 12112 5429 13154
rect 5600 13412 5634 13446
rect 5672 13412 5706 13446
rect 5600 13339 5634 13373
rect 5672 13339 5706 13373
rect 5600 13266 5634 13300
rect 5672 13266 5706 13300
rect 5600 13193 5634 13227
rect 5672 13193 5706 13227
rect 5600 12112 5706 13154
rect 5877 13412 5911 13446
rect 5949 13412 5983 13446
rect 5877 13339 5911 13373
rect 5949 13339 5983 13373
rect 5877 13266 5911 13300
rect 5949 13266 5983 13300
rect 5877 13193 5911 13227
rect 5949 13193 5983 13227
rect 5877 12112 5983 13154
rect 6154 13412 6188 13446
rect 6226 13412 6260 13446
rect 6154 13339 6188 13373
rect 6226 13339 6260 13373
rect 6154 13266 6188 13300
rect 6226 13266 6260 13300
rect 6154 13193 6188 13227
rect 6226 13193 6260 13227
rect 6154 12112 6260 13154
rect 6431 13412 6465 13446
rect 6503 13412 6537 13446
rect 6431 13339 6465 13373
rect 6503 13339 6537 13373
rect 6431 13266 6465 13300
rect 6503 13266 6537 13300
rect 6431 13193 6465 13227
rect 6503 13193 6537 13227
rect 6431 12112 6537 13154
rect 6708 13412 6742 13446
rect 6780 13412 6814 13446
rect 6708 13339 6742 13373
rect 6780 13339 6814 13373
rect 6708 13266 6742 13300
rect 6780 13266 6814 13300
rect 6708 13193 6742 13227
rect 6780 13193 6814 13227
rect 6708 12112 6814 13154
rect 6985 13412 7019 13446
rect 7057 13412 7091 13446
rect 6985 13339 7019 13373
rect 7057 13339 7091 13373
rect 6985 13266 7019 13300
rect 7057 13266 7091 13300
rect 6985 13193 7019 13227
rect 7057 13193 7091 13227
rect 6985 12112 7091 13154
rect 7262 13412 7296 13446
rect 7334 13412 7368 13446
rect 7262 13339 7296 13373
rect 7334 13339 7368 13373
rect 7262 13266 7296 13300
rect 7334 13266 7368 13300
rect 7262 13193 7296 13227
rect 7334 13193 7368 13227
rect 7262 12112 7368 13154
rect 7539 13412 7573 13446
rect 7611 13412 7645 13446
rect 7539 13339 7573 13373
rect 7611 13339 7645 13373
rect 7539 13266 7573 13300
rect 7611 13266 7645 13300
rect 7539 13193 7573 13227
rect 7611 13193 7645 13227
rect 7539 12112 7645 13154
rect 7816 13412 7850 13446
rect 7888 13412 7922 13446
rect 7816 13339 7850 13373
rect 7888 13339 7922 13373
rect 7816 13266 7850 13300
rect 7888 13266 7922 13300
rect 7816 13193 7850 13227
rect 7888 13193 7922 13227
rect 7816 12112 7922 13154
rect 8050 13413 8084 13447
rect 8184 13403 8218 13437
rect 8050 13341 8084 13375
rect 8184 13331 8218 13365
rect 8050 13269 8084 13303
rect 8184 13259 8218 13293
rect 8050 13197 8084 13231
rect 8184 13187 8218 13221
rect 8050 13125 8084 13159
rect 8184 13115 8218 13149
rect 8050 13053 8084 13087
rect 8184 13043 8218 13077
rect 8050 12981 8084 13015
rect 8184 12971 8218 13005
rect 8050 12908 8084 12942
rect 8184 12899 8218 12933
rect 8050 12835 8084 12869
rect 8184 12827 8218 12861
rect 8050 12762 8084 12796
rect 8184 12755 8218 12789
rect 8050 12689 8084 12723
rect 8184 12683 8218 12717
rect 8050 12616 8084 12650
rect 8184 12611 8218 12645
rect 8050 12543 8084 12577
rect 8184 12539 8218 12573
rect 8050 12470 8084 12504
rect 8184 12467 8218 12501
rect 8050 12397 8084 12431
rect 8184 12395 8218 12429
rect 8050 12324 8084 12358
rect 8184 12323 8218 12357
rect 8050 12251 8084 12285
rect 8184 12251 8218 12285
rect 8050 12178 8084 12212
rect 8184 12178 8218 12212
rect 2276 12074 2310 12108
rect 2410 12074 2444 12108
rect 8050 12105 8084 12139
rect 8184 12105 8218 12139
rect 2276 12002 2310 12036
rect 2410 12002 2444 12036
rect 2276 11930 2310 11964
rect 2410 11930 2444 11964
rect 2276 11858 2310 11892
rect 2410 11858 2444 11892
rect 2276 11786 2310 11820
rect 2410 11786 2444 11820
rect 8050 12032 8084 12066
rect 8184 12032 8218 12066
rect 8050 11959 8084 11993
rect 8184 11959 8218 11993
rect 8050 11886 8084 11920
rect 8184 11886 8218 11920
rect 3035 11784 3039 11818
rect 3039 11784 3069 11818
rect 3108 11784 3142 11818
rect 3181 11784 3211 11818
rect 3211 11784 3215 11818
rect 3254 11784 3280 11818
rect 3280 11784 3288 11818
rect 3327 11784 3349 11818
rect 3349 11784 3361 11818
rect 3400 11784 3418 11818
rect 3418 11784 3434 11818
rect 3473 11784 3487 11818
rect 3487 11784 3507 11818
rect 3546 11784 3556 11818
rect 3556 11784 3580 11818
rect 3619 11784 3625 11818
rect 3625 11784 3653 11818
rect 3692 11784 3694 11818
rect 3694 11784 3726 11818
rect 3765 11784 3798 11818
rect 3798 11784 3799 11818
rect 3838 11784 3867 11818
rect 3867 11784 3872 11818
rect 3911 11784 3936 11818
rect 3936 11784 3945 11818
rect 3984 11784 4005 11818
rect 4005 11784 4018 11818
rect 4057 11784 4073 11818
rect 4073 11784 4091 11818
rect 4130 11784 4141 11818
rect 4141 11784 4164 11818
rect 4203 11784 4209 11818
rect 4209 11784 4237 11818
rect 4276 11784 4277 11818
rect 4277 11784 4310 11818
rect 4349 11784 4379 11818
rect 4379 11784 4383 11818
rect 4422 11784 4447 11818
rect 4447 11784 4456 11818
rect 4495 11784 4515 11818
rect 4515 11784 4529 11818
rect 4568 11784 4583 11818
rect 4583 11784 4602 11818
rect 4641 11784 4651 11818
rect 4651 11784 4675 11818
rect 4714 11784 4719 11818
rect 4719 11784 4748 11818
rect 4787 11784 4821 11818
rect 4860 11784 4889 11818
rect 4889 11784 4894 11818
rect 4933 11784 4957 11818
rect 4957 11784 4967 11818
rect 5006 11784 5025 11818
rect 5025 11784 5040 11818
rect 5079 11784 5093 11818
rect 5093 11784 5113 11818
rect 5152 11784 5161 11818
rect 5161 11784 5186 11818
rect 5225 11784 5229 11818
rect 5229 11784 5259 11818
rect 5298 11784 5331 11818
rect 5331 11784 5332 11818
rect 5371 11784 5399 11818
rect 5399 11784 5405 11818
rect 5444 11784 5467 11818
rect 5467 11784 5478 11818
rect 5517 11784 5535 11818
rect 5535 11784 5551 11818
rect 5590 11784 5603 11818
rect 5603 11784 5624 11818
rect 5663 11784 5671 11818
rect 5671 11784 5697 11818
rect 5736 11784 5739 11818
rect 5739 11784 5770 11818
rect 5809 11784 5841 11818
rect 5841 11784 5843 11818
rect 5881 11784 5909 11818
rect 5909 11784 5915 11818
rect 5953 11784 5977 11818
rect 5977 11784 5987 11818
rect 6025 11784 6045 11818
rect 6045 11784 6059 11818
rect 6097 11784 6113 11818
rect 6113 11784 6131 11818
rect 6169 11784 6181 11818
rect 6181 11784 6203 11818
rect 6241 11784 6249 11818
rect 6249 11784 6275 11818
rect 6313 11784 6317 11818
rect 6317 11784 6347 11818
rect 6385 11784 6419 11818
rect 6457 11784 6487 11818
rect 6487 11784 6491 11818
rect 6529 11784 6555 11818
rect 6555 11784 6563 11818
rect 6601 11784 6623 11818
rect 6623 11784 6635 11818
rect 6673 11784 6691 11818
rect 6691 11784 6707 11818
rect 6745 11784 6759 11818
rect 6759 11784 6779 11818
rect 6817 11784 6827 11818
rect 6827 11784 6851 11818
rect 6889 11784 6895 11818
rect 6895 11784 6923 11818
rect 6961 11784 6963 11818
rect 6963 11784 6995 11818
rect 7033 11784 7065 11818
rect 7065 11784 7067 11818
rect 7105 11784 7133 11818
rect 7133 11784 7139 11818
rect 7177 11784 7201 11818
rect 7201 11784 7211 11818
rect 7249 11784 7269 11818
rect 7269 11784 7283 11818
rect 7321 11784 7337 11818
rect 7337 11784 7355 11818
rect 7393 11784 7405 11818
rect 7405 11784 7427 11818
rect 7465 11784 7473 11818
rect 7473 11784 7499 11818
rect 7537 11784 7541 11818
rect 7541 11784 7571 11818
rect 7609 11784 7643 11818
rect 7681 11784 7711 11818
rect 7711 11784 7715 11818
rect 8050 11813 8084 11847
rect 8184 11813 8218 11847
rect 2276 11714 2310 11748
rect 2410 11714 2444 11748
rect 2276 11642 2310 11676
rect 2410 11642 2444 11676
rect 2276 11570 2310 11604
rect 2410 11570 2444 11604
rect 2276 11498 2310 11532
rect 2410 11498 2444 11532
rect 2276 11426 2310 11460
rect 2410 11426 2444 11460
rect 8050 11740 8084 11774
rect 8184 11740 8218 11774
rect 8050 11667 8084 11701
rect 8184 11667 8218 11701
rect 8050 11594 8084 11628
rect 8184 11594 8218 11628
rect 8050 11521 8084 11555
rect 8184 11521 8218 11555
rect 8050 11448 8084 11482
rect 8184 11448 8218 11482
rect 2276 11354 2310 11388
rect 2410 11354 2444 11388
rect 2276 11282 2310 11316
rect 2410 11282 2444 11316
rect 2276 11210 2310 11244
rect 2410 11210 2444 11244
rect 2276 11138 2310 11172
rect 2410 11138 2444 11172
rect 2276 11066 2310 11100
rect 2410 11066 2444 11100
rect 2276 10994 2310 11028
rect 2410 10994 2444 11028
rect 2276 10922 2310 10956
rect 2410 10922 2444 10956
rect 2276 10850 2310 10884
rect 2410 10850 2444 10884
rect 2276 10778 2310 10812
rect 2410 10778 2444 10812
rect 2276 10706 2310 10740
rect 2410 10706 2444 10740
rect 2276 10634 2310 10668
rect 2410 10634 2444 10668
rect 2276 10562 2310 10596
rect 2410 10562 2444 10596
rect 2276 10490 2310 10524
rect 2410 10490 2444 10524
rect 2276 10418 2310 10452
rect 2410 10418 2444 10452
rect 2276 10346 2310 10380
rect 2410 10346 2444 10380
rect 2276 10274 2310 10308
rect 2410 10274 2444 10308
rect 2276 10202 2310 10236
rect 2410 10202 2444 10236
rect 2276 10130 2310 10164
rect 2410 10130 2444 10164
rect 2830 11412 2864 11446
rect 2902 11412 2936 11446
rect 2830 11339 2864 11373
rect 2902 11339 2936 11373
rect 2830 11266 2864 11300
rect 2902 11266 2936 11300
rect 2830 11193 2864 11227
rect 2902 11193 2936 11227
rect 2830 10112 2936 11154
rect 3107 11412 3141 11446
rect 3179 11412 3213 11446
rect 3107 11339 3141 11373
rect 3179 11339 3213 11373
rect 3107 11266 3141 11300
rect 3179 11266 3213 11300
rect 3107 11193 3141 11227
rect 3179 11193 3213 11227
rect 3107 10112 3213 11154
rect 3384 11412 3418 11446
rect 3456 11412 3490 11446
rect 3384 11339 3418 11373
rect 3456 11339 3490 11373
rect 3384 11266 3418 11300
rect 3456 11266 3490 11300
rect 3384 11193 3418 11227
rect 3456 11193 3490 11227
rect 3384 10112 3490 11154
rect 3661 11412 3695 11446
rect 3733 11412 3767 11446
rect 3661 11339 3695 11373
rect 3733 11339 3767 11373
rect 3661 11266 3695 11300
rect 3733 11266 3767 11300
rect 3661 11193 3695 11227
rect 3733 11193 3767 11227
rect 3661 10112 3767 11154
rect 3938 11412 3972 11446
rect 4010 11412 4044 11446
rect 3938 11339 3972 11373
rect 4010 11339 4044 11373
rect 3938 11266 3972 11300
rect 4010 11266 4044 11300
rect 3938 11193 3972 11227
rect 4010 11193 4044 11227
rect 3938 10112 4044 11154
rect 4215 11412 4249 11446
rect 4287 11412 4321 11446
rect 4215 11339 4249 11373
rect 4287 11339 4321 11373
rect 4215 11266 4249 11300
rect 4287 11266 4321 11300
rect 4215 11193 4249 11227
rect 4287 11193 4321 11227
rect 4215 10112 4321 11154
rect 4492 11412 4526 11446
rect 4564 11412 4598 11446
rect 4492 11339 4526 11373
rect 4564 11339 4598 11373
rect 4492 11266 4526 11300
rect 4564 11266 4598 11300
rect 4492 11193 4526 11227
rect 4564 11193 4598 11227
rect 4492 10112 4598 11154
rect 4769 11412 4803 11446
rect 4841 11412 4875 11446
rect 4769 11339 4803 11373
rect 4841 11339 4875 11373
rect 4769 11266 4803 11300
rect 4841 11266 4875 11300
rect 4769 11193 4803 11227
rect 4841 11193 4875 11227
rect 4769 10112 4875 11154
rect 5046 11412 5080 11446
rect 5118 11412 5152 11446
rect 5046 11339 5080 11373
rect 5118 11339 5152 11373
rect 5046 11266 5080 11300
rect 5118 11266 5152 11300
rect 5046 11193 5080 11227
rect 5118 11193 5152 11227
rect 5046 10112 5152 11154
rect 5323 11412 5357 11446
rect 5395 11412 5429 11446
rect 5323 11339 5357 11373
rect 5395 11339 5429 11373
rect 5323 11266 5357 11300
rect 5395 11266 5429 11300
rect 5323 11193 5357 11227
rect 5395 11193 5429 11227
rect 5323 10112 5429 11154
rect 5600 11412 5634 11446
rect 5672 11412 5706 11446
rect 5600 11339 5634 11373
rect 5672 11339 5706 11373
rect 5600 11266 5634 11300
rect 5672 11266 5706 11300
rect 5600 11193 5634 11227
rect 5672 11193 5706 11227
rect 5600 10112 5706 11154
rect 5877 11412 5911 11446
rect 5949 11412 5983 11446
rect 5877 11339 5911 11373
rect 5949 11339 5983 11373
rect 5877 11266 5911 11300
rect 5949 11266 5983 11300
rect 5877 11193 5911 11227
rect 5949 11193 5983 11227
rect 5877 10112 5983 11154
rect 6154 11412 6188 11446
rect 6226 11412 6260 11446
rect 6154 11339 6188 11373
rect 6226 11339 6260 11373
rect 6154 11266 6188 11300
rect 6226 11266 6260 11300
rect 6154 11193 6188 11227
rect 6226 11193 6260 11227
rect 6154 10112 6260 11154
rect 6431 11412 6465 11446
rect 6503 11412 6537 11446
rect 6431 11339 6465 11373
rect 6503 11339 6537 11373
rect 6431 11266 6465 11300
rect 6503 11266 6537 11300
rect 6431 11193 6465 11227
rect 6503 11193 6537 11227
rect 6431 10112 6537 11154
rect 6708 11412 6742 11446
rect 6780 11412 6814 11446
rect 6708 11339 6742 11373
rect 6780 11339 6814 11373
rect 6708 11266 6742 11300
rect 6780 11266 6814 11300
rect 6708 11193 6742 11227
rect 6780 11193 6814 11227
rect 6708 10112 6814 11154
rect 6985 11412 7019 11446
rect 7057 11412 7091 11446
rect 6985 11339 7019 11373
rect 7057 11339 7091 11373
rect 6985 11266 7019 11300
rect 7057 11266 7091 11300
rect 6985 11193 7019 11227
rect 7057 11193 7091 11227
rect 6985 10112 7091 11154
rect 7262 11412 7296 11446
rect 7334 11412 7368 11446
rect 7262 11339 7296 11373
rect 7334 11339 7368 11373
rect 7262 11266 7296 11300
rect 7334 11266 7368 11300
rect 7262 11193 7296 11227
rect 7334 11193 7368 11227
rect 7262 10112 7368 11154
rect 7539 11412 7573 11446
rect 7611 11412 7645 11446
rect 7539 11339 7573 11373
rect 7611 11339 7645 11373
rect 7539 11266 7573 11300
rect 7611 11266 7645 11300
rect 7539 11193 7573 11227
rect 7611 11193 7645 11227
rect 7539 10112 7645 11154
rect 7816 11412 7850 11446
rect 7888 11412 7922 11446
rect 7816 11339 7850 11373
rect 7888 11339 7922 11373
rect 7816 11266 7850 11300
rect 7888 11266 7922 11300
rect 7816 11193 7850 11227
rect 7888 11193 7922 11227
rect 7816 10112 7922 11154
rect 8050 11375 8084 11409
rect 8184 11375 8218 11409
rect 8050 11302 8084 11336
rect 8184 11302 8218 11336
rect 8050 11229 8084 11263
rect 8184 11229 8218 11263
rect 8050 11156 8084 11190
rect 8184 11156 8218 11190
rect 8050 11083 8084 11117
rect 8184 11083 8218 11117
rect 8050 11010 8084 11044
rect 8184 11010 8218 11044
rect 8050 10937 8084 10971
rect 8184 10937 8218 10971
rect 8050 10864 8084 10898
rect 8184 10864 8218 10898
rect 8050 10791 8084 10825
rect 8184 10791 8218 10825
rect 8050 10718 8084 10752
rect 8184 10718 8218 10752
rect 8050 10645 8084 10679
rect 8184 10645 8218 10679
rect 8050 10572 8084 10606
rect 8184 10572 8218 10606
rect 8050 10499 8084 10533
rect 8184 10499 8218 10533
rect 8050 10426 8084 10460
rect 8184 10426 8218 10460
rect 8050 10353 8084 10387
rect 8184 10353 8218 10387
rect 8050 10280 8084 10314
rect 8184 10280 8218 10314
rect 8050 10207 8084 10241
rect 8184 10207 8218 10241
rect 8050 10134 8084 10168
rect 8184 10134 8218 10168
rect 2276 10058 2310 10092
rect 2410 10058 2444 10092
rect 8050 10061 8084 10095
rect 8184 10061 8218 10095
rect 3035 10022 3039 10050
rect 3039 10022 3069 10050
rect 3108 10022 3142 10050
rect 3181 10022 3211 10050
rect 3211 10022 3215 10050
rect 3254 10022 3280 10050
rect 3280 10022 3288 10050
rect 3327 10022 3349 10050
rect 3349 10022 3361 10050
rect 3400 10022 3418 10050
rect 3418 10022 3434 10050
rect 3473 10022 3487 10050
rect 3487 10022 3507 10050
rect 3546 10022 3556 10050
rect 3556 10022 3580 10050
rect 3619 10022 3625 10050
rect 3625 10022 3653 10050
rect 3692 10022 3694 10050
rect 3694 10022 3726 10050
rect 3765 10022 3798 10050
rect 3798 10022 3799 10050
rect 3838 10022 3867 10050
rect 3867 10022 3872 10050
rect 3911 10022 3936 10050
rect 3936 10022 3945 10050
rect 3984 10022 4005 10050
rect 4005 10022 4018 10050
rect 4057 10022 4074 10050
rect 4074 10022 4091 10050
rect 4130 10022 4143 10050
rect 4143 10022 4164 10050
rect 4203 10022 4211 10050
rect 4211 10022 4237 10050
rect 4276 10022 4279 10050
rect 4279 10022 4310 10050
rect 4349 10022 4381 10050
rect 4381 10022 4383 10050
rect 4422 10022 4449 10050
rect 4449 10022 4456 10050
rect 4495 10022 4517 10050
rect 4517 10022 4529 10050
rect 4568 10022 4585 10050
rect 4585 10022 4602 10050
rect 4641 10022 4653 10050
rect 4653 10022 4675 10050
rect 4714 10022 4721 10050
rect 4721 10022 4748 10050
rect 4787 10022 4789 10050
rect 4789 10022 4821 10050
rect 4860 10022 4891 10050
rect 4891 10022 4894 10050
rect 4933 10022 4959 10050
rect 4959 10022 4967 10050
rect 5006 10022 5027 10050
rect 5027 10022 5040 10050
rect 5079 10022 5095 10050
rect 5095 10022 5113 10050
rect 5152 10022 5163 10050
rect 5163 10022 5186 10050
rect 5225 10022 5231 10050
rect 5231 10022 5259 10050
rect 5298 10022 5299 10050
rect 5299 10022 5332 10050
rect 5371 10022 5401 10050
rect 5401 10022 5405 10050
rect 5444 10022 5469 10050
rect 5469 10022 5478 10050
rect 5517 10022 5537 10050
rect 5537 10022 5551 10050
rect 5590 10022 5605 10050
rect 5605 10022 5624 10050
rect 5663 10022 5673 10050
rect 5673 10022 5697 10050
rect 5736 10022 5741 10050
rect 5741 10022 5770 10050
rect 2276 10004 2310 10020
rect 2410 10004 2444 10020
rect 3035 10016 3069 10022
rect 3108 10016 3142 10022
rect 3181 10016 3215 10022
rect 3254 10016 3288 10022
rect 3327 10016 3361 10022
rect 3400 10016 3434 10022
rect 3473 10016 3507 10022
rect 3546 10016 3580 10022
rect 3619 10016 3653 10022
rect 3692 10016 3726 10022
rect 3765 10016 3799 10022
rect 3838 10016 3872 10022
rect 3911 10016 3945 10022
rect 3984 10016 4018 10022
rect 4057 10016 4091 10022
rect 4130 10016 4164 10022
rect 4203 10016 4237 10022
rect 4276 10016 4310 10022
rect 4349 10016 4383 10022
rect 4422 10016 4456 10022
rect 4495 10016 4529 10022
rect 4568 10016 4602 10022
rect 4641 10016 4675 10022
rect 4714 10016 4748 10022
rect 4787 10016 4821 10022
rect 4860 10016 4894 10022
rect 4933 10016 4967 10022
rect 5006 10016 5040 10022
rect 5079 10016 5113 10022
rect 5152 10016 5186 10022
rect 5225 10016 5259 10022
rect 5298 10016 5332 10022
rect 5371 10016 5405 10022
rect 5444 10016 5478 10022
rect 5517 10016 5551 10022
rect 5590 10016 5624 10022
rect 5663 10016 5697 10022
rect 5736 10016 5770 10022
rect 5809 10016 5843 10050
rect 5882 10022 5911 10050
rect 5911 10022 5916 10050
rect 5955 10022 5979 10050
rect 5979 10022 5989 10050
rect 6027 10022 6047 10050
rect 6047 10022 6061 10050
rect 6099 10022 6115 10050
rect 6115 10022 6133 10050
rect 6171 10022 6183 10050
rect 6183 10022 6205 10050
rect 6243 10022 6251 10050
rect 6251 10022 6277 10050
rect 6315 10022 6319 10050
rect 6319 10022 6349 10050
rect 6387 10022 6421 10050
rect 6459 10022 6489 10050
rect 6489 10022 6493 10050
rect 6531 10022 6557 10050
rect 6557 10022 6565 10050
rect 6603 10022 6625 10050
rect 6625 10022 6637 10050
rect 6675 10022 6693 10050
rect 6693 10022 6709 10050
rect 6747 10022 6761 10050
rect 6761 10022 6781 10050
rect 6819 10022 6829 10050
rect 6829 10022 6853 10050
rect 6891 10022 6897 10050
rect 6897 10022 6925 10050
rect 6963 10022 6965 10050
rect 6965 10022 6997 10050
rect 7035 10022 7067 10050
rect 7067 10022 7069 10050
rect 7107 10022 7135 10050
rect 7135 10022 7141 10050
rect 7179 10022 7203 10050
rect 7203 10022 7213 10050
rect 7251 10022 7271 10050
rect 7271 10022 7285 10050
rect 7323 10022 7339 10050
rect 7339 10022 7357 10050
rect 7395 10022 7407 10050
rect 7407 10022 7429 10050
rect 7467 10022 7475 10050
rect 7475 10022 7501 10050
rect 7539 10022 7543 10050
rect 7543 10022 7573 10050
rect 7611 10022 7645 10050
rect 7683 10022 7713 10050
rect 7713 10022 7717 10050
rect 5882 10016 5916 10022
rect 5955 10016 5989 10022
rect 6027 10016 6061 10022
rect 6099 10016 6133 10022
rect 6171 10016 6205 10022
rect 6243 10016 6277 10022
rect 6315 10016 6349 10022
rect 6387 10016 6421 10022
rect 6459 10016 6493 10022
rect 6531 10016 6565 10022
rect 6603 10016 6637 10022
rect 6675 10016 6709 10022
rect 6747 10016 6781 10022
rect 6819 10016 6853 10022
rect 6891 10016 6925 10022
rect 6963 10016 6997 10022
rect 7035 10016 7069 10022
rect 7107 10016 7141 10022
rect 7179 10016 7213 10022
rect 7251 10016 7285 10022
rect 7323 10016 7357 10022
rect 7395 10016 7429 10022
rect 7467 10016 7501 10022
rect 7539 10016 7573 10022
rect 7611 10016 7645 10022
rect 7683 10016 7717 10022
rect 2276 9986 2310 10004
rect 2410 9986 2444 10004
rect 2276 9919 2310 9948
rect 2410 9919 2444 9948
rect 8050 9988 8084 10022
rect 8184 9988 8218 10022
rect 2276 9914 2298 9919
rect 2298 9914 2310 9919
rect 2410 9914 2436 9919
rect 2436 9914 2444 9919
rect 8050 9915 8084 9949
rect 8184 9915 8195 9949
rect 8195 9915 8218 9949
rect 2276 9842 2310 9876
rect 2410 9842 2444 9876
rect 2482 9836 2516 9870
rect 2555 9836 2589 9870
rect 2628 9836 2662 9870
rect 2701 9836 2735 9870
rect 2774 9836 2808 9870
rect 2847 9836 2881 9870
rect 2920 9836 2954 9870
rect 2993 9836 3027 9870
rect 3066 9836 3100 9870
rect 3139 9836 3173 9870
rect 3212 9836 3246 9870
rect 3285 9836 3319 9870
rect 3358 9836 3392 9870
rect 3431 9836 3465 9870
rect 3504 9836 3538 9870
rect 3577 9836 3611 9870
rect 3650 9836 3684 9870
rect 3723 9836 3757 9870
rect 3796 9836 3830 9870
rect 3869 9836 3903 9870
rect 3942 9836 3976 9870
rect 4015 9836 4049 9870
rect 4088 9836 4122 9870
rect 4161 9836 4195 9870
rect 4234 9836 4268 9870
rect 4306 9836 4340 9870
rect 4378 9836 4412 9870
rect 4450 9836 4484 9870
rect 4522 9836 4556 9870
rect 4594 9836 4628 9870
rect 4666 9836 4700 9870
rect 4738 9836 4772 9870
rect 4810 9836 4844 9870
rect 4882 9836 4916 9870
rect 4954 9836 4988 9870
rect 5026 9836 5060 9870
rect 5098 9836 5132 9870
rect 5170 9836 5204 9870
rect 5242 9836 5276 9870
rect 5314 9836 5348 9870
rect 5386 9836 5420 9870
rect 5458 9836 5492 9870
rect 5530 9836 5564 9870
rect 5602 9836 5636 9870
rect 5674 9836 5708 9870
rect 5746 9836 5780 9870
rect 5818 9836 5852 9870
rect 5890 9836 5924 9870
rect 5962 9836 5996 9870
rect 6034 9836 6068 9870
rect 6106 9836 6140 9870
rect 6178 9836 6212 9870
rect 6250 9836 6284 9870
rect 6322 9836 6356 9870
rect 6394 9836 6428 9870
rect 6466 9836 6500 9870
rect 6538 9836 6572 9870
rect 6610 9836 6644 9870
rect 6682 9836 6716 9870
rect 6754 9836 6788 9870
rect 6826 9836 6860 9870
rect 6898 9836 6932 9870
rect 6970 9836 7004 9870
rect 7042 9836 7076 9870
rect 7114 9836 7148 9870
rect 7186 9836 7220 9870
rect 7258 9836 7292 9870
rect 7330 9836 7364 9870
rect 7402 9836 7436 9870
rect 7474 9836 7508 9870
rect 7546 9836 7580 9870
rect 7618 9836 7652 9870
rect 7690 9836 7724 9870
rect 7762 9836 7796 9870
rect 7834 9836 7868 9870
rect 7906 9836 7940 9870
rect 7978 9836 8012 9870
rect 8050 9842 8084 9876
rect 8184 9842 8218 9876
rect 8429 14530 8431 39286
rect 8431 14530 8533 39286
rect 8533 14530 8535 39286
rect 8429 14457 8431 14491
rect 8431 14457 8463 14491
rect 8501 14457 8533 14491
rect 8533 14457 8535 14491
rect 8429 14384 8431 14418
rect 8431 14384 8463 14418
rect 8501 14384 8533 14418
rect 8533 14384 8535 14418
rect 8429 14311 8431 14345
rect 8431 14311 8463 14345
rect 8501 14311 8533 14345
rect 8533 14311 8535 14345
rect 8429 14238 8431 14272
rect 8431 14238 8463 14272
rect 8501 14238 8533 14272
rect 8533 14238 8535 14272
rect 8429 14165 8431 14199
rect 8431 14165 8463 14199
rect 8501 14165 8533 14199
rect 8533 14165 8535 14199
rect 8429 14092 8431 14126
rect 8431 14092 8463 14126
rect 8501 14092 8533 14126
rect 8533 14092 8535 14126
rect 8429 14019 8431 14053
rect 8431 14019 8463 14053
rect 8501 14019 8533 14053
rect 8533 14019 8535 14053
rect 8429 13946 8431 13980
rect 8431 13946 8463 13980
rect 8501 13946 8533 13980
rect 8533 13946 8535 13980
rect 8429 13873 8431 13907
rect 8431 13873 8463 13907
rect 8501 13873 8533 13907
rect 8533 13873 8535 13907
rect 8429 13800 8431 13834
rect 8431 13800 8463 13834
rect 8501 13800 8533 13834
rect 8533 13800 8535 13834
rect 8429 13727 8431 13761
rect 8431 13727 8463 13761
rect 8501 13727 8533 13761
rect 8533 13727 8535 13761
rect 8429 13654 8431 13688
rect 8431 13654 8463 13688
rect 8501 13654 8533 13688
rect 8533 13654 8535 13688
rect 8429 13581 8431 13615
rect 8431 13581 8463 13615
rect 8501 13581 8533 13615
rect 8533 13581 8535 13615
rect 8429 13508 8431 13542
rect 8431 13508 8463 13542
rect 8501 13508 8533 13542
rect 8533 13508 8535 13542
rect 8429 13435 8431 13469
rect 8431 13435 8463 13469
rect 8501 13435 8533 13469
rect 8533 13435 8535 13469
rect 8429 13362 8431 13396
rect 8431 13362 8463 13396
rect 8501 13362 8533 13396
rect 8533 13362 8535 13396
rect 8429 13289 8431 13323
rect 8431 13289 8463 13323
rect 8501 13289 8533 13323
rect 8533 13289 8535 13323
rect 8429 13216 8431 13250
rect 8431 13216 8463 13250
rect 8501 13216 8533 13250
rect 8533 13216 8535 13250
rect 8429 13143 8431 13177
rect 8431 13143 8463 13177
rect 8501 13143 8533 13177
rect 8533 13143 8535 13177
rect 8429 13070 8431 13104
rect 8431 13070 8463 13104
rect 8501 13070 8533 13104
rect 8533 13070 8535 13104
rect 8429 12997 8431 13031
rect 8431 12997 8463 13031
rect 8501 12997 8533 13031
rect 8533 12997 8535 13031
rect 8429 12924 8431 12958
rect 8431 12924 8463 12958
rect 8501 12924 8533 12958
rect 8533 12924 8535 12958
rect 8429 12851 8431 12885
rect 8431 12851 8463 12885
rect 8501 12851 8533 12885
rect 8533 12851 8535 12885
rect 8429 12778 8431 12812
rect 8431 12778 8463 12812
rect 8501 12778 8533 12812
rect 8533 12778 8535 12812
rect 8429 12705 8431 12739
rect 8431 12705 8463 12739
rect 8501 12705 8533 12739
rect 8533 12705 8535 12739
rect 8429 12632 8431 12666
rect 8431 12632 8463 12666
rect 8501 12632 8533 12666
rect 8533 12632 8535 12666
rect 8429 12559 8431 12593
rect 8431 12559 8463 12593
rect 8501 12559 8533 12593
rect 8533 12559 8535 12593
rect 8429 12486 8431 12520
rect 8431 12486 8463 12520
rect 8501 12486 8533 12520
rect 8533 12486 8535 12520
rect 8429 12413 8431 12447
rect 8431 12413 8463 12447
rect 8501 12413 8533 12447
rect 8533 12413 8535 12447
rect 8429 12340 8431 12374
rect 8431 12340 8463 12374
rect 8501 12340 8533 12374
rect 8533 12340 8535 12374
rect 8429 12267 8431 12301
rect 8431 12267 8463 12301
rect 8501 12267 8533 12301
rect 8533 12267 8535 12301
rect 8429 12194 8431 12228
rect 8431 12194 8463 12228
rect 8501 12194 8533 12228
rect 8533 12194 8535 12228
rect 8429 12121 8431 12155
rect 8431 12121 8463 12155
rect 8501 12121 8533 12155
rect 8533 12121 8535 12155
rect 8429 12048 8431 12082
rect 8431 12048 8463 12082
rect 8501 12048 8533 12082
rect 8533 12048 8535 12082
rect 8429 11975 8431 12009
rect 8431 11975 8463 12009
rect 8501 11975 8533 12009
rect 8533 11975 8535 12009
rect 8429 11902 8431 11936
rect 8431 11902 8463 11936
rect 8501 11902 8533 11936
rect 8533 11902 8535 11936
rect 8429 11829 8431 11863
rect 8431 11829 8463 11863
rect 8501 11829 8533 11863
rect 8533 11829 8535 11863
rect 8429 11756 8431 11790
rect 8431 11756 8463 11790
rect 8501 11756 8533 11790
rect 8533 11756 8535 11790
rect 8429 11683 8431 11717
rect 8431 11683 8463 11717
rect 8501 11683 8533 11717
rect 8533 11683 8535 11717
rect 8429 11610 8431 11644
rect 8431 11610 8463 11644
rect 8501 11610 8533 11644
rect 8533 11610 8535 11644
rect 8429 11537 8431 11571
rect 8431 11537 8463 11571
rect 8501 11537 8533 11571
rect 8533 11537 8535 11571
rect 8429 11464 8431 11498
rect 8431 11464 8463 11498
rect 8501 11464 8533 11498
rect 8533 11464 8535 11498
rect 8429 11391 8431 11425
rect 8431 11391 8463 11425
rect 8501 11391 8533 11425
rect 8533 11391 8535 11425
rect 8429 11318 8431 11352
rect 8431 11318 8463 11352
rect 8501 11318 8533 11352
rect 8533 11318 8535 11352
rect 8429 11245 8431 11279
rect 8431 11245 8463 11279
rect 8501 11245 8533 11279
rect 8533 11245 8535 11279
rect 8429 11172 8431 11206
rect 8431 11172 8463 11206
rect 8501 11172 8533 11206
rect 8533 11172 8535 11206
rect 8429 11099 8431 11133
rect 8431 11099 8463 11133
rect 8501 11099 8533 11133
rect 8533 11099 8535 11133
rect 8429 11026 8431 11060
rect 8431 11026 8463 11060
rect 8501 11026 8533 11060
rect 8533 11026 8535 11060
rect 8429 10953 8431 10987
rect 8431 10953 8463 10987
rect 8501 10953 8533 10987
rect 8533 10953 8535 10987
rect 8429 10880 8431 10914
rect 8431 10880 8463 10914
rect 8501 10880 8533 10914
rect 8533 10880 8535 10914
rect 8429 10807 8431 10841
rect 8431 10807 8463 10841
rect 8501 10807 8533 10841
rect 8533 10807 8535 10841
rect 8429 10734 8431 10768
rect 8431 10734 8463 10768
rect 8501 10734 8533 10768
rect 8533 10734 8535 10768
rect 8429 10661 8431 10695
rect 8431 10661 8463 10695
rect 8501 10661 8533 10695
rect 8533 10661 8535 10695
rect 8429 10588 8431 10622
rect 8431 10588 8463 10622
rect 8501 10588 8533 10622
rect 8533 10588 8535 10622
rect 8429 10515 8431 10549
rect 8431 10515 8463 10549
rect 8501 10515 8533 10549
rect 8533 10515 8535 10549
rect 8429 10442 8431 10476
rect 8431 10442 8463 10476
rect 8501 10442 8533 10476
rect 8533 10442 8535 10476
rect 8429 10369 8431 10403
rect 8431 10369 8463 10403
rect 8501 10369 8533 10403
rect 8533 10369 8535 10403
rect 8429 10296 8431 10330
rect 8431 10296 8463 10330
rect 8501 10296 8533 10330
rect 8533 10296 8535 10330
rect 8429 10223 8431 10257
rect 8431 10223 8463 10257
rect 8501 10223 8533 10257
rect 8533 10223 8535 10257
rect 8429 10150 8431 10184
rect 8431 10150 8463 10184
rect 8501 10150 8533 10184
rect 8533 10150 8535 10184
rect 8429 10077 8431 10111
rect 8431 10077 8463 10111
rect 8501 10077 8533 10111
rect 8533 10077 8535 10111
rect 8429 10004 8431 10038
rect 8431 10004 8463 10038
rect 8501 10004 8533 10038
rect 8533 10004 8535 10038
rect 8429 9931 8431 9965
rect 8431 9931 8463 9965
rect 8501 9931 8533 9965
rect 8533 9931 8535 9965
rect 8429 9858 8431 9892
rect 8431 9858 8463 9892
rect 8501 9858 8533 9892
rect 8533 9858 8535 9892
rect 8429 9785 8431 9819
rect 8431 9785 8463 9819
rect 8501 9785 8533 9819
rect 8533 9785 8535 9819
rect 7805 9712 7839 9746
rect 7883 9712 7917 9746
rect 7961 9712 7995 9746
rect 8039 9712 8073 9746
rect 8116 9712 8150 9746
rect 8193 9712 8227 9746
rect 8270 9712 8304 9746
rect 8347 9712 8381 9746
rect 8429 9712 8431 9746
rect 8431 9712 8463 9746
rect 8501 9712 8533 9746
rect 8533 9712 8535 9746
rect 2048 9593 2122 9699
rect 2161 9665 2195 9699
rect 2234 9697 2268 9699
rect 2307 9697 2341 9699
rect 2380 9697 2414 9699
rect 2453 9697 2487 9699
rect 2526 9697 2560 9699
rect 2599 9697 2633 9699
rect 2672 9697 2706 9699
rect 2745 9697 2779 9699
rect 2818 9697 2852 9699
rect 2891 9697 2925 9699
rect 2964 9697 2998 9699
rect 3037 9697 3071 9699
rect 3110 9697 3144 9699
rect 3183 9697 3217 9699
rect 3256 9697 3290 9699
rect 3329 9697 3363 9699
rect 3402 9697 3436 9699
rect 3475 9697 3509 9699
rect 3548 9697 3582 9699
rect 3621 9697 3655 9699
rect 3694 9697 3728 9699
rect 3767 9697 3801 9699
rect 3840 9697 3874 9699
rect 3913 9697 3947 9699
rect 3986 9697 4020 9699
rect 4059 9697 4093 9699
rect 4132 9697 4166 9699
rect 4205 9697 7695 9699
rect 2234 9665 2268 9697
rect 2307 9665 2341 9697
rect 2380 9665 2414 9697
rect 2453 9665 2487 9697
rect 2526 9665 2560 9697
rect 2599 9665 2633 9697
rect 2672 9665 2706 9697
rect 2745 9665 2779 9697
rect 2818 9665 2852 9697
rect 2891 9665 2925 9697
rect 2964 9665 2998 9697
rect 3037 9665 3071 9697
rect 3110 9665 3144 9697
rect 3183 9665 3217 9697
rect 3256 9665 3290 9697
rect 3329 9665 3363 9697
rect 3402 9665 3436 9697
rect 3475 9665 3509 9697
rect 3548 9665 3582 9697
rect 3621 9665 3655 9697
rect 3694 9665 3728 9697
rect 3767 9665 3801 9697
rect 3840 9665 3874 9697
rect 3913 9665 3947 9697
rect 3986 9665 4020 9697
rect 4059 9665 4093 9697
rect 4132 9665 4166 9697
rect 2161 9593 2195 9627
rect 2234 9595 2268 9627
rect 2307 9595 2341 9627
rect 2380 9595 2414 9627
rect 2453 9595 2487 9627
rect 2526 9595 2560 9627
rect 2599 9595 2633 9627
rect 2672 9595 2706 9627
rect 2745 9595 2779 9627
rect 2818 9595 2852 9627
rect 2891 9595 2925 9627
rect 2964 9595 2998 9627
rect 3037 9595 3071 9627
rect 3110 9595 3144 9627
rect 3183 9595 3217 9627
rect 3256 9595 3290 9627
rect 3329 9595 3363 9627
rect 3402 9595 3436 9627
rect 3475 9595 3509 9627
rect 3548 9595 3582 9627
rect 3621 9595 3655 9627
rect 3694 9595 3728 9627
rect 3767 9595 3801 9627
rect 3840 9595 3874 9627
rect 3913 9595 3947 9627
rect 3986 9595 4020 9627
rect 4059 9595 4093 9627
rect 4132 9595 4166 9627
rect 4205 9595 7546 9697
rect 7546 9674 7695 9697
rect 7546 9638 7839 9674
rect 7883 9640 7917 9674
rect 7961 9640 7995 9674
rect 8039 9640 8073 9674
rect 8116 9640 8150 9674
rect 8193 9640 8227 9674
rect 8270 9640 8304 9674
rect 8347 9640 8381 9674
rect 8424 9640 8431 9674
rect 8431 9640 8458 9674
rect 7546 9595 7803 9638
rect 2234 9593 2268 9595
rect 2307 9593 2341 9595
rect 2380 9593 2414 9595
rect 2453 9593 2487 9595
rect 2526 9593 2560 9595
rect 2599 9593 2633 9595
rect 2672 9593 2706 9595
rect 2745 9593 2779 9595
rect 2818 9593 2852 9595
rect 2891 9593 2925 9595
rect 2964 9593 2998 9595
rect 3037 9593 3071 9595
rect 3110 9593 3144 9595
rect 3183 9593 3217 9595
rect 3256 9593 3290 9595
rect 3329 9593 3363 9595
rect 3402 9593 3436 9595
rect 3475 9593 3509 9595
rect 3548 9593 3582 9595
rect 3621 9593 3655 9595
rect 3694 9593 3728 9595
rect 3767 9593 3801 9595
rect 3840 9593 3874 9595
rect 3913 9593 3947 9595
rect 3986 9593 4020 9595
rect 4059 9593 4093 9595
rect 4132 9593 4166 9595
rect 4205 9593 7803 9595
rect 2048 8938 2050 9593
rect 7733 9536 7803 9593
rect 7803 9536 7839 9638
rect 7733 9513 7839 9536
rect 7733 9479 7735 9513
rect 7735 9479 7769 9513
rect 7769 9479 7839 9513
rect 1944 8840 1946 8874
rect 1946 8840 1978 8874
rect 2016 8840 2048 8874
rect 2048 8840 2050 8874
rect 1944 8767 1946 8801
rect 1946 8767 1978 8801
rect 2016 8767 2048 8801
rect 2048 8767 2050 8801
rect 1944 8694 1946 8728
rect 1946 8694 1978 8728
rect 2016 8694 2048 8728
rect 2048 8694 2050 8728
rect 1944 8621 1946 8655
rect 1946 8621 1978 8655
rect 2016 8621 2048 8655
rect 2048 8621 2050 8655
rect 1944 8548 1946 8582
rect 1946 8548 1978 8582
rect 2016 8548 2048 8582
rect 2048 8548 2050 8582
rect 1944 8475 1946 8509
rect 1946 8475 1978 8509
rect 2016 8475 2048 8509
rect 2048 8475 2050 8509
rect 1944 8402 1946 8436
rect 1946 8402 1978 8436
rect 2016 8402 2048 8436
rect 2048 8402 2050 8436
rect 1944 8329 1946 8363
rect 1946 8329 1978 8363
rect 2016 8329 2048 8363
rect 2048 8329 2050 8363
rect 1944 8256 1946 8290
rect 1946 8256 1978 8290
rect 2016 8256 2048 8290
rect 2048 8256 2050 8290
rect 1944 8183 1946 8217
rect 1946 8183 1978 8217
rect 2016 8183 2048 8217
rect 2048 8183 2050 8217
rect 1944 8110 1946 8144
rect 1946 8110 1978 8144
rect 2016 8110 2048 8144
rect 2048 8110 2050 8144
rect 1944 8037 1946 8071
rect 1946 8037 1978 8071
rect 2016 8037 2048 8071
rect 2048 8037 2050 8071
rect 1944 7964 1946 7998
rect 1946 7964 1978 7998
rect 2016 7964 2048 7998
rect 2048 7964 2050 7998
rect 1944 7891 1946 7925
rect 1946 7891 1978 7925
rect 2016 7891 2048 7925
rect 2048 7891 2050 7925
rect 1944 7818 1946 7852
rect 1946 7818 1978 7852
rect 2016 7818 2048 7852
rect 2048 7818 2050 7852
rect 1944 7745 1946 7779
rect 1946 7745 1978 7779
rect 2016 7745 2048 7779
rect 2048 7745 2050 7779
rect 1944 7672 1946 7706
rect 1946 7672 1978 7706
rect 2016 7672 2048 7706
rect 2048 7672 2050 7706
rect 1944 7599 1946 7633
rect 1946 7599 1978 7633
rect 2016 7599 2048 7633
rect 2048 7599 2050 7633
rect 1944 7526 1946 7560
rect 1946 7526 1978 7560
rect 2016 7526 2048 7560
rect 2048 7526 2050 7560
rect 1944 7453 1946 7487
rect 1946 7453 1978 7487
rect 2016 7453 2048 7487
rect 2048 7453 2050 7487
rect 1944 7380 1946 7414
rect 1946 7380 1978 7414
rect 2016 7380 2048 7414
rect 2048 7380 2050 7414
rect 1944 4080 1946 7341
rect 1946 4080 2048 7341
rect 2048 4080 2050 7341
rect 1944 3927 2050 4080
rect 1944 3491 1946 3927
rect 1946 3491 2048 3927
rect 2048 3491 2050 3927
rect 2141 9430 2319 9443
rect 2359 9430 2393 9449
rect 2432 9430 2466 9449
rect 2505 9430 2539 9449
rect 2578 9430 2612 9449
rect 2651 9430 2685 9449
rect 2724 9430 2758 9449
rect 2797 9430 2831 9449
rect 2870 9430 2904 9449
rect 2943 9430 2977 9449
rect 3016 9430 3050 9449
rect 3089 9430 3123 9449
rect 3162 9430 3196 9449
rect 3235 9430 3269 9449
rect 3308 9430 3342 9449
rect 3381 9430 3415 9449
rect 3454 9430 3488 9449
rect 3527 9430 3561 9449
rect 3600 9430 3634 9449
rect 3673 9430 3707 9449
rect 3746 9430 3780 9449
rect 3819 9430 3853 9449
rect 3892 9430 3926 9449
rect 3965 9430 3999 9449
rect 4038 9430 4072 9449
rect 4111 9430 4145 9449
rect 2141 9396 2304 9430
rect 2304 9396 2319 9430
rect 2359 9415 2373 9430
rect 2373 9415 2393 9430
rect 2432 9415 2442 9430
rect 2442 9415 2466 9430
rect 2505 9415 2511 9430
rect 2511 9415 2539 9430
rect 2578 9415 2580 9430
rect 2580 9415 2612 9430
rect 2651 9415 2683 9430
rect 2683 9415 2685 9430
rect 2724 9415 2752 9430
rect 2752 9415 2758 9430
rect 2797 9415 2821 9430
rect 2821 9415 2831 9430
rect 2870 9415 2890 9430
rect 2890 9415 2904 9430
rect 2943 9415 2959 9430
rect 2959 9415 2977 9430
rect 3016 9415 3028 9430
rect 3028 9415 3050 9430
rect 3089 9415 3096 9430
rect 3096 9415 3123 9430
rect 3162 9415 3164 9430
rect 3164 9415 3196 9430
rect 3235 9415 3266 9430
rect 3266 9415 3269 9430
rect 3308 9415 3334 9430
rect 3334 9415 3342 9430
rect 3381 9415 3402 9430
rect 3402 9415 3415 9430
rect 3454 9415 3470 9430
rect 3470 9415 3488 9430
rect 3527 9415 3538 9430
rect 3538 9415 3561 9430
rect 3600 9415 3606 9430
rect 3606 9415 3634 9430
rect 3673 9415 3674 9430
rect 3674 9415 3707 9430
rect 3746 9415 3776 9430
rect 3776 9415 3780 9430
rect 3819 9415 3844 9430
rect 3844 9415 3853 9430
rect 3892 9415 3912 9430
rect 3912 9415 3926 9430
rect 3965 9415 3980 9430
rect 3980 9415 3999 9430
rect 4038 9415 4048 9430
rect 4048 9415 4072 9430
rect 4111 9415 4116 9430
rect 4116 9415 4145 9430
rect 4184 9415 4218 9449
rect 4257 9430 4291 9449
rect 4330 9430 4364 9449
rect 4403 9430 4437 9449
rect 4476 9430 4510 9449
rect 4549 9430 4583 9449
rect 4622 9430 4656 9449
rect 4694 9430 4728 9449
rect 4766 9430 4800 9449
rect 4838 9430 4872 9449
rect 4910 9430 4944 9449
rect 4982 9430 5016 9449
rect 5054 9430 5088 9449
rect 5126 9430 5160 9449
rect 5198 9430 5232 9449
rect 5270 9430 5304 9449
rect 5342 9430 5376 9449
rect 5414 9430 5448 9449
rect 5486 9430 5520 9449
rect 5558 9430 5592 9449
rect 5630 9430 5664 9449
rect 5702 9430 5736 9449
rect 5774 9430 5808 9449
rect 5846 9430 5880 9449
rect 5918 9430 5952 9449
rect 5990 9430 6024 9449
rect 6062 9430 6096 9449
rect 6134 9430 6168 9449
rect 6206 9430 6240 9449
rect 6278 9430 6312 9449
rect 6350 9430 6384 9449
rect 6422 9430 6456 9449
rect 6494 9430 6528 9449
rect 6566 9430 6600 9449
rect 6638 9430 6672 9449
rect 6710 9430 6744 9449
rect 6782 9430 6816 9449
rect 6854 9430 6888 9449
rect 6926 9430 6960 9449
rect 6998 9430 7032 9449
rect 7070 9430 7104 9449
rect 7142 9430 7176 9449
rect 7214 9430 7248 9449
rect 7286 9430 7320 9449
rect 7358 9430 7392 9449
rect 4257 9415 4286 9430
rect 4286 9415 4291 9430
rect 4330 9415 4354 9430
rect 4354 9415 4364 9430
rect 4403 9415 4422 9430
rect 4422 9415 4437 9430
rect 4476 9415 4490 9430
rect 4490 9415 4510 9430
rect 4549 9415 4558 9430
rect 4558 9415 4583 9430
rect 4622 9415 4626 9430
rect 4626 9415 4656 9430
rect 4694 9415 4728 9430
rect 4766 9415 4796 9430
rect 4796 9415 4800 9430
rect 4838 9415 4864 9430
rect 4864 9415 4872 9430
rect 4910 9415 4932 9430
rect 4932 9415 4944 9430
rect 4982 9415 5000 9430
rect 5000 9415 5016 9430
rect 5054 9415 5068 9430
rect 5068 9415 5088 9430
rect 5126 9415 5136 9430
rect 5136 9415 5160 9430
rect 5198 9415 5204 9430
rect 5204 9415 5232 9430
rect 5270 9415 5272 9430
rect 5272 9415 5304 9430
rect 5342 9415 5374 9430
rect 5374 9415 5376 9430
rect 5414 9415 5442 9430
rect 5442 9415 5448 9430
rect 5486 9415 5510 9430
rect 5510 9415 5520 9430
rect 5558 9415 5578 9430
rect 5578 9415 5592 9430
rect 5630 9415 5646 9430
rect 5646 9415 5664 9430
rect 5702 9415 5714 9430
rect 5714 9415 5736 9430
rect 5774 9415 5782 9430
rect 5782 9415 5808 9430
rect 5846 9415 5850 9430
rect 5850 9415 5880 9430
rect 5918 9415 5952 9430
rect 5990 9415 6020 9430
rect 6020 9415 6024 9430
rect 6062 9415 6088 9430
rect 6088 9415 6096 9430
rect 6134 9415 6156 9430
rect 6156 9415 6168 9430
rect 6206 9415 6224 9430
rect 6224 9415 6240 9430
rect 6278 9415 6292 9430
rect 6292 9415 6312 9430
rect 6350 9415 6360 9430
rect 6360 9415 6384 9430
rect 6422 9415 6428 9430
rect 6428 9415 6456 9430
rect 6494 9415 6496 9430
rect 6496 9415 6528 9430
rect 6566 9415 6598 9430
rect 6598 9415 6600 9430
rect 6638 9415 6666 9430
rect 6666 9415 6672 9430
rect 6710 9415 6734 9430
rect 6734 9415 6744 9430
rect 6782 9415 6802 9430
rect 6802 9415 6816 9430
rect 6854 9415 6870 9430
rect 6870 9415 6888 9430
rect 6926 9415 6938 9430
rect 6938 9415 6960 9430
rect 6998 9415 7006 9430
rect 7006 9415 7032 9430
rect 7070 9415 7074 9430
rect 7074 9415 7104 9430
rect 7142 9415 7176 9430
rect 7214 9415 7244 9430
rect 7244 9415 7248 9430
rect 7286 9415 7312 9430
rect 7312 9415 7320 9430
rect 7358 9415 7380 9430
rect 7380 9415 7392 9430
rect 7493 9403 7527 9437
rect 7579 9403 7613 9437
rect 2141 9362 2319 9396
rect 2141 9328 2290 9362
rect 2290 9328 2319 9362
rect 2480 9340 2514 9341
rect 2553 9340 2587 9341
rect 2626 9340 2660 9341
rect 2699 9340 2733 9341
rect 2772 9340 2806 9341
rect 2845 9340 2879 9341
rect 2918 9340 2952 9341
rect 2991 9340 3025 9341
rect 3064 9340 3098 9341
rect 3137 9340 3171 9341
rect 3210 9340 3244 9341
rect 3283 9340 3317 9341
rect 3356 9340 3390 9341
rect 3429 9340 3463 9341
rect 3502 9340 3536 9341
rect 3575 9340 3609 9341
rect 3648 9340 3682 9341
rect 3721 9340 3755 9341
rect 3794 9340 3828 9341
rect 3867 9340 3901 9341
rect 3940 9340 3974 9341
rect 4013 9340 4047 9341
rect 2141 9294 2319 9328
rect 2480 9307 2488 9340
rect 2488 9307 2514 9340
rect 2553 9307 2556 9340
rect 2556 9307 2587 9340
rect 2626 9307 2658 9340
rect 2658 9307 2660 9340
rect 2699 9307 2726 9340
rect 2726 9307 2733 9340
rect 2772 9307 2794 9340
rect 2794 9307 2806 9340
rect 2845 9307 2862 9340
rect 2862 9307 2879 9340
rect 2918 9307 2930 9340
rect 2930 9307 2952 9340
rect 2991 9307 2998 9340
rect 2998 9307 3025 9340
rect 3064 9307 3066 9340
rect 3066 9307 3098 9340
rect 3137 9307 3168 9340
rect 3168 9307 3171 9340
rect 3210 9307 3236 9340
rect 3236 9307 3244 9340
rect 3283 9307 3304 9340
rect 3304 9307 3317 9340
rect 3356 9307 3372 9340
rect 3372 9307 3390 9340
rect 3429 9307 3440 9340
rect 3440 9307 3463 9340
rect 3502 9307 3508 9340
rect 3508 9307 3536 9340
rect 3575 9307 3576 9340
rect 3576 9307 3609 9340
rect 3648 9307 3678 9340
rect 3678 9307 3682 9340
rect 3721 9307 3746 9340
rect 3746 9307 3755 9340
rect 3794 9307 3814 9340
rect 3814 9307 3828 9340
rect 3867 9307 3882 9340
rect 3882 9307 3901 9340
rect 3940 9307 3950 9340
rect 3950 9307 3974 9340
rect 4013 9307 4018 9340
rect 4018 9307 4047 9340
rect 4086 9307 4120 9341
rect 4159 9340 4193 9341
rect 4232 9340 4266 9341
rect 4305 9340 4339 9341
rect 4378 9340 4412 9341
rect 4451 9340 4485 9341
rect 4524 9340 4558 9341
rect 4597 9340 4631 9341
rect 4670 9340 4704 9341
rect 4742 9340 4776 9341
rect 4814 9340 4848 9341
rect 4886 9340 4920 9341
rect 4958 9340 4992 9341
rect 5030 9340 5064 9341
rect 5102 9340 5136 9341
rect 4159 9307 4188 9340
rect 4188 9307 4193 9340
rect 4232 9307 4256 9340
rect 4256 9307 4266 9340
rect 4305 9307 4324 9340
rect 4324 9307 4339 9340
rect 4378 9307 4392 9340
rect 4392 9307 4412 9340
rect 4451 9307 4460 9340
rect 4460 9307 4485 9340
rect 4524 9307 4528 9340
rect 4528 9307 4558 9340
rect 4597 9307 4630 9340
rect 4630 9307 4631 9340
rect 4670 9307 4698 9340
rect 4698 9307 4704 9340
rect 4742 9307 4766 9340
rect 4766 9307 4776 9340
rect 4814 9307 4834 9340
rect 4834 9307 4848 9340
rect 4886 9307 4902 9340
rect 4902 9307 4920 9340
rect 4958 9307 4970 9340
rect 4970 9307 4992 9340
rect 5030 9307 5038 9340
rect 5038 9307 5064 9340
rect 5102 9307 5106 9340
rect 5106 9307 5136 9340
rect 5174 9307 5208 9341
rect 5246 9340 5280 9341
rect 5318 9340 5352 9341
rect 5390 9340 5424 9341
rect 5462 9340 5496 9341
rect 5534 9340 5568 9341
rect 5606 9340 5640 9341
rect 5678 9340 5712 9341
rect 5750 9340 5784 9341
rect 5822 9340 5856 9341
rect 5894 9340 5928 9341
rect 5966 9340 6000 9341
rect 6038 9340 6072 9341
rect 6110 9340 6144 9341
rect 6182 9340 6216 9341
rect 6254 9340 6288 9341
rect 6326 9340 6360 9341
rect 5246 9307 5276 9340
rect 5276 9307 5280 9340
rect 5318 9307 5344 9340
rect 5344 9307 5352 9340
rect 5390 9307 5412 9340
rect 5412 9307 5424 9340
rect 5462 9307 5480 9340
rect 5480 9307 5496 9340
rect 5534 9307 5548 9340
rect 5548 9307 5568 9340
rect 5606 9307 5616 9340
rect 5616 9307 5640 9340
rect 5678 9307 5684 9340
rect 5684 9307 5712 9340
rect 5750 9307 5752 9340
rect 5752 9307 5784 9340
rect 5822 9307 5854 9340
rect 5854 9307 5856 9340
rect 5894 9307 5922 9340
rect 5922 9307 5928 9340
rect 5966 9307 5990 9340
rect 5990 9307 6000 9340
rect 6038 9307 6058 9340
rect 6058 9307 6072 9340
rect 6110 9307 6126 9340
rect 6126 9307 6144 9340
rect 6182 9307 6194 9340
rect 6194 9307 6216 9340
rect 6254 9307 6262 9340
rect 6262 9307 6288 9340
rect 6326 9307 6330 9340
rect 6330 9307 6360 9340
rect 6398 9307 6432 9341
rect 6470 9340 6504 9341
rect 6542 9340 6576 9341
rect 6614 9340 6648 9341
rect 6686 9340 6720 9341
rect 6758 9340 6792 9341
rect 6830 9340 6864 9341
rect 6902 9340 6936 9341
rect 6974 9340 7008 9341
rect 7046 9340 7080 9341
rect 7118 9340 7152 9341
rect 7190 9340 7224 9341
rect 7262 9340 7296 9341
rect 7334 9340 7368 9341
rect 6470 9307 6500 9340
rect 6500 9307 6504 9340
rect 6542 9307 6568 9340
rect 6568 9307 6576 9340
rect 6614 9307 6636 9340
rect 6636 9307 6648 9340
rect 6686 9307 6704 9340
rect 6704 9307 6720 9340
rect 6758 9307 6772 9340
rect 6772 9307 6792 9340
rect 6830 9307 6840 9340
rect 6840 9307 6864 9340
rect 6902 9307 6908 9340
rect 6908 9307 6936 9340
rect 6974 9307 6976 9340
rect 6976 9307 7008 9340
rect 7046 9307 7078 9340
rect 7078 9307 7080 9340
rect 7118 9307 7146 9340
rect 7146 9307 7152 9340
rect 7190 9307 7214 9340
rect 7214 9307 7224 9340
rect 7262 9307 7282 9340
rect 7282 9307 7296 9340
rect 7334 9307 7350 9340
rect 7350 9307 7368 9340
rect 7493 9336 7521 9365
rect 7521 9336 7527 9365
rect 7493 9331 7527 9336
rect 7579 9331 7613 9365
rect 2141 9260 2290 9294
rect 2290 9260 2319 9294
rect 2141 9226 2319 9260
rect 2141 9192 2290 9226
rect 2290 9192 2319 9226
rect 7493 9268 7521 9293
rect 7521 9268 7527 9293
rect 7493 9259 7527 9268
rect 7579 9259 7613 9293
rect 2141 9158 2319 9192
rect 2141 9124 2290 9158
rect 2290 9124 2319 9158
rect 2141 9090 2319 9124
rect 2141 9056 2290 9090
rect 2290 9056 2319 9090
rect 2141 9022 2319 9056
rect 2141 8988 2290 9022
rect 2290 8988 2319 9022
rect 2141 8954 2319 8988
rect 2141 8920 2290 8954
rect 2290 8920 2319 8954
rect 2141 8886 2319 8920
rect 2141 8852 2290 8886
rect 2290 8852 2319 8886
rect 2141 8818 2319 8852
rect 2141 8784 2290 8818
rect 2290 8784 2319 8818
rect 2141 8750 2319 8784
rect 2141 8716 2290 8750
rect 2290 8716 2319 8750
rect 2141 8682 2319 8716
rect 2141 8648 2290 8682
rect 2290 8648 2319 8682
rect 2141 8614 2319 8648
rect 2141 8580 2290 8614
rect 2290 8580 2319 8614
rect 2141 8546 2319 8580
rect 2141 8512 2290 8546
rect 2290 8512 2319 8546
rect 2141 8478 2319 8512
rect 2141 8444 2290 8478
rect 2290 8444 2319 8478
rect 2141 8410 2319 8444
rect 2141 8376 2290 8410
rect 2290 8376 2319 8410
rect 2141 8342 2319 8376
rect 2141 8308 2290 8342
rect 2290 8308 2319 8342
rect 2141 8274 2319 8308
rect 2141 8240 2290 8274
rect 2290 8240 2319 8274
rect 2141 8206 2319 8240
rect 2141 8172 2290 8206
rect 2290 8172 2319 8206
rect 2141 8138 2319 8172
rect 2141 8104 2290 8138
rect 2290 8104 2319 8138
rect 2141 8070 2319 8104
rect 2141 8036 2290 8070
rect 2290 8036 2319 8070
rect 2141 8002 2319 8036
rect 2141 7968 2290 8002
rect 2290 7968 2319 8002
rect 2141 7934 2319 7968
rect 2141 7900 2290 7934
rect 2290 7900 2319 7934
rect 2141 7866 2319 7900
rect 2141 7832 2290 7866
rect 2290 7832 2319 7866
rect 2422 9178 2456 9212
rect 2422 9105 2456 9139
rect 2422 9032 2456 9066
rect 2422 8959 2456 8993
rect 2422 8886 2456 8920
rect 2422 8813 2456 8847
rect 2422 8740 2456 8774
rect 2422 8667 2456 8701
rect 2422 8594 2456 8628
rect 2422 8520 2456 8554
rect 2422 8446 2456 8480
rect 2422 8372 2456 8406
rect 2422 8298 2456 8332
rect 2422 8224 2456 8258
rect 2422 8150 2456 8184
rect 2422 8076 2456 8110
rect 2422 8002 2456 8036
rect 2422 7928 2456 7962
rect 2422 7854 2456 7888
rect 4079 9178 4113 9212
rect 4079 9105 4113 9139
rect 4079 9032 4113 9066
rect 4079 8959 4113 8993
rect 4079 8886 4113 8920
rect 4079 8813 4113 8847
rect 4079 8740 4113 8774
rect 4079 8667 4113 8701
rect 4079 8594 4113 8628
rect 4079 8520 4113 8554
rect 4079 8446 4113 8480
rect 4079 8372 4113 8406
rect 4079 8298 4113 8332
rect 4079 8224 4113 8258
rect 4079 8150 4113 8184
rect 4079 8076 4113 8110
rect 4079 8002 4113 8036
rect 4079 7928 4113 7962
rect 4079 7854 4113 7888
rect 5737 9178 5771 9212
rect 5737 9105 5771 9139
rect 5737 9032 5771 9066
rect 5737 8959 5771 8993
rect 5737 8886 5771 8920
rect 5737 8813 5771 8847
rect 5737 8740 5771 8774
rect 5737 8667 5771 8701
rect 5737 8594 5771 8628
rect 5737 8520 5771 8554
rect 5737 8446 5771 8480
rect 5737 8372 5771 8406
rect 5737 8298 5771 8332
rect 5737 8224 5771 8258
rect 5737 8150 5771 8184
rect 5737 8076 5771 8110
rect 5737 8002 5771 8036
rect 5737 7928 5771 7962
rect 5737 7854 5771 7888
rect 7386 9178 7420 9212
rect 7386 9105 7420 9139
rect 7386 9032 7420 9066
rect 7386 8959 7420 8993
rect 7386 8886 7420 8920
rect 7386 8813 7420 8847
rect 7386 8740 7420 8774
rect 7386 8667 7420 8701
rect 7386 8594 7420 8628
rect 7386 8520 7420 8554
rect 7386 8446 7420 8480
rect 7386 8372 7420 8406
rect 7386 8298 7420 8332
rect 7386 8224 7420 8258
rect 7386 8150 7420 8184
rect 7386 8076 7420 8110
rect 7386 8002 7420 8036
rect 7386 7928 7420 7962
rect 7386 7854 7420 7888
rect 7493 9200 7521 9221
rect 7521 9200 7527 9221
rect 7493 9187 7527 9200
rect 7579 9187 7613 9221
rect 7493 9132 7521 9149
rect 7521 9132 7527 9149
rect 7493 9115 7527 9132
rect 7579 9115 7613 9149
rect 7493 9064 7521 9077
rect 7521 9064 7527 9077
rect 7493 9043 7527 9064
rect 7579 9043 7613 9077
rect 7493 8996 7521 9005
rect 7521 8996 7527 9005
rect 7493 8971 7527 8996
rect 7579 8971 7613 9005
rect 7493 8928 7521 8933
rect 7521 8928 7527 8933
rect 7493 8899 7527 8928
rect 7579 8899 7613 8933
rect 7493 8860 7521 8861
rect 7521 8860 7527 8861
rect 7493 8827 7527 8860
rect 7579 8827 7613 8861
rect 7493 8758 7527 8789
rect 7493 8755 7521 8758
rect 7521 8755 7527 8758
rect 7579 8755 7613 8789
rect 7493 8690 7527 8717
rect 7493 8683 7521 8690
rect 7521 8683 7527 8690
rect 7579 8683 7613 8717
rect 7493 8622 7527 8645
rect 7493 8611 7521 8622
rect 7521 8611 7527 8622
rect 7579 8611 7613 8645
rect 7493 8554 7527 8573
rect 7493 8539 7521 8554
rect 7521 8539 7527 8554
rect 7579 8539 7613 8573
rect 7493 8486 7527 8501
rect 7493 8467 7521 8486
rect 7521 8467 7527 8486
rect 7579 8467 7613 8501
rect 7493 8418 7527 8429
rect 7493 8395 7521 8418
rect 7521 8395 7527 8418
rect 7579 8395 7613 8429
rect 7493 8350 7527 8357
rect 7493 8323 7521 8350
rect 7521 8323 7527 8350
rect 7579 8323 7613 8357
rect 7493 8282 7527 8285
rect 7493 8251 7521 8282
rect 7521 8251 7527 8282
rect 7579 8251 7613 8285
rect 7493 8180 7521 8213
rect 7521 8180 7527 8213
rect 7493 8179 7527 8180
rect 7579 8179 7613 8213
rect 7493 8112 7521 8141
rect 7521 8112 7527 8141
rect 7493 8107 7527 8112
rect 7579 8107 7613 8141
rect 7493 8044 7521 8069
rect 7521 8044 7527 8069
rect 7493 8035 7527 8044
rect 7579 8035 7613 8069
rect 7493 7976 7521 7997
rect 7521 7976 7527 7997
rect 7493 7963 7527 7976
rect 7579 7963 7613 7997
rect 7493 7908 7521 7925
rect 7521 7908 7527 7925
rect 7493 7891 7527 7908
rect 7579 7891 7613 7925
rect 2141 7798 2319 7832
rect 2141 7764 2290 7798
rect 2290 7764 2319 7798
rect 2141 7730 2319 7764
rect 2141 7696 2290 7730
rect 2290 7696 2319 7730
rect 2141 7662 2319 7696
rect 7493 7840 7521 7853
rect 7521 7840 7527 7853
rect 7493 7819 7527 7840
rect 7579 7819 7613 7853
rect 7493 7772 7521 7781
rect 7521 7772 7527 7781
rect 7493 7747 7527 7772
rect 7579 7747 7613 7781
rect 7493 7704 7521 7709
rect 7521 7704 7527 7709
rect 2141 7628 2290 7662
rect 2290 7628 2319 7662
rect 2357 7647 2358 7681
rect 2358 7647 2391 7681
rect 2429 7647 2461 7681
rect 2461 7647 2463 7681
rect 2501 7647 2530 7681
rect 2530 7647 2535 7681
rect 2573 7647 2599 7681
rect 2599 7647 2607 7681
rect 2645 7647 2668 7681
rect 2668 7647 2679 7681
rect 2717 7647 2737 7681
rect 2737 7647 2751 7681
rect 2789 7647 2806 7681
rect 2806 7647 2823 7681
rect 2861 7647 2875 7681
rect 2875 7647 2895 7681
rect 2933 7647 2944 7681
rect 2944 7647 2967 7681
rect 3005 7647 3013 7681
rect 3013 7647 3039 7681
rect 3077 7647 3082 7681
rect 3082 7647 3111 7681
rect 3149 7647 3151 7681
rect 3151 7647 3183 7681
rect 3221 7647 3255 7681
rect 3293 7647 3324 7681
rect 3324 7647 3327 7681
rect 3365 7647 3393 7681
rect 3393 7647 3399 7681
rect 3437 7647 3462 7681
rect 3462 7647 3471 7681
rect 3509 7647 3531 7681
rect 3531 7647 3543 7681
rect 3581 7647 3600 7681
rect 3600 7647 3615 7681
rect 3653 7647 3669 7681
rect 3669 7647 3687 7681
rect 3725 7647 3738 7681
rect 3738 7647 3759 7681
rect 3797 7647 3807 7681
rect 3807 7647 3831 7681
rect 3869 7647 3875 7681
rect 3875 7647 3903 7681
rect 3941 7647 3943 7681
rect 3943 7647 3975 7681
rect 4013 7647 4045 7681
rect 4045 7647 4047 7681
rect 4085 7647 4113 7681
rect 4113 7647 4119 7681
rect 4157 7647 4181 7681
rect 4181 7647 4191 7681
rect 4229 7647 4249 7681
rect 4249 7647 4263 7681
rect 4301 7647 4317 7681
rect 4317 7647 4335 7681
rect 4373 7647 4385 7681
rect 4385 7647 4407 7681
rect 4445 7647 4453 7681
rect 4453 7647 4479 7681
rect 4517 7647 4521 7681
rect 4521 7647 4551 7681
rect 4589 7647 4623 7681
rect 4661 7647 4691 7681
rect 4691 7647 4695 7681
rect 4733 7647 4759 7681
rect 4759 7647 4767 7681
rect 4805 7647 4827 7681
rect 4827 7647 4839 7681
rect 4877 7647 4895 7681
rect 4895 7647 4911 7681
rect 4949 7647 4963 7681
rect 4963 7647 4983 7681
rect 5021 7647 5031 7681
rect 5031 7647 5055 7681
rect 5093 7647 5099 7681
rect 5099 7647 5127 7681
rect 5165 7647 5167 7681
rect 5167 7647 5199 7681
rect 5237 7647 5269 7681
rect 5269 7647 5271 7681
rect 5309 7647 5337 7681
rect 5337 7647 5343 7681
rect 5381 7647 5405 7681
rect 5405 7647 5415 7681
rect 5453 7647 5473 7681
rect 5473 7647 5487 7681
rect 5525 7647 5541 7681
rect 5541 7647 5559 7681
rect 5597 7647 5609 7681
rect 5609 7647 5631 7681
rect 5669 7647 5677 7681
rect 5677 7647 5703 7681
rect 5741 7647 5745 7681
rect 5745 7647 5775 7681
rect 5813 7647 5847 7681
rect 5885 7647 5915 7681
rect 5915 7647 5919 7681
rect 5957 7647 5983 7681
rect 5983 7647 5991 7681
rect 6029 7647 6051 7681
rect 6051 7647 6063 7681
rect 6101 7647 6119 7681
rect 6119 7647 6135 7681
rect 6173 7647 6187 7681
rect 6187 7647 6207 7681
rect 6245 7647 6255 7681
rect 6255 7647 6279 7681
rect 6317 7647 6323 7681
rect 6323 7647 6351 7681
rect 6389 7647 6391 7681
rect 6391 7647 6423 7681
rect 6461 7647 6493 7681
rect 6493 7647 6495 7681
rect 6533 7647 6561 7681
rect 6561 7647 6567 7681
rect 6605 7647 6629 7681
rect 6629 7647 6639 7681
rect 6677 7647 6697 7681
rect 6697 7647 6711 7681
rect 6749 7647 6765 7681
rect 6765 7647 6783 7681
rect 6821 7647 6833 7681
rect 6833 7647 6855 7681
rect 6893 7647 6901 7681
rect 6901 7647 6927 7681
rect 6965 7647 6969 7681
rect 6969 7647 6999 7681
rect 7037 7647 7071 7681
rect 7109 7647 7139 7681
rect 7139 7647 7143 7681
rect 7181 7647 7207 7681
rect 7207 7647 7215 7681
rect 7253 7647 7275 7681
rect 7275 7647 7287 7681
rect 7325 7647 7343 7681
rect 7343 7647 7359 7681
rect 7397 7647 7411 7681
rect 7411 7647 7431 7681
rect 7493 7675 7527 7704
rect 7579 7675 7613 7709
rect 2141 7594 2319 7628
rect 2141 7560 2290 7594
rect 2290 7560 2319 7594
rect 2141 7526 2319 7560
rect 7493 7636 7521 7637
rect 7521 7636 7527 7637
rect 7493 7603 7527 7636
rect 7579 7603 7613 7637
rect 2141 7492 2290 7526
rect 2290 7492 2319 7526
rect 2480 7506 2488 7540
rect 2488 7506 2514 7540
rect 2553 7506 2556 7540
rect 2556 7506 2587 7540
rect 2626 7506 2658 7540
rect 2658 7506 2660 7540
rect 2699 7506 2726 7540
rect 2726 7506 2733 7540
rect 2772 7506 2794 7540
rect 2794 7506 2806 7540
rect 2845 7506 2862 7540
rect 2862 7506 2879 7540
rect 2918 7506 2930 7540
rect 2930 7506 2952 7540
rect 2991 7506 2998 7540
rect 2998 7506 3025 7540
rect 3064 7506 3066 7540
rect 3066 7506 3098 7540
rect 3137 7506 3168 7540
rect 3168 7506 3171 7540
rect 3210 7506 3236 7540
rect 3236 7506 3244 7540
rect 3283 7506 3304 7540
rect 3304 7506 3317 7540
rect 3356 7506 3372 7540
rect 3372 7506 3390 7540
rect 3429 7506 3440 7540
rect 3440 7506 3463 7540
rect 3502 7506 3508 7540
rect 3508 7506 3536 7540
rect 3575 7506 3576 7540
rect 3576 7506 3609 7540
rect 3648 7506 3678 7540
rect 3678 7506 3682 7540
rect 3721 7506 3746 7540
rect 3746 7506 3755 7540
rect 3794 7506 3814 7540
rect 3814 7506 3828 7540
rect 3867 7506 3882 7540
rect 3882 7506 3901 7540
rect 3940 7506 3950 7540
rect 3950 7506 3974 7540
rect 4013 7506 4018 7540
rect 4018 7506 4047 7540
rect 4086 7506 4120 7540
rect 4159 7506 4188 7540
rect 4188 7506 4193 7540
rect 4232 7506 4256 7540
rect 4256 7506 4266 7540
rect 4305 7506 4324 7540
rect 4324 7506 4339 7540
rect 4378 7506 4392 7540
rect 4392 7506 4412 7540
rect 4451 7506 4460 7540
rect 4460 7506 4485 7540
rect 4524 7506 4528 7540
rect 4528 7506 4558 7540
rect 4597 7506 4630 7540
rect 4630 7506 4631 7540
rect 4670 7506 4698 7540
rect 4698 7506 4704 7540
rect 4742 7506 4766 7540
rect 4766 7506 4776 7540
rect 4814 7506 4834 7540
rect 4834 7506 4848 7540
rect 4886 7506 4902 7540
rect 4902 7506 4920 7540
rect 4958 7506 4970 7540
rect 4970 7506 4992 7540
rect 5030 7506 5038 7540
rect 5038 7506 5064 7540
rect 5102 7506 5106 7540
rect 5106 7506 5136 7540
rect 5174 7506 5208 7540
rect 5246 7506 5276 7540
rect 5276 7506 5280 7540
rect 5318 7506 5344 7540
rect 5344 7506 5352 7540
rect 5390 7506 5412 7540
rect 5412 7506 5424 7540
rect 5462 7506 5480 7540
rect 5480 7506 5496 7540
rect 5534 7506 5548 7540
rect 5548 7506 5568 7540
rect 5606 7506 5616 7540
rect 5616 7506 5640 7540
rect 5678 7506 5684 7540
rect 5684 7506 5712 7540
rect 5750 7506 5752 7540
rect 5752 7506 5784 7540
rect 5822 7506 5854 7540
rect 5854 7506 5856 7540
rect 5894 7506 5922 7540
rect 5922 7506 5928 7540
rect 5966 7506 5990 7540
rect 5990 7506 6000 7540
rect 6038 7506 6058 7540
rect 6058 7506 6072 7540
rect 6110 7506 6126 7540
rect 6126 7506 6144 7540
rect 6182 7506 6194 7540
rect 6194 7506 6216 7540
rect 6254 7506 6262 7540
rect 6262 7506 6288 7540
rect 6326 7506 6330 7540
rect 6330 7506 6360 7540
rect 6398 7506 6432 7540
rect 6470 7506 6500 7540
rect 6500 7506 6504 7540
rect 6542 7506 6568 7540
rect 6568 7506 6576 7540
rect 6614 7506 6636 7540
rect 6636 7506 6648 7540
rect 6686 7506 6704 7540
rect 6704 7506 6720 7540
rect 6758 7506 6772 7540
rect 6772 7506 6792 7540
rect 6830 7506 6840 7540
rect 6840 7506 6864 7540
rect 6902 7506 6908 7540
rect 6908 7506 6936 7540
rect 6974 7506 6976 7540
rect 6976 7506 7008 7540
rect 7046 7506 7078 7540
rect 7078 7506 7080 7540
rect 7118 7506 7146 7540
rect 7146 7506 7152 7540
rect 7190 7506 7214 7540
rect 7214 7506 7224 7540
rect 7262 7506 7282 7540
rect 7282 7506 7296 7540
rect 7334 7506 7350 7540
rect 7350 7506 7368 7540
rect 7493 7534 7527 7565
rect 7493 7531 7521 7534
rect 7521 7531 7527 7534
rect 7579 7531 7613 7565
rect 2141 7458 2319 7492
rect 2141 7424 2290 7458
rect 2290 7424 2319 7458
rect 2141 7390 2319 7424
rect 7493 7466 7527 7493
rect 7493 7459 7521 7466
rect 7521 7459 7527 7466
rect 7579 7459 7613 7493
rect 2141 7356 2290 7390
rect 2290 7356 2319 7390
rect 2141 7322 2319 7356
rect 2141 7288 2290 7322
rect 2290 7288 2319 7322
rect 2141 7254 2319 7288
rect 2141 7220 2290 7254
rect 2290 7220 2319 7254
rect 2141 7186 2319 7220
rect 2141 7152 2290 7186
rect 2290 7152 2319 7186
rect 2141 7118 2319 7152
rect 2141 7084 2290 7118
rect 2290 7084 2319 7118
rect 2141 7050 2319 7084
rect 2141 7016 2290 7050
rect 2290 7016 2319 7050
rect 2141 6982 2319 7016
rect 2141 6948 2290 6982
rect 2290 6948 2319 6982
rect 2141 6914 2319 6948
rect 2141 6880 2290 6914
rect 2290 6880 2319 6914
rect 2141 6846 2319 6880
rect 2141 6812 2290 6846
rect 2290 6812 2319 6846
rect 2141 6778 2319 6812
rect 2141 6744 2290 6778
rect 2290 6744 2319 6778
rect 2141 6710 2319 6744
rect 2141 6676 2290 6710
rect 2290 6676 2319 6710
rect 2141 6642 2319 6676
rect 2141 6608 2290 6642
rect 2290 6608 2319 6642
rect 2141 6574 2319 6608
rect 2141 6540 2290 6574
rect 2290 6540 2319 6574
rect 2141 6506 2319 6540
rect 2141 6472 2290 6506
rect 2290 6472 2319 6506
rect 2141 6438 2319 6472
rect 2141 6404 2290 6438
rect 2290 6404 2319 6438
rect 2141 6370 2319 6404
rect 2141 6336 2290 6370
rect 2290 6336 2319 6370
rect 2141 6302 2319 6336
rect 2141 6268 2290 6302
rect 2290 6268 2319 6302
rect 2141 6234 2319 6268
rect 2141 6200 2290 6234
rect 2290 6200 2319 6234
rect 2141 6166 2319 6200
rect 2141 6132 2290 6166
rect 2290 6132 2319 6166
rect 2141 6098 2319 6132
rect 2141 6064 2290 6098
rect 2290 6064 2319 6098
rect 2141 6030 2319 6064
rect 2422 7378 2456 7412
rect 2422 7305 2456 7339
rect 2422 7232 2456 7266
rect 2422 7159 2456 7193
rect 2422 7086 2456 7120
rect 2422 7013 2456 7047
rect 2422 6940 2456 6974
rect 2422 6867 2456 6901
rect 2422 6794 2456 6828
rect 2422 6720 2456 6754
rect 2422 6646 2456 6680
rect 2422 6572 2456 6606
rect 2422 6498 2456 6532
rect 2422 6424 2456 6458
rect 2422 6350 2456 6384
rect 2422 6276 2456 6310
rect 2422 6202 2456 6236
rect 2422 6128 2456 6162
rect 2422 6054 2456 6088
rect 4079 7378 4113 7412
rect 4079 7305 4113 7339
rect 4079 7232 4113 7266
rect 4079 7159 4113 7193
rect 4079 7086 4113 7120
rect 4079 7013 4113 7047
rect 4079 6940 4113 6974
rect 4079 6867 4113 6901
rect 4079 6794 4113 6828
rect 4079 6720 4113 6754
rect 4079 6646 4113 6680
rect 4079 6572 4113 6606
rect 4079 6498 4113 6532
rect 4079 6424 4113 6458
rect 4079 6350 4113 6384
rect 4079 6276 4113 6310
rect 4079 6202 4113 6236
rect 4079 6128 4113 6162
rect 4079 6054 4113 6088
rect 5737 7378 5771 7412
rect 5737 7305 5771 7339
rect 5737 7232 5771 7266
rect 5737 7159 5771 7193
rect 5737 7086 5771 7120
rect 5737 7013 5771 7047
rect 5737 6940 5771 6974
rect 5737 6867 5771 6901
rect 5737 6794 5771 6828
rect 5737 6720 5771 6754
rect 5737 6646 5771 6680
rect 5737 6572 5771 6606
rect 5737 6498 5771 6532
rect 5737 6424 5771 6458
rect 5737 6350 5771 6384
rect 5737 6276 5771 6310
rect 5737 6202 5771 6236
rect 5737 6128 5771 6162
rect 5737 6054 5771 6088
rect 7386 7378 7420 7412
rect 7386 7305 7420 7339
rect 7386 7232 7420 7266
rect 7386 7159 7420 7193
rect 7386 7086 7420 7120
rect 7386 7013 7420 7047
rect 7386 6940 7420 6974
rect 7386 6867 7420 6901
rect 7386 6794 7420 6828
rect 7386 6720 7420 6754
rect 7386 6646 7420 6680
rect 7386 6572 7420 6606
rect 7386 6498 7420 6532
rect 7386 6424 7420 6458
rect 7386 6350 7420 6384
rect 7386 6276 7420 6310
rect 7386 6202 7420 6236
rect 7386 6128 7420 6162
rect 7386 6054 7420 6088
rect 7493 7398 7527 7421
rect 7493 7387 7521 7398
rect 7521 7387 7527 7398
rect 7579 7387 7613 7421
rect 7493 7330 7527 7349
rect 7493 7315 7521 7330
rect 7521 7315 7527 7330
rect 7579 7315 7613 7349
rect 7493 7262 7527 7277
rect 7493 7243 7521 7262
rect 7521 7243 7527 7262
rect 7579 7243 7613 7277
rect 7493 7194 7527 7205
rect 7493 7171 7521 7194
rect 7521 7171 7527 7194
rect 7579 7171 7613 7205
rect 7493 7126 7527 7133
rect 7493 7099 7521 7126
rect 7521 7099 7527 7126
rect 7579 7099 7613 7133
rect 7493 7058 7527 7061
rect 7493 7027 7521 7058
rect 7521 7027 7527 7058
rect 7579 7027 7613 7061
rect 7493 6956 7521 6989
rect 7521 6956 7527 6989
rect 7493 6955 7527 6956
rect 7579 6955 7613 6989
rect 7493 6888 7521 6917
rect 7521 6888 7527 6917
rect 7493 6883 7527 6888
rect 7579 6883 7613 6917
rect 7493 6820 7521 6845
rect 7521 6820 7527 6845
rect 7493 6811 7527 6820
rect 7579 6811 7613 6845
rect 7493 6752 7521 6773
rect 7521 6752 7527 6773
rect 7493 6739 7527 6752
rect 7579 6739 7613 6773
rect 7493 6684 7521 6701
rect 7521 6684 7527 6701
rect 7493 6667 7527 6684
rect 7579 6667 7613 6701
rect 7493 6616 7521 6629
rect 7521 6616 7527 6629
rect 7493 6595 7527 6616
rect 7579 6595 7613 6629
rect 7493 6548 7521 6557
rect 7521 6548 7527 6557
rect 7493 6523 7527 6548
rect 7579 6523 7613 6557
rect 7493 6480 7521 6485
rect 7521 6480 7527 6485
rect 7493 6451 7527 6480
rect 7579 6451 7613 6485
rect 7493 6412 7521 6413
rect 7521 6412 7527 6413
rect 7493 6379 7527 6412
rect 7579 6379 7613 6413
rect 7493 6310 7527 6341
rect 7493 6307 7521 6310
rect 7521 6307 7527 6310
rect 7579 6307 7613 6341
rect 7493 6242 7527 6269
rect 7493 6235 7521 6242
rect 7521 6235 7527 6242
rect 7579 6235 7613 6269
rect 7493 6174 7527 6197
rect 7493 6163 7521 6174
rect 7521 6163 7527 6174
rect 7579 6163 7613 6197
rect 7493 6106 7527 6125
rect 7493 6091 7521 6106
rect 7521 6091 7527 6106
rect 7579 6091 7613 6125
rect 2141 5996 2290 6030
rect 2290 5996 2319 6030
rect 2141 5962 2319 5996
rect 2141 5928 2290 5962
rect 2290 5928 2319 5962
rect 2141 5894 2319 5928
rect 2141 5860 2290 5894
rect 2290 5860 2319 5894
rect 2141 5826 2319 5860
rect 7493 6038 7527 6053
rect 7493 6019 7521 6038
rect 7521 6019 7527 6038
rect 7579 6019 7613 6053
rect 7493 5970 7527 5981
rect 7493 5947 7521 5970
rect 7521 5947 7527 5970
rect 7579 5947 7613 5981
rect 7493 5902 7527 5909
rect 7493 5875 7521 5902
rect 7521 5875 7527 5902
rect 7579 5875 7613 5909
rect 2141 5792 2290 5826
rect 2290 5792 2319 5826
rect 2363 5807 2392 5841
rect 2392 5807 2397 5841
rect 2436 5807 2461 5841
rect 2461 5807 2470 5841
rect 2509 5807 2530 5841
rect 2530 5807 2543 5841
rect 2582 5807 2599 5841
rect 2599 5807 2616 5841
rect 2655 5807 2668 5841
rect 2668 5807 2689 5841
rect 2728 5807 2737 5841
rect 2737 5807 2762 5841
rect 2801 5807 2806 5841
rect 2806 5807 2835 5841
rect 2874 5807 2875 5841
rect 2875 5807 2908 5841
rect 2947 5807 2979 5841
rect 2979 5807 2981 5841
rect 3020 5807 3048 5841
rect 3048 5807 3054 5841
rect 3093 5807 3117 5841
rect 3117 5807 3127 5841
rect 3166 5807 3186 5841
rect 3186 5807 3200 5841
rect 3239 5807 3255 5841
rect 3255 5807 3273 5841
rect 3312 5807 3324 5841
rect 3324 5807 3346 5841
rect 3385 5807 3393 5841
rect 3393 5807 3419 5841
rect 3458 5807 3462 5841
rect 3462 5807 3492 5841
rect 3531 5807 3565 5841
rect 3604 5807 3634 5841
rect 3634 5807 3638 5841
rect 3677 5807 3703 5841
rect 3703 5807 3711 5841
rect 3750 5807 3771 5841
rect 3771 5807 3784 5841
rect 3823 5807 3839 5841
rect 3839 5807 3857 5841
rect 3896 5807 3907 5841
rect 3907 5807 3930 5841
rect 3969 5807 3975 5841
rect 3975 5807 4003 5841
rect 4042 5807 4043 5841
rect 4043 5807 4076 5841
rect 4115 5807 4145 5841
rect 4145 5807 4149 5841
rect 4188 5807 4213 5841
rect 4213 5807 4222 5841
rect 4261 5807 4281 5841
rect 4281 5807 4295 5841
rect 4334 5807 4349 5841
rect 4349 5807 4368 5841
rect 4407 5807 4417 5841
rect 4417 5807 4441 5841
rect 4480 5807 4485 5841
rect 4485 5807 4514 5841
rect 4553 5807 4587 5841
rect 4626 5807 4655 5841
rect 4655 5807 4660 5841
rect 4699 5807 4723 5841
rect 4723 5807 4733 5841
rect 4772 5807 4791 5841
rect 4791 5807 4806 5841
rect 4845 5807 4859 5841
rect 4859 5807 4879 5841
rect 4918 5807 4927 5841
rect 4927 5807 4952 5841
rect 4991 5807 4995 5841
rect 4995 5807 5025 5841
rect 5064 5807 5097 5841
rect 5097 5807 5098 5841
rect 5137 5807 5165 5841
rect 5165 5807 5171 5841
rect 5210 5807 5233 5841
rect 5233 5807 5244 5841
rect 5283 5807 5301 5841
rect 5301 5807 5317 5841
rect 5356 5807 5369 5841
rect 5369 5807 5390 5841
rect 5429 5807 5437 5841
rect 5437 5807 5463 5841
rect 5502 5807 5505 5841
rect 5505 5807 5536 5841
rect 5575 5807 5607 5841
rect 5607 5807 5609 5841
rect 5648 5807 5675 5841
rect 5675 5807 5682 5841
rect 5721 5807 5743 5841
rect 5743 5807 5755 5841
rect 5794 5807 5811 5841
rect 5811 5807 5828 5841
rect 5867 5807 5879 5841
rect 5879 5807 5901 5841
rect 5940 5807 5947 5841
rect 5947 5807 5974 5841
rect 6013 5807 6015 5841
rect 6015 5807 6047 5841
rect 6086 5807 6117 5841
rect 6117 5807 6120 5841
rect 6159 5807 6185 5841
rect 6185 5807 6193 5841
rect 6232 5807 6253 5841
rect 6253 5807 6266 5841
rect 6305 5807 6321 5841
rect 6321 5807 6339 5841
rect 6378 5807 6389 5841
rect 6389 5807 6412 5841
rect 6451 5807 6457 5841
rect 6457 5807 6485 5841
rect 6524 5807 6525 5841
rect 6525 5807 6558 5841
rect 6597 5807 6627 5841
rect 6627 5807 6631 5841
rect 6670 5807 6695 5841
rect 6695 5807 6704 5841
rect 6743 5807 6763 5841
rect 6763 5807 6777 5841
rect 6816 5807 6831 5841
rect 6831 5807 6850 5841
rect 6889 5807 6899 5841
rect 6899 5807 6923 5841
rect 6962 5807 6967 5841
rect 6967 5807 6996 5841
rect 7035 5807 7069 5841
rect 7108 5807 7137 5841
rect 7137 5807 7142 5841
rect 7181 5807 7205 5841
rect 7205 5807 7215 5841
rect 7253 5807 7273 5841
rect 7273 5807 7287 5841
rect 7325 5807 7341 5841
rect 7341 5807 7359 5841
rect 7397 5807 7409 5841
rect 7409 5807 7431 5841
rect 7493 5834 7527 5837
rect 7493 5803 7521 5834
rect 7521 5803 7527 5834
rect 7579 5803 7613 5837
rect 2141 5758 2319 5792
rect 2141 5724 2290 5758
rect 2290 5724 2319 5758
rect 2141 5690 2319 5724
rect 2141 5656 2290 5690
rect 2290 5656 2319 5690
rect 2141 5622 2319 5656
rect 7493 5732 7521 5765
rect 7521 5732 7527 5765
rect 7493 5731 7527 5732
rect 7579 5731 7613 5765
rect 7493 5664 7521 5693
rect 7521 5664 7527 5693
rect 7493 5659 7527 5664
rect 7579 5659 7613 5693
rect 2141 5588 2290 5622
rect 2290 5588 2319 5622
rect 2640 5611 2660 5645
rect 2660 5611 2674 5645
rect 2713 5611 2728 5645
rect 2728 5611 2747 5645
rect 2786 5611 2796 5645
rect 2796 5611 2820 5645
rect 2859 5611 2864 5645
rect 2864 5611 2893 5645
rect 2932 5611 2966 5645
rect 3005 5611 3034 5645
rect 3034 5611 3039 5645
rect 3078 5611 3102 5645
rect 3102 5611 3112 5645
rect 3151 5611 3170 5645
rect 3170 5611 3185 5645
rect 3224 5611 3238 5645
rect 3238 5611 3258 5645
rect 3297 5611 3306 5645
rect 3306 5611 3331 5645
rect 3370 5611 3374 5645
rect 3374 5611 3404 5645
rect 3443 5611 3476 5645
rect 3476 5611 3477 5645
rect 3516 5611 3544 5645
rect 3544 5611 3550 5645
rect 3589 5611 3612 5645
rect 3612 5611 3623 5645
rect 3662 5611 3680 5645
rect 3680 5611 3696 5645
rect 3735 5611 3748 5645
rect 3748 5611 3769 5645
rect 3808 5611 3816 5645
rect 3816 5611 3842 5645
rect 3881 5611 3884 5645
rect 3884 5611 3915 5645
rect 3954 5611 3986 5645
rect 3986 5611 3988 5645
rect 4027 5611 4054 5645
rect 4054 5611 4061 5645
rect 4100 5611 4122 5645
rect 4122 5611 4134 5645
rect 4173 5611 4190 5645
rect 4190 5611 4207 5645
rect 4246 5611 4258 5645
rect 4258 5611 4280 5645
rect 4319 5611 4326 5645
rect 4326 5611 4353 5645
rect 4392 5611 4394 5645
rect 4394 5611 4426 5645
rect 4465 5611 4496 5645
rect 4496 5611 4499 5645
rect 4538 5611 4564 5645
rect 4564 5611 4572 5645
rect 4611 5611 4632 5645
rect 4632 5611 4645 5645
rect 4684 5611 4700 5645
rect 4700 5611 4718 5645
rect 4757 5611 4768 5645
rect 4768 5611 4791 5645
rect 4830 5611 4836 5645
rect 4836 5611 4864 5645
rect 4903 5611 4904 5645
rect 4904 5611 4937 5645
rect 4976 5611 5006 5645
rect 5006 5611 5010 5645
rect 5049 5611 5074 5645
rect 5074 5611 5083 5645
rect 5122 5611 5142 5645
rect 5142 5611 5156 5645
rect 5195 5611 5210 5645
rect 5210 5611 5229 5645
rect 5268 5611 5278 5645
rect 5278 5611 5302 5645
rect 5341 5611 5346 5645
rect 5346 5611 5375 5645
rect 5414 5611 5448 5645
rect 5487 5611 5516 5645
rect 5516 5611 5521 5645
rect 5560 5611 5584 5645
rect 5584 5611 5594 5645
rect 5633 5611 5652 5645
rect 5652 5611 5667 5645
rect 5706 5611 5720 5645
rect 5720 5611 5740 5645
rect 5778 5611 5788 5645
rect 5788 5611 5812 5645
rect 5850 5611 5856 5645
rect 5856 5611 5884 5645
rect 5922 5611 5924 5645
rect 5924 5611 5956 5645
rect 5994 5611 6026 5645
rect 6026 5611 6028 5645
rect 6066 5611 6094 5645
rect 6094 5611 6100 5645
rect 6138 5611 6162 5645
rect 6162 5611 6172 5645
rect 6210 5611 6230 5645
rect 6230 5611 6244 5645
rect 6282 5611 6298 5645
rect 6298 5611 6316 5645
rect 6354 5611 6366 5645
rect 6366 5611 6388 5645
rect 6426 5611 6434 5645
rect 6434 5611 6460 5645
rect 6498 5611 6502 5645
rect 6502 5611 6532 5645
rect 6570 5611 6604 5645
rect 6642 5611 6672 5645
rect 6672 5611 6676 5645
rect 6714 5611 6740 5645
rect 6740 5611 6748 5645
rect 6786 5611 6808 5645
rect 6808 5611 6820 5645
rect 6858 5611 6876 5645
rect 6876 5611 6892 5645
rect 6930 5611 6944 5645
rect 6944 5611 6964 5645
rect 7002 5611 7036 5645
rect 2141 5554 2319 5588
rect 2141 5520 2290 5554
rect 2290 5520 2319 5554
rect 7493 5596 7521 5621
rect 7521 5596 7527 5621
rect 7493 5587 7527 5596
rect 7579 5587 7613 5621
rect 2141 5486 2319 5520
rect 2141 5452 2290 5486
rect 2290 5452 2319 5486
rect 2141 5418 2319 5452
rect 2141 5384 2290 5418
rect 2290 5384 2319 5418
rect 2141 5350 2319 5384
rect 2141 5316 2290 5350
rect 2290 5316 2319 5350
rect 2687 5512 2721 5546
rect 2687 5438 2721 5472
rect 2687 5364 2721 5398
rect 2141 5305 2319 5316
rect 2141 5232 2175 5266
rect 2213 5232 2247 5266
rect 2285 5248 2290 5266
rect 2290 5248 2319 5266
rect 2285 5232 2319 5248
rect 2141 5159 2175 5193
rect 2213 5159 2247 5193
rect 2285 5180 2290 5193
rect 2290 5180 2319 5193
rect 2285 5159 2319 5180
rect 2141 5086 2175 5120
rect 2213 5086 2247 5120
rect 2285 5112 2290 5120
rect 2290 5112 2319 5120
rect 2285 5086 2319 5112
rect 2141 5013 2175 5047
rect 2213 5013 2247 5047
rect 2285 5044 2290 5047
rect 2290 5044 2319 5047
rect 2285 5013 2319 5044
rect 2141 4940 2175 4974
rect 2213 4940 2247 4974
rect 2285 4942 2319 4974
rect 2285 4940 2290 4942
rect 2290 4940 2319 4942
rect 2141 4867 2175 4901
rect 2213 4867 2247 4901
rect 2285 4874 2319 4901
rect 2285 4867 2290 4874
rect 2290 4867 2319 4874
rect 2141 4794 2175 4828
rect 2213 4794 2247 4828
rect 2285 4806 2319 4828
rect 2285 4794 2290 4806
rect 2290 4794 2319 4806
rect 2141 4721 2175 4755
rect 2213 4721 2247 4755
rect 2285 4738 2319 4755
rect 2285 4721 2290 4738
rect 2290 4721 2319 4738
rect 2141 4648 2175 4682
rect 2213 4648 2247 4682
rect 2285 4670 2319 4682
rect 2285 4648 2290 4670
rect 2290 4648 2319 4670
rect 2141 4575 2175 4609
rect 2213 4575 2247 4609
rect 2285 4602 2319 4609
rect 2285 4575 2290 4602
rect 2290 4575 2319 4602
rect 2141 4502 2175 4536
rect 2213 4502 2247 4536
rect 2285 4534 2319 4536
rect 2285 4502 2290 4534
rect 2290 4502 2319 4534
rect 2141 4429 2175 4463
rect 2213 4429 2247 4463
rect 2285 4432 2290 4463
rect 2290 4432 2319 4463
rect 2285 4429 2319 4432
rect 2141 4356 2175 4390
rect 2213 4356 2247 4390
rect 2285 4364 2290 4390
rect 2290 4364 2319 4390
rect 2285 4356 2319 4364
rect 2141 4283 2175 4317
rect 2213 4283 2247 4317
rect 2285 4296 2290 4317
rect 2290 4296 2319 4317
rect 2285 4283 2319 4296
rect 2141 4210 2175 4244
rect 2213 4210 2247 4244
rect 2285 4228 2290 4244
rect 2290 4228 2319 4244
rect 2285 4210 2319 4228
rect 2141 4137 2175 4171
rect 2213 4137 2247 4171
rect 2285 4160 2290 4171
rect 2290 4160 2319 4171
rect 2595 5285 2629 5319
rect 2595 5211 2629 5245
rect 2595 5137 2629 5171
rect 2595 5063 2629 5097
rect 2595 4989 2629 5023
rect 2595 4915 2629 4949
rect 2595 4841 2629 4875
rect 2595 4767 2629 4801
rect 2595 4693 2629 4727
rect 2595 4619 2629 4653
rect 2595 4545 2629 4579
rect 2595 4470 2629 4504
rect 2595 4395 2629 4429
rect 2595 4320 2629 4354
rect 2595 4245 2629 4279
rect 2595 4170 2629 4204
rect 2687 5290 2721 5324
rect 7493 5528 7521 5549
rect 7521 5528 7527 5549
rect 7493 5515 7527 5528
rect 7579 5515 7613 5549
rect 7493 5460 7521 5477
rect 7521 5460 7527 5477
rect 7493 5443 7527 5460
rect 7579 5443 7613 5477
rect 7493 5392 7521 5405
rect 7521 5392 7527 5405
rect 7493 5371 7527 5392
rect 7579 5371 7613 5405
rect 7493 5324 7521 5333
rect 7521 5324 7527 5333
rect 2687 5216 2721 5250
rect 2687 5142 2721 5176
rect 2687 5068 2721 5102
rect 2687 4994 2721 5028
rect 2687 4920 2721 4954
rect 2687 4845 2721 4879
rect 2687 4770 2721 4804
rect 2687 4695 2721 4729
rect 2687 4620 2721 4654
rect 2687 4545 2721 4579
rect 2687 4470 2721 4504
rect 2687 4395 2721 4429
rect 2687 4320 2721 4354
rect 2687 4245 2721 4279
rect 2687 4170 2721 4204
rect 2779 5285 2813 5319
rect 2779 5211 2813 5245
rect 2779 5137 2813 5171
rect 2779 5063 2813 5097
rect 2779 4989 2813 5023
rect 2779 4915 2813 4949
rect 2779 4841 2813 4875
rect 2779 4767 2813 4801
rect 2779 4693 2813 4727
rect 2779 4619 2813 4653
rect 2779 4545 2813 4579
rect 2779 4470 2813 4504
rect 2779 4395 2813 4429
rect 2779 4320 2813 4354
rect 2779 4245 2813 4279
rect 2779 4170 2813 4204
rect 3632 5285 3666 5319
rect 3632 5210 3666 5244
rect 3632 5135 3666 5169
rect 3632 5060 3666 5094
rect 3632 4985 3666 5019
rect 3632 4910 3666 4944
rect 3632 4835 3666 4869
rect 3632 4760 3666 4794
rect 3632 4685 3666 4719
rect 3632 4610 3666 4644
rect 3632 4535 3666 4569
rect 3632 4460 3666 4494
rect 3632 4385 3666 4419
rect 3632 4310 3666 4344
rect 3632 4235 3666 4269
rect 2285 4137 2319 4160
rect 3632 4159 3666 4193
rect 4491 5285 4525 5319
rect 4491 5210 4525 5244
rect 4491 5135 4525 5169
rect 4491 5060 4525 5094
rect 4491 4985 4525 5019
rect 4491 4910 4525 4944
rect 4491 4835 4525 4869
rect 4491 4760 4525 4794
rect 4491 4685 4525 4719
rect 4491 4610 4525 4644
rect 4491 4535 4525 4569
rect 4491 4460 4525 4494
rect 4491 4385 4525 4419
rect 4491 4310 4525 4344
rect 4491 4235 4525 4269
rect 4491 4159 4525 4193
rect 5347 5285 5381 5319
rect 5347 5210 5381 5244
rect 5347 5135 5381 5169
rect 5347 5060 5381 5094
rect 5347 4985 5381 5019
rect 5347 4910 5381 4944
rect 5347 4835 5381 4869
rect 5347 4760 5381 4794
rect 5347 4685 5381 4719
rect 5347 4610 5381 4644
rect 5347 4535 5381 4569
rect 5347 4460 5381 4494
rect 5347 4385 5381 4419
rect 5347 4310 5381 4344
rect 5347 4235 5381 4269
rect 5347 4159 5381 4193
rect 6206 5285 6240 5319
rect 6206 5210 6240 5244
rect 6206 5135 6240 5169
rect 6206 5060 6240 5094
rect 6206 4985 6240 5019
rect 6206 4910 6240 4944
rect 6206 4835 6240 4869
rect 6206 4760 6240 4794
rect 6206 4685 6240 4719
rect 6206 4610 6240 4644
rect 6206 4535 6240 4569
rect 6206 4460 6240 4494
rect 6206 4385 6240 4419
rect 6206 4310 6240 4344
rect 6206 4235 6240 4269
rect 6206 4159 6240 4193
rect 7059 5285 7093 5319
rect 7059 5210 7093 5244
rect 7059 5135 7093 5169
rect 7059 5060 7093 5094
rect 7059 4985 7093 5019
rect 7059 4910 7093 4944
rect 7059 4835 7093 4869
rect 7059 4760 7093 4794
rect 7059 4685 7093 4719
rect 7059 4610 7093 4644
rect 7059 4535 7093 4569
rect 7059 4460 7093 4494
rect 7059 4385 7093 4419
rect 7059 4310 7093 4344
rect 7059 4235 7093 4269
rect 7059 4159 7093 4193
rect 7493 5299 7527 5324
rect 7579 5299 7613 5333
rect 7493 5256 7521 5261
rect 7521 5256 7527 5261
rect 7493 5227 7527 5256
rect 7579 5227 7613 5261
rect 7493 5188 7521 5189
rect 7521 5188 7527 5189
rect 7493 5155 7527 5188
rect 7579 5155 7613 5189
rect 7493 5086 7527 5117
rect 7493 5083 7521 5086
rect 7521 5083 7527 5086
rect 7579 5083 7613 5117
rect 7493 5018 7527 5045
rect 7493 5011 7521 5018
rect 7521 5011 7527 5018
rect 7579 5011 7613 5045
rect 7493 4950 7527 4973
rect 7493 4939 7521 4950
rect 7521 4939 7527 4950
rect 7579 4939 7613 4973
rect 7493 4882 7527 4901
rect 7493 4867 7521 4882
rect 7521 4867 7527 4882
rect 7579 4867 7613 4901
rect 7493 4814 7527 4829
rect 7493 4795 7521 4814
rect 7521 4795 7527 4814
rect 7579 4795 7613 4829
rect 7493 4746 7527 4757
rect 7493 4723 7521 4746
rect 7521 4723 7527 4746
rect 7579 4723 7613 4757
rect 7493 4678 7527 4685
rect 7493 4651 7521 4678
rect 7521 4651 7527 4678
rect 7579 4651 7613 4685
rect 7493 4610 7527 4613
rect 7493 4579 7521 4610
rect 7521 4579 7527 4610
rect 7579 4579 7613 4613
rect 7493 4508 7521 4540
rect 7521 4508 7527 4540
rect 7493 4506 7527 4508
rect 7579 4506 7613 4540
rect 7493 4440 7521 4467
rect 7521 4440 7527 4467
rect 7493 4433 7527 4440
rect 7579 4433 7613 4467
rect 7493 4372 7521 4394
rect 7521 4372 7527 4394
rect 7493 4360 7527 4372
rect 7579 4360 7613 4394
rect 7493 4304 7521 4321
rect 7521 4304 7527 4321
rect 7493 4287 7527 4304
rect 7579 4287 7613 4321
rect 7493 4236 7521 4248
rect 7521 4236 7527 4248
rect 7493 4214 7527 4236
rect 7579 4214 7613 4248
rect 7493 4168 7521 4175
rect 7521 4168 7527 4175
rect 2141 4064 2175 4098
rect 2213 4064 2247 4098
rect 2285 4092 2290 4098
rect 2290 4092 2319 4098
rect 2285 4064 2319 4092
rect 2141 3991 2175 4025
rect 2213 3991 2247 4025
rect 2285 4024 2290 4025
rect 2290 4024 2319 4025
rect 2285 3991 2319 4024
rect 7493 4141 7527 4168
rect 7579 4141 7613 4175
rect 7493 4100 7521 4102
rect 7521 4100 7527 4102
rect 7493 4068 7527 4100
rect 7579 4068 7613 4102
rect 7493 3998 7527 4029
rect 7493 3995 7521 3998
rect 7521 3995 7527 3998
rect 7579 3995 7613 4029
rect 2147 3909 2181 3943
rect 2220 3909 2254 3943
rect 2293 3909 2327 3943
rect 2366 3909 2400 3943
rect 2439 3909 2473 3943
rect 2512 3909 2546 3943
rect 2585 3909 2619 3943
rect 2658 3909 2692 3943
rect 2731 3909 2765 3943
rect 2804 3909 2838 3943
rect 2877 3909 2911 3943
rect 2950 3909 2984 3943
rect 3023 3907 7593 3943
rect 3023 3873 3028 3907
rect 3028 3873 3062 3907
rect 3062 3873 3096 3907
rect 3096 3873 3130 3907
rect 3130 3873 3164 3907
rect 3164 3873 3198 3907
rect 3198 3873 3232 3907
rect 3232 3873 3266 3907
rect 3266 3873 3300 3907
rect 3300 3873 3334 3907
rect 3334 3873 3368 3907
rect 3368 3873 3402 3907
rect 3402 3873 3436 3907
rect 3436 3873 3470 3907
rect 3470 3873 3504 3907
rect 3504 3873 3538 3907
rect 3538 3873 3572 3907
rect 3572 3873 3606 3907
rect 3606 3873 3640 3907
rect 3640 3873 3674 3907
rect 3674 3873 3708 3907
rect 3708 3873 3742 3907
rect 3742 3873 3776 3907
rect 3776 3873 3810 3907
rect 3810 3873 3844 3907
rect 3844 3873 3878 3907
rect 3878 3873 3912 3907
rect 3912 3873 3946 3907
rect 3946 3873 3980 3907
rect 3980 3873 4014 3907
rect 4014 3873 4048 3907
rect 4048 3873 4082 3907
rect 4082 3873 4116 3907
rect 4116 3873 4150 3907
rect 4150 3873 4184 3907
rect 4184 3873 4218 3907
rect 4218 3873 4252 3907
rect 4252 3873 4286 3907
rect 4286 3873 4320 3907
rect 4320 3873 4354 3907
rect 4354 3873 4388 3907
rect 4388 3873 4422 3907
rect 4422 3873 4456 3907
rect 4456 3873 4490 3907
rect 4490 3873 4524 3907
rect 4524 3873 4558 3907
rect 4558 3873 4592 3907
rect 4592 3873 4626 3907
rect 4626 3873 4660 3907
rect 4660 3873 4694 3907
rect 4694 3873 4728 3907
rect 4728 3873 4762 3907
rect 4762 3873 4796 3907
rect 4796 3873 4830 3907
rect 4830 3873 4864 3907
rect 4864 3873 4898 3907
rect 4898 3873 4932 3907
rect 4932 3873 4966 3907
rect 4966 3873 5000 3907
rect 5000 3873 5034 3907
rect 5034 3873 5068 3907
rect 5068 3873 5102 3907
rect 5102 3873 5136 3907
rect 5136 3873 5170 3907
rect 5170 3873 5204 3907
rect 5204 3873 5238 3907
rect 5238 3873 5272 3907
rect 5272 3873 5306 3907
rect 5306 3873 5340 3907
rect 5340 3873 5374 3907
rect 5374 3873 5408 3907
rect 5408 3873 5442 3907
rect 5442 3873 5476 3907
rect 5476 3873 5510 3907
rect 5510 3873 5544 3907
rect 5544 3873 5578 3907
rect 5578 3873 5612 3907
rect 5612 3873 5646 3907
rect 5646 3873 5680 3907
rect 5680 3873 5714 3907
rect 5714 3873 5748 3907
rect 5748 3873 5782 3907
rect 5782 3873 5816 3907
rect 5816 3873 5850 3907
rect 5850 3873 5884 3907
rect 5884 3873 5918 3907
rect 5918 3873 5952 3907
rect 5952 3873 5986 3907
rect 5986 3873 6020 3907
rect 6020 3873 6054 3907
rect 6054 3873 6088 3907
rect 6088 3873 6122 3907
rect 6122 3873 6156 3907
rect 6156 3873 6190 3907
rect 6190 3873 6224 3907
rect 6224 3873 6258 3907
rect 6258 3873 6292 3907
rect 6292 3873 6326 3907
rect 6326 3873 6360 3907
rect 6360 3873 6394 3907
rect 6394 3873 6428 3907
rect 6428 3873 6462 3907
rect 6462 3873 6496 3907
rect 6496 3873 6530 3907
rect 6530 3873 6564 3907
rect 6564 3873 6598 3907
rect 6598 3873 6632 3907
rect 6632 3873 6666 3907
rect 6666 3873 6700 3907
rect 6700 3873 6734 3907
rect 6734 3873 6768 3907
rect 6768 3873 6802 3907
rect 6802 3873 6836 3907
rect 6836 3873 6870 3907
rect 6870 3873 6904 3907
rect 6904 3873 6938 3907
rect 6938 3873 6972 3907
rect 6972 3873 7006 3907
rect 7006 3873 7040 3907
rect 7040 3873 7074 3907
rect 7074 3873 7108 3907
rect 7108 3873 7142 3907
rect 7142 3873 7176 3907
rect 7176 3873 7210 3907
rect 7210 3873 7244 3907
rect 7244 3873 7278 3907
rect 7278 3873 7312 3907
rect 7312 3873 7346 3907
rect 7346 3873 7380 3907
rect 7380 3873 7414 3907
rect 7414 3873 7448 3907
rect 7448 3873 7593 3907
rect 2147 3837 2181 3871
rect 2220 3837 2254 3871
rect 2293 3837 2327 3871
rect 2366 3837 2400 3871
rect 2439 3837 2473 3871
rect 2512 3837 2546 3871
rect 2585 3837 2619 3871
rect 2658 3837 2692 3871
rect 2731 3837 2765 3871
rect 2804 3837 2838 3871
rect 2877 3837 2911 3871
rect 2950 3837 2984 3871
rect 3023 3837 7593 3873
rect 7733 9445 7839 9479
rect 7733 4528 7735 9445
rect 7735 4528 7837 9445
rect 7837 4528 7839 9445
rect 7733 4455 7735 4489
rect 7735 4455 7767 4489
rect 7805 4455 7837 4489
rect 7837 4455 7839 4489
rect 7733 4382 7735 4416
rect 7735 4382 7767 4416
rect 7805 4382 7837 4416
rect 7837 4382 7839 4416
rect 7733 4309 7735 4343
rect 7735 4309 7767 4343
rect 7805 4309 7837 4343
rect 7837 4309 7839 4343
rect 7733 4236 7735 4270
rect 7735 4236 7767 4270
rect 7805 4236 7837 4270
rect 7837 4236 7839 4270
rect 7733 4175 7735 4197
rect 7735 4175 7767 4197
rect 7805 4175 7837 4197
rect 7837 4175 7839 4197
rect 7733 4163 7767 4175
rect 7805 4163 7839 4175
rect 7733 4090 7767 4124
rect 7805 4090 7839 4124
rect 7733 4017 7735 4051
rect 7735 4017 7767 4051
rect 7805 4017 7837 4051
rect 7837 4017 7839 4051
rect 7733 3944 7735 3978
rect 7735 3944 7767 3978
rect 7805 3944 7837 3978
rect 7837 3944 7839 3978
rect 7733 3871 7735 3905
rect 7735 3871 7767 3905
rect 7805 3871 7837 3905
rect 7837 3871 7839 3905
rect 7733 3798 7735 3832
rect 7735 3798 7767 3832
rect 7805 3798 7837 3832
rect 7837 3798 7839 3832
rect 7733 3725 7735 3759
rect 7735 3725 7767 3759
rect 7805 3725 7837 3759
rect 7837 3725 7839 3759
rect 7733 3652 7735 3686
rect 7735 3652 7767 3686
rect 7805 3652 7837 3686
rect 7837 3652 7839 3686
rect 7733 3579 7735 3613
rect 7735 3579 7767 3613
rect 7805 3579 7837 3613
rect 7837 3579 7839 3613
rect 7733 3506 7735 3540
rect 7735 3506 7767 3540
rect 7805 3506 7837 3540
rect 7837 3506 7839 3540
rect 1950 3419 1984 3453
rect 2023 3419 2048 3453
rect 2048 3419 2057 3453
rect 2096 3451 2130 3453
rect 2169 3451 2203 3453
rect 2242 3451 2276 3453
rect 2315 3451 2349 3453
rect 2388 3451 2422 3453
rect 2461 3451 2495 3453
rect 2534 3451 2568 3453
rect 2096 3419 2130 3451
rect 2169 3419 2203 3451
rect 2242 3419 2276 3451
rect 2315 3419 2349 3451
rect 2388 3419 2422 3451
rect 2461 3419 2495 3451
rect 2534 3419 2568 3451
rect 2607 3419 2641 3453
rect 2680 3451 2714 3453
rect 2753 3451 2787 3453
rect 2826 3451 2860 3453
rect 2899 3451 2933 3453
rect 2972 3451 3006 3453
rect 3045 3451 3079 3453
rect 3118 3451 3152 3453
rect 3191 3451 3225 3453
rect 3264 3451 3298 3453
rect 3337 3451 3371 3453
rect 3410 3451 3444 3453
rect 3483 3451 3517 3453
rect 3556 3451 3590 3453
rect 3629 3451 3663 3453
rect 3702 3451 3736 3453
rect 3775 3451 3809 3453
rect 3848 3451 3882 3453
rect 3921 3451 3955 3453
rect 3994 3451 4028 3453
rect 4067 3451 4101 3453
rect 4140 3451 4174 3453
rect 4213 3451 4247 3453
rect 4286 3451 4320 3453
rect 4359 3451 4393 3453
rect 4432 3451 4466 3453
rect 4505 3451 4539 3453
rect 4578 3451 4612 3453
rect 4651 3451 4685 3453
rect 4724 3451 4758 3453
rect 4797 3451 4831 3453
rect 4870 3451 4904 3453
rect 4943 3451 4977 3453
rect 5016 3451 5050 3453
rect 5089 3451 5123 3453
rect 5162 3451 5196 3453
rect 5235 3451 5269 3453
rect 5308 3451 5342 3453
rect 5381 3451 5415 3453
rect 5454 3451 5488 3453
rect 5527 3451 5561 3453
rect 5600 3451 5634 3453
rect 5673 3451 5707 3453
rect 5746 3451 5780 3453
rect 5819 3451 5853 3453
rect 5892 3451 5926 3453
rect 5965 3451 5999 3453
rect 6038 3451 6072 3453
rect 6111 3451 6145 3453
rect 6184 3451 6218 3453
rect 6257 3451 6291 3453
rect 6330 3451 7660 3453
rect 2680 3419 2714 3451
rect 2753 3419 2787 3451
rect 2826 3419 2860 3451
rect 2899 3419 2933 3451
rect 2972 3419 3006 3451
rect 3045 3419 3079 3451
rect 3118 3419 3152 3451
rect 3191 3419 3225 3451
rect 3264 3419 3298 3451
rect 3337 3419 3371 3451
rect 3410 3419 3444 3451
rect 3483 3419 3517 3451
rect 3556 3419 3590 3451
rect 3629 3419 3663 3451
rect 3702 3419 3736 3451
rect 3775 3419 3809 3451
rect 3848 3419 3882 3451
rect 3921 3419 3955 3451
rect 3994 3419 4028 3451
rect 4067 3419 4101 3451
rect 4140 3419 4174 3451
rect 4213 3419 4247 3451
rect 4286 3419 4320 3451
rect 4359 3419 4393 3451
rect 4432 3419 4466 3451
rect 4505 3419 4539 3451
rect 4578 3419 4612 3451
rect 4651 3419 4685 3451
rect 4724 3419 4758 3451
rect 4797 3419 4831 3451
rect 4870 3419 4904 3451
rect 4943 3419 4977 3451
rect 5016 3419 5050 3451
rect 5089 3419 5123 3451
rect 5162 3419 5196 3451
rect 5235 3419 5269 3451
rect 5308 3419 5342 3451
rect 5381 3419 5415 3451
rect 5454 3419 5488 3451
rect 5527 3419 5561 3451
rect 5600 3419 5634 3451
rect 5673 3419 5707 3451
rect 5746 3419 5780 3451
rect 5819 3419 5853 3451
rect 5892 3419 5926 3451
rect 5965 3419 5999 3451
rect 6038 3419 6072 3451
rect 6111 3419 6145 3451
rect 6184 3419 6218 3451
rect 6257 3419 6291 3451
rect 1950 3347 1984 3381
rect 2023 3349 2054 3381
rect 2054 3349 2057 3381
rect 2096 3349 2130 3381
rect 2169 3349 2203 3381
rect 2242 3349 2276 3381
rect 2315 3349 2349 3381
rect 2388 3349 2422 3381
rect 2461 3349 2495 3381
rect 2534 3349 2568 3381
rect 2023 3347 2057 3349
rect 2096 3347 2130 3349
rect 2169 3347 2203 3349
rect 2242 3347 2276 3349
rect 2315 3347 2349 3349
rect 2388 3347 2422 3349
rect 2461 3347 2495 3349
rect 2534 3347 2568 3349
rect 2607 3347 2641 3381
rect 2680 3349 2714 3381
rect 2753 3349 2787 3381
rect 2826 3349 2860 3381
rect 2899 3349 2933 3381
rect 2972 3349 3006 3381
rect 3045 3349 3079 3381
rect 3118 3349 3152 3381
rect 3191 3349 3225 3381
rect 3264 3349 3298 3381
rect 3337 3349 3371 3381
rect 3410 3349 3444 3381
rect 3483 3349 3517 3381
rect 3556 3349 3590 3381
rect 3629 3349 3663 3381
rect 3702 3349 3736 3381
rect 3775 3349 3809 3381
rect 3848 3349 3882 3381
rect 3921 3349 3955 3381
rect 3994 3349 4028 3381
rect 4067 3349 4101 3381
rect 4140 3349 4174 3381
rect 4213 3349 4247 3381
rect 4286 3349 4320 3381
rect 4359 3349 4393 3381
rect 4432 3349 4466 3381
rect 4505 3349 4539 3381
rect 4578 3349 4612 3381
rect 4651 3349 4685 3381
rect 4724 3349 4758 3381
rect 4797 3349 4831 3381
rect 4870 3349 4904 3381
rect 4943 3349 4977 3381
rect 5016 3349 5050 3381
rect 5089 3349 5123 3381
rect 5162 3349 5196 3381
rect 5235 3349 5269 3381
rect 5308 3349 5342 3381
rect 5381 3349 5415 3381
rect 5454 3349 5488 3381
rect 5527 3349 5561 3381
rect 5600 3349 5634 3381
rect 5673 3349 5707 3381
rect 5746 3349 5780 3381
rect 5819 3349 5853 3381
rect 5892 3349 5926 3381
rect 5965 3349 5999 3381
rect 6038 3349 6072 3381
rect 6111 3349 6145 3381
rect 6184 3349 6218 3381
rect 6257 3349 6291 3381
rect 6330 3349 7120 3451
rect 7120 3349 7235 3451
rect 7235 3349 7660 3451
rect 7733 3433 7735 3467
rect 7735 3433 7767 3467
rect 7805 3433 7837 3467
rect 7837 3433 7839 3467
rect 7733 3383 7767 3394
rect 7733 3360 7745 3383
rect 7745 3360 7767 3383
rect 7805 3360 7839 3394
rect 2680 3347 2714 3349
rect 2753 3347 2787 3349
rect 2826 3347 2860 3349
rect 2899 3347 2933 3349
rect 2972 3347 3006 3349
rect 3045 3347 3079 3349
rect 3118 3347 3152 3349
rect 3191 3347 3225 3349
rect 3264 3347 3298 3349
rect 3337 3347 3371 3349
rect 3410 3347 3444 3349
rect 3483 3347 3517 3349
rect 3556 3347 3590 3349
rect 3629 3347 3663 3349
rect 3702 3347 3736 3349
rect 3775 3347 3809 3349
rect 3848 3347 3882 3349
rect 3921 3347 3955 3349
rect 3994 3347 4028 3349
rect 4067 3347 4101 3349
rect 4140 3347 4174 3349
rect 4213 3347 4247 3349
rect 4286 3347 4320 3349
rect 4359 3347 4393 3349
rect 4432 3347 4466 3349
rect 4505 3347 4539 3349
rect 4578 3347 4612 3349
rect 4651 3347 4685 3349
rect 4724 3347 4758 3349
rect 4797 3347 4831 3349
rect 4870 3347 4904 3349
rect 4943 3347 4977 3349
rect 5016 3347 5050 3349
rect 5089 3347 5123 3349
rect 5162 3347 5196 3349
rect 5235 3347 5269 3349
rect 5308 3347 5342 3349
rect 5381 3347 5415 3349
rect 5454 3347 5488 3349
rect 5527 3347 5561 3349
rect 5600 3347 5634 3349
rect 5673 3347 5707 3349
rect 5746 3347 5780 3349
rect 5819 3347 5853 3349
rect 5892 3347 5926 3349
rect 5965 3347 5999 3349
rect 6038 3347 6072 3349
rect 6111 3347 6145 3349
rect 6184 3347 6218 3349
rect 6257 3347 6291 3349
rect 6330 3347 7660 3349
rect 1935 3015 1969 3049
rect 2008 3015 2042 3049
rect 2081 3015 2115 3049
rect 2154 3015 2188 3049
rect 2227 3015 2261 3049
rect 2300 3015 2334 3049
rect 2373 3015 2407 3049
rect 2446 3015 2480 3049
rect 2519 3015 2553 3049
rect 2592 3015 2626 3049
rect 2665 3015 2699 3049
rect 2738 3015 2772 3049
rect 2811 3015 2845 3049
rect 2884 3015 2918 3049
rect 2957 3015 2991 3049
rect 3030 3015 3064 3049
rect 3103 3015 3137 3049
rect 3176 3015 3210 3049
rect 3249 3015 3283 3049
rect 3322 3015 3356 3049
rect 3395 3015 3429 3049
rect 3468 3015 3502 3049
rect 3541 3015 3575 3049
rect 3614 3015 3648 3049
rect 3687 3015 3721 3049
rect 3760 3015 3794 3049
rect 3833 3015 3867 3049
rect 3906 3015 3940 3049
rect 3979 3015 4013 3049
rect 4052 3015 4086 3049
rect 4125 3015 4159 3049
rect 4198 3015 4232 3049
rect 4271 3015 4305 3049
rect 4344 3015 4378 3049
rect 4417 3015 4451 3049
rect 4490 3015 4524 3049
rect 4563 3015 4597 3049
rect 4636 3015 4670 3049
rect 4709 3015 4743 3049
rect 4782 3015 4816 3049
rect 4855 3015 4889 3049
rect 4928 3015 4962 3049
rect 5001 3015 5035 3049
rect 5074 3015 5108 3049
rect 5147 3015 5181 3049
rect 5220 3015 5254 3049
rect 5293 3015 5327 3049
rect 5366 3015 5400 3049
rect 5439 3015 5473 3049
rect 5511 3015 5545 3049
rect 5583 3015 5617 3049
rect 5655 3015 5689 3049
rect 5727 3015 5761 3049
rect 5799 3015 5833 3049
rect 5871 3015 5905 3049
rect 5943 3015 5977 3049
rect 6015 3015 6049 3049
rect 6087 3015 6121 3049
rect 6159 3015 6193 3049
rect 6231 3015 6265 3049
rect 6303 3015 6337 3049
rect 6375 3015 6409 3049
rect 6447 3015 6481 3049
rect 6519 3015 6553 3049
rect 6591 3015 6625 3049
rect 6663 3015 6697 3049
rect 6735 3015 6769 3049
rect 6807 3015 6841 3049
rect 6879 3015 6913 3049
rect 6951 3015 6985 3049
rect 7023 3015 7057 3049
rect 7095 3015 7129 3049
rect 7167 3015 7201 3049
rect 7239 3015 7273 3049
rect 7311 3015 7345 3049
rect 7383 3015 7417 3049
rect 7455 3015 7489 3049
rect 7527 3015 7561 3049
rect 1935 2937 1969 2971
rect 2008 2937 2042 2971
rect 2081 2937 2115 2971
rect 2154 2937 2188 2971
rect 2227 2937 2261 2971
rect 2300 2937 2334 2971
rect 2373 2937 2407 2971
rect 2446 2937 2480 2971
rect 2519 2937 2553 2971
rect 2592 2937 2626 2971
rect 2665 2937 2699 2971
rect 2738 2937 2772 2971
rect 2811 2937 2845 2971
rect 2884 2937 2918 2971
rect 2957 2937 2991 2971
rect 3030 2937 3064 2971
rect 3103 2937 3137 2971
rect 3176 2937 3210 2971
rect 3249 2937 3283 2971
rect 3322 2937 3356 2971
rect 3395 2937 3429 2971
rect 3468 2937 3502 2971
rect 3541 2937 3575 2971
rect 3614 2937 3648 2971
rect 3687 2937 3721 2971
rect 3760 2937 3794 2971
rect 3833 2937 3867 2971
rect 3906 2937 3940 2971
rect 3979 2937 4013 2971
rect 4052 2937 4086 2971
rect 4125 2937 4159 2971
rect 4198 2937 4232 2971
rect 4271 2937 4305 2971
rect 4344 2937 4378 2971
rect 4417 2937 4451 2971
rect 4490 2937 4524 2971
rect 4563 2937 4597 2971
rect 4636 2937 4670 2971
rect 4709 2937 4743 2971
rect 4782 2937 4816 2971
rect 4855 2937 4889 2971
rect 4928 2937 4962 2971
rect 5001 2937 5035 2971
rect 5074 2937 5108 2971
rect 5147 2937 5181 2971
rect 5220 2937 5254 2971
rect 5293 2937 5327 2971
rect 5366 2937 5400 2971
rect 5439 2937 5473 2971
rect 5511 2937 5545 2971
rect 5583 2937 5617 2971
rect 5655 2937 5689 2971
rect 5727 2937 5761 2971
rect 5799 2937 5833 2971
rect 5871 2937 5905 2971
rect 5943 2937 5977 2971
rect 6015 2937 6049 2971
rect 6087 2937 6121 2971
rect 6159 2937 6193 2971
rect 6231 2937 6265 2971
rect 6303 2937 6337 2971
rect 6375 2937 6409 2971
rect 6447 2937 6481 2971
rect 6519 2937 6553 2971
rect 6591 2937 6625 2971
rect 6663 2937 6697 2971
rect 6735 2937 6769 2971
rect 6807 2937 6841 2971
rect 6879 2937 6913 2971
rect 6951 2937 6985 2971
rect 7023 2937 7057 2971
rect 7095 2937 7129 2971
rect 7167 2937 7201 2971
rect 7239 2937 7273 2971
rect 7311 2937 7345 2971
rect 7383 2937 7417 2971
rect 7455 2937 7489 2971
rect 7527 2937 7561 2971
rect 1935 2859 1969 2893
rect 2008 2860 2026 2893
rect 2026 2860 2042 2893
rect 2008 2859 2042 2860
rect 2081 2859 2115 2893
rect 2154 2860 2163 2893
rect 2163 2860 2188 2893
rect 2154 2859 2188 2860
rect 2227 2859 2261 2893
rect 2300 2859 2334 2893
rect 2373 2860 2403 2893
rect 2403 2860 2407 2893
rect 2373 2859 2407 2860
rect 2446 2859 2480 2893
rect 2519 2860 2540 2893
rect 2540 2860 2553 2893
rect 2519 2859 2553 2860
rect 2592 2859 2626 2893
rect 2665 2860 2677 2893
rect 2677 2860 2699 2893
rect 2665 2859 2699 2860
rect 2738 2859 2772 2893
rect 2811 2860 2814 2893
rect 2814 2860 2845 2893
rect 2811 2859 2845 2860
rect 2884 2859 2918 2893
rect 2957 2860 2984 2893
rect 2984 2860 2991 2893
rect 2957 2859 2991 2860
rect 3030 2859 3064 2893
rect 3103 2860 3120 2893
rect 3120 2860 3137 2893
rect 3103 2859 3137 2860
rect 3176 2859 3210 2893
rect 3249 2860 3256 2893
rect 3256 2860 3283 2893
rect 3249 2859 3283 2860
rect 3322 2859 3356 2893
rect 3395 2859 3429 2893
rect 3468 2860 3494 2893
rect 3494 2860 3502 2893
rect 3468 2859 3502 2860
rect 3541 2859 3575 2893
rect 3614 2860 3630 2893
rect 3630 2860 3648 2893
rect 3614 2859 3648 2860
rect 3687 2859 3721 2893
rect 3760 2860 3766 2893
rect 3766 2860 3794 2893
rect 3760 2859 3794 2860
rect 3833 2859 3867 2893
rect 3906 2860 3936 2893
rect 3936 2860 3940 2893
rect 3906 2859 3940 2860
rect 3979 2859 4013 2893
rect 4052 2860 4072 2893
rect 4072 2860 4086 2893
rect 4052 2859 4086 2860
rect 4125 2859 4159 2893
rect 4198 2860 4208 2893
rect 4208 2860 4232 2893
rect 4198 2859 4232 2860
rect 4271 2859 4305 2893
rect 4344 2859 4378 2893
rect 4417 2860 4446 2893
rect 4446 2860 4451 2893
rect 4417 2859 4451 2860
rect 4490 2859 4524 2893
rect 4563 2860 4582 2893
rect 4582 2860 4597 2893
rect 4563 2859 4597 2860
rect 4636 2859 4670 2893
rect 4709 2860 4718 2893
rect 4718 2860 4743 2893
rect 4709 2859 4743 2860
rect 4782 2859 4816 2893
rect 4855 2860 4888 2893
rect 4888 2860 4889 2893
rect 4855 2859 4889 2860
rect 4928 2859 4962 2893
rect 5001 2860 5024 2893
rect 5024 2860 5035 2893
rect 5001 2859 5035 2860
rect 5074 2859 5108 2893
rect 5147 2860 5160 2893
rect 5160 2860 5181 2893
rect 5147 2859 5181 2860
rect 5220 2859 5254 2893
rect 5293 2860 5296 2893
rect 5296 2860 5327 2893
rect 5293 2859 5327 2860
rect 5366 2860 5398 2893
rect 5398 2860 5400 2893
rect 5366 2859 5400 2860
rect 5439 2859 5473 2893
rect 5511 2860 5534 2893
rect 5534 2860 5545 2893
rect 5511 2859 5545 2860
rect 5583 2859 5617 2893
rect 5655 2860 5670 2893
rect 5670 2860 5689 2893
rect 5655 2859 5689 2860
rect 5727 2859 5761 2893
rect 5799 2860 5806 2893
rect 5806 2860 5833 2893
rect 5799 2859 5833 2860
rect 5871 2859 5905 2893
rect 5943 2860 5976 2893
rect 5976 2860 5977 2893
rect 5943 2859 5977 2860
rect 6015 2859 6049 2893
rect 6087 2860 6112 2893
rect 6112 2860 6121 2893
rect 6087 2859 6121 2860
rect 6159 2859 6193 2893
rect 6231 2860 6248 2893
rect 6248 2860 6265 2893
rect 6231 2859 6265 2860
rect 6303 2859 6337 2893
rect 6375 2860 6384 2893
rect 6384 2860 6409 2893
rect 6375 2859 6409 2860
rect 6447 2859 6481 2893
rect 6519 2860 6520 2893
rect 6520 2860 6553 2893
rect 6519 2859 6553 2860
rect 6591 2860 6622 2893
rect 6622 2860 6625 2893
rect 6591 2859 6625 2860
rect 6663 2859 6697 2893
rect 6735 2860 6758 2893
rect 6758 2860 6769 2893
rect 6735 2859 6769 2860
rect 6807 2859 6841 2893
rect 6879 2860 6894 2893
rect 6894 2860 6913 2893
rect 6879 2859 6913 2860
rect 6951 2859 6985 2893
rect 7023 2860 7030 2893
rect 7030 2860 7057 2893
rect 7023 2859 7057 2860
rect 7095 2859 7129 2893
rect 7167 2860 7200 2893
rect 7200 2860 7201 2893
rect 7167 2859 7201 2860
rect 7239 2859 7273 2893
rect 7311 2860 7336 2893
rect 7336 2860 7345 2893
rect 7311 2859 7345 2860
rect 7383 2859 7417 2893
rect 7455 2860 7472 2893
rect 7472 2860 7489 2893
rect 7455 2859 7489 2860
rect 7527 2859 7561 2893
rect 1935 2781 1969 2815
rect 2008 2781 2042 2815
rect 2081 2781 2115 2815
rect 2154 2781 2188 2815
rect 2227 2781 2261 2815
rect 2300 2781 2334 2815
rect 2373 2781 2407 2815
rect 2446 2781 2480 2815
rect 2519 2781 2553 2815
rect 2592 2781 2626 2815
rect 2665 2781 2699 2815
rect 2738 2781 2772 2815
rect 2811 2781 2845 2815
rect 2884 2781 2918 2815
rect 2957 2781 2991 2815
rect 3030 2781 3064 2815
rect 3103 2781 3137 2815
rect 3176 2781 3210 2815
rect 3249 2781 3283 2815
rect 3322 2781 3356 2815
rect 3395 2781 3429 2815
rect 3468 2781 3502 2815
rect 3541 2781 3575 2815
rect 3614 2781 3648 2815
rect 3687 2781 3721 2815
rect 3760 2781 3794 2815
rect 3833 2781 3867 2815
rect 3906 2781 3940 2815
rect 3979 2781 4013 2815
rect 4052 2781 4086 2815
rect 4125 2781 4159 2815
rect 4198 2781 4232 2815
rect 4271 2781 4305 2815
rect 4344 2781 4378 2815
rect 4417 2781 4451 2815
rect 4490 2781 4524 2815
rect 4563 2781 4597 2815
rect 4636 2781 4670 2815
rect 4709 2781 4743 2815
rect 4782 2781 4816 2815
rect 4855 2781 4889 2815
rect 4928 2781 4962 2815
rect 5001 2781 5035 2815
rect 5074 2781 5108 2815
rect 5147 2781 5181 2815
rect 5220 2781 5254 2815
rect 5293 2781 5327 2815
rect 5366 2781 5400 2815
rect 5439 2781 5473 2815
rect 5511 2781 5545 2815
rect 5583 2781 5617 2815
rect 5655 2781 5689 2815
rect 5727 2781 5761 2815
rect 5799 2781 5833 2815
rect 5871 2781 5905 2815
rect 5943 2781 5977 2815
rect 6015 2781 6049 2815
rect 6087 2781 6121 2815
rect 6159 2781 6193 2815
rect 6231 2781 6265 2815
rect 6303 2781 6337 2815
rect 6375 2781 6409 2815
rect 6447 2781 6481 2815
rect 6519 2781 6553 2815
rect 6591 2781 6625 2815
rect 6663 2781 6697 2815
rect 6735 2781 6769 2815
rect 6807 2781 6841 2815
rect 6879 2781 6913 2815
rect 6951 2781 6985 2815
rect 7023 2781 7057 2815
rect 7095 2781 7129 2815
rect 7167 2781 7201 2815
rect 7239 2781 7273 2815
rect 7311 2781 7345 2815
rect 7383 2781 7417 2815
rect 7455 2781 7489 2815
rect 7527 2781 7561 2815
rect 1935 2703 1969 2737
rect 2008 2703 2042 2737
rect 2081 2703 2115 2737
rect 2154 2703 2188 2737
rect 2227 2703 2261 2737
rect 2300 2703 2334 2737
rect 2373 2703 2407 2737
rect 2446 2703 2480 2737
rect 2519 2703 2553 2737
rect 2592 2703 2626 2737
rect 2665 2703 2699 2737
rect 2738 2703 2772 2737
rect 2811 2703 2845 2737
rect 2884 2703 2918 2737
rect 2957 2703 2991 2737
rect 3030 2703 3064 2737
rect 3103 2703 3137 2737
rect 3176 2703 3210 2737
rect 3249 2703 3283 2737
rect 3322 2703 3356 2737
rect 3395 2703 3429 2737
rect 3468 2703 3502 2737
rect 3541 2703 3575 2737
rect 3614 2703 3648 2737
rect 3687 2703 3721 2737
rect 3760 2703 3794 2737
rect 3833 2703 3867 2737
rect 3906 2703 3940 2737
rect 3979 2703 4013 2737
rect 4052 2703 4086 2737
rect 4125 2703 4159 2737
rect 4198 2703 4232 2737
rect 4271 2703 4305 2737
rect 4344 2703 4378 2737
rect 4417 2703 4451 2737
rect 4490 2703 4524 2737
rect 4563 2703 4597 2737
rect 4636 2703 4670 2737
rect 4709 2703 4743 2737
rect 4782 2703 4816 2737
rect 4855 2703 4889 2737
rect 4928 2703 4962 2737
rect 5001 2703 5035 2737
rect 5074 2703 5108 2737
rect 5147 2703 5181 2737
rect 5220 2703 5254 2737
rect 5293 2703 5327 2737
rect 5366 2703 5400 2737
rect 5439 2703 5473 2737
rect 5511 2703 5545 2737
rect 5583 2703 5617 2737
rect 5655 2703 5689 2737
rect 5727 2703 5761 2737
rect 5799 2703 5833 2737
rect 5871 2703 5905 2737
rect 5943 2703 5977 2737
rect 6015 2703 6049 2737
rect 6087 2703 6121 2737
rect 6159 2703 6193 2737
rect 6231 2703 6265 2737
rect 6303 2703 6337 2737
rect 6375 2703 6409 2737
rect 6447 2703 6481 2737
rect 6519 2703 6553 2737
rect 6591 2703 6625 2737
rect 6663 2703 6697 2737
rect 6735 2703 6769 2737
rect 6807 2703 6841 2737
rect 6879 2703 6913 2737
rect 6951 2703 6985 2737
rect 7023 2703 7057 2737
rect 7095 2703 7129 2737
rect 7167 2703 7201 2737
rect 7239 2703 7273 2737
rect 7311 2703 7345 2737
rect 7383 2703 7417 2737
rect 7455 2703 7489 2737
rect 7527 2703 7561 2737
rect 1935 2625 1969 2659
rect 2008 2628 2026 2659
rect 2026 2628 2042 2659
rect 2008 2625 2042 2628
rect 2081 2625 2115 2659
rect 2154 2628 2163 2659
rect 2163 2628 2188 2659
rect 2154 2625 2188 2628
rect 2227 2625 2261 2659
rect 2300 2625 2334 2659
rect 2373 2628 2403 2659
rect 2403 2628 2407 2659
rect 2373 2625 2407 2628
rect 2446 2625 2480 2659
rect 2519 2628 2540 2659
rect 2540 2628 2553 2659
rect 2519 2625 2553 2628
rect 2592 2625 2626 2659
rect 2665 2628 2677 2659
rect 2677 2628 2699 2659
rect 2665 2625 2699 2628
rect 2738 2625 2772 2659
rect 2811 2628 2814 2659
rect 2814 2628 2845 2659
rect 2811 2625 2845 2628
rect 2884 2625 2918 2659
rect 2957 2628 2984 2659
rect 2984 2628 2991 2659
rect 2957 2625 2991 2628
rect 3030 2625 3064 2659
rect 3103 2628 3120 2659
rect 3120 2628 3137 2659
rect 3103 2625 3137 2628
rect 3176 2625 3210 2659
rect 3249 2628 3256 2659
rect 3256 2628 3283 2659
rect 3249 2625 3283 2628
rect 3322 2625 3356 2659
rect 3395 2625 3429 2659
rect 3468 2628 3494 2659
rect 3494 2628 3502 2659
rect 3468 2625 3502 2628
rect 3541 2625 3575 2659
rect 3614 2628 3630 2659
rect 3630 2628 3648 2659
rect 3614 2625 3648 2628
rect 3687 2625 3721 2659
rect 3760 2628 3766 2659
rect 3766 2628 3794 2659
rect 3760 2625 3794 2628
rect 3833 2625 3867 2659
rect 3906 2628 3936 2659
rect 3936 2628 3940 2659
rect 3906 2625 3940 2628
rect 3979 2625 4013 2659
rect 4052 2628 4072 2659
rect 4072 2628 4086 2659
rect 4052 2625 4086 2628
rect 4125 2625 4159 2659
rect 4198 2628 4208 2659
rect 4208 2628 4232 2659
rect 4198 2625 4232 2628
rect 4271 2625 4305 2659
rect 4344 2625 4378 2659
rect 4417 2628 4446 2659
rect 4446 2628 4451 2659
rect 4417 2625 4451 2628
rect 4490 2625 4524 2659
rect 4563 2628 4582 2659
rect 4582 2628 4597 2659
rect 4563 2625 4597 2628
rect 4636 2625 4670 2659
rect 4709 2628 4718 2659
rect 4718 2628 4743 2659
rect 4709 2625 4743 2628
rect 4782 2625 4816 2659
rect 4855 2628 4888 2659
rect 4888 2628 4889 2659
rect 4855 2625 4889 2628
rect 4928 2625 4962 2659
rect 5001 2628 5024 2659
rect 5024 2628 5035 2659
rect 5001 2625 5035 2628
rect 5074 2625 5108 2659
rect 5147 2628 5160 2659
rect 5160 2628 5181 2659
rect 5147 2625 5181 2628
rect 5220 2625 5254 2659
rect 5293 2628 5296 2659
rect 5296 2628 5327 2659
rect 5293 2625 5327 2628
rect 5366 2628 5398 2659
rect 5398 2628 5400 2659
rect 5366 2625 5400 2628
rect 5439 2625 5473 2659
rect 5511 2628 5534 2659
rect 5534 2628 5545 2659
rect 5511 2625 5545 2628
rect 5583 2625 5617 2659
rect 5655 2628 5670 2659
rect 5670 2628 5689 2659
rect 5655 2625 5689 2628
rect 5727 2625 5761 2659
rect 5799 2628 5806 2659
rect 5806 2628 5833 2659
rect 5799 2625 5833 2628
rect 5871 2625 5905 2659
rect 5943 2628 5976 2659
rect 5976 2628 5977 2659
rect 5943 2625 5977 2628
rect 6015 2625 6049 2659
rect 6087 2628 6112 2659
rect 6112 2628 6121 2659
rect 6087 2625 6121 2628
rect 6159 2625 6193 2659
rect 6231 2628 6248 2659
rect 6248 2628 6265 2659
rect 6231 2625 6265 2628
rect 6303 2625 6337 2659
rect 6375 2628 6384 2659
rect 6384 2628 6409 2659
rect 6375 2625 6409 2628
rect 6447 2625 6481 2659
rect 6519 2628 6520 2659
rect 6520 2628 6553 2659
rect 6519 2625 6553 2628
rect 6591 2628 6622 2659
rect 6622 2628 6625 2659
rect 6591 2625 6625 2628
rect 6663 2625 6697 2659
rect 6735 2628 6758 2659
rect 6758 2628 6769 2659
rect 6735 2625 6769 2628
rect 6807 2625 6841 2659
rect 6879 2628 6894 2659
rect 6894 2628 6913 2659
rect 6879 2625 6913 2628
rect 6951 2625 6985 2659
rect 7023 2628 7030 2659
rect 7030 2628 7057 2659
rect 7023 2625 7057 2628
rect 7095 2625 7129 2659
rect 7167 2628 7200 2659
rect 7200 2628 7201 2659
rect 7167 2625 7201 2628
rect 7239 2625 7273 2659
rect 7311 2628 7336 2659
rect 7336 2628 7345 2659
rect 7311 2625 7345 2628
rect 7383 2625 7417 2659
rect 7455 2628 7472 2659
rect 7472 2628 7489 2659
rect 7455 2625 7489 2628
rect 7527 2625 7561 2659
rect 1935 2547 1969 2581
rect 2008 2547 2042 2581
rect 2081 2547 2115 2581
rect 2154 2547 2188 2581
rect 2227 2547 2261 2581
rect 2300 2547 2334 2581
rect 2373 2547 2407 2581
rect 2446 2547 2480 2581
rect 2519 2547 2553 2581
rect 2592 2547 2626 2581
rect 2665 2547 2699 2581
rect 2738 2547 2772 2581
rect 2811 2547 2845 2581
rect 2884 2547 2918 2581
rect 2957 2547 2991 2581
rect 3030 2547 3064 2581
rect 3103 2547 3137 2581
rect 3176 2547 3210 2581
rect 3249 2547 3283 2581
rect 3322 2547 3356 2581
rect 3395 2547 3429 2581
rect 3468 2547 3502 2581
rect 3541 2547 3575 2581
rect 3614 2547 3648 2581
rect 3687 2547 3721 2581
rect 3760 2547 3794 2581
rect 3833 2547 3867 2581
rect 3906 2547 3940 2581
rect 3979 2547 4013 2581
rect 4052 2547 4086 2581
rect 4125 2547 4159 2581
rect 4198 2547 4232 2581
rect 4271 2547 4305 2581
rect 4344 2547 4378 2581
rect 4417 2547 4451 2581
rect 4490 2547 4524 2581
rect 4563 2547 4597 2581
rect 4636 2547 4670 2581
rect 4709 2547 4743 2581
rect 4782 2547 4816 2581
rect 4855 2547 4889 2581
rect 4928 2547 4962 2581
rect 5001 2547 5035 2581
rect 5074 2547 5108 2581
rect 5147 2547 5181 2581
rect 5220 2547 5254 2581
rect 5293 2547 5327 2581
rect 5366 2547 5400 2581
rect 5439 2547 5473 2581
rect 5511 2547 5545 2581
rect 5583 2547 5617 2581
rect 5655 2547 5689 2581
rect 5727 2547 5761 2581
rect 5799 2547 5833 2581
rect 5871 2547 5905 2581
rect 5943 2547 5977 2581
rect 6015 2547 6049 2581
rect 6087 2547 6121 2581
rect 6159 2547 6193 2581
rect 6231 2547 6265 2581
rect 6303 2547 6337 2581
rect 6375 2547 6409 2581
rect 6447 2547 6481 2581
rect 6519 2547 6553 2581
rect 6591 2547 6625 2581
rect 6663 2547 6697 2581
rect 6735 2547 6769 2581
rect 6807 2547 6841 2581
rect 6879 2547 6913 2581
rect 6951 2547 6985 2581
rect 7023 2547 7057 2581
rect 7095 2547 7129 2581
rect 7167 2547 7201 2581
rect 7239 2547 7273 2581
rect 7311 2547 7345 2581
rect 7383 2547 7417 2581
rect 7455 2547 7489 2581
rect 7527 2547 7561 2581
rect 1935 2469 1969 2503
rect 2008 2469 2042 2503
rect 2081 2469 2115 2503
rect 2154 2469 2188 2503
rect 2227 2469 2261 2503
rect 2300 2469 2334 2503
rect 2373 2469 2407 2503
rect 2446 2469 2480 2503
rect 2519 2469 2553 2503
rect 2592 2469 2626 2503
rect 2665 2469 2699 2503
rect 2738 2469 2772 2503
rect 2811 2469 2845 2503
rect 2884 2469 2918 2503
rect 2957 2469 2991 2503
rect 3030 2469 3064 2503
rect 3103 2469 3137 2503
rect 3176 2469 3210 2503
rect 3249 2469 3283 2503
rect 3322 2469 3356 2503
rect 3395 2469 3429 2503
rect 3468 2469 3502 2503
rect 3541 2469 3575 2503
rect 3614 2469 3648 2503
rect 3687 2469 3721 2503
rect 3760 2469 3794 2503
rect 3833 2469 3867 2503
rect 3906 2469 3940 2503
rect 3979 2469 4013 2503
rect 4052 2469 4086 2503
rect 4125 2469 4159 2503
rect 4198 2469 4232 2503
rect 4271 2469 4305 2503
rect 4344 2469 4378 2503
rect 4417 2469 4451 2503
rect 4490 2469 4524 2503
rect 4563 2469 4597 2503
rect 4636 2469 4670 2503
rect 4709 2469 4743 2503
rect 4782 2469 4816 2503
rect 4855 2469 4889 2503
rect 4928 2469 4962 2503
rect 5001 2469 5035 2503
rect 5074 2469 5108 2503
rect 5147 2469 5181 2503
rect 5220 2469 5254 2503
rect 5293 2469 5327 2503
rect 5366 2469 5400 2503
rect 5439 2469 5473 2503
rect 5511 2469 5545 2503
rect 5583 2469 5617 2503
rect 5655 2469 5689 2503
rect 5727 2469 5761 2503
rect 5799 2469 5833 2503
rect 5871 2469 5905 2503
rect 5943 2469 5977 2503
rect 6015 2469 6049 2503
rect 6087 2469 6121 2503
rect 6159 2469 6193 2503
rect 6231 2469 6265 2503
rect 6303 2469 6337 2503
rect 6375 2469 6409 2503
rect 6447 2469 6481 2503
rect 6519 2469 6553 2503
rect 6591 2469 6625 2503
rect 6663 2469 6697 2503
rect 6735 2469 6769 2503
rect 6807 2469 6841 2503
rect 6879 2469 6913 2503
rect 6951 2469 6985 2503
rect 7023 2469 7057 2503
rect 7095 2469 7129 2503
rect 7167 2469 7201 2503
rect 7239 2469 7273 2503
rect 7311 2469 7345 2503
rect 7383 2469 7417 2503
rect 7455 2469 7489 2503
rect 7527 2469 7561 2503
rect 5414 2235 5448 2269
rect 5486 2235 5520 2269
rect 5558 2235 5592 2269
rect 5630 2235 5664 2269
rect 5702 2235 5736 2269
rect 5774 2235 5808 2269
rect 5846 2235 5880 2269
rect 5918 2235 5952 2269
rect 5990 2235 6024 2269
rect 6062 2235 6096 2269
rect 6134 2235 6168 2269
rect 6206 2235 6240 2269
rect 6278 2235 6312 2269
rect 6350 2235 6384 2269
rect 6595 2235 6629 2269
rect 6667 2235 6701 2269
rect 6739 2235 6773 2269
rect 6811 2235 6845 2269
rect 6883 2235 6917 2269
rect 6955 2235 6989 2269
rect 7027 2235 7061 2269
rect 7099 2235 7133 2269
rect 7171 2235 7205 2269
rect 7243 2235 7277 2269
rect 7315 2235 7349 2269
rect 7387 2235 7421 2269
rect 7459 2235 7493 2269
rect 7531 2235 7565 2269
rect 5414 2161 5448 2195
rect 5486 2189 5518 2195
rect 5518 2189 5520 2195
rect 5486 2161 5520 2189
rect 5558 2161 5592 2195
rect 5630 2189 5656 2195
rect 5656 2189 5664 2195
rect 5630 2161 5664 2189
rect 5702 2161 5736 2195
rect 5774 2189 5794 2195
rect 5794 2189 5808 2195
rect 5774 2161 5808 2189
rect 5846 2161 5880 2195
rect 5918 2189 5932 2195
rect 5932 2189 5952 2195
rect 5918 2161 5952 2189
rect 5990 2161 6024 2195
rect 6062 2189 6070 2195
rect 6070 2189 6096 2195
rect 6062 2161 6096 2189
rect 6134 2161 6168 2195
rect 6206 2189 6208 2195
rect 6208 2189 6240 2195
rect 6206 2161 6240 2189
rect 6278 2161 6312 2195
rect 6350 2161 6384 2195
rect 6595 2189 6622 2195
rect 6622 2189 6629 2195
rect 6595 2161 6629 2189
rect 6667 2161 6701 2195
rect 6739 2189 6760 2195
rect 6760 2189 6773 2195
rect 6739 2161 6773 2189
rect 6811 2161 6845 2195
rect 6883 2189 6898 2195
rect 6898 2189 6917 2195
rect 6883 2161 6917 2189
rect 6955 2161 6989 2195
rect 7027 2189 7036 2195
rect 7036 2189 7061 2195
rect 7027 2161 7061 2189
rect 7099 2161 7133 2195
rect 7171 2189 7174 2195
rect 7174 2189 7205 2195
rect 7171 2161 7205 2189
rect 7243 2161 7277 2195
rect 7315 2161 7349 2195
rect 7387 2189 7416 2195
rect 7416 2189 7421 2195
rect 7387 2161 7421 2189
rect 7459 2161 7493 2195
rect 7531 2189 7554 2195
rect 7554 2189 7565 2195
rect 7531 2161 7565 2189
rect 5414 2087 5448 2121
rect 5486 2087 5520 2121
rect 5558 2087 5592 2121
rect 5630 2087 5664 2121
rect 5702 2087 5736 2121
rect 5774 2087 5808 2121
rect 5846 2087 5880 2121
rect 5918 2087 5952 2121
rect 5990 2087 6024 2121
rect 6062 2087 6096 2121
rect 6134 2087 6168 2121
rect 6206 2087 6240 2121
rect 6278 2087 6312 2121
rect 6350 2087 6384 2121
rect 6595 2087 6629 2121
rect 6667 2087 6701 2121
rect 6739 2087 6773 2121
rect 6811 2087 6845 2121
rect 6883 2087 6917 2121
rect 6955 2087 6989 2121
rect 7027 2087 7061 2121
rect 7099 2087 7133 2121
rect 7171 2087 7205 2121
rect 7243 2087 7277 2121
rect 7315 2087 7349 2121
rect 7387 2087 7421 2121
rect 7459 2087 7493 2121
rect 7531 2087 7565 2121
rect 2253 1982 2277 2016
rect 2277 1982 2287 2016
rect 2326 1982 2345 2016
rect 2345 1982 2360 2016
rect 2399 1982 2413 2016
rect 2413 1982 2433 2016
rect 2472 1982 2481 2016
rect 2481 1982 2506 2016
rect 2545 1982 2549 2016
rect 2549 1982 2579 2016
rect 2618 1982 2651 2016
rect 2651 1982 2652 2016
rect 2691 1982 2719 2016
rect 2719 1982 2725 2016
rect 2764 1982 2787 2016
rect 2787 1982 2798 2016
rect 2837 1982 2855 2016
rect 2855 1982 2871 2016
rect 2910 1982 2923 2016
rect 2923 1982 2944 2016
rect 2983 1982 2991 2016
rect 2991 1982 3017 2016
rect 3056 1982 3059 2016
rect 3059 1982 3090 2016
rect 3129 1982 3161 2016
rect 3161 1982 3163 2016
rect 3202 1982 3229 2016
rect 3229 1982 3236 2016
rect 3275 1982 3297 2016
rect 3297 1982 3309 2016
rect 3348 1982 3365 2016
rect 3365 1982 3382 2016
rect 3421 1982 3433 2016
rect 3433 1982 3455 2016
rect 3493 1982 3501 2016
rect 3501 1982 3527 2016
rect 3565 1982 3569 2016
rect 3569 1982 3599 2016
rect 3637 1982 3671 2016
rect 3709 1982 3739 2016
rect 3739 1982 3743 2016
rect 3781 1982 3807 2016
rect 3807 1982 3815 2016
rect 3853 1982 3875 2016
rect 3875 1982 3887 2016
rect 3925 1982 3943 2016
rect 3943 1982 3959 2016
rect 3997 1982 4011 2016
rect 4011 1982 4031 2016
rect 4069 1982 4079 2016
rect 4079 1982 4103 2016
rect 4141 1982 4147 2016
rect 4147 1982 4175 2016
rect 4213 1982 4215 2016
rect 4215 1982 4247 2016
rect 4285 1982 4317 2016
rect 4317 1982 4319 2016
rect 4357 1982 4385 2016
rect 4385 1982 4391 2016
rect 4429 1982 4453 2016
rect 4453 1982 4463 2016
rect 4501 1982 4521 2016
rect 4521 1982 4535 2016
rect 4573 1982 4589 2016
rect 4589 1982 4607 2016
rect 4645 1982 4657 2016
rect 4657 1982 4679 2016
rect 4717 1982 4725 2016
rect 4725 1982 4751 2016
rect 4789 1982 4793 2016
rect 4793 1982 4823 2016
rect 4861 1982 4895 2016
rect 4933 1982 4963 2016
rect 4963 1982 4967 2016
rect 2009 1883 2043 1917
rect 2084 1883 2118 1917
rect 2159 1883 2193 1917
rect 2234 1883 2268 1917
rect 2309 1883 2343 1917
rect 2384 1883 2418 1917
rect 2459 1883 2493 1917
rect 2534 1883 2568 1917
rect 2609 1883 2643 1917
rect 2684 1883 2718 1917
rect 2759 1883 2793 1917
rect 2834 1883 2868 1917
rect 2909 1883 2943 1917
rect 2984 1883 3018 1917
rect 3059 1883 3093 1917
rect 3133 1883 3167 1917
rect 3207 1883 3241 1917
rect 3281 1883 3315 1917
rect 3355 1883 3389 1917
rect 3539 1883 3573 1917
rect 3614 1883 3648 1917
rect 3689 1883 3723 1917
rect 3764 1883 3798 1917
rect 3839 1883 3873 1917
rect 3914 1883 3948 1917
rect 3989 1883 4023 1917
rect 4064 1883 4098 1917
rect 4139 1883 4173 1917
rect 4214 1883 4248 1917
rect 4289 1883 4323 1917
rect 4364 1883 4398 1917
rect 4439 1883 4473 1917
rect 4514 1883 4548 1917
rect 4589 1883 4623 1917
rect 4663 1883 4697 1917
rect 4737 1883 4771 1917
rect 4811 1883 4845 1917
rect 4885 1883 4919 1917
rect 5005 1914 5039 1944
rect 5005 1910 5039 1914
rect 1919 1856 1953 1860
rect 1919 1826 1953 1856
rect 2095 1791 2129 1825
rect 2170 1791 2204 1825
rect 2245 1791 2279 1825
rect 2319 1791 2353 1825
rect 2393 1791 2427 1825
rect 2467 1791 2501 1825
rect 2541 1791 2575 1825
rect 2615 1791 2649 1825
rect 2689 1791 2723 1825
rect 2763 1791 2797 1825
rect 2837 1791 2871 1825
rect 2911 1791 2945 1825
rect 2985 1791 3019 1825
rect 3059 1791 3093 1825
rect 3133 1791 3167 1825
rect 3207 1791 3241 1825
rect 3281 1791 3315 1825
rect 3355 1791 3389 1825
rect 5005 1846 5039 1869
rect 5005 1835 5039 1846
rect 1919 1784 1953 1787
rect 1919 1753 1953 1784
rect 3625 1791 3659 1825
rect 3699 1791 3733 1825
rect 3773 1791 3807 1825
rect 3847 1791 3881 1825
rect 3921 1791 3955 1825
rect 3994 1791 4028 1825
rect 4067 1791 4101 1825
rect 4140 1791 4174 1825
rect 4213 1791 4247 1825
rect 4286 1791 4320 1825
rect 4359 1791 4393 1825
rect 4432 1791 4466 1825
rect 4505 1791 4539 1825
rect 4578 1791 4612 1825
rect 4651 1791 4685 1825
rect 1919 1712 1953 1714
rect 1919 1680 1953 1712
rect 2241 1699 2275 1733
rect 2316 1699 2350 1733
rect 2391 1699 2425 1733
rect 2466 1699 2500 1733
rect 2541 1699 2575 1733
rect 2615 1699 2649 1733
rect 2689 1699 2723 1733
rect 2763 1699 2797 1733
rect 2837 1699 2871 1733
rect 2911 1699 2945 1733
rect 2985 1699 3019 1733
rect 3059 1699 3093 1733
rect 3133 1699 3167 1733
rect 3207 1699 3241 1733
rect 3281 1699 3315 1733
rect 3355 1699 3389 1733
rect 5005 1778 5039 1794
rect 5005 1760 5039 1778
rect 3539 1699 3573 1733
rect 3614 1699 3648 1733
rect 3689 1699 3723 1733
rect 3764 1699 3798 1733
rect 3839 1699 3873 1733
rect 3914 1699 3948 1733
rect 3989 1699 4023 1733
rect 4064 1699 4098 1733
rect 4139 1699 4173 1733
rect 4214 1699 4248 1733
rect 4289 1699 4323 1733
rect 4364 1699 4398 1733
rect 4439 1699 4473 1733
rect 4514 1699 4548 1733
rect 4589 1699 4623 1733
rect 4663 1699 4697 1733
rect 4737 1699 4771 1733
rect 4811 1699 4845 1733
rect 4885 1699 4919 1733
rect 5005 1710 5039 1719
rect 1919 1640 1953 1641
rect 1919 1607 1953 1640
rect 2095 1607 2129 1641
rect 2170 1607 2204 1641
rect 2245 1607 2279 1641
rect 2319 1607 2353 1641
rect 2393 1607 2427 1641
rect 2467 1607 2501 1641
rect 2541 1607 2575 1641
rect 2615 1607 2649 1641
rect 2689 1607 2723 1641
rect 2763 1607 2797 1641
rect 2837 1607 2871 1641
rect 2911 1607 2945 1641
rect 2985 1607 3019 1641
rect 3059 1607 3093 1641
rect 3133 1607 3167 1641
rect 3207 1607 3241 1641
rect 3281 1607 3315 1641
rect 3355 1607 3389 1641
rect 5005 1685 5039 1710
rect 5005 1642 5039 1644
rect 1919 1534 1953 1568
rect 3625 1607 3659 1641
rect 3699 1607 3733 1641
rect 3773 1607 3807 1641
rect 3847 1607 3881 1641
rect 3921 1607 3955 1641
rect 3994 1607 4028 1641
rect 4067 1607 4101 1641
rect 4140 1607 4174 1641
rect 4213 1607 4247 1641
rect 4286 1607 4320 1641
rect 4359 1607 4393 1641
rect 4432 1607 4466 1641
rect 4505 1607 4539 1641
rect 4578 1607 4612 1641
rect 4651 1607 4685 1641
rect 5005 1610 5039 1642
rect 2241 1515 2275 1549
rect 2316 1515 2350 1549
rect 2391 1515 2425 1549
rect 2466 1515 2500 1549
rect 2541 1515 2575 1549
rect 2615 1515 2649 1549
rect 2689 1515 2723 1549
rect 2763 1515 2797 1549
rect 2837 1515 2871 1549
rect 2911 1515 2945 1549
rect 2985 1515 3019 1549
rect 3059 1515 3093 1549
rect 3133 1515 3167 1549
rect 3207 1515 3241 1549
rect 3281 1515 3315 1549
rect 3355 1515 3389 1549
rect 1919 1462 1953 1495
rect 1919 1461 1953 1462
rect 3539 1515 3573 1549
rect 3614 1515 3648 1549
rect 3689 1515 3723 1549
rect 3764 1515 3798 1549
rect 3839 1515 3873 1549
rect 3914 1515 3948 1549
rect 3989 1515 4023 1549
rect 4064 1515 4098 1549
rect 4139 1515 4173 1549
rect 4214 1515 4248 1549
rect 4289 1515 4323 1549
rect 4364 1515 4398 1549
rect 4439 1515 4473 1549
rect 4514 1515 4548 1549
rect 4589 1515 4623 1549
rect 4663 1515 4697 1549
rect 4737 1515 4771 1549
rect 4811 1515 4845 1549
rect 4885 1515 4919 1549
rect 5005 1540 5039 1569
rect 5005 1535 5039 1540
rect 2095 1423 2129 1457
rect 2170 1423 2204 1457
rect 2245 1423 2279 1457
rect 2319 1423 2353 1457
rect 2393 1423 2427 1457
rect 2467 1423 2501 1457
rect 2541 1423 2575 1457
rect 2615 1423 2649 1457
rect 2689 1423 2723 1457
rect 2763 1423 2797 1457
rect 2837 1423 2871 1457
rect 2911 1423 2945 1457
rect 2985 1423 3019 1457
rect 3059 1423 3093 1457
rect 3133 1423 3167 1457
rect 3207 1423 3241 1457
rect 3281 1423 3315 1457
rect 3355 1423 3389 1457
rect 5005 1472 5039 1494
rect 5005 1460 5039 1472
rect 3625 1423 3659 1457
rect 3699 1423 3733 1457
rect 3773 1423 3807 1457
rect 3847 1423 3881 1457
rect 3921 1423 3955 1457
rect 3994 1423 4028 1457
rect 4067 1423 4101 1457
rect 4140 1423 4174 1457
rect 4213 1423 4247 1457
rect 4286 1423 4320 1457
rect 4359 1423 4393 1457
rect 4432 1423 4466 1457
rect 4505 1423 4539 1457
rect 4578 1423 4612 1457
rect 4651 1423 4685 1457
rect 1919 1389 1953 1422
rect 1919 1388 1953 1389
rect 1919 1316 1953 1349
rect 2241 1331 2275 1365
rect 2316 1331 2350 1365
rect 2391 1331 2425 1365
rect 2466 1331 2500 1365
rect 2541 1331 2575 1365
rect 2615 1331 2649 1365
rect 2689 1331 2723 1365
rect 2763 1331 2797 1365
rect 2837 1331 2871 1365
rect 2911 1331 2945 1365
rect 2985 1331 3019 1365
rect 3059 1331 3093 1365
rect 3133 1331 3167 1365
rect 3207 1331 3241 1365
rect 3281 1331 3315 1365
rect 3355 1331 3389 1365
rect 5005 1404 5039 1419
rect 5005 1385 5039 1404
rect 1919 1315 1953 1316
rect 1919 1243 1953 1276
rect 3539 1331 3573 1365
rect 3614 1331 3648 1365
rect 3689 1331 3723 1365
rect 3764 1331 3798 1365
rect 3839 1331 3873 1365
rect 3914 1331 3948 1365
rect 3989 1331 4023 1365
rect 4064 1331 4098 1365
rect 4139 1331 4173 1365
rect 4214 1331 4248 1365
rect 4289 1331 4323 1365
rect 4364 1331 4398 1365
rect 4439 1331 4473 1365
rect 4514 1331 4548 1365
rect 4589 1331 4623 1365
rect 4663 1331 4697 1365
rect 4737 1331 4771 1365
rect 4811 1331 4845 1365
rect 4885 1331 4919 1365
rect 5005 1336 5039 1344
rect 1919 1242 1953 1243
rect 2095 1239 2129 1273
rect 2170 1239 2204 1273
rect 2245 1239 2279 1273
rect 2319 1239 2353 1273
rect 2393 1239 2427 1273
rect 2467 1239 2501 1273
rect 2541 1239 2575 1273
rect 2615 1239 2649 1273
rect 2689 1239 2723 1273
rect 2763 1239 2797 1273
rect 2837 1239 2871 1273
rect 2911 1239 2945 1273
rect 2985 1239 3019 1273
rect 3059 1239 3093 1273
rect 3133 1239 3167 1273
rect 3207 1239 3241 1273
rect 3281 1239 3315 1273
rect 3355 1239 3389 1273
rect 5005 1310 5039 1336
rect 1919 1170 1953 1202
rect 3625 1239 3659 1273
rect 3699 1239 3733 1273
rect 3773 1239 3807 1273
rect 3847 1239 3881 1273
rect 3921 1239 3955 1273
rect 3994 1239 4028 1273
rect 4067 1239 4101 1273
rect 4140 1239 4174 1273
rect 4213 1239 4247 1273
rect 4286 1239 4320 1273
rect 4359 1239 4393 1273
rect 4432 1239 4466 1273
rect 4505 1239 4539 1273
rect 4578 1239 4612 1273
rect 4651 1239 4685 1273
rect 5005 1268 5039 1270
rect 1919 1168 1953 1170
rect 2241 1147 2275 1181
rect 2316 1147 2350 1181
rect 2391 1147 2425 1181
rect 2466 1147 2500 1181
rect 2541 1147 2575 1181
rect 2615 1147 2649 1181
rect 2689 1147 2723 1181
rect 2763 1147 2797 1181
rect 2837 1147 2871 1181
rect 2911 1147 2945 1181
rect 2985 1147 3019 1181
rect 3059 1147 3093 1181
rect 3133 1147 3167 1181
rect 3207 1147 3241 1181
rect 3281 1147 3315 1181
rect 3355 1147 3389 1181
rect 5005 1236 5039 1268
rect 1919 1097 1953 1128
rect 1919 1094 1953 1097
rect 3539 1147 3573 1181
rect 3614 1147 3648 1181
rect 3689 1147 3723 1181
rect 3764 1147 3798 1181
rect 3839 1147 3873 1181
rect 3914 1147 3948 1181
rect 3989 1147 4023 1181
rect 4064 1147 4098 1181
rect 4139 1147 4173 1181
rect 4214 1147 4248 1181
rect 4289 1147 4323 1181
rect 4364 1147 4398 1181
rect 4439 1147 4473 1181
rect 4514 1147 4548 1181
rect 4589 1147 4623 1181
rect 4663 1147 4697 1181
rect 4737 1147 4771 1181
rect 4811 1147 4845 1181
rect 4885 1147 4919 1181
rect 5005 1166 5039 1196
rect 5005 1162 5039 1166
rect 2095 1055 2129 1089
rect 2170 1055 2204 1089
rect 2245 1055 2279 1089
rect 2319 1055 2353 1089
rect 2393 1055 2427 1089
rect 2467 1055 2501 1089
rect 2541 1055 2575 1089
rect 2615 1055 2649 1089
rect 2689 1055 2723 1089
rect 2763 1055 2797 1089
rect 2837 1055 2871 1089
rect 2911 1055 2945 1089
rect 2985 1055 3019 1089
rect 3059 1055 3093 1089
rect 3133 1055 3167 1089
rect 3207 1055 3241 1089
rect 3281 1055 3315 1089
rect 3355 1055 3389 1089
rect 5005 1098 5039 1122
rect 1919 1024 1953 1054
rect 1919 1020 1953 1024
rect 3625 1055 3659 1089
rect 3699 1055 3733 1089
rect 3773 1055 3807 1089
rect 3847 1055 3881 1089
rect 3921 1055 3955 1089
rect 3994 1055 4028 1089
rect 4067 1055 4101 1089
rect 4140 1055 4174 1089
rect 4213 1055 4247 1089
rect 4286 1055 4320 1089
rect 4359 1055 4393 1089
rect 4432 1055 4466 1089
rect 4505 1055 4539 1089
rect 4578 1055 4612 1089
rect 4651 1055 4685 1089
rect 5005 1088 5039 1098
rect 2241 963 2275 997
rect 2316 963 2350 997
rect 2391 963 2425 997
rect 2466 963 2500 997
rect 2541 963 2575 997
rect 2615 963 2649 997
rect 2689 963 2723 997
rect 2763 963 2797 997
rect 2837 963 2871 997
rect 2911 963 2945 997
rect 2985 963 3019 997
rect 3059 963 3093 997
rect 3133 963 3167 997
rect 3207 963 3241 997
rect 3281 963 3315 997
rect 3355 963 3389 997
rect 3539 963 3573 997
rect 3614 963 3648 997
rect 3689 963 3723 997
rect 3764 963 3798 997
rect 3839 963 3873 997
rect 3914 963 3948 997
rect 3989 963 4023 997
rect 4064 963 4098 997
rect 4139 963 4173 997
rect 4214 963 4248 997
rect 4289 963 4323 997
rect 4364 963 4398 997
rect 4439 963 4473 997
rect 4514 963 4548 997
rect 4589 963 4623 997
rect 4663 963 4697 997
rect 4737 963 4771 997
rect 4811 963 4845 997
rect 4885 963 4919 997
rect 5005 996 5039 998
rect 5005 964 5039 996
rect 2471 864 2489 898
rect 2489 864 2505 898
rect 2543 864 2557 898
rect 2557 864 2577 898
rect 2615 864 2625 898
rect 2625 864 2649 898
rect 2687 864 2693 898
rect 2693 864 2721 898
rect 2759 864 2761 898
rect 2761 864 2793 898
rect 2831 864 2863 898
rect 2863 864 2865 898
rect 2903 864 2931 898
rect 2931 864 2937 898
rect 2975 864 2999 898
rect 2999 864 3009 898
rect 3047 864 3067 898
rect 3067 864 3081 898
rect 3119 864 3135 898
rect 3135 864 3153 898
rect 3191 864 3203 898
rect 3203 864 3225 898
rect 3263 864 3271 898
rect 3271 864 3297 898
rect 3335 864 3339 898
rect 3339 864 3369 898
rect 3407 864 3441 898
rect 3479 864 3509 898
rect 3509 864 3513 898
rect 3551 864 3577 898
rect 3577 864 3585 898
rect 3623 864 3645 898
rect 3645 864 3657 898
rect 3695 864 3713 898
rect 3713 864 3729 898
rect 3767 864 3781 898
rect 3781 864 3801 898
rect 3839 864 3849 898
rect 3849 864 3873 898
rect 3911 864 3917 898
rect 3917 864 3945 898
rect 3984 864 3985 898
rect 3985 864 4018 898
rect 4057 864 4087 898
rect 4087 864 4091 898
rect 4130 864 4155 898
rect 4155 864 4164 898
rect 4203 864 4223 898
rect 4223 864 4237 898
rect 4276 864 4291 898
rect 4291 864 4310 898
rect 4349 864 4359 898
rect 4359 864 4383 898
rect 4422 864 4427 898
rect 4427 864 4456 898
rect 4495 864 4529 898
rect 4568 864 4597 898
rect 4597 864 4602 898
rect 4641 864 4665 898
rect 4665 864 4675 898
rect 4714 864 4733 898
rect 4733 864 4748 898
rect 4787 864 4801 898
rect 4801 864 4821 898
rect 4860 864 4869 898
rect 4869 864 4894 898
rect 4933 864 4937 898
rect 4937 864 4967 898
rect 5414 2013 5448 2047
rect 5486 2013 5520 2047
rect 5558 2013 5592 2047
rect 5630 2013 5664 2047
rect 5702 2013 5736 2047
rect 5774 2013 5808 2047
rect 5846 2013 5880 2047
rect 5918 2013 5952 2047
rect 5990 2013 6024 2047
rect 6062 2013 6096 2047
rect 6134 2013 6168 2047
rect 6206 2013 6240 2047
rect 6278 2013 6312 2047
rect 6350 2013 6384 2047
rect 6595 2013 6629 2047
rect 6667 2013 6701 2047
rect 6739 2013 6773 2047
rect 6811 2013 6845 2047
rect 6883 2013 6917 2047
rect 6955 2013 6989 2047
rect 7027 2013 7061 2047
rect 7099 2013 7133 2047
rect 7171 2013 7205 2047
rect 7243 2013 7277 2047
rect 7315 2013 7349 2047
rect 7387 2013 7421 2047
rect 7459 2013 7493 2047
rect 7531 2013 7565 2047
rect 5414 1939 5448 1973
rect 5486 1947 5520 1973
rect 5486 1939 5518 1947
rect 5518 1939 5520 1947
rect 5558 1939 5592 1973
rect 5630 1947 5664 1973
rect 5630 1939 5656 1947
rect 5656 1939 5664 1947
rect 5702 1939 5736 1973
rect 5774 1947 5808 1973
rect 5774 1939 5794 1947
rect 5794 1939 5808 1947
rect 5846 1939 5880 1973
rect 5918 1947 5952 1973
rect 5918 1939 5932 1947
rect 5932 1939 5952 1947
rect 5990 1939 6024 1973
rect 6062 1947 6096 1973
rect 6062 1939 6070 1947
rect 6070 1939 6096 1947
rect 6134 1939 6168 1973
rect 6206 1947 6240 1973
rect 6206 1939 6208 1947
rect 6208 1939 6240 1947
rect 6278 1939 6312 1973
rect 6350 1939 6384 1973
rect 6595 1947 6629 1973
rect 6595 1939 6622 1947
rect 6622 1939 6629 1947
rect 6667 1939 6701 1973
rect 6739 1947 6773 1973
rect 6739 1939 6760 1947
rect 6760 1939 6773 1947
rect 6811 1939 6845 1973
rect 6883 1947 6917 1973
rect 6883 1939 6898 1947
rect 6898 1939 6917 1947
rect 6955 1939 6989 1973
rect 7027 1947 7061 1973
rect 7027 1939 7036 1947
rect 7036 1939 7061 1947
rect 7099 1939 7133 1973
rect 7171 1947 7205 1973
rect 7171 1939 7174 1947
rect 7174 1939 7205 1947
rect 7243 1939 7277 1973
rect 7315 1939 7349 1973
rect 7387 1947 7421 1973
rect 7387 1939 7416 1947
rect 7416 1939 7421 1947
rect 7459 1939 7493 1973
rect 7531 1947 7565 1973
rect 7531 1939 7554 1947
rect 7554 1939 7565 1947
rect 5414 1865 5448 1899
rect 5486 1865 5520 1899
rect 5558 1865 5592 1899
rect 5630 1865 5664 1899
rect 5702 1865 5736 1899
rect 5774 1865 5808 1899
rect 5846 1865 5880 1899
rect 5918 1865 5952 1899
rect 5990 1865 6024 1899
rect 6062 1865 6096 1899
rect 6134 1865 6168 1899
rect 6206 1865 6240 1899
rect 6278 1865 6312 1899
rect 6350 1865 6384 1899
rect 6595 1865 6629 1899
rect 6667 1865 6701 1899
rect 6739 1865 6773 1899
rect 6811 1865 6845 1899
rect 6883 1865 6917 1899
rect 6955 1865 6989 1899
rect 7027 1865 7061 1899
rect 7099 1865 7133 1899
rect 7171 1865 7205 1899
rect 7243 1865 7277 1899
rect 7315 1865 7349 1899
rect 7387 1865 7421 1899
rect 7459 1865 7493 1899
rect 7531 1865 7565 1899
rect 5414 1791 5448 1825
rect 5486 1809 5520 1825
rect 5486 1791 5518 1809
rect 5518 1791 5520 1809
rect 5558 1791 5592 1825
rect 5630 1809 5664 1825
rect 5630 1791 5656 1809
rect 5656 1791 5664 1809
rect 5702 1791 5736 1825
rect 5774 1809 5808 1825
rect 5774 1791 5794 1809
rect 5794 1791 5808 1809
rect 5846 1791 5880 1825
rect 5918 1809 5952 1825
rect 5918 1791 5932 1809
rect 5932 1791 5952 1809
rect 5990 1791 6024 1825
rect 6062 1809 6096 1825
rect 6062 1791 6070 1809
rect 6070 1791 6096 1809
rect 6134 1791 6168 1825
rect 6206 1809 6240 1825
rect 6206 1791 6208 1809
rect 6208 1791 6240 1809
rect 6278 1791 6312 1825
rect 6350 1791 6384 1825
rect 6595 1809 6629 1825
rect 6595 1791 6622 1809
rect 6622 1791 6629 1809
rect 6667 1791 6701 1825
rect 6739 1809 6773 1825
rect 6739 1791 6760 1809
rect 6760 1791 6773 1809
rect 6811 1791 6845 1825
rect 6883 1809 6917 1825
rect 6883 1791 6898 1809
rect 6898 1791 6917 1809
rect 6955 1791 6989 1825
rect 7027 1809 7061 1825
rect 7027 1791 7036 1809
rect 7036 1791 7061 1809
rect 7099 1791 7133 1825
rect 7171 1809 7205 1825
rect 7171 1791 7174 1809
rect 7174 1791 7205 1809
rect 7243 1791 7277 1825
rect 7315 1791 7349 1825
rect 7387 1809 7421 1825
rect 7387 1791 7416 1809
rect 7416 1791 7421 1809
rect 7459 1791 7493 1825
rect 7531 1809 7565 1825
rect 7531 1791 7554 1809
rect 7554 1791 7565 1809
rect 5414 1717 5448 1751
rect 5486 1717 5520 1751
rect 5558 1717 5592 1751
rect 5630 1717 5664 1751
rect 5702 1717 5736 1751
rect 5774 1717 5808 1751
rect 5846 1717 5880 1751
rect 5918 1717 5952 1751
rect 5990 1717 6024 1751
rect 6062 1717 6096 1751
rect 6134 1717 6168 1751
rect 6206 1717 6240 1751
rect 6278 1717 6312 1751
rect 6350 1717 6384 1751
rect 6595 1717 6629 1751
rect 6667 1717 6701 1751
rect 6739 1717 6773 1751
rect 6811 1717 6845 1751
rect 6883 1717 6917 1751
rect 6955 1717 6989 1751
rect 7027 1717 7061 1751
rect 7099 1717 7133 1751
rect 7171 1717 7205 1751
rect 7243 1717 7277 1751
rect 7315 1717 7349 1751
rect 7387 1717 7421 1751
rect 7459 1717 7493 1751
rect 7531 1717 7565 1751
rect 5414 1642 5448 1676
rect 5486 1671 5520 1676
rect 5486 1642 5518 1671
rect 5518 1642 5520 1671
rect 5558 1642 5592 1676
rect 5630 1671 5664 1676
rect 5630 1642 5656 1671
rect 5656 1642 5664 1671
rect 5702 1642 5736 1676
rect 5774 1671 5808 1676
rect 5774 1642 5794 1671
rect 5794 1642 5808 1671
rect 5846 1642 5880 1676
rect 5918 1671 5952 1676
rect 5918 1642 5932 1671
rect 5932 1642 5952 1671
rect 5990 1642 6024 1676
rect 6062 1671 6096 1676
rect 6062 1642 6070 1671
rect 6070 1642 6096 1671
rect 6134 1642 6168 1676
rect 6206 1671 6240 1676
rect 6206 1642 6208 1671
rect 6208 1642 6240 1671
rect 6278 1642 6312 1676
rect 6350 1642 6384 1676
rect 6595 1671 6629 1676
rect 6595 1642 6622 1671
rect 6622 1642 6629 1671
rect 6667 1642 6701 1676
rect 6739 1671 6773 1676
rect 6739 1642 6760 1671
rect 6760 1642 6773 1671
rect 6811 1642 6845 1676
rect 6883 1671 6917 1676
rect 6883 1642 6898 1671
rect 6898 1642 6917 1671
rect 6955 1642 6989 1676
rect 7027 1671 7061 1676
rect 7027 1642 7036 1671
rect 7036 1642 7061 1671
rect 7099 1642 7133 1676
rect 7171 1671 7205 1676
rect 7171 1642 7174 1671
rect 7174 1642 7205 1671
rect 7243 1642 7277 1676
rect 7315 1642 7349 1676
rect 7387 1671 7421 1676
rect 7387 1642 7416 1671
rect 7416 1642 7421 1671
rect 7459 1642 7493 1676
rect 7531 1671 7565 1676
rect 7531 1642 7554 1671
rect 7554 1642 7565 1671
rect 5414 1567 5448 1601
rect 5486 1567 5520 1601
rect 5558 1567 5592 1601
rect 5630 1567 5664 1601
rect 5702 1567 5736 1601
rect 5774 1567 5808 1601
rect 5846 1567 5880 1601
rect 5918 1567 5952 1601
rect 5990 1567 6024 1601
rect 6062 1567 6096 1601
rect 6134 1567 6168 1601
rect 6206 1567 6240 1601
rect 6278 1567 6312 1601
rect 6350 1567 6384 1601
rect 6595 1567 6629 1601
rect 6667 1567 6701 1601
rect 6739 1567 6773 1601
rect 6811 1567 6845 1601
rect 6883 1567 6917 1601
rect 6955 1567 6989 1601
rect 7027 1567 7061 1601
rect 7099 1567 7133 1601
rect 7171 1567 7205 1601
rect 7243 1567 7277 1601
rect 7315 1567 7349 1601
rect 7387 1567 7421 1601
rect 7459 1567 7493 1601
rect 7531 1567 7565 1601
rect 5414 1492 5448 1526
rect 5486 1498 5518 1526
rect 5518 1498 5520 1526
rect 5486 1492 5520 1498
rect 5558 1492 5592 1526
rect 5630 1498 5656 1526
rect 5656 1498 5664 1526
rect 5630 1492 5664 1498
rect 5702 1492 5736 1526
rect 5774 1498 5794 1526
rect 5794 1498 5808 1526
rect 5774 1492 5808 1498
rect 5846 1492 5880 1526
rect 5918 1498 5932 1526
rect 5932 1498 5952 1526
rect 5918 1492 5952 1498
rect 5990 1492 6024 1526
rect 6062 1498 6070 1526
rect 6070 1498 6096 1526
rect 6062 1492 6096 1498
rect 6134 1492 6168 1526
rect 6206 1498 6208 1526
rect 6208 1498 6240 1526
rect 6206 1492 6240 1498
rect 6278 1492 6312 1526
rect 6350 1492 6384 1526
rect 6595 1498 6622 1526
rect 6622 1498 6629 1526
rect 6595 1492 6629 1498
rect 6667 1492 6701 1526
rect 6739 1498 6760 1526
rect 6760 1498 6773 1526
rect 6739 1492 6773 1498
rect 6811 1492 6845 1526
rect 6883 1498 6898 1526
rect 6898 1498 6917 1526
rect 6883 1492 6917 1498
rect 6955 1492 6989 1526
rect 7027 1498 7036 1526
rect 7036 1498 7061 1526
rect 7027 1492 7061 1498
rect 7099 1492 7133 1526
rect 7171 1498 7174 1526
rect 7174 1498 7205 1526
rect 7171 1492 7205 1498
rect 7243 1492 7277 1526
rect 7315 1492 7349 1526
rect 7387 1498 7416 1526
rect 7416 1498 7421 1526
rect 7387 1492 7421 1498
rect 7459 1492 7493 1526
rect 7531 1498 7554 1526
rect 7554 1498 7565 1526
rect 7531 1492 7565 1498
rect 5414 1417 5448 1451
rect 5486 1417 5520 1451
rect 5558 1417 5592 1451
rect 5630 1417 5664 1451
rect 5702 1417 5736 1451
rect 5774 1417 5808 1451
rect 5846 1417 5880 1451
rect 5918 1417 5952 1451
rect 5990 1417 6024 1451
rect 6062 1417 6096 1451
rect 6134 1417 6168 1451
rect 6206 1417 6240 1451
rect 6278 1417 6312 1451
rect 6350 1417 6384 1451
rect 6595 1417 6629 1451
rect 6667 1417 6701 1451
rect 6739 1417 6773 1451
rect 6811 1417 6845 1451
rect 6883 1417 6917 1451
rect 6955 1417 6989 1451
rect 7027 1417 7061 1451
rect 7099 1417 7133 1451
rect 7171 1417 7205 1451
rect 7243 1417 7277 1451
rect 7315 1417 7349 1451
rect 7387 1417 7421 1451
rect 7459 1417 7493 1451
rect 7531 1417 7565 1451
rect 5414 1342 5448 1376
rect 5486 1359 5518 1376
rect 5518 1359 5520 1376
rect 5486 1342 5520 1359
rect 5558 1342 5592 1376
rect 5630 1359 5656 1376
rect 5656 1359 5664 1376
rect 5630 1342 5664 1359
rect 5702 1342 5736 1376
rect 5774 1359 5794 1376
rect 5794 1359 5808 1376
rect 5774 1342 5808 1359
rect 5846 1342 5880 1376
rect 5918 1359 5932 1376
rect 5932 1359 5952 1376
rect 5918 1342 5952 1359
rect 5990 1342 6024 1376
rect 6062 1359 6070 1376
rect 6070 1359 6096 1376
rect 6062 1342 6096 1359
rect 6134 1342 6168 1376
rect 6206 1359 6208 1376
rect 6208 1359 6240 1376
rect 6206 1342 6240 1359
rect 6278 1342 6312 1376
rect 6350 1342 6384 1376
rect 6595 1359 6622 1376
rect 6622 1359 6629 1376
rect 6595 1342 6629 1359
rect 6667 1342 6701 1376
rect 6739 1359 6760 1376
rect 6760 1359 6773 1376
rect 6739 1342 6773 1359
rect 6811 1342 6845 1376
rect 6883 1359 6898 1376
rect 6898 1359 6917 1376
rect 6883 1342 6917 1359
rect 6955 1342 6989 1376
rect 7027 1359 7036 1376
rect 7036 1359 7061 1376
rect 7027 1342 7061 1359
rect 7099 1342 7133 1376
rect 7171 1359 7174 1376
rect 7174 1359 7205 1376
rect 7171 1342 7205 1359
rect 7243 1342 7277 1376
rect 7315 1342 7349 1376
rect 7387 1359 7416 1376
rect 7416 1359 7421 1376
rect 7387 1342 7421 1359
rect 7459 1342 7493 1376
rect 7531 1359 7554 1376
rect 7554 1359 7565 1376
rect 7531 1342 7565 1359
rect 5414 1267 5448 1301
rect 5486 1267 5520 1301
rect 5558 1267 5592 1301
rect 5630 1267 5664 1301
rect 5702 1267 5736 1301
rect 5774 1267 5808 1301
rect 5846 1267 5880 1301
rect 5918 1267 5952 1301
rect 5990 1267 6024 1301
rect 6062 1267 6096 1301
rect 6134 1267 6168 1301
rect 6206 1267 6240 1301
rect 6278 1267 6312 1301
rect 6350 1267 6384 1301
rect 6595 1267 6629 1301
rect 6667 1267 6701 1301
rect 6739 1267 6773 1301
rect 6811 1267 6845 1301
rect 6883 1267 6917 1301
rect 6955 1267 6989 1301
rect 7027 1267 7061 1301
rect 7099 1267 7133 1301
rect 7171 1267 7205 1301
rect 7243 1267 7277 1301
rect 7315 1267 7349 1301
rect 7387 1267 7421 1301
rect 7459 1267 7493 1301
rect 7531 1267 7565 1301
rect 5414 1192 5448 1226
rect 5486 1220 5518 1226
rect 5518 1220 5520 1226
rect 5486 1192 5520 1220
rect 5558 1192 5592 1226
rect 5630 1220 5656 1226
rect 5656 1220 5664 1226
rect 5630 1192 5664 1220
rect 5702 1192 5736 1226
rect 5774 1220 5794 1226
rect 5794 1220 5808 1226
rect 5774 1192 5808 1220
rect 5846 1192 5880 1226
rect 5918 1220 5932 1226
rect 5932 1220 5952 1226
rect 5918 1192 5952 1220
rect 5990 1192 6024 1226
rect 6062 1220 6070 1226
rect 6070 1220 6096 1226
rect 6062 1192 6096 1220
rect 6134 1192 6168 1226
rect 6206 1220 6208 1226
rect 6208 1220 6240 1226
rect 6206 1192 6240 1220
rect 6278 1192 6312 1226
rect 6350 1192 6384 1226
rect 6595 1220 6622 1226
rect 6622 1220 6629 1226
rect 6595 1192 6629 1220
rect 6667 1192 6701 1226
rect 6739 1220 6760 1226
rect 6760 1220 6773 1226
rect 6739 1192 6773 1220
rect 6811 1192 6845 1226
rect 6883 1220 6898 1226
rect 6898 1220 6917 1226
rect 6883 1192 6917 1220
rect 6955 1192 6989 1226
rect 7027 1220 7036 1226
rect 7036 1220 7061 1226
rect 7027 1192 7061 1220
rect 7099 1192 7133 1226
rect 7171 1220 7174 1226
rect 7174 1220 7205 1226
rect 7171 1192 7205 1220
rect 7243 1192 7277 1226
rect 7315 1192 7349 1226
rect 7387 1220 7416 1226
rect 7416 1220 7421 1226
rect 7387 1192 7421 1220
rect 7459 1192 7493 1226
rect 7531 1220 7554 1226
rect 7554 1220 7565 1226
rect 7531 1192 7565 1220
rect 5414 1117 5448 1151
rect 5486 1117 5520 1151
rect 5558 1117 5592 1151
rect 5630 1117 5664 1151
rect 5702 1117 5736 1151
rect 5774 1117 5808 1151
rect 5846 1117 5880 1151
rect 5918 1117 5952 1151
rect 5990 1117 6024 1151
rect 6062 1117 6096 1151
rect 6134 1117 6168 1151
rect 6206 1117 6240 1151
rect 6278 1117 6312 1151
rect 6350 1117 6384 1151
rect 6595 1117 6629 1151
rect 6667 1117 6701 1151
rect 6739 1117 6773 1151
rect 6811 1117 6845 1151
rect 6883 1117 6917 1151
rect 6955 1117 6989 1151
rect 7027 1117 7061 1151
rect 7099 1117 7133 1151
rect 7171 1117 7205 1151
rect 7243 1117 7277 1151
rect 7315 1117 7349 1151
rect 7387 1117 7421 1151
rect 7459 1117 7493 1151
rect 7531 1117 7565 1151
rect 5414 1042 5448 1076
rect 5486 1042 5520 1076
rect 5558 1042 5592 1076
rect 5630 1042 5664 1076
rect 5702 1042 5736 1076
rect 5774 1042 5808 1076
rect 5846 1042 5880 1076
rect 5918 1042 5952 1076
rect 5990 1042 6024 1076
rect 6062 1042 6096 1076
rect 6134 1042 6168 1076
rect 6206 1042 6240 1076
rect 6278 1042 6312 1076
rect 6350 1042 6384 1076
rect 6595 1042 6629 1076
rect 6667 1042 6701 1076
rect 6739 1042 6773 1076
rect 6811 1042 6845 1076
rect 6883 1042 6917 1076
rect 6955 1042 6989 1076
rect 7027 1042 7061 1076
rect 7099 1042 7133 1076
rect 7171 1042 7205 1076
rect 7243 1042 7277 1076
rect 7315 1042 7349 1076
rect 7387 1042 7421 1076
rect 7459 1042 7493 1076
rect 7531 1042 7565 1076
rect 5414 967 5448 1001
rect 5486 976 5520 1001
rect 5486 967 5518 976
rect 5518 967 5520 976
rect 5558 967 5592 1001
rect 5630 976 5664 1001
rect 5630 967 5656 976
rect 5656 967 5664 976
rect 5702 967 5736 1001
rect 5774 976 5808 1001
rect 5774 967 5794 976
rect 5794 967 5808 976
rect 5846 967 5880 1001
rect 5918 976 5952 1001
rect 5918 967 5932 976
rect 5932 967 5952 976
rect 5990 967 6024 1001
rect 6062 976 6096 1001
rect 6062 967 6070 976
rect 6070 967 6096 976
rect 6134 967 6168 1001
rect 6206 976 6240 1001
rect 6206 967 6208 976
rect 6208 967 6240 976
rect 6278 967 6312 1001
rect 6350 967 6384 1001
rect 6595 976 6629 1001
rect 6595 967 6622 976
rect 6622 967 6629 976
rect 6667 967 6701 1001
rect 6739 976 6773 1001
rect 6739 967 6760 976
rect 6760 967 6773 976
rect 6811 967 6845 1001
rect 6883 976 6917 1001
rect 6883 967 6898 976
rect 6898 967 6917 976
rect 6955 967 6989 1001
rect 7027 976 7061 1001
rect 7027 967 7036 976
rect 7036 967 7061 976
rect 7099 967 7133 1001
rect 7171 976 7205 1001
rect 7171 967 7174 976
rect 7174 967 7205 976
rect 7243 967 7277 1001
rect 7315 967 7349 1001
rect 7387 976 7421 1001
rect 7387 967 7416 976
rect 7416 967 7421 976
rect 7459 967 7493 1001
rect 7531 976 7565 1001
rect 7531 967 7554 976
rect 7554 967 7565 976
rect 5414 892 5448 926
rect 5486 892 5520 926
rect 5558 892 5592 926
rect 5630 892 5664 926
rect 5702 892 5736 926
rect 5774 892 5808 926
rect 5846 892 5880 926
rect 5918 892 5952 926
rect 5990 892 6024 926
rect 6062 892 6096 926
rect 6134 892 6168 926
rect 6206 892 6240 926
rect 6278 892 6312 926
rect 6350 892 6384 926
rect 6595 892 6629 926
rect 6667 892 6701 926
rect 6739 892 6773 926
rect 6811 892 6845 926
rect 6883 892 6917 926
rect 6955 892 6989 926
rect 7027 892 7061 926
rect 7099 892 7133 926
rect 7171 892 7205 926
rect 7243 892 7277 926
rect 7315 892 7349 926
rect 7387 892 7421 926
rect 7459 892 7493 926
rect 7531 892 7565 926
rect 5414 817 5448 851
rect 5486 837 5520 851
rect 5486 817 5518 837
rect 5518 817 5520 837
rect 5558 817 5592 851
rect 5630 837 5664 851
rect 5630 817 5656 837
rect 5656 817 5664 837
rect 5702 817 5736 851
rect 5774 837 5808 851
rect 5774 817 5794 837
rect 5794 817 5808 837
rect 5846 817 5880 851
rect 5918 837 5952 851
rect 5918 817 5932 837
rect 5932 817 5952 837
rect 5990 817 6024 851
rect 6062 837 6096 851
rect 6062 817 6070 837
rect 6070 817 6096 837
rect 6134 817 6168 851
rect 6206 837 6240 851
rect 6206 817 6208 837
rect 6208 817 6240 837
rect 6278 817 6312 851
rect 6350 817 6384 851
rect 6595 837 6629 851
rect 6595 817 6622 837
rect 6622 817 6629 837
rect 6667 817 6701 851
rect 6739 837 6773 851
rect 6739 817 6760 837
rect 6760 817 6773 837
rect 6811 817 6845 851
rect 6883 837 6917 851
rect 6883 817 6898 837
rect 6898 817 6917 837
rect 6955 817 6989 851
rect 7027 837 7061 851
rect 7027 817 7036 837
rect 7036 817 7061 837
rect 7099 817 7133 851
rect 7171 837 7205 851
rect 7171 817 7174 837
rect 7174 817 7205 837
rect 7243 817 7277 851
rect 7315 817 7349 851
rect 7387 837 7421 851
rect 7387 817 7416 837
rect 7416 817 7421 837
rect 7459 817 7493 851
rect 7531 837 7565 851
rect 7531 817 7554 837
rect 7554 817 7565 837
rect 5414 742 5448 776
rect 5486 742 5520 776
rect 5558 742 5592 776
rect 5630 742 5664 776
rect 5702 742 5736 776
rect 5774 742 5808 776
rect 5846 742 5880 776
rect 5918 742 5952 776
rect 5990 742 6024 776
rect 6062 742 6096 776
rect 6134 742 6168 776
rect 6206 742 6240 776
rect 6278 742 6312 776
rect 6350 742 6384 776
rect 6595 742 6629 776
rect 6667 742 6701 776
rect 6739 742 6773 776
rect 6811 742 6845 776
rect 6883 742 6917 776
rect 6955 742 6989 776
rect 7027 742 7061 776
rect 7099 742 7133 776
rect 7171 742 7205 776
rect 7243 742 7277 776
rect 7315 742 7349 776
rect 7387 742 7421 776
rect 7459 742 7493 776
rect 7531 742 7565 776
rect 5414 667 5448 701
rect 5486 698 5520 701
rect 5486 667 5518 698
rect 5518 667 5520 698
rect 5558 667 5592 701
rect 5630 698 5664 701
rect 5630 667 5656 698
rect 5656 667 5664 698
rect 5702 667 5736 701
rect 5774 698 5808 701
rect 5774 667 5794 698
rect 5794 667 5808 698
rect 5846 667 5880 701
rect 5918 698 5952 701
rect 5918 667 5932 698
rect 5932 667 5952 698
rect 5990 667 6024 701
rect 6062 698 6096 701
rect 6062 667 6070 698
rect 6070 667 6096 698
rect 6134 667 6168 701
rect 6206 698 6240 701
rect 6206 667 6208 698
rect 6208 667 6240 698
rect 6278 667 6312 701
rect 6350 667 6384 701
rect 6595 698 6629 701
rect 6595 667 6622 698
rect 6622 667 6629 698
rect 6667 667 6701 701
rect 6739 698 6773 701
rect 6739 667 6760 698
rect 6760 667 6773 698
rect 6811 667 6845 701
rect 6883 698 6917 701
rect 6883 667 6898 698
rect 6898 667 6917 698
rect 6955 667 6989 701
rect 7027 698 7061 701
rect 7027 667 7036 698
rect 7036 667 7061 698
rect 7099 667 7133 701
rect 7171 698 7205 701
rect 7171 667 7174 698
rect 7174 667 7205 698
rect 7243 667 7277 701
rect 7315 667 7349 701
rect 7387 698 7421 701
rect 7387 667 7416 698
rect 7416 667 7421 698
rect 7459 667 7493 701
rect 7531 698 7565 701
rect 7531 667 7554 698
rect 7554 667 7565 698
rect 5414 592 5448 626
rect 5486 592 5520 626
rect 5558 592 5592 626
rect 5630 592 5664 626
rect 5702 592 5736 626
rect 5774 592 5808 626
rect 5846 592 5880 626
rect 5918 592 5952 626
rect 5990 592 6024 626
rect 6062 592 6096 626
rect 6134 592 6168 626
rect 6206 592 6240 626
rect 6278 592 6312 626
rect 6350 592 6384 626
rect 6595 592 6629 626
rect 6667 592 6701 626
rect 6739 592 6773 626
rect 6811 592 6845 626
rect 6883 592 6917 626
rect 6955 592 6989 626
rect 7027 592 7061 626
rect 7099 592 7133 626
rect 7171 592 7205 626
rect 7243 592 7277 626
rect 7315 592 7349 626
rect 7387 592 7421 626
rect 7459 592 7493 626
rect 7531 592 7565 626
rect 5414 517 5448 551
rect 5486 525 5518 551
rect 5518 525 5520 551
rect 5486 517 5520 525
rect 5558 517 5592 551
rect 5630 525 5656 551
rect 5656 525 5664 551
rect 5630 517 5664 525
rect 5702 517 5736 551
rect 5774 525 5794 551
rect 5794 525 5808 551
rect 5774 517 5808 525
rect 5846 517 5880 551
rect 5918 525 5932 551
rect 5932 525 5952 551
rect 5918 517 5952 525
rect 5990 517 6024 551
rect 6062 525 6070 551
rect 6070 525 6096 551
rect 6062 517 6096 525
rect 6134 517 6168 551
rect 6206 525 6208 551
rect 6208 525 6240 551
rect 6206 517 6240 525
rect 6278 517 6312 551
rect 6350 517 6384 551
rect 6595 525 6622 551
rect 6622 525 6629 551
rect 6595 517 6629 525
rect 6667 517 6701 551
rect 6739 525 6760 551
rect 6760 525 6773 551
rect 6739 517 6773 525
rect 6811 517 6845 551
rect 6883 525 6898 551
rect 6898 525 6917 551
rect 6883 517 6917 525
rect 6955 517 6989 551
rect 7027 525 7036 551
rect 7036 525 7061 551
rect 7027 517 7061 525
rect 7099 517 7133 551
rect 7171 525 7174 551
rect 7174 525 7205 551
rect 7171 517 7205 525
rect 7243 517 7277 551
rect 7315 517 7349 551
rect 7387 525 7416 551
rect 7416 525 7421 551
rect 7387 517 7421 525
rect 7459 517 7493 551
rect 7531 525 7554 551
rect 7554 525 7565 551
rect 7531 517 7565 525
rect 5414 442 5448 476
rect 5486 442 5520 476
rect 5558 442 5592 476
rect 5630 442 5664 476
rect 5702 442 5736 476
rect 5774 442 5808 476
rect 5846 442 5880 476
rect 5918 442 5952 476
rect 5990 442 6024 476
rect 6062 442 6096 476
rect 6134 442 6168 476
rect 6206 442 6240 476
rect 6278 442 6312 476
rect 6350 442 6384 476
rect 6595 442 6629 476
rect 6667 442 6701 476
rect 6739 442 6773 476
rect 6811 442 6845 476
rect 6883 442 6917 476
rect 6955 442 6989 476
rect 7027 442 7061 476
rect 7099 442 7133 476
rect 7171 442 7205 476
rect 7243 442 7277 476
rect 7315 442 7349 476
rect 7387 442 7421 476
rect 7459 442 7493 476
rect 7531 442 7565 476
rect 1358 307 1392 341
rect 1451 307 1485 341
rect 1543 307 1577 341
rect 1635 307 1669 341
rect 81 262 115 296
rect 175 262 209 296
rect 81 179 115 213
rect 175 187 204 213
rect 204 187 209 213
rect 175 179 209 187
rect 81 96 115 130
rect 175 119 204 130
rect 204 119 209 130
rect 175 96 209 119
rect 1358 235 1392 269
rect 1451 235 1485 269
rect 1543 235 1577 269
rect 1635 235 1669 269
<< metal1 >>
rect 1938 39476 8573 39482
rect 1938 39470 2163 39476
rect 1938 34108 1944 39470
rect 2050 39370 2163 39470
rect 2989 39442 3028 39476
rect 3062 39442 3101 39476
rect 3135 39442 3174 39476
rect 3208 39442 3247 39476
rect 3281 39442 3320 39476
rect 3354 39442 3393 39476
rect 3427 39442 3466 39476
rect 3500 39442 3539 39476
rect 3573 39442 3612 39476
rect 3646 39442 3685 39476
rect 3719 39442 3758 39476
rect 3792 39442 3831 39476
rect 3865 39442 3904 39476
rect 3938 39442 3977 39476
rect 4011 39442 4050 39476
rect 4084 39442 4123 39476
rect 4157 39442 4196 39476
rect 4230 39442 4269 39476
rect 4303 39442 4342 39476
rect 4376 39442 4415 39476
rect 4449 39442 4488 39476
rect 4522 39442 4561 39476
rect 4595 39442 4634 39476
rect 4668 39442 4707 39476
rect 4741 39442 4780 39476
rect 4814 39442 4853 39476
rect 4887 39442 4926 39476
rect 4960 39442 4999 39476
rect 5033 39442 5072 39476
rect 5106 39442 5145 39476
rect 5179 39442 5218 39476
rect 5252 39442 5291 39476
rect 5325 39442 5364 39476
rect 5398 39442 5437 39476
rect 5471 39442 5510 39476
rect 5544 39442 5583 39476
rect 5617 39442 5656 39476
rect 5690 39442 5729 39476
rect 5763 39442 5802 39476
rect 5836 39442 5875 39476
rect 5909 39442 5948 39476
rect 5982 39442 6021 39476
rect 6055 39442 6094 39476
rect 6128 39442 6167 39476
rect 6201 39442 6240 39476
rect 6274 39442 6313 39476
rect 6347 39442 6386 39476
rect 6420 39442 6459 39476
rect 6493 39442 6532 39476
rect 6566 39442 6605 39476
rect 6639 39442 6678 39476
rect 6712 39442 6751 39476
rect 6785 39442 6824 39476
rect 6858 39442 6897 39476
rect 6931 39442 6970 39476
rect 7004 39442 7043 39476
rect 7077 39442 7116 39476
rect 7150 39442 7189 39476
rect 7223 39442 7262 39476
rect 7296 39442 7335 39476
rect 7369 39442 7408 39476
rect 7442 39442 7481 39476
rect 7515 39442 7554 39476
rect 7588 39442 7627 39476
rect 7661 39442 7786 39476
rect 7820 39442 7866 39476
rect 7900 39442 7946 39476
rect 7980 39442 8026 39476
rect 8060 39442 8106 39476
rect 8140 39442 8186 39476
rect 8220 39442 8267 39476
rect 8301 39442 8348 39476
rect 8382 39442 8429 39476
rect 8463 39442 8573 39476
rect 2989 39404 8573 39442
rect 2989 39370 3028 39404
rect 3062 39370 3101 39404
rect 3135 39370 3174 39404
rect 3208 39370 3247 39404
rect 3281 39370 3320 39404
rect 3354 39370 3393 39404
rect 3427 39370 3466 39404
rect 3500 39370 3539 39404
rect 3573 39370 3612 39404
rect 3646 39370 3685 39404
rect 3719 39370 3758 39404
rect 3792 39370 3831 39404
rect 3865 39370 3904 39404
rect 3938 39370 3977 39404
rect 4011 39370 4050 39404
rect 4084 39370 4123 39404
rect 4157 39370 4196 39404
rect 4230 39370 4269 39404
rect 4303 39370 4342 39404
rect 4376 39370 4415 39404
rect 4449 39370 4488 39404
rect 4522 39370 4561 39404
rect 4595 39370 4634 39404
rect 4668 39370 4707 39404
rect 4741 39370 4780 39404
rect 4814 39370 4853 39404
rect 4887 39370 4926 39404
rect 4960 39370 4999 39404
rect 5033 39370 5072 39404
rect 5106 39370 5145 39404
rect 5179 39370 5218 39404
rect 5252 39370 5291 39404
rect 5325 39370 5364 39404
rect 5398 39370 5437 39404
rect 5471 39370 5510 39404
rect 5544 39370 5583 39404
rect 5617 39370 5656 39404
rect 5690 39370 5729 39404
rect 5763 39370 5802 39404
rect 5836 39370 5875 39404
rect 5909 39370 5948 39404
rect 5982 39370 6021 39404
rect 6055 39370 6094 39404
rect 6128 39370 6167 39404
rect 6201 39370 6240 39404
rect 6274 39370 6313 39404
rect 6347 39370 6386 39404
rect 6420 39370 6459 39404
rect 6493 39370 6532 39404
rect 6566 39370 6605 39404
rect 6639 39370 6678 39404
rect 6712 39370 6751 39404
rect 6785 39370 6824 39404
rect 6858 39370 6897 39404
rect 6931 39370 6970 39404
rect 7004 39370 7043 39404
rect 7077 39370 7116 39404
rect 7150 39370 7189 39404
rect 7223 39370 7262 39404
rect 7296 39370 7335 39404
rect 7369 39370 7408 39404
rect 7442 39370 7481 39404
rect 7515 39370 7554 39404
rect 7588 39370 7627 39404
rect 7661 39370 7786 39404
rect 7820 39370 7866 39404
rect 7900 39370 7946 39404
rect 7980 39370 8026 39404
rect 8060 39370 8106 39404
rect 8140 39370 8186 39404
rect 8220 39370 8267 39404
rect 8301 39370 8348 39404
rect 8382 39370 8429 39404
rect 2050 39364 8429 39370
rect 2050 34108 2056 39364
tri 2056 39330 2090 39364 nw
tri 8375 39330 8409 39364 ne
rect 8409 39330 8429 39364
tri 8409 39316 8423 39330 ne
rect 1938 34069 2056 34108
rect 1938 34035 1944 34069
rect 1978 34035 2016 34069
rect 2050 34035 2056 34069
rect 1938 33996 2056 34035
rect 1938 33962 1944 33996
rect 1978 33962 2016 33996
rect 2050 33962 2056 33996
rect 1938 33923 2056 33962
rect 1938 33889 1944 33923
rect 1978 33889 2016 33923
rect 2050 33889 2056 33923
rect 1938 33850 2056 33889
rect 1938 33816 1944 33850
rect 1978 33816 2016 33850
rect 2050 33816 2056 33850
rect 1938 33777 2056 33816
rect 1938 33743 1944 33777
rect 1978 33743 2016 33777
rect 2050 33743 2056 33777
rect 1938 33704 2056 33743
rect 1938 33670 1944 33704
rect 1978 33670 2016 33704
rect 2050 33670 2056 33704
rect 1938 33607 2056 33670
rect 1938 27020 1944 33607
rect 2050 27020 2056 33607
rect 1938 26956 1944 26968
rect 2050 26956 2056 26968
rect 1938 11037 1944 26904
rect 2050 11037 2056 26904
rect 1938 10998 2056 11037
rect 1938 10964 1944 10998
rect 1978 10964 2016 10998
rect 2050 10964 2056 10998
rect 1938 10925 2056 10964
rect 1938 10891 1944 10925
rect 1978 10891 2016 10925
rect 2050 10891 2056 10925
rect 1938 10847 2056 10891
rect 1938 10813 1944 10847
rect 1978 10813 2016 10847
rect 2050 10813 2056 10847
rect 1938 10774 2056 10813
rect 1938 10740 1944 10774
rect 1978 10740 2016 10774
rect 2050 10740 2056 10774
rect 1938 10701 2056 10740
rect 1938 10667 1944 10701
rect 1978 10667 2016 10701
rect 2050 10667 2056 10701
rect 1938 10628 2056 10667
rect 1938 8938 1944 10628
rect 2050 9785 2056 10628
rect 2270 39141 8224 39147
rect 2270 39107 2348 39141
rect 2382 39107 2420 39141
rect 2454 39107 2492 39141
rect 2526 39107 2564 39141
rect 2598 39107 2636 39141
rect 2670 39107 2708 39141
rect 2742 39107 2780 39141
rect 2814 39107 2852 39141
rect 2886 39107 2924 39141
rect 2958 39107 2996 39141
rect 3030 39107 3068 39141
rect 3102 39107 3140 39141
rect 3174 39107 3212 39141
rect 3246 39107 3284 39141
rect 3318 39107 3356 39141
rect 3390 39107 3428 39141
rect 3462 39107 3500 39141
rect 3534 39107 3572 39141
rect 3606 39107 3644 39141
rect 3678 39107 3716 39141
rect 3750 39107 3788 39141
rect 3822 39107 3860 39141
rect 3894 39107 3932 39141
rect 3966 39107 4004 39141
rect 4038 39107 4076 39141
rect 4110 39107 4148 39141
rect 4182 39107 4220 39141
rect 4254 39107 4292 39141
rect 4326 39107 4364 39141
rect 4398 39107 4436 39141
rect 4470 39107 4508 39141
rect 4542 39107 4580 39141
rect 4614 39107 4652 39141
rect 4686 39107 4724 39141
rect 4758 39107 4796 39141
rect 4830 39107 4868 39141
rect 4902 39107 4940 39141
rect 4974 39107 5012 39141
rect 5046 39107 5084 39141
rect 5118 39107 5156 39141
rect 5190 39107 5228 39141
rect 5262 39107 5300 39141
rect 5334 39107 5372 39141
rect 5406 39107 5444 39141
rect 5478 39107 5516 39141
rect 5550 39107 5588 39141
rect 5622 39107 5660 39141
rect 5694 39107 5732 39141
rect 5766 39107 5804 39141
rect 5838 39107 5877 39141
rect 5911 39107 5950 39141
rect 5984 39107 6023 39141
rect 6057 39107 6096 39141
rect 6130 39107 6169 39141
rect 6203 39107 6242 39141
rect 6276 39107 6315 39141
rect 6349 39107 6388 39141
rect 6422 39107 6461 39141
rect 6495 39107 6534 39141
rect 6568 39107 6607 39141
rect 6641 39107 6680 39141
rect 6714 39107 6753 39141
rect 6787 39107 6826 39141
rect 6860 39107 6963 39141
rect 6997 39107 7039 39141
rect 7073 39107 7115 39141
rect 7149 39107 7191 39141
rect 7225 39107 7267 39141
rect 7301 39107 7343 39141
rect 7377 39107 7419 39141
rect 7453 39107 7496 39141
rect 7530 39107 7573 39141
rect 7607 39107 7650 39141
rect 7684 39107 7727 39141
rect 7761 39107 7804 39141
rect 7838 39107 7881 39141
rect 7915 39107 7958 39141
rect 7992 39107 8035 39141
rect 8069 39107 8112 39141
rect 8146 39107 8224 39141
rect 2270 39069 8224 39107
rect 2270 39035 2276 39069
rect 2310 39035 8184 39069
rect 8218 39035 8224 39069
rect 2270 39007 8224 39035
rect 2270 38996 2410 39007
rect 2270 38962 2276 38996
rect 2310 38973 2410 38996
rect 2444 38973 2482 39007
rect 2516 38973 2554 39007
rect 2588 38973 2626 39007
rect 2660 38973 2698 39007
rect 2732 38973 2770 39007
rect 2804 38973 2842 39007
rect 2876 38973 2914 39007
rect 2948 38973 2986 39007
rect 3020 38973 3058 39007
rect 3092 38973 3130 39007
rect 3164 38973 3202 39007
rect 3236 38973 3274 39007
rect 3308 38973 3346 39007
rect 3380 38973 3418 39007
rect 3452 38973 3490 39007
rect 3524 38973 3562 39007
rect 3596 38973 3634 39007
rect 3668 38973 3706 39007
rect 3740 38973 3778 39007
rect 3812 38973 3850 39007
rect 3884 38973 3922 39007
rect 3956 38973 3994 39007
rect 4028 38973 4066 39007
rect 4100 38973 4138 39007
rect 4172 38973 4210 39007
rect 4244 38973 4282 39007
rect 4316 38973 4354 39007
rect 4388 38973 4426 39007
rect 4460 38973 4498 39007
rect 4532 38973 4570 39007
rect 4604 38973 4642 39007
rect 4676 38973 4714 39007
rect 4748 38973 4786 39007
rect 4820 38973 4858 39007
rect 4892 38973 4930 39007
rect 4964 38973 5002 39007
rect 5036 38973 5074 39007
rect 5108 38973 5147 39007
rect 5181 38973 5220 39007
rect 5254 38973 5293 39007
rect 5327 38973 5366 39007
rect 5400 38973 5439 39007
rect 5473 38973 5512 39007
rect 5546 38973 5585 39007
rect 5619 38973 5658 39007
rect 5692 38973 5731 39007
rect 5765 38973 5804 39007
rect 5838 38973 5877 39007
rect 5911 38973 5950 39007
rect 5984 38973 6023 39007
rect 6057 38973 6096 39007
rect 6130 38973 6169 39007
rect 6203 38973 6242 39007
rect 6276 38973 6315 39007
rect 6349 38973 6388 39007
rect 6422 38973 6461 39007
rect 6495 38973 6534 39007
rect 6568 38973 6607 39007
rect 6641 38973 6680 39007
rect 6714 38973 6753 39007
rect 6787 38973 6826 39007
rect 6860 38973 6963 39007
rect 6997 38973 7035 39007
rect 7069 38973 7107 39007
rect 7141 38973 7179 39007
rect 7213 38973 7251 39007
rect 7285 38973 7323 39007
rect 7357 38973 7395 39007
rect 7429 38973 7467 39007
rect 7501 38973 7539 39007
rect 7573 38973 7612 39007
rect 7646 38973 7685 39007
rect 7719 38973 7758 39007
rect 7792 38973 7831 39007
rect 7865 38973 7904 39007
rect 7938 38973 7977 39007
rect 8011 38973 8050 39007
rect 8084 38997 8224 39007
rect 8084 38973 8184 38997
rect 2310 38967 8184 38973
rect 2310 38963 2480 38967
tri 2480 38963 2484 38967 nw
tri 8018 38963 8022 38967 ne
rect 8022 38963 8184 38967
rect 8218 38963 8224 38997
rect 2310 38962 2452 38963
rect 2270 38935 2452 38962
tri 2452 38935 2480 38963 nw
tri 8022 38941 8044 38963 ne
rect 8044 38935 8224 38963
rect 2270 38934 2450 38935
rect 2270 38923 2410 38934
rect 2270 38889 2276 38923
rect 2310 38900 2410 38923
rect 2444 38900 2450 38934
tri 2450 38933 2452 38935 nw
rect 2310 38889 2450 38900
rect 2270 38861 2450 38889
rect 8044 38901 8050 38935
rect 8084 38925 8224 38935
rect 8084 38901 8184 38925
rect 8044 38891 8184 38901
rect 8218 38891 8224 38925
rect 2270 38850 2410 38861
rect 2270 38816 2276 38850
rect 2310 38827 2410 38850
rect 2444 38827 2450 38861
rect 2310 38816 2450 38827
rect 2270 38788 2450 38816
rect 2270 38777 2410 38788
rect 2270 38743 2276 38777
rect 2310 38754 2410 38777
rect 2444 38754 2450 38788
rect 2310 38743 2450 38754
rect 2270 38724 2450 38743
rect 2322 38672 2392 38724
rect 2444 38672 2450 38724
rect 2270 38670 2276 38672
rect 2310 38670 2450 38672
rect 2270 38655 2450 38670
rect 2322 38603 2392 38655
rect 2444 38603 2450 38655
rect 2270 38597 2276 38603
rect 2310 38597 2450 38603
rect 2270 38586 2450 38597
rect 2322 38534 2392 38586
rect 2444 38534 2450 38586
rect 2270 38524 2276 38534
rect 2310 38524 2450 38534
rect 2270 38517 2450 38524
rect 2322 38465 2392 38517
rect 2270 38451 2276 38465
rect 2310 38462 2410 38465
rect 2444 38462 2450 38517
rect 2310 38451 2450 38462
rect 2270 38448 2450 38451
rect 2322 38396 2392 38448
rect 2270 38378 2276 38396
rect 2310 38389 2410 38396
rect 2444 38389 2450 38448
rect 2310 38378 2450 38389
rect 2322 38326 2392 38378
rect 2270 38308 2276 38326
rect 2310 38316 2410 38326
rect 2444 38316 2450 38378
rect 2310 38308 2450 38316
rect 2322 38256 2392 38308
rect 2270 38238 2276 38256
rect 2310 38243 2410 38256
rect 2444 38243 2450 38308
rect 2310 38238 2450 38243
rect 2322 38186 2392 38238
rect 2270 38168 2276 38186
rect 2310 38170 2410 38186
rect 2444 38170 2450 38238
rect 2310 38168 2450 38170
rect 2322 38116 2392 38168
rect 2270 38086 2276 38116
rect 2310 38097 2410 38116
rect 2444 38097 2450 38168
rect 2310 38086 2450 38097
rect 2270 38058 2450 38086
rect 2270 38047 2410 38058
rect 2270 38013 2276 38047
rect 2310 38024 2410 38047
rect 2444 38024 2450 38058
rect 2310 38013 2450 38024
rect 2270 37985 2450 38013
rect 2270 37974 2410 37985
rect 2270 37940 2276 37974
rect 2310 37951 2410 37974
rect 2444 37951 2450 37985
rect 2310 37940 2450 37951
rect 2270 37912 2450 37940
rect 2270 37901 2410 37912
rect 2270 37867 2276 37901
rect 2310 37878 2410 37901
rect 2444 37878 2450 37912
rect 2310 37867 2450 37878
rect 2270 37839 2450 37867
rect 2270 37828 2410 37839
rect 2270 37794 2276 37828
rect 2310 37805 2410 37828
rect 2444 37805 2450 37839
rect 2310 37794 2450 37805
rect 2270 37766 2450 37794
rect 2270 37755 2410 37766
rect 2270 37721 2276 37755
rect 2310 37732 2410 37755
rect 2444 37732 2450 37766
rect 2310 37721 2450 37732
rect 2270 37693 2450 37721
rect 2270 37682 2410 37693
rect 2270 37648 2276 37682
rect 2310 37659 2410 37682
rect 2444 37659 2450 37693
rect 2310 37648 2450 37659
rect 2270 37620 2450 37648
rect 2270 37609 2410 37620
rect 2270 37575 2276 37609
rect 2310 37586 2410 37609
rect 2444 37586 2450 37620
rect 2310 37575 2450 37586
rect 2270 37547 2450 37575
rect 2270 37536 2410 37547
rect 2270 37502 2276 37536
rect 2310 37513 2410 37536
rect 2444 37513 2450 37547
rect 2310 37502 2450 37513
rect 2270 37474 2450 37502
rect 2270 37463 2410 37474
rect 2270 37429 2276 37463
rect 2310 37440 2410 37463
rect 2444 37440 2450 37474
rect 2310 37429 2450 37440
rect 2270 37401 2450 37429
rect 2270 37390 2410 37401
rect 2270 37356 2276 37390
rect 2310 37367 2410 37390
rect 2444 37367 2450 37401
rect 2310 37356 2450 37367
rect 2270 37328 2450 37356
rect 2270 37317 2410 37328
rect 2270 37283 2276 37317
rect 2310 37294 2410 37317
rect 2444 37294 2450 37328
rect 2310 37283 2450 37294
rect 2270 37255 2450 37283
rect 2270 37244 2410 37255
rect 2270 37210 2276 37244
rect 2310 37221 2410 37244
rect 2444 37221 2450 37255
rect 2310 37210 2450 37221
rect 2270 37182 2450 37210
rect 2270 37171 2410 37182
rect 2270 37137 2276 37171
rect 2310 37148 2410 37171
rect 2444 37148 2450 37182
rect 2310 37137 2450 37148
rect 2270 37109 2450 37137
rect 2270 37098 2410 37109
rect 2270 37064 2276 37098
rect 2310 37075 2410 37098
rect 2444 37075 2450 37109
rect 2310 37064 2450 37075
rect 2270 37036 2450 37064
rect 2270 37025 2410 37036
rect 2270 36991 2276 37025
rect 2310 37002 2410 37025
rect 2444 37002 2450 37036
rect 2310 36991 2450 37002
rect 2270 36963 2450 36991
rect 2270 36952 2410 36963
rect 2270 36918 2276 36952
rect 2310 36929 2410 36952
rect 2444 36929 2450 36963
rect 2310 36918 2450 36929
rect 2270 36890 2450 36918
rect 2270 36879 2410 36890
rect 2270 36845 2276 36879
rect 2310 36856 2410 36879
rect 2444 36856 2450 36890
rect 2310 36845 2450 36856
rect 2270 36817 2450 36845
rect 2270 36806 2410 36817
rect 2270 36772 2276 36806
rect 2310 36783 2410 36806
rect 2444 36783 2450 36817
rect 2310 36772 2450 36783
rect 2270 36744 2450 36772
rect 2270 36733 2410 36744
rect 2270 36724 2276 36733
rect 2310 36724 2410 36733
rect 2322 36672 2392 36724
rect 2444 36672 2450 36744
rect 2270 36671 2450 36672
rect 2270 36660 2410 36671
rect 2270 36655 2276 36660
rect 2310 36655 2410 36660
rect 2322 36603 2392 36655
rect 2444 36603 2450 36671
rect 2270 36598 2450 36603
rect 2270 36588 2410 36598
rect 2270 36586 2276 36588
rect 2310 36586 2410 36588
rect 2322 36534 2392 36586
rect 2444 36534 2450 36598
rect 2270 36525 2450 36534
rect 2270 36517 2410 36525
rect 2322 36465 2392 36517
rect 2444 36465 2450 36525
rect 2270 36452 2450 36465
rect 2270 36448 2410 36452
rect 2322 36396 2392 36448
rect 2444 36396 2450 36452
rect 2270 36379 2450 36396
rect 2270 36378 2410 36379
rect 2322 36326 2392 36378
rect 2444 36326 2450 36379
rect 2270 36308 2450 36326
rect 2322 36256 2392 36308
rect 2444 36256 2450 36308
rect 2270 36238 2450 36256
rect 2322 36186 2392 36238
rect 2444 36186 2450 36238
rect 2270 36168 2450 36186
rect 2322 36116 2392 36168
rect 2444 36116 2450 36168
rect 2270 36087 2450 36116
rect 2270 36084 2410 36087
rect 2270 36050 2276 36084
rect 2310 36053 2410 36084
rect 2444 36053 2450 36087
rect 2310 36050 2450 36053
rect 2270 36014 2450 36050
rect 2270 36012 2410 36014
rect 2270 35978 2276 36012
rect 2310 35980 2410 36012
rect 2444 35980 2450 36014
rect 2310 35978 2450 35980
rect 2270 35941 2450 35978
rect 2270 35940 2410 35941
rect 2270 35906 2276 35940
rect 2310 35907 2410 35940
rect 2444 35907 2450 35941
rect 2310 35906 2450 35907
rect 2270 35868 2450 35906
rect 2270 35834 2276 35868
rect 2310 35834 2410 35868
rect 2444 35834 2450 35868
rect 2270 35796 2450 35834
rect 2270 35762 2276 35796
rect 2310 35762 2410 35796
rect 2444 35762 2450 35796
rect 2270 35724 2450 35762
rect 2270 35690 2276 35724
rect 2310 35690 2410 35724
rect 2444 35690 2450 35724
rect 2270 35652 2450 35690
rect 2270 35618 2276 35652
rect 2310 35618 2410 35652
rect 2444 35618 2450 35652
rect 2270 35580 2450 35618
rect 2270 35546 2276 35580
rect 2310 35546 2410 35580
rect 2444 35546 2450 35580
rect 2270 35508 2450 35546
rect 2270 35474 2276 35508
rect 2310 35474 2410 35508
rect 2444 35474 2450 35508
rect 2270 35436 2450 35474
rect 2270 35402 2276 35436
rect 2310 35402 2410 35436
rect 2444 35402 2450 35436
rect 2270 35364 2450 35402
rect 2270 35330 2276 35364
rect 2310 35330 2410 35364
rect 2444 35330 2450 35364
rect 2270 35292 2450 35330
rect 2270 35258 2276 35292
rect 2310 35258 2410 35292
rect 2444 35258 2450 35292
rect 2270 35220 2450 35258
rect 2270 35186 2276 35220
rect 2310 35186 2410 35220
rect 2444 35186 2450 35220
rect 2270 35148 2450 35186
rect 2270 35114 2276 35148
rect 2310 35114 2410 35148
rect 2444 35114 2450 35148
rect 2270 35076 2450 35114
rect 2270 35042 2276 35076
rect 2310 35042 2410 35076
rect 2444 35042 2450 35076
rect 2270 35004 2450 35042
rect 2270 34970 2276 35004
rect 2310 34970 2410 35004
rect 2444 34970 2450 35004
rect 2270 34932 2450 34970
rect 2270 34898 2276 34932
rect 2310 34898 2410 34932
rect 2444 34898 2450 34932
rect 2270 34860 2450 34898
rect 2270 34826 2276 34860
rect 2310 34826 2410 34860
rect 2444 34826 2450 34860
rect 2270 34788 2450 34826
rect 2270 34754 2276 34788
rect 2310 34754 2410 34788
rect 2444 34754 2450 34788
rect 2270 34724 2450 34754
rect 2322 34672 2392 34724
rect 2444 34672 2450 34724
rect 2270 34655 2450 34672
rect 2322 34603 2392 34655
rect 2444 34603 2450 34655
rect 2270 34586 2450 34603
rect 2322 34534 2392 34586
rect 2444 34534 2450 34586
rect 2270 34517 2450 34534
rect 2322 34465 2392 34517
rect 2444 34465 2450 34517
rect 2270 34448 2450 34465
rect 2322 34396 2392 34448
rect 2270 34394 2276 34396
rect 2310 34394 2410 34396
rect 2444 34394 2450 34448
rect 2270 34378 2450 34394
rect 2322 34326 2392 34378
rect 2270 34322 2276 34326
rect 2310 34322 2410 34326
rect 2444 34322 2450 34378
rect 2270 34308 2450 34322
rect 2322 34256 2392 34308
rect 2270 34250 2276 34256
rect 2310 34250 2410 34256
rect 2444 34250 2450 34308
rect 2270 34238 2450 34250
rect 2322 34186 2392 34238
rect 2270 34178 2276 34186
rect 2310 34178 2410 34186
rect 2444 34178 2450 34238
rect 2270 34168 2450 34178
rect 2322 34116 2392 34168
rect 2270 34106 2276 34116
rect 2310 34106 2410 34116
rect 2444 34106 2450 34168
rect 2270 34068 2450 34106
rect 2270 34034 2276 34068
rect 2310 34034 2410 34068
rect 2444 34034 2450 34068
rect 2270 33996 2450 34034
rect 2270 33962 2276 33996
rect 2310 33962 2410 33996
rect 2444 33962 2450 33996
rect 2270 33924 2450 33962
rect 2270 33890 2276 33924
rect 2310 33890 2410 33924
rect 2444 33890 2450 33924
rect 2270 33852 2450 33890
rect 2270 33818 2276 33852
rect 2310 33818 2410 33852
rect 2444 33818 2450 33852
rect 2270 33780 2450 33818
rect 2270 33746 2276 33780
rect 2310 33746 2410 33780
rect 2444 33746 2450 33780
rect 2270 33708 2450 33746
rect 2270 33674 2276 33708
rect 2310 33674 2410 33708
rect 2444 33674 2450 33708
rect 2270 33636 2450 33674
rect 2270 33602 2276 33636
rect 2310 33602 2410 33636
rect 2444 33602 2450 33636
rect 2270 33564 2450 33602
rect 2270 33530 2276 33564
rect 2310 33530 2410 33564
rect 2444 33530 2450 33564
rect 2270 33492 2450 33530
rect 2270 33458 2276 33492
rect 2310 33458 2410 33492
rect 2444 33458 2450 33492
rect 2270 33420 2450 33458
rect 2270 33386 2276 33420
rect 2310 33386 2410 33420
rect 2444 33386 2450 33420
rect 2270 33348 2450 33386
rect 2270 33314 2276 33348
rect 2310 33314 2410 33348
rect 2444 33314 2450 33348
rect 2270 33276 2450 33314
rect 2270 33242 2276 33276
rect 2310 33242 2410 33276
rect 2444 33242 2450 33276
rect 2270 33204 2450 33242
rect 2270 33170 2276 33204
rect 2310 33170 2410 33204
rect 2444 33170 2450 33204
rect 2270 33132 2450 33170
rect 2270 33098 2276 33132
rect 2310 33098 2410 33132
rect 2444 33098 2450 33132
rect 2270 33060 2450 33098
rect 2270 33026 2276 33060
rect 2310 33026 2410 33060
rect 2444 33026 2450 33060
rect 2270 32988 2450 33026
rect 2270 32954 2276 32988
rect 2310 32954 2410 32988
rect 2444 32954 2450 32988
rect 2270 32916 2450 32954
rect 2270 32882 2276 32916
rect 2310 32882 2410 32916
rect 2444 32882 2450 32916
rect 2270 32844 2450 32882
rect 2270 32810 2276 32844
rect 2310 32810 2410 32844
rect 2444 32810 2450 32844
rect 2270 32772 2450 32810
rect 2270 32738 2276 32772
rect 2310 32738 2410 32772
rect 2444 32738 2450 32772
rect 2270 32724 2450 32738
rect 2322 32672 2392 32724
rect 2270 32666 2276 32672
rect 2310 32666 2410 32672
rect 2444 32666 2450 32724
rect 2270 32655 2450 32666
rect 2322 32603 2392 32655
rect 2270 32594 2276 32603
rect 2310 32594 2410 32603
rect 2444 32594 2450 32655
rect 2270 32586 2450 32594
rect 2322 32534 2392 32586
rect 2270 32522 2276 32534
rect 2310 32522 2410 32534
rect 2444 32522 2450 32586
rect 2270 32517 2450 32522
rect 2322 32465 2392 32517
rect 2270 32450 2276 32465
rect 2310 32450 2410 32465
rect 2444 32450 2450 32517
rect 2270 32448 2450 32450
rect 2322 32396 2392 32448
rect 2270 32378 2276 32396
rect 2310 32378 2410 32396
rect 2322 32326 2392 32378
rect 2270 32308 2276 32326
rect 2310 32308 2410 32326
rect 2322 32256 2392 32308
rect 2270 32238 2276 32256
rect 2310 32238 2410 32256
rect 2322 32186 2392 32238
rect 2270 32168 2276 32186
rect 2310 32168 2410 32186
rect 2322 32116 2392 32168
rect 2270 32090 2276 32116
rect 2310 32090 2410 32116
rect 2444 32090 2450 32448
rect 2270 32052 2450 32090
rect 2270 32018 2276 32052
rect 2310 32018 2410 32052
rect 2444 32018 2450 32052
rect 2270 31980 2450 32018
rect 2270 31946 2276 31980
rect 2310 31946 2410 31980
rect 2444 31946 2450 31980
rect 2270 31908 2450 31946
rect 2270 31874 2276 31908
rect 2310 31874 2410 31908
rect 2444 31874 2450 31908
rect 2270 31836 2450 31874
rect 2270 31802 2276 31836
rect 2310 31802 2410 31836
rect 2444 31802 2450 31836
rect 2270 31764 2450 31802
rect 2270 31730 2276 31764
rect 2310 31730 2410 31764
rect 2444 31730 2450 31764
rect 2270 31692 2450 31730
rect 2270 31658 2276 31692
rect 2310 31658 2410 31692
rect 2444 31658 2450 31692
rect 2270 31620 2450 31658
rect 2270 31586 2276 31620
rect 2310 31586 2410 31620
rect 2444 31586 2450 31620
rect 2270 31548 2450 31586
rect 2270 31514 2276 31548
rect 2310 31514 2410 31548
rect 2444 31514 2450 31548
rect 2270 31476 2450 31514
rect 2270 31442 2276 31476
rect 2310 31442 2410 31476
rect 2444 31442 2450 31476
rect 2270 31404 2450 31442
rect 2270 31370 2276 31404
rect 2310 31370 2410 31404
rect 2444 31370 2450 31404
rect 2270 31332 2450 31370
rect 2270 31298 2276 31332
rect 2310 31298 2410 31332
rect 2444 31298 2450 31332
rect 2270 31260 2450 31298
rect 2270 31226 2276 31260
rect 2310 31226 2410 31260
rect 2444 31226 2450 31260
rect 2270 31188 2450 31226
rect 2270 31154 2276 31188
rect 2310 31154 2410 31188
rect 2444 31154 2450 31188
rect 2270 31116 2450 31154
rect 2270 31082 2276 31116
rect 2310 31082 2410 31116
rect 2444 31082 2450 31116
rect 2270 31044 2450 31082
rect 2270 31010 2276 31044
rect 2310 31010 2410 31044
rect 2444 31010 2450 31044
rect 2270 30972 2450 31010
rect 2270 30938 2276 30972
rect 2310 30938 2410 30972
rect 2444 30938 2450 30972
rect 2270 30900 2450 30938
rect 2270 30866 2276 30900
rect 2310 30866 2410 30900
rect 2444 30866 2450 30900
rect 2270 30828 2450 30866
rect 2270 30794 2276 30828
rect 2310 30794 2410 30828
rect 2444 30794 2450 30828
rect 2270 30756 2450 30794
rect 2270 30724 2276 30756
rect 2310 30724 2410 30756
rect 2322 30672 2392 30724
rect 2270 30655 2276 30672
rect 2310 30655 2410 30672
rect 2322 30603 2392 30655
rect 2270 30586 2276 30603
rect 2310 30586 2410 30603
rect 2322 30534 2392 30586
rect 2270 30517 2276 30534
rect 2310 30517 2410 30534
rect 2322 30465 2392 30517
rect 2270 30448 2276 30465
rect 2310 30448 2410 30465
rect 2322 30396 2392 30448
rect 2270 30378 2276 30396
rect 2310 30378 2410 30396
rect 2322 30326 2392 30378
rect 2444 30326 2450 30756
rect 2270 30324 2450 30326
rect 2270 30308 2276 30324
rect 2310 30308 2410 30324
rect 2322 30256 2392 30308
rect 2444 30256 2450 30324
rect 2270 30252 2450 30256
rect 2270 30238 2276 30252
rect 2310 30238 2410 30252
rect 2322 30186 2392 30238
rect 2444 30186 2450 30252
rect 2270 30180 2450 30186
rect 2270 30168 2276 30180
rect 2310 30168 2410 30180
rect 2322 30116 2392 30168
rect 2444 30116 2450 30180
rect 2270 30108 2450 30116
rect 2270 30074 2276 30108
rect 2310 30074 2410 30108
rect 2444 30074 2450 30108
rect 2270 30036 2450 30074
rect 2270 30002 2276 30036
rect 2310 30002 2410 30036
rect 2444 30002 2450 30036
rect 2270 29964 2450 30002
rect 2270 29930 2276 29964
rect 2310 29930 2410 29964
rect 2444 29930 2450 29964
rect 2270 29892 2450 29930
rect 2270 29858 2276 29892
rect 2310 29858 2410 29892
rect 2444 29858 2450 29892
rect 2270 29820 2450 29858
rect 2270 29786 2276 29820
rect 2310 29786 2410 29820
rect 2444 29786 2450 29820
rect 2270 29748 2450 29786
rect 2270 29714 2276 29748
rect 2310 29714 2410 29748
rect 2444 29714 2450 29748
rect 2270 29676 2450 29714
rect 2270 29642 2276 29676
rect 2310 29642 2410 29676
rect 2444 29642 2450 29676
rect 2270 29604 2450 29642
rect 2270 29570 2276 29604
rect 2310 29570 2410 29604
rect 2444 29570 2450 29604
rect 2270 29532 2450 29570
rect 2270 29498 2276 29532
rect 2310 29498 2410 29532
rect 2444 29498 2450 29532
rect 2270 29460 2450 29498
rect 2270 29426 2276 29460
rect 2310 29426 2410 29460
rect 2444 29426 2450 29460
rect 2270 29388 2450 29426
rect 2270 29354 2276 29388
rect 2310 29354 2410 29388
rect 2444 29354 2450 29388
rect 2270 29316 2450 29354
rect 2270 29282 2276 29316
rect 2310 29282 2410 29316
rect 2444 29282 2450 29316
rect 2270 29244 2450 29282
rect 2270 29210 2276 29244
rect 2310 29210 2410 29244
rect 2444 29210 2450 29244
rect 2270 29172 2450 29210
rect 2270 29138 2276 29172
rect 2310 29138 2410 29172
rect 2444 29138 2450 29172
rect 2270 29100 2450 29138
rect 2543 38854 7729 38886
rect 2543 38820 3035 38854
rect 3069 38820 3108 38854
rect 3142 38820 3181 38854
rect 3215 38820 3254 38854
rect 3288 38820 3327 38854
rect 3361 38820 3400 38854
rect 3434 38820 3473 38854
rect 3507 38820 3546 38854
rect 3580 38820 3619 38854
rect 3653 38820 3692 38854
rect 3726 38820 3765 38854
rect 3799 38820 3838 38854
rect 3872 38820 3911 38854
rect 3945 38820 3984 38854
rect 4018 38820 4057 38854
rect 4091 38820 4130 38854
rect 4164 38820 4203 38854
rect 4237 38820 4276 38854
rect 4310 38820 4349 38854
rect 4383 38820 4422 38854
rect 4456 38820 4495 38854
rect 4529 38820 4568 38854
rect 4602 38820 4641 38854
rect 4675 38820 4714 38854
rect 4748 38820 4787 38854
rect 4821 38820 4860 38854
rect 4894 38820 4933 38854
rect 4967 38820 5006 38854
rect 5040 38820 5079 38854
rect 5113 38820 5152 38854
rect 5186 38820 5225 38854
rect 5259 38820 5298 38854
rect 5332 38820 5371 38854
rect 5405 38820 5444 38854
rect 5478 38820 5517 38854
rect 5551 38820 5590 38854
rect 5624 38820 5663 38854
rect 5697 38820 5736 38854
rect 5770 38820 5809 38854
rect 5843 38820 5882 38854
rect 5916 38820 5955 38854
rect 5989 38820 6027 38854
rect 6061 38820 6099 38854
rect 6133 38820 6171 38854
rect 6205 38820 6243 38854
rect 6277 38820 6315 38854
rect 6349 38820 6387 38854
rect 6421 38820 6459 38854
rect 6493 38820 6531 38854
rect 6565 38820 6603 38854
rect 6637 38820 6675 38854
rect 6709 38820 6747 38854
rect 6781 38820 6819 38854
rect 6853 38820 6891 38854
rect 6925 38820 6963 38854
rect 6997 38820 7035 38854
rect 7069 38820 7107 38854
rect 7141 38820 7179 38854
rect 7213 38820 7251 38854
rect 7285 38820 7323 38854
rect 7357 38820 7395 38854
rect 7429 38820 7467 38854
rect 7501 38820 7539 38854
rect 7573 38820 7611 38854
rect 7645 38820 7683 38854
rect 7717 38820 7729 38854
rect 2543 38814 7729 38820
rect 8044 38863 8224 38891
rect 8044 38829 8050 38863
rect 8084 38853 8224 38863
rect 8084 38829 8184 38853
rect 8044 38819 8184 38829
rect 8218 38819 8224 38853
rect 2543 38791 2767 38814
tri 2767 38791 2790 38814 nw
rect 8044 38791 8224 38819
rect 2543 38757 2733 38791
tri 2733 38757 2767 38791 nw
rect 8044 38757 8050 38791
rect 8084 38781 8224 38791
rect 8084 38757 8184 38781
rect 2543 38747 2723 38757
tri 2723 38747 2733 38757 nw
rect 8044 38747 8184 38757
rect 8218 38747 8224 38781
rect 2543 37207 2712 38747
tri 2712 38736 2723 38747 nw
rect 2824 38720 2942 38726
rect 2876 38668 2890 38720
rect 2824 38651 2942 38668
rect 2876 38599 2890 38651
rect 2824 38582 2942 38599
rect 2876 38530 2890 38582
rect 2824 38513 2942 38530
rect 2876 38461 2890 38513
rect 2824 38444 2942 38461
rect 2876 38422 2890 38444
rect 2824 38375 2830 38392
rect 2936 38375 2942 38392
rect 2824 38306 2830 38323
rect 2936 38306 2942 38323
rect 2824 38236 2830 38254
rect 2936 38236 2942 38254
rect 2824 38166 2830 38184
rect 2936 38166 2942 38184
rect 2824 37380 2830 38114
rect 2936 37380 2942 38114
rect 2824 37368 2942 37380
rect 3101 38714 3219 38726
rect 3101 38680 3107 38714
rect 3141 38680 3179 38714
rect 3213 38680 3219 38714
rect 3101 38641 3219 38680
rect 3101 38607 3107 38641
rect 3141 38607 3179 38641
rect 3213 38607 3219 38641
rect 3101 38568 3219 38607
rect 3101 38534 3107 38568
rect 3141 38534 3179 38568
rect 3213 38534 3219 38568
rect 3101 38495 3219 38534
rect 3101 38461 3107 38495
rect 3141 38461 3179 38495
rect 3213 38461 3219 38495
rect 3101 38422 3219 38461
rect 3101 37982 3107 38422
rect 3213 37982 3219 38422
rect 3101 37913 3107 37930
rect 3213 37913 3219 37930
rect 3101 37844 3107 37861
rect 3213 37844 3219 37861
rect 3101 37775 3107 37792
rect 3213 37775 3219 37792
rect 3101 37706 3107 37723
rect 3213 37706 3219 37723
rect 3101 37636 3107 37654
rect 3213 37636 3219 37654
rect 3101 37566 3107 37584
rect 3213 37566 3219 37584
rect 3101 37496 3107 37514
rect 3213 37496 3219 37514
rect 3101 37426 3107 37444
rect 3213 37426 3219 37444
rect 3153 37374 3167 37380
rect 3101 37368 3219 37374
rect 3378 38720 3496 38726
rect 3430 38668 3444 38720
rect 3378 38651 3496 38668
rect 3430 38599 3444 38651
rect 3378 38582 3496 38599
rect 3430 38530 3444 38582
rect 3378 38513 3496 38530
rect 3430 38461 3444 38513
rect 3378 38444 3496 38461
rect 3430 38422 3444 38444
rect 3378 38375 3384 38392
rect 3490 38375 3496 38392
rect 3378 38306 3384 38323
rect 3490 38306 3496 38323
rect 3378 38236 3384 38254
rect 3490 38236 3496 38254
rect 3378 38166 3384 38184
rect 3490 38166 3496 38184
rect 3378 37380 3384 38114
rect 3490 37380 3496 38114
rect 3378 37368 3496 37380
rect 3655 38714 3773 38726
rect 3655 38680 3661 38714
rect 3695 38680 3733 38714
rect 3767 38680 3773 38714
rect 3655 38641 3773 38680
rect 3655 38607 3661 38641
rect 3695 38607 3733 38641
rect 3767 38607 3773 38641
rect 3655 38568 3773 38607
rect 3655 38534 3661 38568
rect 3695 38534 3733 38568
rect 3767 38534 3773 38568
rect 3655 38495 3773 38534
rect 3655 38461 3661 38495
rect 3695 38461 3733 38495
rect 3767 38461 3773 38495
rect 3655 38422 3773 38461
rect 3655 37982 3661 38422
rect 3767 37982 3773 38422
rect 3655 37913 3661 37930
rect 3767 37913 3773 37930
rect 3655 37844 3661 37861
rect 3767 37844 3773 37861
rect 3655 37775 3661 37792
rect 3767 37775 3773 37792
rect 3655 37706 3661 37723
rect 3767 37706 3773 37723
rect 3655 37636 3661 37654
rect 3767 37636 3773 37654
rect 3655 37566 3661 37584
rect 3767 37566 3773 37584
rect 3655 37496 3661 37514
rect 3767 37496 3773 37514
rect 3655 37426 3661 37444
rect 3767 37426 3773 37444
rect 3707 37374 3721 37380
rect 3655 37368 3773 37374
rect 3932 38720 4050 38726
rect 3984 38668 3998 38720
rect 3932 38651 4050 38668
rect 3984 38599 3998 38651
rect 3932 38582 4050 38599
rect 3984 38530 3998 38582
rect 3932 38513 4050 38530
rect 3984 38461 3998 38513
rect 3932 38444 4050 38461
rect 3984 38422 3998 38444
rect 3932 38375 3938 38392
rect 4044 38375 4050 38392
rect 3932 38306 3938 38323
rect 4044 38306 4050 38323
rect 3932 38236 3938 38254
rect 4044 38236 4050 38254
rect 3932 38166 3938 38184
rect 4044 38166 4050 38184
rect 3932 37380 3938 38114
rect 4044 37380 4050 38114
rect 3932 37368 4050 37380
rect 4209 38714 4327 38726
rect 4209 38680 4215 38714
rect 4249 38680 4287 38714
rect 4321 38680 4327 38714
rect 4209 38641 4327 38680
rect 4209 38607 4215 38641
rect 4249 38607 4287 38641
rect 4321 38607 4327 38641
rect 4209 38568 4327 38607
rect 4209 38534 4215 38568
rect 4249 38534 4287 38568
rect 4321 38534 4327 38568
rect 4209 38495 4327 38534
rect 4209 38461 4215 38495
rect 4249 38461 4287 38495
rect 4321 38461 4327 38495
rect 4209 38422 4327 38461
rect 4209 37982 4215 38422
rect 4321 37982 4327 38422
rect 4209 37913 4215 37930
rect 4321 37913 4327 37930
rect 4209 37844 4215 37861
rect 4321 37844 4327 37861
rect 4209 37775 4215 37792
rect 4321 37775 4327 37792
rect 4209 37706 4215 37723
rect 4321 37706 4327 37723
rect 4209 37636 4215 37654
rect 4321 37636 4327 37654
rect 4209 37566 4215 37584
rect 4321 37566 4327 37584
rect 4209 37496 4215 37514
rect 4321 37496 4327 37514
rect 4209 37426 4215 37444
rect 4321 37426 4327 37444
rect 4261 37374 4275 37380
rect 4209 37368 4327 37374
rect 4486 38720 4604 38726
rect 4538 38668 4552 38720
rect 4486 38651 4604 38668
rect 4538 38599 4552 38651
rect 4486 38582 4604 38599
rect 4538 38530 4552 38582
rect 4486 38513 4604 38530
rect 4538 38461 4552 38513
rect 4486 38444 4604 38461
rect 4538 38422 4552 38444
rect 4486 38375 4492 38392
rect 4598 38375 4604 38392
rect 4486 38306 4492 38323
rect 4598 38306 4604 38323
rect 4486 38236 4492 38254
rect 4598 38236 4604 38254
rect 4486 38166 4492 38184
rect 4598 38166 4604 38184
rect 4486 37380 4492 38114
rect 4598 37380 4604 38114
rect 4486 37368 4604 37380
rect 4763 38714 4881 38726
rect 4763 38680 4769 38714
rect 4803 38680 4841 38714
rect 4875 38680 4881 38714
rect 4763 38641 4881 38680
rect 4763 38607 4769 38641
rect 4803 38607 4841 38641
rect 4875 38607 4881 38641
rect 4763 38568 4881 38607
rect 4763 38534 4769 38568
rect 4803 38534 4841 38568
rect 4875 38534 4881 38568
rect 4763 38495 4881 38534
rect 4763 38461 4769 38495
rect 4803 38461 4841 38495
rect 4875 38461 4881 38495
rect 4763 38422 4881 38461
rect 4763 37982 4769 38422
rect 4875 37982 4881 38422
rect 4763 37913 4769 37930
rect 4875 37913 4881 37930
rect 4763 37844 4769 37861
rect 4875 37844 4881 37861
rect 4763 37775 4769 37792
rect 4875 37775 4881 37792
rect 4763 37706 4769 37723
rect 4875 37706 4881 37723
rect 4763 37636 4769 37654
rect 4875 37636 4881 37654
rect 4763 37566 4769 37584
rect 4875 37566 4881 37584
rect 4763 37496 4769 37514
rect 4875 37496 4881 37514
rect 4763 37426 4769 37444
rect 4875 37426 4881 37444
rect 4815 37374 4829 37380
rect 4763 37368 4881 37374
rect 5040 38720 5158 38726
rect 5092 38668 5106 38720
rect 5040 38651 5158 38668
rect 5092 38599 5106 38651
rect 5040 38582 5158 38599
rect 5092 38530 5106 38582
rect 5040 38513 5158 38530
rect 5092 38461 5106 38513
rect 5040 38444 5158 38461
rect 5092 38422 5106 38444
rect 5040 38375 5046 38392
rect 5152 38375 5158 38392
rect 5040 38306 5046 38323
rect 5152 38306 5158 38323
rect 5040 38236 5046 38254
rect 5152 38236 5158 38254
rect 5040 38166 5046 38184
rect 5152 38166 5158 38184
rect 5040 37380 5046 38114
rect 5152 37380 5158 38114
rect 5040 37368 5158 37380
rect 5317 38714 5435 38726
rect 5317 38680 5323 38714
rect 5357 38680 5395 38714
rect 5429 38680 5435 38714
rect 5317 38641 5435 38680
rect 5317 38607 5323 38641
rect 5357 38607 5395 38641
rect 5429 38607 5435 38641
rect 5317 38568 5435 38607
rect 5317 38534 5323 38568
rect 5357 38534 5395 38568
rect 5429 38534 5435 38568
rect 5317 38495 5435 38534
rect 5317 38461 5323 38495
rect 5357 38461 5395 38495
rect 5429 38461 5435 38495
rect 5317 38422 5435 38461
rect 5317 37982 5323 38422
rect 5429 37982 5435 38422
rect 5317 37913 5323 37930
rect 5429 37913 5435 37930
rect 5317 37844 5323 37861
rect 5429 37844 5435 37861
rect 5317 37775 5323 37792
rect 5429 37775 5435 37792
rect 5317 37706 5323 37723
rect 5429 37706 5435 37723
rect 5317 37636 5323 37654
rect 5429 37636 5435 37654
rect 5317 37566 5323 37584
rect 5429 37566 5435 37584
rect 5317 37496 5323 37514
rect 5429 37496 5435 37514
rect 5317 37426 5323 37444
rect 5429 37426 5435 37444
rect 5369 37374 5383 37380
rect 5317 37368 5435 37374
rect 5594 38720 5712 38726
rect 5646 38668 5660 38720
rect 5594 38651 5712 38668
rect 5646 38599 5660 38651
rect 5594 38582 5712 38599
rect 5646 38530 5660 38582
rect 5594 38513 5712 38530
rect 5646 38461 5660 38513
rect 5594 38444 5712 38461
rect 5646 38422 5660 38444
rect 5594 38375 5600 38392
rect 5706 38375 5712 38392
rect 5594 38306 5600 38323
rect 5706 38306 5712 38323
rect 5594 38236 5600 38254
rect 5706 38236 5712 38254
rect 5594 38166 5600 38184
rect 5706 38166 5712 38184
rect 5594 37380 5600 38114
rect 5706 37380 5712 38114
rect 5594 37368 5712 37380
rect 5871 38714 5989 38726
rect 5871 38680 5877 38714
rect 5911 38680 5949 38714
rect 5983 38680 5989 38714
rect 5871 38641 5989 38680
rect 5871 38607 5877 38641
rect 5911 38607 5949 38641
rect 5983 38607 5989 38641
rect 5871 38568 5989 38607
rect 5871 38534 5877 38568
rect 5911 38534 5949 38568
rect 5983 38534 5989 38568
rect 5871 38495 5989 38534
rect 5871 38461 5877 38495
rect 5911 38461 5949 38495
rect 5983 38461 5989 38495
rect 5871 38422 5989 38461
rect 5871 37982 5877 38422
rect 5983 37982 5989 38422
rect 5871 37913 5877 37930
rect 5983 37913 5989 37930
rect 5871 37844 5877 37861
rect 5983 37844 5989 37861
rect 5871 37775 5877 37792
rect 5983 37775 5989 37792
rect 5871 37706 5877 37723
rect 5983 37706 5989 37723
rect 5871 37636 5877 37654
rect 5983 37636 5989 37654
rect 5871 37566 5877 37584
rect 5983 37566 5989 37584
rect 5871 37496 5877 37514
rect 5983 37496 5989 37514
rect 5871 37426 5877 37444
rect 5983 37426 5989 37444
rect 5923 37374 5937 37380
rect 5871 37368 5989 37374
rect 6148 38720 6266 38726
rect 6200 38668 6214 38720
rect 6148 38651 6266 38668
rect 6200 38599 6214 38651
rect 6148 38582 6266 38599
rect 6200 38530 6214 38582
rect 6148 38513 6266 38530
rect 6200 38461 6214 38513
rect 6148 38444 6266 38461
rect 6200 38422 6214 38444
rect 6148 38375 6154 38392
rect 6260 38375 6266 38392
rect 6148 38306 6154 38323
rect 6260 38306 6266 38323
rect 6148 38236 6154 38254
rect 6260 38236 6266 38254
rect 6148 38166 6154 38184
rect 6260 38166 6266 38184
rect 6148 37380 6154 38114
rect 6260 37380 6266 38114
rect 6148 37368 6266 37380
rect 6425 38714 6543 38726
rect 6425 38680 6431 38714
rect 6465 38680 6503 38714
rect 6537 38680 6543 38714
rect 6425 38641 6543 38680
rect 6425 38607 6431 38641
rect 6465 38607 6503 38641
rect 6537 38607 6543 38641
rect 6425 38568 6543 38607
rect 6425 38534 6431 38568
rect 6465 38534 6503 38568
rect 6537 38534 6543 38568
rect 6425 38495 6543 38534
rect 6425 38461 6431 38495
rect 6465 38461 6503 38495
rect 6537 38461 6543 38495
rect 6425 38422 6543 38461
rect 6425 37982 6431 38422
rect 6537 37982 6543 38422
rect 6425 37913 6431 37930
rect 6537 37913 6543 37930
rect 6425 37844 6431 37861
rect 6537 37844 6543 37861
rect 6425 37775 6431 37792
rect 6537 37775 6543 37792
rect 6425 37706 6431 37723
rect 6537 37706 6543 37723
rect 6425 37636 6431 37654
rect 6537 37636 6543 37654
rect 6425 37566 6431 37584
rect 6537 37566 6543 37584
rect 6425 37496 6431 37514
rect 6537 37496 6543 37514
rect 6425 37426 6431 37444
rect 6537 37426 6543 37444
rect 6477 37374 6491 37380
rect 6425 37368 6543 37374
rect 6702 38720 6820 38726
rect 6754 38668 6768 38720
rect 6702 38651 6820 38668
rect 6754 38599 6768 38651
rect 6702 38582 6820 38599
rect 6754 38530 6768 38582
rect 6702 38513 6820 38530
rect 6754 38461 6768 38513
rect 6702 38444 6820 38461
rect 6754 38422 6768 38444
rect 6702 38375 6708 38392
rect 6814 38375 6820 38392
rect 6702 38306 6708 38323
rect 6814 38306 6820 38323
rect 6702 38236 6708 38254
rect 6814 38236 6820 38254
rect 6702 38166 6708 38184
rect 6814 38166 6820 38184
rect 6702 37380 6708 38114
rect 6814 37380 6820 38114
rect 6702 37368 6820 37380
rect 6979 38714 7097 38726
rect 6979 38680 6985 38714
rect 7019 38680 7057 38714
rect 7091 38680 7097 38714
rect 6979 38641 7097 38680
rect 6979 38607 6985 38641
rect 7019 38607 7057 38641
rect 7091 38607 7097 38641
rect 6979 38568 7097 38607
rect 6979 38534 6985 38568
rect 7019 38534 7057 38568
rect 7091 38534 7097 38568
rect 6979 38495 7097 38534
rect 6979 38461 6985 38495
rect 7019 38461 7057 38495
rect 7091 38461 7097 38495
rect 6979 38422 7097 38461
rect 6979 37982 6985 38422
rect 7091 37982 7097 38422
rect 6979 37913 6985 37930
rect 7091 37913 7097 37930
rect 6979 37844 6985 37861
rect 7091 37844 7097 37861
rect 6979 37775 6985 37792
rect 7091 37775 7097 37792
rect 6979 37706 6985 37723
rect 7091 37706 7097 37723
rect 6979 37636 6985 37654
rect 7091 37636 7097 37654
rect 6979 37566 6985 37584
rect 7091 37566 7097 37584
rect 6979 37496 6985 37514
rect 7091 37496 7097 37514
rect 6979 37426 6985 37444
rect 7091 37426 7097 37444
rect 7031 37374 7045 37380
rect 6979 37368 7097 37374
rect 7256 38720 7374 38726
rect 7308 38668 7322 38720
rect 7256 38651 7374 38668
rect 7308 38599 7322 38651
rect 7256 38582 7374 38599
rect 7308 38530 7322 38582
rect 7256 38513 7374 38530
rect 7308 38461 7322 38513
rect 7256 38444 7374 38461
rect 7308 38422 7322 38444
rect 7256 38375 7262 38392
rect 7368 38375 7374 38392
rect 7256 38306 7262 38323
rect 7368 38306 7374 38323
rect 7256 38236 7262 38254
rect 7368 38236 7374 38254
rect 7256 38166 7262 38184
rect 7368 38166 7374 38184
rect 7256 37380 7262 38114
rect 7368 37380 7374 38114
rect 7256 37368 7374 37380
rect 7533 38714 7651 38726
rect 7533 38680 7539 38714
rect 7573 38680 7611 38714
rect 7645 38680 7651 38714
rect 7533 38641 7651 38680
rect 7533 38607 7539 38641
rect 7573 38607 7611 38641
rect 7645 38607 7651 38641
rect 7533 38568 7651 38607
rect 7533 38534 7539 38568
rect 7573 38534 7611 38568
rect 7645 38534 7651 38568
rect 7533 38495 7651 38534
rect 7533 38461 7539 38495
rect 7573 38461 7611 38495
rect 7645 38461 7651 38495
rect 7533 38422 7651 38461
rect 7533 37982 7539 38422
rect 7645 37982 7651 38422
rect 7533 37913 7539 37930
rect 7645 37913 7651 37930
rect 7533 37844 7539 37861
rect 7645 37844 7651 37861
rect 7533 37775 7539 37792
rect 7645 37775 7651 37792
rect 7533 37706 7539 37723
rect 7645 37706 7651 37723
rect 7533 37636 7539 37654
rect 7645 37636 7651 37654
rect 7533 37566 7539 37584
rect 7645 37566 7651 37584
rect 7533 37496 7539 37514
rect 7645 37496 7651 37514
rect 7533 37426 7539 37444
rect 7645 37426 7651 37444
rect 7585 37374 7599 37380
rect 7533 37368 7651 37374
rect 7810 38720 7928 38726
rect 7862 38668 7876 38720
rect 7810 38651 7928 38668
rect 7862 38599 7876 38651
rect 7810 38582 7928 38599
rect 7862 38530 7876 38582
rect 7810 38513 7928 38530
rect 7862 38461 7876 38513
rect 7810 38444 7928 38461
rect 7862 38422 7876 38444
rect 7810 38375 7816 38392
rect 7922 38375 7928 38392
rect 7810 38306 7816 38323
rect 7922 38306 7928 38323
rect 7810 38236 7816 38254
rect 7922 38236 7928 38254
rect 7810 38166 7816 38184
rect 7922 38166 7928 38184
rect 7810 37380 7816 38114
rect 7922 37380 7928 38114
rect 7810 37368 7928 37380
rect 8044 38724 8224 38747
rect 8044 38672 8047 38724
rect 8099 38672 8169 38724
rect 8221 38672 8224 38724
rect 8044 38655 8224 38672
rect 8044 38603 8047 38655
rect 8099 38603 8169 38655
rect 8221 38603 8224 38655
rect 8044 38586 8224 38603
rect 8044 38534 8047 38586
rect 8099 38534 8169 38586
rect 8221 38534 8224 38586
rect 8044 38531 8184 38534
rect 8218 38531 8224 38534
rect 8044 38517 8224 38531
rect 8044 38465 8047 38517
rect 8099 38465 8169 38517
rect 8221 38465 8224 38517
rect 8044 38459 8184 38465
rect 8218 38459 8224 38465
rect 8044 38448 8224 38459
rect 8044 38396 8047 38448
rect 8099 38396 8169 38448
rect 8221 38396 8224 38448
rect 8044 38387 8184 38396
rect 8218 38387 8224 38396
rect 8044 38378 8224 38387
rect 8044 38326 8047 38378
rect 8099 38326 8169 38378
rect 8221 38326 8224 38378
rect 8044 38325 8050 38326
rect 8084 38325 8184 38326
rect 8044 38315 8184 38325
rect 8218 38315 8224 38326
rect 8044 38308 8224 38315
rect 8044 38256 8047 38308
rect 8099 38256 8169 38308
rect 8221 38256 8224 38308
rect 8044 38253 8050 38256
rect 8084 38253 8184 38256
rect 8044 38243 8184 38253
rect 8218 38243 8224 38256
rect 8044 38238 8224 38243
rect 8044 38186 8047 38238
rect 8099 38186 8169 38238
rect 8221 38186 8224 38238
rect 8044 38181 8050 38186
rect 8084 38181 8184 38186
rect 8044 38171 8184 38181
rect 8218 38171 8224 38186
rect 8044 38168 8224 38171
rect 8044 38116 8047 38168
rect 8099 38116 8169 38168
rect 8221 38116 8224 38168
rect 8044 38109 8050 38116
rect 8084 38109 8184 38116
rect 8044 38099 8184 38109
rect 8218 38099 8224 38116
rect 8044 38071 8224 38099
rect 8044 38037 8050 38071
rect 8084 38061 8224 38071
rect 8084 38037 8184 38061
rect 8044 38027 8184 38037
rect 8218 38027 8224 38061
rect 8044 37999 8224 38027
rect 8044 37965 8050 37999
rect 8084 37989 8224 37999
rect 8084 37965 8184 37989
rect 8044 37955 8184 37965
rect 8218 37955 8224 37989
rect 8044 37927 8224 37955
rect 8044 37893 8050 37927
rect 8084 37917 8224 37927
rect 8084 37893 8184 37917
rect 8044 37883 8184 37893
rect 8218 37883 8224 37917
rect 8044 37855 8224 37883
rect 8044 37821 8050 37855
rect 8084 37845 8224 37855
rect 8084 37821 8184 37845
rect 8044 37811 8184 37821
rect 8218 37811 8224 37845
rect 8044 37783 8224 37811
rect 8044 37749 8050 37783
rect 8084 37773 8224 37783
rect 8084 37749 8184 37773
rect 8044 37739 8184 37749
rect 8218 37739 8224 37773
rect 8044 37711 8224 37739
rect 8044 37677 8050 37711
rect 8084 37701 8224 37711
rect 8084 37677 8184 37701
rect 8044 37667 8184 37677
rect 8218 37667 8224 37701
rect 8044 37639 8224 37667
rect 8044 37605 8050 37639
rect 8084 37629 8224 37639
rect 8084 37605 8184 37629
rect 8044 37595 8184 37605
rect 8218 37595 8224 37629
rect 8044 37567 8224 37595
rect 8044 37533 8050 37567
rect 8084 37557 8224 37567
rect 8084 37533 8184 37557
rect 8044 37523 8184 37533
rect 8218 37523 8224 37557
rect 8044 37495 8224 37523
rect 8044 37461 8050 37495
rect 8084 37485 8224 37495
rect 8084 37461 8184 37485
rect 8044 37451 8184 37461
rect 8218 37451 8224 37485
rect 8044 37423 8224 37451
rect 8044 37389 8050 37423
rect 8084 37413 8224 37423
rect 8084 37389 8184 37413
rect 8044 37379 8184 37389
rect 8218 37379 8224 37413
rect 8044 37351 8224 37379
rect 8044 37317 8050 37351
rect 8084 37341 8224 37351
rect 8084 37317 8184 37341
rect 8044 37307 8184 37317
rect 8218 37307 8224 37341
rect 8044 37279 8224 37307
rect 8044 37245 8050 37279
rect 8084 37269 8224 37279
rect 8084 37245 8184 37269
rect 8044 37235 8184 37245
rect 8218 37235 8224 37269
tri 2712 37207 2723 37218 sw
rect 8044 37207 8224 37235
rect 2543 37173 2723 37207
tri 2723 37173 2757 37207 sw
rect 8044 37173 8050 37207
rect 8084 37197 8224 37207
rect 8084 37173 8184 37197
rect 2543 37163 2757 37173
tri 2757 37163 2767 37173 sw
rect 8044 37163 8184 37173
rect 8218 37163 8224 37197
rect 2543 37135 2767 37163
tri 2767 37135 2795 37163 sw
rect 8044 37135 8224 37163
rect 2543 37129 2795 37135
tri 2795 37129 2801 37135 sw
rect 2543 37065 7750 37129
rect 2543 37031 3035 37065
rect 3069 37031 3108 37065
rect 3142 37031 3181 37065
rect 3215 37031 3254 37065
rect 3288 37031 3327 37065
rect 3361 37031 3400 37065
rect 3434 37031 3473 37065
rect 3507 37031 3546 37065
rect 3580 37031 3619 37065
rect 3653 37031 3692 37065
rect 3726 37031 3765 37065
rect 3799 37031 3838 37065
rect 3872 37031 3911 37065
rect 3945 37031 3984 37065
rect 4018 37031 4057 37065
rect 4091 37031 4130 37065
rect 4164 37031 4203 37065
rect 4237 37031 4276 37065
rect 4310 37031 4349 37065
rect 4383 37031 4422 37065
rect 4456 37031 4495 37065
rect 4529 37031 4568 37065
rect 4602 37031 4641 37065
rect 4675 37031 4714 37065
rect 4748 37031 4787 37065
rect 4821 37031 4860 37065
rect 4894 37031 4933 37065
rect 4967 37031 5006 37065
rect 5040 37031 5079 37065
rect 5113 37031 5152 37065
rect 5186 37031 5225 37065
rect 5259 37031 5298 37065
rect 5332 37031 5371 37065
rect 5405 37031 5444 37065
rect 5478 37031 5517 37065
rect 5551 37031 5590 37065
rect 5624 37031 5663 37065
rect 5697 37031 5736 37065
rect 5770 37031 5809 37065
rect 5843 37031 5882 37065
rect 5916 37031 5955 37065
rect 5989 37031 6027 37065
rect 6061 37031 6099 37065
rect 6133 37031 6171 37065
rect 6205 37031 6243 37065
rect 6277 37031 6315 37065
rect 6349 37031 6387 37065
rect 6421 37031 6459 37065
rect 6493 37031 6531 37065
rect 6565 37031 6603 37065
rect 6637 37031 6675 37065
rect 6709 37031 6747 37065
rect 6781 37031 6819 37065
rect 6853 37031 6891 37065
rect 6925 37031 6963 37065
rect 6997 37031 7035 37065
rect 7069 37031 7107 37065
rect 7141 37031 7179 37065
rect 7213 37031 7251 37065
rect 7285 37031 7323 37065
rect 7357 37031 7395 37065
rect 7429 37031 7467 37065
rect 7501 37031 7539 37065
rect 7573 37031 7611 37065
rect 7645 37031 7683 37065
rect 7717 37031 7750 37065
rect 2543 36962 7750 37031
rect 8044 37101 8050 37135
rect 8084 37125 8224 37135
rect 8084 37101 8184 37125
rect 8044 37091 8184 37101
rect 8218 37091 8224 37125
rect 8044 37063 8224 37091
rect 8044 37029 8050 37063
rect 8084 37053 8224 37063
rect 8084 37029 8184 37053
rect 8044 37019 8184 37029
rect 8218 37019 8224 37053
rect 8044 36991 8224 37019
rect 2543 36957 2795 36962
tri 2795 36957 2800 36962 nw
rect 8044 36957 8050 36991
rect 8084 36981 8224 36991
rect 8084 36957 8184 36981
rect 2543 36947 2785 36957
tri 2785 36947 2795 36957 nw
rect 8044 36947 8184 36957
rect 8218 36947 8224 36981
rect 2543 36919 2757 36947
tri 2757 36919 2785 36947 nw
rect 8044 36919 8224 36947
rect 2543 36885 2723 36919
tri 2723 36885 2757 36919 nw
rect 8044 36885 8050 36919
rect 8084 36909 8224 36919
rect 8084 36885 8184 36909
rect 2543 36875 2713 36885
tri 2713 36875 2723 36885 nw
rect 8044 36875 8184 36885
rect 8218 36875 8224 36909
rect 2543 35157 2712 36875
tri 2712 36874 2713 36875 nw
rect 8044 36847 8224 36875
rect 8044 36813 8050 36847
rect 8084 36837 8224 36847
rect 8084 36813 8184 36837
rect 8044 36803 8184 36813
rect 8218 36803 8224 36837
rect 8044 36775 8224 36803
rect 8044 36741 8050 36775
rect 8084 36765 8224 36775
rect 8084 36741 8184 36765
rect 8044 36731 8184 36741
rect 8218 36731 8224 36765
rect 2824 36720 2942 36726
rect 2876 36668 2890 36720
rect 2824 36651 2942 36668
rect 2876 36599 2890 36651
rect 2824 36582 2942 36599
rect 2876 36530 2890 36582
rect 2824 36513 2942 36530
rect 2876 36461 2890 36513
rect 2824 36444 2942 36461
rect 2876 36422 2890 36444
rect 2824 36375 2830 36392
rect 2936 36375 2942 36392
rect 2824 36306 2830 36323
rect 2936 36306 2942 36323
rect 2824 36236 2830 36254
rect 2936 36236 2942 36254
rect 2824 36166 2830 36184
rect 2936 36166 2942 36184
rect 2824 35380 2830 36114
rect 2936 35380 2942 36114
rect 2824 35368 2942 35380
rect 3101 36714 3219 36726
rect 3101 36680 3107 36714
rect 3141 36680 3179 36714
rect 3213 36680 3219 36714
rect 3101 36641 3219 36680
rect 3101 36607 3107 36641
rect 3141 36607 3179 36641
rect 3213 36607 3219 36641
rect 3101 36568 3219 36607
rect 3101 36534 3107 36568
rect 3141 36534 3179 36568
rect 3213 36534 3219 36568
rect 3101 36495 3219 36534
rect 3101 36461 3107 36495
rect 3141 36461 3179 36495
rect 3213 36461 3219 36495
rect 3101 36422 3219 36461
rect 3101 35982 3107 36422
rect 3213 35982 3219 36422
rect 3101 35913 3107 35930
rect 3213 35913 3219 35930
rect 3101 35844 3107 35861
rect 3213 35844 3219 35861
rect 3101 35775 3107 35792
rect 3213 35775 3219 35792
rect 3101 35706 3107 35723
rect 3213 35706 3219 35723
rect 3101 35636 3107 35654
rect 3213 35636 3219 35654
rect 3101 35566 3107 35584
rect 3213 35566 3219 35584
rect 3101 35496 3107 35514
rect 3213 35496 3219 35514
rect 3101 35426 3107 35444
rect 3213 35426 3219 35444
rect 3153 35374 3167 35380
rect 3101 35368 3219 35374
rect 3378 36720 3496 36726
rect 3430 36668 3444 36720
rect 3378 36651 3496 36668
rect 3430 36599 3444 36651
rect 3378 36582 3496 36599
rect 3430 36530 3444 36582
rect 3378 36513 3496 36530
rect 3430 36461 3444 36513
rect 3378 36444 3496 36461
rect 3430 36422 3444 36444
rect 3378 36375 3384 36392
rect 3490 36375 3496 36392
rect 3378 36306 3384 36323
rect 3490 36306 3496 36323
rect 3378 36236 3384 36254
rect 3490 36236 3496 36254
rect 3378 36166 3384 36184
rect 3490 36166 3496 36184
rect 3378 35380 3384 36114
rect 3490 35380 3496 36114
rect 3378 35368 3496 35380
rect 3655 36714 3773 36726
rect 3655 36680 3661 36714
rect 3695 36680 3733 36714
rect 3767 36680 3773 36714
rect 3655 36641 3773 36680
rect 3655 36607 3661 36641
rect 3695 36607 3733 36641
rect 3767 36607 3773 36641
rect 3655 36568 3773 36607
rect 3655 36534 3661 36568
rect 3695 36534 3733 36568
rect 3767 36534 3773 36568
rect 3655 36495 3773 36534
rect 3655 36461 3661 36495
rect 3695 36461 3733 36495
rect 3767 36461 3773 36495
rect 3655 36422 3773 36461
rect 3655 35982 3661 36422
rect 3767 35982 3773 36422
rect 3655 35913 3661 35930
rect 3767 35913 3773 35930
rect 3655 35844 3661 35861
rect 3767 35844 3773 35861
rect 3655 35775 3661 35792
rect 3767 35775 3773 35792
rect 3655 35706 3661 35723
rect 3767 35706 3773 35723
rect 3655 35636 3661 35654
rect 3767 35636 3773 35654
rect 3655 35566 3661 35584
rect 3767 35566 3773 35584
rect 3655 35496 3661 35514
rect 3767 35496 3773 35514
rect 3655 35426 3661 35444
rect 3767 35426 3773 35444
rect 3707 35374 3721 35380
rect 3655 35368 3773 35374
rect 3932 36720 4050 36726
rect 3984 36668 3998 36720
rect 3932 36651 4050 36668
rect 3984 36599 3998 36651
rect 3932 36582 4050 36599
rect 3984 36530 3998 36582
rect 3932 36513 4050 36530
rect 3984 36461 3998 36513
rect 3932 36444 4050 36461
rect 3984 36422 3998 36444
rect 3932 36375 3938 36392
rect 4044 36375 4050 36392
rect 3932 36306 3938 36323
rect 4044 36306 4050 36323
rect 3932 36236 3938 36254
rect 4044 36236 4050 36254
rect 3932 36166 3938 36184
rect 4044 36166 4050 36184
rect 3932 35380 3938 36114
rect 4044 35380 4050 36114
rect 3932 35368 4050 35380
rect 4209 36714 4327 36726
rect 4209 36680 4215 36714
rect 4249 36680 4287 36714
rect 4321 36680 4327 36714
rect 4209 36641 4327 36680
rect 4209 36607 4215 36641
rect 4249 36607 4287 36641
rect 4321 36607 4327 36641
rect 4209 36568 4327 36607
rect 4209 36534 4215 36568
rect 4249 36534 4287 36568
rect 4321 36534 4327 36568
rect 4209 36495 4327 36534
rect 4209 36461 4215 36495
rect 4249 36461 4287 36495
rect 4321 36461 4327 36495
rect 4209 36422 4327 36461
rect 4209 35982 4215 36422
rect 4321 35982 4327 36422
rect 4209 35913 4215 35930
rect 4321 35913 4327 35930
rect 4209 35844 4215 35861
rect 4321 35844 4327 35861
rect 4209 35775 4215 35792
rect 4321 35775 4327 35792
rect 4209 35706 4215 35723
rect 4321 35706 4327 35723
rect 4209 35636 4215 35654
rect 4321 35636 4327 35654
rect 4209 35566 4215 35584
rect 4321 35566 4327 35584
rect 4209 35496 4215 35514
rect 4321 35496 4327 35514
rect 4209 35426 4215 35444
rect 4321 35426 4327 35444
rect 4261 35374 4275 35380
rect 4209 35368 4327 35374
rect 4486 36720 4604 36726
rect 4538 36668 4552 36720
rect 4486 36651 4604 36668
rect 4538 36599 4552 36651
rect 4486 36582 4604 36599
rect 4538 36530 4552 36582
rect 4486 36513 4604 36530
rect 4538 36461 4552 36513
rect 4486 36444 4604 36461
rect 4538 36422 4552 36444
rect 4486 36375 4492 36392
rect 4598 36375 4604 36392
rect 4486 36306 4492 36323
rect 4598 36306 4604 36323
rect 4486 36236 4492 36254
rect 4598 36236 4604 36254
rect 4486 36166 4492 36184
rect 4598 36166 4604 36184
rect 4486 35380 4492 36114
rect 4598 35380 4604 36114
rect 4486 35368 4604 35380
rect 4763 36714 4881 36726
rect 4763 36680 4769 36714
rect 4803 36680 4841 36714
rect 4875 36680 4881 36714
rect 4763 36641 4881 36680
rect 4763 36607 4769 36641
rect 4803 36607 4841 36641
rect 4875 36607 4881 36641
rect 4763 36568 4881 36607
rect 4763 36534 4769 36568
rect 4803 36534 4841 36568
rect 4875 36534 4881 36568
rect 4763 36495 4881 36534
rect 4763 36461 4769 36495
rect 4803 36461 4841 36495
rect 4875 36461 4881 36495
rect 4763 36422 4881 36461
rect 4763 35982 4769 36422
rect 4875 35982 4881 36422
rect 4763 35913 4769 35930
rect 4875 35913 4881 35930
rect 4763 35844 4769 35861
rect 4875 35844 4881 35861
rect 4763 35775 4769 35792
rect 4875 35775 4881 35792
rect 4763 35706 4769 35723
rect 4875 35706 4881 35723
rect 4763 35636 4769 35654
rect 4875 35636 4881 35654
rect 4763 35566 4769 35584
rect 4875 35566 4881 35584
rect 4763 35496 4769 35514
rect 4875 35496 4881 35514
rect 4763 35426 4769 35444
rect 4875 35426 4881 35444
rect 4815 35374 4829 35380
rect 4763 35368 4881 35374
rect 5040 36720 5158 36726
rect 5092 36668 5106 36720
rect 5040 36651 5158 36668
rect 5092 36599 5106 36651
rect 5040 36582 5158 36599
rect 5092 36530 5106 36582
rect 5040 36513 5158 36530
rect 5092 36461 5106 36513
rect 5040 36444 5158 36461
rect 5092 36422 5106 36444
rect 5040 36375 5046 36392
rect 5152 36375 5158 36392
rect 5040 36306 5046 36323
rect 5152 36306 5158 36323
rect 5040 36236 5046 36254
rect 5152 36236 5158 36254
rect 5040 36166 5046 36184
rect 5152 36166 5158 36184
rect 5040 35380 5046 36114
rect 5152 35380 5158 36114
rect 5040 35368 5158 35380
rect 5317 36714 5435 36726
rect 5317 36680 5323 36714
rect 5357 36680 5395 36714
rect 5429 36680 5435 36714
rect 5317 36641 5435 36680
rect 5317 36607 5323 36641
rect 5357 36607 5395 36641
rect 5429 36607 5435 36641
rect 5317 36568 5435 36607
rect 5317 36534 5323 36568
rect 5357 36534 5395 36568
rect 5429 36534 5435 36568
rect 5317 36495 5435 36534
rect 5317 36461 5323 36495
rect 5357 36461 5395 36495
rect 5429 36461 5435 36495
rect 5317 36422 5435 36461
rect 5317 35982 5323 36422
rect 5429 35982 5435 36422
rect 5317 35913 5323 35930
rect 5429 35913 5435 35930
rect 5317 35844 5323 35861
rect 5429 35844 5435 35861
rect 5317 35775 5323 35792
rect 5429 35775 5435 35792
rect 5317 35706 5323 35723
rect 5429 35706 5435 35723
rect 5317 35636 5323 35654
rect 5429 35636 5435 35654
rect 5317 35566 5323 35584
rect 5429 35566 5435 35584
rect 5317 35496 5323 35514
rect 5429 35496 5435 35514
rect 5317 35426 5323 35444
rect 5429 35426 5435 35444
rect 5369 35374 5383 35380
rect 5317 35368 5435 35374
rect 5594 36720 5712 36726
rect 5646 36668 5660 36720
rect 5594 36651 5712 36668
rect 5646 36599 5660 36651
rect 5594 36582 5712 36599
rect 5646 36530 5660 36582
rect 5594 36513 5712 36530
rect 5646 36461 5660 36513
rect 5594 36444 5712 36461
rect 5646 36422 5660 36444
rect 5594 36375 5600 36392
rect 5706 36375 5712 36392
rect 5594 36306 5600 36323
rect 5706 36306 5712 36323
rect 5594 36236 5600 36254
rect 5706 36236 5712 36254
rect 5594 36166 5600 36184
rect 5706 36166 5712 36184
rect 5594 35380 5600 36114
rect 5706 35380 5712 36114
rect 5594 35368 5712 35380
rect 5871 36714 5989 36726
rect 5871 36680 5877 36714
rect 5911 36680 5949 36714
rect 5983 36680 5989 36714
rect 5871 36641 5989 36680
rect 5871 36607 5877 36641
rect 5911 36607 5949 36641
rect 5983 36607 5989 36641
rect 5871 36568 5989 36607
rect 5871 36534 5877 36568
rect 5911 36534 5949 36568
rect 5983 36534 5989 36568
rect 5871 36495 5989 36534
rect 5871 36461 5877 36495
rect 5911 36461 5949 36495
rect 5983 36461 5989 36495
rect 5871 36422 5989 36461
rect 5871 35982 5877 36422
rect 5983 35982 5989 36422
rect 5871 35913 5877 35930
rect 5983 35913 5989 35930
rect 5871 35844 5877 35861
rect 5983 35844 5989 35861
rect 5871 35775 5877 35792
rect 5983 35775 5989 35792
rect 5871 35706 5877 35723
rect 5983 35706 5989 35723
rect 5871 35636 5877 35654
rect 5983 35636 5989 35654
rect 5871 35566 5877 35584
rect 5983 35566 5989 35584
rect 5871 35496 5877 35514
rect 5983 35496 5989 35514
rect 5871 35426 5877 35444
rect 5983 35426 5989 35444
rect 5923 35374 5937 35380
rect 5871 35368 5989 35374
rect 6148 36720 6266 36726
rect 6200 36668 6214 36720
rect 6148 36651 6266 36668
rect 6200 36599 6214 36651
rect 6148 36582 6266 36599
rect 6200 36530 6214 36582
rect 6148 36513 6266 36530
rect 6200 36461 6214 36513
rect 6148 36444 6266 36461
rect 6200 36422 6214 36444
rect 6148 36375 6154 36392
rect 6260 36375 6266 36392
rect 6148 36306 6154 36323
rect 6260 36306 6266 36323
rect 6148 36236 6154 36254
rect 6260 36236 6266 36254
rect 6148 36166 6154 36184
rect 6260 36166 6266 36184
rect 6148 35380 6154 36114
rect 6260 35380 6266 36114
rect 6148 35368 6266 35380
rect 6425 36714 6543 36726
rect 6425 36680 6431 36714
rect 6465 36680 6503 36714
rect 6537 36680 6543 36714
rect 6425 36641 6543 36680
rect 6425 36607 6431 36641
rect 6465 36607 6503 36641
rect 6537 36607 6543 36641
rect 6425 36568 6543 36607
rect 6425 36534 6431 36568
rect 6465 36534 6503 36568
rect 6537 36534 6543 36568
rect 6425 36495 6543 36534
rect 6425 36461 6431 36495
rect 6465 36461 6503 36495
rect 6537 36461 6543 36495
rect 6425 36422 6543 36461
rect 6425 35982 6431 36422
rect 6537 35982 6543 36422
rect 6425 35913 6431 35930
rect 6537 35913 6543 35930
rect 6425 35844 6431 35861
rect 6537 35844 6543 35861
rect 6425 35775 6431 35792
rect 6537 35775 6543 35792
rect 6425 35706 6431 35723
rect 6537 35706 6543 35723
rect 6425 35636 6431 35654
rect 6537 35636 6543 35654
rect 6425 35566 6431 35584
rect 6537 35566 6543 35584
rect 6425 35496 6431 35514
rect 6537 35496 6543 35514
rect 6425 35426 6431 35444
rect 6537 35426 6543 35444
rect 6477 35374 6491 35380
rect 6425 35368 6543 35374
rect 6702 36720 6820 36726
rect 6754 36668 6768 36720
rect 6702 36651 6820 36668
rect 6754 36599 6768 36651
rect 6702 36582 6820 36599
rect 6754 36530 6768 36582
rect 6702 36513 6820 36530
rect 6754 36461 6768 36513
rect 6702 36444 6820 36461
rect 6754 36422 6768 36444
rect 6702 36375 6708 36392
rect 6814 36375 6820 36392
rect 6702 36306 6708 36323
rect 6814 36306 6820 36323
rect 6702 36236 6708 36254
rect 6814 36236 6820 36254
rect 6702 36166 6708 36184
rect 6814 36166 6820 36184
rect 6702 35380 6708 36114
rect 6814 35380 6820 36114
rect 6702 35368 6820 35380
rect 6979 36714 7097 36726
rect 6979 36680 6985 36714
rect 7019 36680 7057 36714
rect 7091 36680 7097 36714
rect 6979 36641 7097 36680
rect 6979 36607 6985 36641
rect 7019 36607 7057 36641
rect 7091 36607 7097 36641
rect 6979 36568 7097 36607
rect 6979 36534 6985 36568
rect 7019 36534 7057 36568
rect 7091 36534 7097 36568
rect 6979 36495 7097 36534
rect 6979 36461 6985 36495
rect 7019 36461 7057 36495
rect 7091 36461 7097 36495
rect 6979 36422 7097 36461
rect 6979 35982 6985 36422
rect 7091 35982 7097 36422
rect 6979 35913 6985 35930
rect 7091 35913 7097 35930
rect 6979 35844 6985 35861
rect 7091 35844 7097 35861
rect 6979 35775 6985 35792
rect 7091 35775 7097 35792
rect 6979 35706 6985 35723
rect 7091 35706 7097 35723
rect 6979 35636 6985 35654
rect 7091 35636 7097 35654
rect 6979 35566 6985 35584
rect 7091 35566 7097 35584
rect 6979 35496 6985 35514
rect 7091 35496 7097 35514
rect 6979 35426 6985 35444
rect 7091 35426 7097 35444
rect 7031 35374 7045 35380
rect 6979 35368 7097 35374
rect 7256 36720 7374 36726
rect 7308 36668 7322 36720
rect 7256 36651 7374 36668
rect 7308 36599 7322 36651
rect 7256 36582 7374 36599
rect 7308 36530 7322 36582
rect 7256 36513 7374 36530
rect 7308 36461 7322 36513
rect 7256 36444 7374 36461
rect 7308 36422 7322 36444
rect 7256 36375 7262 36392
rect 7368 36375 7374 36392
rect 7256 36306 7262 36323
rect 7368 36306 7374 36323
rect 7256 36236 7262 36254
rect 7368 36236 7374 36254
rect 7256 36166 7262 36184
rect 7368 36166 7374 36184
rect 7256 35380 7262 36114
rect 7368 35380 7374 36114
rect 7256 35368 7374 35380
rect 7533 36714 7651 36726
rect 7533 36680 7539 36714
rect 7573 36680 7611 36714
rect 7645 36680 7651 36714
rect 7533 36641 7651 36680
rect 7533 36607 7539 36641
rect 7573 36607 7611 36641
rect 7645 36607 7651 36641
rect 7533 36568 7651 36607
rect 7533 36534 7539 36568
rect 7573 36534 7611 36568
rect 7645 36534 7651 36568
rect 7533 36495 7651 36534
rect 7533 36461 7539 36495
rect 7573 36461 7611 36495
rect 7645 36461 7651 36495
rect 7533 36422 7651 36461
rect 7533 35982 7539 36422
rect 7645 35982 7651 36422
rect 7533 35913 7539 35930
rect 7645 35913 7651 35930
rect 7533 35844 7539 35861
rect 7645 35844 7651 35861
rect 7533 35775 7539 35792
rect 7645 35775 7651 35792
rect 7533 35706 7539 35723
rect 7645 35706 7651 35723
rect 7533 35636 7539 35654
rect 7645 35636 7651 35654
rect 7533 35566 7539 35584
rect 7645 35566 7651 35584
rect 7533 35496 7539 35514
rect 7645 35496 7651 35514
rect 7533 35426 7539 35444
rect 7645 35426 7651 35444
rect 7585 35374 7599 35380
rect 7533 35368 7651 35374
rect 7810 36720 7928 36726
rect 7862 36668 7876 36720
rect 7810 36651 7928 36668
rect 7862 36599 7876 36651
rect 7810 36582 7928 36599
rect 7862 36530 7876 36582
rect 7810 36513 7928 36530
rect 7862 36461 7876 36513
rect 7810 36444 7928 36461
rect 7862 36422 7876 36444
rect 7810 36375 7816 36392
rect 7922 36375 7928 36392
rect 7810 36306 7816 36323
rect 7922 36306 7928 36323
rect 7810 36236 7816 36254
rect 7922 36236 7928 36254
rect 7810 36166 7816 36184
rect 7922 36166 7928 36184
rect 7810 35380 7816 36114
rect 7922 35380 7928 36114
rect 7810 35368 7928 35380
rect 8044 36724 8224 36731
rect 8044 36672 8047 36724
rect 8099 36672 8169 36724
rect 8221 36672 8224 36724
rect 8044 36669 8050 36672
rect 8084 36669 8184 36672
rect 8044 36659 8184 36669
rect 8218 36659 8224 36672
rect 8044 36655 8224 36659
rect 8044 36603 8047 36655
rect 8099 36603 8169 36655
rect 8221 36603 8224 36655
rect 8044 36597 8050 36603
rect 8084 36597 8184 36603
rect 8044 36587 8184 36597
rect 8218 36587 8224 36603
rect 8044 36586 8224 36587
rect 8044 36534 8047 36586
rect 8099 36534 8169 36586
rect 8221 36534 8224 36586
rect 8044 36525 8050 36534
rect 8084 36525 8184 36534
rect 8044 36517 8184 36525
rect 8218 36517 8224 36534
rect 8044 36465 8047 36517
rect 8099 36465 8169 36517
rect 8221 36465 8224 36517
rect 8044 36453 8050 36465
rect 8084 36453 8184 36465
rect 8044 36448 8184 36453
rect 8218 36448 8224 36465
rect 8044 36396 8047 36448
rect 8099 36396 8169 36448
rect 8221 36396 8224 36448
rect 8044 36381 8050 36396
rect 8084 36381 8184 36396
rect 8044 36378 8184 36381
rect 8218 36378 8224 36396
rect 8044 36326 8047 36378
rect 8099 36326 8169 36378
rect 8221 36326 8224 36378
rect 8044 36309 8050 36326
rect 8084 36309 8184 36326
rect 8044 36308 8184 36309
rect 8218 36308 8224 36326
rect 8044 36256 8047 36308
rect 8099 36256 8169 36308
rect 8221 36256 8224 36308
rect 8044 36238 8050 36256
rect 8084 36238 8184 36256
rect 8218 36238 8224 36256
rect 8044 36186 8047 36238
rect 8099 36186 8169 36238
rect 8221 36186 8224 36238
rect 8044 36168 8050 36186
rect 8084 36168 8184 36186
rect 8218 36168 8224 36186
rect 8044 36116 8047 36168
rect 8099 36116 8169 36168
rect 8221 36116 8224 36168
rect 8044 36093 8050 36116
rect 8084 36093 8184 36116
rect 8044 36083 8184 36093
rect 8218 36083 8224 36116
rect 8044 36055 8224 36083
rect 8044 36021 8050 36055
rect 8084 36045 8224 36055
rect 8084 36021 8184 36045
rect 8044 36011 8184 36021
rect 8218 36011 8224 36045
rect 8044 35983 8224 36011
rect 8044 35949 8050 35983
rect 8084 35973 8224 35983
rect 8084 35949 8184 35973
rect 8044 35939 8184 35949
rect 8218 35939 8224 35973
rect 8044 35911 8224 35939
rect 8044 35877 8050 35911
rect 8084 35901 8224 35911
rect 8084 35877 8184 35901
rect 8044 35867 8184 35877
rect 8218 35867 8224 35901
rect 8044 35839 8224 35867
rect 8044 35805 8050 35839
rect 8084 35829 8224 35839
rect 8084 35805 8184 35829
rect 8044 35795 8184 35805
rect 8218 35795 8224 35829
rect 8044 35767 8224 35795
rect 8044 35733 8050 35767
rect 8084 35757 8224 35767
rect 8084 35733 8184 35757
rect 8044 35723 8184 35733
rect 8218 35723 8224 35757
rect 8044 35695 8224 35723
rect 8044 35661 8050 35695
rect 8084 35685 8224 35695
rect 8084 35661 8184 35685
rect 8044 35651 8184 35661
rect 8218 35651 8224 35685
rect 8044 35623 8224 35651
rect 8044 35589 8050 35623
rect 8084 35613 8224 35623
rect 8084 35589 8184 35613
rect 8044 35579 8184 35589
rect 8218 35579 8224 35613
rect 8044 35551 8224 35579
rect 8044 35517 8050 35551
rect 8084 35541 8224 35551
rect 8084 35517 8184 35541
rect 8044 35507 8184 35517
rect 8218 35507 8224 35541
rect 8044 35479 8224 35507
rect 8044 35445 8050 35479
rect 8084 35469 8224 35479
rect 8084 35445 8184 35469
rect 8044 35435 8184 35445
rect 8218 35435 8224 35469
rect 8044 35407 8224 35435
rect 8044 35373 8050 35407
rect 8084 35397 8224 35407
rect 8084 35373 8184 35397
rect 8044 35363 8184 35373
rect 8218 35363 8224 35397
rect 8044 35335 8224 35363
rect 8044 35301 8050 35335
rect 8084 35325 8224 35335
rect 8084 35301 8184 35325
rect 8044 35291 8184 35301
rect 8218 35291 8224 35325
rect 8044 35263 8224 35291
rect 8044 35229 8050 35263
rect 8084 35253 8224 35263
rect 8084 35229 8184 35253
rect 8044 35219 8184 35229
rect 8218 35219 8224 35253
rect 8044 35191 8224 35219
tri 2712 35157 2721 35166 sw
rect 8044 35157 8050 35191
rect 8084 35181 8224 35191
rect 8084 35157 8184 35181
rect 2543 35147 2721 35157
tri 2721 35147 2731 35157 sw
rect 8044 35147 8184 35157
rect 8218 35147 8224 35181
rect 2543 35134 2731 35147
tri 2731 35134 2744 35147 sw
rect 2543 35099 7750 35134
rect 2543 35065 3035 35099
rect 3069 35065 3108 35099
rect 3142 35065 3181 35099
rect 3215 35065 3254 35099
rect 3288 35065 3327 35099
rect 3361 35065 3400 35099
rect 3434 35065 3473 35099
rect 3507 35065 3546 35099
rect 3580 35065 3619 35099
rect 3653 35065 3692 35099
rect 3726 35065 3765 35099
rect 3799 35065 3838 35099
rect 3872 35065 3911 35099
rect 3945 35065 3984 35099
rect 4018 35065 4057 35099
rect 4091 35065 4130 35099
rect 4164 35065 4203 35099
rect 4237 35065 4276 35099
rect 4310 35065 4349 35099
rect 4383 35065 4422 35099
rect 4456 35065 4495 35099
rect 4529 35065 4568 35099
rect 4602 35065 4641 35099
rect 4675 35065 4714 35099
rect 4748 35065 4787 35099
rect 4821 35065 4860 35099
rect 4894 35065 4933 35099
rect 4967 35065 5006 35099
rect 5040 35065 5079 35099
rect 5113 35065 5152 35099
rect 5186 35065 5225 35099
rect 5259 35065 5298 35099
rect 5332 35065 5371 35099
rect 5405 35065 5444 35099
rect 5478 35065 5517 35099
rect 5551 35065 5590 35099
rect 5624 35065 5663 35099
rect 5697 35065 5736 35099
rect 5770 35065 5809 35099
rect 5843 35065 5882 35099
rect 5916 35065 5955 35099
rect 5989 35065 6027 35099
rect 6061 35065 6099 35099
rect 6133 35065 6171 35099
rect 6205 35065 6243 35099
rect 6277 35065 6315 35099
rect 6349 35065 6387 35099
rect 6421 35065 6459 35099
rect 6493 35065 6531 35099
rect 6565 35065 6603 35099
rect 6637 35065 6675 35099
rect 6709 35065 6747 35099
rect 6781 35065 6819 35099
rect 6853 35065 6891 35099
rect 6925 35065 6963 35099
rect 6997 35065 7035 35099
rect 7069 35065 7107 35099
rect 7141 35065 7179 35099
rect 7213 35065 7251 35099
rect 7285 35065 7323 35099
rect 7357 35065 7395 35099
rect 7429 35065 7467 35099
rect 7501 35065 7539 35099
rect 7573 35065 7611 35099
rect 7645 35065 7683 35099
rect 7717 35065 7750 35099
rect 2543 35028 7750 35065
rect 8044 35119 8224 35147
rect 8044 35085 8050 35119
rect 8084 35109 8224 35119
rect 8084 35085 8184 35109
rect 8044 35075 8184 35085
rect 8218 35075 8224 35109
rect 8044 35047 8224 35075
rect 2543 35013 2751 35028
tri 2751 35013 2766 35028 nw
rect 8044 35013 8050 35047
rect 8084 35037 8224 35047
rect 8084 35013 8184 35037
rect 2543 35003 2741 35013
tri 2741 35003 2751 35013 nw
rect 8044 35003 8184 35013
rect 8218 35003 8224 35037
rect 2543 34975 2713 35003
tri 2713 34975 2741 35003 nw
rect 8044 34975 8224 35003
rect 2543 33141 2712 34975
tri 2712 34974 2713 34975 nw
rect 8044 34941 8050 34975
rect 8084 34965 8224 34975
rect 8084 34941 8184 34965
rect 8044 34931 8184 34941
rect 8218 34931 8224 34965
rect 8044 34903 8224 34931
rect 8044 34869 8050 34903
rect 8084 34893 8224 34903
rect 8084 34869 8184 34893
rect 8044 34859 8184 34869
rect 8218 34859 8224 34893
rect 8044 34831 8224 34859
rect 8044 34797 8050 34831
rect 8084 34821 8224 34831
rect 8084 34797 8184 34821
rect 8044 34787 8184 34797
rect 8218 34787 8224 34821
rect 8044 34759 8224 34787
rect 2824 34720 2942 34726
rect 2876 34668 2890 34720
rect 2824 34651 2942 34668
rect 2876 34599 2890 34651
rect 2824 34582 2942 34599
rect 2876 34530 2890 34582
rect 2824 34513 2942 34530
rect 2876 34461 2890 34513
rect 2824 34444 2942 34461
rect 2876 34422 2890 34444
rect 2824 34375 2830 34392
rect 2936 34375 2942 34392
rect 2824 34306 2830 34323
rect 2936 34306 2942 34323
rect 2824 34236 2830 34254
rect 2936 34236 2942 34254
rect 2824 34166 2830 34184
rect 2936 34166 2942 34184
rect 2824 33380 2830 34114
rect 2936 33380 2942 34114
rect 2824 33368 2942 33380
rect 3101 34714 3219 34726
rect 3101 34680 3107 34714
rect 3141 34680 3179 34714
rect 3213 34680 3219 34714
rect 3101 34641 3219 34680
rect 3101 34607 3107 34641
rect 3141 34607 3179 34641
rect 3213 34607 3219 34641
rect 3101 34568 3219 34607
rect 3101 34534 3107 34568
rect 3141 34534 3179 34568
rect 3213 34534 3219 34568
rect 3101 34495 3219 34534
rect 3101 34461 3107 34495
rect 3141 34461 3179 34495
rect 3213 34461 3219 34495
rect 3101 34422 3219 34461
rect 3101 33982 3107 34422
rect 3213 33982 3219 34422
rect 3101 33913 3107 33930
rect 3213 33913 3219 33930
rect 3101 33844 3107 33861
rect 3213 33844 3219 33861
rect 3101 33775 3107 33792
rect 3213 33775 3219 33792
rect 3101 33706 3107 33723
rect 3213 33706 3219 33723
rect 3101 33636 3107 33654
rect 3213 33636 3219 33654
rect 3101 33566 3107 33584
rect 3213 33566 3219 33584
rect 3101 33496 3107 33514
rect 3213 33496 3219 33514
rect 3101 33426 3107 33444
rect 3213 33426 3219 33444
rect 3153 33374 3167 33380
rect 3101 33368 3219 33374
rect 3378 34720 3496 34726
rect 3430 34668 3444 34720
rect 3378 34651 3496 34668
rect 3430 34599 3444 34651
rect 3378 34582 3496 34599
rect 3430 34530 3444 34582
rect 3378 34513 3496 34530
rect 3430 34461 3444 34513
rect 3378 34444 3496 34461
rect 3430 34422 3444 34444
rect 3378 34375 3384 34392
rect 3490 34375 3496 34392
rect 3378 34306 3384 34323
rect 3490 34306 3496 34323
rect 3378 34236 3384 34254
rect 3490 34236 3496 34254
rect 3378 34166 3384 34184
rect 3490 34166 3496 34184
rect 3378 33380 3384 34114
rect 3490 33380 3496 34114
rect 3378 33368 3496 33380
rect 3655 34714 3773 34726
rect 3655 34680 3661 34714
rect 3695 34680 3733 34714
rect 3767 34680 3773 34714
rect 3655 34641 3773 34680
rect 3655 34607 3661 34641
rect 3695 34607 3733 34641
rect 3767 34607 3773 34641
rect 3655 34568 3773 34607
rect 3655 34534 3661 34568
rect 3695 34534 3733 34568
rect 3767 34534 3773 34568
rect 3655 34495 3773 34534
rect 3655 34461 3661 34495
rect 3695 34461 3733 34495
rect 3767 34461 3773 34495
rect 3655 34422 3773 34461
rect 3655 33982 3661 34422
rect 3767 33982 3773 34422
rect 3655 33913 3661 33930
rect 3767 33913 3773 33930
rect 3655 33844 3661 33861
rect 3767 33844 3773 33861
rect 3655 33775 3661 33792
rect 3767 33775 3773 33792
rect 3655 33706 3661 33723
rect 3767 33706 3773 33723
rect 3655 33636 3661 33654
rect 3767 33636 3773 33654
rect 3655 33566 3661 33584
rect 3767 33566 3773 33584
rect 3655 33496 3661 33514
rect 3767 33496 3773 33514
rect 3655 33426 3661 33444
rect 3767 33426 3773 33444
rect 3707 33374 3721 33380
rect 3655 33368 3773 33374
rect 3932 34720 4050 34726
rect 3984 34668 3998 34720
rect 3932 34651 4050 34668
rect 3984 34599 3998 34651
rect 3932 34582 4050 34599
rect 3984 34530 3998 34582
rect 3932 34513 4050 34530
rect 3984 34461 3998 34513
rect 3932 34444 4050 34461
rect 3984 34422 3998 34444
rect 3932 34375 3938 34392
rect 4044 34375 4050 34392
rect 3932 34306 3938 34323
rect 4044 34306 4050 34323
rect 3932 34236 3938 34254
rect 4044 34236 4050 34254
rect 3932 34166 3938 34184
rect 4044 34166 4050 34184
rect 3932 33380 3938 34114
rect 4044 33380 4050 34114
rect 3932 33368 4050 33380
rect 4209 34714 4327 34726
rect 4209 34680 4215 34714
rect 4249 34680 4287 34714
rect 4321 34680 4327 34714
rect 4209 34641 4327 34680
rect 4209 34607 4215 34641
rect 4249 34607 4287 34641
rect 4321 34607 4327 34641
rect 4209 34568 4327 34607
rect 4209 34534 4215 34568
rect 4249 34534 4287 34568
rect 4321 34534 4327 34568
rect 4209 34495 4327 34534
rect 4209 34461 4215 34495
rect 4249 34461 4287 34495
rect 4321 34461 4327 34495
rect 4209 34422 4327 34461
rect 4209 33982 4215 34422
rect 4321 33982 4327 34422
rect 4209 33913 4215 33930
rect 4321 33913 4327 33930
rect 4209 33844 4215 33861
rect 4321 33844 4327 33861
rect 4209 33775 4215 33792
rect 4321 33775 4327 33792
rect 4209 33706 4215 33723
rect 4321 33706 4327 33723
rect 4209 33636 4215 33654
rect 4321 33636 4327 33654
rect 4209 33566 4215 33584
rect 4321 33566 4327 33584
rect 4209 33496 4215 33514
rect 4321 33496 4327 33514
rect 4209 33426 4215 33444
rect 4321 33426 4327 33444
rect 4261 33374 4275 33380
rect 4209 33368 4327 33374
rect 4486 34720 4604 34726
rect 4538 34668 4552 34720
rect 4486 34651 4604 34668
rect 4538 34599 4552 34651
rect 4486 34582 4604 34599
rect 4538 34530 4552 34582
rect 4486 34513 4604 34530
rect 4538 34461 4552 34513
rect 4486 34444 4604 34461
rect 4538 34422 4552 34444
rect 4486 34375 4492 34392
rect 4598 34375 4604 34392
rect 4486 34306 4492 34323
rect 4598 34306 4604 34323
rect 4486 34236 4492 34254
rect 4598 34236 4604 34254
rect 4486 34166 4492 34184
rect 4598 34166 4604 34184
rect 4486 33380 4492 34114
rect 4598 33380 4604 34114
rect 4486 33368 4604 33380
rect 4763 34714 4881 34726
rect 4763 34680 4769 34714
rect 4803 34680 4841 34714
rect 4875 34680 4881 34714
rect 4763 34641 4881 34680
rect 4763 34607 4769 34641
rect 4803 34607 4841 34641
rect 4875 34607 4881 34641
rect 4763 34568 4881 34607
rect 4763 34534 4769 34568
rect 4803 34534 4841 34568
rect 4875 34534 4881 34568
rect 4763 34495 4881 34534
rect 4763 34461 4769 34495
rect 4803 34461 4841 34495
rect 4875 34461 4881 34495
rect 4763 34422 4881 34461
rect 4763 33982 4769 34422
rect 4875 33982 4881 34422
rect 4763 33913 4769 33930
rect 4875 33913 4881 33930
rect 4763 33844 4769 33861
rect 4875 33844 4881 33861
rect 4763 33775 4769 33792
rect 4875 33775 4881 33792
rect 4763 33706 4769 33723
rect 4875 33706 4881 33723
rect 4763 33636 4769 33654
rect 4875 33636 4881 33654
rect 4763 33566 4769 33584
rect 4875 33566 4881 33584
rect 4763 33496 4769 33514
rect 4875 33496 4881 33514
rect 4763 33426 4769 33444
rect 4875 33426 4881 33444
rect 4815 33374 4829 33380
rect 4763 33368 4881 33374
rect 5040 34720 5158 34726
rect 5092 34668 5106 34720
rect 5040 34651 5158 34668
rect 5092 34599 5106 34651
rect 5040 34582 5158 34599
rect 5092 34530 5106 34582
rect 5040 34513 5158 34530
rect 5092 34461 5106 34513
rect 5040 34444 5158 34461
rect 5092 34422 5106 34444
rect 5040 34375 5046 34392
rect 5152 34375 5158 34392
rect 5040 34306 5046 34323
rect 5152 34306 5158 34323
rect 5040 34236 5046 34254
rect 5152 34236 5158 34254
rect 5040 34166 5046 34184
rect 5152 34166 5158 34184
rect 5040 33380 5046 34114
rect 5152 33380 5158 34114
rect 5040 33368 5158 33380
rect 5317 34714 5435 34726
rect 5317 34680 5323 34714
rect 5357 34680 5395 34714
rect 5429 34680 5435 34714
rect 5317 34641 5435 34680
rect 5317 34607 5323 34641
rect 5357 34607 5395 34641
rect 5429 34607 5435 34641
rect 5317 34568 5435 34607
rect 5317 34534 5323 34568
rect 5357 34534 5395 34568
rect 5429 34534 5435 34568
rect 5317 34495 5435 34534
rect 5317 34461 5323 34495
rect 5357 34461 5395 34495
rect 5429 34461 5435 34495
rect 5317 34422 5435 34461
rect 5317 33982 5323 34422
rect 5429 33982 5435 34422
rect 5317 33913 5323 33930
rect 5429 33913 5435 33930
rect 5317 33844 5323 33861
rect 5429 33844 5435 33861
rect 5317 33775 5323 33792
rect 5429 33775 5435 33792
rect 5317 33706 5323 33723
rect 5429 33706 5435 33723
rect 5317 33636 5323 33654
rect 5429 33636 5435 33654
rect 5317 33566 5323 33584
rect 5429 33566 5435 33584
rect 5317 33496 5323 33514
rect 5429 33496 5435 33514
rect 5317 33426 5323 33444
rect 5429 33426 5435 33444
rect 5369 33374 5383 33380
rect 5317 33368 5435 33374
rect 5594 34720 5712 34726
rect 5646 34668 5660 34720
rect 5594 34651 5712 34668
rect 5646 34599 5660 34651
rect 5594 34582 5712 34599
rect 5646 34530 5660 34582
rect 5594 34513 5712 34530
rect 5646 34461 5660 34513
rect 5594 34444 5712 34461
rect 5646 34422 5660 34444
rect 5594 34375 5600 34392
rect 5706 34375 5712 34392
rect 5594 34306 5600 34323
rect 5706 34306 5712 34323
rect 5594 34236 5600 34254
rect 5706 34236 5712 34254
rect 5594 34166 5600 34184
rect 5706 34166 5712 34184
rect 5594 33380 5600 34114
rect 5706 33380 5712 34114
rect 5594 33368 5712 33380
rect 5871 34714 5989 34726
rect 5871 34680 5877 34714
rect 5911 34680 5949 34714
rect 5983 34680 5989 34714
rect 5871 34641 5989 34680
rect 5871 34607 5877 34641
rect 5911 34607 5949 34641
rect 5983 34607 5989 34641
rect 5871 34568 5989 34607
rect 5871 34534 5877 34568
rect 5911 34534 5949 34568
rect 5983 34534 5989 34568
rect 5871 34495 5989 34534
rect 5871 34461 5877 34495
rect 5911 34461 5949 34495
rect 5983 34461 5989 34495
rect 5871 34422 5989 34461
rect 5871 33982 5877 34422
rect 5983 33982 5989 34422
rect 5871 33913 5877 33930
rect 5983 33913 5989 33930
rect 5871 33844 5877 33861
rect 5983 33844 5989 33861
rect 5871 33775 5877 33792
rect 5983 33775 5989 33792
rect 5871 33706 5877 33723
rect 5983 33706 5989 33723
rect 5871 33636 5877 33654
rect 5983 33636 5989 33654
rect 5871 33566 5877 33584
rect 5983 33566 5989 33584
rect 5871 33496 5877 33514
rect 5983 33496 5989 33514
rect 5871 33426 5877 33444
rect 5983 33426 5989 33444
rect 5923 33374 5937 33380
rect 5871 33368 5989 33374
rect 6148 34720 6266 34726
rect 6200 34668 6214 34720
rect 6148 34651 6266 34668
rect 6200 34599 6214 34651
rect 6148 34582 6266 34599
rect 6200 34530 6214 34582
rect 6148 34513 6266 34530
rect 6200 34461 6214 34513
rect 6148 34444 6266 34461
rect 6200 34422 6214 34444
rect 6148 34375 6154 34392
rect 6260 34375 6266 34392
rect 6148 34306 6154 34323
rect 6260 34306 6266 34323
rect 6148 34236 6154 34254
rect 6260 34236 6266 34254
rect 6148 34166 6154 34184
rect 6260 34166 6266 34184
rect 6148 33380 6154 34114
rect 6260 33380 6266 34114
rect 6148 33368 6266 33380
rect 6425 34714 6543 34726
rect 6425 34680 6431 34714
rect 6465 34680 6503 34714
rect 6537 34680 6543 34714
rect 6425 34641 6543 34680
rect 6425 34607 6431 34641
rect 6465 34607 6503 34641
rect 6537 34607 6543 34641
rect 6425 34568 6543 34607
rect 6425 34534 6431 34568
rect 6465 34534 6503 34568
rect 6537 34534 6543 34568
rect 6425 34495 6543 34534
rect 6425 34461 6431 34495
rect 6465 34461 6503 34495
rect 6537 34461 6543 34495
rect 6425 34422 6543 34461
rect 6425 33982 6431 34422
rect 6537 33982 6543 34422
rect 6425 33913 6431 33930
rect 6537 33913 6543 33930
rect 6425 33844 6431 33861
rect 6537 33844 6543 33861
rect 6425 33775 6431 33792
rect 6537 33775 6543 33792
rect 6425 33706 6431 33723
rect 6537 33706 6543 33723
rect 6425 33636 6431 33654
rect 6537 33636 6543 33654
rect 6425 33566 6431 33584
rect 6537 33566 6543 33584
rect 6425 33496 6431 33514
rect 6537 33496 6543 33514
rect 6425 33426 6431 33444
rect 6537 33426 6543 33444
rect 6477 33374 6491 33380
rect 6425 33368 6543 33374
rect 6702 34720 6820 34726
rect 6754 34668 6768 34720
rect 6702 34651 6820 34668
rect 6754 34599 6768 34651
rect 6702 34582 6820 34599
rect 6754 34530 6768 34582
rect 6702 34513 6820 34530
rect 6754 34461 6768 34513
rect 6702 34444 6820 34461
rect 6754 34422 6768 34444
rect 6702 34375 6708 34392
rect 6814 34375 6820 34392
rect 6702 34306 6708 34323
rect 6814 34306 6820 34323
rect 6702 34236 6708 34254
rect 6814 34236 6820 34254
rect 6702 34166 6708 34184
rect 6814 34166 6820 34184
rect 6702 33380 6708 34114
rect 6814 33380 6820 34114
rect 6702 33368 6820 33380
rect 6979 34714 7097 34726
rect 6979 34680 6985 34714
rect 7019 34680 7057 34714
rect 7091 34680 7097 34714
rect 6979 34641 7097 34680
rect 6979 34607 6985 34641
rect 7019 34607 7057 34641
rect 7091 34607 7097 34641
rect 6979 34568 7097 34607
rect 6979 34534 6985 34568
rect 7019 34534 7057 34568
rect 7091 34534 7097 34568
rect 6979 34495 7097 34534
rect 6979 34461 6985 34495
rect 7019 34461 7057 34495
rect 7091 34461 7097 34495
rect 6979 34422 7097 34461
rect 6979 33982 6985 34422
rect 7091 33982 7097 34422
rect 6979 33913 6985 33930
rect 7091 33913 7097 33930
rect 6979 33844 6985 33861
rect 7091 33844 7097 33861
rect 6979 33775 6985 33792
rect 7091 33775 7097 33792
rect 6979 33706 6985 33723
rect 7091 33706 7097 33723
rect 6979 33636 6985 33654
rect 7091 33636 7097 33654
rect 6979 33566 6985 33584
rect 7091 33566 7097 33584
rect 6979 33496 6985 33514
rect 7091 33496 7097 33514
rect 6979 33426 6985 33444
rect 7091 33426 7097 33444
rect 7031 33374 7045 33380
rect 6979 33368 7097 33374
rect 7256 34720 7374 34726
rect 7308 34668 7322 34720
rect 7256 34651 7374 34668
rect 7308 34599 7322 34651
rect 7256 34582 7374 34599
rect 7308 34530 7322 34582
rect 7256 34513 7374 34530
rect 7308 34461 7322 34513
rect 7256 34444 7374 34461
rect 7308 34422 7322 34444
rect 7256 34375 7262 34392
rect 7368 34375 7374 34392
rect 7256 34306 7262 34323
rect 7368 34306 7374 34323
rect 7256 34236 7262 34254
rect 7368 34236 7374 34254
rect 7256 34166 7262 34184
rect 7368 34166 7374 34184
rect 7256 33380 7262 34114
rect 7368 33380 7374 34114
rect 7256 33368 7374 33380
rect 7533 34714 7651 34726
rect 7533 34680 7539 34714
rect 7573 34680 7611 34714
rect 7645 34680 7651 34714
rect 7533 34641 7651 34680
rect 7533 34607 7539 34641
rect 7573 34607 7611 34641
rect 7645 34607 7651 34641
rect 7533 34568 7651 34607
rect 7533 34534 7539 34568
rect 7573 34534 7611 34568
rect 7645 34534 7651 34568
rect 7533 34495 7651 34534
rect 7533 34461 7539 34495
rect 7573 34461 7611 34495
rect 7645 34461 7651 34495
rect 7533 34422 7651 34461
rect 7533 33982 7539 34422
rect 7645 33982 7651 34422
rect 7533 33913 7539 33930
rect 7645 33913 7651 33930
rect 7533 33844 7539 33861
rect 7645 33844 7651 33861
rect 7533 33775 7539 33792
rect 7645 33775 7651 33792
rect 7533 33706 7539 33723
rect 7645 33706 7651 33723
rect 7533 33636 7539 33654
rect 7645 33636 7651 33654
rect 7533 33566 7539 33584
rect 7645 33566 7651 33584
rect 7533 33496 7539 33514
rect 7645 33496 7651 33514
rect 7533 33426 7539 33444
rect 7645 33426 7651 33444
rect 7585 33374 7599 33380
rect 7533 33368 7651 33374
rect 7810 34720 7928 34726
rect 7862 34668 7876 34720
rect 7810 34651 7928 34668
rect 7862 34599 7876 34651
rect 7810 34582 7928 34599
rect 7862 34530 7876 34582
rect 7810 34513 7928 34530
rect 7862 34461 7876 34513
rect 7810 34444 7928 34461
rect 7862 34422 7876 34444
rect 7810 34375 7816 34392
rect 7922 34375 7928 34392
rect 7810 34306 7816 34323
rect 7922 34306 7928 34323
rect 7810 34236 7816 34254
rect 7922 34236 7928 34254
rect 7810 34166 7816 34184
rect 7922 34166 7928 34184
rect 7810 33380 7816 34114
rect 7922 33380 7928 34114
rect 7810 33368 7928 33380
rect 8044 34725 8050 34759
rect 8084 34749 8224 34759
rect 8084 34725 8184 34749
rect 8044 34724 8184 34725
rect 8218 34724 8224 34749
rect 8044 34672 8047 34724
rect 8099 34672 8169 34724
rect 8221 34672 8224 34724
rect 8044 34655 8050 34672
rect 8084 34655 8184 34672
rect 8218 34655 8224 34672
rect 8044 34603 8047 34655
rect 8099 34603 8169 34655
rect 8221 34603 8224 34655
rect 8044 34586 8050 34603
rect 8084 34586 8184 34603
rect 8218 34586 8224 34603
rect 8044 34534 8047 34586
rect 8099 34534 8169 34586
rect 8221 34534 8224 34586
rect 8044 34517 8050 34534
rect 8084 34533 8224 34534
rect 8084 34517 8184 34533
rect 8218 34517 8224 34533
rect 8044 34465 8047 34517
rect 8099 34465 8169 34517
rect 8221 34465 8224 34517
rect 8044 34448 8050 34465
rect 8084 34461 8224 34465
rect 8084 34448 8184 34461
rect 8218 34448 8224 34461
rect 8044 34396 8047 34448
rect 8099 34396 8169 34448
rect 8221 34396 8224 34448
rect 8044 34378 8050 34396
rect 8084 34389 8224 34396
rect 8084 34378 8184 34389
rect 8218 34378 8224 34389
rect 8044 34326 8047 34378
rect 8099 34326 8169 34378
rect 8221 34326 8224 34378
rect 8044 34308 8050 34326
rect 8084 34317 8224 34326
rect 8084 34308 8184 34317
rect 8218 34308 8224 34317
rect 8044 34256 8047 34308
rect 8099 34256 8169 34308
rect 8221 34256 8224 34308
rect 8044 34255 8224 34256
rect 8044 34238 8050 34255
rect 8084 34245 8224 34255
rect 8084 34238 8184 34245
rect 8218 34238 8224 34245
rect 8044 34186 8047 34238
rect 8099 34186 8169 34238
rect 8221 34186 8224 34238
rect 8044 34183 8224 34186
rect 8044 34168 8050 34183
rect 8084 34173 8224 34183
rect 8084 34168 8184 34173
rect 8218 34168 8224 34173
rect 8044 34116 8047 34168
rect 8099 34116 8169 34168
rect 8221 34116 8224 34168
rect 8044 34111 8224 34116
rect 8044 34077 8050 34111
rect 8084 34101 8224 34111
rect 8084 34077 8184 34101
rect 8044 34067 8184 34077
rect 8218 34067 8224 34101
rect 8044 34039 8224 34067
rect 8044 34005 8050 34039
rect 8084 34029 8224 34039
rect 8084 34005 8184 34029
rect 8044 33995 8184 34005
rect 8218 33995 8224 34029
rect 8044 33967 8224 33995
rect 8044 33933 8050 33967
rect 8084 33957 8224 33967
rect 8084 33933 8184 33957
rect 8044 33923 8184 33933
rect 8218 33923 8224 33957
rect 8044 33895 8224 33923
rect 8044 33861 8050 33895
rect 8084 33885 8224 33895
rect 8084 33861 8184 33885
rect 8044 33851 8184 33861
rect 8218 33851 8224 33885
rect 8044 33823 8224 33851
rect 8044 33789 8050 33823
rect 8084 33813 8224 33823
rect 8084 33789 8184 33813
rect 8044 33779 8184 33789
rect 8218 33779 8224 33813
rect 8044 33751 8224 33779
rect 8044 33717 8050 33751
rect 8084 33741 8224 33751
rect 8084 33717 8184 33741
rect 8044 33707 8184 33717
rect 8218 33707 8224 33741
rect 8044 33679 8224 33707
rect 8044 33645 8050 33679
rect 8084 33669 8224 33679
rect 8084 33645 8184 33669
rect 8044 33635 8184 33645
rect 8218 33635 8224 33669
rect 8044 33607 8224 33635
rect 8044 33573 8050 33607
rect 8084 33597 8224 33607
rect 8084 33573 8184 33597
rect 8044 33563 8184 33573
rect 8218 33563 8224 33597
rect 8044 33535 8224 33563
rect 8044 33501 8050 33535
rect 8084 33525 8224 33535
rect 8084 33501 8184 33525
rect 8044 33491 8184 33501
rect 8218 33491 8224 33525
rect 8044 33463 8224 33491
rect 8044 33429 8050 33463
rect 8084 33453 8224 33463
rect 8084 33429 8184 33453
rect 8044 33419 8184 33429
rect 8218 33419 8224 33453
rect 8044 33391 8224 33419
rect 8044 33357 8050 33391
rect 8084 33381 8224 33391
rect 8084 33357 8184 33381
rect 8044 33347 8184 33357
rect 8218 33347 8224 33381
rect 8044 33319 8224 33347
rect 8044 33285 8050 33319
rect 8084 33309 8224 33319
rect 8084 33285 8184 33309
rect 8044 33275 8184 33285
rect 8218 33275 8224 33309
rect 8044 33247 8224 33275
rect 8044 33213 8050 33247
rect 8084 33237 8224 33247
rect 8084 33213 8184 33237
rect 8044 33203 8184 33213
rect 8218 33203 8224 33237
rect 8044 33175 8224 33203
tri 2712 33141 2736 33165 sw
rect 8044 33141 8050 33175
rect 8084 33165 8224 33175
rect 8084 33141 8184 33165
rect 2543 33133 2736 33141
tri 2736 33133 2744 33141 sw
rect 2543 33100 7750 33133
rect 2543 33066 3035 33100
rect 3069 33066 3108 33100
rect 3142 33066 3181 33100
rect 3215 33066 3254 33100
rect 3288 33066 3327 33100
rect 3361 33066 3400 33100
rect 3434 33066 3473 33100
rect 3507 33066 3546 33100
rect 3580 33066 3619 33100
rect 3653 33066 3692 33100
rect 3726 33066 3765 33100
rect 3799 33066 3838 33100
rect 3872 33066 3911 33100
rect 3945 33066 3984 33100
rect 4018 33066 4057 33100
rect 4091 33066 4130 33100
rect 4164 33066 4203 33100
rect 4237 33066 4276 33100
rect 4310 33066 4349 33100
rect 4383 33066 4422 33100
rect 4456 33066 4495 33100
rect 4529 33066 4568 33100
rect 4602 33066 4641 33100
rect 4675 33066 4714 33100
rect 4748 33066 4787 33100
rect 4821 33066 4860 33100
rect 4894 33066 4933 33100
rect 4967 33066 5006 33100
rect 5040 33066 5079 33100
rect 5113 33066 5152 33100
rect 5186 33066 5225 33100
rect 5259 33066 5298 33100
rect 5332 33066 5371 33100
rect 5405 33066 5444 33100
rect 5478 33066 5517 33100
rect 5551 33066 5590 33100
rect 5624 33066 5663 33100
rect 5697 33066 5736 33100
rect 5770 33066 5809 33100
rect 5843 33066 5882 33100
rect 5916 33066 5955 33100
rect 5989 33066 6027 33100
rect 6061 33066 6099 33100
rect 6133 33066 6171 33100
rect 6205 33066 6243 33100
rect 6277 33066 6315 33100
rect 6349 33066 6387 33100
rect 6421 33066 6459 33100
rect 6493 33066 6531 33100
rect 6565 33066 6603 33100
rect 6637 33066 6675 33100
rect 6709 33066 6747 33100
rect 6781 33066 6819 33100
rect 6853 33066 6891 33100
rect 6925 33066 6963 33100
rect 6997 33066 7035 33100
rect 7069 33066 7107 33100
rect 7141 33066 7179 33100
rect 7213 33066 7251 33100
rect 7285 33066 7323 33100
rect 7357 33066 7395 33100
rect 7429 33066 7467 33100
rect 7501 33066 7539 33100
rect 7573 33066 7611 33100
rect 7645 33066 7683 33100
rect 7717 33066 7750 33100
rect 2543 33046 7750 33066
rect 8044 33131 8184 33141
rect 8218 33131 8224 33165
rect 8044 33103 8224 33131
rect 8044 33069 8050 33103
rect 8084 33093 8224 33103
rect 8084 33069 8184 33093
rect 8044 33059 8184 33069
rect 8218 33059 8224 33093
rect 2543 33031 2740 33046
tri 2740 33031 2755 33046 nw
rect 8044 33031 8224 33059
rect 2543 31187 2712 33031
tri 2712 33003 2740 33031 nw
rect 8044 32997 8050 33031
rect 8084 33021 8224 33031
rect 8084 32997 8184 33021
rect 8044 32987 8184 32997
rect 8218 32987 8224 33021
rect 8044 32959 8224 32987
rect 8044 32925 8050 32959
rect 8084 32949 8224 32959
rect 8084 32925 8184 32949
rect 8044 32915 8184 32925
rect 8218 32915 8224 32949
rect 8044 32887 8224 32915
rect 8044 32853 8050 32887
rect 8084 32877 8224 32887
rect 8084 32853 8184 32877
rect 8044 32843 8184 32853
rect 8218 32843 8224 32877
rect 8044 32815 8224 32843
rect 8044 32781 8050 32815
rect 8084 32805 8224 32815
rect 8084 32781 8184 32805
rect 8044 32771 8184 32781
rect 8218 32771 8224 32805
rect 8044 32743 8224 32771
rect 2824 32720 2942 32726
rect 2876 32668 2890 32720
rect 2824 32651 2942 32668
rect 2876 32599 2890 32651
rect 2824 32582 2942 32599
rect 2876 32530 2890 32582
rect 2824 32513 2942 32530
rect 2876 32461 2890 32513
rect 2824 32444 2942 32461
rect 2876 32422 2890 32444
rect 2824 32375 2830 32392
rect 2936 32375 2942 32392
rect 2824 32306 2830 32323
rect 2936 32306 2942 32323
rect 2824 32236 2830 32254
rect 2936 32236 2942 32254
rect 2824 32166 2830 32184
rect 2936 32166 2942 32184
rect 2824 31380 2830 32114
rect 2936 31380 2942 32114
rect 2824 31368 2942 31380
rect 3101 32714 3219 32726
rect 3101 32680 3107 32714
rect 3141 32680 3179 32714
rect 3213 32680 3219 32714
rect 3101 32641 3219 32680
rect 3101 32607 3107 32641
rect 3141 32607 3179 32641
rect 3213 32607 3219 32641
rect 3101 32568 3219 32607
rect 3101 32534 3107 32568
rect 3141 32534 3179 32568
rect 3213 32534 3219 32568
rect 3101 32495 3219 32534
rect 3101 32461 3107 32495
rect 3141 32461 3179 32495
rect 3213 32461 3219 32495
rect 3101 32422 3219 32461
rect 3101 31982 3107 32422
rect 3213 31982 3219 32422
rect 3101 31913 3107 31930
rect 3213 31913 3219 31930
rect 3101 31844 3107 31861
rect 3213 31844 3219 31861
rect 3101 31775 3107 31792
rect 3213 31775 3219 31792
rect 3101 31706 3107 31723
rect 3213 31706 3219 31723
rect 3101 31636 3107 31654
rect 3213 31636 3219 31654
rect 3101 31566 3107 31584
rect 3213 31566 3219 31584
rect 3101 31496 3107 31514
rect 3213 31496 3219 31514
rect 3101 31426 3107 31444
rect 3213 31426 3219 31444
rect 3153 31374 3167 31380
rect 3101 31368 3219 31374
rect 3378 32720 3496 32726
rect 3430 32668 3444 32720
rect 3378 32651 3496 32668
rect 3430 32599 3444 32651
rect 3378 32582 3496 32599
rect 3430 32530 3444 32582
rect 3378 32513 3496 32530
rect 3430 32461 3444 32513
rect 3378 32444 3496 32461
rect 3430 32422 3444 32444
rect 3378 32375 3384 32392
rect 3490 32375 3496 32392
rect 3378 32306 3384 32323
rect 3490 32306 3496 32323
rect 3378 32236 3384 32254
rect 3490 32236 3496 32254
rect 3378 32166 3384 32184
rect 3490 32166 3496 32184
rect 3378 31380 3384 32114
rect 3490 31380 3496 32114
rect 3378 31368 3496 31380
rect 3655 32714 3773 32726
rect 3655 32680 3661 32714
rect 3695 32680 3733 32714
rect 3767 32680 3773 32714
rect 3655 32641 3773 32680
rect 3655 32607 3661 32641
rect 3695 32607 3733 32641
rect 3767 32607 3773 32641
rect 3655 32568 3773 32607
rect 3655 32534 3661 32568
rect 3695 32534 3733 32568
rect 3767 32534 3773 32568
rect 3655 32495 3773 32534
rect 3655 32461 3661 32495
rect 3695 32461 3733 32495
rect 3767 32461 3773 32495
rect 3655 32422 3773 32461
rect 3655 31982 3661 32422
rect 3767 31982 3773 32422
rect 3655 31913 3661 31930
rect 3767 31913 3773 31930
rect 3655 31844 3661 31861
rect 3767 31844 3773 31861
rect 3655 31775 3661 31792
rect 3767 31775 3773 31792
rect 3655 31706 3661 31723
rect 3767 31706 3773 31723
rect 3655 31636 3661 31654
rect 3767 31636 3773 31654
rect 3655 31566 3661 31584
rect 3767 31566 3773 31584
rect 3655 31496 3661 31514
rect 3767 31496 3773 31514
rect 3655 31426 3661 31444
rect 3767 31426 3773 31444
rect 3707 31374 3721 31380
rect 3655 31368 3773 31374
rect 3932 32720 4050 32726
rect 3984 32668 3998 32720
rect 3932 32651 4050 32668
rect 3984 32599 3998 32651
rect 3932 32582 4050 32599
rect 3984 32530 3998 32582
rect 3932 32513 4050 32530
rect 3984 32461 3998 32513
rect 3932 32444 4050 32461
rect 3984 32422 3998 32444
rect 3932 32375 3938 32392
rect 4044 32375 4050 32392
rect 3932 32306 3938 32323
rect 4044 32306 4050 32323
rect 3932 32236 3938 32254
rect 4044 32236 4050 32254
rect 3932 32166 3938 32184
rect 4044 32166 4050 32184
rect 3932 31380 3938 32114
rect 4044 31380 4050 32114
rect 3932 31368 4050 31380
rect 4209 32714 4327 32726
rect 4209 32680 4215 32714
rect 4249 32680 4287 32714
rect 4321 32680 4327 32714
rect 4209 32641 4327 32680
rect 4209 32607 4215 32641
rect 4249 32607 4287 32641
rect 4321 32607 4327 32641
rect 4209 32568 4327 32607
rect 4209 32534 4215 32568
rect 4249 32534 4287 32568
rect 4321 32534 4327 32568
rect 4209 32495 4327 32534
rect 4209 32461 4215 32495
rect 4249 32461 4287 32495
rect 4321 32461 4327 32495
rect 4209 32422 4327 32461
rect 4209 31982 4215 32422
rect 4321 31982 4327 32422
rect 4209 31913 4215 31930
rect 4321 31913 4327 31930
rect 4209 31844 4215 31861
rect 4321 31844 4327 31861
rect 4209 31775 4215 31792
rect 4321 31775 4327 31792
rect 4209 31706 4215 31723
rect 4321 31706 4327 31723
rect 4209 31636 4215 31654
rect 4321 31636 4327 31654
rect 4209 31566 4215 31584
rect 4321 31566 4327 31584
rect 4209 31496 4215 31514
rect 4321 31496 4327 31514
rect 4209 31426 4215 31444
rect 4321 31426 4327 31444
rect 4261 31374 4275 31380
rect 4209 31368 4327 31374
rect 4486 32720 4604 32726
rect 4538 32668 4552 32720
rect 4486 32651 4604 32668
rect 4538 32599 4552 32651
rect 4486 32582 4604 32599
rect 4538 32530 4552 32582
rect 4486 32513 4604 32530
rect 4538 32461 4552 32513
rect 4486 32444 4604 32461
rect 4538 32422 4552 32444
rect 4486 32375 4492 32392
rect 4598 32375 4604 32392
rect 4486 32306 4492 32323
rect 4598 32306 4604 32323
rect 4486 32236 4492 32254
rect 4598 32236 4604 32254
rect 4486 32166 4492 32184
rect 4598 32166 4604 32184
rect 4486 31380 4492 32114
rect 4598 31380 4604 32114
rect 4486 31368 4604 31380
rect 4763 32714 4881 32726
rect 4763 32680 4769 32714
rect 4803 32680 4841 32714
rect 4875 32680 4881 32714
rect 4763 32641 4881 32680
rect 4763 32607 4769 32641
rect 4803 32607 4841 32641
rect 4875 32607 4881 32641
rect 4763 32568 4881 32607
rect 4763 32534 4769 32568
rect 4803 32534 4841 32568
rect 4875 32534 4881 32568
rect 4763 32495 4881 32534
rect 4763 32461 4769 32495
rect 4803 32461 4841 32495
rect 4875 32461 4881 32495
rect 4763 32422 4881 32461
rect 4763 31982 4769 32422
rect 4875 31982 4881 32422
rect 4763 31913 4769 31930
rect 4875 31913 4881 31930
rect 4763 31844 4769 31861
rect 4875 31844 4881 31861
rect 4763 31775 4769 31792
rect 4875 31775 4881 31792
rect 4763 31706 4769 31723
rect 4875 31706 4881 31723
rect 4763 31636 4769 31654
rect 4875 31636 4881 31654
rect 4763 31566 4769 31584
rect 4875 31566 4881 31584
rect 4763 31496 4769 31514
rect 4875 31496 4881 31514
rect 4763 31426 4769 31444
rect 4875 31426 4881 31444
rect 4815 31374 4829 31380
rect 4763 31368 4881 31374
rect 5040 32720 5158 32726
rect 5092 32668 5106 32720
rect 5040 32651 5158 32668
rect 5092 32599 5106 32651
rect 5040 32582 5158 32599
rect 5092 32530 5106 32582
rect 5040 32513 5158 32530
rect 5092 32461 5106 32513
rect 5040 32444 5158 32461
rect 5092 32422 5106 32444
rect 5040 32375 5046 32392
rect 5152 32375 5158 32392
rect 5040 32306 5046 32323
rect 5152 32306 5158 32323
rect 5040 32236 5046 32254
rect 5152 32236 5158 32254
rect 5040 32166 5046 32184
rect 5152 32166 5158 32184
rect 5040 31380 5046 32114
rect 5152 31380 5158 32114
rect 5040 31368 5158 31380
rect 5317 32714 5435 32726
rect 5317 32680 5323 32714
rect 5357 32680 5395 32714
rect 5429 32680 5435 32714
rect 5317 32641 5435 32680
rect 5317 32607 5323 32641
rect 5357 32607 5395 32641
rect 5429 32607 5435 32641
rect 5317 32568 5435 32607
rect 5317 32534 5323 32568
rect 5357 32534 5395 32568
rect 5429 32534 5435 32568
rect 5317 32495 5435 32534
rect 5317 32461 5323 32495
rect 5357 32461 5395 32495
rect 5429 32461 5435 32495
rect 5317 32422 5435 32461
rect 5317 31982 5323 32422
rect 5429 31982 5435 32422
rect 5317 31913 5323 31930
rect 5429 31913 5435 31930
rect 5317 31844 5323 31861
rect 5429 31844 5435 31861
rect 5317 31775 5323 31792
rect 5429 31775 5435 31792
rect 5317 31706 5323 31723
rect 5429 31706 5435 31723
rect 5317 31636 5323 31654
rect 5429 31636 5435 31654
rect 5317 31566 5323 31584
rect 5429 31566 5435 31584
rect 5317 31496 5323 31514
rect 5429 31496 5435 31514
rect 5317 31426 5323 31444
rect 5429 31426 5435 31444
rect 5369 31374 5383 31380
rect 5317 31368 5435 31374
rect 5594 32720 5712 32726
rect 5646 32668 5660 32720
rect 5594 32651 5712 32668
rect 5646 32599 5660 32651
rect 5594 32582 5712 32599
rect 5646 32530 5660 32582
rect 5594 32513 5712 32530
rect 5646 32461 5660 32513
rect 5594 32444 5712 32461
rect 5646 32422 5660 32444
rect 5594 32375 5600 32392
rect 5706 32375 5712 32392
rect 5594 32306 5600 32323
rect 5706 32306 5712 32323
rect 5594 32236 5600 32254
rect 5706 32236 5712 32254
rect 5594 32166 5600 32184
rect 5706 32166 5712 32184
rect 5594 31380 5600 32114
rect 5706 31380 5712 32114
rect 5594 31368 5712 31380
rect 5871 32714 5989 32726
rect 5871 32680 5877 32714
rect 5911 32680 5949 32714
rect 5983 32680 5989 32714
rect 5871 32641 5989 32680
rect 5871 32607 5877 32641
rect 5911 32607 5949 32641
rect 5983 32607 5989 32641
rect 5871 32568 5989 32607
rect 5871 32534 5877 32568
rect 5911 32534 5949 32568
rect 5983 32534 5989 32568
rect 5871 32495 5989 32534
rect 5871 32461 5877 32495
rect 5911 32461 5949 32495
rect 5983 32461 5989 32495
rect 5871 32422 5989 32461
rect 5871 31982 5877 32422
rect 5983 31982 5989 32422
rect 5871 31913 5877 31930
rect 5983 31913 5989 31930
rect 5871 31844 5877 31861
rect 5983 31844 5989 31861
rect 5871 31775 5877 31792
rect 5983 31775 5989 31792
rect 5871 31706 5877 31723
rect 5983 31706 5989 31723
rect 5871 31636 5877 31654
rect 5983 31636 5989 31654
rect 5871 31566 5877 31584
rect 5983 31566 5989 31584
rect 5871 31496 5877 31514
rect 5983 31496 5989 31514
rect 5871 31426 5877 31444
rect 5983 31426 5989 31444
rect 5923 31374 5937 31380
rect 5871 31368 5989 31374
rect 6148 32720 6266 32726
rect 6200 32668 6214 32720
rect 6148 32651 6266 32668
rect 6200 32599 6214 32651
rect 6148 32582 6266 32599
rect 6200 32530 6214 32582
rect 6148 32513 6266 32530
rect 6200 32461 6214 32513
rect 6148 32444 6266 32461
rect 6200 32422 6214 32444
rect 6148 32375 6154 32392
rect 6260 32375 6266 32392
rect 6148 32306 6154 32323
rect 6260 32306 6266 32323
rect 6148 32236 6154 32254
rect 6260 32236 6266 32254
rect 6148 32166 6154 32184
rect 6260 32166 6266 32184
rect 6148 31380 6154 32114
rect 6260 31380 6266 32114
rect 6148 31368 6266 31380
rect 6425 32714 6543 32726
rect 6425 32680 6431 32714
rect 6465 32680 6503 32714
rect 6537 32680 6543 32714
rect 6425 32641 6543 32680
rect 6425 32607 6431 32641
rect 6465 32607 6503 32641
rect 6537 32607 6543 32641
rect 6425 32568 6543 32607
rect 6425 32534 6431 32568
rect 6465 32534 6503 32568
rect 6537 32534 6543 32568
rect 6425 32495 6543 32534
rect 6425 32461 6431 32495
rect 6465 32461 6503 32495
rect 6537 32461 6543 32495
rect 6425 32422 6543 32461
rect 6425 31982 6431 32422
rect 6537 31982 6543 32422
rect 6425 31913 6431 31930
rect 6537 31913 6543 31930
rect 6425 31844 6431 31861
rect 6537 31844 6543 31861
rect 6425 31775 6431 31792
rect 6537 31775 6543 31792
rect 6425 31706 6431 31723
rect 6537 31706 6543 31723
rect 6425 31636 6431 31654
rect 6537 31636 6543 31654
rect 6425 31566 6431 31584
rect 6537 31566 6543 31584
rect 6425 31496 6431 31514
rect 6537 31496 6543 31514
rect 6425 31426 6431 31444
rect 6537 31426 6543 31444
rect 6477 31374 6491 31380
rect 6425 31368 6543 31374
rect 6702 32720 6820 32726
rect 6754 32668 6768 32720
rect 6702 32651 6820 32668
rect 6754 32599 6768 32651
rect 6702 32582 6820 32599
rect 6754 32530 6768 32582
rect 6702 32513 6820 32530
rect 6754 32461 6768 32513
rect 6702 32444 6820 32461
rect 6754 32422 6768 32444
rect 6702 32375 6708 32392
rect 6814 32375 6820 32392
rect 6702 32306 6708 32323
rect 6814 32306 6820 32323
rect 6702 32236 6708 32254
rect 6814 32236 6820 32254
rect 6702 32166 6708 32184
rect 6814 32166 6820 32184
rect 6702 31380 6708 32114
rect 6814 31380 6820 32114
rect 6702 31368 6820 31380
rect 6979 32714 7097 32726
rect 6979 32680 6985 32714
rect 7019 32680 7057 32714
rect 7091 32680 7097 32714
rect 6979 32641 7097 32680
rect 6979 32607 6985 32641
rect 7019 32607 7057 32641
rect 7091 32607 7097 32641
rect 6979 32568 7097 32607
rect 6979 32534 6985 32568
rect 7019 32534 7057 32568
rect 7091 32534 7097 32568
rect 6979 32495 7097 32534
rect 6979 32461 6985 32495
rect 7019 32461 7057 32495
rect 7091 32461 7097 32495
rect 6979 32422 7097 32461
rect 6979 31982 6985 32422
rect 7091 31982 7097 32422
rect 6979 31913 6985 31930
rect 7091 31913 7097 31930
rect 6979 31844 6985 31861
rect 7091 31844 7097 31861
rect 6979 31775 6985 31792
rect 7091 31775 7097 31792
rect 6979 31706 6985 31723
rect 7091 31706 7097 31723
rect 6979 31636 6985 31654
rect 7091 31636 7097 31654
rect 6979 31566 6985 31584
rect 7091 31566 7097 31584
rect 6979 31496 6985 31514
rect 7091 31496 7097 31514
rect 6979 31426 6985 31444
rect 7091 31426 7097 31444
rect 7031 31374 7045 31380
rect 6979 31368 7097 31374
rect 7256 32720 7374 32726
rect 7308 32668 7322 32720
rect 7256 32651 7374 32668
rect 7308 32599 7322 32651
rect 7256 32582 7374 32599
rect 7308 32530 7322 32582
rect 7256 32513 7374 32530
rect 7308 32461 7322 32513
rect 7256 32444 7374 32461
rect 7308 32422 7322 32444
rect 7256 32375 7262 32392
rect 7368 32375 7374 32392
rect 7256 32306 7262 32323
rect 7368 32306 7374 32323
rect 7256 32236 7262 32254
rect 7368 32236 7374 32254
rect 7256 32166 7262 32184
rect 7368 32166 7374 32184
rect 7256 31380 7262 32114
rect 7368 31380 7374 32114
rect 7256 31368 7374 31380
rect 7533 32714 7651 32726
rect 7533 32680 7539 32714
rect 7573 32680 7611 32714
rect 7645 32680 7651 32714
rect 7533 32641 7651 32680
rect 7533 32607 7539 32641
rect 7573 32607 7611 32641
rect 7645 32607 7651 32641
rect 7533 32568 7651 32607
rect 7533 32534 7539 32568
rect 7573 32534 7611 32568
rect 7645 32534 7651 32568
rect 7533 32495 7651 32534
rect 7533 32461 7539 32495
rect 7573 32461 7611 32495
rect 7645 32461 7651 32495
rect 7533 32422 7651 32461
rect 7533 31982 7539 32422
rect 7645 31982 7651 32422
rect 7533 31913 7539 31930
rect 7645 31913 7651 31930
rect 7533 31844 7539 31861
rect 7645 31844 7651 31861
rect 7533 31775 7539 31792
rect 7645 31775 7651 31792
rect 7533 31706 7539 31723
rect 7645 31706 7651 31723
rect 7533 31636 7539 31654
rect 7645 31636 7651 31654
rect 7533 31566 7539 31584
rect 7645 31566 7651 31584
rect 7533 31496 7539 31514
rect 7645 31496 7651 31514
rect 7533 31426 7539 31444
rect 7645 31426 7651 31444
rect 7585 31374 7599 31380
rect 7533 31368 7651 31374
rect 7810 32720 7928 32726
rect 7862 32668 7876 32720
rect 7810 32651 7928 32668
rect 7862 32599 7876 32651
rect 7810 32582 7928 32599
rect 7862 32530 7876 32582
rect 7810 32513 7928 32530
rect 7862 32461 7876 32513
rect 7810 32444 7928 32461
rect 7862 32422 7876 32444
rect 7810 32375 7816 32392
rect 7922 32375 7928 32392
rect 7810 32306 7816 32323
rect 7922 32306 7928 32323
rect 7810 32236 7816 32254
rect 7922 32236 7928 32254
rect 7810 32166 7816 32184
rect 7922 32166 7928 32184
rect 7810 31380 7816 32114
rect 7922 31380 7928 32114
rect 7810 31368 7928 31380
rect 8044 32724 8050 32743
rect 8084 32733 8224 32743
rect 8084 32724 8184 32733
rect 8218 32724 8224 32733
rect 8044 32672 8047 32724
rect 8099 32672 8169 32724
rect 8221 32672 8224 32724
rect 8044 32671 8224 32672
rect 8044 32655 8050 32671
rect 8084 32661 8224 32671
rect 8084 32655 8184 32661
rect 8218 32655 8224 32661
rect 8044 32603 8047 32655
rect 8099 32603 8169 32655
rect 8221 32603 8224 32655
rect 8044 32599 8224 32603
rect 8044 32586 8050 32599
rect 8084 32589 8224 32599
rect 8084 32586 8184 32589
rect 8218 32586 8224 32589
rect 8044 32534 8047 32586
rect 8099 32534 8169 32586
rect 8221 32534 8224 32586
rect 8044 32527 8224 32534
rect 8044 32517 8050 32527
rect 8084 32517 8224 32527
rect 8044 32465 8047 32517
rect 8099 32465 8169 32517
rect 8221 32465 8224 32517
rect 8044 32455 8224 32465
rect 8044 32448 8050 32455
rect 8084 32448 8224 32455
rect 8044 32396 8047 32448
rect 8099 32396 8169 32448
rect 8221 32396 8224 32448
rect 8044 32383 8224 32396
rect 8044 32378 8050 32383
rect 8084 32378 8224 32383
rect 8044 32326 8047 32378
rect 8099 32326 8169 32378
rect 8221 32326 8224 32378
rect 8044 32311 8224 32326
rect 8044 32308 8050 32311
rect 8084 32308 8224 32311
rect 8044 32256 8047 32308
rect 8099 32256 8169 32308
rect 8221 32256 8224 32308
rect 8044 32239 8224 32256
rect 8044 32238 8050 32239
rect 8084 32238 8224 32239
rect 8044 32186 8047 32238
rect 8099 32186 8169 32238
rect 8221 32186 8224 32238
rect 8044 32168 8224 32186
rect 8044 32116 8047 32168
rect 8099 32116 8169 32168
rect 8221 32116 8224 32168
rect 8044 32095 8224 32116
rect 8044 32061 8050 32095
rect 8084 32085 8224 32095
rect 8084 32061 8184 32085
rect 8044 32051 8184 32061
rect 8218 32051 8224 32085
rect 8044 32023 8224 32051
rect 8044 31989 8050 32023
rect 8084 32013 8224 32023
rect 8084 31989 8184 32013
rect 8044 31979 8184 31989
rect 8218 31979 8224 32013
rect 8044 31951 8224 31979
rect 8044 31917 8050 31951
rect 8084 31941 8224 31951
rect 8084 31917 8184 31941
rect 8044 31907 8184 31917
rect 8218 31907 8224 31941
rect 8044 31879 8224 31907
rect 8044 31845 8050 31879
rect 8084 31869 8224 31879
rect 8084 31845 8184 31869
rect 8044 31835 8184 31845
rect 8218 31835 8224 31869
rect 8044 31807 8224 31835
rect 8044 31773 8050 31807
rect 8084 31797 8224 31807
rect 8084 31773 8184 31797
rect 8044 31763 8184 31773
rect 8218 31763 8224 31797
rect 8044 31735 8224 31763
rect 8044 31701 8050 31735
rect 8084 31725 8224 31735
rect 8084 31701 8184 31725
rect 8044 31691 8184 31701
rect 8218 31691 8224 31725
rect 8044 31663 8224 31691
rect 8044 31629 8050 31663
rect 8084 31653 8224 31663
rect 8084 31629 8184 31653
rect 8044 31619 8184 31629
rect 8218 31619 8224 31653
rect 8044 31591 8224 31619
rect 8044 31557 8050 31591
rect 8084 31581 8224 31591
rect 8084 31557 8184 31581
rect 8044 31547 8184 31557
rect 8218 31547 8224 31581
rect 8044 31519 8224 31547
rect 8044 31485 8050 31519
rect 8084 31509 8224 31519
rect 8084 31485 8184 31509
rect 8044 31475 8184 31485
rect 8218 31475 8224 31509
rect 8044 31447 8224 31475
rect 8044 31413 8050 31447
rect 8084 31437 8224 31447
rect 8084 31413 8184 31437
rect 8044 31403 8184 31413
rect 8218 31403 8224 31437
rect 8044 31375 8224 31403
rect 8044 31341 8050 31375
rect 8084 31365 8224 31375
rect 8084 31341 8184 31365
rect 8044 31331 8184 31341
rect 8218 31331 8224 31365
rect 8044 31303 8224 31331
rect 8044 31269 8050 31303
rect 8084 31293 8224 31303
rect 8084 31269 8184 31293
rect 8044 31259 8184 31269
rect 8218 31259 8224 31293
rect 8044 31231 8224 31259
rect 8044 31197 8050 31231
rect 8084 31221 8224 31231
rect 8084 31197 8184 31221
tri 2712 31187 2714 31189 sw
rect 8044 31187 8184 31197
rect 8218 31187 8224 31221
rect 2543 31159 2714 31187
tri 2714 31159 2742 31187 sw
rect 8044 31159 8224 31187
rect 2543 31157 2742 31159
tri 2742 31157 2744 31159 sw
rect 2543 31077 7729 31157
rect 2543 31043 3035 31077
rect 3069 31043 3108 31077
rect 3142 31043 3181 31077
rect 3215 31043 3254 31077
rect 3288 31043 3327 31077
rect 3361 31043 3400 31077
rect 3434 31043 3473 31077
rect 3507 31043 3546 31077
rect 3580 31043 3619 31077
rect 3653 31043 3692 31077
rect 3726 31043 3765 31077
rect 3799 31043 3838 31077
rect 3872 31043 3911 31077
rect 3945 31043 3984 31077
rect 4018 31043 4057 31077
rect 4091 31043 4130 31077
rect 4164 31043 4203 31077
rect 4237 31043 4276 31077
rect 4310 31043 4349 31077
rect 4383 31043 4422 31077
rect 4456 31043 4495 31077
rect 4529 31043 4568 31077
rect 4602 31043 4641 31077
rect 4675 31043 4714 31077
rect 4748 31043 4787 31077
rect 4821 31043 4860 31077
rect 4894 31043 4933 31077
rect 4967 31043 5006 31077
rect 5040 31043 5079 31077
rect 5113 31043 5152 31077
rect 5186 31043 5225 31077
rect 5259 31043 5298 31077
rect 5332 31043 5371 31077
rect 5405 31043 5444 31077
rect 5478 31043 5517 31077
rect 5551 31043 5590 31077
rect 5624 31043 5663 31077
rect 5697 31043 5736 31077
rect 5770 31043 5809 31077
rect 5843 31043 5882 31077
rect 5916 31043 5955 31077
rect 5989 31043 6027 31077
rect 6061 31043 6099 31077
rect 6133 31043 6171 31077
rect 6205 31043 6243 31077
rect 6277 31043 6315 31077
rect 6349 31043 6387 31077
rect 6421 31043 6459 31077
rect 6493 31043 6531 31077
rect 6565 31043 6603 31077
rect 6637 31043 6675 31077
rect 6709 31043 6747 31077
rect 6781 31043 6819 31077
rect 6853 31043 6891 31077
rect 6925 31043 6963 31077
rect 6997 31043 7035 31077
rect 7069 31043 7107 31077
rect 7141 31043 7179 31077
rect 7213 31043 7251 31077
rect 7285 31043 7323 31077
rect 7357 31043 7395 31077
rect 7429 31043 7467 31077
rect 7501 31043 7539 31077
rect 7573 31043 7611 31077
rect 7645 31043 7683 31077
rect 7717 31043 7729 31077
rect 2543 31037 7729 31043
rect 8044 31125 8050 31159
rect 8084 31149 8224 31159
rect 8084 31125 8184 31149
rect 8044 31115 8184 31125
rect 8218 31115 8224 31149
rect 8044 31087 8224 31115
rect 8044 31053 8050 31087
rect 8084 31077 8224 31087
rect 8084 31053 8184 31077
rect 8044 31043 8184 31053
rect 8218 31043 8224 31077
rect 2543 31015 2740 31037
tri 2740 31015 2762 31037 nw
rect 8044 31015 8224 31043
rect 2543 29359 2712 31015
tri 2712 30987 2740 31015 nw
rect 8044 30981 8050 31015
rect 8084 31005 8224 31015
rect 8084 30981 8184 31005
rect 8044 30971 8184 30981
rect 8218 30971 8224 31005
rect 8044 30943 8224 30971
rect 8044 30909 8050 30943
rect 8084 30933 8224 30943
rect 8084 30909 8184 30933
rect 8044 30899 8184 30909
rect 8218 30899 8224 30933
rect 8044 30871 8224 30899
rect 8044 30837 8050 30871
rect 8084 30861 8224 30871
rect 8084 30837 8184 30861
rect 8044 30827 8184 30837
rect 8218 30827 8224 30861
rect 8044 30799 8224 30827
rect 8044 30765 8050 30799
rect 8084 30789 8224 30799
rect 8084 30765 8184 30789
rect 8044 30755 8184 30765
rect 8218 30755 8224 30789
rect 8044 30727 8224 30755
rect 2824 30720 2942 30726
rect 2876 30668 2890 30720
rect 2824 30651 2942 30668
rect 2876 30599 2890 30651
rect 2824 30582 2942 30599
rect 2876 30530 2890 30582
rect 2824 30513 2942 30530
rect 2876 30461 2890 30513
rect 2824 30444 2942 30461
rect 2876 30422 2890 30444
rect 2824 30375 2830 30392
rect 2936 30375 2942 30392
rect 2824 30306 2830 30323
rect 2936 30306 2942 30323
rect 2824 30236 2830 30254
rect 2936 30236 2942 30254
rect 2824 30166 2830 30184
rect 2936 30166 2942 30184
rect 2824 29380 2830 30114
rect 2936 29380 2942 30114
tri 2712 29359 2729 29376 sw
rect 2824 29368 2942 29380
rect 3101 30714 3219 30726
rect 3101 30680 3107 30714
rect 3141 30680 3179 30714
rect 3213 30680 3219 30714
rect 3101 30641 3219 30680
rect 3101 30607 3107 30641
rect 3141 30607 3179 30641
rect 3213 30607 3219 30641
rect 3101 30568 3219 30607
rect 3101 30534 3107 30568
rect 3141 30534 3179 30568
rect 3213 30534 3219 30568
rect 3101 30495 3219 30534
rect 3101 30461 3107 30495
rect 3141 30461 3179 30495
rect 3213 30461 3219 30495
rect 3101 30422 3219 30461
rect 3101 29982 3107 30422
rect 3213 29982 3219 30422
rect 3101 29913 3107 29930
rect 3213 29913 3219 29930
rect 3101 29844 3107 29861
rect 3213 29844 3219 29861
rect 3101 29775 3107 29792
rect 3213 29775 3219 29792
rect 3101 29706 3107 29723
rect 3213 29706 3219 29723
rect 3101 29636 3107 29654
rect 3213 29636 3219 29654
rect 3101 29566 3107 29584
rect 3213 29566 3219 29584
rect 3101 29496 3107 29514
rect 3213 29496 3219 29514
rect 3101 29426 3107 29444
rect 3213 29426 3219 29444
rect 3153 29374 3167 29380
rect 3101 29368 3219 29374
rect 3378 30720 3496 30726
rect 3430 30668 3444 30720
rect 3378 30651 3496 30668
rect 3430 30599 3444 30651
rect 3378 30582 3496 30599
rect 3430 30530 3444 30582
rect 3378 30513 3496 30530
rect 3430 30461 3444 30513
rect 3378 30444 3496 30461
rect 3430 30422 3444 30444
rect 3378 30375 3384 30392
rect 3490 30375 3496 30392
rect 3378 30306 3384 30323
rect 3490 30306 3496 30323
rect 3378 30236 3384 30254
rect 3490 30236 3496 30254
rect 3378 30166 3384 30184
rect 3490 30166 3496 30184
rect 3378 29380 3384 30114
rect 3490 29380 3496 30114
rect 3378 29368 3496 29380
rect 3655 30714 3773 30726
rect 3655 30680 3661 30714
rect 3695 30680 3733 30714
rect 3767 30680 3773 30714
rect 3655 30641 3773 30680
rect 3655 30607 3661 30641
rect 3695 30607 3733 30641
rect 3767 30607 3773 30641
rect 3655 30568 3773 30607
rect 3655 30534 3661 30568
rect 3695 30534 3733 30568
rect 3767 30534 3773 30568
rect 3655 30495 3773 30534
rect 3655 30461 3661 30495
rect 3695 30461 3733 30495
rect 3767 30461 3773 30495
rect 3655 30422 3773 30461
rect 3655 29982 3661 30422
rect 3767 29982 3773 30422
rect 3655 29913 3661 29930
rect 3767 29913 3773 29930
rect 3655 29844 3661 29861
rect 3767 29844 3773 29861
rect 3655 29775 3661 29792
rect 3767 29775 3773 29792
rect 3655 29706 3661 29723
rect 3767 29706 3773 29723
rect 3655 29636 3661 29654
rect 3767 29636 3773 29654
rect 3655 29566 3661 29584
rect 3767 29566 3773 29584
rect 3655 29496 3661 29514
rect 3767 29496 3773 29514
rect 3655 29426 3661 29444
rect 3767 29426 3773 29444
rect 3707 29374 3721 29380
rect 3655 29368 3773 29374
rect 3932 30720 4050 30726
rect 3984 30668 3998 30720
rect 3932 30651 4050 30668
rect 3984 30599 3998 30651
rect 3932 30582 4050 30599
rect 3984 30530 3998 30582
rect 3932 30513 4050 30530
rect 3984 30461 3998 30513
rect 3932 30444 4050 30461
rect 3984 30422 3998 30444
rect 3932 30375 3938 30392
rect 4044 30375 4050 30392
rect 3932 30306 3938 30323
rect 4044 30306 4050 30323
rect 3932 30236 3938 30254
rect 4044 30236 4050 30254
rect 3932 30166 3938 30184
rect 4044 30166 4050 30184
rect 3932 29380 3938 30114
rect 4044 29380 4050 30114
rect 3932 29368 4050 29380
rect 4209 30714 4327 30726
rect 4209 30680 4215 30714
rect 4249 30680 4287 30714
rect 4321 30680 4327 30714
rect 4209 30641 4327 30680
rect 4209 30607 4215 30641
rect 4249 30607 4287 30641
rect 4321 30607 4327 30641
rect 4209 30568 4327 30607
rect 4209 30534 4215 30568
rect 4249 30534 4287 30568
rect 4321 30534 4327 30568
rect 4209 30495 4327 30534
rect 4209 30461 4215 30495
rect 4249 30461 4287 30495
rect 4321 30461 4327 30495
rect 4209 30422 4327 30461
rect 4209 29982 4215 30422
rect 4321 29982 4327 30422
rect 4209 29913 4215 29930
rect 4321 29913 4327 29930
rect 4209 29844 4215 29861
rect 4321 29844 4327 29861
rect 4209 29775 4215 29792
rect 4321 29775 4327 29792
rect 4209 29706 4215 29723
rect 4321 29706 4327 29723
rect 4209 29636 4215 29654
rect 4321 29636 4327 29654
rect 4209 29566 4215 29584
rect 4321 29566 4327 29584
rect 4209 29496 4215 29514
rect 4321 29496 4327 29514
rect 4209 29426 4215 29444
rect 4321 29426 4327 29444
rect 4261 29374 4275 29380
rect 4209 29368 4327 29374
rect 4486 30720 4604 30726
rect 4538 30668 4552 30720
rect 4486 30651 4604 30668
rect 4538 30599 4552 30651
rect 4486 30582 4604 30599
rect 4538 30530 4552 30582
rect 4486 30513 4604 30530
rect 4538 30461 4552 30513
rect 4486 30444 4604 30461
rect 4538 30422 4552 30444
rect 4486 30375 4492 30392
rect 4598 30375 4604 30392
rect 4486 30306 4492 30323
rect 4598 30306 4604 30323
rect 4486 30236 4492 30254
rect 4598 30236 4604 30254
rect 4486 30166 4492 30184
rect 4598 30166 4604 30184
rect 4486 29380 4492 30114
rect 4598 29380 4604 30114
rect 4486 29368 4604 29380
rect 4763 30714 4881 30726
rect 4763 30680 4769 30714
rect 4803 30680 4841 30714
rect 4875 30680 4881 30714
rect 4763 30641 4881 30680
rect 4763 30607 4769 30641
rect 4803 30607 4841 30641
rect 4875 30607 4881 30641
rect 4763 30568 4881 30607
rect 4763 30534 4769 30568
rect 4803 30534 4841 30568
rect 4875 30534 4881 30568
rect 4763 30495 4881 30534
rect 4763 30461 4769 30495
rect 4803 30461 4841 30495
rect 4875 30461 4881 30495
rect 4763 30422 4881 30461
rect 4763 29982 4769 30422
rect 4875 29982 4881 30422
rect 4763 29913 4769 29930
rect 4875 29913 4881 29930
rect 4763 29844 4769 29861
rect 4875 29844 4881 29861
rect 4763 29775 4769 29792
rect 4875 29775 4881 29792
rect 4763 29706 4769 29723
rect 4875 29706 4881 29723
rect 4763 29636 4769 29654
rect 4875 29636 4881 29654
rect 4763 29566 4769 29584
rect 4875 29566 4881 29584
rect 4763 29496 4769 29514
rect 4875 29496 4881 29514
rect 4763 29426 4769 29444
rect 4875 29426 4881 29444
rect 4815 29374 4829 29380
rect 4763 29368 4881 29374
rect 5040 30720 5158 30726
rect 5092 30668 5106 30720
rect 5040 30651 5158 30668
rect 5092 30599 5106 30651
rect 5040 30582 5158 30599
rect 5092 30530 5106 30582
rect 5040 30513 5158 30530
rect 5092 30461 5106 30513
rect 5040 30444 5158 30461
rect 5092 30422 5106 30444
rect 5040 30375 5046 30392
rect 5152 30375 5158 30392
rect 5040 30306 5046 30323
rect 5152 30306 5158 30323
rect 5040 30236 5046 30254
rect 5152 30236 5158 30254
rect 5040 30166 5046 30184
rect 5152 30166 5158 30184
rect 5040 29380 5046 30114
rect 5152 29380 5158 30114
rect 5040 29368 5158 29380
rect 5317 30714 5435 30726
rect 5317 30680 5323 30714
rect 5357 30680 5395 30714
rect 5429 30680 5435 30714
rect 5317 30641 5435 30680
rect 5317 30607 5323 30641
rect 5357 30607 5395 30641
rect 5429 30607 5435 30641
rect 5317 30568 5435 30607
rect 5317 30534 5323 30568
rect 5357 30534 5395 30568
rect 5429 30534 5435 30568
rect 5317 30495 5435 30534
rect 5317 30461 5323 30495
rect 5357 30461 5395 30495
rect 5429 30461 5435 30495
rect 5317 30422 5435 30461
rect 5317 29982 5323 30422
rect 5429 29982 5435 30422
rect 5317 29913 5323 29930
rect 5429 29913 5435 29930
rect 5317 29844 5323 29861
rect 5429 29844 5435 29861
rect 5317 29775 5323 29792
rect 5429 29775 5435 29792
rect 5317 29706 5323 29723
rect 5429 29706 5435 29723
rect 5317 29636 5323 29654
rect 5429 29636 5435 29654
rect 5317 29566 5323 29584
rect 5429 29566 5435 29584
rect 5317 29496 5323 29514
rect 5429 29496 5435 29514
rect 5317 29426 5323 29444
rect 5429 29426 5435 29444
rect 5369 29374 5383 29380
rect 5317 29368 5435 29374
rect 5594 30720 5712 30726
rect 5646 30668 5660 30720
rect 5594 30651 5712 30668
rect 5646 30599 5660 30651
rect 5594 30582 5712 30599
rect 5646 30530 5660 30582
rect 5594 30513 5712 30530
rect 5646 30461 5660 30513
rect 5594 30444 5712 30461
rect 5646 30422 5660 30444
rect 5594 30375 5600 30392
rect 5706 30375 5712 30392
rect 5594 30306 5600 30323
rect 5706 30306 5712 30323
rect 5594 30236 5600 30254
rect 5706 30236 5712 30254
rect 5594 30166 5600 30184
rect 5706 30166 5712 30184
rect 5594 29380 5600 30114
rect 5706 29380 5712 30114
rect 5594 29368 5712 29380
rect 5871 30714 5989 30726
rect 5871 30680 5877 30714
rect 5911 30680 5949 30714
rect 5983 30680 5989 30714
rect 5871 30641 5989 30680
rect 5871 30607 5877 30641
rect 5911 30607 5949 30641
rect 5983 30607 5989 30641
rect 5871 30568 5989 30607
rect 5871 30534 5877 30568
rect 5911 30534 5949 30568
rect 5983 30534 5989 30568
rect 5871 30495 5989 30534
rect 5871 30461 5877 30495
rect 5911 30461 5949 30495
rect 5983 30461 5989 30495
rect 5871 30422 5989 30461
rect 5871 29982 5877 30422
rect 5983 29982 5989 30422
rect 5871 29913 5877 29930
rect 5983 29913 5989 29930
rect 5871 29844 5877 29861
rect 5983 29844 5989 29861
rect 5871 29775 5877 29792
rect 5983 29775 5989 29792
rect 5871 29706 5877 29723
rect 5983 29706 5989 29723
rect 5871 29636 5877 29654
rect 5983 29636 5989 29654
rect 5871 29566 5877 29584
rect 5983 29566 5989 29584
rect 5871 29496 5877 29514
rect 5983 29496 5989 29514
rect 5871 29426 5877 29444
rect 5983 29426 5989 29444
rect 5923 29374 5937 29380
rect 5871 29368 5989 29374
rect 6148 30720 6266 30726
rect 6200 30668 6214 30720
rect 6148 30651 6266 30668
rect 6200 30599 6214 30651
rect 6148 30582 6266 30599
rect 6200 30530 6214 30582
rect 6148 30513 6266 30530
rect 6200 30461 6214 30513
rect 6148 30444 6266 30461
rect 6200 30422 6214 30444
rect 6148 30375 6154 30392
rect 6260 30375 6266 30392
rect 6148 30306 6154 30323
rect 6260 30306 6266 30323
rect 6148 30236 6154 30254
rect 6260 30236 6266 30254
rect 6148 30166 6154 30184
rect 6260 30166 6266 30184
rect 6148 29380 6154 30114
rect 6260 29380 6266 30114
rect 6148 29368 6266 29380
rect 6425 30714 6543 30726
rect 6425 30680 6431 30714
rect 6465 30680 6503 30714
rect 6537 30680 6543 30714
rect 6425 30641 6543 30680
rect 6425 30607 6431 30641
rect 6465 30607 6503 30641
rect 6537 30607 6543 30641
rect 6425 30568 6543 30607
rect 6425 30534 6431 30568
rect 6465 30534 6503 30568
rect 6537 30534 6543 30568
rect 6425 30495 6543 30534
rect 6425 30461 6431 30495
rect 6465 30461 6503 30495
rect 6537 30461 6543 30495
rect 6425 30422 6543 30461
rect 6425 29982 6431 30422
rect 6537 29982 6543 30422
rect 6425 29913 6431 29930
rect 6537 29913 6543 29930
rect 6425 29844 6431 29861
rect 6537 29844 6543 29861
rect 6425 29775 6431 29792
rect 6537 29775 6543 29792
rect 6425 29706 6431 29723
rect 6537 29706 6543 29723
rect 6425 29636 6431 29654
rect 6537 29636 6543 29654
rect 6425 29566 6431 29584
rect 6537 29566 6543 29584
rect 6425 29496 6431 29514
rect 6537 29496 6543 29514
rect 6425 29426 6431 29444
rect 6537 29426 6543 29444
rect 6477 29374 6491 29380
rect 6425 29368 6543 29374
rect 6702 30720 6820 30726
rect 6754 30668 6768 30720
rect 6702 30651 6820 30668
rect 6754 30599 6768 30651
rect 6702 30582 6820 30599
rect 6754 30530 6768 30582
rect 6702 30513 6820 30530
rect 6754 30461 6768 30513
rect 6702 30444 6820 30461
rect 6754 30422 6768 30444
rect 6702 30375 6708 30392
rect 6814 30375 6820 30392
rect 6702 30306 6708 30323
rect 6814 30306 6820 30323
rect 6702 30236 6708 30254
rect 6814 30236 6820 30254
rect 6702 30166 6708 30184
rect 6814 30166 6820 30184
rect 6702 29380 6708 30114
rect 6814 29380 6820 30114
rect 6702 29368 6820 29380
rect 6979 30714 7097 30726
rect 6979 30680 6985 30714
rect 7019 30680 7057 30714
rect 7091 30680 7097 30714
rect 6979 30641 7097 30680
rect 6979 30607 6985 30641
rect 7019 30607 7057 30641
rect 7091 30607 7097 30641
rect 6979 30568 7097 30607
rect 6979 30534 6985 30568
rect 7019 30534 7057 30568
rect 7091 30534 7097 30568
rect 6979 30495 7097 30534
rect 6979 30461 6985 30495
rect 7019 30461 7057 30495
rect 7091 30461 7097 30495
rect 6979 30422 7097 30461
rect 6979 29982 6985 30422
rect 7091 29982 7097 30422
rect 6979 29913 6985 29930
rect 7091 29913 7097 29930
rect 6979 29844 6985 29861
rect 7091 29844 7097 29861
rect 6979 29775 6985 29792
rect 7091 29775 7097 29792
rect 6979 29706 6985 29723
rect 7091 29706 7097 29723
rect 6979 29636 6985 29654
rect 7091 29636 7097 29654
rect 6979 29566 6985 29584
rect 7091 29566 7097 29584
rect 6979 29496 6985 29514
rect 7091 29496 7097 29514
rect 6979 29426 6985 29444
rect 7091 29426 7097 29444
rect 7031 29374 7045 29380
rect 6979 29368 7097 29374
rect 7256 30720 7374 30726
rect 7308 30668 7322 30720
rect 7256 30651 7374 30668
rect 7308 30599 7322 30651
rect 7256 30582 7374 30599
rect 7308 30530 7322 30582
rect 7256 30513 7374 30530
rect 7308 30461 7322 30513
rect 7256 30444 7374 30461
rect 7308 30422 7322 30444
rect 7256 30375 7262 30392
rect 7368 30375 7374 30392
rect 7256 30306 7262 30323
rect 7368 30306 7374 30323
rect 7256 30236 7262 30254
rect 7368 30236 7374 30254
rect 7256 30166 7262 30184
rect 7368 30166 7374 30184
rect 7256 29380 7262 30114
rect 7368 29380 7374 30114
rect 7256 29368 7374 29380
rect 7533 30714 7651 30726
rect 7533 30680 7539 30714
rect 7573 30680 7611 30714
rect 7645 30680 7651 30714
rect 7533 30641 7651 30680
rect 7533 30607 7539 30641
rect 7573 30607 7611 30641
rect 7645 30607 7651 30641
rect 7533 30568 7651 30607
rect 7533 30534 7539 30568
rect 7573 30534 7611 30568
rect 7645 30534 7651 30568
rect 7533 30495 7651 30534
rect 7533 30461 7539 30495
rect 7573 30461 7611 30495
rect 7645 30461 7651 30495
rect 7533 30422 7651 30461
rect 7533 29982 7539 30422
rect 7645 29982 7651 30422
rect 7533 29913 7539 29930
rect 7645 29913 7651 29930
rect 7533 29844 7539 29861
rect 7645 29844 7651 29861
rect 7533 29775 7539 29792
rect 7645 29775 7651 29792
rect 7533 29706 7539 29723
rect 7645 29706 7651 29723
rect 7533 29636 7539 29654
rect 7645 29636 7651 29654
rect 7533 29566 7539 29584
rect 7645 29566 7651 29584
rect 7533 29496 7539 29514
rect 7645 29496 7651 29514
rect 7533 29426 7539 29444
rect 7645 29426 7651 29444
rect 7585 29374 7599 29380
rect 7533 29368 7651 29374
rect 7810 30720 7928 30726
rect 7862 30668 7876 30720
rect 7810 30651 7928 30668
rect 7862 30599 7876 30651
rect 7810 30582 7928 30599
rect 7862 30530 7876 30582
rect 7810 30513 7928 30530
rect 7862 30461 7876 30513
rect 7810 30444 7928 30461
rect 7862 30422 7876 30444
rect 7810 30375 7816 30392
rect 7922 30375 7928 30392
rect 7810 30306 7816 30323
rect 7922 30306 7928 30323
rect 7810 30236 7816 30254
rect 7922 30236 7928 30254
rect 7810 30166 7816 30184
rect 7922 30166 7928 30184
rect 7810 29380 7816 30114
rect 7922 29380 7928 30114
rect 7810 29368 7928 29380
rect 8044 30724 8050 30727
rect 8084 30724 8224 30727
rect 8044 30672 8047 30724
rect 8099 30672 8169 30724
rect 8221 30672 8224 30724
rect 8044 30655 8224 30672
rect 8044 30603 8047 30655
rect 8099 30603 8169 30655
rect 8221 30603 8224 30655
rect 8044 30586 8224 30603
rect 8044 30534 8047 30586
rect 8099 30534 8169 30586
rect 8221 30534 8224 30586
rect 8044 30517 8224 30534
rect 8044 30465 8047 30517
rect 8099 30465 8169 30517
rect 8221 30465 8224 30517
rect 8044 30448 8224 30465
rect 8044 30396 8047 30448
rect 8099 30396 8169 30448
rect 8221 30396 8224 30448
rect 8044 30395 8184 30396
rect 8218 30395 8224 30396
rect 8044 30378 8224 30395
rect 8044 30326 8047 30378
rect 8099 30326 8169 30378
rect 8221 30326 8224 30378
rect 8044 30323 8184 30326
rect 8218 30323 8224 30326
rect 8044 30308 8224 30323
rect 8044 30256 8047 30308
rect 8099 30256 8169 30308
rect 8221 30256 8224 30308
rect 8044 30251 8184 30256
rect 8218 30251 8224 30256
rect 8044 30238 8224 30251
rect 8044 30186 8047 30238
rect 8099 30186 8169 30238
rect 8221 30186 8224 30238
rect 8044 30179 8184 30186
rect 8218 30179 8224 30186
rect 8044 30168 8224 30179
rect 8044 30116 8047 30168
rect 8099 30116 8169 30168
rect 8221 30116 8224 30168
rect 8044 30107 8184 30116
rect 8218 30107 8224 30116
rect 8044 30079 8224 30107
rect 8044 30045 8050 30079
rect 8084 30069 8224 30079
rect 8084 30045 8184 30069
rect 8044 30035 8184 30045
rect 8218 30035 8224 30069
rect 8044 30007 8224 30035
rect 8044 29973 8050 30007
rect 8084 29997 8224 30007
rect 8084 29973 8184 29997
rect 8044 29963 8184 29973
rect 8218 29963 8224 29997
rect 8044 29935 8224 29963
rect 8044 29901 8050 29935
rect 8084 29925 8224 29935
rect 8084 29901 8184 29925
rect 8044 29891 8184 29901
rect 8218 29891 8224 29925
rect 8044 29863 8224 29891
rect 8044 29829 8050 29863
rect 8084 29853 8224 29863
rect 8084 29829 8184 29853
rect 8044 29819 8184 29829
rect 8218 29819 8224 29853
rect 8044 29791 8224 29819
rect 8044 29757 8050 29791
rect 8084 29781 8224 29791
rect 8084 29757 8184 29781
rect 8044 29747 8184 29757
rect 8218 29747 8224 29781
rect 8044 29719 8224 29747
rect 8044 29685 8050 29719
rect 8084 29709 8224 29719
rect 8084 29685 8184 29709
rect 8044 29675 8184 29685
rect 8218 29675 8224 29709
rect 8044 29647 8224 29675
rect 8044 29613 8050 29647
rect 8084 29637 8224 29647
rect 8084 29613 8184 29637
rect 8044 29603 8184 29613
rect 8218 29603 8224 29637
rect 8044 29575 8224 29603
rect 8044 29541 8050 29575
rect 8084 29565 8224 29575
rect 8084 29541 8184 29565
rect 8044 29531 8184 29541
rect 8218 29531 8224 29565
rect 8044 29503 8224 29531
rect 8044 29469 8050 29503
rect 8084 29493 8224 29503
rect 8084 29469 8184 29493
rect 8044 29459 8184 29469
rect 8218 29459 8224 29493
rect 8044 29431 8224 29459
rect 8044 29397 8050 29431
rect 8084 29421 8224 29431
rect 8084 29397 8184 29421
rect 8044 29387 8184 29397
rect 8218 29387 8224 29421
rect 8044 29359 8224 29387
rect 2543 29325 2729 29359
tri 2729 29325 2763 29359 sw
rect 8044 29325 8050 29359
rect 8084 29349 8224 29359
rect 8084 29325 8184 29349
rect 2543 29315 2763 29325
tri 2763 29315 2773 29325 sw
rect 8044 29315 8184 29325
rect 8218 29315 8224 29349
rect 2543 29310 2773 29315
tri 2773 29310 2778 29315 sw
rect 2543 29250 7729 29310
rect 2543 29216 3035 29250
rect 3069 29216 3108 29250
rect 3142 29216 3181 29250
rect 3215 29216 3254 29250
rect 3288 29216 3327 29250
rect 3361 29216 3400 29250
rect 3434 29216 3473 29250
rect 3507 29216 3546 29250
rect 3580 29216 3619 29250
rect 3653 29216 3692 29250
rect 3726 29216 3765 29250
rect 3799 29216 3838 29250
rect 3872 29216 3911 29250
rect 3945 29216 3984 29250
rect 4018 29216 4057 29250
rect 4091 29216 4130 29250
rect 4164 29216 4203 29250
rect 4237 29216 4276 29250
rect 4310 29216 4349 29250
rect 4383 29216 4422 29250
rect 4456 29216 4495 29250
rect 4529 29216 4568 29250
rect 4602 29216 4641 29250
rect 4675 29216 4714 29250
rect 4748 29216 4787 29250
rect 4821 29216 4860 29250
rect 4894 29216 4933 29250
rect 4967 29216 5006 29250
rect 5040 29216 5079 29250
rect 5113 29216 5152 29250
rect 5186 29216 5225 29250
rect 5259 29216 5298 29250
rect 5332 29216 5371 29250
rect 5405 29216 5444 29250
rect 5478 29216 5517 29250
rect 5551 29216 5590 29250
rect 5624 29216 5663 29250
rect 5697 29216 5736 29250
rect 5770 29216 5809 29250
rect 5843 29216 5882 29250
rect 5916 29216 5955 29250
rect 5989 29216 6027 29250
rect 6061 29216 6099 29250
rect 6133 29216 6171 29250
rect 6205 29216 6243 29250
rect 6277 29216 6315 29250
rect 6349 29216 6387 29250
rect 6421 29216 6459 29250
rect 6493 29216 6531 29250
rect 6565 29216 6603 29250
rect 6637 29216 6675 29250
rect 6709 29216 6747 29250
rect 6781 29216 6819 29250
rect 6853 29216 6891 29250
rect 6925 29216 6963 29250
rect 6997 29216 7035 29250
rect 7069 29216 7107 29250
rect 7141 29216 7179 29250
rect 7213 29216 7251 29250
rect 7285 29216 7323 29250
rect 7357 29216 7395 29250
rect 7429 29216 7467 29250
rect 7501 29216 7539 29250
rect 7573 29216 7611 29250
rect 7645 29216 7683 29250
rect 7717 29216 7729 29250
rect 2543 29190 7729 29216
rect 8044 29287 8224 29315
rect 8044 29253 8050 29287
rect 8084 29277 8224 29287
rect 8084 29253 8184 29277
rect 8044 29243 8184 29253
rect 8218 29243 8224 29277
rect 8044 29215 8224 29243
rect 2543 29181 4985 29190
tri 4985 29181 4994 29190 nw
rect 8044 29181 8050 29215
rect 8084 29205 8224 29215
rect 8084 29181 8184 29205
rect 2543 29171 4975 29181
tri 4975 29171 4985 29181 nw
rect 8044 29171 8184 29181
rect 8218 29171 8224 29205
rect 2543 29143 4947 29171
tri 4947 29143 4975 29171 nw
rect 8044 29143 8224 29171
rect 2543 29103 4928 29143
tri 4928 29124 4947 29143 nw
rect 2270 29066 2276 29100
rect 2310 29066 2410 29100
rect 2444 29066 2450 29100
tri 4723 29099 4727 29103 ne
rect 4727 29099 4928 29103
tri 4727 29071 4755 29099 ne
rect 4755 29071 4928 29099
rect 2270 29028 2450 29066
tri 4755 29053 4773 29071 ne
rect 2270 28994 2276 29028
rect 2310 28994 2410 29028
rect 2444 28994 2450 29028
rect 2270 28956 2450 28994
rect 2270 28922 2276 28956
rect 2310 28922 2410 28956
rect 2444 28922 2450 28956
rect 2270 28884 2450 28922
rect 2270 28850 2276 28884
rect 2310 28850 2410 28884
rect 2444 28850 2450 28884
rect 2270 28812 2450 28850
rect 2270 28778 2276 28812
rect 2310 28778 2410 28812
rect 2444 28778 2450 28812
rect 2270 28740 2450 28778
rect 2270 28724 2276 28740
rect 2310 28724 2410 28740
rect 2322 28672 2392 28724
rect 2444 28672 2450 28740
rect 2270 28668 2450 28672
rect 2270 28655 2276 28668
rect 2310 28655 2410 28668
rect 2322 28603 2392 28655
rect 2444 28603 2450 28668
rect 2270 28596 2450 28603
rect 2270 28586 2276 28596
rect 2310 28586 2410 28596
rect 2322 28534 2392 28586
rect 2444 28534 2450 28596
rect 2270 28524 2450 28534
rect 2270 28517 2276 28524
rect 2310 28517 2410 28524
rect 2322 28465 2392 28517
rect 2444 28465 2450 28524
rect 2270 28452 2450 28465
rect 2270 28448 2276 28452
rect 2310 28448 2410 28452
rect 2322 28396 2392 28448
rect 2444 28396 2450 28452
rect 2270 28380 2450 28396
rect 2270 28378 2276 28380
rect 2310 28378 2410 28380
rect 2322 28326 2392 28378
rect 2444 28326 2450 28380
rect 2270 28308 2450 28326
rect 2322 28256 2392 28308
rect 2444 28256 2450 28308
rect 2270 28238 2450 28256
rect 2322 28186 2392 28238
rect 2444 28186 2450 28238
rect 2270 28168 2450 28186
rect 2322 28116 2392 28168
rect 2444 28116 2450 28168
rect 2270 28092 2450 28116
rect 2270 28058 2276 28092
rect 2310 28058 2410 28092
rect 2444 28058 2450 28092
rect 2270 28020 2450 28058
rect 2270 27986 2276 28020
rect 2310 27986 2410 28020
rect 2444 27986 2450 28020
rect 2270 27948 2450 27986
rect 2270 27914 2276 27948
rect 2310 27914 2410 27948
rect 2444 27914 2450 27948
rect 2270 27876 2450 27914
rect 2270 27842 2276 27876
rect 2310 27842 2410 27876
rect 2444 27842 2450 27876
rect 2270 27804 2450 27842
rect 2270 27770 2276 27804
rect 2310 27770 2410 27804
rect 2444 27770 2450 27804
rect 2270 27732 2450 27770
rect 2270 27698 2276 27732
rect 2310 27698 2410 27732
rect 2444 27698 2450 27732
rect 2270 27660 2450 27698
rect 2270 27626 2276 27660
rect 2310 27626 2410 27660
rect 2444 27626 2450 27660
rect 2270 27588 2450 27626
rect 2270 27554 2276 27588
rect 2310 27554 2410 27588
rect 2444 27554 2450 27588
rect 2270 27516 2450 27554
rect 2270 27482 2276 27516
rect 2310 27482 2410 27516
rect 2444 27482 2450 27516
rect 2270 27444 2450 27482
rect 2270 27410 2276 27444
rect 2310 27410 2410 27444
rect 2444 27410 2450 27444
rect 2270 27372 2450 27410
rect 2270 27338 2276 27372
rect 2310 27338 2410 27372
rect 2444 27338 2450 27372
rect 2270 27300 2450 27338
rect 2270 27266 2276 27300
rect 2310 27266 2410 27300
rect 2444 27266 2450 27300
rect 2270 27228 2450 27266
rect 2270 27194 2276 27228
rect 2310 27194 2410 27228
rect 2444 27194 2450 27228
rect 2270 27156 2450 27194
rect 2270 27122 2276 27156
rect 2310 27122 2410 27156
rect 2444 27122 2450 27156
rect 2270 27084 2450 27122
rect 2270 27050 2276 27084
rect 2310 27050 2410 27084
rect 2444 27050 2450 27084
rect 2270 27012 2450 27050
rect 2270 26978 2276 27012
rect 2310 26978 2410 27012
rect 2444 26978 2450 27012
rect 2270 26940 2450 26978
rect 2270 26906 2276 26940
rect 2310 26906 2410 26940
rect 2444 26906 2450 26940
rect 2270 26868 2450 26906
rect 2270 26834 2276 26868
rect 2310 26834 2410 26868
rect 2444 26834 2450 26868
rect 2270 26796 2450 26834
rect 2270 26762 2276 26796
rect 2310 26762 2410 26796
rect 2444 26762 2450 26796
rect 2270 26724 2450 26762
rect 2322 26672 2392 26724
rect 2444 26672 2450 26724
rect 2270 26655 2450 26672
rect 2322 26603 2392 26655
rect 2444 26603 2450 26655
rect 2270 26586 2450 26603
rect 2322 26534 2392 26586
rect 2444 26534 2450 26586
rect 2270 26517 2450 26534
rect 2322 26465 2392 26517
rect 2444 26465 2450 26517
rect 2270 26448 2450 26465
rect 2322 26396 2392 26448
rect 2444 26396 2450 26448
rect 2270 26378 2450 26396
rect 2322 26326 2392 26378
rect 2444 26326 2450 26378
rect 2270 26308 2450 26326
rect 2322 26256 2392 26308
rect 2444 26256 2450 26308
rect 2270 26238 2450 26256
rect 2322 26186 2392 26238
rect 2444 26186 2450 26238
rect 2270 26168 2450 26186
rect 2322 26116 2392 26168
rect 2270 26114 2276 26116
rect 2310 26114 2410 26116
rect 2444 26114 2450 26168
rect 2270 26076 2450 26114
rect 2270 26042 2276 26076
rect 2310 26042 2410 26076
rect 2444 26042 2450 26076
rect 2270 26004 2450 26042
rect 2270 25970 2276 26004
rect 2310 25970 2410 26004
rect 2444 25970 2450 26004
rect 2270 25932 2450 25970
rect 2270 25898 2276 25932
rect 2310 25898 2410 25932
rect 2444 25898 2450 25932
rect 2270 25860 2450 25898
rect 2270 25826 2276 25860
rect 2310 25826 2410 25860
rect 2444 25826 2450 25860
rect 2270 25788 2450 25826
rect 2270 25754 2276 25788
rect 2310 25754 2410 25788
rect 2444 25754 2450 25788
rect 2270 25716 2450 25754
rect 2270 25682 2276 25716
rect 2310 25682 2410 25716
rect 2444 25682 2450 25716
rect 2270 25644 2450 25682
rect 2270 25610 2276 25644
rect 2310 25610 2410 25644
rect 2444 25610 2450 25644
rect 2270 25572 2450 25610
rect 2270 25538 2276 25572
rect 2310 25538 2410 25572
rect 2444 25538 2450 25572
rect 2270 25500 2450 25538
rect 2270 25466 2276 25500
rect 2310 25466 2410 25500
rect 2444 25466 2450 25500
rect 2270 25428 2450 25466
rect 2270 25394 2276 25428
rect 2310 25394 2410 25428
rect 2444 25394 2450 25428
rect 2270 25356 2450 25394
rect 2270 25322 2276 25356
rect 2310 25322 2410 25356
rect 2444 25322 2450 25356
rect 2270 25284 2450 25322
rect 2270 25250 2276 25284
rect 2310 25250 2410 25284
rect 2444 25250 2450 25284
rect 2270 25212 2450 25250
rect 2270 25178 2276 25212
rect 2310 25178 2410 25212
rect 2444 25178 2450 25212
rect 2270 25140 2450 25178
rect 2270 25106 2276 25140
rect 2310 25106 2410 25140
rect 2444 25106 2450 25140
rect 2270 25068 2450 25106
rect 2270 25034 2276 25068
rect 2310 25034 2410 25068
rect 2444 25034 2450 25068
rect 2270 24996 2450 25034
rect 2270 24962 2276 24996
rect 2310 24962 2410 24996
rect 2444 24962 2450 24996
rect 2270 24924 2450 24962
rect 2270 24890 2276 24924
rect 2310 24890 2410 24924
rect 2444 24890 2450 24924
rect 2270 24852 2450 24890
rect 2270 24818 2276 24852
rect 2310 24818 2410 24852
rect 2444 24818 2450 24852
rect 2270 24780 2450 24818
rect 2270 24746 2276 24780
rect 2310 24746 2410 24780
rect 2444 24746 2450 24780
rect 2270 24724 2450 24746
rect 2322 24672 2392 24724
rect 2444 24672 2450 24724
rect 2270 24655 2450 24672
rect 2322 24603 2392 24655
rect 2270 24602 2276 24603
rect 2310 24602 2410 24603
rect 2444 24602 2450 24655
rect 2270 24586 2450 24602
rect 2322 24534 2392 24586
rect 2270 24530 2276 24534
rect 2310 24530 2410 24534
rect 2444 24530 2450 24586
rect 2270 24517 2450 24530
rect 2322 24465 2392 24517
rect 2270 24458 2276 24465
rect 2310 24458 2410 24465
rect 2444 24458 2450 24517
rect 2270 24448 2450 24458
rect 2322 24396 2392 24448
rect 2270 24386 2276 24396
rect 2310 24386 2410 24396
rect 2444 24386 2450 24448
rect 2270 24378 2450 24386
rect 2322 24326 2392 24378
rect 2270 24314 2276 24326
rect 2310 24314 2410 24326
rect 2444 24314 2450 24378
rect 2270 24308 2450 24314
rect 2322 24256 2392 24308
rect 2270 24242 2276 24256
rect 2310 24242 2410 24256
rect 2444 24242 2450 24308
rect 2270 24238 2450 24242
rect 2322 24186 2392 24238
rect 2270 24170 2276 24186
rect 2310 24170 2410 24186
rect 2444 24170 2450 24238
rect 2270 24168 2450 24170
rect 2322 24116 2392 24168
rect 2270 24098 2276 24116
rect 2310 24098 2410 24116
rect 2444 24098 2450 24168
rect 2270 24060 2450 24098
rect 2270 24026 2276 24060
rect 2310 24026 2410 24060
rect 2444 24026 2450 24060
rect 2270 23988 2450 24026
rect 2270 23954 2276 23988
rect 2310 23954 2410 23988
rect 2444 23954 2450 23988
rect 2270 23916 2450 23954
rect 2270 23882 2276 23916
rect 2310 23882 2410 23916
rect 2444 23882 2450 23916
rect 2270 23844 2450 23882
rect 2270 23810 2276 23844
rect 2310 23810 2410 23844
rect 2444 23810 2450 23844
rect 2270 23772 2450 23810
rect 2270 23738 2276 23772
rect 2310 23738 2410 23772
rect 2444 23738 2450 23772
rect 2270 23700 2450 23738
rect 2270 23666 2276 23700
rect 2310 23666 2410 23700
rect 2444 23666 2450 23700
rect 2270 23628 2450 23666
rect 2270 23594 2276 23628
rect 2310 23594 2410 23628
rect 2444 23594 2450 23628
rect 2270 23556 2450 23594
rect 2270 23522 2276 23556
rect 2310 23522 2410 23556
rect 2444 23522 2450 23556
rect 2270 23484 2450 23522
rect 2270 23450 2276 23484
rect 2310 23450 2410 23484
rect 2444 23450 2450 23484
rect 2270 23412 2450 23450
rect 2270 23378 2276 23412
rect 2310 23378 2410 23412
rect 2444 23378 2450 23412
rect 2270 23340 2450 23378
rect 2270 23306 2276 23340
rect 2310 23306 2410 23340
rect 2444 23306 2450 23340
rect 2270 23268 2450 23306
rect 2270 23234 2276 23268
rect 2310 23234 2410 23268
rect 2444 23234 2450 23268
rect 2270 23196 2450 23234
rect 2270 23162 2276 23196
rect 2310 23162 2410 23196
rect 2444 23162 2450 23196
rect 2270 23124 2450 23162
rect 2270 23090 2276 23124
rect 2310 23090 2410 23124
rect 2444 23090 2450 23124
rect 2270 23052 2450 23090
rect 2270 23018 2276 23052
rect 2310 23018 2410 23052
rect 2444 23018 2450 23052
rect 2270 22980 2450 23018
rect 2270 22946 2276 22980
rect 2310 22946 2410 22980
rect 2444 22946 2450 22980
rect 2270 22908 2450 22946
rect 2270 22874 2276 22908
rect 2310 22874 2410 22908
rect 2444 22874 2450 22908
rect 2270 22836 2450 22874
rect 2270 22802 2276 22836
rect 2310 22802 2410 22836
rect 2444 22802 2450 22836
rect 2270 22764 2450 22802
rect 2270 22730 2276 22764
rect 2310 22730 2410 22764
rect 2444 22730 2450 22764
rect 2270 22724 2450 22730
rect 2322 22672 2392 22724
rect 2270 22658 2276 22672
rect 2310 22658 2410 22672
rect 2444 22658 2450 22724
rect 2270 22655 2450 22658
rect 2322 22603 2392 22655
rect 2270 22586 2276 22603
rect 2310 22586 2410 22603
rect 2322 22534 2392 22586
rect 2270 22517 2276 22534
rect 2310 22517 2410 22534
rect 2322 22465 2392 22517
rect 2270 22448 2276 22465
rect 2310 22448 2410 22465
rect 2322 22396 2392 22448
rect 2270 22378 2276 22396
rect 2310 22378 2410 22396
rect 2322 22326 2392 22378
rect 2270 22308 2276 22326
rect 2310 22308 2410 22326
rect 2322 22256 2392 22308
rect 2270 22238 2276 22256
rect 2310 22238 2410 22256
rect 2322 22186 2392 22238
rect 2270 22168 2276 22186
rect 2310 22168 2410 22186
rect 2322 22116 2392 22168
rect 2270 22082 2276 22116
rect 2310 22082 2410 22116
rect 2444 22082 2450 22655
rect 2270 22044 2450 22082
rect 2270 22010 2276 22044
rect 2310 22010 2410 22044
rect 2444 22010 2450 22044
rect 2270 21972 2450 22010
rect 2270 21938 2276 21972
rect 2310 21938 2410 21972
rect 2444 21938 2450 21972
rect 2270 21900 2450 21938
rect 2270 21866 2276 21900
rect 2310 21866 2410 21900
rect 2444 21866 2450 21900
rect 2270 21828 2450 21866
rect 2270 21794 2276 21828
rect 2310 21794 2410 21828
rect 2444 21794 2450 21828
rect 2270 21756 2450 21794
rect 2270 21722 2276 21756
rect 2310 21722 2410 21756
rect 2444 21722 2450 21756
rect 2270 21684 2450 21722
rect 2270 21650 2276 21684
rect 2310 21650 2410 21684
rect 2444 21650 2450 21684
rect 2270 21612 2450 21650
rect 2270 21578 2276 21612
rect 2310 21578 2410 21612
rect 2444 21578 2450 21612
rect 2270 21540 2450 21578
rect 2270 21506 2276 21540
rect 2310 21506 2410 21540
rect 2444 21506 2450 21540
rect 2270 21468 2450 21506
rect 2270 21434 2276 21468
rect 2310 21434 2410 21468
rect 2444 21434 2450 21468
rect 2270 21396 2450 21434
rect 2270 21362 2276 21396
rect 2310 21362 2410 21396
rect 2444 21362 2450 21396
rect 2270 21324 2450 21362
rect 2270 21290 2276 21324
rect 2310 21290 2410 21324
rect 2444 21290 2450 21324
rect 2270 21252 2450 21290
rect 2270 21218 2276 21252
rect 2310 21218 2410 21252
rect 2444 21218 2450 21252
rect 2270 21180 2450 21218
rect 2270 21146 2276 21180
rect 2310 21146 2410 21180
rect 2444 21146 2450 21180
rect 2270 21108 2450 21146
rect 2270 21074 2276 21108
rect 2310 21074 2410 21108
rect 2444 21074 2450 21108
rect 2270 21036 2450 21074
rect 2270 21002 2276 21036
rect 2310 21002 2410 21036
rect 2444 21002 2450 21036
rect 2270 20964 2450 21002
rect 2270 20930 2276 20964
rect 2310 20930 2410 20964
rect 2444 20930 2450 20964
rect 2270 20892 2450 20930
rect 2270 20858 2276 20892
rect 2310 20858 2410 20892
rect 2444 20858 2450 20892
rect 2270 20820 2450 20858
rect 2270 20786 2276 20820
rect 2310 20786 2410 20820
rect 2444 20786 2450 20820
rect 2270 20748 2450 20786
rect 2270 20724 2276 20748
rect 2310 20724 2410 20748
rect 2322 20672 2392 20724
rect 2270 20655 2276 20672
rect 2310 20655 2410 20672
rect 2322 20603 2392 20655
rect 2270 20586 2276 20603
rect 2310 20586 2410 20603
rect 2322 20534 2392 20586
rect 2444 20534 2450 20748
rect 2270 20532 2450 20534
rect 2270 20517 2276 20532
rect 2310 20517 2410 20532
rect 2322 20465 2392 20517
rect 2444 20465 2450 20532
rect 2270 20460 2450 20465
rect 2270 20448 2276 20460
rect 2310 20448 2410 20460
rect 2322 20396 2392 20448
rect 2444 20396 2450 20460
rect 2270 20388 2450 20396
rect 2270 20378 2276 20388
rect 2310 20378 2410 20388
rect 2322 20326 2392 20378
rect 2444 20326 2450 20388
rect 2270 20316 2450 20326
rect 2270 20308 2276 20316
rect 2310 20308 2410 20316
rect 2322 20256 2392 20308
rect 2444 20256 2450 20316
rect 2270 20244 2450 20256
rect 2270 20238 2276 20244
rect 2310 20238 2410 20244
rect 2322 20186 2392 20238
rect 2444 20186 2450 20244
rect 2270 20172 2450 20186
rect 2270 20168 2276 20172
rect 2310 20168 2410 20172
rect 2322 20116 2392 20168
rect 2444 20116 2450 20172
rect 2270 20100 2450 20116
rect 2270 20066 2276 20100
rect 2310 20066 2410 20100
rect 2444 20066 2450 20100
rect 2270 20028 2450 20066
rect 2270 19994 2276 20028
rect 2310 19994 2410 20028
rect 2444 19994 2450 20028
rect 2270 19956 2450 19994
rect 2270 19922 2276 19956
rect 2310 19922 2410 19956
rect 2444 19922 2450 19956
rect 2270 19884 2450 19922
rect 2270 19850 2276 19884
rect 2310 19850 2410 19884
rect 2444 19850 2450 19884
rect 2270 19812 2450 19850
rect 2270 19778 2276 19812
rect 2310 19778 2410 19812
rect 2444 19778 2450 19812
rect 2270 19740 2450 19778
rect 2270 19706 2276 19740
rect 2310 19706 2410 19740
rect 2444 19706 2450 19740
rect 2270 19668 2450 19706
rect 2270 19634 2276 19668
rect 2310 19634 2410 19668
rect 2444 19634 2450 19668
rect 2270 19596 2450 19634
rect 2270 19562 2276 19596
rect 2310 19562 2410 19596
rect 2444 19562 2450 19596
rect 2270 19524 2450 19562
rect 2270 19490 2276 19524
rect 2310 19490 2410 19524
rect 2444 19490 2450 19524
rect 2270 19452 2450 19490
rect 2270 19418 2276 19452
rect 2310 19418 2410 19452
rect 2444 19418 2450 19452
rect 2270 19380 2450 19418
rect 2270 19346 2276 19380
rect 2310 19346 2410 19380
rect 2444 19346 2450 19380
rect 2270 19308 2450 19346
rect 2270 19274 2276 19308
rect 2310 19274 2410 19308
rect 2444 19274 2450 19308
rect 2270 19236 2450 19274
rect 2270 19202 2276 19236
rect 2310 19202 2410 19236
rect 2444 19202 2450 19236
rect 2270 19164 2450 19202
rect 2270 19130 2276 19164
rect 2310 19130 2410 19164
rect 2444 19130 2450 19164
rect 2270 19092 2450 19130
rect 2270 19058 2276 19092
rect 2310 19058 2410 19092
rect 2444 19058 2450 19092
rect 2270 19020 2450 19058
rect 2270 18986 2276 19020
rect 2310 18986 2410 19020
rect 2444 18986 2450 19020
rect 2270 18948 2450 18986
rect 2270 18914 2276 18948
rect 2310 18914 2410 18948
rect 2444 18914 2450 18948
rect 2270 18876 2450 18914
rect 2270 18842 2276 18876
rect 2310 18842 2410 18876
rect 2444 18842 2450 18876
rect 2270 18804 2450 18842
rect 2270 18770 2276 18804
rect 2310 18770 2410 18804
rect 2444 18770 2450 18804
rect 2270 18732 2450 18770
rect 2270 18724 2276 18732
rect 2310 18724 2410 18732
rect 2322 18672 2392 18724
rect 2444 18672 2450 18732
rect 2270 18660 2450 18672
rect 2270 18655 2276 18660
rect 2310 18655 2410 18660
rect 2322 18603 2392 18655
rect 2444 18603 2450 18660
rect 2270 18588 2450 18603
rect 2270 18586 2276 18588
rect 2310 18586 2410 18588
rect 2322 18534 2392 18586
rect 2444 18534 2450 18588
rect 2270 18517 2450 18534
rect 2322 18465 2392 18517
rect 2444 18465 2450 18517
rect 2270 18448 2450 18465
rect 2322 18396 2392 18448
rect 2444 18396 2450 18448
rect 2270 18378 2450 18396
rect 2322 18326 2392 18378
rect 2444 18326 2450 18378
rect 2270 18308 2450 18326
rect 2322 18256 2392 18308
rect 2444 18256 2450 18308
rect 2270 18238 2450 18256
rect 2322 18186 2392 18238
rect 2444 18186 2450 18238
rect 2270 18168 2450 18186
rect 2322 18116 2392 18168
rect 2444 18116 2450 18168
rect 2270 18084 2450 18116
rect 2270 18050 2276 18084
rect 2310 18050 2410 18084
rect 2444 18050 2450 18084
rect 2270 18012 2450 18050
rect 2270 17978 2276 18012
rect 2310 17978 2410 18012
rect 2444 17978 2450 18012
rect 2270 17940 2450 17978
rect 2270 17906 2276 17940
rect 2310 17906 2410 17940
rect 2444 17906 2450 17940
rect 2270 17868 2450 17906
rect 2270 17834 2276 17868
rect 2310 17834 2410 17868
rect 2444 17834 2450 17868
rect 2270 17796 2450 17834
rect 2270 17762 2276 17796
rect 2310 17762 2410 17796
rect 2444 17762 2450 17796
rect 2270 17724 2450 17762
rect 2270 17690 2276 17724
rect 2310 17690 2410 17724
rect 2444 17690 2450 17724
rect 2270 17652 2450 17690
rect 2270 17618 2276 17652
rect 2310 17618 2410 17652
rect 2444 17618 2450 17652
rect 2270 17580 2450 17618
rect 2270 17546 2276 17580
rect 2310 17546 2410 17580
rect 2444 17546 2450 17580
rect 2270 17508 2450 17546
rect 2270 17474 2276 17508
rect 2310 17474 2410 17508
rect 2444 17474 2450 17508
rect 2270 17436 2450 17474
rect 2270 17402 2276 17436
rect 2310 17402 2410 17436
rect 2444 17402 2450 17436
rect 2270 17364 2450 17402
rect 2270 17330 2276 17364
rect 2310 17330 2410 17364
rect 2444 17330 2450 17364
rect 2270 17292 2450 17330
rect 2270 17258 2276 17292
rect 2310 17258 2410 17292
rect 2444 17258 2450 17292
rect 2270 17220 2450 17258
rect 2270 17186 2276 17220
rect 2310 17186 2410 17220
rect 2444 17186 2450 17220
rect 2270 17148 2450 17186
rect 2270 17114 2276 17148
rect 2310 17114 2410 17148
rect 2444 17114 2450 17148
rect 2270 17076 2450 17114
rect 2270 17042 2276 17076
rect 2310 17042 2410 17076
rect 2444 17042 2450 17076
rect 2270 17004 2450 17042
rect 2270 16973 2276 17004
rect 2310 16973 2410 17004
rect 2322 16921 2392 16973
rect 2270 16907 2276 16921
rect 2310 16907 2410 16921
rect 2322 16855 2392 16907
rect 2270 16841 2276 16855
rect 2310 16841 2410 16855
rect 2322 16789 2392 16841
rect 2444 16789 2450 17004
rect 2270 16788 2450 16789
rect 2270 16775 2276 16788
rect 2310 16775 2410 16788
rect 2322 16723 2392 16775
rect 2444 16723 2450 16788
rect 2270 16716 2450 16723
rect 2270 16709 2276 16716
rect 2310 16709 2410 16716
rect 2322 16657 2392 16709
rect 2444 16657 2450 16716
rect 2270 16644 2450 16657
rect 2270 16643 2276 16644
rect 2310 16643 2410 16644
rect 2322 16591 2392 16643
rect 2444 16591 2450 16644
rect 2270 16577 2450 16591
rect 2322 16525 2392 16577
rect 2444 16525 2450 16577
rect 2270 16511 2450 16525
rect 2322 16459 2392 16511
rect 2444 16459 2450 16511
rect 2270 16445 2450 16459
rect 2322 16393 2392 16445
rect 2444 16393 2450 16445
rect 2270 16378 2450 16393
rect 2322 16326 2392 16378
rect 2270 16322 2276 16326
rect 2310 16322 2410 16326
rect 2444 16322 2450 16378
rect 2270 16311 2450 16322
rect 2322 16259 2392 16311
rect 2270 16250 2276 16259
rect 2310 16250 2410 16259
rect 2444 16250 2450 16311
rect 2270 16244 2450 16250
rect 2322 16192 2392 16244
rect 2270 16178 2276 16192
rect 2310 16178 2410 16192
rect 2444 16178 2450 16244
rect 2270 16177 2450 16178
rect 2322 16125 2392 16177
rect 2270 16110 2276 16125
rect 2310 16110 2410 16125
rect 2322 16058 2392 16110
rect 2270 16043 2276 16058
rect 2310 16043 2410 16058
rect 2322 15991 2392 16043
rect 2270 15962 2276 15991
rect 2310 15962 2410 15991
rect 2444 15962 2450 16177
rect 2270 15924 2450 15962
rect 2270 15890 2276 15924
rect 2310 15890 2410 15924
rect 2444 15890 2450 15924
rect 2642 28965 4590 28977
rect 2642 26728 2663 28965
rect 4569 26728 4590 28965
rect 2642 26676 2648 26728
rect 4584 26676 4590 26728
rect 2642 26660 2663 26676
rect 4569 26660 4590 26676
rect 2642 26608 2648 26660
rect 4584 26608 4590 26660
rect 2642 26592 2663 26608
rect 4569 26592 4590 26608
rect 2642 26540 2648 26592
rect 4584 26540 4590 26592
rect 2642 26524 2663 26540
rect 4569 26524 4590 26540
rect 2642 26472 2648 26524
rect 4584 26472 4590 26524
rect 2642 26456 2663 26472
rect 4569 26456 4590 26472
rect 2642 26404 2648 26456
rect 4584 26404 4590 26456
rect 2642 26388 2663 26404
rect 4569 26388 4590 26404
rect 2642 26336 2648 26388
rect 4584 26336 4590 26388
rect 2642 26320 2663 26336
rect 4569 26320 4590 26336
rect 2642 26268 2648 26320
rect 4584 26268 4590 26320
rect 2642 26252 2663 26268
rect 4569 26252 4590 26268
rect 2642 26200 2648 26252
rect 4584 26200 4590 26252
rect 2642 24728 2663 26200
rect 4569 24728 4590 26200
rect 2642 24676 2648 24728
rect 4584 24676 4590 24728
rect 2642 24660 2663 24676
rect 4569 24660 4590 24676
rect 2642 24608 2648 24660
rect 4584 24608 4590 24660
rect 2642 24592 2663 24608
rect 4569 24592 4590 24608
rect 2642 24540 2648 24592
rect 4584 24540 4590 24592
rect 2642 24524 2663 24540
rect 4569 24524 4590 24540
rect 2642 24472 2648 24524
rect 4584 24472 4590 24524
rect 2642 24456 2663 24472
rect 4569 24456 4590 24472
rect 2642 24404 2648 24456
rect 4584 24404 4590 24456
rect 2642 24388 2663 24404
rect 4569 24388 4590 24404
rect 2642 24336 2648 24388
rect 4584 24336 4590 24388
rect 2642 24320 2663 24336
rect 4569 24320 4590 24336
rect 2642 24268 2648 24320
rect 4584 24268 4590 24320
rect 2642 24252 2663 24268
rect 4569 24252 4590 24268
rect 2642 24200 2648 24252
rect 4584 24200 4590 24252
rect 2642 22728 2663 24200
rect 4569 22728 4590 24200
rect 2642 22676 2648 22728
rect 4584 22676 4590 22728
rect 2642 22660 2663 22676
rect 4569 22660 4590 22676
rect 2642 22608 2648 22660
rect 4584 22608 4590 22660
rect 2642 22592 2663 22608
rect 4569 22592 4590 22608
rect 2642 22540 2648 22592
rect 4584 22540 4590 22592
rect 2642 22524 2663 22540
rect 4569 22524 4590 22540
rect 2642 22472 2648 22524
rect 4584 22472 4590 22524
rect 2642 22456 2663 22472
rect 4569 22456 4590 22472
rect 2642 22404 2648 22456
rect 4584 22404 4590 22456
rect 2642 22388 2663 22404
rect 4569 22388 4590 22404
rect 2642 22336 2648 22388
rect 4584 22336 4590 22388
rect 2642 22320 2663 22336
rect 4569 22320 4590 22336
rect 2642 22268 2648 22320
rect 4584 22268 4590 22320
rect 2642 22252 2663 22268
rect 4569 22252 4590 22268
rect 2642 22200 2648 22252
rect 4584 22200 4590 22252
rect 2642 20728 2663 22200
rect 4569 20728 4590 22200
rect 2642 20676 2648 20728
rect 4584 20676 4590 20728
rect 2642 20660 2663 20676
rect 4569 20660 4590 20676
rect 2642 20608 2648 20660
rect 4584 20608 4590 20660
rect 2642 20592 2663 20608
rect 4569 20592 4590 20608
rect 2642 20540 2648 20592
rect 4584 20540 4590 20592
rect 2642 20524 2663 20540
rect 4569 20524 4590 20540
rect 2642 20472 2648 20524
rect 4584 20472 4590 20524
rect 2642 20456 2663 20472
rect 4569 20456 4590 20472
rect 2642 20404 2648 20456
rect 4584 20404 4590 20456
rect 2642 20388 2663 20404
rect 4569 20388 4590 20404
rect 2642 20336 2648 20388
rect 4584 20336 4590 20388
rect 2642 20320 2663 20336
rect 4569 20320 4590 20336
rect 2642 20268 2648 20320
rect 4584 20268 4590 20320
rect 2642 20252 2663 20268
rect 4569 20252 4590 20268
rect 2642 20200 2648 20252
rect 4584 20200 4590 20252
rect 2642 18728 2663 20200
rect 4569 18728 4590 20200
rect 2642 18676 2648 18728
rect 4584 18676 4590 18728
rect 2642 18660 2663 18676
rect 4569 18660 4590 18676
rect 2642 18608 2648 18660
rect 4584 18608 4590 18660
rect 2642 18592 2663 18608
rect 4569 18592 4590 18608
rect 2642 18540 2648 18592
rect 2700 18540 2713 18563
rect 2765 18540 2778 18563
rect 2830 18540 2843 18563
rect 2895 18540 2908 18563
rect 2960 18540 2973 18563
rect 3025 18540 3038 18563
rect 3090 18540 3103 18563
rect 3155 18540 3168 18563
rect 3220 18540 3233 18563
rect 3285 18540 3298 18563
rect 3350 18540 3363 18563
rect 3415 18540 3428 18563
rect 3480 18540 3493 18563
rect 3545 18540 3558 18563
rect 3610 18540 3623 18563
rect 3675 18540 3688 18563
rect 3740 18540 3753 18563
rect 3805 18540 3818 18563
rect 3870 18540 3883 18563
rect 3935 18540 3948 18563
rect 4000 18540 4013 18563
rect 4065 18540 4078 18563
rect 4130 18540 4143 18563
rect 4195 18540 4208 18563
rect 4260 18540 4273 18563
rect 4325 18540 4338 18563
rect 4390 18540 4403 18563
rect 4455 18540 4468 18563
rect 4520 18540 4532 18563
rect 4584 18540 4590 18592
rect 2642 18524 4590 18540
rect 2642 18472 2648 18524
rect 2700 18472 2713 18524
rect 2769 18490 2778 18524
rect 2841 18490 2843 18524
rect 3090 18490 3095 18524
rect 3155 18490 3167 18524
rect 2765 18472 2778 18490
rect 2830 18472 2843 18490
rect 2895 18472 2908 18490
rect 2960 18472 2973 18490
rect 3025 18472 3038 18490
rect 3090 18472 3103 18490
rect 3155 18472 3168 18490
rect 3220 18472 3233 18524
rect 3285 18472 3298 18524
rect 3350 18472 3363 18524
rect 3417 18490 3428 18524
rect 3489 18490 3493 18524
rect 3740 18490 3743 18524
rect 3805 18490 3815 18524
rect 3415 18472 3428 18490
rect 3480 18472 3493 18490
rect 3545 18472 3558 18490
rect 3610 18472 3623 18490
rect 3675 18472 3688 18490
rect 3740 18472 3753 18490
rect 3805 18472 3818 18490
rect 3870 18472 3883 18524
rect 3935 18472 3948 18524
rect 4000 18472 4013 18524
rect 4065 18472 4078 18524
rect 4137 18490 4143 18524
rect 4390 18490 4391 18524
rect 4455 18490 4463 18524
rect 4130 18472 4143 18490
rect 4195 18472 4208 18490
rect 4260 18472 4273 18490
rect 4325 18472 4338 18490
rect 4390 18472 4403 18490
rect 4455 18472 4468 18490
rect 4520 18472 4532 18524
rect 4584 18472 4590 18524
rect 2642 18456 4590 18472
rect 2642 18404 2648 18456
rect 2700 18404 2713 18456
rect 2765 18451 2778 18456
rect 2830 18451 2843 18456
rect 2895 18451 2908 18456
rect 2960 18451 2973 18456
rect 3025 18451 3038 18456
rect 3090 18451 3103 18456
rect 3155 18451 3168 18456
rect 2769 18417 2778 18451
rect 2841 18417 2843 18451
rect 3090 18417 3095 18451
rect 3155 18417 3167 18451
rect 2765 18404 2778 18417
rect 2830 18404 2843 18417
rect 2895 18404 2908 18417
rect 2960 18404 2973 18417
rect 3025 18404 3038 18417
rect 3090 18404 3103 18417
rect 3155 18404 3168 18417
rect 3220 18404 3233 18456
rect 3285 18404 3298 18456
rect 3350 18404 3363 18456
rect 3415 18451 3428 18456
rect 3480 18451 3493 18456
rect 3545 18451 3558 18456
rect 3610 18451 3623 18456
rect 3675 18451 3688 18456
rect 3740 18451 3753 18456
rect 3805 18451 3818 18456
rect 3417 18417 3428 18451
rect 3489 18417 3493 18451
rect 3740 18417 3743 18451
rect 3805 18417 3815 18451
rect 3415 18404 3428 18417
rect 3480 18404 3493 18417
rect 3545 18404 3558 18417
rect 3610 18404 3623 18417
rect 3675 18404 3688 18417
rect 3740 18404 3753 18417
rect 3805 18404 3818 18417
rect 3870 18404 3883 18456
rect 3935 18404 3948 18456
rect 4000 18404 4013 18456
rect 4065 18404 4078 18456
rect 4130 18451 4143 18456
rect 4195 18451 4208 18456
rect 4260 18451 4273 18456
rect 4325 18451 4338 18456
rect 4390 18451 4403 18456
rect 4455 18451 4468 18456
rect 4137 18417 4143 18451
rect 4390 18417 4391 18451
rect 4455 18417 4463 18451
rect 4130 18404 4143 18417
rect 4195 18404 4208 18417
rect 4260 18404 4273 18417
rect 4325 18404 4338 18417
rect 4390 18404 4403 18417
rect 4455 18404 4468 18417
rect 4520 18404 4532 18456
rect 4584 18404 4590 18456
rect 2642 18388 4590 18404
rect 2642 18336 2648 18388
rect 2700 18336 2713 18388
rect 2765 18378 2778 18388
rect 2830 18378 2843 18388
rect 2895 18378 2908 18388
rect 2960 18378 2973 18388
rect 3025 18378 3038 18388
rect 3090 18378 3103 18388
rect 3155 18378 3168 18388
rect 2769 18344 2778 18378
rect 2841 18344 2843 18378
rect 3090 18344 3095 18378
rect 3155 18344 3167 18378
rect 2765 18336 2778 18344
rect 2830 18336 2843 18344
rect 2895 18336 2908 18344
rect 2960 18336 2973 18344
rect 3025 18336 3038 18344
rect 3090 18336 3103 18344
rect 3155 18336 3168 18344
rect 3220 18336 3233 18388
rect 3285 18336 3298 18388
rect 3350 18336 3363 18388
rect 3415 18378 3428 18388
rect 3480 18378 3493 18388
rect 3545 18378 3558 18388
rect 3610 18378 3623 18388
rect 3675 18378 3688 18388
rect 3740 18378 3753 18388
rect 3805 18378 3818 18388
rect 3417 18344 3428 18378
rect 3489 18344 3493 18378
rect 3740 18344 3743 18378
rect 3805 18344 3815 18378
rect 3415 18336 3428 18344
rect 3480 18336 3493 18344
rect 3545 18336 3558 18344
rect 3610 18336 3623 18344
rect 3675 18336 3688 18344
rect 3740 18336 3753 18344
rect 3805 18336 3818 18344
rect 3870 18336 3883 18388
rect 3935 18336 3948 18388
rect 4000 18336 4013 18388
rect 4065 18336 4078 18388
rect 4130 18378 4143 18388
rect 4195 18378 4208 18388
rect 4260 18378 4273 18388
rect 4325 18378 4338 18388
rect 4390 18378 4403 18388
rect 4455 18378 4468 18388
rect 4137 18344 4143 18378
rect 4390 18344 4391 18378
rect 4455 18344 4463 18378
rect 4130 18336 4143 18344
rect 4195 18336 4208 18344
rect 4260 18336 4273 18344
rect 4325 18336 4338 18344
rect 4390 18336 4403 18344
rect 4455 18336 4468 18344
rect 4520 18336 4532 18388
rect 4584 18336 4590 18388
rect 2642 18320 4590 18336
rect 2642 18268 2648 18320
rect 2700 18268 2713 18320
rect 2765 18305 2778 18320
rect 2830 18305 2843 18320
rect 2895 18305 2908 18320
rect 2960 18305 2973 18320
rect 3025 18305 3038 18320
rect 3090 18305 3103 18320
rect 3155 18305 3168 18320
rect 2769 18271 2778 18305
rect 2841 18271 2843 18305
rect 3090 18271 3095 18305
rect 3155 18271 3167 18305
rect 2765 18268 2778 18271
rect 2830 18268 2843 18271
rect 2895 18268 2908 18271
rect 2960 18268 2973 18271
rect 3025 18268 3038 18271
rect 3090 18268 3103 18271
rect 3155 18268 3168 18271
rect 3220 18268 3233 18320
rect 3285 18268 3298 18320
rect 3350 18268 3363 18320
rect 3415 18305 3428 18320
rect 3480 18305 3493 18320
rect 3545 18305 3558 18320
rect 3610 18305 3623 18320
rect 3675 18305 3688 18320
rect 3740 18305 3753 18320
rect 3805 18305 3818 18320
rect 3417 18271 3428 18305
rect 3489 18271 3493 18305
rect 3740 18271 3743 18305
rect 3805 18271 3815 18305
rect 3415 18268 3428 18271
rect 3480 18268 3493 18271
rect 3545 18268 3558 18271
rect 3610 18268 3623 18271
rect 3675 18268 3688 18271
rect 3740 18268 3753 18271
rect 3805 18268 3818 18271
rect 3870 18268 3883 18320
rect 3935 18268 3948 18320
rect 4000 18268 4013 18320
rect 4065 18268 4078 18320
rect 4130 18305 4143 18320
rect 4195 18305 4208 18320
rect 4260 18305 4273 18320
rect 4325 18305 4338 18320
rect 4390 18305 4403 18320
rect 4455 18305 4468 18320
rect 4137 18271 4143 18305
rect 4390 18271 4391 18305
rect 4455 18271 4463 18305
rect 4130 18268 4143 18271
rect 4195 18268 4208 18271
rect 4260 18268 4273 18271
rect 4325 18268 4338 18271
rect 4390 18268 4403 18271
rect 4455 18268 4468 18271
rect 4520 18268 4532 18320
rect 4584 18268 4590 18320
rect 2642 18252 4590 18268
rect 2642 18200 2648 18252
rect 2700 18200 2713 18252
rect 2765 18232 2778 18252
rect 2830 18232 2843 18252
rect 2895 18232 2908 18252
rect 2960 18232 2973 18252
rect 3025 18232 3038 18252
rect 3090 18232 3103 18252
rect 3155 18232 3168 18252
rect 2769 18200 2778 18232
rect 2841 18200 2843 18232
rect 3090 18200 3095 18232
rect 3155 18200 3167 18232
rect 3220 18200 3233 18252
rect 3285 18200 3298 18252
rect 3350 18200 3363 18252
rect 3415 18232 3428 18252
rect 3480 18232 3493 18252
rect 3545 18232 3558 18252
rect 3610 18232 3623 18252
rect 3675 18232 3688 18252
rect 3740 18232 3753 18252
rect 3805 18232 3818 18252
rect 3417 18200 3428 18232
rect 3489 18200 3493 18232
rect 3740 18200 3743 18232
rect 3805 18200 3815 18232
rect 3870 18200 3883 18252
rect 3935 18200 3948 18252
rect 4000 18200 4013 18252
rect 4065 18200 4078 18252
rect 4130 18232 4143 18252
rect 4195 18232 4208 18252
rect 4260 18232 4273 18252
rect 4325 18232 4338 18252
rect 4390 18232 4403 18252
rect 4455 18232 4468 18252
rect 4137 18200 4143 18232
rect 4390 18200 4391 18232
rect 4455 18200 4463 18232
rect 4520 18200 4532 18252
rect 4584 18200 4590 18252
rect 2642 18198 2663 18200
rect 2697 18198 2735 18200
rect 2769 18198 2807 18200
rect 2841 18198 2879 18200
rect 2913 18198 2951 18200
rect 2985 18198 3023 18200
rect 3057 18198 3095 18200
rect 3129 18198 3167 18200
rect 3201 18198 3239 18200
rect 3273 18198 3311 18200
rect 3345 18198 3383 18200
rect 3417 18198 3455 18200
rect 3489 18198 3527 18200
rect 3561 18198 3599 18200
rect 3633 18198 3671 18200
rect 3705 18198 3743 18200
rect 3777 18198 3815 18200
rect 3849 18198 3887 18200
rect 3921 18198 3959 18200
rect 3993 18198 4031 18200
rect 4065 18198 4103 18200
rect 4137 18198 4175 18200
rect 4209 18198 4247 18200
rect 4281 18198 4319 18200
rect 4353 18198 4391 18200
rect 4425 18198 4463 18200
rect 4497 18198 4535 18200
rect 4569 18198 4590 18200
rect 2642 18159 4590 18198
rect 2642 18125 2663 18159
rect 2697 18125 2735 18159
rect 2769 18125 2807 18159
rect 2841 18125 2879 18159
rect 2913 18125 2951 18159
rect 2985 18125 3023 18159
rect 3057 18125 3095 18159
rect 3129 18125 3167 18159
rect 3201 18125 3239 18159
rect 3273 18125 3311 18159
rect 3345 18125 3383 18159
rect 3417 18125 3455 18159
rect 3489 18125 3527 18159
rect 3561 18125 3599 18159
rect 3633 18125 3671 18159
rect 3705 18125 3743 18159
rect 3777 18125 3815 18159
rect 3849 18125 3887 18159
rect 3921 18125 3959 18159
rect 3993 18125 4031 18159
rect 4065 18125 4103 18159
rect 4137 18125 4175 18159
rect 4209 18125 4247 18159
rect 4281 18125 4319 18159
rect 4353 18125 4391 18159
rect 4425 18125 4463 18159
rect 4497 18125 4535 18159
rect 4569 18125 4590 18159
rect 2642 18086 4590 18125
rect 2642 18052 2663 18086
rect 2697 18052 2735 18086
rect 2769 18052 2807 18086
rect 2841 18052 2879 18086
rect 2913 18052 2951 18086
rect 2985 18052 3023 18086
rect 3057 18052 3095 18086
rect 3129 18052 3167 18086
rect 3201 18052 3239 18086
rect 3273 18052 3311 18086
rect 3345 18052 3383 18086
rect 3417 18052 3455 18086
rect 3489 18052 3527 18086
rect 3561 18052 3599 18086
rect 3633 18052 3671 18086
rect 3705 18052 3743 18086
rect 3777 18052 3815 18086
rect 3849 18052 3887 18086
rect 3921 18052 3959 18086
rect 3993 18052 4031 18086
rect 4065 18052 4103 18086
rect 4137 18052 4175 18086
rect 4209 18052 4247 18086
rect 4281 18052 4319 18086
rect 4353 18052 4391 18086
rect 4425 18052 4463 18086
rect 4497 18052 4535 18086
rect 4569 18052 4590 18086
rect 2642 18013 4590 18052
rect 2642 17979 2663 18013
rect 2697 17979 2735 18013
rect 2769 17979 2807 18013
rect 2841 17979 2879 18013
rect 2913 17979 2951 18013
rect 2985 17979 3023 18013
rect 3057 17979 3095 18013
rect 3129 17979 3167 18013
rect 3201 17979 3239 18013
rect 3273 17979 3311 18013
rect 3345 17979 3383 18013
rect 3417 17979 3455 18013
rect 3489 17979 3527 18013
rect 3561 17979 3599 18013
rect 3633 17979 3671 18013
rect 3705 17979 3743 18013
rect 3777 17979 3815 18013
rect 3849 17979 3887 18013
rect 3921 17979 3959 18013
rect 3993 17979 4031 18013
rect 4065 17979 4103 18013
rect 4137 17979 4175 18013
rect 4209 17979 4247 18013
rect 4281 17979 4319 18013
rect 4353 17979 4391 18013
rect 4425 17979 4463 18013
rect 4497 17979 4535 18013
rect 4569 17979 4590 18013
rect 2642 17940 4590 17979
rect 2642 17906 2663 17940
rect 2697 17906 2735 17940
rect 2769 17906 2807 17940
rect 2841 17906 2879 17940
rect 2913 17906 2951 17940
rect 2985 17906 3023 17940
rect 3057 17906 3095 17940
rect 3129 17906 3167 17940
rect 3201 17906 3239 17940
rect 3273 17906 3311 17940
rect 3345 17906 3383 17940
rect 3417 17906 3455 17940
rect 3489 17906 3527 17940
rect 3561 17906 3599 17940
rect 3633 17906 3671 17940
rect 3705 17906 3743 17940
rect 3777 17906 3815 17940
rect 3849 17906 3887 17940
rect 3921 17906 3959 17940
rect 3993 17906 4031 17940
rect 4065 17906 4103 17940
rect 4137 17906 4175 17940
rect 4209 17906 4247 17940
rect 4281 17906 4319 17940
rect 4353 17906 4391 17940
rect 4425 17906 4463 17940
rect 4497 17906 4535 17940
rect 4569 17906 4590 17940
rect 2642 17867 4590 17906
rect 2642 17833 2663 17867
rect 2697 17833 2735 17867
rect 2769 17833 2807 17867
rect 2841 17833 2879 17867
rect 2913 17833 2951 17867
rect 2985 17833 3023 17867
rect 3057 17833 3095 17867
rect 3129 17833 3167 17867
rect 3201 17833 3239 17867
rect 3273 17833 3311 17867
rect 3345 17833 3383 17867
rect 3417 17833 3455 17867
rect 3489 17833 3527 17867
rect 3561 17833 3599 17867
rect 3633 17833 3671 17867
rect 3705 17833 3743 17867
rect 3777 17833 3815 17867
rect 3849 17833 3887 17867
rect 3921 17833 3959 17867
rect 3993 17833 4031 17867
rect 4065 17833 4103 17867
rect 4137 17833 4175 17867
rect 4209 17833 4247 17867
rect 4281 17833 4319 17867
rect 4353 17833 4391 17867
rect 4425 17833 4463 17867
rect 4497 17833 4535 17867
rect 4569 17833 4590 17867
rect 2642 17794 4590 17833
rect 2642 17760 2663 17794
rect 2697 17760 2735 17794
rect 2769 17760 2807 17794
rect 2841 17760 2879 17794
rect 2913 17760 2951 17794
rect 2985 17760 3023 17794
rect 3057 17760 3095 17794
rect 3129 17760 3167 17794
rect 3201 17760 3239 17794
rect 3273 17760 3311 17794
rect 3345 17760 3383 17794
rect 3417 17760 3455 17794
rect 3489 17760 3527 17794
rect 3561 17760 3599 17794
rect 3633 17760 3671 17794
rect 3705 17760 3743 17794
rect 3777 17760 3815 17794
rect 3849 17760 3887 17794
rect 3921 17760 3959 17794
rect 3993 17760 4031 17794
rect 4065 17760 4103 17794
rect 4137 17760 4175 17794
rect 4209 17760 4247 17794
rect 4281 17760 4319 17794
rect 4353 17760 4391 17794
rect 4425 17760 4463 17794
rect 4497 17760 4535 17794
rect 4569 17760 4590 17794
rect 2642 17721 4590 17760
rect 2642 17687 2663 17721
rect 2697 17687 2735 17721
rect 2769 17687 2807 17721
rect 2841 17687 2879 17721
rect 2913 17687 2951 17721
rect 2985 17687 3023 17721
rect 3057 17687 3095 17721
rect 3129 17687 3167 17721
rect 3201 17687 3239 17721
rect 3273 17687 3311 17721
rect 3345 17687 3383 17721
rect 3417 17687 3455 17721
rect 3489 17687 3527 17721
rect 3561 17687 3599 17721
rect 3633 17687 3671 17721
rect 3705 17687 3743 17721
rect 3777 17687 3815 17721
rect 3849 17687 3887 17721
rect 3921 17687 3959 17721
rect 3993 17687 4031 17721
rect 4065 17687 4103 17721
rect 4137 17687 4175 17721
rect 4209 17687 4247 17721
rect 4281 17687 4319 17721
rect 4353 17687 4391 17721
rect 4425 17687 4463 17721
rect 4497 17687 4535 17721
rect 4569 17687 4590 17721
rect 2642 17648 4590 17687
rect 2642 17614 2663 17648
rect 2697 17614 2735 17648
rect 2769 17614 2807 17648
rect 2841 17614 2879 17648
rect 2913 17614 2951 17648
rect 2985 17614 3023 17648
rect 3057 17614 3095 17648
rect 3129 17614 3167 17648
rect 3201 17614 3239 17648
rect 3273 17614 3311 17648
rect 3345 17614 3383 17648
rect 3417 17614 3455 17648
rect 3489 17614 3527 17648
rect 3561 17614 3599 17648
rect 3633 17614 3671 17648
rect 3705 17614 3743 17648
rect 3777 17614 3815 17648
rect 3849 17614 3887 17648
rect 3921 17614 3959 17648
rect 3993 17614 4031 17648
rect 4065 17614 4103 17648
rect 4137 17614 4175 17648
rect 4209 17614 4247 17648
rect 4281 17614 4319 17648
rect 4353 17614 4391 17648
rect 4425 17614 4463 17648
rect 4497 17614 4535 17648
rect 4569 17614 4590 17648
rect 2642 17575 4590 17614
rect 2642 17541 2663 17575
rect 2697 17541 2735 17575
rect 2769 17541 2807 17575
rect 2841 17541 2879 17575
rect 2913 17541 2951 17575
rect 2985 17541 3023 17575
rect 3057 17541 3095 17575
rect 3129 17541 3167 17575
rect 3201 17541 3239 17575
rect 3273 17541 3311 17575
rect 3345 17541 3383 17575
rect 3417 17541 3455 17575
rect 3489 17541 3527 17575
rect 3561 17541 3599 17575
rect 3633 17541 3671 17575
rect 3705 17541 3743 17575
rect 3777 17541 3815 17575
rect 3849 17541 3887 17575
rect 3921 17541 3959 17575
rect 3993 17541 4031 17575
rect 4065 17541 4103 17575
rect 4137 17541 4175 17575
rect 4209 17541 4247 17575
rect 4281 17541 4319 17575
rect 4353 17541 4391 17575
rect 4425 17541 4463 17575
rect 4497 17541 4535 17575
rect 4569 17541 4590 17575
rect 2642 17502 4590 17541
rect 2642 17468 2663 17502
rect 2697 17468 2735 17502
rect 2769 17468 2807 17502
rect 2841 17468 2879 17502
rect 2913 17468 2951 17502
rect 2985 17468 3023 17502
rect 3057 17468 3095 17502
rect 3129 17468 3167 17502
rect 3201 17468 3239 17502
rect 3273 17468 3311 17502
rect 3345 17468 3383 17502
rect 3417 17468 3455 17502
rect 3489 17468 3527 17502
rect 3561 17468 3599 17502
rect 3633 17468 3671 17502
rect 3705 17468 3743 17502
rect 3777 17468 3815 17502
rect 3849 17468 3887 17502
rect 3921 17468 3959 17502
rect 3993 17468 4031 17502
rect 4065 17468 4103 17502
rect 4137 17468 4175 17502
rect 4209 17468 4247 17502
rect 4281 17468 4319 17502
rect 4353 17468 4391 17502
rect 4425 17468 4463 17502
rect 4497 17468 4535 17502
rect 4569 17468 4590 17502
rect 2642 17429 4590 17468
rect 2642 17395 2663 17429
rect 2697 17395 2735 17429
rect 2769 17395 2807 17429
rect 2841 17395 2879 17429
rect 2913 17395 2951 17429
rect 2985 17395 3023 17429
rect 3057 17395 3095 17429
rect 3129 17395 3167 17429
rect 3201 17395 3239 17429
rect 3273 17395 3311 17429
rect 3345 17395 3383 17429
rect 3417 17395 3455 17429
rect 3489 17395 3527 17429
rect 3561 17395 3599 17429
rect 3633 17395 3671 17429
rect 3705 17395 3743 17429
rect 3777 17395 3815 17429
rect 3849 17395 3887 17429
rect 3921 17395 3959 17429
rect 3993 17395 4031 17429
rect 4065 17395 4103 17429
rect 4137 17395 4175 17429
rect 4209 17395 4247 17429
rect 4281 17395 4319 17429
rect 4353 17395 4391 17429
rect 4425 17395 4463 17429
rect 4497 17395 4535 17429
rect 4569 17395 4590 17429
rect 2642 17356 4590 17395
rect 2642 17322 2663 17356
rect 2697 17322 2735 17356
rect 2769 17322 2807 17356
rect 2841 17322 2879 17356
rect 2913 17322 2951 17356
rect 2985 17322 3023 17356
rect 3057 17322 3095 17356
rect 3129 17322 3167 17356
rect 3201 17322 3239 17356
rect 3273 17322 3311 17356
rect 3345 17322 3383 17356
rect 3417 17322 3455 17356
rect 3489 17322 3527 17356
rect 3561 17322 3599 17356
rect 3633 17322 3671 17356
rect 3705 17322 3743 17356
rect 3777 17322 3815 17356
rect 3849 17322 3887 17356
rect 3921 17322 3959 17356
rect 3993 17322 4031 17356
rect 4065 17322 4103 17356
rect 4137 17322 4175 17356
rect 4209 17322 4247 17356
rect 4281 17322 4319 17356
rect 4353 17322 4391 17356
rect 4425 17322 4463 17356
rect 4497 17322 4535 17356
rect 4569 17322 4590 17356
rect 2642 17283 4590 17322
rect 2642 17249 2663 17283
rect 2697 17249 2735 17283
rect 2769 17249 2807 17283
rect 2841 17249 2879 17283
rect 2913 17249 2951 17283
rect 2985 17249 3023 17283
rect 3057 17249 3095 17283
rect 3129 17249 3167 17283
rect 3201 17249 3239 17283
rect 3273 17249 3311 17283
rect 3345 17249 3383 17283
rect 3417 17249 3455 17283
rect 3489 17249 3527 17283
rect 3561 17249 3599 17283
rect 3633 17249 3671 17283
rect 3705 17249 3743 17283
rect 3777 17249 3815 17283
rect 3849 17249 3887 17283
rect 3921 17249 3959 17283
rect 3993 17249 4031 17283
rect 4065 17249 4103 17283
rect 4137 17249 4175 17283
rect 4209 17249 4247 17283
rect 4281 17249 4319 17283
rect 4353 17249 4391 17283
rect 4425 17249 4463 17283
rect 4497 17249 4535 17283
rect 4569 17249 4590 17283
rect 2642 17210 4590 17249
rect 2642 17176 2663 17210
rect 2697 17176 2735 17210
rect 2769 17176 2807 17210
rect 2841 17176 2879 17210
rect 2913 17176 2951 17210
rect 2985 17176 3023 17210
rect 3057 17176 3095 17210
rect 3129 17176 3167 17210
rect 3201 17176 3239 17210
rect 3273 17176 3311 17210
rect 3345 17176 3383 17210
rect 3417 17176 3455 17210
rect 3489 17176 3527 17210
rect 3561 17176 3599 17210
rect 3633 17176 3671 17210
rect 3705 17176 3743 17210
rect 3777 17176 3815 17210
rect 3849 17176 3887 17210
rect 3921 17176 3959 17210
rect 3993 17176 4031 17210
rect 4065 17176 4103 17210
rect 4137 17176 4175 17210
rect 4209 17176 4247 17210
rect 4281 17176 4319 17210
rect 4353 17176 4391 17210
rect 4425 17176 4463 17210
rect 4497 17176 4535 17210
rect 4569 17176 4590 17210
rect 2642 17137 4590 17176
rect 2642 17103 2663 17137
rect 2697 17103 2735 17137
rect 2769 17103 2807 17137
rect 2841 17103 2879 17137
rect 2913 17103 2951 17137
rect 2985 17103 3023 17137
rect 3057 17103 3095 17137
rect 3129 17103 3167 17137
rect 3201 17103 3239 17137
rect 3273 17103 3311 17137
rect 3345 17103 3383 17137
rect 3417 17103 3455 17137
rect 3489 17103 3527 17137
rect 3561 17103 3599 17137
rect 3633 17103 3671 17137
rect 3705 17103 3743 17137
rect 3777 17103 3815 17137
rect 3849 17103 3887 17137
rect 3921 17103 3959 17137
rect 3993 17103 4031 17137
rect 4065 17103 4103 17137
rect 4137 17103 4175 17137
rect 4209 17103 4247 17137
rect 4281 17103 4319 17137
rect 4353 17103 4391 17137
rect 4425 17103 4463 17137
rect 4497 17103 4535 17137
rect 4569 17103 4590 17137
rect 2642 17064 4590 17103
rect 2642 17030 2663 17064
rect 2697 17030 2735 17064
rect 2769 17030 2807 17064
rect 2841 17030 2879 17064
rect 2913 17030 2951 17064
rect 2985 17030 3023 17064
rect 3057 17030 3095 17064
rect 3129 17030 3167 17064
rect 3201 17030 3239 17064
rect 3273 17030 3311 17064
rect 3345 17030 3383 17064
rect 3417 17030 3455 17064
rect 3489 17030 3527 17064
rect 3561 17030 3599 17064
rect 3633 17030 3671 17064
rect 3705 17030 3743 17064
rect 3777 17030 3815 17064
rect 3849 17030 3887 17064
rect 3921 17030 3959 17064
rect 3993 17030 4031 17064
rect 4065 17030 4103 17064
rect 4137 17030 4175 17064
rect 4209 17030 4247 17064
rect 4281 17030 4319 17064
rect 4353 17030 4391 17064
rect 4425 17030 4463 17064
rect 4497 17030 4535 17064
rect 4569 17030 4590 17064
rect 2642 16991 4590 17030
rect 2642 16957 2663 16991
rect 2697 16957 2735 16991
rect 2769 16970 2807 16991
rect 2841 16970 2879 16991
rect 2913 16970 2951 16991
rect 2985 16970 3023 16991
rect 3057 16970 3095 16991
rect 3129 16970 3167 16991
rect 3201 16970 3239 16991
rect 3273 16970 3311 16991
rect 3345 16970 3383 16991
rect 3417 16970 3455 16991
rect 3489 16970 3527 16991
rect 3561 16970 3599 16991
rect 3633 16970 3671 16991
rect 3705 16970 3743 16991
rect 3777 16970 3815 16991
rect 3849 16970 3887 16991
rect 3921 16970 3959 16991
rect 3993 16970 4031 16991
rect 4065 16970 4103 16991
rect 4137 16970 4175 16991
rect 4209 16970 4247 16991
rect 4281 16970 4319 16991
rect 4353 16970 4391 16991
rect 4425 16970 4463 16991
rect 4497 16970 4535 16991
rect 2798 16957 2807 16970
rect 2865 16957 2879 16970
rect 2642 16918 2746 16957
rect 2798 16918 2813 16957
rect 2865 16918 2880 16957
rect 2932 16918 2946 16970
rect 2998 16918 3012 16970
rect 3064 16918 3078 16970
rect 3130 16918 3144 16970
rect 3201 16957 3210 16970
rect 3273 16957 3276 16970
rect 3526 16957 3527 16970
rect 3592 16957 3599 16970
rect 3658 16957 3671 16970
rect 3196 16918 3210 16957
rect 3262 16918 3276 16957
rect 3328 16918 3342 16957
rect 3394 16918 3408 16957
rect 3460 16918 3474 16957
rect 3526 16918 3540 16957
rect 3592 16918 3606 16957
rect 3658 16918 3672 16957
rect 3724 16918 3738 16970
rect 3790 16918 3804 16970
rect 3856 16918 3870 16970
rect 3922 16918 3936 16970
rect 3993 16957 4002 16970
rect 4065 16957 4068 16970
rect 4318 16957 4319 16970
rect 4384 16957 4391 16970
rect 4450 16957 4463 16970
rect 4516 16957 4535 16970
rect 4569 16957 4590 16991
rect 3988 16918 4002 16957
rect 4054 16918 4068 16957
rect 4120 16918 4134 16957
rect 4186 16918 4200 16957
rect 4252 16918 4266 16957
rect 4318 16918 4332 16957
rect 4384 16918 4398 16957
rect 4450 16918 4464 16957
rect 4516 16918 4590 16957
rect 2642 16884 2663 16918
rect 2697 16884 2735 16918
rect 2769 16904 2807 16918
rect 2841 16904 2879 16918
rect 2913 16904 2951 16918
rect 2985 16904 3023 16918
rect 3057 16904 3095 16918
rect 3129 16904 3167 16918
rect 3201 16904 3239 16918
rect 3273 16904 3311 16918
rect 3345 16904 3383 16918
rect 3417 16904 3455 16918
rect 3489 16904 3527 16918
rect 3561 16904 3599 16918
rect 3633 16904 3671 16918
rect 3705 16904 3743 16918
rect 3777 16904 3815 16918
rect 3849 16904 3887 16918
rect 3921 16904 3959 16918
rect 3993 16904 4031 16918
rect 4065 16904 4103 16918
rect 4137 16904 4175 16918
rect 4209 16904 4247 16918
rect 4281 16904 4319 16918
rect 4353 16904 4391 16918
rect 4425 16904 4463 16918
rect 4497 16904 4535 16918
rect 2798 16884 2807 16904
rect 2865 16884 2879 16904
rect 2642 16852 2746 16884
rect 2798 16852 2813 16884
rect 2865 16852 2880 16884
rect 2932 16852 2946 16904
rect 2998 16852 3012 16904
rect 3064 16852 3078 16904
rect 3130 16852 3144 16904
rect 3201 16884 3210 16904
rect 3273 16884 3276 16904
rect 3526 16884 3527 16904
rect 3592 16884 3599 16904
rect 3658 16884 3671 16904
rect 3196 16852 3210 16884
rect 3262 16852 3276 16884
rect 3328 16852 3342 16884
rect 3394 16852 3408 16884
rect 3460 16852 3474 16884
rect 3526 16852 3540 16884
rect 3592 16852 3606 16884
rect 3658 16852 3672 16884
rect 3724 16852 3738 16904
rect 3790 16852 3804 16904
rect 3856 16852 3870 16904
rect 3922 16852 3936 16904
rect 3993 16884 4002 16904
rect 4065 16884 4068 16904
rect 4318 16884 4319 16904
rect 4384 16884 4391 16904
rect 4450 16884 4463 16904
rect 4516 16884 4535 16904
rect 4569 16884 4590 16918
rect 3988 16852 4002 16884
rect 4054 16852 4068 16884
rect 4120 16852 4134 16884
rect 4186 16852 4200 16884
rect 4252 16852 4266 16884
rect 4318 16852 4332 16884
rect 4384 16852 4398 16884
rect 4450 16852 4464 16884
rect 4516 16852 4590 16884
rect 2642 16845 4590 16852
rect 2642 16811 2663 16845
rect 2697 16811 2735 16845
rect 2769 16838 2807 16845
rect 2841 16838 2879 16845
rect 2913 16838 2951 16845
rect 2985 16838 3023 16845
rect 3057 16838 3095 16845
rect 3129 16838 3167 16845
rect 3201 16838 3239 16845
rect 3273 16838 3311 16845
rect 3345 16838 3383 16845
rect 3417 16838 3455 16845
rect 3489 16838 3527 16845
rect 3561 16838 3599 16845
rect 3633 16838 3671 16845
rect 3705 16838 3743 16845
rect 3777 16838 3815 16845
rect 3849 16838 3887 16845
rect 3921 16838 3959 16845
rect 3993 16838 4031 16845
rect 4065 16838 4103 16845
rect 4137 16838 4175 16845
rect 4209 16838 4247 16845
rect 4281 16838 4319 16845
rect 4353 16838 4391 16845
rect 4425 16838 4463 16845
rect 4497 16838 4535 16845
rect 2798 16811 2807 16838
rect 2865 16811 2879 16838
rect 2642 16786 2746 16811
rect 2798 16786 2813 16811
rect 2865 16786 2880 16811
rect 2932 16786 2946 16838
rect 2998 16786 3012 16838
rect 3064 16786 3078 16838
rect 3130 16786 3144 16838
rect 3201 16811 3210 16838
rect 3273 16811 3276 16838
rect 3526 16811 3527 16838
rect 3592 16811 3599 16838
rect 3658 16811 3671 16838
rect 3196 16786 3210 16811
rect 3262 16786 3276 16811
rect 3328 16786 3342 16811
rect 3394 16786 3408 16811
rect 3460 16786 3474 16811
rect 3526 16786 3540 16811
rect 3592 16786 3606 16811
rect 3658 16786 3672 16811
rect 3724 16786 3738 16838
rect 3790 16786 3804 16838
rect 3856 16786 3870 16838
rect 3922 16786 3936 16838
rect 3993 16811 4002 16838
rect 4065 16811 4068 16838
rect 4318 16811 4319 16838
rect 4384 16811 4391 16838
rect 4450 16811 4463 16838
rect 4516 16811 4535 16838
rect 4569 16811 4590 16845
rect 3988 16786 4002 16811
rect 4054 16786 4068 16811
rect 4120 16786 4134 16811
rect 4186 16786 4200 16811
rect 4252 16786 4266 16811
rect 4318 16786 4332 16811
rect 4384 16786 4398 16811
rect 4450 16786 4464 16811
rect 4516 16786 4590 16811
rect 2642 16772 4590 16786
rect 2642 16738 2663 16772
rect 2697 16738 2735 16772
rect 2798 16738 2807 16772
rect 2865 16738 2879 16772
rect 2642 16720 2746 16738
rect 2798 16720 2813 16738
rect 2865 16720 2880 16738
rect 2932 16720 2946 16772
rect 2998 16720 3012 16772
rect 3064 16720 3078 16772
rect 3130 16720 3144 16772
rect 3201 16738 3210 16772
rect 3273 16738 3276 16772
rect 3526 16738 3527 16772
rect 3592 16738 3599 16772
rect 3658 16738 3671 16772
rect 3196 16720 3210 16738
rect 3262 16720 3276 16738
rect 3328 16720 3342 16738
rect 3394 16720 3408 16738
rect 3460 16720 3474 16738
rect 3526 16720 3540 16738
rect 3592 16720 3606 16738
rect 3658 16720 3672 16738
rect 3724 16720 3738 16772
rect 3790 16720 3804 16772
rect 3856 16720 3870 16772
rect 3922 16720 3936 16772
rect 3993 16738 4002 16772
rect 4065 16738 4068 16772
rect 4318 16738 4319 16772
rect 4384 16738 4391 16772
rect 4450 16738 4463 16772
rect 4516 16738 4535 16772
rect 4569 16738 4590 16772
rect 3988 16720 4002 16738
rect 4054 16720 4068 16738
rect 4120 16720 4134 16738
rect 4186 16720 4200 16738
rect 4252 16720 4266 16738
rect 4318 16720 4332 16738
rect 4384 16720 4398 16738
rect 4450 16720 4464 16738
rect 4516 16720 4590 16738
rect 2642 16706 4590 16720
rect 2642 16699 2746 16706
rect 2798 16699 2813 16706
rect 2865 16699 2880 16706
rect 2642 16665 2663 16699
rect 2697 16665 2735 16699
rect 2798 16665 2807 16699
rect 2865 16665 2879 16699
rect 2642 16654 2746 16665
rect 2798 16654 2813 16665
rect 2865 16654 2880 16665
rect 2932 16654 2946 16706
rect 2998 16654 3012 16706
rect 3064 16654 3078 16706
rect 3130 16654 3144 16706
rect 3196 16699 3210 16706
rect 3262 16699 3276 16706
rect 3328 16699 3342 16706
rect 3394 16699 3408 16706
rect 3460 16699 3474 16706
rect 3526 16699 3540 16706
rect 3592 16699 3606 16706
rect 3658 16699 3672 16706
rect 3201 16665 3210 16699
rect 3273 16665 3276 16699
rect 3526 16665 3527 16699
rect 3592 16665 3599 16699
rect 3658 16665 3671 16699
rect 3196 16654 3210 16665
rect 3262 16654 3276 16665
rect 3328 16654 3342 16665
rect 3394 16654 3408 16665
rect 3460 16654 3474 16665
rect 3526 16654 3540 16665
rect 3592 16654 3606 16665
rect 3658 16654 3672 16665
rect 3724 16654 3738 16706
rect 3790 16654 3804 16706
rect 3856 16654 3870 16706
rect 3922 16654 3936 16706
rect 3988 16699 4002 16706
rect 4054 16699 4068 16706
rect 4120 16699 4134 16706
rect 4186 16699 4200 16706
rect 4252 16699 4266 16706
rect 4318 16699 4332 16706
rect 4384 16699 4398 16706
rect 4450 16699 4464 16706
rect 4516 16699 4590 16706
rect 3993 16665 4002 16699
rect 4065 16665 4068 16699
rect 4318 16665 4319 16699
rect 4384 16665 4391 16699
rect 4450 16665 4463 16699
rect 4516 16665 4535 16699
rect 4569 16665 4590 16699
rect 3988 16654 4002 16665
rect 4054 16654 4068 16665
rect 4120 16654 4134 16665
rect 4186 16654 4200 16665
rect 4252 16654 4266 16665
rect 4318 16654 4332 16665
rect 4384 16654 4398 16665
rect 4450 16654 4464 16665
rect 4516 16654 4590 16665
rect 2642 16640 4590 16654
rect 2642 16626 2746 16640
rect 2798 16626 2813 16640
rect 2865 16626 2880 16640
rect 2642 16592 2663 16626
rect 2697 16592 2735 16626
rect 2798 16592 2807 16626
rect 2865 16592 2879 16626
rect 2642 16588 2746 16592
rect 2798 16588 2813 16592
rect 2865 16588 2880 16592
rect 2932 16588 2946 16640
rect 2998 16588 3012 16640
rect 3064 16588 3078 16640
rect 3130 16588 3144 16640
rect 3196 16626 3210 16640
rect 3262 16626 3276 16640
rect 3328 16626 3342 16640
rect 3394 16626 3408 16640
rect 3460 16626 3474 16640
rect 3526 16626 3540 16640
rect 3592 16626 3606 16640
rect 3658 16626 3672 16640
rect 3201 16592 3210 16626
rect 3273 16592 3276 16626
rect 3526 16592 3527 16626
rect 3592 16592 3599 16626
rect 3658 16592 3671 16626
rect 3196 16588 3210 16592
rect 3262 16588 3276 16592
rect 3328 16588 3342 16592
rect 3394 16588 3408 16592
rect 3460 16588 3474 16592
rect 3526 16588 3540 16592
rect 3592 16588 3606 16592
rect 3658 16588 3672 16592
rect 3724 16588 3738 16640
rect 3790 16588 3804 16640
rect 3856 16588 3870 16640
rect 3922 16588 3936 16640
rect 3988 16626 4002 16640
rect 4054 16626 4068 16640
rect 4120 16626 4134 16640
rect 4186 16626 4200 16640
rect 4252 16626 4266 16640
rect 4318 16626 4332 16640
rect 4384 16626 4398 16640
rect 4450 16626 4464 16640
rect 4516 16626 4590 16640
rect 3993 16592 4002 16626
rect 4065 16592 4068 16626
rect 4318 16592 4319 16626
rect 4384 16592 4391 16626
rect 4450 16592 4463 16626
rect 4516 16592 4535 16626
rect 4569 16592 4590 16626
rect 3988 16588 4002 16592
rect 4054 16588 4068 16592
rect 4120 16588 4134 16592
rect 4186 16588 4200 16592
rect 4252 16588 4266 16592
rect 4318 16588 4332 16592
rect 4384 16588 4398 16592
rect 4450 16588 4464 16592
rect 4516 16588 4590 16592
rect 2642 16574 4590 16588
rect 2642 16553 2746 16574
rect 2798 16553 2813 16574
rect 2865 16553 2880 16574
rect 2642 16519 2663 16553
rect 2697 16519 2735 16553
rect 2798 16522 2807 16553
rect 2865 16522 2879 16553
rect 2932 16522 2946 16574
rect 2998 16522 3012 16574
rect 3064 16522 3078 16574
rect 3130 16522 3144 16574
rect 3196 16553 3210 16574
rect 3262 16553 3276 16574
rect 3328 16553 3342 16574
rect 3394 16553 3408 16574
rect 3460 16553 3474 16574
rect 3526 16553 3540 16574
rect 3592 16553 3606 16574
rect 3658 16553 3672 16574
rect 3201 16522 3210 16553
rect 3273 16522 3276 16553
rect 3526 16522 3527 16553
rect 3592 16522 3599 16553
rect 3658 16522 3671 16553
rect 3724 16522 3738 16574
rect 3790 16522 3804 16574
rect 3856 16522 3870 16574
rect 3922 16522 3936 16574
rect 3988 16553 4002 16574
rect 4054 16553 4068 16574
rect 4120 16553 4134 16574
rect 4186 16553 4200 16574
rect 4252 16553 4266 16574
rect 4318 16553 4332 16574
rect 4384 16553 4398 16574
rect 4450 16553 4464 16574
rect 4516 16553 4590 16574
rect 3993 16522 4002 16553
rect 4065 16522 4068 16553
rect 4318 16522 4319 16553
rect 4384 16522 4391 16553
rect 4450 16522 4463 16553
rect 4516 16522 4535 16553
rect 2769 16519 2807 16522
rect 2841 16519 2879 16522
rect 2913 16519 2951 16522
rect 2985 16519 3023 16522
rect 3057 16519 3095 16522
rect 3129 16519 3167 16522
rect 3201 16519 3239 16522
rect 3273 16519 3311 16522
rect 3345 16519 3383 16522
rect 3417 16519 3455 16522
rect 3489 16519 3527 16522
rect 3561 16519 3599 16522
rect 3633 16519 3671 16522
rect 3705 16519 3743 16522
rect 3777 16519 3815 16522
rect 3849 16519 3887 16522
rect 3921 16519 3959 16522
rect 3993 16519 4031 16522
rect 4065 16519 4103 16522
rect 4137 16519 4175 16522
rect 4209 16519 4247 16522
rect 4281 16519 4319 16522
rect 4353 16519 4391 16522
rect 4425 16519 4463 16522
rect 4497 16519 4535 16522
rect 4569 16519 4590 16553
rect 2642 16508 4590 16519
rect 2642 16480 2746 16508
rect 2798 16480 2813 16508
rect 2865 16480 2880 16508
rect 2642 16446 2663 16480
rect 2697 16446 2735 16480
rect 2798 16456 2807 16480
rect 2865 16456 2879 16480
rect 2932 16456 2946 16508
rect 2998 16456 3012 16508
rect 3064 16456 3078 16508
rect 3130 16456 3144 16508
rect 3196 16480 3210 16508
rect 3262 16480 3276 16508
rect 3328 16480 3342 16508
rect 3394 16480 3408 16508
rect 3460 16480 3474 16508
rect 3526 16480 3540 16508
rect 3592 16480 3606 16508
rect 3658 16480 3672 16508
rect 3201 16456 3210 16480
rect 3273 16456 3276 16480
rect 3526 16456 3527 16480
rect 3592 16456 3599 16480
rect 3658 16456 3671 16480
rect 3724 16456 3738 16508
rect 3790 16456 3804 16508
rect 3856 16456 3870 16508
rect 3922 16456 3936 16508
rect 3988 16480 4002 16508
rect 4054 16480 4068 16508
rect 4120 16480 4134 16508
rect 4186 16480 4200 16508
rect 4252 16480 4266 16508
rect 4318 16480 4332 16508
rect 4384 16480 4398 16508
rect 4450 16480 4464 16508
rect 4516 16480 4590 16508
rect 3993 16456 4002 16480
rect 4065 16456 4068 16480
rect 4318 16456 4319 16480
rect 4384 16456 4391 16480
rect 4450 16456 4463 16480
rect 4516 16456 4535 16480
rect 2769 16446 2807 16456
rect 2841 16446 2879 16456
rect 2913 16446 2951 16456
rect 2985 16446 3023 16456
rect 3057 16446 3095 16456
rect 3129 16446 3167 16456
rect 3201 16446 3239 16456
rect 3273 16446 3311 16456
rect 3345 16446 3383 16456
rect 3417 16446 3455 16456
rect 3489 16446 3527 16456
rect 3561 16446 3599 16456
rect 3633 16446 3671 16456
rect 3705 16446 3743 16456
rect 3777 16446 3815 16456
rect 3849 16446 3887 16456
rect 3921 16446 3959 16456
rect 3993 16446 4031 16456
rect 4065 16446 4103 16456
rect 4137 16446 4175 16456
rect 4209 16446 4247 16456
rect 4281 16446 4319 16456
rect 4353 16446 4391 16456
rect 4425 16446 4463 16456
rect 4497 16446 4535 16456
rect 4569 16446 4590 16480
rect 2642 16442 4590 16446
rect 2642 16407 2746 16442
rect 2798 16407 2813 16442
rect 2865 16407 2880 16442
rect 2642 16373 2663 16407
rect 2697 16373 2735 16407
rect 2798 16390 2807 16407
rect 2865 16390 2879 16407
rect 2932 16390 2946 16442
rect 2998 16390 3012 16442
rect 3064 16390 3078 16442
rect 3130 16390 3144 16442
rect 3196 16407 3210 16442
rect 3262 16407 3276 16442
rect 3328 16407 3342 16442
rect 3394 16407 3408 16442
rect 3460 16407 3474 16442
rect 3526 16407 3540 16442
rect 3592 16407 3606 16442
rect 3658 16407 3672 16442
rect 3201 16390 3210 16407
rect 3273 16390 3276 16407
rect 3526 16390 3527 16407
rect 3592 16390 3599 16407
rect 3658 16390 3671 16407
rect 3724 16390 3738 16442
rect 3790 16390 3804 16442
rect 3856 16390 3870 16442
rect 3922 16390 3936 16442
rect 3988 16407 4002 16442
rect 4054 16407 4068 16442
rect 4120 16407 4134 16442
rect 4186 16407 4200 16442
rect 4252 16407 4266 16442
rect 4318 16407 4332 16442
rect 4384 16407 4398 16442
rect 4450 16407 4464 16442
rect 4516 16407 4590 16442
rect 3993 16390 4002 16407
rect 4065 16390 4068 16407
rect 4318 16390 4319 16407
rect 4384 16390 4391 16407
rect 4450 16390 4463 16407
rect 4516 16390 4535 16407
rect 2769 16376 2807 16390
rect 2841 16376 2879 16390
rect 2913 16376 2951 16390
rect 2985 16376 3023 16390
rect 3057 16376 3095 16390
rect 3129 16376 3167 16390
rect 3201 16376 3239 16390
rect 3273 16376 3311 16390
rect 3345 16376 3383 16390
rect 3417 16376 3455 16390
rect 3489 16376 3527 16390
rect 3561 16376 3599 16390
rect 3633 16376 3671 16390
rect 3705 16376 3743 16390
rect 3777 16376 3815 16390
rect 3849 16376 3887 16390
rect 3921 16376 3959 16390
rect 3993 16376 4031 16390
rect 4065 16376 4103 16390
rect 4137 16376 4175 16390
rect 4209 16376 4247 16390
rect 4281 16376 4319 16390
rect 4353 16376 4391 16390
rect 4425 16376 4463 16390
rect 4497 16376 4535 16390
rect 2798 16373 2807 16376
rect 2865 16373 2879 16376
rect 2642 16334 2746 16373
rect 2798 16334 2813 16373
rect 2865 16334 2880 16373
rect 2642 16300 2663 16334
rect 2697 16300 2735 16334
rect 2798 16324 2807 16334
rect 2865 16324 2879 16334
rect 2932 16324 2946 16376
rect 2998 16324 3012 16376
rect 3064 16324 3078 16376
rect 3130 16324 3144 16376
rect 3201 16373 3210 16376
rect 3273 16373 3276 16376
rect 3526 16373 3527 16376
rect 3592 16373 3599 16376
rect 3658 16373 3671 16376
rect 3196 16334 3210 16373
rect 3262 16334 3276 16373
rect 3328 16334 3342 16373
rect 3394 16334 3408 16373
rect 3460 16334 3474 16373
rect 3526 16334 3540 16373
rect 3592 16334 3606 16373
rect 3658 16334 3672 16373
rect 3201 16324 3210 16334
rect 3273 16324 3276 16334
rect 3526 16324 3527 16334
rect 3592 16324 3599 16334
rect 3658 16324 3671 16334
rect 3724 16324 3738 16376
rect 3790 16324 3804 16376
rect 3856 16324 3870 16376
rect 3922 16324 3936 16376
rect 3993 16373 4002 16376
rect 4065 16373 4068 16376
rect 4318 16373 4319 16376
rect 4384 16373 4391 16376
rect 4450 16373 4463 16376
rect 4516 16373 4535 16376
rect 4569 16373 4590 16407
rect 3988 16334 4002 16373
rect 4054 16334 4068 16373
rect 4120 16334 4134 16373
rect 4186 16334 4200 16373
rect 4252 16334 4266 16373
rect 4318 16334 4332 16373
rect 4384 16334 4398 16373
rect 4450 16334 4464 16373
rect 4516 16334 4590 16373
rect 3993 16324 4002 16334
rect 4065 16324 4068 16334
rect 4318 16324 4319 16334
rect 4384 16324 4391 16334
rect 4450 16324 4463 16334
rect 4516 16324 4535 16334
rect 2769 16310 2807 16324
rect 2841 16310 2879 16324
rect 2913 16310 2951 16324
rect 2985 16310 3023 16324
rect 3057 16310 3095 16324
rect 3129 16310 3167 16324
rect 3201 16310 3239 16324
rect 3273 16310 3311 16324
rect 3345 16310 3383 16324
rect 3417 16310 3455 16324
rect 3489 16310 3527 16324
rect 3561 16310 3599 16324
rect 3633 16310 3671 16324
rect 3705 16310 3743 16324
rect 3777 16310 3815 16324
rect 3849 16310 3887 16324
rect 3921 16310 3959 16324
rect 3993 16310 4031 16324
rect 4065 16310 4103 16324
rect 4137 16310 4175 16324
rect 4209 16310 4247 16324
rect 4281 16310 4319 16324
rect 4353 16310 4391 16324
rect 4425 16310 4463 16324
rect 4497 16310 4535 16324
rect 2798 16300 2807 16310
rect 2865 16300 2879 16310
rect 2642 16261 2746 16300
rect 2798 16261 2813 16300
rect 2865 16261 2880 16300
rect 2642 16227 2663 16261
rect 2697 16227 2735 16261
rect 2798 16258 2807 16261
rect 2865 16258 2879 16261
rect 2932 16258 2946 16310
rect 2998 16258 3012 16310
rect 3064 16258 3078 16310
rect 3130 16258 3144 16310
rect 3201 16300 3210 16310
rect 3273 16300 3276 16310
rect 3526 16300 3527 16310
rect 3592 16300 3599 16310
rect 3658 16300 3671 16310
rect 3196 16261 3210 16300
rect 3262 16261 3276 16300
rect 3328 16261 3342 16300
rect 3394 16261 3408 16300
rect 3460 16261 3474 16300
rect 3526 16261 3540 16300
rect 3592 16261 3606 16300
rect 3658 16261 3672 16300
rect 3201 16258 3210 16261
rect 3273 16258 3276 16261
rect 3526 16258 3527 16261
rect 3592 16258 3599 16261
rect 3658 16258 3671 16261
rect 3724 16258 3738 16310
rect 3790 16258 3804 16310
rect 3856 16258 3870 16310
rect 3922 16258 3936 16310
rect 3993 16300 4002 16310
rect 4065 16300 4068 16310
rect 4318 16300 4319 16310
rect 4384 16300 4391 16310
rect 4450 16300 4463 16310
rect 4516 16300 4535 16310
rect 4569 16300 4590 16334
rect 3988 16261 4002 16300
rect 4054 16261 4068 16300
rect 4120 16261 4134 16300
rect 4186 16261 4200 16300
rect 4252 16261 4266 16300
rect 4318 16261 4332 16300
rect 4384 16261 4398 16300
rect 4450 16261 4464 16300
rect 4516 16261 4590 16300
rect 3993 16258 4002 16261
rect 4065 16258 4068 16261
rect 4318 16258 4319 16261
rect 4384 16258 4391 16261
rect 4450 16258 4463 16261
rect 4516 16258 4535 16261
rect 2769 16244 2807 16258
rect 2841 16244 2879 16258
rect 2913 16244 2951 16258
rect 2985 16244 3023 16258
rect 3057 16244 3095 16258
rect 3129 16244 3167 16258
rect 3201 16244 3239 16258
rect 3273 16244 3311 16258
rect 3345 16244 3383 16258
rect 3417 16244 3455 16258
rect 3489 16244 3527 16258
rect 3561 16244 3599 16258
rect 3633 16244 3671 16258
rect 3705 16244 3743 16258
rect 3777 16244 3815 16258
rect 3849 16244 3887 16258
rect 3921 16244 3959 16258
rect 3993 16244 4031 16258
rect 4065 16244 4103 16258
rect 4137 16244 4175 16258
rect 4209 16244 4247 16258
rect 4281 16244 4319 16258
rect 4353 16244 4391 16258
rect 4425 16244 4463 16258
rect 4497 16244 4535 16258
rect 2798 16227 2807 16244
rect 2865 16227 2879 16244
rect 2642 16192 2746 16227
rect 2798 16192 2813 16227
rect 2865 16192 2880 16227
rect 2932 16192 2946 16244
rect 2998 16192 3012 16244
rect 3064 16192 3078 16244
rect 3130 16192 3144 16244
rect 3201 16227 3210 16244
rect 3273 16227 3276 16244
rect 3526 16227 3527 16244
rect 3592 16227 3599 16244
rect 3658 16227 3671 16244
rect 3196 16192 3210 16227
rect 3262 16192 3276 16227
rect 3328 16192 3342 16227
rect 3394 16192 3408 16227
rect 3460 16192 3474 16227
rect 3526 16192 3540 16227
rect 3592 16192 3606 16227
rect 3658 16192 3672 16227
rect 3724 16192 3738 16244
rect 3790 16192 3804 16244
rect 3856 16192 3870 16244
rect 3922 16192 3936 16244
rect 3993 16227 4002 16244
rect 4065 16227 4068 16244
rect 4318 16227 4319 16244
rect 4384 16227 4391 16244
rect 4450 16227 4463 16244
rect 4516 16227 4535 16244
rect 4569 16227 4590 16261
rect 3988 16192 4002 16227
rect 4054 16192 4068 16227
rect 4120 16192 4134 16227
rect 4186 16192 4200 16227
rect 4252 16192 4266 16227
rect 4318 16192 4332 16227
rect 4384 16192 4398 16227
rect 4450 16192 4464 16227
rect 4516 16192 4590 16227
rect 2642 16188 4590 16192
rect 2642 16154 2663 16188
rect 2697 16154 2735 16188
rect 2769 16178 2807 16188
rect 2841 16178 2879 16188
rect 2913 16178 2951 16188
rect 2985 16178 3023 16188
rect 3057 16178 3095 16188
rect 3129 16178 3167 16188
rect 3201 16178 3239 16188
rect 3273 16178 3311 16188
rect 3345 16178 3383 16188
rect 3417 16178 3455 16188
rect 3489 16178 3527 16188
rect 3561 16178 3599 16188
rect 3633 16178 3671 16188
rect 3705 16178 3743 16188
rect 3777 16178 3815 16188
rect 3849 16178 3887 16188
rect 3921 16178 3959 16188
rect 3993 16178 4031 16188
rect 4065 16178 4103 16188
rect 4137 16178 4175 16188
rect 4209 16178 4247 16188
rect 4281 16178 4319 16188
rect 4353 16178 4391 16188
rect 4425 16178 4463 16188
rect 4497 16178 4535 16188
rect 2798 16154 2807 16178
rect 2865 16154 2879 16178
rect 2642 16126 2746 16154
rect 2798 16126 2813 16154
rect 2865 16126 2880 16154
rect 2932 16126 2946 16178
rect 2998 16126 3012 16178
rect 3064 16126 3078 16178
rect 3130 16126 3144 16178
rect 3201 16154 3210 16178
rect 3273 16154 3276 16178
rect 3526 16154 3527 16178
rect 3592 16154 3599 16178
rect 3658 16154 3671 16178
rect 3196 16126 3210 16154
rect 3262 16126 3276 16154
rect 3328 16126 3342 16154
rect 3394 16126 3408 16154
rect 3460 16126 3474 16154
rect 3526 16126 3540 16154
rect 3592 16126 3606 16154
rect 3658 16126 3672 16154
rect 3724 16126 3738 16178
rect 3790 16126 3804 16178
rect 3856 16126 3870 16178
rect 3922 16126 3936 16178
rect 3993 16154 4002 16178
rect 4065 16154 4068 16178
rect 4318 16154 4319 16178
rect 4384 16154 4391 16178
rect 4450 16154 4463 16178
rect 4516 16154 4535 16178
rect 4569 16154 4590 16188
rect 3988 16126 4002 16154
rect 4054 16126 4068 16154
rect 4120 16126 4134 16154
rect 4186 16126 4200 16154
rect 4252 16126 4266 16154
rect 4318 16126 4332 16154
rect 4384 16126 4398 16154
rect 4450 16126 4464 16154
rect 4516 16126 4590 16154
rect 2642 16115 4590 16126
rect 2642 16081 2663 16115
rect 2697 16081 2735 16115
rect 2769 16112 2807 16115
rect 2841 16112 2879 16115
rect 2913 16112 2951 16115
rect 2985 16112 3023 16115
rect 3057 16112 3095 16115
rect 3129 16112 3167 16115
rect 3201 16112 3239 16115
rect 3273 16112 3311 16115
rect 3345 16112 3383 16115
rect 3417 16112 3455 16115
rect 3489 16112 3527 16115
rect 3561 16112 3599 16115
rect 3633 16112 3671 16115
rect 3705 16112 3743 16115
rect 3777 16112 3815 16115
rect 3849 16112 3887 16115
rect 3921 16112 3959 16115
rect 3993 16112 4031 16115
rect 4065 16112 4103 16115
rect 4137 16112 4175 16115
rect 4209 16112 4247 16115
rect 4281 16112 4319 16115
rect 4353 16112 4391 16115
rect 4425 16112 4463 16115
rect 4497 16112 4535 16115
rect 2798 16081 2807 16112
rect 2865 16081 2879 16112
rect 2642 16060 2746 16081
rect 2798 16060 2813 16081
rect 2865 16060 2880 16081
rect 2932 16060 2946 16112
rect 2998 16060 3012 16112
rect 3064 16060 3078 16112
rect 3130 16060 3144 16112
rect 3201 16081 3210 16112
rect 3273 16081 3276 16112
rect 3526 16081 3527 16112
rect 3592 16081 3599 16112
rect 3658 16081 3671 16112
rect 3196 16060 3210 16081
rect 3262 16060 3276 16081
rect 3328 16060 3342 16081
rect 3394 16060 3408 16081
rect 3460 16060 3474 16081
rect 3526 16060 3540 16081
rect 3592 16060 3606 16081
rect 3658 16060 3672 16081
rect 3724 16060 3738 16112
rect 3790 16060 3804 16112
rect 3856 16060 3870 16112
rect 3922 16060 3936 16112
rect 3993 16081 4002 16112
rect 4065 16081 4068 16112
rect 4318 16081 4319 16112
rect 4384 16081 4391 16112
rect 4450 16081 4463 16112
rect 4516 16081 4535 16112
rect 4569 16081 4590 16115
rect 3988 16060 4002 16081
rect 4054 16060 4068 16081
rect 4120 16060 4134 16081
rect 4186 16060 4200 16081
rect 4252 16060 4266 16081
rect 4318 16060 4332 16081
rect 4384 16060 4398 16081
rect 4450 16060 4464 16081
rect 4516 16060 4590 16081
rect 2642 16046 4590 16060
rect 2642 16042 2746 16046
rect 2798 16042 2813 16046
rect 2865 16042 2880 16046
rect 2642 16008 2663 16042
rect 2697 16008 2735 16042
rect 2798 16008 2807 16042
rect 2865 16008 2879 16042
rect 2642 15994 2746 16008
rect 2798 15994 2813 16008
rect 2865 15994 2880 16008
rect 2932 15994 2946 16046
rect 2998 15994 3012 16046
rect 3064 15994 3078 16046
rect 3130 15994 3144 16046
rect 3196 16042 3210 16046
rect 3262 16042 3276 16046
rect 3328 16042 3342 16046
rect 3394 16042 3408 16046
rect 3460 16042 3474 16046
rect 3526 16042 3540 16046
rect 3592 16042 3606 16046
rect 3658 16042 3672 16046
rect 3201 16008 3210 16042
rect 3273 16008 3276 16042
rect 3526 16008 3527 16042
rect 3592 16008 3599 16042
rect 3658 16008 3671 16042
rect 3196 15994 3210 16008
rect 3262 15994 3276 16008
rect 3328 15994 3342 16008
rect 3394 15994 3408 16008
rect 3460 15994 3474 16008
rect 3526 15994 3540 16008
rect 3592 15994 3606 16008
rect 3658 15994 3672 16008
rect 3724 15994 3738 16046
rect 3790 15994 3804 16046
rect 3856 15994 3870 16046
rect 3922 15994 3936 16046
rect 3988 16042 4002 16046
rect 4054 16042 4068 16046
rect 4120 16042 4134 16046
rect 4186 16042 4200 16046
rect 4252 16042 4266 16046
rect 4318 16042 4332 16046
rect 4384 16042 4398 16046
rect 4450 16042 4464 16046
rect 4516 16042 4590 16046
rect 3993 16008 4002 16042
rect 4065 16008 4068 16042
rect 4318 16008 4319 16042
rect 4384 16008 4391 16042
rect 4450 16008 4463 16042
rect 4516 16008 4535 16042
rect 4569 16008 4590 16042
rect 3988 15994 4002 16008
rect 4054 15994 4068 16008
rect 4120 15994 4134 16008
rect 4186 15994 4200 16008
rect 4252 15994 4266 16008
rect 4318 15994 4332 16008
rect 4384 15994 4398 16008
rect 4450 15994 4464 16008
rect 4516 15994 4590 16008
rect 2642 15969 4590 15994
rect 2642 15935 2663 15969
rect 2697 15935 2735 15969
rect 2769 15935 2807 15969
rect 2841 15935 2879 15969
rect 2913 15935 2951 15969
rect 2985 15935 3023 15969
rect 3057 15935 3095 15969
rect 3129 15935 3167 15969
rect 3201 15935 3239 15969
rect 3273 15935 3311 15969
rect 3345 15935 3383 15969
rect 3417 15935 3455 15969
rect 3489 15935 3527 15969
rect 3561 15935 3599 15969
rect 3633 15935 3671 15969
rect 3705 15935 3743 15969
rect 3777 15935 3815 15969
rect 3849 15935 3887 15969
rect 3921 15935 3959 15969
rect 3993 15935 4031 15969
rect 4065 15935 4103 15969
rect 4137 15935 4175 15969
rect 4209 15935 4247 15969
rect 4281 15935 4319 15969
rect 4353 15935 4391 15969
rect 4425 15935 4463 15969
rect 4497 15935 4535 15969
rect 4569 15935 4590 15969
rect 2642 15923 4590 15935
rect 4773 27165 4928 29071
rect 8044 29109 8050 29143
rect 8084 29133 8224 29143
rect 8084 29109 8184 29133
rect 8044 29099 8184 29109
rect 8218 29099 8224 29133
rect 8044 29071 8224 29099
rect 8044 29037 8050 29071
rect 8084 29061 8224 29071
rect 8084 29037 8184 29061
rect 8044 29027 8184 29037
rect 8218 29027 8224 29061
rect 8044 28999 8224 29027
rect 8044 28965 8050 28999
rect 8084 28989 8224 28999
rect 8084 28965 8184 28989
rect 8044 28955 8184 28965
rect 8218 28955 8224 28989
rect 8044 28927 8224 28955
rect 8044 28893 8050 28927
rect 8084 28917 8224 28927
rect 8084 28893 8184 28917
rect 8044 28883 8184 28893
rect 8218 28883 8224 28917
rect 8044 28855 8224 28883
rect 8044 28821 8050 28855
rect 8084 28845 8224 28855
rect 8084 28821 8184 28845
rect 8044 28811 8184 28821
rect 8218 28811 8224 28845
rect 8044 28783 8224 28811
rect 8044 28749 8050 28783
rect 8084 28773 8224 28783
rect 8084 28749 8184 28773
rect 8044 28739 8184 28749
rect 8218 28739 8224 28773
rect 5040 28720 5158 28726
rect 5092 28668 5106 28720
rect 5040 28651 5158 28668
rect 5092 28599 5106 28651
rect 5040 28582 5158 28599
rect 5092 28530 5106 28582
rect 5040 28513 5158 28530
rect 5092 28461 5106 28513
rect 5040 28444 5158 28461
rect 5092 28422 5106 28444
rect 5040 28375 5046 28392
rect 5152 28375 5158 28392
rect 5040 28306 5046 28323
rect 5152 28306 5158 28323
rect 5040 28236 5046 28254
rect 5152 28236 5158 28254
rect 5040 28166 5046 28184
rect 5152 28166 5158 28184
rect 5040 27380 5046 28114
rect 5152 27380 5158 28114
rect 5040 27368 5158 27380
rect 5317 28714 5435 28726
rect 5317 28680 5323 28714
rect 5357 28680 5395 28714
rect 5429 28680 5435 28714
rect 5317 28641 5435 28680
rect 5317 28607 5323 28641
rect 5357 28607 5395 28641
rect 5429 28607 5435 28641
rect 5317 28568 5435 28607
rect 5317 28534 5323 28568
rect 5357 28534 5395 28568
rect 5429 28534 5435 28568
rect 5317 28495 5435 28534
rect 5317 28461 5323 28495
rect 5357 28461 5395 28495
rect 5429 28461 5435 28495
rect 5317 28422 5435 28461
rect 5317 27982 5323 28422
rect 5429 27982 5435 28422
rect 5317 27913 5323 27930
rect 5429 27913 5435 27930
rect 5317 27844 5323 27861
rect 5429 27844 5435 27861
rect 5317 27775 5323 27792
rect 5429 27775 5435 27792
rect 5317 27706 5323 27723
rect 5429 27706 5435 27723
rect 5317 27636 5323 27654
rect 5429 27636 5435 27654
rect 5317 27566 5323 27584
rect 5429 27566 5435 27584
rect 5317 27496 5323 27514
rect 5429 27496 5435 27514
rect 5317 27426 5323 27444
rect 5429 27426 5435 27444
rect 5369 27374 5383 27380
rect 5317 27368 5435 27374
rect 5594 28720 5712 28726
rect 5646 28668 5660 28720
rect 5594 28651 5712 28668
rect 5646 28599 5660 28651
rect 5594 28582 5712 28599
rect 5646 28530 5660 28582
rect 5594 28513 5712 28530
rect 5646 28461 5660 28513
rect 5594 28444 5712 28461
rect 5646 28422 5660 28444
rect 5594 28375 5600 28392
rect 5706 28375 5712 28392
rect 5594 28306 5600 28323
rect 5706 28306 5712 28323
rect 5594 28236 5600 28254
rect 5706 28236 5712 28254
rect 5594 28166 5600 28184
rect 5706 28166 5712 28184
rect 5594 27380 5600 28114
rect 5706 27380 5712 28114
rect 5594 27368 5712 27380
rect 5871 28714 5989 28726
rect 5871 28680 5877 28714
rect 5911 28680 5949 28714
rect 5983 28680 5989 28714
rect 5871 28641 5989 28680
rect 5871 28607 5877 28641
rect 5911 28607 5949 28641
rect 5983 28607 5989 28641
rect 5871 28568 5989 28607
rect 5871 28534 5877 28568
rect 5911 28534 5949 28568
rect 5983 28534 5989 28568
rect 5871 28495 5989 28534
rect 5871 28461 5877 28495
rect 5911 28461 5949 28495
rect 5983 28461 5989 28495
rect 5871 28422 5989 28461
rect 5871 27982 5877 28422
rect 5983 27982 5989 28422
rect 5871 27913 5877 27930
rect 5983 27913 5989 27930
rect 5871 27844 5877 27861
rect 5983 27844 5989 27861
rect 5871 27775 5877 27792
rect 5983 27775 5989 27792
rect 5871 27706 5877 27723
rect 5983 27706 5989 27723
rect 5871 27636 5877 27654
rect 5983 27636 5989 27654
rect 5871 27566 5877 27584
rect 5983 27566 5989 27584
rect 5871 27496 5877 27514
rect 5983 27496 5989 27514
rect 5871 27426 5877 27444
rect 5983 27426 5989 27444
rect 5923 27374 5937 27380
rect 5871 27368 5989 27374
rect 6148 28720 6266 28726
rect 6200 28668 6214 28720
rect 6148 28651 6266 28668
rect 6200 28599 6214 28651
rect 6148 28582 6266 28599
rect 6200 28530 6214 28582
rect 6148 28513 6266 28530
rect 6200 28461 6214 28513
rect 6148 28444 6266 28461
rect 6200 28422 6214 28444
rect 6148 28375 6154 28392
rect 6260 28375 6266 28392
rect 6148 28306 6154 28323
rect 6260 28306 6266 28323
rect 6148 28236 6154 28254
rect 6260 28236 6266 28254
rect 6148 28166 6154 28184
rect 6260 28166 6266 28184
rect 6148 27380 6154 28114
rect 6260 27380 6266 28114
rect 6148 27368 6266 27380
rect 6425 28714 6543 28726
rect 6425 28680 6431 28714
rect 6465 28680 6503 28714
rect 6537 28680 6543 28714
rect 6425 28641 6543 28680
rect 6425 28607 6431 28641
rect 6465 28607 6503 28641
rect 6537 28607 6543 28641
rect 6425 28568 6543 28607
rect 6425 28534 6431 28568
rect 6465 28534 6503 28568
rect 6537 28534 6543 28568
rect 6425 28495 6543 28534
rect 6425 28461 6431 28495
rect 6465 28461 6503 28495
rect 6537 28461 6543 28495
rect 6425 28422 6543 28461
rect 6425 27982 6431 28422
rect 6537 27982 6543 28422
rect 6425 27913 6431 27930
rect 6537 27913 6543 27930
rect 6425 27844 6431 27861
rect 6537 27844 6543 27861
rect 6425 27775 6431 27792
rect 6537 27775 6543 27792
rect 6425 27706 6431 27723
rect 6537 27706 6543 27723
rect 6425 27636 6431 27654
rect 6537 27636 6543 27654
rect 6425 27566 6431 27584
rect 6537 27566 6543 27584
rect 6425 27496 6431 27514
rect 6537 27496 6543 27514
rect 6425 27426 6431 27444
rect 6537 27426 6543 27444
rect 6477 27374 6491 27380
rect 6425 27368 6543 27374
rect 6702 28720 6820 28726
rect 6754 28668 6768 28720
rect 6702 28651 6820 28668
rect 6754 28599 6768 28651
rect 6702 28582 6820 28599
rect 6754 28530 6768 28582
rect 6702 28513 6820 28530
rect 6754 28461 6768 28513
rect 6702 28444 6820 28461
rect 6754 28422 6768 28444
rect 6702 28375 6708 28392
rect 6814 28375 6820 28392
rect 6702 28306 6708 28323
rect 6814 28306 6820 28323
rect 6702 28236 6708 28254
rect 6814 28236 6820 28254
rect 6702 28166 6708 28184
rect 6814 28166 6820 28184
rect 6702 27380 6708 28114
rect 6814 27380 6820 28114
rect 6702 27368 6820 27380
rect 6979 28714 7097 28726
rect 6979 28680 6985 28714
rect 7019 28680 7057 28714
rect 7091 28680 7097 28714
rect 6979 28641 7097 28680
rect 6979 28607 6985 28641
rect 7019 28607 7057 28641
rect 7091 28607 7097 28641
rect 6979 28568 7097 28607
rect 6979 28534 6985 28568
rect 7019 28534 7057 28568
rect 7091 28534 7097 28568
rect 6979 28495 7097 28534
rect 6979 28461 6985 28495
rect 7019 28461 7057 28495
rect 7091 28461 7097 28495
rect 6979 28422 7097 28461
rect 6979 27982 6985 28422
rect 7091 27982 7097 28422
rect 6979 27913 6985 27930
rect 7091 27913 7097 27930
rect 6979 27844 6985 27861
rect 7091 27844 7097 27861
rect 6979 27775 6985 27792
rect 7091 27775 7097 27792
rect 6979 27706 6985 27723
rect 7091 27706 7097 27723
rect 6979 27636 6985 27654
rect 7091 27636 7097 27654
rect 6979 27566 6985 27584
rect 7091 27566 7097 27584
rect 6979 27496 6985 27514
rect 7091 27496 7097 27514
rect 6979 27426 6985 27444
rect 7091 27426 7097 27444
rect 7031 27374 7045 27380
rect 6979 27368 7097 27374
rect 7256 28720 7374 28726
rect 7308 28668 7322 28720
rect 7256 28651 7374 28668
rect 7308 28599 7322 28651
rect 7256 28582 7374 28599
rect 7308 28530 7322 28582
rect 7256 28513 7374 28530
rect 7308 28461 7322 28513
rect 7256 28444 7374 28461
rect 7308 28422 7322 28444
rect 7256 28375 7262 28392
rect 7368 28375 7374 28392
rect 7256 28306 7262 28323
rect 7368 28306 7374 28323
rect 7256 28236 7262 28254
rect 7368 28236 7374 28254
rect 7256 28166 7262 28184
rect 7368 28166 7374 28184
rect 7256 27380 7262 28114
rect 7368 27380 7374 28114
rect 7256 27368 7374 27380
rect 7533 28714 7651 28726
rect 7533 28680 7539 28714
rect 7573 28680 7611 28714
rect 7645 28680 7651 28714
rect 7533 28641 7651 28680
rect 7533 28607 7539 28641
rect 7573 28607 7611 28641
rect 7645 28607 7651 28641
rect 7533 28568 7651 28607
rect 7533 28534 7539 28568
rect 7573 28534 7611 28568
rect 7645 28534 7651 28568
rect 7533 28495 7651 28534
rect 7533 28461 7539 28495
rect 7573 28461 7611 28495
rect 7645 28461 7651 28495
rect 7533 28422 7651 28461
rect 7533 27982 7539 28422
rect 7645 27982 7651 28422
rect 7533 27913 7539 27930
rect 7645 27913 7651 27930
rect 7533 27844 7539 27861
rect 7645 27844 7651 27861
rect 7533 27775 7539 27792
rect 7645 27775 7651 27792
rect 7533 27706 7539 27723
rect 7645 27706 7651 27723
rect 7533 27636 7539 27654
rect 7645 27636 7651 27654
rect 7533 27566 7539 27584
rect 7645 27566 7651 27584
rect 7533 27496 7539 27514
rect 7645 27496 7651 27514
rect 7533 27426 7539 27444
rect 7645 27426 7651 27444
rect 7585 27374 7599 27380
rect 7533 27368 7651 27374
rect 7810 28720 7928 28726
rect 7862 28668 7876 28720
rect 7810 28651 7928 28668
rect 7862 28599 7876 28651
rect 7810 28582 7928 28599
rect 7862 28530 7876 28582
rect 7810 28513 7928 28530
rect 7862 28461 7876 28513
rect 7810 28444 7928 28461
rect 7862 28422 7876 28444
rect 7810 28375 7816 28392
rect 7922 28375 7928 28392
rect 7810 28306 7816 28323
rect 7922 28306 7928 28323
rect 7810 28236 7816 28254
rect 7922 28236 7928 28254
rect 7810 28166 7816 28184
rect 7922 28166 7928 28184
rect 7810 27380 7816 28114
rect 7922 27380 7928 28114
rect 7810 27368 7928 27380
rect 8044 28724 8224 28739
rect 8044 28672 8047 28724
rect 8099 28672 8169 28724
rect 8221 28672 8224 28724
rect 8044 28667 8184 28672
rect 8218 28667 8224 28672
rect 8044 28655 8224 28667
rect 8044 28603 8047 28655
rect 8099 28603 8169 28655
rect 8221 28603 8224 28655
rect 8044 28595 8184 28603
rect 8218 28595 8224 28603
rect 8044 28586 8224 28595
rect 8044 28534 8047 28586
rect 8099 28534 8169 28586
rect 8221 28534 8224 28586
rect 8044 28533 8050 28534
rect 8084 28533 8184 28534
rect 8044 28523 8184 28533
rect 8218 28523 8224 28534
rect 8044 28517 8224 28523
rect 8044 28465 8047 28517
rect 8099 28465 8169 28517
rect 8221 28465 8224 28517
rect 8044 28461 8050 28465
rect 8084 28461 8184 28465
rect 8044 28451 8184 28461
rect 8218 28451 8224 28465
rect 8044 28448 8224 28451
rect 8044 28396 8047 28448
rect 8099 28396 8169 28448
rect 8221 28396 8224 28448
rect 8044 28389 8050 28396
rect 8084 28389 8184 28396
rect 8044 28379 8184 28389
rect 8218 28379 8224 28396
rect 8044 28378 8224 28379
rect 8044 28326 8047 28378
rect 8099 28326 8169 28378
rect 8221 28326 8224 28378
rect 8044 28317 8050 28326
rect 8084 28317 8184 28326
rect 8044 28308 8184 28317
rect 8218 28308 8224 28326
rect 8044 28256 8047 28308
rect 8099 28256 8169 28308
rect 8221 28256 8224 28308
rect 8044 28245 8050 28256
rect 8084 28245 8184 28256
rect 8044 28238 8184 28245
rect 8218 28238 8224 28256
rect 8044 28186 8047 28238
rect 8099 28186 8169 28238
rect 8221 28186 8224 28238
rect 8044 28173 8050 28186
rect 8084 28173 8184 28186
rect 8044 28168 8184 28173
rect 8218 28168 8224 28186
rect 8044 28116 8047 28168
rect 8099 28116 8169 28168
rect 8221 28116 8224 28168
rect 8044 28101 8050 28116
rect 8084 28101 8184 28116
rect 8044 28091 8184 28101
rect 8218 28091 8224 28116
rect 8044 28063 8224 28091
rect 8044 28029 8050 28063
rect 8084 28053 8224 28063
rect 8084 28029 8184 28053
rect 8044 28019 8184 28029
rect 8218 28019 8224 28053
rect 8044 27991 8224 28019
rect 8044 27957 8050 27991
rect 8084 27981 8224 27991
rect 8084 27957 8184 27981
rect 8044 27947 8184 27957
rect 8218 27947 8224 27981
rect 8044 27919 8224 27947
rect 8044 27885 8050 27919
rect 8084 27909 8224 27919
rect 8084 27885 8184 27909
rect 8044 27875 8184 27885
rect 8218 27875 8224 27909
rect 8044 27847 8224 27875
rect 8044 27813 8050 27847
rect 8084 27837 8224 27847
rect 8084 27813 8184 27837
rect 8044 27803 8184 27813
rect 8218 27803 8224 27837
rect 8044 27775 8224 27803
rect 8044 27741 8050 27775
rect 8084 27765 8224 27775
rect 8084 27741 8184 27765
rect 8044 27731 8184 27741
rect 8218 27731 8224 27765
rect 8044 27703 8224 27731
rect 8044 27669 8050 27703
rect 8084 27693 8224 27703
rect 8084 27669 8184 27693
rect 8044 27659 8184 27669
rect 8218 27659 8224 27693
rect 8044 27631 8224 27659
rect 8044 27597 8050 27631
rect 8084 27621 8224 27631
rect 8084 27597 8184 27621
rect 8044 27587 8184 27597
rect 8218 27587 8224 27621
rect 8044 27559 8224 27587
rect 8044 27525 8050 27559
rect 8084 27549 8224 27559
rect 8084 27525 8184 27549
rect 8044 27515 8184 27525
rect 8218 27515 8224 27549
rect 8044 27487 8224 27515
rect 8044 27453 8050 27487
rect 8084 27477 8224 27487
rect 8084 27453 8184 27477
rect 8044 27443 8184 27453
rect 8218 27443 8224 27477
rect 8044 27415 8224 27443
rect 8044 27381 8050 27415
rect 8084 27405 8224 27415
rect 8084 27381 8184 27405
rect 8044 27371 8184 27381
rect 8218 27371 8224 27405
rect 8044 27343 8224 27371
rect 8044 27309 8050 27343
rect 8084 27333 8224 27343
rect 8084 27309 8184 27333
rect 8044 27299 8184 27309
rect 8218 27299 8224 27333
rect 8044 27271 8224 27299
rect 8044 27237 8050 27271
rect 8084 27261 8224 27271
rect 8084 27237 8184 27261
rect 8044 27227 8184 27237
rect 8218 27227 8224 27261
rect 8044 27199 8224 27227
tri 4928 27165 4947 27184 sw
rect 8044 27165 8050 27199
rect 8084 27189 8224 27199
rect 8084 27165 8184 27189
rect 4773 27155 4947 27165
tri 4947 27155 4957 27165 sw
rect 8044 27155 8184 27165
rect 8218 27155 8224 27189
rect 4773 27152 4957 27155
tri 4957 27152 4960 27155 sw
rect 4773 27105 7729 27152
rect 4773 27071 5251 27105
rect 5285 27071 5326 27105
rect 5360 27071 5401 27105
rect 5435 27071 5476 27105
rect 5510 27071 5551 27105
rect 5585 27071 5626 27105
rect 5660 27071 5701 27105
rect 5735 27071 5776 27105
rect 5810 27071 5851 27105
rect 5885 27071 5926 27105
rect 5960 27071 6001 27105
rect 6035 27071 6076 27105
rect 6110 27071 6151 27105
rect 6185 27071 6225 27105
rect 6259 27071 6299 27105
rect 6333 27071 6373 27105
rect 6407 27071 6447 27105
rect 6481 27071 6521 27105
rect 6555 27071 6595 27105
rect 6629 27071 6669 27105
rect 6703 27071 6743 27105
rect 6777 27071 6817 27105
rect 6851 27071 6891 27105
rect 6925 27071 7729 27105
rect 4773 27032 7729 27071
rect 8044 27127 8224 27155
rect 8044 27093 8050 27127
rect 8084 27117 8224 27127
rect 8084 27093 8184 27117
rect 8044 27083 8184 27093
rect 8218 27083 8224 27117
rect 8044 27055 8224 27083
rect 4773 27021 4977 27032
tri 4977 27021 4988 27032 nw
rect 8044 27021 8050 27055
rect 8084 27045 8224 27055
rect 8084 27021 8184 27045
rect 4773 27011 4967 27021
tri 4967 27011 4977 27021 nw
rect 8044 27011 8184 27021
rect 8218 27011 8224 27045
rect 4773 26983 4939 27011
tri 4939 26983 4967 27011 nw
rect 8044 26983 8224 27011
rect 4773 25183 4928 26983
tri 4928 26972 4939 26983 nw
rect 8044 26949 8050 26983
rect 8084 26973 8224 26983
rect 8084 26949 8184 26973
rect 8044 26939 8184 26949
rect 8218 26939 8224 26973
rect 8044 26911 8224 26939
rect 8044 26877 8050 26911
rect 8084 26901 8224 26911
rect 8084 26877 8184 26901
rect 8044 26867 8184 26877
rect 8218 26867 8224 26901
rect 8044 26839 8224 26867
rect 8044 26805 8050 26839
rect 8084 26829 8224 26839
rect 8084 26805 8184 26829
rect 8044 26795 8184 26805
rect 8218 26795 8224 26829
rect 8044 26767 8224 26795
rect 8044 26733 8050 26767
rect 8084 26757 8224 26767
rect 8084 26733 8184 26757
rect 5040 26720 5158 26726
rect 5092 26668 5106 26720
rect 5040 26651 5158 26668
rect 5092 26599 5106 26651
rect 5040 26582 5158 26599
rect 5092 26530 5106 26582
rect 5040 26513 5158 26530
rect 5092 26461 5106 26513
rect 5040 26444 5158 26461
rect 5092 26422 5106 26444
rect 5040 26375 5046 26392
rect 5152 26375 5158 26392
rect 5040 26306 5046 26323
rect 5152 26306 5158 26323
rect 5040 26236 5046 26254
rect 5152 26236 5158 26254
rect 5040 26166 5046 26184
rect 5152 26166 5158 26184
rect 5040 25380 5046 26114
rect 5152 25380 5158 26114
rect 5040 25368 5158 25380
rect 5317 26714 5435 26726
rect 5317 26680 5323 26714
rect 5357 26680 5395 26714
rect 5429 26680 5435 26714
rect 5317 26641 5435 26680
rect 5317 26607 5323 26641
rect 5357 26607 5395 26641
rect 5429 26607 5435 26641
rect 5317 26568 5435 26607
rect 5317 26534 5323 26568
rect 5357 26534 5395 26568
rect 5429 26534 5435 26568
rect 5317 26495 5435 26534
rect 5317 26461 5323 26495
rect 5357 26461 5395 26495
rect 5429 26461 5435 26495
rect 5317 26422 5435 26461
rect 5317 25982 5323 26422
rect 5429 25982 5435 26422
rect 5317 25913 5323 25930
rect 5429 25913 5435 25930
rect 5317 25844 5323 25861
rect 5429 25844 5435 25861
rect 5317 25775 5323 25792
rect 5429 25775 5435 25792
rect 5317 25706 5323 25723
rect 5429 25706 5435 25723
rect 5317 25636 5323 25654
rect 5429 25636 5435 25654
rect 5317 25566 5323 25584
rect 5429 25566 5435 25584
rect 5317 25496 5323 25514
rect 5429 25496 5435 25514
rect 5317 25426 5323 25444
rect 5429 25426 5435 25444
rect 5369 25374 5383 25380
rect 5317 25368 5435 25374
rect 5594 26720 5712 26726
rect 5646 26668 5660 26720
rect 5594 26651 5712 26668
rect 5646 26599 5660 26651
rect 5594 26582 5712 26599
rect 5646 26530 5660 26582
rect 5594 26513 5712 26530
rect 5646 26461 5660 26513
rect 5594 26444 5712 26461
rect 5646 26422 5660 26444
rect 5594 26375 5600 26392
rect 5706 26375 5712 26392
rect 5594 26306 5600 26323
rect 5706 26306 5712 26323
rect 5594 26236 5600 26254
rect 5706 26236 5712 26254
rect 5594 26166 5600 26184
rect 5706 26166 5712 26184
rect 5594 25380 5600 26114
rect 5706 25380 5712 26114
rect 5594 25368 5712 25380
rect 5871 26714 5989 26726
rect 5871 26680 5877 26714
rect 5911 26680 5949 26714
rect 5983 26680 5989 26714
rect 5871 26641 5989 26680
rect 5871 26607 5877 26641
rect 5911 26607 5949 26641
rect 5983 26607 5989 26641
rect 5871 26568 5989 26607
rect 5871 26534 5877 26568
rect 5911 26534 5949 26568
rect 5983 26534 5989 26568
rect 5871 26495 5989 26534
rect 5871 26461 5877 26495
rect 5911 26461 5949 26495
rect 5983 26461 5989 26495
rect 5871 26422 5989 26461
rect 5871 25982 5877 26422
rect 5983 25982 5989 26422
rect 5871 25913 5877 25930
rect 5983 25913 5989 25930
rect 5871 25844 5877 25861
rect 5983 25844 5989 25861
rect 5871 25775 5877 25792
rect 5983 25775 5989 25792
rect 5871 25706 5877 25723
rect 5983 25706 5989 25723
rect 5871 25636 5877 25654
rect 5983 25636 5989 25654
rect 5871 25566 5877 25584
rect 5983 25566 5989 25584
rect 5871 25496 5877 25514
rect 5983 25496 5989 25514
rect 5871 25426 5877 25444
rect 5983 25426 5989 25444
rect 5923 25374 5937 25380
rect 5871 25368 5989 25374
rect 6148 26720 6266 26726
rect 6200 26668 6214 26720
rect 6148 26651 6266 26668
rect 6200 26599 6214 26651
rect 6148 26582 6266 26599
rect 6200 26530 6214 26582
rect 6148 26513 6266 26530
rect 6200 26461 6214 26513
rect 6148 26444 6266 26461
rect 6200 26422 6214 26444
rect 6148 26375 6154 26392
rect 6260 26375 6266 26392
rect 6148 26306 6154 26323
rect 6260 26306 6266 26323
rect 6148 26236 6154 26254
rect 6260 26236 6266 26254
rect 6148 26166 6154 26184
rect 6260 26166 6266 26184
rect 6148 25380 6154 26114
rect 6260 25380 6266 26114
rect 6148 25368 6266 25380
rect 6425 26714 6543 26726
rect 6425 26680 6431 26714
rect 6465 26680 6503 26714
rect 6537 26680 6543 26714
rect 6425 26641 6543 26680
rect 6425 26607 6431 26641
rect 6465 26607 6503 26641
rect 6537 26607 6543 26641
rect 6425 26568 6543 26607
rect 6425 26534 6431 26568
rect 6465 26534 6503 26568
rect 6537 26534 6543 26568
rect 6425 26495 6543 26534
rect 6425 26461 6431 26495
rect 6465 26461 6503 26495
rect 6537 26461 6543 26495
rect 6425 26422 6543 26461
rect 6425 25982 6431 26422
rect 6537 25982 6543 26422
rect 6425 25913 6431 25930
rect 6537 25913 6543 25930
rect 6425 25844 6431 25861
rect 6537 25844 6543 25861
rect 6425 25775 6431 25792
rect 6537 25775 6543 25792
rect 6425 25706 6431 25723
rect 6537 25706 6543 25723
rect 6425 25636 6431 25654
rect 6537 25636 6543 25654
rect 6425 25566 6431 25584
rect 6537 25566 6543 25584
rect 6425 25496 6431 25514
rect 6537 25496 6543 25514
rect 6425 25426 6431 25444
rect 6537 25426 6543 25444
rect 6477 25374 6491 25380
rect 6425 25368 6543 25374
rect 6702 26720 6820 26726
rect 6754 26668 6768 26720
rect 6702 26651 6820 26668
rect 6754 26599 6768 26651
rect 6702 26582 6820 26599
rect 6754 26530 6768 26582
rect 6702 26513 6820 26530
rect 6754 26461 6768 26513
rect 6702 26444 6820 26461
rect 6754 26422 6768 26444
rect 6702 26375 6708 26392
rect 6814 26375 6820 26392
rect 6702 26306 6708 26323
rect 6814 26306 6820 26323
rect 6702 26236 6708 26254
rect 6814 26236 6820 26254
rect 6702 26166 6708 26184
rect 6814 26166 6820 26184
rect 6702 25380 6708 26114
rect 6814 25380 6820 26114
rect 6702 25368 6820 25380
rect 6979 26714 7097 26726
rect 6979 26680 6985 26714
rect 7019 26680 7057 26714
rect 7091 26680 7097 26714
rect 6979 26641 7097 26680
rect 6979 26607 6985 26641
rect 7019 26607 7057 26641
rect 7091 26607 7097 26641
rect 6979 26568 7097 26607
rect 6979 26534 6985 26568
rect 7019 26534 7057 26568
rect 7091 26534 7097 26568
rect 6979 26495 7097 26534
rect 6979 26461 6985 26495
rect 7019 26461 7057 26495
rect 7091 26461 7097 26495
rect 6979 26422 7097 26461
rect 6979 25982 6985 26422
rect 7091 25982 7097 26422
rect 6979 25913 6985 25930
rect 7091 25913 7097 25930
rect 6979 25844 6985 25861
rect 7091 25844 7097 25861
rect 6979 25775 6985 25792
rect 7091 25775 7097 25792
rect 6979 25706 6985 25723
rect 7091 25706 7097 25723
rect 6979 25636 6985 25654
rect 7091 25636 7097 25654
rect 6979 25566 6985 25584
rect 7091 25566 7097 25584
rect 6979 25496 6985 25514
rect 7091 25496 7097 25514
rect 6979 25426 6985 25444
rect 7091 25426 7097 25444
rect 7031 25374 7045 25380
rect 6979 25368 7097 25374
rect 7256 26720 7374 26726
rect 7308 26668 7322 26720
rect 7256 26651 7374 26668
rect 7308 26599 7322 26651
rect 7256 26582 7374 26599
rect 7308 26530 7322 26582
rect 7256 26513 7374 26530
rect 7308 26461 7322 26513
rect 7256 26444 7374 26461
rect 7308 26422 7322 26444
rect 7256 26375 7262 26392
rect 7368 26375 7374 26392
rect 7256 26306 7262 26323
rect 7368 26306 7374 26323
rect 7256 26236 7262 26254
rect 7368 26236 7374 26254
rect 7256 26166 7262 26184
rect 7368 26166 7374 26184
rect 7256 25380 7262 26114
rect 7368 25380 7374 26114
rect 7256 25368 7374 25380
rect 7533 26714 7651 26726
rect 7533 26680 7539 26714
rect 7573 26680 7611 26714
rect 7645 26680 7651 26714
rect 7533 26641 7651 26680
rect 7533 26607 7539 26641
rect 7573 26607 7611 26641
rect 7645 26607 7651 26641
rect 7533 26568 7651 26607
rect 7533 26534 7539 26568
rect 7573 26534 7611 26568
rect 7645 26534 7651 26568
rect 7533 26495 7651 26534
rect 7533 26461 7539 26495
rect 7573 26461 7611 26495
rect 7645 26461 7651 26495
rect 7533 26422 7651 26461
rect 7533 25982 7539 26422
rect 7645 25982 7651 26422
rect 7533 25913 7539 25930
rect 7645 25913 7651 25930
rect 7533 25844 7539 25861
rect 7645 25844 7651 25861
rect 7533 25775 7539 25792
rect 7645 25775 7651 25792
rect 7533 25706 7539 25723
rect 7645 25706 7651 25723
rect 7533 25636 7539 25654
rect 7645 25636 7651 25654
rect 7533 25566 7539 25584
rect 7645 25566 7651 25584
rect 7533 25496 7539 25514
rect 7645 25496 7651 25514
rect 7533 25426 7539 25444
rect 7645 25426 7651 25444
rect 7585 25374 7599 25380
rect 7533 25368 7651 25374
rect 7810 26720 7928 26726
rect 7862 26668 7876 26720
rect 7810 26651 7928 26668
rect 7862 26599 7876 26651
rect 7810 26582 7928 26599
rect 7862 26530 7876 26582
rect 7810 26513 7928 26530
rect 7862 26461 7876 26513
rect 7810 26444 7928 26461
rect 7862 26422 7876 26444
rect 7810 26375 7816 26392
rect 7922 26375 7928 26392
rect 7810 26306 7816 26323
rect 7922 26306 7928 26323
rect 7810 26236 7816 26254
rect 7922 26236 7928 26254
rect 7810 26166 7816 26184
rect 7922 26166 7928 26184
rect 7810 25380 7816 26114
rect 7922 25380 7928 26114
rect 7810 25368 7928 25380
rect 8044 26724 8184 26733
rect 8218 26724 8224 26757
rect 8044 26672 8047 26724
rect 8099 26672 8169 26724
rect 8221 26672 8224 26724
rect 8044 26661 8050 26672
rect 8084 26661 8184 26672
rect 8044 26655 8184 26661
rect 8218 26655 8224 26672
rect 8044 26603 8047 26655
rect 8099 26603 8169 26655
rect 8221 26603 8224 26655
rect 8044 26589 8050 26603
rect 8084 26589 8184 26603
rect 8044 26586 8184 26589
rect 8218 26586 8224 26603
rect 8044 26534 8047 26586
rect 8099 26534 8169 26586
rect 8221 26534 8224 26586
rect 8044 26517 8050 26534
rect 8084 26517 8184 26534
rect 8218 26517 8224 26534
rect 8044 26465 8047 26517
rect 8099 26465 8169 26517
rect 8221 26465 8224 26517
rect 8044 26448 8050 26465
rect 8084 26448 8184 26465
rect 8218 26448 8224 26465
rect 8044 26396 8047 26448
rect 8099 26396 8169 26448
rect 8221 26396 8224 26448
rect 8044 26378 8050 26396
rect 8084 26378 8184 26396
rect 8218 26378 8224 26396
rect 8044 26326 8047 26378
rect 8099 26326 8169 26378
rect 8221 26326 8224 26378
rect 8044 26308 8050 26326
rect 8084 26325 8224 26326
rect 8084 26308 8184 26325
rect 8218 26308 8224 26325
rect 8044 26256 8047 26308
rect 8099 26256 8169 26308
rect 8221 26256 8224 26308
rect 8044 26238 8050 26256
rect 8084 26253 8224 26256
rect 8084 26238 8184 26253
rect 8218 26238 8224 26253
rect 8044 26186 8047 26238
rect 8099 26186 8169 26238
rect 8221 26186 8224 26238
rect 8044 26168 8050 26186
rect 8084 26181 8224 26186
rect 8084 26168 8184 26181
rect 8218 26168 8224 26181
rect 8044 26116 8047 26168
rect 8099 26116 8169 26168
rect 8221 26116 8224 26168
rect 8044 26085 8050 26116
rect 8084 26109 8224 26116
rect 8084 26085 8184 26109
rect 8044 26075 8184 26085
rect 8218 26075 8224 26109
rect 8044 26047 8224 26075
rect 8044 26013 8050 26047
rect 8084 26037 8224 26047
rect 8084 26013 8184 26037
rect 8044 26003 8184 26013
rect 8218 26003 8224 26037
rect 8044 25975 8224 26003
rect 8044 25941 8050 25975
rect 8084 25965 8224 25975
rect 8084 25941 8184 25965
rect 8044 25931 8184 25941
rect 8218 25931 8224 25965
rect 8044 25903 8224 25931
rect 8044 25869 8050 25903
rect 8084 25893 8224 25903
rect 8084 25869 8184 25893
rect 8044 25859 8184 25869
rect 8218 25859 8224 25893
rect 8044 25831 8224 25859
rect 8044 25797 8050 25831
rect 8084 25821 8224 25831
rect 8084 25797 8184 25821
rect 8044 25787 8184 25797
rect 8218 25787 8224 25821
rect 8044 25759 8224 25787
rect 8044 25725 8050 25759
rect 8084 25749 8224 25759
rect 8084 25725 8184 25749
rect 8044 25715 8184 25725
rect 8218 25715 8224 25749
rect 8044 25687 8224 25715
rect 8044 25653 8050 25687
rect 8084 25677 8224 25687
rect 8084 25653 8184 25677
rect 8044 25643 8184 25653
rect 8218 25643 8224 25677
rect 8044 25615 8224 25643
rect 8044 25581 8050 25615
rect 8084 25605 8224 25615
rect 8084 25581 8184 25605
rect 8044 25571 8184 25581
rect 8218 25571 8224 25605
rect 8044 25543 8224 25571
rect 8044 25509 8050 25543
rect 8084 25533 8224 25543
rect 8084 25509 8184 25533
rect 8044 25499 8184 25509
rect 8218 25499 8224 25533
rect 8044 25471 8224 25499
rect 8044 25437 8050 25471
rect 8084 25461 8224 25471
rect 8084 25437 8184 25461
rect 8044 25427 8184 25437
rect 8218 25427 8224 25461
rect 8044 25399 8224 25427
rect 8044 25365 8050 25399
rect 8084 25389 8224 25399
rect 8084 25365 8184 25389
rect 8044 25355 8184 25365
rect 8218 25355 8224 25389
rect 8044 25327 8224 25355
rect 8044 25293 8050 25327
rect 8084 25317 8224 25327
rect 8084 25293 8184 25317
rect 8044 25283 8184 25293
rect 8218 25283 8224 25317
rect 8044 25255 8224 25283
rect 8044 25221 8050 25255
rect 8084 25245 8224 25255
rect 8084 25221 8184 25245
rect 8044 25211 8184 25221
rect 8218 25211 8224 25245
tri 4928 25183 4944 25199 sw
rect 8044 25183 8224 25211
rect 4773 25167 4944 25183
tri 4944 25167 4960 25183 sw
rect 4773 25112 7729 25167
rect 4773 25078 5251 25112
rect 5285 25078 5325 25112
rect 5359 25078 5399 25112
rect 5433 25078 5473 25112
rect 5507 25078 5547 25112
rect 5581 25078 5621 25112
rect 5655 25078 5695 25112
rect 5729 25078 5769 25112
rect 5803 25078 5843 25112
rect 5877 25078 5917 25112
rect 5951 25078 5991 25112
rect 6025 25078 6065 25112
rect 6099 25078 6139 25112
rect 6173 25078 6213 25112
rect 6247 25078 6287 25112
rect 6321 25078 6361 25112
rect 6395 25078 6435 25112
rect 6469 25078 6509 25112
rect 6543 25078 6583 25112
rect 6617 25078 6657 25112
rect 6691 25078 6731 25112
rect 6765 25078 6805 25112
rect 6839 25078 6879 25112
rect 6913 25078 6953 25112
rect 6987 25078 7026 25112
rect 7060 25078 7099 25112
rect 7133 25078 7172 25112
rect 7206 25078 7245 25112
rect 7279 25078 7318 25112
rect 7352 25078 7391 25112
rect 7425 25078 7464 25112
rect 7498 25078 7537 25112
rect 7571 25078 7610 25112
rect 7644 25078 7683 25112
rect 7717 25078 7729 25112
rect 4773 25047 7729 25078
rect 8044 25149 8050 25183
rect 8084 25173 8224 25183
rect 8084 25149 8184 25173
rect 8044 25139 8184 25149
rect 8218 25139 8224 25173
rect 8044 25111 8224 25139
rect 8044 25077 8050 25111
rect 8084 25101 8224 25111
rect 8084 25077 8184 25101
rect 8044 25067 8184 25077
rect 8218 25067 8224 25101
rect 4773 25039 5016 25047
tri 5016 25039 5024 25047 nw
rect 8044 25039 8224 25067
rect 4773 25005 4982 25039
tri 4982 25005 5016 25039 nw
rect 8044 25005 8050 25039
rect 8084 25029 8224 25039
rect 8084 25005 8184 25029
rect 4773 24995 4972 25005
tri 4972 24995 4982 25005 nw
rect 8044 24995 8184 25005
rect 8218 24995 8224 25029
rect 4773 24967 4944 24995
tri 4944 24967 4972 24995 nw
rect 8044 24967 8224 24995
rect 4773 23195 4928 24967
tri 4928 24951 4944 24967 nw
rect 8044 24933 8050 24967
rect 8084 24957 8224 24967
rect 8084 24933 8184 24957
rect 8044 24923 8184 24933
rect 8218 24923 8224 24957
rect 8044 24895 8224 24923
rect 8044 24861 8050 24895
rect 8084 24885 8224 24895
rect 8084 24861 8184 24885
rect 8044 24851 8184 24861
rect 8218 24851 8224 24885
rect 8044 24823 8224 24851
rect 8044 24789 8050 24823
rect 8084 24813 8224 24823
rect 8084 24789 8184 24813
rect 8044 24779 8184 24789
rect 8218 24779 8224 24813
rect 8044 24751 8224 24779
rect 5040 24720 5158 24726
rect 5092 24668 5106 24720
rect 5040 24651 5158 24668
rect 5092 24599 5106 24651
rect 5040 24582 5158 24599
rect 5092 24530 5106 24582
rect 5040 24513 5158 24530
rect 5092 24461 5106 24513
rect 5040 24444 5158 24461
rect 5092 24422 5106 24444
rect 5040 24375 5046 24392
rect 5152 24375 5158 24392
rect 5040 24306 5046 24323
rect 5152 24306 5158 24323
rect 5040 24236 5046 24254
rect 5152 24236 5158 24254
rect 5040 24166 5046 24184
rect 5152 24166 5158 24184
rect 5040 23380 5046 24114
rect 5152 23380 5158 24114
rect 5040 23368 5158 23380
rect 5317 24714 5435 24726
rect 5317 24680 5323 24714
rect 5357 24680 5395 24714
rect 5429 24680 5435 24714
rect 5317 24641 5435 24680
rect 5317 24607 5323 24641
rect 5357 24607 5395 24641
rect 5429 24607 5435 24641
rect 5317 24568 5435 24607
rect 5317 24534 5323 24568
rect 5357 24534 5395 24568
rect 5429 24534 5435 24568
rect 5317 24495 5435 24534
rect 5317 24461 5323 24495
rect 5357 24461 5395 24495
rect 5429 24461 5435 24495
rect 5317 24422 5435 24461
rect 5317 23982 5323 24422
rect 5429 23982 5435 24422
rect 5317 23913 5323 23930
rect 5429 23913 5435 23930
rect 5317 23844 5323 23861
rect 5429 23844 5435 23861
rect 5317 23775 5323 23792
rect 5429 23775 5435 23792
rect 5317 23706 5323 23723
rect 5429 23706 5435 23723
rect 5317 23636 5323 23654
rect 5429 23636 5435 23654
rect 5317 23566 5323 23584
rect 5429 23566 5435 23584
rect 5317 23496 5323 23514
rect 5429 23496 5435 23514
rect 5317 23426 5323 23444
rect 5429 23426 5435 23444
rect 5369 23374 5383 23380
rect 5317 23368 5435 23374
rect 5594 24720 5712 24726
rect 5646 24668 5660 24720
rect 5594 24651 5712 24668
rect 5646 24599 5660 24651
rect 5594 24582 5712 24599
rect 5646 24530 5660 24582
rect 5594 24513 5712 24530
rect 5646 24461 5660 24513
rect 5594 24444 5712 24461
rect 5646 24422 5660 24444
rect 5594 24375 5600 24392
rect 5706 24375 5712 24392
rect 5594 24306 5600 24323
rect 5706 24306 5712 24323
rect 5594 24236 5600 24254
rect 5706 24236 5712 24254
rect 5594 24166 5600 24184
rect 5706 24166 5712 24184
rect 5594 23380 5600 24114
rect 5706 23380 5712 24114
rect 5594 23368 5712 23380
rect 5871 24714 5989 24726
rect 5871 24680 5877 24714
rect 5911 24680 5949 24714
rect 5983 24680 5989 24714
rect 5871 24641 5989 24680
rect 5871 24607 5877 24641
rect 5911 24607 5949 24641
rect 5983 24607 5989 24641
rect 5871 24568 5989 24607
rect 5871 24534 5877 24568
rect 5911 24534 5949 24568
rect 5983 24534 5989 24568
rect 5871 24495 5989 24534
rect 5871 24461 5877 24495
rect 5911 24461 5949 24495
rect 5983 24461 5989 24495
rect 5871 24422 5989 24461
rect 5871 23982 5877 24422
rect 5983 23982 5989 24422
rect 5871 23913 5877 23930
rect 5983 23913 5989 23930
rect 5871 23844 5877 23861
rect 5983 23844 5989 23861
rect 5871 23775 5877 23792
rect 5983 23775 5989 23792
rect 5871 23706 5877 23723
rect 5983 23706 5989 23723
rect 5871 23636 5877 23654
rect 5983 23636 5989 23654
rect 5871 23566 5877 23584
rect 5983 23566 5989 23584
rect 5871 23496 5877 23514
rect 5983 23496 5989 23514
rect 5871 23426 5877 23444
rect 5983 23426 5989 23444
rect 5923 23374 5937 23380
rect 5871 23368 5989 23374
rect 6148 24720 6266 24726
rect 6200 24668 6214 24720
rect 6148 24651 6266 24668
rect 6200 24599 6214 24651
rect 6148 24582 6266 24599
rect 6200 24530 6214 24582
rect 6148 24513 6266 24530
rect 6200 24461 6214 24513
rect 6148 24444 6266 24461
rect 6200 24422 6214 24444
rect 6148 24375 6154 24392
rect 6260 24375 6266 24392
rect 6148 24306 6154 24323
rect 6260 24306 6266 24323
rect 6148 24236 6154 24254
rect 6260 24236 6266 24254
rect 6148 24166 6154 24184
rect 6260 24166 6266 24184
rect 6148 23380 6154 24114
rect 6260 23380 6266 24114
rect 6148 23368 6266 23380
rect 6425 24714 6543 24726
rect 6425 24680 6431 24714
rect 6465 24680 6503 24714
rect 6537 24680 6543 24714
rect 6425 24641 6543 24680
rect 6425 24607 6431 24641
rect 6465 24607 6503 24641
rect 6537 24607 6543 24641
rect 6425 24568 6543 24607
rect 6425 24534 6431 24568
rect 6465 24534 6503 24568
rect 6537 24534 6543 24568
rect 6425 24495 6543 24534
rect 6425 24461 6431 24495
rect 6465 24461 6503 24495
rect 6537 24461 6543 24495
rect 6425 24422 6543 24461
rect 6425 23982 6431 24422
rect 6537 23982 6543 24422
rect 6425 23913 6431 23930
rect 6537 23913 6543 23930
rect 6425 23844 6431 23861
rect 6537 23844 6543 23861
rect 6425 23775 6431 23792
rect 6537 23775 6543 23792
rect 6425 23706 6431 23723
rect 6537 23706 6543 23723
rect 6425 23636 6431 23654
rect 6537 23636 6543 23654
rect 6425 23566 6431 23584
rect 6537 23566 6543 23584
rect 6425 23496 6431 23514
rect 6537 23496 6543 23514
rect 6425 23426 6431 23444
rect 6537 23426 6543 23444
rect 6477 23374 6491 23380
rect 6425 23368 6543 23374
rect 6702 24720 6820 24726
rect 6754 24668 6768 24720
rect 6702 24651 6820 24668
rect 6754 24599 6768 24651
rect 6702 24582 6820 24599
rect 6754 24530 6768 24582
rect 6702 24513 6820 24530
rect 6754 24461 6768 24513
rect 6702 24444 6820 24461
rect 6754 24422 6768 24444
rect 6702 24375 6708 24392
rect 6814 24375 6820 24392
rect 6702 24306 6708 24323
rect 6814 24306 6820 24323
rect 6702 24236 6708 24254
rect 6814 24236 6820 24254
rect 6702 24166 6708 24184
rect 6814 24166 6820 24184
rect 6702 23380 6708 24114
rect 6814 23380 6820 24114
rect 6702 23368 6820 23380
rect 6979 24714 7097 24726
rect 6979 24680 6985 24714
rect 7019 24680 7057 24714
rect 7091 24680 7097 24714
rect 6979 24641 7097 24680
rect 6979 24607 6985 24641
rect 7019 24607 7057 24641
rect 7091 24607 7097 24641
rect 6979 24568 7097 24607
rect 6979 24534 6985 24568
rect 7019 24534 7057 24568
rect 7091 24534 7097 24568
rect 6979 24495 7097 24534
rect 6979 24461 6985 24495
rect 7019 24461 7057 24495
rect 7091 24461 7097 24495
rect 6979 24422 7097 24461
rect 6979 23982 6985 24422
rect 7091 23982 7097 24422
rect 6979 23913 6985 23930
rect 7091 23913 7097 23930
rect 6979 23844 6985 23861
rect 7091 23844 7097 23861
rect 6979 23775 6985 23792
rect 7091 23775 7097 23792
rect 6979 23706 6985 23723
rect 7091 23706 7097 23723
rect 6979 23636 6985 23654
rect 7091 23636 7097 23654
rect 6979 23566 6985 23584
rect 7091 23566 7097 23584
rect 6979 23496 6985 23514
rect 7091 23496 7097 23514
rect 6979 23426 6985 23444
rect 7091 23426 7097 23444
rect 7031 23374 7045 23380
rect 6979 23368 7097 23374
rect 7256 24720 7374 24726
rect 7308 24668 7322 24720
rect 7256 24651 7374 24668
rect 7308 24599 7322 24651
rect 7256 24582 7374 24599
rect 7308 24530 7322 24582
rect 7256 24513 7374 24530
rect 7308 24461 7322 24513
rect 7256 24444 7374 24461
rect 7308 24422 7322 24444
rect 7256 24375 7262 24392
rect 7368 24375 7374 24392
rect 7256 24306 7262 24323
rect 7368 24306 7374 24323
rect 7256 24236 7262 24254
rect 7368 24236 7374 24254
rect 7256 24166 7262 24184
rect 7368 24166 7374 24184
rect 7256 23380 7262 24114
rect 7368 23380 7374 24114
rect 7256 23368 7374 23380
rect 7533 24714 7651 24726
rect 7533 24680 7539 24714
rect 7573 24680 7611 24714
rect 7645 24680 7651 24714
rect 7533 24641 7651 24680
rect 7533 24607 7539 24641
rect 7573 24607 7611 24641
rect 7645 24607 7651 24641
rect 7533 24568 7651 24607
rect 7533 24534 7539 24568
rect 7573 24534 7611 24568
rect 7645 24534 7651 24568
rect 7533 24495 7651 24534
rect 7533 24461 7539 24495
rect 7573 24461 7611 24495
rect 7645 24461 7651 24495
rect 7533 24422 7651 24461
rect 7533 23982 7539 24422
rect 7645 23982 7651 24422
rect 7533 23913 7539 23930
rect 7645 23913 7651 23930
rect 7533 23844 7539 23861
rect 7645 23844 7651 23861
rect 7533 23775 7539 23792
rect 7645 23775 7651 23792
rect 7533 23706 7539 23723
rect 7645 23706 7651 23723
rect 7533 23636 7539 23654
rect 7645 23636 7651 23654
rect 7533 23566 7539 23584
rect 7645 23566 7651 23584
rect 7533 23496 7539 23514
rect 7645 23496 7651 23514
rect 7533 23426 7539 23444
rect 7645 23426 7651 23444
rect 7585 23374 7599 23380
rect 7533 23368 7651 23374
rect 7810 24720 7928 24726
rect 7862 24668 7876 24720
rect 7810 24651 7928 24668
rect 7862 24599 7876 24651
rect 7810 24582 7928 24599
rect 7862 24530 7876 24582
rect 7810 24513 7928 24530
rect 7862 24461 7876 24513
rect 7810 24444 7928 24461
rect 7862 24422 7876 24444
rect 7810 24375 7816 24392
rect 7922 24375 7928 24392
rect 7810 24306 7816 24323
rect 7922 24306 7928 24323
rect 7810 24236 7816 24254
rect 7922 24236 7928 24254
rect 7810 24166 7816 24184
rect 7922 24166 7928 24184
rect 7810 23380 7816 24114
rect 7922 23380 7928 24114
rect 7810 23368 7928 23380
rect 8044 24724 8050 24751
rect 8084 24741 8224 24751
rect 8084 24724 8184 24741
rect 8218 24724 8224 24741
rect 8044 24672 8047 24724
rect 8099 24672 8169 24724
rect 8221 24672 8224 24724
rect 8044 24655 8050 24672
rect 8084 24669 8224 24672
rect 8084 24655 8184 24669
rect 8218 24655 8224 24669
rect 8044 24603 8047 24655
rect 8099 24603 8169 24655
rect 8221 24603 8224 24655
rect 8044 24586 8050 24603
rect 8084 24597 8224 24603
rect 8084 24586 8184 24597
rect 8218 24586 8224 24597
rect 8044 24534 8047 24586
rect 8099 24534 8169 24586
rect 8221 24534 8224 24586
rect 8044 24517 8050 24534
rect 8084 24525 8224 24534
rect 8084 24517 8184 24525
rect 8218 24517 8224 24525
rect 8044 24465 8047 24517
rect 8099 24465 8169 24517
rect 8221 24465 8224 24517
rect 8044 24463 8224 24465
rect 8044 24448 8050 24463
rect 8084 24453 8224 24463
rect 8084 24448 8184 24453
rect 8218 24448 8224 24453
rect 8044 24396 8047 24448
rect 8099 24396 8169 24448
rect 8221 24396 8224 24448
rect 8044 24391 8224 24396
rect 8044 24378 8050 24391
rect 8084 24381 8224 24391
rect 8084 24378 8184 24381
rect 8218 24378 8224 24381
rect 8044 24326 8047 24378
rect 8099 24326 8169 24378
rect 8221 24326 8224 24378
rect 8044 24319 8224 24326
rect 8044 24308 8050 24319
rect 8084 24309 8224 24319
rect 8084 24308 8184 24309
rect 8218 24308 8224 24309
rect 8044 24256 8047 24308
rect 8099 24256 8169 24308
rect 8221 24256 8224 24308
rect 8044 24247 8224 24256
rect 8044 24238 8050 24247
rect 8084 24238 8224 24247
rect 8044 24186 8047 24238
rect 8099 24186 8169 24238
rect 8221 24186 8224 24238
rect 8044 24175 8224 24186
rect 8044 24168 8050 24175
rect 8084 24168 8224 24175
rect 8044 24116 8047 24168
rect 8099 24116 8169 24168
rect 8221 24116 8224 24168
rect 8044 24103 8224 24116
rect 8044 24069 8050 24103
rect 8084 24093 8224 24103
rect 8084 24069 8184 24093
rect 8044 24059 8184 24069
rect 8218 24059 8224 24093
rect 8044 24031 8224 24059
rect 8044 23997 8050 24031
rect 8084 24021 8224 24031
rect 8084 23997 8184 24021
rect 8044 23987 8184 23997
rect 8218 23987 8224 24021
rect 8044 23959 8224 23987
rect 8044 23925 8050 23959
rect 8084 23949 8224 23959
rect 8084 23925 8184 23949
rect 8044 23915 8184 23925
rect 8218 23915 8224 23949
rect 8044 23887 8224 23915
rect 8044 23853 8050 23887
rect 8084 23877 8224 23887
rect 8084 23853 8184 23877
rect 8044 23843 8184 23853
rect 8218 23843 8224 23877
rect 8044 23815 8224 23843
rect 8044 23781 8050 23815
rect 8084 23805 8224 23815
rect 8084 23781 8184 23805
rect 8044 23771 8184 23781
rect 8218 23771 8224 23805
rect 8044 23743 8224 23771
rect 8044 23709 8050 23743
rect 8084 23733 8224 23743
rect 8084 23709 8184 23733
rect 8044 23699 8184 23709
rect 8218 23699 8224 23733
rect 8044 23671 8224 23699
rect 8044 23637 8050 23671
rect 8084 23661 8224 23671
rect 8084 23637 8184 23661
rect 8044 23627 8184 23637
rect 8218 23627 8224 23661
rect 8044 23599 8224 23627
rect 8044 23565 8050 23599
rect 8084 23589 8224 23599
rect 8084 23565 8184 23589
rect 8044 23555 8184 23565
rect 8218 23555 8224 23589
rect 8044 23527 8224 23555
rect 8044 23493 8050 23527
rect 8084 23517 8224 23527
rect 8084 23493 8184 23517
rect 8044 23483 8184 23493
rect 8218 23483 8224 23517
rect 8044 23455 8224 23483
rect 8044 23421 8050 23455
rect 8084 23445 8224 23455
rect 8084 23421 8184 23445
rect 8044 23411 8184 23421
rect 8218 23411 8224 23445
rect 8044 23383 8224 23411
rect 8044 23349 8050 23383
rect 8084 23373 8224 23383
rect 8084 23349 8184 23373
rect 8044 23339 8184 23349
rect 8218 23339 8224 23373
rect 8044 23311 8224 23339
rect 8044 23277 8050 23311
rect 8084 23301 8224 23311
rect 8084 23277 8184 23301
rect 8044 23267 8184 23277
rect 8218 23267 8224 23301
rect 8044 23239 8224 23267
rect 8044 23205 8050 23239
rect 8084 23229 8224 23239
rect 8084 23205 8184 23229
tri 4928 23195 4932 23199 sw
rect 8044 23195 8184 23205
rect 8218 23195 8224 23229
rect 4773 23167 4932 23195
tri 4932 23167 4960 23195 sw
rect 8044 23167 8224 23195
rect 4773 23124 7729 23167
rect 4773 23090 5251 23124
rect 5285 23090 5325 23124
rect 5359 23090 5399 23124
rect 5433 23090 5473 23124
rect 5507 23090 5547 23124
rect 5581 23090 5621 23124
rect 5655 23090 5695 23124
rect 5729 23090 5769 23124
rect 5803 23090 5843 23124
rect 5877 23090 5917 23124
rect 5951 23090 5991 23124
rect 6025 23090 6065 23124
rect 6099 23090 6139 23124
rect 6173 23090 6213 23124
rect 6247 23090 6287 23124
rect 6321 23090 6361 23124
rect 6395 23090 6435 23124
rect 6469 23090 6509 23124
rect 6543 23090 6583 23124
rect 6617 23090 6657 23124
rect 6691 23090 6731 23124
rect 6765 23090 6805 23124
rect 6839 23090 6879 23124
rect 6913 23090 6953 23124
rect 6987 23090 7026 23124
rect 7060 23090 7099 23124
rect 7133 23090 7172 23124
rect 7206 23090 7245 23124
rect 7279 23090 7318 23124
rect 7352 23090 7391 23124
rect 7425 23090 7464 23124
rect 7498 23090 7537 23124
rect 7571 23090 7610 23124
rect 7644 23090 7683 23124
rect 7717 23090 7729 23124
rect 4773 23047 7729 23090
rect 8044 23133 8050 23167
rect 8084 23157 8224 23167
rect 8084 23133 8184 23157
rect 8044 23123 8184 23133
rect 8218 23123 8224 23157
rect 8044 23095 8224 23123
rect 8044 23061 8050 23095
rect 8084 23085 8224 23095
rect 8084 23061 8184 23085
rect 8044 23051 8184 23061
rect 8218 23051 8224 23085
rect 4773 23023 4962 23047
tri 4962 23023 4986 23047 nw
rect 8044 23023 8224 23051
rect 4773 21151 4928 23023
tri 4928 22989 4962 23023 nw
rect 8044 22989 8050 23023
rect 8084 23013 8224 23023
rect 8084 22989 8184 23013
rect 8044 22979 8184 22989
rect 8218 22979 8224 23013
rect 8044 22951 8224 22979
rect 8044 22917 8050 22951
rect 8084 22941 8224 22951
rect 8084 22917 8184 22941
rect 8044 22907 8184 22917
rect 8218 22907 8224 22941
rect 8044 22879 8224 22907
rect 8044 22845 8050 22879
rect 8084 22869 8224 22879
rect 8084 22845 8184 22869
rect 8044 22835 8184 22845
rect 8218 22835 8224 22869
rect 8044 22807 8224 22835
rect 8044 22773 8050 22807
rect 8084 22797 8224 22807
rect 8084 22773 8184 22797
rect 8044 22763 8184 22773
rect 8218 22763 8224 22797
rect 8044 22735 8224 22763
rect 5040 22720 5158 22726
rect 5092 22668 5106 22720
rect 5040 22651 5158 22668
rect 5092 22599 5106 22651
rect 5040 22582 5158 22599
rect 5092 22530 5106 22582
rect 5040 22513 5158 22530
rect 5092 22461 5106 22513
rect 5040 22444 5158 22461
rect 5092 22422 5106 22444
rect 5040 22375 5046 22392
rect 5152 22375 5158 22392
rect 5040 22306 5046 22323
rect 5152 22306 5158 22323
rect 5040 22236 5046 22254
rect 5152 22236 5158 22254
rect 5040 22166 5046 22184
rect 5152 22166 5158 22184
rect 5040 21380 5046 22114
rect 5152 21380 5158 22114
rect 5040 21368 5158 21380
rect 5317 22714 5435 22726
rect 5317 22680 5323 22714
rect 5357 22680 5395 22714
rect 5429 22680 5435 22714
rect 5317 22641 5435 22680
rect 5317 22607 5323 22641
rect 5357 22607 5395 22641
rect 5429 22607 5435 22641
rect 5317 22568 5435 22607
rect 5317 22534 5323 22568
rect 5357 22534 5395 22568
rect 5429 22534 5435 22568
rect 5317 22495 5435 22534
rect 5317 22461 5323 22495
rect 5357 22461 5395 22495
rect 5429 22461 5435 22495
rect 5317 22422 5435 22461
rect 5317 21982 5323 22422
rect 5429 21982 5435 22422
rect 5317 21913 5323 21930
rect 5429 21913 5435 21930
rect 5317 21844 5323 21861
rect 5429 21844 5435 21861
rect 5317 21775 5323 21792
rect 5429 21775 5435 21792
rect 5317 21706 5323 21723
rect 5429 21706 5435 21723
rect 5317 21636 5323 21654
rect 5429 21636 5435 21654
rect 5317 21566 5323 21584
rect 5429 21566 5435 21584
rect 5317 21496 5323 21514
rect 5429 21496 5435 21514
rect 5317 21426 5323 21444
rect 5429 21426 5435 21444
rect 5369 21374 5383 21380
rect 5317 21368 5435 21374
rect 5594 22720 5712 22726
rect 5646 22668 5660 22720
rect 5594 22651 5712 22668
rect 5646 22599 5660 22651
rect 5594 22582 5712 22599
rect 5646 22530 5660 22582
rect 5594 22513 5712 22530
rect 5646 22461 5660 22513
rect 5594 22444 5712 22461
rect 5646 22422 5660 22444
rect 5594 22375 5600 22392
rect 5706 22375 5712 22392
rect 5594 22306 5600 22323
rect 5706 22306 5712 22323
rect 5594 22236 5600 22254
rect 5706 22236 5712 22254
rect 5594 22166 5600 22184
rect 5706 22166 5712 22184
rect 5594 21380 5600 22114
rect 5706 21380 5712 22114
rect 5594 21368 5712 21380
rect 5871 22714 5989 22726
rect 5871 22680 5877 22714
rect 5911 22680 5949 22714
rect 5983 22680 5989 22714
rect 5871 22641 5989 22680
rect 5871 22607 5877 22641
rect 5911 22607 5949 22641
rect 5983 22607 5989 22641
rect 5871 22568 5989 22607
rect 5871 22534 5877 22568
rect 5911 22534 5949 22568
rect 5983 22534 5989 22568
rect 5871 22495 5989 22534
rect 5871 22461 5877 22495
rect 5911 22461 5949 22495
rect 5983 22461 5989 22495
rect 5871 22422 5989 22461
rect 5871 21982 5877 22422
rect 5983 21982 5989 22422
rect 5871 21913 5877 21930
rect 5983 21913 5989 21930
rect 5871 21844 5877 21861
rect 5983 21844 5989 21861
rect 5871 21775 5877 21792
rect 5983 21775 5989 21792
rect 5871 21706 5877 21723
rect 5983 21706 5989 21723
rect 5871 21636 5877 21654
rect 5983 21636 5989 21654
rect 5871 21566 5877 21584
rect 5983 21566 5989 21584
rect 5871 21496 5877 21514
rect 5983 21496 5989 21514
rect 5871 21426 5877 21444
rect 5983 21426 5989 21444
rect 5923 21374 5937 21380
rect 5871 21368 5989 21374
rect 6148 22720 6266 22726
rect 6200 22668 6214 22720
rect 6148 22651 6266 22668
rect 6200 22599 6214 22651
rect 6148 22582 6266 22599
rect 6200 22530 6214 22582
rect 6148 22513 6266 22530
rect 6200 22461 6214 22513
rect 6148 22444 6266 22461
rect 6200 22422 6214 22444
rect 6148 22375 6154 22392
rect 6260 22375 6266 22392
rect 6148 22306 6154 22323
rect 6260 22306 6266 22323
rect 6148 22236 6154 22254
rect 6260 22236 6266 22254
rect 6148 22166 6154 22184
rect 6260 22166 6266 22184
rect 6148 21380 6154 22114
rect 6260 21380 6266 22114
rect 6148 21368 6266 21380
rect 6425 22714 6543 22726
rect 6425 22680 6431 22714
rect 6465 22680 6503 22714
rect 6537 22680 6543 22714
rect 6425 22641 6543 22680
rect 6425 22607 6431 22641
rect 6465 22607 6503 22641
rect 6537 22607 6543 22641
rect 6425 22568 6543 22607
rect 6425 22534 6431 22568
rect 6465 22534 6503 22568
rect 6537 22534 6543 22568
rect 6425 22495 6543 22534
rect 6425 22461 6431 22495
rect 6465 22461 6503 22495
rect 6537 22461 6543 22495
rect 6425 22422 6543 22461
rect 6425 21982 6431 22422
rect 6537 21982 6543 22422
rect 6425 21913 6431 21930
rect 6537 21913 6543 21930
rect 6425 21844 6431 21861
rect 6537 21844 6543 21861
rect 6425 21775 6431 21792
rect 6537 21775 6543 21792
rect 6425 21706 6431 21723
rect 6537 21706 6543 21723
rect 6425 21636 6431 21654
rect 6537 21636 6543 21654
rect 6425 21566 6431 21584
rect 6537 21566 6543 21584
rect 6425 21496 6431 21514
rect 6537 21496 6543 21514
rect 6425 21426 6431 21444
rect 6537 21426 6543 21444
rect 6477 21374 6491 21380
rect 6425 21368 6543 21374
rect 6702 22720 6820 22726
rect 6754 22668 6768 22720
rect 6702 22651 6820 22668
rect 6754 22599 6768 22651
rect 6702 22582 6820 22599
rect 6754 22530 6768 22582
rect 6702 22513 6820 22530
rect 6754 22461 6768 22513
rect 6702 22444 6820 22461
rect 6754 22422 6768 22444
rect 6702 22375 6708 22392
rect 6814 22375 6820 22392
rect 6702 22306 6708 22323
rect 6814 22306 6820 22323
rect 6702 22236 6708 22254
rect 6814 22236 6820 22254
rect 6702 22166 6708 22184
rect 6814 22166 6820 22184
rect 6702 21380 6708 22114
rect 6814 21380 6820 22114
rect 6702 21368 6820 21380
rect 6979 22714 7097 22726
rect 6979 22680 6985 22714
rect 7019 22680 7057 22714
rect 7091 22680 7097 22714
rect 6979 22641 7097 22680
rect 6979 22607 6985 22641
rect 7019 22607 7057 22641
rect 7091 22607 7097 22641
rect 6979 22568 7097 22607
rect 6979 22534 6985 22568
rect 7019 22534 7057 22568
rect 7091 22534 7097 22568
rect 6979 22495 7097 22534
rect 6979 22461 6985 22495
rect 7019 22461 7057 22495
rect 7091 22461 7097 22495
rect 6979 22422 7097 22461
rect 6979 21982 6985 22422
rect 7091 21982 7097 22422
rect 6979 21913 6985 21930
rect 7091 21913 7097 21930
rect 6979 21844 6985 21861
rect 7091 21844 7097 21861
rect 6979 21775 6985 21792
rect 7091 21775 7097 21792
rect 6979 21706 6985 21723
rect 7091 21706 7097 21723
rect 6979 21636 6985 21654
rect 7091 21636 7097 21654
rect 6979 21566 6985 21584
rect 7091 21566 7097 21584
rect 6979 21496 6985 21514
rect 7091 21496 7097 21514
rect 6979 21426 6985 21444
rect 7091 21426 7097 21444
rect 7031 21374 7045 21380
rect 6979 21368 7097 21374
rect 7256 22720 7374 22726
rect 7308 22668 7322 22720
rect 7256 22651 7374 22668
rect 7308 22599 7322 22651
rect 7256 22582 7374 22599
rect 7308 22530 7322 22582
rect 7256 22513 7374 22530
rect 7308 22461 7322 22513
rect 7256 22444 7374 22461
rect 7308 22422 7322 22444
rect 7256 22375 7262 22392
rect 7368 22375 7374 22392
rect 7256 22306 7262 22323
rect 7368 22306 7374 22323
rect 7256 22236 7262 22254
rect 7368 22236 7374 22254
rect 7256 22166 7262 22184
rect 7368 22166 7374 22184
rect 7256 21380 7262 22114
rect 7368 21380 7374 22114
rect 7256 21368 7374 21380
rect 7533 22714 7651 22726
rect 7533 22680 7539 22714
rect 7573 22680 7611 22714
rect 7645 22680 7651 22714
rect 7533 22641 7651 22680
rect 7533 22607 7539 22641
rect 7573 22607 7611 22641
rect 7645 22607 7651 22641
rect 7533 22568 7651 22607
rect 7533 22534 7539 22568
rect 7573 22534 7611 22568
rect 7645 22534 7651 22568
rect 7533 22495 7651 22534
rect 7533 22461 7539 22495
rect 7573 22461 7611 22495
rect 7645 22461 7651 22495
rect 7533 22422 7651 22461
rect 7533 21982 7539 22422
rect 7645 21982 7651 22422
rect 7533 21913 7539 21930
rect 7645 21913 7651 21930
rect 7533 21844 7539 21861
rect 7645 21844 7651 21861
rect 7533 21775 7539 21792
rect 7645 21775 7651 21792
rect 7533 21706 7539 21723
rect 7645 21706 7651 21723
rect 7533 21636 7539 21654
rect 7645 21636 7651 21654
rect 7533 21566 7539 21584
rect 7645 21566 7651 21584
rect 7533 21496 7539 21514
rect 7645 21496 7651 21514
rect 7533 21426 7539 21444
rect 7645 21426 7651 21444
rect 7585 21374 7599 21380
rect 7533 21368 7651 21374
rect 7810 22720 7928 22726
rect 7862 22668 7876 22720
rect 7810 22651 7928 22668
rect 7862 22599 7876 22651
rect 7810 22582 7928 22599
rect 7862 22530 7876 22582
rect 7810 22513 7928 22530
rect 7862 22461 7876 22513
rect 7810 22444 7928 22461
rect 7862 22422 7876 22444
rect 7810 22375 7816 22392
rect 7922 22375 7928 22392
rect 7810 22306 7816 22323
rect 7922 22306 7928 22323
rect 7810 22236 7816 22254
rect 7922 22236 7928 22254
rect 7810 22166 7816 22184
rect 7922 22166 7928 22184
rect 7810 21380 7816 22114
rect 7922 21380 7928 22114
rect 7810 21368 7928 21380
rect 8044 22724 8050 22735
rect 8084 22725 8224 22735
rect 8084 22724 8184 22725
rect 8218 22724 8224 22725
rect 8044 22672 8047 22724
rect 8099 22672 8169 22724
rect 8221 22672 8224 22724
rect 8044 22663 8224 22672
rect 8044 22655 8050 22663
rect 8084 22655 8224 22663
rect 8044 22603 8047 22655
rect 8099 22603 8169 22655
rect 8221 22603 8224 22655
rect 8044 22591 8224 22603
rect 8044 22586 8050 22591
rect 8084 22586 8224 22591
rect 8044 22534 8047 22586
rect 8099 22534 8169 22586
rect 8221 22534 8224 22586
rect 8044 22519 8224 22534
rect 8044 22517 8050 22519
rect 8084 22517 8224 22519
rect 8044 22465 8047 22517
rect 8099 22465 8169 22517
rect 8221 22465 8224 22517
rect 8044 22448 8224 22465
rect 8044 22396 8047 22448
rect 8099 22396 8169 22448
rect 8221 22396 8224 22448
rect 8044 22378 8224 22396
rect 8044 22326 8047 22378
rect 8099 22326 8169 22378
rect 8221 22326 8224 22378
rect 8044 22308 8224 22326
rect 8044 22256 8047 22308
rect 8099 22256 8169 22308
rect 8221 22256 8224 22308
rect 8044 22238 8224 22256
rect 8044 22186 8047 22238
rect 8099 22186 8169 22238
rect 8221 22186 8224 22238
rect 8044 22168 8224 22186
rect 8044 22116 8047 22168
rect 8099 22116 8169 22168
rect 8221 22116 8224 22168
rect 8044 22115 8184 22116
rect 8218 22115 8224 22116
rect 8044 22087 8224 22115
rect 8044 22053 8050 22087
rect 8084 22077 8224 22087
rect 8084 22053 8184 22077
rect 8044 22043 8184 22053
rect 8218 22043 8224 22077
rect 8044 22015 8224 22043
rect 8044 21981 8050 22015
rect 8084 22005 8224 22015
rect 8084 21981 8184 22005
rect 8044 21971 8184 21981
rect 8218 21971 8224 22005
rect 8044 21943 8224 21971
rect 8044 21909 8050 21943
rect 8084 21933 8224 21943
rect 8084 21909 8184 21933
rect 8044 21899 8184 21909
rect 8218 21899 8224 21933
rect 8044 21871 8224 21899
rect 8044 21837 8050 21871
rect 8084 21861 8224 21871
rect 8084 21837 8184 21861
rect 8044 21827 8184 21837
rect 8218 21827 8224 21861
rect 8044 21799 8224 21827
rect 8044 21765 8050 21799
rect 8084 21789 8224 21799
rect 8084 21765 8184 21789
rect 8044 21755 8184 21765
rect 8218 21755 8224 21789
rect 8044 21727 8224 21755
rect 8044 21693 8050 21727
rect 8084 21717 8224 21727
rect 8084 21693 8184 21717
rect 8044 21683 8184 21693
rect 8218 21683 8224 21717
rect 8044 21655 8224 21683
rect 8044 21621 8050 21655
rect 8084 21645 8224 21655
rect 8084 21621 8184 21645
rect 8044 21611 8184 21621
rect 8218 21611 8224 21645
rect 8044 21583 8224 21611
rect 8044 21549 8050 21583
rect 8084 21573 8224 21583
rect 8084 21549 8184 21573
rect 8044 21539 8184 21549
rect 8218 21539 8224 21573
rect 8044 21511 8224 21539
rect 8044 21477 8050 21511
rect 8084 21501 8224 21511
rect 8084 21477 8184 21501
rect 8044 21467 8184 21477
rect 8218 21467 8224 21501
rect 8044 21439 8224 21467
rect 8044 21405 8050 21439
rect 8084 21429 8224 21439
rect 8084 21405 8184 21429
rect 8044 21395 8184 21405
rect 8218 21395 8224 21429
rect 8044 21367 8224 21395
rect 8044 21333 8050 21367
rect 8084 21357 8224 21367
rect 8084 21333 8184 21357
rect 8044 21323 8184 21333
rect 8218 21323 8224 21357
rect 8044 21295 8224 21323
rect 8044 21261 8050 21295
rect 8084 21285 8224 21295
rect 8084 21261 8184 21285
rect 8044 21251 8184 21261
rect 8218 21251 8224 21285
rect 8044 21223 8224 21251
rect 8044 21189 8050 21223
rect 8084 21213 8224 21223
rect 8084 21189 8184 21213
rect 8044 21179 8184 21189
rect 8218 21179 8224 21213
tri 4928 21151 4940 21163 sw
rect 8044 21151 8224 21179
rect 4773 21131 4940 21151
tri 4940 21131 4960 21151 sw
rect 4773 21083 7729 21131
rect 4773 21049 5251 21083
rect 5285 21049 5326 21083
rect 5360 21049 5401 21083
rect 5435 21049 5476 21083
rect 5510 21049 5551 21083
rect 5585 21049 5626 21083
rect 5660 21049 5701 21083
rect 5735 21049 5776 21083
rect 5810 21049 5851 21083
rect 5885 21049 5926 21083
rect 5960 21049 6001 21083
rect 6035 21049 6076 21083
rect 6110 21049 6151 21083
rect 6185 21049 6225 21083
rect 6259 21049 6299 21083
rect 6333 21049 6373 21083
rect 6407 21049 6447 21083
rect 6481 21049 6521 21083
rect 6555 21049 6595 21083
rect 6629 21049 6669 21083
rect 6703 21049 6743 21083
rect 6777 21049 6817 21083
rect 6851 21049 6891 21083
rect 6925 21049 7729 21083
rect 4773 21011 7729 21049
rect 8044 21117 8050 21151
rect 8084 21141 8224 21151
rect 8084 21117 8184 21141
rect 8044 21107 8184 21117
rect 8218 21107 8224 21141
rect 8044 21079 8224 21107
rect 8044 21045 8050 21079
rect 8084 21069 8224 21079
rect 8084 21045 8184 21069
rect 8044 21035 8184 21045
rect 8218 21035 8224 21069
rect 4773 21007 4978 21011
tri 4978 21007 4982 21011 nw
rect 8044 21007 8224 21035
rect 4773 20973 4944 21007
tri 4944 20973 4978 21007 nw
rect 8044 20973 8050 21007
rect 8084 20997 8224 21007
rect 8084 20973 8184 20997
rect 4773 20963 4934 20973
tri 4934 20963 4944 20973 nw
rect 8044 20963 8184 20973
rect 8218 20963 8224 20997
rect 4773 19173 4928 20963
tri 4928 20957 4934 20963 nw
rect 8044 20935 8224 20963
rect 8044 20901 8050 20935
rect 8084 20925 8224 20935
rect 8084 20901 8184 20925
rect 8044 20891 8184 20901
rect 8218 20891 8224 20925
rect 8044 20863 8224 20891
rect 8044 20829 8050 20863
rect 8084 20853 8224 20863
rect 8084 20829 8184 20853
rect 8044 20819 8184 20829
rect 8218 20819 8224 20853
rect 8044 20791 8224 20819
rect 8044 20757 8050 20791
rect 8084 20781 8224 20791
rect 8084 20757 8184 20781
rect 8044 20747 8184 20757
rect 8218 20747 8224 20781
rect 5040 20720 5158 20726
rect 5092 20668 5106 20720
rect 5040 20651 5158 20668
rect 5092 20599 5106 20651
rect 5040 20582 5158 20599
rect 5092 20530 5106 20582
rect 5040 20513 5158 20530
rect 5092 20461 5106 20513
rect 5040 20444 5158 20461
rect 5092 20422 5106 20444
rect 5040 20375 5046 20392
rect 5152 20375 5158 20392
rect 5040 20306 5046 20323
rect 5152 20306 5158 20323
rect 5040 20236 5046 20254
rect 5152 20236 5158 20254
rect 5040 20166 5046 20184
rect 5152 20166 5158 20184
rect 5040 19380 5046 20114
rect 5152 19380 5158 20114
rect 5040 19368 5158 19380
rect 5317 20714 5435 20726
rect 5317 20680 5323 20714
rect 5357 20680 5395 20714
rect 5429 20680 5435 20714
rect 5317 20641 5435 20680
rect 5317 20607 5323 20641
rect 5357 20607 5395 20641
rect 5429 20607 5435 20641
rect 5317 20568 5435 20607
rect 5317 20534 5323 20568
rect 5357 20534 5395 20568
rect 5429 20534 5435 20568
rect 5317 20495 5435 20534
rect 5317 20461 5323 20495
rect 5357 20461 5395 20495
rect 5429 20461 5435 20495
rect 5317 20422 5435 20461
rect 5317 19982 5323 20422
rect 5429 19982 5435 20422
rect 5317 19913 5323 19930
rect 5429 19913 5435 19930
rect 5317 19844 5323 19861
rect 5429 19844 5435 19861
rect 5317 19775 5323 19792
rect 5429 19775 5435 19792
rect 5317 19706 5323 19723
rect 5429 19706 5435 19723
rect 5317 19636 5323 19654
rect 5429 19636 5435 19654
rect 5317 19566 5323 19584
rect 5429 19566 5435 19584
rect 5317 19496 5323 19514
rect 5429 19496 5435 19514
rect 5317 19426 5323 19444
rect 5429 19426 5435 19444
rect 5369 19374 5383 19380
rect 5317 19368 5435 19374
rect 5594 20720 5712 20726
rect 5646 20668 5660 20720
rect 5594 20651 5712 20668
rect 5646 20599 5660 20651
rect 5594 20582 5712 20599
rect 5646 20530 5660 20582
rect 5594 20513 5712 20530
rect 5646 20461 5660 20513
rect 5594 20444 5712 20461
rect 5646 20422 5660 20444
rect 5594 20375 5600 20392
rect 5706 20375 5712 20392
rect 5594 20306 5600 20323
rect 5706 20306 5712 20323
rect 5594 20236 5600 20254
rect 5706 20236 5712 20254
rect 5594 20166 5600 20184
rect 5706 20166 5712 20184
rect 5594 19380 5600 20114
rect 5706 19380 5712 20114
rect 5594 19368 5712 19380
rect 5871 20714 5989 20726
rect 5871 20680 5877 20714
rect 5911 20680 5949 20714
rect 5983 20680 5989 20714
rect 5871 20641 5989 20680
rect 5871 20607 5877 20641
rect 5911 20607 5949 20641
rect 5983 20607 5989 20641
rect 5871 20568 5989 20607
rect 5871 20534 5877 20568
rect 5911 20534 5949 20568
rect 5983 20534 5989 20568
rect 5871 20495 5989 20534
rect 5871 20461 5877 20495
rect 5911 20461 5949 20495
rect 5983 20461 5989 20495
rect 5871 20422 5989 20461
rect 5871 19982 5877 20422
rect 5983 19982 5989 20422
rect 5871 19913 5877 19930
rect 5983 19913 5989 19930
rect 5871 19844 5877 19861
rect 5983 19844 5989 19861
rect 5871 19775 5877 19792
rect 5983 19775 5989 19792
rect 5871 19706 5877 19723
rect 5983 19706 5989 19723
rect 5871 19636 5877 19654
rect 5983 19636 5989 19654
rect 5871 19566 5877 19584
rect 5983 19566 5989 19584
rect 5871 19496 5877 19514
rect 5983 19496 5989 19514
rect 5871 19426 5877 19444
rect 5983 19426 5989 19444
rect 5923 19374 5937 19380
rect 5871 19368 5989 19374
rect 6148 20720 6266 20726
rect 6200 20668 6214 20720
rect 6148 20651 6266 20668
rect 6200 20599 6214 20651
rect 6148 20582 6266 20599
rect 6200 20530 6214 20582
rect 6148 20513 6266 20530
rect 6200 20461 6214 20513
rect 6148 20444 6266 20461
rect 6200 20422 6214 20444
rect 6148 20375 6154 20392
rect 6260 20375 6266 20392
rect 6148 20306 6154 20323
rect 6260 20306 6266 20323
rect 6148 20236 6154 20254
rect 6260 20236 6266 20254
rect 6148 20166 6154 20184
rect 6260 20166 6266 20184
rect 6148 19380 6154 20114
rect 6260 19380 6266 20114
rect 6148 19368 6266 19380
rect 6425 20714 6543 20726
rect 6425 20680 6431 20714
rect 6465 20680 6503 20714
rect 6537 20680 6543 20714
rect 6425 20641 6543 20680
rect 6425 20607 6431 20641
rect 6465 20607 6503 20641
rect 6537 20607 6543 20641
rect 6425 20568 6543 20607
rect 6425 20534 6431 20568
rect 6465 20534 6503 20568
rect 6537 20534 6543 20568
rect 6425 20495 6543 20534
rect 6425 20461 6431 20495
rect 6465 20461 6503 20495
rect 6537 20461 6543 20495
rect 6425 20422 6543 20461
rect 6425 19982 6431 20422
rect 6537 19982 6543 20422
rect 6425 19913 6431 19930
rect 6537 19913 6543 19930
rect 6425 19844 6431 19861
rect 6537 19844 6543 19861
rect 6425 19775 6431 19792
rect 6537 19775 6543 19792
rect 6425 19706 6431 19723
rect 6537 19706 6543 19723
rect 6425 19636 6431 19654
rect 6537 19636 6543 19654
rect 6425 19566 6431 19584
rect 6537 19566 6543 19584
rect 6425 19496 6431 19514
rect 6537 19496 6543 19514
rect 6425 19426 6431 19444
rect 6537 19426 6543 19444
rect 6477 19374 6491 19380
rect 6425 19368 6543 19374
rect 6702 20720 6820 20726
rect 6754 20668 6768 20720
rect 6702 20651 6820 20668
rect 6754 20599 6768 20651
rect 6702 20582 6820 20599
rect 6754 20530 6768 20582
rect 6702 20513 6820 20530
rect 6754 20461 6768 20513
rect 6702 20444 6820 20461
rect 6754 20422 6768 20444
rect 6702 20375 6708 20392
rect 6814 20375 6820 20392
rect 6702 20306 6708 20323
rect 6814 20306 6820 20323
rect 6702 20236 6708 20254
rect 6814 20236 6820 20254
rect 6702 20166 6708 20184
rect 6814 20166 6820 20184
rect 6702 19380 6708 20114
rect 6814 19380 6820 20114
rect 6702 19368 6820 19380
rect 6979 20714 7097 20726
rect 6979 20680 6985 20714
rect 7019 20680 7057 20714
rect 7091 20680 7097 20714
rect 6979 20641 7097 20680
rect 6979 20607 6985 20641
rect 7019 20607 7057 20641
rect 7091 20607 7097 20641
rect 6979 20568 7097 20607
rect 6979 20534 6985 20568
rect 7019 20534 7057 20568
rect 7091 20534 7097 20568
rect 6979 20495 7097 20534
rect 6979 20461 6985 20495
rect 7019 20461 7057 20495
rect 7091 20461 7097 20495
rect 6979 20422 7097 20461
rect 6979 19982 6985 20422
rect 7091 19982 7097 20422
rect 6979 19913 6985 19930
rect 7091 19913 7097 19930
rect 6979 19844 6985 19861
rect 7091 19844 7097 19861
rect 6979 19775 6985 19792
rect 7091 19775 7097 19792
rect 6979 19706 6985 19723
rect 7091 19706 7097 19723
rect 6979 19636 6985 19654
rect 7091 19636 7097 19654
rect 6979 19566 6985 19584
rect 7091 19566 7097 19584
rect 6979 19496 6985 19514
rect 7091 19496 7097 19514
rect 6979 19426 6985 19444
rect 7091 19426 7097 19444
rect 7031 19374 7045 19380
rect 6979 19368 7097 19374
rect 7256 20720 7374 20726
rect 7308 20668 7322 20720
rect 7256 20651 7374 20668
rect 7308 20599 7322 20651
rect 7256 20582 7374 20599
rect 7308 20530 7322 20582
rect 7256 20513 7374 20530
rect 7308 20461 7322 20513
rect 7256 20444 7374 20461
rect 7308 20422 7322 20444
rect 7256 20375 7262 20392
rect 7368 20375 7374 20392
rect 7256 20306 7262 20323
rect 7368 20306 7374 20323
rect 7256 20236 7262 20254
rect 7368 20236 7374 20254
rect 7256 20166 7262 20184
rect 7368 20166 7374 20184
rect 7256 19380 7262 20114
rect 7368 19380 7374 20114
rect 7256 19368 7374 19380
rect 7533 20714 7651 20726
rect 7533 20680 7539 20714
rect 7573 20680 7611 20714
rect 7645 20680 7651 20714
rect 7533 20641 7651 20680
rect 7533 20607 7539 20641
rect 7573 20607 7611 20641
rect 7645 20607 7651 20641
rect 7533 20568 7651 20607
rect 7533 20534 7539 20568
rect 7573 20534 7611 20568
rect 7645 20534 7651 20568
rect 7533 20495 7651 20534
rect 7533 20461 7539 20495
rect 7573 20461 7611 20495
rect 7645 20461 7651 20495
rect 7533 20422 7651 20461
rect 7533 19982 7539 20422
rect 7645 19982 7651 20422
rect 7533 19913 7539 19930
rect 7645 19913 7651 19930
rect 7533 19844 7539 19861
rect 7645 19844 7651 19861
rect 7533 19775 7539 19792
rect 7645 19775 7651 19792
rect 7533 19706 7539 19723
rect 7645 19706 7651 19723
rect 7533 19636 7539 19654
rect 7645 19636 7651 19654
rect 7533 19566 7539 19584
rect 7645 19566 7651 19584
rect 7533 19496 7539 19514
rect 7645 19496 7651 19514
rect 7533 19426 7539 19444
rect 7645 19426 7651 19444
rect 7585 19374 7599 19380
rect 7533 19368 7651 19374
rect 7810 20720 7928 20726
rect 7862 20668 7876 20720
rect 7810 20651 7928 20668
rect 7862 20599 7876 20651
rect 7810 20582 7928 20599
rect 7862 20530 7876 20582
rect 7810 20513 7928 20530
rect 7862 20461 7876 20513
rect 7810 20444 7928 20461
rect 7862 20422 7876 20444
rect 7810 20375 7816 20392
rect 7922 20375 7928 20392
rect 7810 20306 7816 20323
rect 7922 20306 7928 20323
rect 7810 20236 7816 20254
rect 7922 20236 7928 20254
rect 7810 20166 7816 20184
rect 7922 20166 7928 20184
rect 7810 19380 7816 20114
rect 7922 19380 7928 20114
rect 7810 19368 7928 19380
rect 8044 20724 8224 20747
rect 8044 20672 8047 20724
rect 8099 20672 8169 20724
rect 8221 20672 8224 20724
rect 8044 20655 8224 20672
rect 8044 20603 8047 20655
rect 8099 20603 8169 20655
rect 8221 20603 8224 20655
rect 8044 20586 8224 20603
rect 8044 20534 8047 20586
rect 8099 20534 8169 20586
rect 8221 20534 8224 20586
rect 8044 20531 8184 20534
rect 8218 20531 8224 20534
rect 8044 20517 8224 20531
rect 8044 20465 8047 20517
rect 8099 20465 8169 20517
rect 8221 20465 8224 20517
rect 8044 20459 8184 20465
rect 8218 20459 8224 20465
rect 8044 20448 8224 20459
rect 8044 20396 8047 20448
rect 8099 20396 8169 20448
rect 8221 20396 8224 20448
rect 8044 20387 8184 20396
rect 8218 20387 8224 20396
rect 8044 20378 8224 20387
rect 8044 20326 8047 20378
rect 8099 20326 8169 20378
rect 8221 20326 8224 20378
rect 8044 20325 8050 20326
rect 8084 20325 8184 20326
rect 8044 20315 8184 20325
rect 8218 20315 8224 20326
rect 8044 20308 8224 20315
rect 8044 20256 8047 20308
rect 8099 20256 8169 20308
rect 8221 20256 8224 20308
rect 8044 20253 8050 20256
rect 8084 20253 8184 20256
rect 8044 20243 8184 20253
rect 8218 20243 8224 20256
rect 8044 20238 8224 20243
rect 8044 20186 8047 20238
rect 8099 20186 8169 20238
rect 8221 20186 8224 20238
rect 8044 20181 8050 20186
rect 8084 20181 8184 20186
rect 8044 20171 8184 20181
rect 8218 20171 8224 20186
rect 8044 20168 8224 20171
rect 8044 20116 8047 20168
rect 8099 20116 8169 20168
rect 8221 20116 8224 20168
rect 8044 20109 8050 20116
rect 8084 20109 8184 20116
rect 8044 20099 8184 20109
rect 8218 20099 8224 20116
rect 8044 20071 8224 20099
rect 8044 20037 8050 20071
rect 8084 20061 8224 20071
rect 8084 20037 8184 20061
rect 8044 20027 8184 20037
rect 8218 20027 8224 20061
rect 8044 19999 8224 20027
rect 8044 19965 8050 19999
rect 8084 19989 8224 19999
rect 8084 19965 8184 19989
rect 8044 19955 8184 19965
rect 8218 19955 8224 19989
rect 8044 19927 8224 19955
rect 8044 19893 8050 19927
rect 8084 19917 8224 19927
rect 8084 19893 8184 19917
rect 8044 19883 8184 19893
rect 8218 19883 8224 19917
rect 8044 19855 8224 19883
rect 8044 19821 8050 19855
rect 8084 19845 8224 19855
rect 8084 19821 8184 19845
rect 8044 19811 8184 19821
rect 8218 19811 8224 19845
rect 8044 19783 8224 19811
rect 8044 19749 8050 19783
rect 8084 19773 8224 19783
rect 8084 19749 8184 19773
rect 8044 19739 8184 19749
rect 8218 19739 8224 19773
rect 8044 19711 8224 19739
rect 8044 19677 8050 19711
rect 8084 19701 8224 19711
rect 8084 19677 8184 19701
rect 8044 19667 8184 19677
rect 8218 19667 8224 19701
rect 8044 19639 8224 19667
rect 8044 19605 8050 19639
rect 8084 19629 8224 19639
rect 8084 19605 8184 19629
rect 8044 19595 8184 19605
rect 8218 19595 8224 19629
rect 8044 19567 8224 19595
rect 8044 19533 8050 19567
rect 8084 19557 8224 19567
rect 8084 19533 8184 19557
rect 8044 19523 8184 19533
rect 8218 19523 8224 19557
rect 8044 19495 8224 19523
rect 8044 19461 8050 19495
rect 8084 19485 8224 19495
rect 8084 19461 8184 19485
rect 8044 19451 8184 19461
rect 8218 19451 8224 19485
rect 8044 19423 8224 19451
rect 8044 19389 8050 19423
rect 8084 19413 8224 19423
rect 8084 19389 8184 19413
rect 8044 19379 8184 19389
rect 8218 19379 8224 19413
rect 8044 19351 8224 19379
rect 8044 19317 8050 19351
rect 8084 19341 8224 19351
rect 8084 19317 8184 19341
rect 8044 19307 8184 19317
rect 8218 19307 8224 19341
rect 8044 19279 8224 19307
rect 8044 19245 8050 19279
rect 8084 19269 8224 19279
rect 8084 19245 8184 19269
rect 8044 19235 8184 19245
rect 8218 19235 8224 19269
rect 8044 19207 8224 19235
tri 4928 19173 4954 19199 sw
rect 8044 19173 8050 19207
rect 8084 19197 8224 19207
rect 8084 19173 8184 19197
rect 4773 19167 4954 19173
tri 4954 19167 4960 19173 sw
rect 4773 19119 7729 19167
rect 4773 19085 5251 19119
rect 5285 19085 5325 19119
rect 5359 19085 5399 19119
rect 5433 19085 5473 19119
rect 5507 19085 5547 19119
rect 5581 19085 5621 19119
rect 5655 19085 5695 19119
rect 5729 19085 5769 19119
rect 5803 19085 5843 19119
rect 5877 19085 5917 19119
rect 5951 19085 5991 19119
rect 6025 19085 6065 19119
rect 6099 19085 6139 19119
rect 6173 19085 6213 19119
rect 6247 19085 6287 19119
rect 6321 19085 6361 19119
rect 6395 19085 6435 19119
rect 6469 19085 6509 19119
rect 6543 19085 6583 19119
rect 6617 19085 6657 19119
rect 6691 19085 6731 19119
rect 6765 19085 6805 19119
rect 6839 19085 6879 19119
rect 6913 19085 6953 19119
rect 6987 19085 7026 19119
rect 7060 19085 7099 19119
rect 7133 19085 7172 19119
rect 7206 19085 7245 19119
rect 7279 19085 7318 19119
rect 7352 19085 7391 19119
rect 7425 19085 7464 19119
rect 7498 19085 7537 19119
rect 7571 19085 7610 19119
rect 7644 19085 7683 19119
rect 7717 19085 7729 19119
rect 4773 19047 7729 19085
rect 8044 19163 8184 19173
rect 8218 19163 8224 19197
rect 8044 19135 8224 19163
rect 8044 19101 8050 19135
rect 8084 19125 8224 19135
rect 8084 19101 8184 19125
rect 8044 19091 8184 19101
rect 8218 19091 8224 19125
rect 8044 19063 8224 19091
rect 4773 19029 4974 19047
tri 4974 19029 4992 19047 nw
rect 8044 19029 8050 19063
rect 8084 19053 8224 19063
rect 8084 19029 8184 19053
rect 4773 19019 4964 19029
tri 4964 19019 4974 19029 nw
rect 8044 19019 8184 19029
rect 8218 19019 8224 19053
rect 4773 18991 4936 19019
tri 4936 18991 4964 19019 nw
rect 8044 18991 8224 19019
rect 4773 17291 4928 18991
tri 4928 18983 4936 18991 nw
rect 8044 18957 8050 18991
rect 8084 18981 8224 18991
rect 8084 18957 8184 18981
rect 8044 18947 8184 18957
rect 8218 18947 8224 18981
rect 8044 18919 8224 18947
rect 8044 18885 8050 18919
rect 8084 18909 8224 18919
rect 8084 18885 8184 18909
rect 8044 18875 8184 18885
rect 8218 18875 8224 18909
rect 8044 18847 8224 18875
rect 8044 18813 8050 18847
rect 8084 18837 8224 18847
rect 8084 18813 8184 18837
rect 8044 18803 8184 18813
rect 8218 18803 8224 18837
rect 8044 18775 8224 18803
rect 8044 18741 8050 18775
rect 8084 18765 8224 18775
rect 8084 18741 8184 18765
rect 8044 18731 8184 18741
rect 8218 18731 8224 18765
rect 5040 18720 5158 18726
rect 5092 18668 5106 18720
rect 5040 18651 5158 18668
rect 5092 18599 5106 18651
rect 5040 18582 5158 18599
rect 5092 18530 5106 18582
rect 5040 18513 5158 18530
rect 5092 18461 5106 18513
rect 5040 18444 5158 18461
rect 5092 18422 5106 18444
rect 5040 18375 5046 18392
rect 5152 18375 5158 18392
rect 5040 18306 5046 18323
rect 5152 18306 5158 18323
rect 5040 18236 5046 18254
rect 5152 18236 5158 18254
rect 5040 18166 5046 18184
rect 5152 18166 5158 18184
rect 5040 17380 5046 18114
rect 5152 17380 5158 18114
rect 5040 17368 5158 17380
rect 5317 18714 5435 18726
rect 5317 18680 5323 18714
rect 5357 18680 5395 18714
rect 5429 18680 5435 18714
rect 5317 18641 5435 18680
rect 5317 18607 5323 18641
rect 5357 18607 5395 18641
rect 5429 18607 5435 18641
rect 5317 18568 5435 18607
rect 5317 18534 5323 18568
rect 5357 18534 5395 18568
rect 5429 18534 5435 18568
rect 5317 18495 5435 18534
rect 5317 18461 5323 18495
rect 5357 18461 5395 18495
rect 5429 18461 5435 18495
rect 5317 18422 5435 18461
rect 5317 17982 5323 18422
rect 5429 17982 5435 18422
rect 5317 17913 5323 17930
rect 5429 17913 5435 17930
rect 5317 17844 5323 17861
rect 5429 17844 5435 17861
rect 5317 17775 5323 17792
rect 5429 17775 5435 17792
rect 5317 17706 5323 17723
rect 5429 17706 5435 17723
rect 5317 17636 5323 17654
rect 5429 17636 5435 17654
rect 5317 17566 5323 17584
rect 5429 17566 5435 17584
rect 5317 17496 5323 17514
rect 5429 17496 5435 17514
rect 5317 17426 5323 17444
rect 5429 17426 5435 17444
rect 5369 17374 5383 17380
rect 5317 17368 5435 17374
rect 5594 18720 5712 18726
rect 5646 18668 5660 18720
rect 5594 18651 5712 18668
rect 5646 18599 5660 18651
rect 5594 18582 5712 18599
rect 5646 18530 5660 18582
rect 5594 18513 5712 18530
rect 5646 18461 5660 18513
rect 5594 18444 5712 18461
rect 5646 18422 5660 18444
rect 5594 18375 5600 18392
rect 5706 18375 5712 18392
rect 5594 18306 5600 18323
rect 5706 18306 5712 18323
rect 5594 18236 5600 18254
rect 5706 18236 5712 18254
rect 5594 18166 5600 18184
rect 5706 18166 5712 18184
rect 5594 17380 5600 18114
rect 5706 17380 5712 18114
rect 5594 17368 5712 17380
rect 5871 18714 5989 18726
rect 5871 18680 5877 18714
rect 5911 18680 5949 18714
rect 5983 18680 5989 18714
rect 5871 18641 5989 18680
rect 5871 18607 5877 18641
rect 5911 18607 5949 18641
rect 5983 18607 5989 18641
rect 5871 18568 5989 18607
rect 5871 18534 5877 18568
rect 5911 18534 5949 18568
rect 5983 18534 5989 18568
rect 5871 18495 5989 18534
rect 5871 18461 5877 18495
rect 5911 18461 5949 18495
rect 5983 18461 5989 18495
rect 5871 18422 5989 18461
rect 5871 17982 5877 18422
rect 5983 17982 5989 18422
rect 5871 17913 5877 17930
rect 5983 17913 5989 17930
rect 5871 17844 5877 17861
rect 5983 17844 5989 17861
rect 5871 17775 5877 17792
rect 5983 17775 5989 17792
rect 5871 17706 5877 17723
rect 5983 17706 5989 17723
rect 5871 17636 5877 17654
rect 5983 17636 5989 17654
rect 5871 17566 5877 17584
rect 5983 17566 5989 17584
rect 5871 17496 5877 17514
rect 5983 17496 5989 17514
rect 5871 17426 5877 17444
rect 5983 17426 5989 17444
rect 5923 17374 5937 17380
rect 5871 17368 5989 17374
rect 6148 18720 6266 18726
rect 6200 18668 6214 18720
rect 6148 18651 6266 18668
rect 6200 18599 6214 18651
rect 6148 18582 6266 18599
rect 6200 18530 6214 18582
rect 6148 18513 6266 18530
rect 6200 18461 6214 18513
rect 6148 18444 6266 18461
rect 6200 18422 6214 18444
rect 6148 18375 6154 18392
rect 6260 18375 6266 18392
rect 6148 18306 6154 18323
rect 6260 18306 6266 18323
rect 6148 18236 6154 18254
rect 6260 18236 6266 18254
rect 6148 18166 6154 18184
rect 6260 18166 6266 18184
rect 6148 17380 6154 18114
rect 6260 17380 6266 18114
rect 6148 17368 6266 17380
rect 6425 18714 6543 18726
rect 6425 18680 6431 18714
rect 6465 18680 6503 18714
rect 6537 18680 6543 18714
rect 6425 18641 6543 18680
rect 6425 18607 6431 18641
rect 6465 18607 6503 18641
rect 6537 18607 6543 18641
rect 6425 18568 6543 18607
rect 6425 18534 6431 18568
rect 6465 18534 6503 18568
rect 6537 18534 6543 18568
rect 6425 18495 6543 18534
rect 6425 18461 6431 18495
rect 6465 18461 6503 18495
rect 6537 18461 6543 18495
rect 6425 18422 6543 18461
rect 6425 17982 6431 18422
rect 6537 17982 6543 18422
rect 6425 17913 6431 17930
rect 6537 17913 6543 17930
rect 6425 17844 6431 17861
rect 6537 17844 6543 17861
rect 6425 17775 6431 17792
rect 6537 17775 6543 17792
rect 6425 17706 6431 17723
rect 6537 17706 6543 17723
rect 6425 17636 6431 17654
rect 6537 17636 6543 17654
rect 6425 17566 6431 17584
rect 6537 17566 6543 17584
rect 6425 17496 6431 17514
rect 6537 17496 6543 17514
rect 6425 17426 6431 17444
rect 6537 17426 6543 17444
rect 6477 17374 6491 17380
rect 6425 17368 6543 17374
rect 6702 18720 6820 18726
rect 6754 18668 6768 18720
rect 6702 18651 6820 18668
rect 6754 18599 6768 18651
rect 6702 18582 6820 18599
rect 6754 18530 6768 18582
rect 6702 18513 6820 18530
rect 6754 18461 6768 18513
rect 6702 18444 6820 18461
rect 6754 18422 6768 18444
rect 6702 18375 6708 18392
rect 6814 18375 6820 18392
rect 6702 18306 6708 18323
rect 6814 18306 6820 18323
rect 6702 18236 6708 18254
rect 6814 18236 6820 18254
rect 6702 18166 6708 18184
rect 6814 18166 6820 18184
rect 6702 17380 6708 18114
rect 6814 17380 6820 18114
rect 6702 17368 6820 17380
rect 6979 18714 7097 18726
rect 6979 18680 6985 18714
rect 7019 18680 7057 18714
rect 7091 18680 7097 18714
rect 6979 18641 7097 18680
rect 6979 18607 6985 18641
rect 7019 18607 7057 18641
rect 7091 18607 7097 18641
rect 6979 18568 7097 18607
rect 6979 18534 6985 18568
rect 7019 18534 7057 18568
rect 7091 18534 7097 18568
rect 6979 18495 7097 18534
rect 6979 18461 6985 18495
rect 7019 18461 7057 18495
rect 7091 18461 7097 18495
rect 6979 18422 7097 18461
rect 6979 17982 6985 18422
rect 7091 17982 7097 18422
rect 6979 17913 6985 17930
rect 7091 17913 7097 17930
rect 6979 17844 6985 17861
rect 7091 17844 7097 17861
rect 6979 17775 6985 17792
rect 7091 17775 7097 17792
rect 6979 17706 6985 17723
rect 7091 17706 7097 17723
rect 6979 17636 6985 17654
rect 7091 17636 7097 17654
rect 6979 17566 6985 17584
rect 7091 17566 7097 17584
rect 6979 17496 6985 17514
rect 7091 17496 7097 17514
rect 6979 17426 6985 17444
rect 7091 17426 7097 17444
rect 7031 17374 7045 17380
rect 6979 17368 7097 17374
rect 7256 18720 7374 18726
rect 7308 18668 7322 18720
rect 7256 18651 7374 18668
rect 7308 18599 7322 18651
rect 7256 18582 7374 18599
rect 7308 18530 7322 18582
rect 7256 18513 7374 18530
rect 7308 18461 7322 18513
rect 7256 18444 7374 18461
rect 7308 18422 7322 18444
rect 7256 18375 7262 18392
rect 7368 18375 7374 18392
rect 7256 18306 7262 18323
rect 7368 18306 7374 18323
rect 7256 18236 7262 18254
rect 7368 18236 7374 18254
rect 7256 18166 7262 18184
rect 7368 18166 7374 18184
rect 7256 17380 7262 18114
rect 7368 17380 7374 18114
rect 7256 17368 7374 17380
rect 7533 18714 7651 18726
rect 7533 18680 7539 18714
rect 7573 18680 7611 18714
rect 7645 18680 7651 18714
rect 7533 18641 7651 18680
rect 7533 18607 7539 18641
rect 7573 18607 7611 18641
rect 7645 18607 7651 18641
rect 7533 18568 7651 18607
rect 7533 18534 7539 18568
rect 7573 18534 7611 18568
rect 7645 18534 7651 18568
rect 7533 18495 7651 18534
rect 7533 18461 7539 18495
rect 7573 18461 7611 18495
rect 7645 18461 7651 18495
rect 7533 18422 7651 18461
rect 7533 17982 7539 18422
rect 7645 17982 7651 18422
rect 7533 17913 7539 17930
rect 7645 17913 7651 17930
rect 7533 17844 7539 17861
rect 7645 17844 7651 17861
rect 7533 17775 7539 17792
rect 7645 17775 7651 17792
rect 7533 17706 7539 17723
rect 7645 17706 7651 17723
rect 7533 17636 7539 17654
rect 7645 17636 7651 17654
rect 7533 17566 7539 17584
rect 7645 17566 7651 17584
rect 7533 17496 7539 17514
rect 7645 17496 7651 17514
rect 7533 17426 7539 17444
rect 7645 17426 7651 17444
rect 7585 17374 7599 17380
rect 7533 17368 7651 17374
rect 7810 18720 7928 18726
rect 7862 18668 7876 18720
rect 7810 18651 7928 18668
rect 7862 18599 7876 18651
rect 7810 18582 7928 18599
rect 7862 18530 7876 18582
rect 7810 18513 7928 18530
rect 7862 18461 7876 18513
rect 7810 18444 7928 18461
rect 7862 18422 7876 18444
rect 7810 18375 7816 18392
rect 7922 18375 7928 18392
rect 7810 18306 7816 18323
rect 7922 18306 7928 18323
rect 7810 18236 7816 18254
rect 7922 18236 7928 18254
rect 7810 18166 7816 18184
rect 7922 18166 7928 18184
rect 7810 17380 7816 18114
rect 7922 17380 7928 18114
rect 7810 17368 7928 17380
rect 8044 18724 8224 18731
rect 8044 18672 8047 18724
rect 8099 18672 8169 18724
rect 8221 18672 8224 18724
rect 8044 18669 8050 18672
rect 8084 18669 8184 18672
rect 8044 18659 8184 18669
rect 8218 18659 8224 18672
rect 8044 18655 8224 18659
rect 8044 18603 8047 18655
rect 8099 18603 8169 18655
rect 8221 18603 8224 18655
rect 8044 18597 8050 18603
rect 8084 18597 8184 18603
rect 8044 18587 8184 18597
rect 8218 18587 8224 18603
rect 8044 18586 8224 18587
rect 8044 18534 8047 18586
rect 8099 18534 8169 18586
rect 8221 18534 8224 18586
rect 8044 18525 8050 18534
rect 8084 18525 8184 18534
rect 8044 18517 8184 18525
rect 8218 18517 8224 18534
rect 8044 18465 8047 18517
rect 8099 18465 8169 18517
rect 8221 18465 8224 18517
rect 8044 18453 8050 18465
rect 8084 18453 8184 18465
rect 8044 18448 8184 18453
rect 8218 18448 8224 18465
rect 8044 18396 8047 18448
rect 8099 18396 8169 18448
rect 8221 18396 8224 18448
rect 8044 18381 8050 18396
rect 8084 18381 8184 18396
rect 8044 18378 8184 18381
rect 8218 18378 8224 18396
rect 8044 18326 8047 18378
rect 8099 18326 8169 18378
rect 8221 18326 8224 18378
rect 8044 18309 8050 18326
rect 8084 18309 8184 18326
rect 8044 18308 8184 18309
rect 8218 18308 8224 18326
rect 8044 18256 8047 18308
rect 8099 18256 8169 18308
rect 8221 18256 8224 18308
rect 8044 18238 8050 18256
rect 8084 18238 8184 18256
rect 8218 18238 8224 18256
rect 8044 18186 8047 18238
rect 8099 18186 8169 18238
rect 8221 18186 8224 18238
rect 8044 18168 8050 18186
rect 8084 18168 8184 18186
rect 8218 18168 8224 18186
rect 8044 18116 8047 18168
rect 8099 18116 8169 18168
rect 8221 18116 8224 18168
rect 8044 18093 8050 18116
rect 8084 18093 8184 18116
rect 8044 18083 8184 18093
rect 8218 18083 8224 18116
rect 8044 18055 8224 18083
rect 8044 18021 8050 18055
rect 8084 18045 8224 18055
rect 8084 18021 8184 18045
rect 8044 18011 8184 18021
rect 8218 18011 8224 18045
rect 8044 17983 8224 18011
rect 8044 17949 8050 17983
rect 8084 17973 8224 17983
rect 8084 17949 8184 17973
rect 8044 17939 8184 17949
rect 8218 17939 8224 17973
rect 8044 17911 8224 17939
rect 8044 17877 8050 17911
rect 8084 17901 8224 17911
rect 8084 17877 8184 17901
rect 8044 17867 8184 17877
rect 8218 17867 8224 17901
rect 8044 17839 8224 17867
rect 8044 17805 8050 17839
rect 8084 17829 8224 17839
rect 8084 17805 8184 17829
rect 8044 17795 8184 17805
rect 8218 17795 8224 17829
rect 8044 17767 8224 17795
rect 8044 17733 8050 17767
rect 8084 17757 8224 17767
rect 8084 17733 8184 17757
rect 8044 17723 8184 17733
rect 8218 17723 8224 17757
rect 8044 17695 8224 17723
rect 8044 17661 8050 17695
rect 8084 17685 8224 17695
rect 8084 17661 8184 17685
rect 8044 17651 8184 17661
rect 8218 17651 8224 17685
rect 8044 17623 8224 17651
rect 8044 17589 8050 17623
rect 8084 17613 8224 17623
rect 8084 17589 8184 17613
rect 8044 17579 8184 17589
rect 8218 17579 8224 17613
rect 8044 17551 8224 17579
rect 8044 17517 8050 17551
rect 8084 17541 8224 17551
rect 8084 17517 8184 17541
rect 8044 17507 8184 17517
rect 8218 17507 8224 17541
rect 8044 17479 8224 17507
rect 8044 17445 8050 17479
rect 8084 17469 8224 17479
rect 8084 17445 8184 17469
rect 8044 17435 8184 17445
rect 8218 17435 8224 17469
rect 8044 17407 8224 17435
rect 8044 17373 8050 17407
rect 8084 17397 8224 17407
rect 8084 17373 8184 17397
rect 8044 17363 8184 17373
rect 8218 17363 8224 17397
rect 8044 17335 8224 17363
rect 8044 17301 8050 17335
rect 8084 17325 8224 17335
rect 8084 17301 8184 17325
tri 4928 17291 4938 17301 sw
rect 8044 17291 8184 17301
rect 8218 17291 8224 17325
rect 4773 17275 4938 17291
tri 4938 17275 4954 17291 sw
rect 4773 17245 7729 17275
rect 4773 17211 5251 17245
rect 5285 17211 5325 17245
rect 5359 17211 5399 17245
rect 5433 17211 5473 17245
rect 5507 17211 5547 17245
rect 5581 17211 5621 17245
rect 5655 17211 5695 17245
rect 5729 17211 5769 17245
rect 5803 17211 5843 17245
rect 5877 17211 5917 17245
rect 5951 17211 5991 17245
rect 6025 17211 6065 17245
rect 6099 17211 6139 17245
rect 6173 17211 6213 17245
rect 6247 17211 6287 17245
rect 6321 17211 6361 17245
rect 6395 17211 6435 17245
rect 6469 17211 6509 17245
rect 6543 17211 6583 17245
rect 6617 17211 6657 17245
rect 6691 17211 6731 17245
rect 6765 17211 6805 17245
rect 6839 17211 6879 17245
rect 6913 17211 6953 17245
rect 6987 17211 7026 17245
rect 7060 17211 7099 17245
rect 7133 17211 7172 17245
rect 7206 17211 7245 17245
rect 7279 17211 7318 17245
rect 7352 17211 7391 17245
rect 7425 17211 7464 17245
rect 7498 17211 7537 17245
rect 7571 17211 7610 17245
rect 7644 17211 7683 17245
rect 7717 17211 7729 17245
rect 4773 17155 7729 17211
rect 8044 17263 8224 17291
rect 8044 17229 8050 17263
rect 8084 17253 8224 17263
rect 8084 17229 8184 17253
rect 8044 17219 8184 17229
rect 8218 17219 8224 17253
rect 8044 17191 8224 17219
rect 8044 17157 8050 17191
rect 8084 17181 8224 17191
rect 8084 17157 8184 17181
rect 4773 17147 4974 17155
tri 4974 17147 4982 17155 nw
rect 8044 17147 8184 17157
rect 8218 17147 8224 17181
rect 4773 17119 4946 17147
tri 4946 17119 4974 17147 nw
rect 8044 17119 8224 17147
rect 2270 15852 2450 15890
rect 2270 15818 2276 15852
rect 2310 15818 2410 15852
rect 2444 15818 2450 15852
rect 2270 15780 2450 15818
rect 2270 15746 2276 15780
rect 2310 15746 2410 15780
rect 2444 15746 2450 15780
rect 2270 15708 2450 15746
rect 2270 15674 2276 15708
rect 2310 15674 2410 15708
rect 2444 15674 2450 15708
tri 4757 15679 4773 15695 se
rect 4773 15679 4928 17119
tri 4928 17101 4946 17119 nw
rect 8044 17085 8050 17119
rect 8084 17109 8224 17119
rect 8084 17085 8184 17109
rect 8044 17075 8184 17085
rect 8218 17075 8224 17109
rect 8044 17047 8224 17075
rect 8044 17013 8050 17047
rect 8084 17037 8224 17047
rect 8084 17013 8184 17037
rect 5077 16989 7884 17004
rect 5077 16955 5089 16989
rect 5123 16970 5162 16989
rect 5196 16970 5235 16989
rect 5269 16970 5308 16989
rect 5342 16970 5381 16989
rect 5415 16970 5454 16989
rect 5488 16970 5527 16989
rect 5561 16970 5600 16989
rect 5634 16970 5673 16989
rect 5707 16970 5746 16989
rect 5780 16970 5819 16989
rect 5853 16970 5892 16989
rect 5926 16970 5965 16989
rect 5999 16970 6038 16989
rect 6072 16970 6110 16989
rect 6144 16970 6182 16989
rect 6216 16970 6254 16989
rect 6288 16970 6326 16989
rect 6360 16970 6398 16989
rect 6432 16970 6470 16989
rect 6504 16970 6542 16989
rect 6576 16970 6614 16989
rect 6648 16970 6686 16989
rect 6720 16970 6758 16989
rect 6792 16970 6830 16989
rect 6864 16970 6902 16989
rect 6936 16970 6974 16989
rect 7008 16970 7046 16989
rect 7080 16970 7118 16989
rect 7152 16970 7190 16989
rect 7224 16970 7262 16989
rect 7296 16970 7334 16989
rect 7368 16970 7406 16989
rect 7440 16970 7478 16989
rect 7512 16970 7550 16989
rect 7584 16970 7622 16989
rect 7656 16970 7694 16989
rect 7728 16970 7766 16989
rect 7800 16970 7838 16989
rect 5234 16955 5235 16970
rect 5300 16955 5308 16970
rect 5077 16918 5116 16955
rect 5168 16918 5182 16955
rect 5234 16918 5248 16955
rect 5300 16918 5314 16955
rect 5366 16918 5380 16970
rect 5432 16918 5446 16970
rect 5498 16918 5512 16970
rect 5564 16918 5578 16970
rect 5634 16955 5644 16970
rect 5707 16955 5710 16970
rect 5960 16955 5965 16970
rect 6026 16955 6038 16970
rect 5630 16918 5644 16955
rect 5696 16918 5710 16955
rect 5762 16918 5776 16955
rect 5828 16918 5842 16955
rect 5894 16918 5908 16955
rect 5960 16918 5974 16955
rect 6026 16918 6040 16955
rect 6092 16918 6106 16970
rect 6158 16918 6172 16970
rect 6224 16918 6238 16970
rect 6290 16918 6304 16970
rect 6360 16955 6370 16970
rect 6432 16955 6436 16970
rect 6683 16955 6686 16970
rect 6748 16955 6758 16970
rect 6356 16918 6370 16955
rect 6422 16918 6436 16955
rect 6488 16918 6501 16955
rect 6553 16918 6566 16955
rect 6618 16918 6631 16955
rect 6683 16918 6696 16955
rect 6748 16918 6761 16955
rect 6813 16918 6826 16970
rect 6878 16918 6891 16970
rect 6943 16918 6956 16970
rect 7008 16918 7021 16970
rect 7080 16955 7086 16970
rect 7333 16955 7334 16970
rect 7398 16955 7406 16970
rect 7073 16918 7086 16955
rect 7138 16918 7151 16955
rect 7203 16918 7216 16955
rect 7268 16918 7281 16955
rect 7333 16918 7346 16955
rect 7398 16918 7411 16955
rect 7463 16918 7476 16970
rect 7528 16918 7541 16970
rect 7593 16918 7606 16970
rect 7658 16918 7671 16970
rect 7728 16955 7736 16970
rect 7800 16955 7801 16970
rect 7872 16955 7884 16989
rect 7723 16918 7736 16955
rect 7788 16918 7801 16955
rect 7853 16918 7884 16955
rect 5077 16913 7884 16918
rect 5077 16879 5089 16913
rect 5123 16904 5162 16913
rect 5196 16904 5235 16913
rect 5269 16904 5308 16913
rect 5342 16904 5381 16913
rect 5415 16904 5454 16913
rect 5488 16904 5527 16913
rect 5561 16904 5600 16913
rect 5634 16904 5673 16913
rect 5707 16904 5746 16913
rect 5780 16904 5819 16913
rect 5853 16904 5892 16913
rect 5926 16904 5965 16913
rect 5999 16904 6038 16913
rect 6072 16904 6110 16913
rect 6144 16904 6182 16913
rect 6216 16904 6254 16913
rect 6288 16904 6326 16913
rect 6360 16904 6398 16913
rect 6432 16904 6470 16913
rect 6504 16904 6542 16913
rect 6576 16904 6614 16913
rect 6648 16904 6686 16913
rect 6720 16904 6758 16913
rect 6792 16904 6830 16913
rect 6864 16904 6902 16913
rect 6936 16904 6974 16913
rect 7008 16904 7046 16913
rect 7080 16904 7118 16913
rect 7152 16904 7190 16913
rect 7224 16904 7262 16913
rect 7296 16904 7334 16913
rect 7368 16904 7406 16913
rect 7440 16904 7478 16913
rect 7512 16904 7550 16913
rect 7584 16904 7622 16913
rect 7656 16904 7694 16913
rect 7728 16904 7766 16913
rect 7800 16904 7838 16913
rect 5234 16879 5235 16904
rect 5300 16879 5308 16904
rect 5077 16852 5116 16879
rect 5168 16852 5182 16879
rect 5234 16852 5248 16879
rect 5300 16852 5314 16879
rect 5366 16852 5380 16904
rect 5432 16852 5446 16904
rect 5498 16852 5512 16904
rect 5564 16852 5578 16904
rect 5634 16879 5644 16904
rect 5707 16879 5710 16904
rect 5960 16879 5965 16904
rect 6026 16879 6038 16904
rect 5630 16852 5644 16879
rect 5696 16852 5710 16879
rect 5762 16852 5776 16879
rect 5828 16852 5842 16879
rect 5894 16852 5908 16879
rect 5960 16852 5974 16879
rect 6026 16852 6040 16879
rect 6092 16852 6106 16904
rect 6158 16852 6172 16904
rect 6224 16852 6238 16904
rect 6290 16852 6304 16904
rect 6360 16879 6370 16904
rect 6432 16879 6436 16904
rect 6683 16879 6686 16904
rect 6748 16879 6758 16904
rect 6356 16852 6370 16879
rect 6422 16852 6436 16879
rect 6488 16852 6501 16879
rect 6553 16852 6566 16879
rect 6618 16852 6631 16879
rect 6683 16852 6696 16879
rect 6748 16852 6761 16879
rect 6813 16852 6826 16904
rect 6878 16852 6891 16904
rect 6943 16852 6956 16904
rect 7008 16852 7021 16904
rect 7080 16879 7086 16904
rect 7333 16879 7334 16904
rect 7398 16879 7406 16904
rect 7073 16852 7086 16879
rect 7138 16852 7151 16879
rect 7203 16852 7216 16879
rect 7268 16852 7281 16879
rect 7333 16852 7346 16879
rect 7398 16852 7411 16879
rect 7463 16852 7476 16904
rect 7528 16852 7541 16904
rect 7593 16852 7606 16904
rect 7658 16852 7671 16904
rect 7728 16879 7736 16904
rect 7800 16879 7801 16904
rect 7872 16879 7884 16913
rect 7723 16852 7736 16879
rect 7788 16852 7801 16879
rect 7853 16852 7884 16879
rect 5077 16838 7884 16852
rect 5077 16837 5116 16838
rect 5168 16837 5182 16838
rect 5234 16837 5248 16838
rect 5300 16837 5314 16838
rect 5077 16803 5089 16837
rect 5234 16803 5235 16837
rect 5300 16803 5308 16837
rect 5077 16786 5116 16803
rect 5168 16786 5182 16803
rect 5234 16786 5248 16803
rect 5300 16786 5314 16803
rect 5366 16786 5380 16838
rect 5432 16786 5446 16838
rect 5498 16786 5512 16838
rect 5564 16786 5578 16838
rect 5630 16837 5644 16838
rect 5696 16837 5710 16838
rect 5762 16837 5776 16838
rect 5828 16837 5842 16838
rect 5894 16837 5908 16838
rect 5960 16837 5974 16838
rect 6026 16837 6040 16838
rect 5634 16803 5644 16837
rect 5707 16803 5710 16837
rect 5960 16803 5965 16837
rect 6026 16803 6038 16837
rect 5630 16786 5644 16803
rect 5696 16786 5710 16803
rect 5762 16786 5776 16803
rect 5828 16786 5842 16803
rect 5894 16786 5908 16803
rect 5960 16786 5974 16803
rect 6026 16786 6040 16803
rect 6092 16786 6106 16838
rect 6158 16786 6172 16838
rect 6224 16786 6238 16838
rect 6290 16786 6304 16838
rect 6356 16837 6370 16838
rect 6422 16837 6436 16838
rect 6488 16837 6501 16838
rect 6553 16837 6566 16838
rect 6618 16837 6631 16838
rect 6683 16837 6696 16838
rect 6748 16837 6761 16838
rect 6360 16803 6370 16837
rect 6432 16803 6436 16837
rect 6683 16803 6686 16837
rect 6748 16803 6758 16837
rect 6356 16786 6370 16803
rect 6422 16786 6436 16803
rect 6488 16786 6501 16803
rect 6553 16786 6566 16803
rect 6618 16786 6631 16803
rect 6683 16786 6696 16803
rect 6748 16786 6761 16803
rect 6813 16786 6826 16838
rect 6878 16786 6891 16838
rect 6943 16786 6956 16838
rect 7008 16786 7021 16838
rect 7073 16837 7086 16838
rect 7138 16837 7151 16838
rect 7203 16837 7216 16838
rect 7268 16837 7281 16838
rect 7333 16837 7346 16838
rect 7398 16837 7411 16838
rect 7080 16803 7086 16837
rect 7333 16803 7334 16837
rect 7398 16803 7406 16837
rect 7073 16786 7086 16803
rect 7138 16786 7151 16803
rect 7203 16786 7216 16803
rect 7268 16786 7281 16803
rect 7333 16786 7346 16803
rect 7398 16786 7411 16803
rect 7463 16786 7476 16838
rect 7528 16786 7541 16838
rect 7593 16786 7606 16838
rect 7658 16786 7671 16838
rect 7723 16837 7736 16838
rect 7788 16837 7801 16838
rect 7853 16837 7884 16838
rect 7728 16803 7736 16837
rect 7800 16803 7801 16837
rect 7872 16803 7884 16837
rect 7723 16786 7736 16803
rect 7788 16786 7801 16803
rect 7853 16786 7884 16803
rect 5077 16772 7884 16786
rect 5077 16761 5116 16772
rect 5168 16761 5182 16772
rect 5234 16761 5248 16772
rect 5300 16761 5314 16772
rect 5077 16727 5089 16761
rect 5234 16727 5235 16761
rect 5300 16727 5308 16761
rect 5077 16720 5116 16727
rect 5168 16720 5182 16727
rect 5234 16720 5248 16727
rect 5300 16720 5314 16727
rect 5366 16720 5380 16772
rect 5432 16720 5446 16772
rect 5498 16720 5512 16772
rect 5564 16720 5578 16772
rect 5630 16761 5644 16772
rect 5696 16761 5710 16772
rect 5762 16761 5776 16772
rect 5828 16761 5842 16772
rect 5894 16761 5908 16772
rect 5960 16761 5974 16772
rect 6026 16761 6040 16772
rect 5634 16727 5644 16761
rect 5707 16727 5710 16761
rect 5960 16727 5965 16761
rect 6026 16727 6038 16761
rect 5630 16720 5644 16727
rect 5696 16720 5710 16727
rect 5762 16720 5776 16727
rect 5828 16720 5842 16727
rect 5894 16720 5908 16727
rect 5960 16720 5974 16727
rect 6026 16720 6040 16727
rect 6092 16720 6106 16772
rect 6158 16720 6172 16772
rect 6224 16720 6238 16772
rect 6290 16720 6304 16772
rect 6356 16761 6370 16772
rect 6422 16761 6436 16772
rect 6488 16761 6501 16772
rect 6553 16761 6566 16772
rect 6618 16761 6631 16772
rect 6683 16761 6696 16772
rect 6748 16761 6761 16772
rect 6360 16727 6370 16761
rect 6432 16727 6436 16761
rect 6683 16727 6686 16761
rect 6748 16727 6758 16761
rect 6356 16720 6370 16727
rect 6422 16720 6436 16727
rect 6488 16720 6501 16727
rect 6553 16720 6566 16727
rect 6618 16720 6631 16727
rect 6683 16720 6696 16727
rect 6748 16720 6761 16727
rect 6813 16720 6826 16772
rect 6878 16720 6891 16772
rect 6943 16720 6956 16772
rect 7008 16720 7021 16772
rect 7073 16761 7086 16772
rect 7138 16761 7151 16772
rect 7203 16761 7216 16772
rect 7268 16761 7281 16772
rect 7333 16761 7346 16772
rect 7398 16761 7411 16772
rect 7080 16727 7086 16761
rect 7333 16727 7334 16761
rect 7398 16727 7406 16761
rect 7073 16720 7086 16727
rect 7138 16720 7151 16727
rect 7203 16720 7216 16727
rect 7268 16720 7281 16727
rect 7333 16720 7346 16727
rect 7398 16720 7411 16727
rect 7463 16720 7476 16772
rect 7528 16720 7541 16772
rect 7593 16720 7606 16772
rect 7658 16720 7671 16772
rect 7723 16761 7736 16772
rect 7788 16761 7801 16772
rect 7853 16761 7884 16772
rect 7728 16727 7736 16761
rect 7800 16727 7801 16761
rect 7872 16727 7884 16761
rect 7723 16720 7736 16727
rect 7788 16720 7801 16727
rect 7853 16720 7884 16727
rect 5077 16706 7884 16720
rect 5077 16685 5116 16706
rect 5168 16685 5182 16706
rect 5234 16685 5248 16706
rect 5300 16685 5314 16706
rect 5077 16651 5089 16685
rect 5234 16654 5235 16685
rect 5300 16654 5308 16685
rect 5366 16654 5380 16706
rect 5432 16654 5446 16706
rect 5498 16654 5512 16706
rect 5564 16654 5578 16706
rect 5630 16685 5644 16706
rect 5696 16685 5710 16706
rect 5762 16685 5776 16706
rect 5828 16685 5842 16706
rect 5894 16685 5908 16706
rect 5960 16685 5974 16706
rect 6026 16685 6040 16706
rect 5634 16654 5644 16685
rect 5707 16654 5710 16685
rect 5960 16654 5965 16685
rect 6026 16654 6038 16685
rect 6092 16654 6106 16706
rect 6158 16654 6172 16706
rect 6224 16654 6238 16706
rect 6290 16654 6304 16706
rect 6356 16685 6370 16706
rect 6422 16685 6436 16706
rect 6488 16685 6501 16706
rect 6553 16685 6566 16706
rect 6618 16685 6631 16706
rect 6683 16685 6696 16706
rect 6748 16685 6761 16706
rect 6360 16654 6370 16685
rect 6432 16654 6436 16685
rect 6683 16654 6686 16685
rect 6748 16654 6758 16685
rect 6813 16654 6826 16706
rect 6878 16654 6891 16706
rect 6943 16654 6956 16706
rect 7008 16654 7021 16706
rect 7073 16685 7086 16706
rect 7138 16685 7151 16706
rect 7203 16685 7216 16706
rect 7268 16685 7281 16706
rect 7333 16685 7346 16706
rect 7398 16685 7411 16706
rect 7080 16654 7086 16685
rect 7333 16654 7334 16685
rect 7398 16654 7406 16685
rect 7463 16654 7476 16706
rect 7528 16654 7541 16706
rect 7593 16654 7606 16706
rect 7658 16654 7671 16706
rect 7723 16685 7736 16706
rect 7788 16685 7801 16706
rect 7853 16685 7884 16706
rect 7728 16654 7736 16685
rect 7800 16654 7801 16685
rect 5123 16651 5162 16654
rect 5196 16651 5235 16654
rect 5269 16651 5308 16654
rect 5342 16651 5381 16654
rect 5415 16651 5454 16654
rect 5488 16651 5527 16654
rect 5561 16651 5600 16654
rect 5634 16651 5673 16654
rect 5707 16651 5746 16654
rect 5780 16651 5819 16654
rect 5853 16651 5892 16654
rect 5926 16651 5965 16654
rect 5999 16651 6038 16654
rect 6072 16651 6110 16654
rect 6144 16651 6182 16654
rect 6216 16651 6254 16654
rect 6288 16651 6326 16654
rect 6360 16651 6398 16654
rect 6432 16651 6470 16654
rect 6504 16651 6542 16654
rect 6576 16651 6614 16654
rect 6648 16651 6686 16654
rect 6720 16651 6758 16654
rect 6792 16651 6830 16654
rect 6864 16651 6902 16654
rect 6936 16651 6974 16654
rect 7008 16651 7046 16654
rect 7080 16651 7118 16654
rect 7152 16651 7190 16654
rect 7224 16651 7262 16654
rect 7296 16651 7334 16654
rect 7368 16651 7406 16654
rect 7440 16651 7478 16654
rect 7512 16651 7550 16654
rect 7584 16651 7622 16654
rect 7656 16651 7694 16654
rect 7728 16651 7766 16654
rect 7800 16651 7838 16654
rect 7872 16651 7884 16685
rect 5077 16640 7884 16651
rect 5077 16609 5116 16640
rect 5168 16609 5182 16640
rect 5234 16609 5248 16640
rect 5300 16609 5314 16640
rect 5077 16575 5089 16609
rect 5234 16588 5235 16609
rect 5300 16588 5308 16609
rect 5366 16588 5380 16640
rect 5432 16588 5446 16640
rect 5498 16588 5512 16640
rect 5564 16588 5578 16640
rect 5630 16609 5644 16640
rect 5696 16609 5710 16640
rect 5762 16609 5776 16640
rect 5828 16609 5842 16640
rect 5894 16609 5908 16640
rect 5960 16609 5974 16640
rect 6026 16609 6040 16640
rect 5634 16588 5644 16609
rect 5707 16588 5710 16609
rect 5960 16588 5965 16609
rect 6026 16588 6038 16609
rect 6092 16588 6106 16640
rect 6158 16588 6172 16640
rect 6224 16588 6238 16640
rect 6290 16588 6304 16640
rect 6356 16609 6370 16640
rect 6422 16609 6436 16640
rect 6488 16609 6501 16640
rect 6553 16609 6566 16640
rect 6618 16609 6631 16640
rect 6683 16609 6696 16640
rect 6748 16609 6761 16640
rect 6360 16588 6370 16609
rect 6432 16588 6436 16609
rect 6683 16588 6686 16609
rect 6748 16588 6758 16609
rect 6813 16588 6826 16640
rect 6878 16588 6891 16640
rect 6943 16588 6956 16640
rect 7008 16588 7021 16640
rect 7073 16609 7086 16640
rect 7138 16609 7151 16640
rect 7203 16609 7216 16640
rect 7268 16609 7281 16640
rect 7333 16609 7346 16640
rect 7398 16609 7411 16640
rect 7080 16588 7086 16609
rect 7333 16588 7334 16609
rect 7398 16588 7406 16609
rect 7463 16588 7476 16640
rect 7528 16588 7541 16640
rect 7593 16588 7606 16640
rect 7658 16588 7671 16640
rect 7723 16609 7736 16640
rect 7788 16609 7801 16640
rect 7853 16609 7884 16640
rect 7728 16588 7736 16609
rect 7800 16588 7801 16609
rect 5123 16575 5162 16588
rect 5196 16575 5235 16588
rect 5269 16575 5308 16588
rect 5342 16575 5381 16588
rect 5415 16575 5454 16588
rect 5488 16575 5527 16588
rect 5561 16575 5600 16588
rect 5634 16575 5673 16588
rect 5707 16575 5746 16588
rect 5780 16575 5819 16588
rect 5853 16575 5892 16588
rect 5926 16575 5965 16588
rect 5999 16575 6038 16588
rect 6072 16575 6110 16588
rect 6144 16575 6182 16588
rect 6216 16575 6254 16588
rect 6288 16575 6326 16588
rect 6360 16575 6398 16588
rect 6432 16575 6470 16588
rect 6504 16575 6542 16588
rect 6576 16575 6614 16588
rect 6648 16575 6686 16588
rect 6720 16575 6758 16588
rect 6792 16575 6830 16588
rect 6864 16575 6902 16588
rect 6936 16575 6974 16588
rect 7008 16575 7046 16588
rect 7080 16575 7118 16588
rect 7152 16575 7190 16588
rect 7224 16575 7262 16588
rect 7296 16575 7334 16588
rect 7368 16575 7406 16588
rect 7440 16575 7478 16588
rect 7512 16575 7550 16588
rect 7584 16575 7622 16588
rect 7656 16575 7694 16588
rect 7728 16575 7766 16588
rect 7800 16575 7838 16588
rect 7872 16575 7884 16609
rect 5077 16574 7884 16575
rect 5077 16533 5116 16574
rect 5168 16533 5182 16574
rect 5234 16533 5248 16574
rect 5300 16533 5314 16574
rect 5077 16499 5089 16533
rect 5234 16522 5235 16533
rect 5300 16522 5308 16533
rect 5366 16522 5380 16574
rect 5432 16522 5446 16574
rect 5498 16522 5512 16574
rect 5564 16522 5578 16574
rect 5630 16533 5644 16574
rect 5696 16533 5710 16574
rect 5762 16533 5776 16574
rect 5828 16533 5842 16574
rect 5894 16533 5908 16574
rect 5960 16533 5974 16574
rect 6026 16533 6040 16574
rect 5634 16522 5644 16533
rect 5707 16522 5710 16533
rect 5960 16522 5965 16533
rect 6026 16522 6038 16533
rect 6092 16522 6106 16574
rect 6158 16522 6172 16574
rect 6224 16522 6238 16574
rect 6290 16522 6304 16574
rect 6356 16533 6370 16574
rect 6422 16533 6436 16574
rect 6488 16533 6501 16574
rect 6553 16533 6566 16574
rect 6618 16533 6631 16574
rect 6683 16533 6696 16574
rect 6748 16533 6761 16574
rect 6360 16522 6370 16533
rect 6432 16522 6436 16533
rect 6683 16522 6686 16533
rect 6748 16522 6758 16533
rect 6813 16522 6826 16574
rect 6878 16522 6891 16574
rect 6943 16522 6956 16574
rect 7008 16522 7021 16574
rect 7073 16533 7086 16574
rect 7138 16533 7151 16574
rect 7203 16533 7216 16574
rect 7268 16533 7281 16574
rect 7333 16533 7346 16574
rect 7398 16533 7411 16574
rect 7080 16522 7086 16533
rect 7333 16522 7334 16533
rect 7398 16522 7406 16533
rect 7463 16522 7476 16574
rect 7528 16522 7541 16574
rect 7593 16522 7606 16574
rect 7658 16522 7671 16574
rect 7723 16533 7736 16574
rect 7788 16533 7801 16574
rect 7853 16533 7884 16574
rect 7728 16522 7736 16533
rect 7800 16522 7801 16533
rect 5123 16508 5162 16522
rect 5196 16508 5235 16522
rect 5269 16508 5308 16522
rect 5342 16508 5381 16522
rect 5415 16508 5454 16522
rect 5488 16508 5527 16522
rect 5561 16508 5600 16522
rect 5634 16508 5673 16522
rect 5707 16508 5746 16522
rect 5780 16508 5819 16522
rect 5853 16508 5892 16522
rect 5926 16508 5965 16522
rect 5999 16508 6038 16522
rect 6072 16508 6110 16522
rect 6144 16508 6182 16522
rect 6216 16508 6254 16522
rect 6288 16508 6326 16522
rect 6360 16508 6398 16522
rect 6432 16508 6470 16522
rect 6504 16508 6542 16522
rect 6576 16508 6614 16522
rect 6648 16508 6686 16522
rect 6720 16508 6758 16522
rect 6792 16508 6830 16522
rect 6864 16508 6902 16522
rect 6936 16508 6974 16522
rect 7008 16508 7046 16522
rect 7080 16508 7118 16522
rect 7152 16508 7190 16522
rect 7224 16508 7262 16522
rect 7296 16508 7334 16522
rect 7368 16508 7406 16522
rect 7440 16508 7478 16522
rect 7512 16508 7550 16522
rect 7584 16508 7622 16522
rect 7656 16508 7694 16522
rect 7728 16508 7766 16522
rect 7800 16508 7838 16522
rect 5234 16499 5235 16508
rect 5300 16499 5308 16508
rect 5077 16457 5116 16499
rect 5168 16457 5182 16499
rect 5234 16457 5248 16499
rect 5300 16457 5314 16499
rect 5077 16423 5089 16457
rect 5234 16456 5235 16457
rect 5300 16456 5308 16457
rect 5366 16456 5380 16508
rect 5432 16456 5446 16508
rect 5498 16456 5512 16508
rect 5564 16456 5578 16508
rect 5634 16499 5644 16508
rect 5707 16499 5710 16508
rect 5960 16499 5965 16508
rect 6026 16499 6038 16508
rect 5630 16457 5644 16499
rect 5696 16457 5710 16499
rect 5762 16457 5776 16499
rect 5828 16457 5842 16499
rect 5894 16457 5908 16499
rect 5960 16457 5974 16499
rect 6026 16457 6040 16499
rect 5634 16456 5644 16457
rect 5707 16456 5710 16457
rect 5960 16456 5965 16457
rect 6026 16456 6038 16457
rect 6092 16456 6106 16508
rect 6158 16456 6172 16508
rect 6224 16456 6238 16508
rect 6290 16456 6304 16508
rect 6360 16499 6370 16508
rect 6432 16499 6436 16508
rect 6683 16499 6686 16508
rect 6748 16499 6758 16508
rect 6356 16457 6370 16499
rect 6422 16457 6436 16499
rect 6488 16457 6501 16499
rect 6553 16457 6566 16499
rect 6618 16457 6631 16499
rect 6683 16457 6696 16499
rect 6748 16457 6761 16499
rect 6360 16456 6370 16457
rect 6432 16456 6436 16457
rect 6683 16456 6686 16457
rect 6748 16456 6758 16457
rect 6813 16456 6826 16508
rect 6878 16456 6891 16508
rect 6943 16456 6956 16508
rect 7008 16456 7021 16508
rect 7080 16499 7086 16508
rect 7333 16499 7334 16508
rect 7398 16499 7406 16508
rect 7073 16457 7086 16499
rect 7138 16457 7151 16499
rect 7203 16457 7216 16499
rect 7268 16457 7281 16499
rect 7333 16457 7346 16499
rect 7398 16457 7411 16499
rect 7080 16456 7086 16457
rect 7333 16456 7334 16457
rect 7398 16456 7406 16457
rect 7463 16456 7476 16508
rect 7528 16456 7541 16508
rect 7593 16456 7606 16508
rect 7658 16456 7671 16508
rect 7728 16499 7736 16508
rect 7800 16499 7801 16508
rect 7872 16499 7884 16533
rect 7723 16457 7736 16499
rect 7788 16457 7801 16499
rect 7853 16457 7884 16499
rect 7728 16456 7736 16457
rect 7800 16456 7801 16457
rect 5123 16442 5162 16456
rect 5196 16442 5235 16456
rect 5269 16442 5308 16456
rect 5342 16442 5381 16456
rect 5415 16442 5454 16456
rect 5488 16442 5527 16456
rect 5561 16442 5600 16456
rect 5634 16442 5673 16456
rect 5707 16442 5746 16456
rect 5780 16442 5819 16456
rect 5853 16442 5892 16456
rect 5926 16442 5965 16456
rect 5999 16442 6038 16456
rect 6072 16442 6110 16456
rect 6144 16442 6182 16456
rect 6216 16442 6254 16456
rect 6288 16442 6326 16456
rect 6360 16442 6398 16456
rect 6432 16442 6470 16456
rect 6504 16442 6542 16456
rect 6576 16442 6614 16456
rect 6648 16442 6686 16456
rect 6720 16442 6758 16456
rect 6792 16442 6830 16456
rect 6864 16442 6902 16456
rect 6936 16442 6974 16456
rect 7008 16442 7046 16456
rect 7080 16442 7118 16456
rect 7152 16442 7190 16456
rect 7224 16442 7262 16456
rect 7296 16442 7334 16456
rect 7368 16442 7406 16456
rect 7440 16442 7478 16456
rect 7512 16442 7550 16456
rect 7584 16442 7622 16456
rect 7656 16442 7694 16456
rect 7728 16442 7766 16456
rect 7800 16442 7838 16456
rect 5234 16423 5235 16442
rect 5300 16423 5308 16442
rect 5077 16390 5116 16423
rect 5168 16390 5182 16423
rect 5234 16390 5248 16423
rect 5300 16390 5314 16423
rect 5366 16390 5380 16442
rect 5432 16390 5446 16442
rect 5498 16390 5512 16442
rect 5564 16390 5578 16442
rect 5634 16423 5644 16442
rect 5707 16423 5710 16442
rect 5960 16423 5965 16442
rect 6026 16423 6038 16442
rect 5630 16390 5644 16423
rect 5696 16390 5710 16423
rect 5762 16390 5776 16423
rect 5828 16390 5842 16423
rect 5894 16390 5908 16423
rect 5960 16390 5974 16423
rect 6026 16390 6040 16423
rect 6092 16390 6106 16442
rect 6158 16390 6172 16442
rect 6224 16390 6238 16442
rect 6290 16390 6304 16442
rect 6360 16423 6370 16442
rect 6432 16423 6436 16442
rect 6683 16423 6686 16442
rect 6748 16423 6758 16442
rect 6356 16390 6370 16423
rect 6422 16390 6436 16423
rect 6488 16390 6501 16423
rect 6553 16390 6566 16423
rect 6618 16390 6631 16423
rect 6683 16390 6696 16423
rect 6748 16390 6761 16423
rect 6813 16390 6826 16442
rect 6878 16390 6891 16442
rect 6943 16390 6956 16442
rect 7008 16390 7021 16442
rect 7080 16423 7086 16442
rect 7333 16423 7334 16442
rect 7398 16423 7406 16442
rect 7073 16390 7086 16423
rect 7138 16390 7151 16423
rect 7203 16390 7216 16423
rect 7268 16390 7281 16423
rect 7333 16390 7346 16423
rect 7398 16390 7411 16423
rect 7463 16390 7476 16442
rect 7528 16390 7541 16442
rect 7593 16390 7606 16442
rect 7658 16390 7671 16442
rect 7728 16423 7736 16442
rect 7800 16423 7801 16442
rect 7872 16423 7884 16457
rect 7723 16390 7736 16423
rect 7788 16390 7801 16423
rect 7853 16390 7884 16423
rect 5077 16381 7884 16390
rect 5077 16347 5089 16381
rect 5123 16376 5162 16381
rect 5196 16376 5235 16381
rect 5269 16376 5308 16381
rect 5342 16376 5381 16381
rect 5415 16376 5454 16381
rect 5488 16376 5527 16381
rect 5561 16376 5600 16381
rect 5634 16376 5673 16381
rect 5707 16376 5746 16381
rect 5780 16376 5819 16381
rect 5853 16376 5892 16381
rect 5926 16376 5965 16381
rect 5999 16376 6038 16381
rect 6072 16376 6110 16381
rect 6144 16376 6182 16381
rect 6216 16376 6254 16381
rect 6288 16376 6326 16381
rect 6360 16376 6398 16381
rect 6432 16376 6470 16381
rect 6504 16376 6542 16381
rect 6576 16376 6614 16381
rect 6648 16376 6686 16381
rect 6720 16376 6758 16381
rect 6792 16376 6830 16381
rect 6864 16376 6902 16381
rect 6936 16376 6974 16381
rect 7008 16376 7046 16381
rect 7080 16376 7118 16381
rect 7152 16376 7190 16381
rect 7224 16376 7262 16381
rect 7296 16376 7334 16381
rect 7368 16376 7406 16381
rect 7440 16376 7478 16381
rect 7512 16376 7550 16381
rect 7584 16376 7622 16381
rect 7656 16376 7694 16381
rect 7728 16376 7766 16381
rect 7800 16376 7838 16381
rect 5234 16347 5235 16376
rect 5300 16347 5308 16376
rect 5077 16324 5116 16347
rect 5168 16324 5182 16347
rect 5234 16324 5248 16347
rect 5300 16324 5314 16347
rect 5366 16324 5380 16376
rect 5432 16324 5446 16376
rect 5498 16324 5512 16376
rect 5564 16324 5578 16376
rect 5634 16347 5644 16376
rect 5707 16347 5710 16376
rect 5960 16347 5965 16376
rect 6026 16347 6038 16376
rect 5630 16324 5644 16347
rect 5696 16324 5710 16347
rect 5762 16324 5776 16347
rect 5828 16324 5842 16347
rect 5894 16324 5908 16347
rect 5960 16324 5974 16347
rect 6026 16324 6040 16347
rect 6092 16324 6106 16376
rect 6158 16324 6172 16376
rect 6224 16324 6238 16376
rect 6290 16324 6304 16376
rect 6360 16347 6370 16376
rect 6432 16347 6436 16376
rect 6683 16347 6686 16376
rect 6748 16347 6758 16376
rect 6356 16324 6370 16347
rect 6422 16324 6436 16347
rect 6488 16324 6501 16347
rect 6553 16324 6566 16347
rect 6618 16324 6631 16347
rect 6683 16324 6696 16347
rect 6748 16324 6761 16347
rect 6813 16324 6826 16376
rect 6878 16324 6891 16376
rect 6943 16324 6956 16376
rect 7008 16324 7021 16376
rect 7080 16347 7086 16376
rect 7333 16347 7334 16376
rect 7398 16347 7406 16376
rect 7073 16324 7086 16347
rect 7138 16324 7151 16347
rect 7203 16324 7216 16347
rect 7268 16324 7281 16347
rect 7333 16324 7346 16347
rect 7398 16324 7411 16347
rect 7463 16324 7476 16376
rect 7528 16324 7541 16376
rect 7593 16324 7606 16376
rect 7658 16324 7671 16376
rect 7728 16347 7736 16376
rect 7800 16347 7801 16376
rect 7872 16347 7884 16381
rect 7723 16324 7736 16347
rect 7788 16324 7801 16347
rect 7853 16324 7884 16347
rect 5077 16310 7884 16324
rect 5077 16305 5116 16310
rect 5168 16305 5182 16310
rect 5234 16305 5248 16310
rect 5300 16305 5314 16310
rect 5077 16271 5089 16305
rect 5234 16271 5235 16305
rect 5300 16271 5308 16305
rect 5077 16258 5116 16271
rect 5168 16258 5182 16271
rect 5234 16258 5248 16271
rect 5300 16258 5314 16271
rect 5366 16258 5380 16310
rect 5432 16258 5446 16310
rect 5498 16258 5512 16310
rect 5564 16258 5578 16310
rect 5630 16305 5644 16310
rect 5696 16305 5710 16310
rect 5762 16305 5776 16310
rect 5828 16305 5842 16310
rect 5894 16305 5908 16310
rect 5960 16305 5974 16310
rect 6026 16305 6040 16310
rect 5634 16271 5644 16305
rect 5707 16271 5710 16305
rect 5960 16271 5965 16305
rect 6026 16271 6038 16305
rect 5630 16258 5644 16271
rect 5696 16258 5710 16271
rect 5762 16258 5776 16271
rect 5828 16258 5842 16271
rect 5894 16258 5908 16271
rect 5960 16258 5974 16271
rect 6026 16258 6040 16271
rect 6092 16258 6106 16310
rect 6158 16258 6172 16310
rect 6224 16258 6238 16310
rect 6290 16258 6304 16310
rect 6356 16305 6370 16310
rect 6422 16305 6436 16310
rect 6488 16305 6501 16310
rect 6553 16305 6566 16310
rect 6618 16305 6631 16310
rect 6683 16305 6696 16310
rect 6748 16305 6761 16310
rect 6360 16271 6370 16305
rect 6432 16271 6436 16305
rect 6683 16271 6686 16305
rect 6748 16271 6758 16305
rect 6356 16258 6370 16271
rect 6422 16258 6436 16271
rect 6488 16258 6501 16271
rect 6553 16258 6566 16271
rect 6618 16258 6631 16271
rect 6683 16258 6696 16271
rect 6748 16258 6761 16271
rect 6813 16258 6826 16310
rect 6878 16258 6891 16310
rect 6943 16258 6956 16310
rect 7008 16258 7021 16310
rect 7073 16305 7086 16310
rect 7138 16305 7151 16310
rect 7203 16305 7216 16310
rect 7268 16305 7281 16310
rect 7333 16305 7346 16310
rect 7398 16305 7411 16310
rect 7080 16271 7086 16305
rect 7333 16271 7334 16305
rect 7398 16271 7406 16305
rect 7073 16258 7086 16271
rect 7138 16258 7151 16271
rect 7203 16258 7216 16271
rect 7268 16258 7281 16271
rect 7333 16258 7346 16271
rect 7398 16258 7411 16271
rect 7463 16258 7476 16310
rect 7528 16258 7541 16310
rect 7593 16258 7606 16310
rect 7658 16258 7671 16310
rect 7723 16305 7736 16310
rect 7788 16305 7801 16310
rect 7853 16305 7884 16310
rect 7728 16271 7736 16305
rect 7800 16271 7801 16305
rect 7872 16271 7884 16305
rect 7723 16258 7736 16271
rect 7788 16258 7801 16271
rect 7853 16258 7884 16271
rect 5077 16244 7884 16258
rect 5077 16229 5116 16244
rect 5168 16229 5182 16244
rect 5234 16229 5248 16244
rect 5300 16229 5314 16244
rect 5077 16195 5089 16229
rect 5234 16195 5235 16229
rect 5300 16195 5308 16229
rect 5077 16192 5116 16195
rect 5168 16192 5182 16195
rect 5234 16192 5248 16195
rect 5300 16192 5314 16195
rect 5366 16192 5380 16244
rect 5432 16192 5446 16244
rect 5498 16192 5512 16244
rect 5564 16192 5578 16244
rect 5630 16229 5644 16244
rect 5696 16229 5710 16244
rect 5762 16229 5776 16244
rect 5828 16229 5842 16244
rect 5894 16229 5908 16244
rect 5960 16229 5974 16244
rect 6026 16229 6040 16244
rect 5634 16195 5644 16229
rect 5707 16195 5710 16229
rect 5960 16195 5965 16229
rect 6026 16195 6038 16229
rect 5630 16192 5644 16195
rect 5696 16192 5710 16195
rect 5762 16192 5776 16195
rect 5828 16192 5842 16195
rect 5894 16192 5908 16195
rect 5960 16192 5974 16195
rect 6026 16192 6040 16195
rect 6092 16192 6106 16244
rect 6158 16192 6172 16244
rect 6224 16192 6238 16244
rect 6290 16192 6304 16244
rect 6356 16229 6370 16244
rect 6422 16229 6436 16244
rect 6488 16229 6501 16244
rect 6553 16229 6566 16244
rect 6618 16229 6631 16244
rect 6683 16229 6696 16244
rect 6748 16229 6761 16244
rect 6360 16195 6370 16229
rect 6432 16195 6436 16229
rect 6683 16195 6686 16229
rect 6748 16195 6758 16229
rect 6356 16192 6370 16195
rect 6422 16192 6436 16195
rect 6488 16192 6501 16195
rect 6553 16192 6566 16195
rect 6618 16192 6631 16195
rect 6683 16192 6696 16195
rect 6748 16192 6761 16195
rect 6813 16192 6826 16244
rect 6878 16192 6891 16244
rect 6943 16192 6956 16244
rect 7008 16192 7021 16244
rect 7073 16229 7086 16244
rect 7138 16229 7151 16244
rect 7203 16229 7216 16244
rect 7268 16229 7281 16244
rect 7333 16229 7346 16244
rect 7398 16229 7411 16244
rect 7080 16195 7086 16229
rect 7333 16195 7334 16229
rect 7398 16195 7406 16229
rect 7073 16192 7086 16195
rect 7138 16192 7151 16195
rect 7203 16192 7216 16195
rect 7268 16192 7281 16195
rect 7333 16192 7346 16195
rect 7398 16192 7411 16195
rect 7463 16192 7476 16244
rect 7528 16192 7541 16244
rect 7593 16192 7606 16244
rect 7658 16192 7671 16244
rect 7723 16229 7736 16244
rect 7788 16229 7801 16244
rect 7853 16229 7884 16244
rect 7728 16195 7736 16229
rect 7800 16195 7801 16229
rect 7872 16195 7884 16229
rect 7723 16192 7736 16195
rect 7788 16192 7801 16195
rect 7853 16192 7884 16195
rect 5077 16178 7884 16192
rect 5077 16153 5116 16178
rect 5168 16153 5182 16178
rect 5234 16153 5248 16178
rect 5300 16153 5314 16178
rect 5077 16119 5089 16153
rect 5234 16126 5235 16153
rect 5300 16126 5308 16153
rect 5366 16126 5380 16178
rect 5432 16126 5446 16178
rect 5498 16126 5512 16178
rect 5564 16126 5578 16178
rect 5630 16153 5644 16178
rect 5696 16153 5710 16178
rect 5762 16153 5776 16178
rect 5828 16153 5842 16178
rect 5894 16153 5908 16178
rect 5960 16153 5974 16178
rect 6026 16153 6040 16178
rect 5634 16126 5644 16153
rect 5707 16126 5710 16153
rect 5960 16126 5965 16153
rect 6026 16126 6038 16153
rect 6092 16126 6106 16178
rect 6158 16126 6172 16178
rect 6224 16126 6238 16178
rect 6290 16126 6304 16178
rect 6356 16153 6370 16178
rect 6422 16153 6436 16178
rect 6488 16153 6501 16178
rect 6553 16153 6566 16178
rect 6618 16153 6631 16178
rect 6683 16153 6696 16178
rect 6748 16153 6761 16178
rect 6360 16126 6370 16153
rect 6432 16126 6436 16153
rect 6683 16126 6686 16153
rect 6748 16126 6758 16153
rect 6813 16126 6826 16178
rect 6878 16126 6891 16178
rect 6943 16126 6956 16178
rect 7008 16126 7021 16178
rect 7073 16153 7086 16178
rect 7138 16153 7151 16178
rect 7203 16153 7216 16178
rect 7268 16153 7281 16178
rect 7333 16153 7346 16178
rect 7398 16153 7411 16178
rect 7080 16126 7086 16153
rect 7333 16126 7334 16153
rect 7398 16126 7406 16153
rect 7463 16126 7476 16178
rect 7528 16126 7541 16178
rect 7593 16126 7606 16178
rect 7658 16126 7671 16178
rect 7723 16153 7736 16178
rect 7788 16153 7801 16178
rect 7853 16153 7884 16178
rect 7728 16126 7736 16153
rect 7800 16126 7801 16153
rect 5123 16119 5162 16126
rect 5196 16119 5235 16126
rect 5269 16119 5308 16126
rect 5342 16119 5381 16126
rect 5415 16119 5454 16126
rect 5488 16119 5527 16126
rect 5561 16119 5600 16126
rect 5634 16119 5673 16126
rect 5707 16119 5746 16126
rect 5780 16119 5819 16126
rect 5853 16119 5892 16126
rect 5926 16119 5965 16126
rect 5999 16119 6038 16126
rect 6072 16119 6110 16126
rect 6144 16119 6182 16126
rect 6216 16119 6254 16126
rect 6288 16119 6326 16126
rect 6360 16119 6398 16126
rect 6432 16119 6470 16126
rect 6504 16119 6542 16126
rect 6576 16119 6614 16126
rect 6648 16119 6686 16126
rect 6720 16119 6758 16126
rect 6792 16119 6830 16126
rect 6864 16119 6902 16126
rect 6936 16119 6974 16126
rect 7008 16119 7046 16126
rect 7080 16119 7118 16126
rect 7152 16119 7190 16126
rect 7224 16119 7262 16126
rect 7296 16119 7334 16126
rect 7368 16119 7406 16126
rect 7440 16119 7478 16126
rect 7512 16119 7550 16126
rect 7584 16119 7622 16126
rect 7656 16119 7694 16126
rect 7728 16119 7766 16126
rect 7800 16119 7838 16126
rect 7872 16119 7884 16153
rect 5077 16112 7884 16119
rect 5077 16077 5116 16112
rect 5168 16077 5182 16112
rect 5234 16077 5248 16112
rect 5300 16077 5314 16112
rect 5077 16043 5089 16077
rect 5234 16060 5235 16077
rect 5300 16060 5308 16077
rect 5366 16060 5380 16112
rect 5432 16060 5446 16112
rect 5498 16060 5512 16112
rect 5564 16060 5578 16112
rect 5630 16077 5644 16112
rect 5696 16077 5710 16112
rect 5762 16077 5776 16112
rect 5828 16077 5842 16112
rect 5894 16077 5908 16112
rect 5960 16077 5974 16112
rect 6026 16077 6040 16112
rect 5634 16060 5644 16077
rect 5707 16060 5710 16077
rect 5960 16060 5965 16077
rect 6026 16060 6038 16077
rect 6092 16060 6106 16112
rect 6158 16060 6172 16112
rect 6224 16060 6238 16112
rect 6290 16060 6304 16112
rect 6356 16077 6370 16112
rect 6422 16077 6436 16112
rect 6488 16077 6501 16112
rect 6553 16077 6566 16112
rect 6618 16077 6631 16112
rect 6683 16077 6696 16112
rect 6748 16077 6761 16112
rect 6360 16060 6370 16077
rect 6432 16060 6436 16077
rect 6683 16060 6686 16077
rect 6748 16060 6758 16077
rect 6813 16060 6826 16112
rect 6878 16060 6891 16112
rect 6943 16060 6956 16112
rect 7008 16060 7021 16112
rect 7073 16077 7086 16112
rect 7138 16077 7151 16112
rect 7203 16077 7216 16112
rect 7268 16077 7281 16112
rect 7333 16077 7346 16112
rect 7398 16077 7411 16112
rect 7080 16060 7086 16077
rect 7333 16060 7334 16077
rect 7398 16060 7406 16077
rect 7463 16060 7476 16112
rect 7528 16060 7541 16112
rect 7593 16060 7606 16112
rect 7658 16060 7671 16112
rect 7723 16077 7736 16112
rect 7788 16077 7801 16112
rect 7853 16077 7884 16112
rect 7728 16060 7736 16077
rect 7800 16060 7801 16077
rect 5123 16046 5162 16060
rect 5196 16046 5235 16060
rect 5269 16046 5308 16060
rect 5342 16046 5381 16060
rect 5415 16046 5454 16060
rect 5488 16046 5527 16060
rect 5561 16046 5600 16060
rect 5634 16046 5673 16060
rect 5707 16046 5746 16060
rect 5780 16046 5819 16060
rect 5853 16046 5892 16060
rect 5926 16046 5965 16060
rect 5999 16046 6038 16060
rect 6072 16046 6110 16060
rect 6144 16046 6182 16060
rect 6216 16046 6254 16060
rect 6288 16046 6326 16060
rect 6360 16046 6398 16060
rect 6432 16046 6470 16060
rect 6504 16046 6542 16060
rect 6576 16046 6614 16060
rect 6648 16046 6686 16060
rect 6720 16046 6758 16060
rect 6792 16046 6830 16060
rect 6864 16046 6902 16060
rect 6936 16046 6974 16060
rect 7008 16046 7046 16060
rect 7080 16046 7118 16060
rect 7152 16046 7190 16060
rect 7224 16046 7262 16060
rect 7296 16046 7334 16060
rect 7368 16046 7406 16060
rect 7440 16046 7478 16060
rect 7512 16046 7550 16060
rect 7584 16046 7622 16060
rect 7656 16046 7694 16060
rect 7728 16046 7766 16060
rect 7800 16046 7838 16060
rect 5234 16043 5235 16046
rect 5300 16043 5308 16046
rect 5077 16001 5116 16043
rect 5168 16001 5182 16043
rect 5234 16001 5248 16043
rect 5300 16001 5314 16043
rect 5077 15967 5089 16001
rect 5234 15994 5235 16001
rect 5300 15994 5308 16001
rect 5366 15994 5380 16046
rect 5432 15994 5446 16046
rect 5498 15994 5512 16046
rect 5564 15994 5578 16046
rect 5634 16043 5644 16046
rect 5707 16043 5710 16046
rect 5960 16043 5965 16046
rect 6026 16043 6038 16046
rect 5630 16001 5644 16043
rect 5696 16001 5710 16043
rect 5762 16001 5776 16043
rect 5828 16001 5842 16043
rect 5894 16001 5908 16043
rect 5960 16001 5974 16043
rect 6026 16001 6040 16043
rect 5634 15994 5644 16001
rect 5707 15994 5710 16001
rect 5960 15994 5965 16001
rect 6026 15994 6038 16001
rect 6092 15994 6106 16046
rect 6158 15994 6172 16046
rect 6224 15994 6238 16046
rect 6290 15994 6304 16046
rect 6360 16043 6370 16046
rect 6432 16043 6436 16046
rect 6683 16043 6686 16046
rect 6748 16043 6758 16046
rect 6356 16001 6370 16043
rect 6422 16001 6436 16043
rect 6488 16001 6501 16043
rect 6553 16001 6566 16043
rect 6618 16001 6631 16043
rect 6683 16001 6696 16043
rect 6748 16001 6761 16043
rect 6360 15994 6370 16001
rect 6432 15994 6436 16001
rect 6683 15994 6686 16001
rect 6748 15994 6758 16001
rect 6813 15994 6826 16046
rect 6878 15994 6891 16046
rect 6943 15994 6956 16046
rect 7008 15994 7021 16046
rect 7080 16043 7086 16046
rect 7333 16043 7334 16046
rect 7398 16043 7406 16046
rect 7073 16001 7086 16043
rect 7138 16001 7151 16043
rect 7203 16001 7216 16043
rect 7268 16001 7281 16043
rect 7333 16001 7346 16043
rect 7398 16001 7411 16043
rect 7080 15994 7086 16001
rect 7333 15994 7334 16001
rect 7398 15994 7406 16001
rect 7463 15994 7476 16046
rect 7528 15994 7541 16046
rect 7593 15994 7606 16046
rect 7658 15994 7671 16046
rect 7728 16043 7736 16046
rect 7800 16043 7801 16046
rect 7872 16043 7884 16077
rect 7723 16001 7736 16043
rect 7788 16001 7801 16043
rect 7853 16001 7884 16043
rect 7728 15994 7736 16001
rect 7800 15994 7801 16001
rect 5123 15967 5162 15994
rect 5196 15967 5235 15994
rect 5269 15967 5308 15994
rect 5342 15967 5381 15994
rect 5415 15967 5454 15994
rect 5488 15967 5527 15994
rect 5561 15967 5600 15994
rect 5634 15967 5673 15994
rect 5707 15967 5746 15994
rect 5780 15967 5819 15994
rect 5853 15967 5892 15994
rect 5926 15967 5965 15994
rect 5999 15967 6038 15994
rect 6072 15967 6110 15994
rect 6144 15967 6182 15994
rect 6216 15967 6254 15994
rect 6288 15967 6326 15994
rect 6360 15967 6398 15994
rect 6432 15967 6470 15994
rect 6504 15967 6542 15994
rect 6576 15967 6614 15994
rect 6648 15967 6686 15994
rect 6720 15967 6758 15994
rect 6792 15967 6830 15994
rect 6864 15967 6902 15994
rect 6936 15967 6974 15994
rect 7008 15967 7046 15994
rect 7080 15967 7118 15994
rect 7152 15967 7190 15994
rect 7224 15967 7262 15994
rect 7296 15967 7334 15994
rect 7368 15967 7406 15994
rect 7440 15967 7478 15994
rect 7512 15967 7550 15994
rect 7584 15967 7622 15994
rect 7656 15967 7694 15994
rect 7728 15967 7766 15994
rect 7800 15967 7838 15994
rect 7872 15967 7884 16001
rect 5077 15952 7884 15967
rect 8044 17003 8184 17013
rect 8218 17003 8224 17037
rect 8044 16975 8224 17003
rect 8044 16973 8050 16975
rect 8084 16973 8224 16975
rect 8044 16921 8047 16973
rect 8099 16921 8169 16973
rect 8221 16921 8224 16973
rect 8044 16907 8224 16921
rect 8044 16855 8047 16907
rect 8099 16855 8169 16907
rect 8221 16855 8224 16907
rect 8044 16841 8224 16855
rect 8044 16789 8047 16841
rect 8099 16789 8169 16841
rect 8221 16789 8224 16841
rect 8044 16787 8184 16789
rect 8218 16787 8224 16789
rect 8044 16775 8224 16787
rect 8044 16723 8047 16775
rect 8099 16723 8169 16775
rect 8221 16723 8224 16775
rect 8044 16715 8184 16723
rect 8218 16715 8224 16723
rect 8044 16709 8224 16715
rect 8044 16657 8047 16709
rect 8099 16657 8169 16709
rect 8221 16657 8224 16709
rect 8044 16653 8050 16657
rect 8084 16653 8184 16657
rect 8044 16643 8184 16653
rect 8218 16643 8224 16657
rect 8044 16591 8047 16643
rect 8099 16591 8169 16643
rect 8221 16591 8224 16643
rect 8044 16581 8050 16591
rect 8084 16581 8184 16591
rect 8044 16577 8184 16581
rect 8218 16577 8224 16591
rect 8044 16525 8047 16577
rect 8099 16525 8169 16577
rect 8221 16525 8224 16577
rect 8044 16511 8050 16525
rect 8084 16511 8184 16525
rect 8218 16511 8224 16525
rect 8044 16459 8047 16511
rect 8099 16459 8169 16511
rect 8221 16459 8224 16511
rect 8044 16445 8050 16459
rect 8084 16445 8184 16459
rect 8218 16445 8224 16459
rect 8044 16393 8047 16445
rect 8099 16393 8169 16445
rect 8221 16393 8224 16445
rect 8044 16378 8050 16393
rect 8084 16389 8224 16393
rect 8084 16378 8184 16389
rect 8218 16378 8224 16389
rect 8044 16326 8047 16378
rect 8099 16326 8169 16378
rect 8221 16326 8224 16378
rect 8044 16311 8050 16326
rect 8084 16317 8224 16326
rect 8084 16311 8184 16317
rect 8218 16311 8224 16317
rect 8044 16259 8047 16311
rect 8099 16259 8169 16311
rect 8221 16259 8224 16311
rect 8044 16255 8224 16259
rect 8044 16244 8050 16255
rect 8084 16245 8224 16255
rect 8084 16244 8184 16245
rect 8218 16244 8224 16245
rect 8044 16192 8047 16244
rect 8099 16192 8169 16244
rect 8221 16192 8224 16244
rect 8044 16183 8224 16192
rect 8044 16177 8050 16183
rect 8084 16177 8224 16183
rect 8044 16125 8047 16177
rect 8099 16125 8169 16177
rect 8221 16125 8224 16177
rect 8044 16111 8224 16125
rect 8044 16110 8050 16111
rect 8084 16110 8224 16111
rect 8044 16058 8047 16110
rect 8099 16058 8169 16110
rect 8221 16058 8224 16110
rect 8044 16043 8224 16058
rect 8044 15991 8047 16043
rect 8099 15991 8169 16043
rect 8221 15991 8224 16043
rect 8044 15967 8224 15991
rect 8044 15933 8050 15967
rect 8084 15957 8224 15967
rect 8084 15933 8184 15957
rect 8044 15923 8184 15933
rect 8218 15923 8224 15957
rect 8044 15895 8224 15923
rect 8044 15861 8050 15895
rect 8084 15885 8224 15895
rect 8084 15861 8184 15885
rect 8044 15851 8184 15861
rect 8218 15851 8224 15885
rect 8044 15823 8224 15851
rect 8044 15789 8050 15823
rect 8084 15813 8224 15823
rect 8084 15789 8184 15813
rect 8044 15779 8184 15789
rect 8218 15779 8224 15813
rect 8044 15751 8224 15779
rect 8044 15717 8050 15751
rect 8084 15741 8224 15751
rect 8084 15717 8184 15741
rect 8044 15707 8184 15717
rect 8218 15707 8224 15741
tri 4928 15679 4940 15691 sw
rect 8044 15679 8224 15707
rect 2270 15636 2450 15674
tri 4738 15660 4757 15679 se
rect 4757 15665 4940 15679
tri 4940 15665 4954 15679 sw
rect 4757 15660 7729 15665
rect 2270 15602 2276 15636
rect 2310 15602 2410 15636
rect 2444 15602 2450 15636
rect 2270 15564 2450 15602
rect 2270 15530 2276 15564
rect 2310 15530 2410 15564
rect 2444 15530 2450 15564
rect 2270 15492 2450 15530
rect 2270 15458 2276 15492
rect 2310 15458 2410 15492
rect 2444 15458 2450 15492
rect 2270 15456 2450 15458
rect 2322 15404 2392 15456
rect 2270 15387 2276 15404
rect 2310 15387 2410 15404
rect 2322 15335 2392 15387
rect 2270 15318 2276 15335
rect 2310 15318 2410 15335
rect 2322 15266 2392 15318
rect 2270 15249 2276 15266
rect 2310 15249 2410 15266
rect 2322 15197 2392 15249
rect 2270 15180 2276 15197
rect 2310 15180 2410 15197
rect 2322 15128 2392 15180
rect 2270 15110 2276 15128
rect 2310 15110 2410 15128
rect 2322 15058 2392 15110
rect 2270 15040 2276 15058
rect 2310 15040 2410 15058
rect 2322 14988 2392 15040
rect 2270 14970 2276 14988
rect 2310 14970 2410 14988
rect 2322 14918 2392 14970
rect 2444 14918 2450 15456
rect 2270 14916 2450 14918
rect 2270 14900 2276 14916
rect 2310 14900 2410 14916
rect 2322 14848 2392 14900
rect 2444 14848 2450 14916
rect 2270 14844 2450 14848
rect 2270 14810 2276 14844
rect 2310 14810 2410 14844
rect 2444 14810 2450 14844
rect 2270 14772 2450 14810
rect 2270 14738 2276 14772
rect 2310 14738 2410 14772
rect 2444 14738 2450 14772
rect 2270 14700 2450 14738
rect 2270 14666 2276 14700
rect 2310 14666 2410 14700
rect 2444 14666 2450 14700
rect 2270 14628 2450 14666
rect 2270 14594 2276 14628
rect 2310 14594 2410 14628
rect 2444 14594 2450 14628
rect 2270 14556 2450 14594
rect 2270 14522 2276 14556
rect 2310 14522 2410 14556
rect 2444 14522 2450 14556
rect 2270 14484 2450 14522
rect 2270 14450 2276 14484
rect 2310 14450 2410 14484
rect 2444 14450 2450 14484
rect 2270 14412 2450 14450
rect 2270 14378 2276 14412
rect 2310 14378 2410 14412
rect 2444 14378 2450 14412
rect 2270 14340 2450 14378
rect 2270 14306 2276 14340
rect 2310 14306 2410 14340
rect 2444 14306 2450 14340
rect 2270 14268 2450 14306
rect 2270 14234 2276 14268
rect 2310 14234 2410 14268
rect 2444 14234 2450 14268
rect 2270 14196 2450 14234
rect 2270 14162 2276 14196
rect 2310 14162 2410 14196
rect 2444 14162 2450 14196
rect 2270 14124 2450 14162
rect 2270 14090 2276 14124
rect 2310 14090 2410 14124
rect 2444 14090 2450 14124
rect 2270 14052 2450 14090
rect 2270 14018 2276 14052
rect 2310 14018 2410 14052
rect 2444 14018 2450 14052
rect 2270 13980 2450 14018
rect 2270 13946 2276 13980
rect 2310 13946 2410 13980
rect 2444 13946 2450 13980
rect 2270 13908 2450 13946
rect 2270 13874 2276 13908
rect 2310 13874 2410 13908
rect 2444 13874 2450 13908
rect 2270 13836 2450 13874
rect 2270 13802 2276 13836
rect 2310 13802 2410 13836
rect 2444 13802 2450 13836
rect 2270 13764 2450 13802
rect 2270 13730 2276 13764
rect 2310 13730 2410 13764
rect 2444 13730 2450 13764
rect 2270 13692 2450 13730
rect 2270 13658 2276 13692
rect 2310 13658 2410 13692
rect 2444 13658 2450 13692
rect 2270 13620 2450 13658
rect 2270 13586 2276 13620
rect 2310 13586 2410 13620
rect 2444 13586 2450 13620
rect 2270 13548 2450 13586
rect 2270 13514 2276 13548
rect 2310 13514 2410 13548
rect 2444 13514 2450 13548
rect 2270 13476 2450 13514
rect 2270 13456 2276 13476
rect 2310 13456 2410 13476
rect 2322 13404 2392 13456
rect 2270 13387 2276 13404
rect 2310 13387 2410 13404
rect 2322 13335 2392 13387
rect 2444 13335 2450 13476
rect 2270 13332 2450 13335
rect 2270 13318 2276 13332
rect 2310 13318 2410 13332
rect 2322 13266 2392 13318
rect 2444 13266 2450 13332
rect 2270 13260 2450 13266
rect 2270 13249 2276 13260
rect 2310 13249 2410 13260
rect 2322 13197 2392 13249
rect 2444 13197 2450 13260
rect 2270 13188 2450 13197
rect 2270 13180 2276 13188
rect 2310 13180 2410 13188
rect 2322 13128 2392 13180
rect 2444 13128 2450 13188
rect 2270 13116 2450 13128
rect 2270 13110 2276 13116
rect 2310 13110 2410 13116
rect 2322 13058 2392 13110
rect 2444 13058 2450 13116
rect 2270 13044 2450 13058
rect 2270 13040 2276 13044
rect 2310 13040 2410 13044
rect 2322 12988 2392 13040
rect 2444 12988 2450 13044
rect 2270 12972 2450 12988
rect 2270 12970 2276 12972
rect 2310 12970 2410 12972
rect 2322 12918 2392 12970
rect 2444 12918 2450 12972
rect 2270 12900 2450 12918
rect 2322 12848 2392 12900
rect 2444 12848 2450 12900
rect 2270 12828 2450 12848
rect 2270 12794 2276 12828
rect 2310 12794 2410 12828
rect 2444 12794 2450 12828
rect 2270 12756 2450 12794
rect 2270 12722 2276 12756
rect 2310 12722 2410 12756
rect 2444 12722 2450 12756
rect 2270 12684 2450 12722
rect 2270 12650 2276 12684
rect 2310 12650 2410 12684
rect 2444 12650 2450 12684
rect 2270 12612 2450 12650
rect 2270 12578 2276 12612
rect 2310 12578 2410 12612
rect 2444 12578 2450 12612
rect 2270 12540 2450 12578
rect 2270 12506 2276 12540
rect 2310 12506 2410 12540
rect 2444 12506 2450 12540
rect 2270 12468 2450 12506
rect 2270 12434 2276 12468
rect 2310 12434 2410 12468
rect 2444 12434 2450 12468
rect 2270 12396 2450 12434
rect 2270 12362 2276 12396
rect 2310 12362 2410 12396
rect 2444 12362 2450 12396
rect 2270 12324 2450 12362
rect 2270 12290 2276 12324
rect 2310 12290 2410 12324
rect 2444 12290 2450 12324
rect 2270 12252 2450 12290
rect 2270 12218 2276 12252
rect 2310 12218 2410 12252
rect 2444 12218 2450 12252
rect 2270 12180 2450 12218
rect 2270 12146 2276 12180
rect 2310 12146 2410 12180
rect 2444 12146 2450 12180
rect 2270 12108 2450 12146
rect 2270 12074 2276 12108
rect 2310 12074 2410 12108
rect 2444 12074 2450 12108
rect 2270 12036 2450 12074
rect 2270 12002 2276 12036
rect 2310 12002 2410 12036
rect 2444 12002 2450 12036
rect 2270 11964 2450 12002
rect 2270 11930 2276 11964
rect 2310 11930 2410 11964
rect 2444 11930 2450 11964
rect 2270 11892 2450 11930
rect 2270 11858 2276 11892
rect 2310 11858 2410 11892
rect 2444 11858 2450 11892
rect 2270 11820 2450 11858
rect 2270 11786 2276 11820
rect 2310 11786 2410 11820
rect 2444 11786 2450 11820
rect 2270 11748 2450 11786
rect 2270 11714 2276 11748
rect 2310 11714 2410 11748
rect 2444 11714 2450 11748
rect 2270 11676 2450 11714
rect 2270 11642 2276 11676
rect 2310 11642 2410 11676
rect 2444 11642 2450 11676
rect 2270 11604 2450 11642
rect 2270 11570 2276 11604
rect 2310 11570 2410 11604
rect 2444 11570 2450 11604
rect 2270 11532 2450 11570
rect 2270 11498 2276 11532
rect 2310 11498 2410 11532
rect 2444 11498 2450 11532
rect 2270 11460 2450 11498
rect 2270 11456 2276 11460
rect 2310 11456 2410 11460
rect 2322 11404 2392 11456
rect 2444 11404 2450 11460
rect 2270 11388 2450 11404
rect 2270 11387 2276 11388
rect 2310 11387 2410 11388
rect 2322 11335 2392 11387
rect 2444 11335 2450 11388
rect 2270 11318 2450 11335
rect 2322 11266 2392 11318
rect 2444 11266 2450 11318
rect 2270 11249 2450 11266
rect 2322 11197 2392 11249
rect 2444 11197 2450 11249
rect 2270 11180 2450 11197
rect 2322 11128 2392 11180
rect 2444 11128 2450 11180
rect 2270 11110 2450 11128
rect 2322 11058 2392 11110
rect 2444 11058 2450 11110
rect 2270 11040 2450 11058
rect 2322 10988 2392 11040
rect 2444 10988 2450 11040
rect 2270 10970 2450 10988
rect 2322 10918 2392 10970
rect 2444 10918 2450 10970
rect 2270 10900 2450 10918
rect 2322 10848 2392 10900
rect 2444 10848 2450 10900
rect 2270 10812 2450 10848
rect 2270 10778 2276 10812
rect 2310 10778 2410 10812
rect 2444 10778 2450 10812
rect 2270 10740 2450 10778
rect 2270 10706 2276 10740
rect 2310 10706 2410 10740
rect 2444 10706 2450 10740
rect 2270 10668 2450 10706
rect 2270 10634 2276 10668
rect 2310 10634 2410 10668
rect 2444 10634 2450 10668
rect 2270 10596 2450 10634
rect 2270 10562 2276 10596
rect 2310 10562 2410 10596
rect 2444 10562 2450 10596
rect 2270 10524 2450 10562
rect 2270 10490 2276 10524
rect 2310 10490 2410 10524
rect 2444 10490 2450 10524
rect 2270 10452 2450 10490
rect 2270 10418 2276 10452
rect 2310 10418 2410 10452
rect 2444 10418 2450 10452
rect 2270 10380 2450 10418
rect 2270 10346 2276 10380
rect 2310 10346 2410 10380
rect 2444 10346 2450 10380
rect 2270 10308 2450 10346
rect 2270 10274 2276 10308
rect 2310 10274 2410 10308
rect 2444 10274 2450 10308
rect 2270 10236 2450 10274
rect 2270 10202 2276 10236
rect 2310 10202 2410 10236
rect 2444 10202 2450 10236
rect 2270 10164 2450 10202
rect 2270 10130 2276 10164
rect 2310 10130 2410 10164
rect 2444 10130 2450 10164
rect 2270 10092 2450 10130
rect 2270 10058 2276 10092
rect 2310 10058 2410 10092
rect 2444 10058 2450 10092
rect 2270 10020 2450 10058
rect 2270 9986 2276 10020
rect 2310 9986 2410 10020
rect 2444 9986 2450 10020
rect 2580 15586 7729 15660
rect 2580 15552 3035 15586
rect 3069 15552 3108 15586
rect 3142 15552 3181 15586
rect 3215 15552 3254 15586
rect 3288 15552 3327 15586
rect 3361 15552 3400 15586
rect 3434 15552 3473 15586
rect 3507 15552 3546 15586
rect 3580 15552 3619 15586
rect 3653 15552 3692 15586
rect 3726 15552 3765 15586
rect 3799 15552 3838 15586
rect 3872 15552 3911 15586
rect 3945 15552 3984 15586
rect 4018 15552 4057 15586
rect 4091 15552 4130 15586
rect 4164 15552 4203 15586
rect 4237 15552 4276 15586
rect 4310 15552 4349 15586
rect 4383 15552 4422 15586
rect 4456 15552 4495 15586
rect 4529 15552 4568 15586
rect 4602 15552 4641 15586
rect 4675 15552 4714 15586
rect 4748 15552 4787 15586
rect 4821 15552 4860 15586
rect 4894 15552 4933 15586
rect 4967 15552 5006 15586
rect 5040 15552 5079 15586
rect 5113 15552 5152 15586
rect 5186 15552 5225 15586
rect 5259 15552 5298 15586
rect 5332 15552 5371 15586
rect 5405 15552 5444 15586
rect 5478 15552 5517 15586
rect 5551 15552 5590 15586
rect 5624 15552 5663 15586
rect 5697 15552 5736 15586
rect 5770 15552 5809 15586
rect 5843 15552 5881 15586
rect 5915 15552 5953 15586
rect 5987 15552 6025 15586
rect 6059 15552 6097 15586
rect 6131 15552 6169 15586
rect 6203 15552 6241 15586
rect 6275 15552 6313 15586
rect 6347 15552 6385 15586
rect 6419 15552 6457 15586
rect 6491 15552 6529 15586
rect 6563 15552 6601 15586
rect 6635 15552 6673 15586
rect 6707 15552 6745 15586
rect 6779 15552 6817 15586
rect 6851 15552 6889 15586
rect 6923 15552 6961 15586
rect 6995 15552 7033 15586
rect 7067 15552 7105 15586
rect 7139 15552 7177 15586
rect 7211 15552 7249 15586
rect 7283 15552 7321 15586
rect 7355 15552 7393 15586
rect 7427 15552 7465 15586
rect 7499 15552 7537 15586
rect 7571 15552 7609 15586
rect 7643 15552 7681 15586
rect 7715 15552 7729 15586
rect 2580 15546 7729 15552
rect 8044 15645 8050 15679
rect 8084 15669 8224 15679
rect 8084 15645 8184 15669
rect 8044 15635 8184 15645
rect 8218 15635 8224 15669
rect 8044 15607 8224 15635
rect 8044 15573 8050 15607
rect 8084 15597 8224 15607
rect 8084 15573 8184 15597
rect 8044 15563 8184 15573
rect 8218 15563 8224 15597
rect 2580 15535 2761 15546
tri 2761 15535 2772 15546 nw
rect 8044 15535 8224 15563
rect 2580 15501 2727 15535
tri 2727 15501 2761 15535 nw
rect 8044 15501 8050 15535
rect 8084 15525 8224 15535
rect 8084 15501 8184 15525
rect 2580 15491 2717 15501
tri 2717 15491 2727 15501 nw
rect 8044 15491 8184 15501
rect 8218 15491 8224 15525
rect 2580 13917 2712 15491
tri 2712 15486 2717 15491 nw
rect 8044 15463 8224 15491
rect 2824 15452 2942 15458
rect 2876 15400 2890 15452
rect 2824 15383 2942 15400
rect 2876 15331 2890 15383
rect 2824 15314 2942 15331
rect 2876 15262 2890 15314
rect 2824 15245 2942 15262
rect 2876 15193 2890 15245
rect 2824 15176 2942 15193
rect 2876 15154 2890 15176
rect 2824 15107 2830 15124
rect 2936 15107 2942 15124
rect 2824 15038 2830 15055
rect 2936 15038 2942 15055
rect 2824 14968 2830 14986
rect 2936 14968 2942 14986
rect 2824 14898 2830 14916
rect 2936 14898 2942 14916
rect 2824 14112 2830 14846
rect 2936 14112 2942 14846
rect 2824 14100 2942 14112
rect 3101 15446 3219 15458
rect 3101 15412 3107 15446
rect 3141 15412 3179 15446
rect 3213 15412 3219 15446
rect 3101 15373 3219 15412
rect 3101 15339 3107 15373
rect 3141 15339 3179 15373
rect 3213 15339 3219 15373
rect 3101 15300 3219 15339
rect 3101 15266 3107 15300
rect 3141 15266 3179 15300
rect 3213 15266 3219 15300
rect 3101 15227 3219 15266
rect 3101 15193 3107 15227
rect 3141 15193 3179 15227
rect 3213 15193 3219 15227
rect 3101 15154 3219 15193
rect 3101 14714 3107 15154
rect 3213 14714 3219 15154
rect 3101 14645 3107 14662
rect 3213 14645 3219 14662
rect 3101 14576 3107 14593
rect 3213 14576 3219 14593
rect 3101 14507 3107 14524
rect 3213 14507 3219 14524
rect 3101 14438 3107 14455
rect 3213 14438 3219 14455
rect 3101 14368 3107 14386
rect 3213 14368 3219 14386
rect 3101 14298 3107 14316
rect 3213 14298 3219 14316
rect 3101 14228 3107 14246
rect 3213 14228 3219 14246
rect 3101 14158 3107 14176
rect 3213 14158 3219 14176
rect 3153 14106 3167 14112
rect 3101 14100 3219 14106
rect 3378 15452 3496 15458
rect 3430 15400 3444 15452
rect 3378 15383 3496 15400
rect 3430 15331 3444 15383
rect 3378 15314 3496 15331
rect 3430 15262 3444 15314
rect 3378 15245 3496 15262
rect 3430 15193 3444 15245
rect 3378 15176 3496 15193
rect 3430 15154 3444 15176
rect 3378 15107 3384 15124
rect 3490 15107 3496 15124
rect 3378 15038 3384 15055
rect 3490 15038 3496 15055
rect 3378 14968 3384 14986
rect 3490 14968 3496 14986
rect 3378 14898 3384 14916
rect 3490 14898 3496 14916
rect 3378 14112 3384 14846
rect 3490 14112 3496 14846
rect 3378 14100 3496 14112
rect 3655 15446 3773 15458
rect 3655 15412 3661 15446
rect 3695 15412 3733 15446
rect 3767 15412 3773 15446
rect 3655 15373 3773 15412
rect 3655 15339 3661 15373
rect 3695 15339 3733 15373
rect 3767 15339 3773 15373
rect 3655 15300 3773 15339
rect 3655 15266 3661 15300
rect 3695 15266 3733 15300
rect 3767 15266 3773 15300
rect 3655 15227 3773 15266
rect 3655 15193 3661 15227
rect 3695 15193 3733 15227
rect 3767 15193 3773 15227
rect 3655 15154 3773 15193
rect 3655 14714 3661 15154
rect 3767 14714 3773 15154
rect 3655 14645 3661 14662
rect 3767 14645 3773 14662
rect 3655 14576 3661 14593
rect 3767 14576 3773 14593
rect 3655 14507 3661 14524
rect 3767 14507 3773 14524
rect 3655 14438 3661 14455
rect 3767 14438 3773 14455
rect 3655 14368 3661 14386
rect 3767 14368 3773 14386
rect 3655 14298 3661 14316
rect 3767 14298 3773 14316
rect 3655 14228 3661 14246
rect 3767 14228 3773 14246
rect 3655 14158 3661 14176
rect 3767 14158 3773 14176
rect 3707 14106 3721 14112
rect 3655 14100 3773 14106
rect 3932 15452 4050 15458
rect 3984 15400 3998 15452
rect 3932 15383 4050 15400
rect 3984 15331 3998 15383
rect 3932 15314 4050 15331
rect 3984 15262 3998 15314
rect 3932 15245 4050 15262
rect 3984 15193 3998 15245
rect 3932 15176 4050 15193
rect 3984 15154 3998 15176
rect 3932 15107 3938 15124
rect 4044 15107 4050 15124
rect 3932 15038 3938 15055
rect 4044 15038 4050 15055
rect 3932 14968 3938 14986
rect 4044 14968 4050 14986
rect 3932 14898 3938 14916
rect 4044 14898 4050 14916
rect 3932 14112 3938 14846
rect 4044 14112 4050 14846
rect 3932 14100 4050 14112
rect 4209 15446 4327 15458
rect 4209 15412 4215 15446
rect 4249 15412 4287 15446
rect 4321 15412 4327 15446
rect 4209 15373 4327 15412
rect 4209 15339 4215 15373
rect 4249 15339 4287 15373
rect 4321 15339 4327 15373
rect 4209 15300 4327 15339
rect 4209 15266 4215 15300
rect 4249 15266 4287 15300
rect 4321 15266 4327 15300
rect 4209 15227 4327 15266
rect 4209 15193 4215 15227
rect 4249 15193 4287 15227
rect 4321 15193 4327 15227
rect 4209 15154 4327 15193
rect 4209 14714 4215 15154
rect 4321 14714 4327 15154
rect 4209 14645 4215 14662
rect 4321 14645 4327 14662
rect 4209 14576 4215 14593
rect 4321 14576 4327 14593
rect 4209 14507 4215 14524
rect 4321 14507 4327 14524
rect 4209 14438 4215 14455
rect 4321 14438 4327 14455
rect 4209 14368 4215 14386
rect 4321 14368 4327 14386
rect 4209 14298 4215 14316
rect 4321 14298 4327 14316
rect 4209 14228 4215 14246
rect 4321 14228 4327 14246
rect 4209 14158 4215 14176
rect 4321 14158 4327 14176
rect 4261 14106 4275 14112
rect 4209 14100 4327 14106
rect 4486 15452 4604 15458
rect 4538 15400 4552 15452
rect 4486 15383 4604 15400
rect 4538 15331 4552 15383
rect 4486 15314 4604 15331
rect 4538 15262 4552 15314
rect 4486 15245 4604 15262
rect 4538 15193 4552 15245
rect 4486 15176 4604 15193
rect 4538 15154 4552 15176
rect 4486 15107 4492 15124
rect 4598 15107 4604 15124
rect 4486 15038 4492 15055
rect 4598 15038 4604 15055
rect 4486 14968 4492 14986
rect 4598 14968 4604 14986
rect 4486 14898 4492 14916
rect 4598 14898 4604 14916
rect 4486 14112 4492 14846
rect 4598 14112 4604 14846
rect 4486 14100 4604 14112
rect 4763 15446 4881 15458
rect 4763 15412 4769 15446
rect 4803 15412 4841 15446
rect 4875 15412 4881 15446
rect 4763 15373 4881 15412
rect 4763 15339 4769 15373
rect 4803 15339 4841 15373
rect 4875 15339 4881 15373
rect 4763 15300 4881 15339
rect 4763 15266 4769 15300
rect 4803 15266 4841 15300
rect 4875 15266 4881 15300
rect 4763 15227 4881 15266
rect 4763 15193 4769 15227
rect 4803 15193 4841 15227
rect 4875 15193 4881 15227
rect 4763 15154 4881 15193
rect 4763 14714 4769 15154
rect 4875 14714 4881 15154
rect 4763 14645 4769 14662
rect 4875 14645 4881 14662
rect 4763 14576 4769 14593
rect 4875 14576 4881 14593
rect 4763 14507 4769 14524
rect 4875 14507 4881 14524
rect 4763 14438 4769 14455
rect 4875 14438 4881 14455
rect 4763 14368 4769 14386
rect 4875 14368 4881 14386
rect 4763 14298 4769 14316
rect 4875 14298 4881 14316
rect 4763 14228 4769 14246
rect 4875 14228 4881 14246
rect 4763 14158 4769 14176
rect 4875 14158 4881 14176
rect 4815 14106 4829 14112
rect 4763 14100 4881 14106
rect 5040 15452 5158 15458
rect 5092 15400 5106 15452
rect 5040 15383 5158 15400
rect 5092 15331 5106 15383
rect 5040 15314 5158 15331
rect 5092 15262 5106 15314
rect 5040 15245 5158 15262
rect 5092 15193 5106 15245
rect 5040 15176 5158 15193
rect 5092 15154 5106 15176
rect 5040 15107 5046 15124
rect 5152 15107 5158 15124
rect 5040 15038 5046 15055
rect 5152 15038 5158 15055
rect 5040 14968 5046 14986
rect 5152 14968 5158 14986
rect 5040 14898 5046 14916
rect 5152 14898 5158 14916
rect 5040 14112 5046 14846
rect 5152 14112 5158 14846
rect 5040 14100 5158 14112
rect 5317 15446 5435 15458
rect 5317 15412 5323 15446
rect 5357 15412 5395 15446
rect 5429 15412 5435 15446
rect 5317 15373 5435 15412
rect 5317 15339 5323 15373
rect 5357 15339 5395 15373
rect 5429 15339 5435 15373
rect 5317 15300 5435 15339
rect 5317 15266 5323 15300
rect 5357 15266 5395 15300
rect 5429 15266 5435 15300
rect 5317 15227 5435 15266
rect 5317 15193 5323 15227
rect 5357 15193 5395 15227
rect 5429 15193 5435 15227
rect 5317 15154 5435 15193
rect 5317 14714 5323 15154
rect 5429 14714 5435 15154
rect 5317 14645 5323 14662
rect 5429 14645 5435 14662
rect 5317 14576 5323 14593
rect 5429 14576 5435 14593
rect 5317 14507 5323 14524
rect 5429 14507 5435 14524
rect 5317 14438 5323 14455
rect 5429 14438 5435 14455
rect 5317 14368 5323 14386
rect 5429 14368 5435 14386
rect 5317 14298 5323 14316
rect 5429 14298 5435 14316
rect 5317 14228 5323 14246
rect 5429 14228 5435 14246
rect 5317 14158 5323 14176
rect 5429 14158 5435 14176
rect 5369 14106 5383 14112
rect 5317 14100 5435 14106
rect 5594 15452 5712 15458
rect 5646 15400 5660 15452
rect 5594 15383 5712 15400
rect 5646 15331 5660 15383
rect 5594 15314 5712 15331
rect 5646 15262 5660 15314
rect 5594 15245 5712 15262
rect 5646 15193 5660 15245
rect 5594 15176 5712 15193
rect 5646 15154 5660 15176
rect 5594 15107 5600 15124
rect 5706 15107 5712 15124
rect 5594 15038 5600 15055
rect 5706 15038 5712 15055
rect 5594 14968 5600 14986
rect 5706 14968 5712 14986
rect 5594 14898 5600 14916
rect 5706 14898 5712 14916
rect 5594 14112 5600 14846
rect 5706 14112 5712 14846
rect 5594 14100 5712 14112
rect 5871 15446 5989 15458
rect 5871 15412 5877 15446
rect 5911 15412 5949 15446
rect 5983 15412 5989 15446
rect 5871 15373 5989 15412
rect 5871 15339 5877 15373
rect 5911 15339 5949 15373
rect 5983 15339 5989 15373
rect 5871 15300 5989 15339
rect 5871 15266 5877 15300
rect 5911 15266 5949 15300
rect 5983 15266 5989 15300
rect 5871 15227 5989 15266
rect 5871 15193 5877 15227
rect 5911 15193 5949 15227
rect 5983 15193 5989 15227
rect 5871 15154 5989 15193
rect 5871 14714 5877 15154
rect 5983 14714 5989 15154
rect 5871 14645 5877 14662
rect 5983 14645 5989 14662
rect 5871 14576 5877 14593
rect 5983 14576 5989 14593
rect 5871 14507 5877 14524
rect 5983 14507 5989 14524
rect 5871 14438 5877 14455
rect 5983 14438 5989 14455
rect 5871 14368 5877 14386
rect 5983 14368 5989 14386
rect 5871 14298 5877 14316
rect 5983 14298 5989 14316
rect 5871 14228 5877 14246
rect 5983 14228 5989 14246
rect 5871 14158 5877 14176
rect 5983 14158 5989 14176
rect 5923 14106 5937 14112
rect 5871 14100 5989 14106
rect 6148 15452 6266 15458
rect 6200 15400 6214 15452
rect 6148 15383 6266 15400
rect 6200 15331 6214 15383
rect 6148 15314 6266 15331
rect 6200 15262 6214 15314
rect 6148 15245 6266 15262
rect 6200 15193 6214 15245
rect 6148 15176 6266 15193
rect 6200 15154 6214 15176
rect 6148 15107 6154 15124
rect 6260 15107 6266 15124
rect 6148 15038 6154 15055
rect 6260 15038 6266 15055
rect 6148 14968 6154 14986
rect 6260 14968 6266 14986
rect 6148 14898 6154 14916
rect 6260 14898 6266 14916
rect 6148 14112 6154 14846
rect 6260 14112 6266 14846
rect 6148 14100 6266 14112
rect 6425 15446 6543 15458
rect 6425 15412 6431 15446
rect 6465 15412 6503 15446
rect 6537 15412 6543 15446
rect 6425 15373 6543 15412
rect 6425 15339 6431 15373
rect 6465 15339 6503 15373
rect 6537 15339 6543 15373
rect 6425 15300 6543 15339
rect 6425 15266 6431 15300
rect 6465 15266 6503 15300
rect 6537 15266 6543 15300
rect 6425 15227 6543 15266
rect 6425 15193 6431 15227
rect 6465 15193 6503 15227
rect 6537 15193 6543 15227
rect 6425 15154 6543 15193
rect 6425 14714 6431 15154
rect 6537 14714 6543 15154
rect 6425 14645 6431 14662
rect 6537 14645 6543 14662
rect 6425 14576 6431 14593
rect 6537 14576 6543 14593
rect 6425 14507 6431 14524
rect 6537 14507 6543 14524
rect 6425 14438 6431 14455
rect 6537 14438 6543 14455
rect 6425 14368 6431 14386
rect 6537 14368 6543 14386
rect 6425 14298 6431 14316
rect 6537 14298 6543 14316
rect 6425 14228 6431 14246
rect 6537 14228 6543 14246
rect 6425 14158 6431 14176
rect 6537 14158 6543 14176
rect 6477 14106 6491 14112
rect 6425 14100 6543 14106
rect 6702 15452 6820 15458
rect 6754 15400 6768 15452
rect 6702 15383 6820 15400
rect 6754 15331 6768 15383
rect 6702 15314 6820 15331
rect 6754 15262 6768 15314
rect 6702 15245 6820 15262
rect 6754 15193 6768 15245
rect 6702 15176 6820 15193
rect 6754 15154 6768 15176
rect 6702 15107 6708 15124
rect 6814 15107 6820 15124
rect 6702 15038 6708 15055
rect 6814 15038 6820 15055
rect 6702 14968 6708 14986
rect 6814 14968 6820 14986
rect 6702 14898 6708 14916
rect 6814 14898 6820 14916
rect 6702 14112 6708 14846
rect 6814 14112 6820 14846
rect 6702 14100 6820 14112
rect 6979 15446 7097 15458
rect 6979 15412 6985 15446
rect 7019 15412 7057 15446
rect 7091 15412 7097 15446
rect 6979 15373 7097 15412
rect 6979 15339 6985 15373
rect 7019 15339 7057 15373
rect 7091 15339 7097 15373
rect 6979 15300 7097 15339
rect 6979 15266 6985 15300
rect 7019 15266 7057 15300
rect 7091 15266 7097 15300
rect 6979 15227 7097 15266
rect 6979 15193 6985 15227
rect 7019 15193 7057 15227
rect 7091 15193 7097 15227
rect 6979 15154 7097 15193
rect 6979 14714 6985 15154
rect 7091 14714 7097 15154
rect 6979 14645 6985 14662
rect 7091 14645 7097 14662
rect 6979 14576 6985 14593
rect 7091 14576 7097 14593
rect 6979 14507 6985 14524
rect 7091 14507 7097 14524
rect 6979 14438 6985 14455
rect 7091 14438 7097 14455
rect 6979 14368 6985 14386
rect 7091 14368 7097 14386
rect 6979 14298 6985 14316
rect 7091 14298 7097 14316
rect 6979 14228 6985 14246
rect 7091 14228 7097 14246
rect 6979 14158 6985 14176
rect 7091 14158 7097 14176
rect 7031 14106 7045 14112
rect 6979 14100 7097 14106
rect 7256 15452 7374 15458
rect 7308 15400 7322 15452
rect 7256 15383 7374 15400
rect 7308 15331 7322 15383
rect 7256 15314 7374 15331
rect 7308 15262 7322 15314
rect 7256 15245 7374 15262
rect 7308 15193 7322 15245
rect 7256 15176 7374 15193
rect 7308 15154 7322 15176
rect 7256 15107 7262 15124
rect 7368 15107 7374 15124
rect 7256 15038 7262 15055
rect 7368 15038 7374 15055
rect 7256 14968 7262 14986
rect 7368 14968 7374 14986
rect 7256 14898 7262 14916
rect 7368 14898 7374 14916
rect 7256 14112 7262 14846
rect 7368 14112 7374 14846
rect 7256 14100 7374 14112
rect 7533 15446 7651 15458
rect 7533 15412 7539 15446
rect 7573 15412 7611 15446
rect 7645 15412 7651 15446
rect 7533 15373 7651 15412
rect 7533 15339 7539 15373
rect 7573 15339 7611 15373
rect 7645 15339 7651 15373
rect 7533 15300 7651 15339
rect 7533 15266 7539 15300
rect 7573 15266 7611 15300
rect 7645 15266 7651 15300
rect 7533 15227 7651 15266
rect 7533 15193 7539 15227
rect 7573 15193 7611 15227
rect 7645 15193 7651 15227
rect 7533 15154 7651 15193
rect 7533 14714 7539 15154
rect 7645 14714 7651 15154
rect 7533 14645 7539 14662
rect 7645 14645 7651 14662
rect 7533 14576 7539 14593
rect 7645 14576 7651 14593
rect 7533 14507 7539 14524
rect 7645 14507 7651 14524
rect 7533 14438 7539 14455
rect 7645 14438 7651 14455
rect 7533 14368 7539 14386
rect 7645 14368 7651 14386
rect 7533 14298 7539 14316
rect 7645 14298 7651 14316
rect 7533 14228 7539 14246
rect 7645 14228 7651 14246
rect 7533 14158 7539 14176
rect 7645 14158 7651 14176
rect 7585 14106 7599 14112
rect 7533 14100 7651 14106
rect 7810 15452 7928 15458
rect 7862 15400 7876 15452
rect 7810 15383 7928 15400
rect 7862 15331 7876 15383
rect 7810 15314 7928 15331
rect 7862 15262 7876 15314
rect 7810 15245 7928 15262
rect 7862 15193 7876 15245
rect 7810 15176 7928 15193
rect 7862 15154 7876 15176
rect 7810 15107 7816 15124
rect 7922 15107 7928 15124
rect 7810 15038 7816 15055
rect 7922 15038 7928 15055
rect 7810 14968 7816 14986
rect 7922 14968 7928 14986
rect 7810 14898 7816 14916
rect 7922 14898 7928 14916
rect 7810 14112 7816 14846
rect 7922 14112 7928 14846
rect 7810 14100 7928 14112
rect 8044 15456 8050 15463
rect 8084 15456 8224 15463
rect 8044 15404 8047 15456
rect 8099 15404 8169 15456
rect 8221 15404 8224 15456
rect 8044 15391 8224 15404
rect 8044 15387 8050 15391
rect 8084 15387 8224 15391
rect 8044 15335 8047 15387
rect 8099 15335 8169 15387
rect 8221 15335 8224 15387
rect 8044 15319 8224 15335
rect 8044 15318 8050 15319
rect 8084 15318 8224 15319
rect 8044 15266 8047 15318
rect 8099 15266 8169 15318
rect 8221 15266 8224 15318
rect 8044 15249 8224 15266
rect 8044 15197 8047 15249
rect 8099 15197 8169 15249
rect 8221 15197 8224 15249
rect 8044 15180 8224 15197
rect 8044 15128 8047 15180
rect 8099 15128 8169 15180
rect 8221 15128 8224 15180
rect 8044 15110 8224 15128
rect 8044 15058 8047 15110
rect 8099 15058 8169 15110
rect 8221 15058 8224 15110
rect 8044 15040 8224 15058
rect 8044 14988 8047 15040
rect 8099 14988 8169 15040
rect 8221 14988 8224 15040
rect 8044 14987 8184 14988
rect 8218 14987 8224 14988
rect 8044 14970 8224 14987
rect 8044 14918 8047 14970
rect 8099 14918 8169 14970
rect 8221 14918 8224 14970
rect 8044 14915 8184 14918
rect 8218 14915 8224 14918
rect 8044 14900 8224 14915
rect 8044 14848 8047 14900
rect 8099 14848 8169 14900
rect 8221 14848 8224 14900
rect 8044 14843 8184 14848
rect 8218 14843 8224 14848
rect 8044 14815 8224 14843
rect 8044 14781 8050 14815
rect 8084 14805 8224 14815
rect 8084 14781 8184 14805
rect 8044 14771 8184 14781
rect 8218 14771 8224 14805
rect 8044 14743 8224 14771
rect 8044 14709 8050 14743
rect 8084 14733 8224 14743
rect 8084 14709 8184 14733
rect 8044 14699 8184 14709
rect 8218 14699 8224 14733
rect 8044 14671 8224 14699
rect 8044 14637 8050 14671
rect 8084 14661 8224 14671
rect 8084 14637 8184 14661
rect 8044 14627 8184 14637
rect 8218 14627 8224 14661
rect 8044 14599 8224 14627
rect 8044 14565 8050 14599
rect 8084 14589 8224 14599
rect 8084 14565 8184 14589
rect 8044 14555 8184 14565
rect 8218 14555 8224 14589
rect 8044 14527 8224 14555
rect 8044 14493 8050 14527
rect 8084 14517 8224 14527
rect 8084 14493 8184 14517
rect 8044 14483 8184 14493
rect 8218 14483 8224 14517
rect 8044 14455 8224 14483
rect 8044 14421 8050 14455
rect 8084 14445 8224 14455
rect 8084 14421 8184 14445
rect 8044 14411 8184 14421
rect 8218 14411 8224 14445
rect 8044 14383 8224 14411
rect 8044 14349 8050 14383
rect 8084 14373 8224 14383
rect 8084 14349 8184 14373
rect 8044 14339 8184 14349
rect 8218 14339 8224 14373
rect 8044 14311 8224 14339
rect 8044 14277 8050 14311
rect 8084 14301 8224 14311
rect 8084 14277 8184 14301
rect 8044 14267 8184 14277
rect 8218 14267 8224 14301
rect 8044 14239 8224 14267
rect 8044 14205 8050 14239
rect 8084 14229 8224 14239
rect 8084 14205 8184 14229
rect 8044 14195 8184 14205
rect 8218 14195 8224 14229
rect 8044 14167 8224 14195
rect 8044 14133 8050 14167
rect 8084 14157 8224 14167
rect 8084 14133 8184 14157
rect 8044 14123 8184 14133
rect 8218 14123 8224 14157
rect 8044 14095 8224 14123
rect 8044 14061 8050 14095
rect 8084 14085 8224 14095
rect 8084 14061 8184 14085
rect 8044 14051 8184 14061
rect 8218 14051 8224 14085
rect 8044 14023 8224 14051
rect 8044 13989 8050 14023
rect 8084 14013 8224 14023
rect 8084 13989 8184 14013
rect 8044 13979 8184 13989
rect 8218 13979 8224 14013
rect 8044 13951 8224 13979
tri 2712 13917 2741 13946 sw
rect 8044 13917 8050 13951
rect 8084 13941 8224 13951
rect 8084 13917 8184 13941
rect 2580 13914 2741 13917
tri 2741 13914 2744 13917 sw
rect 2580 13856 7748 13914
rect 2580 13822 3035 13856
rect 3069 13822 3108 13856
rect 3142 13822 3181 13856
rect 3215 13822 3254 13856
rect 3288 13822 3327 13856
rect 3361 13822 3400 13856
rect 3434 13822 3473 13856
rect 3507 13822 3546 13856
rect 3580 13822 3619 13856
rect 3653 13822 3692 13856
rect 3726 13822 3765 13856
rect 3799 13822 3838 13856
rect 3872 13822 3911 13856
rect 3945 13822 3984 13856
rect 4018 13822 4057 13856
rect 4091 13822 4130 13856
rect 4164 13822 4203 13856
rect 4237 13822 4276 13856
rect 4310 13822 4349 13856
rect 4383 13822 4422 13856
rect 4456 13822 4495 13856
rect 4529 13822 4568 13856
rect 4602 13822 4641 13856
rect 4675 13822 4714 13856
rect 4748 13822 4787 13856
rect 4821 13822 4860 13856
rect 4894 13822 4933 13856
rect 4967 13822 5006 13856
rect 5040 13822 5079 13856
rect 5113 13822 5152 13856
rect 5186 13822 5225 13856
rect 5259 13822 5298 13856
rect 5332 13822 5371 13856
rect 5405 13822 5444 13856
rect 5478 13822 5517 13856
rect 5551 13822 5590 13856
rect 5624 13822 5663 13856
rect 5697 13822 5736 13856
rect 5770 13822 5809 13856
rect 5843 13822 5881 13856
rect 5915 13822 5953 13856
rect 5987 13822 6025 13856
rect 6059 13822 6097 13856
rect 6131 13822 6169 13856
rect 6203 13822 6241 13856
rect 6275 13822 6313 13856
rect 6347 13822 6385 13856
rect 6419 13822 6457 13856
rect 6491 13822 6529 13856
rect 6563 13822 6601 13856
rect 6635 13822 6673 13856
rect 6707 13822 6745 13856
rect 6779 13822 6817 13856
rect 6851 13822 6889 13856
rect 6923 13822 6961 13856
rect 6995 13822 7033 13856
rect 7067 13822 7105 13856
rect 7139 13822 7177 13856
rect 7211 13822 7249 13856
rect 7283 13822 7321 13856
rect 7355 13822 7393 13856
rect 7427 13822 7465 13856
rect 7499 13822 7537 13856
rect 7571 13822 7609 13856
rect 7643 13822 7681 13856
rect 7715 13822 7748 13856
rect 2580 13751 7748 13822
rect 8044 13907 8184 13917
rect 8218 13907 8224 13941
rect 8044 13879 8224 13907
rect 8044 13845 8050 13879
rect 8084 13869 8224 13879
rect 8084 13845 8184 13869
rect 8044 13835 8184 13845
rect 8218 13835 8224 13869
rect 8044 13807 8224 13835
rect 8044 13773 8050 13807
rect 8084 13797 8224 13807
rect 8084 13773 8184 13797
rect 8044 13763 8184 13773
rect 8218 13763 8224 13797
rect 2580 13735 2740 13751
tri 2740 13735 2756 13751 nw
rect 8044 13735 8224 13763
rect 2580 11959 2712 13735
tri 2712 13707 2740 13735 nw
rect 8044 13701 8050 13735
rect 8084 13725 8224 13735
rect 8084 13701 8184 13725
rect 8044 13691 8184 13701
rect 8218 13691 8224 13725
rect 8044 13663 8224 13691
rect 8044 13629 8050 13663
rect 8084 13653 8224 13663
rect 8084 13629 8184 13653
rect 8044 13619 8184 13629
rect 8218 13619 8224 13653
rect 8044 13591 8224 13619
rect 8044 13557 8050 13591
rect 8084 13581 8224 13591
rect 8084 13557 8184 13581
rect 8044 13547 8184 13557
rect 8218 13547 8224 13581
rect 8044 13519 8224 13547
rect 8044 13485 8050 13519
rect 8084 13509 8224 13519
rect 8084 13485 8184 13509
rect 8044 13475 8184 13485
rect 8218 13475 8224 13509
rect 2824 13452 2942 13458
rect 2876 13400 2890 13452
rect 2824 13383 2942 13400
rect 2876 13331 2890 13383
rect 2824 13314 2942 13331
rect 2876 13262 2890 13314
rect 2824 13245 2942 13262
rect 2876 13193 2890 13245
rect 2824 13176 2942 13193
rect 2876 13154 2890 13176
rect 2824 13107 2830 13124
rect 2936 13107 2942 13124
rect 2824 13038 2830 13055
rect 2936 13038 2942 13055
rect 2824 12968 2830 12986
rect 2936 12968 2942 12986
rect 2824 12898 2830 12916
rect 2936 12898 2942 12916
rect 2824 12112 2830 12846
rect 2936 12112 2942 12846
rect 2824 12100 2942 12112
rect 3101 13446 3219 13458
rect 3101 13412 3107 13446
rect 3141 13412 3179 13446
rect 3213 13412 3219 13446
rect 3101 13373 3219 13412
rect 3101 13339 3107 13373
rect 3141 13339 3179 13373
rect 3213 13339 3219 13373
rect 3101 13300 3219 13339
rect 3101 13266 3107 13300
rect 3141 13266 3179 13300
rect 3213 13266 3219 13300
rect 3101 13227 3219 13266
rect 3101 13193 3107 13227
rect 3141 13193 3179 13227
rect 3213 13193 3219 13227
rect 3101 13154 3219 13193
rect 3101 12714 3107 13154
rect 3213 12714 3219 13154
rect 3101 12645 3107 12662
rect 3213 12645 3219 12662
rect 3101 12576 3107 12593
rect 3213 12576 3219 12593
rect 3101 12507 3107 12524
rect 3213 12507 3219 12524
rect 3101 12438 3107 12455
rect 3213 12438 3219 12455
rect 3101 12368 3107 12386
rect 3213 12368 3219 12386
rect 3101 12298 3107 12316
rect 3213 12298 3219 12316
rect 3101 12228 3107 12246
rect 3213 12228 3219 12246
rect 3101 12158 3107 12176
rect 3213 12158 3219 12176
rect 3153 12106 3167 12112
rect 3101 12100 3219 12106
rect 3378 13452 3496 13458
rect 3430 13400 3444 13452
rect 3378 13383 3496 13400
rect 3430 13331 3444 13383
rect 3378 13314 3496 13331
rect 3430 13262 3444 13314
rect 3378 13245 3496 13262
rect 3430 13193 3444 13245
rect 3378 13176 3496 13193
rect 3430 13154 3444 13176
rect 3378 13107 3384 13124
rect 3490 13107 3496 13124
rect 3378 13038 3384 13055
rect 3490 13038 3496 13055
rect 3378 12968 3384 12986
rect 3490 12968 3496 12986
rect 3378 12898 3384 12916
rect 3490 12898 3496 12916
rect 3378 12112 3384 12846
rect 3490 12112 3496 12846
rect 3378 12100 3496 12112
rect 3655 13446 3773 13458
rect 3655 13412 3661 13446
rect 3695 13412 3733 13446
rect 3767 13412 3773 13446
rect 3655 13373 3773 13412
rect 3655 13339 3661 13373
rect 3695 13339 3733 13373
rect 3767 13339 3773 13373
rect 3655 13300 3773 13339
rect 3655 13266 3661 13300
rect 3695 13266 3733 13300
rect 3767 13266 3773 13300
rect 3655 13227 3773 13266
rect 3655 13193 3661 13227
rect 3695 13193 3733 13227
rect 3767 13193 3773 13227
rect 3655 13154 3773 13193
rect 3655 12714 3661 13154
rect 3767 12714 3773 13154
rect 3655 12645 3661 12662
rect 3767 12645 3773 12662
rect 3655 12576 3661 12593
rect 3767 12576 3773 12593
rect 3655 12507 3661 12524
rect 3767 12507 3773 12524
rect 3655 12438 3661 12455
rect 3767 12438 3773 12455
rect 3655 12368 3661 12386
rect 3767 12368 3773 12386
rect 3655 12298 3661 12316
rect 3767 12298 3773 12316
rect 3655 12228 3661 12246
rect 3767 12228 3773 12246
rect 3655 12158 3661 12176
rect 3767 12158 3773 12176
rect 3707 12106 3721 12112
rect 3655 12100 3773 12106
rect 3932 13452 4050 13458
rect 3984 13400 3998 13452
rect 3932 13383 4050 13400
rect 3984 13331 3998 13383
rect 3932 13314 4050 13331
rect 3984 13262 3998 13314
rect 3932 13245 4050 13262
rect 3984 13193 3998 13245
rect 3932 13176 4050 13193
rect 3984 13154 3998 13176
rect 3932 13107 3938 13124
rect 4044 13107 4050 13124
rect 3932 13038 3938 13055
rect 4044 13038 4050 13055
rect 3932 12968 3938 12986
rect 4044 12968 4050 12986
rect 3932 12898 3938 12916
rect 4044 12898 4050 12916
rect 3932 12112 3938 12846
rect 4044 12112 4050 12846
rect 3932 12100 4050 12112
rect 4209 13446 4327 13458
rect 4209 13412 4215 13446
rect 4249 13412 4287 13446
rect 4321 13412 4327 13446
rect 4209 13373 4327 13412
rect 4209 13339 4215 13373
rect 4249 13339 4287 13373
rect 4321 13339 4327 13373
rect 4209 13300 4327 13339
rect 4209 13266 4215 13300
rect 4249 13266 4287 13300
rect 4321 13266 4327 13300
rect 4209 13227 4327 13266
rect 4209 13193 4215 13227
rect 4249 13193 4287 13227
rect 4321 13193 4327 13227
rect 4209 13154 4327 13193
rect 4209 12714 4215 13154
rect 4321 12714 4327 13154
rect 4209 12645 4215 12662
rect 4321 12645 4327 12662
rect 4209 12576 4215 12593
rect 4321 12576 4327 12593
rect 4209 12507 4215 12524
rect 4321 12507 4327 12524
rect 4209 12438 4215 12455
rect 4321 12438 4327 12455
rect 4209 12368 4215 12386
rect 4321 12368 4327 12386
rect 4209 12298 4215 12316
rect 4321 12298 4327 12316
rect 4209 12228 4215 12246
rect 4321 12228 4327 12246
rect 4209 12158 4215 12176
rect 4321 12158 4327 12176
rect 4261 12106 4275 12112
rect 4209 12100 4327 12106
rect 4486 13452 4604 13458
rect 4538 13400 4552 13452
rect 4486 13383 4604 13400
rect 4538 13331 4552 13383
rect 4486 13314 4604 13331
rect 4538 13262 4552 13314
rect 4486 13245 4604 13262
rect 4538 13193 4552 13245
rect 4486 13176 4604 13193
rect 4538 13154 4552 13176
rect 4486 13107 4492 13124
rect 4598 13107 4604 13124
rect 4486 13038 4492 13055
rect 4598 13038 4604 13055
rect 4486 12968 4492 12986
rect 4598 12968 4604 12986
rect 4486 12898 4492 12916
rect 4598 12898 4604 12916
rect 4486 12112 4492 12846
rect 4598 12112 4604 12846
rect 4486 12100 4604 12112
rect 4763 13446 4881 13458
rect 4763 13412 4769 13446
rect 4803 13412 4841 13446
rect 4875 13412 4881 13446
rect 4763 13373 4881 13412
rect 4763 13339 4769 13373
rect 4803 13339 4841 13373
rect 4875 13339 4881 13373
rect 4763 13300 4881 13339
rect 4763 13266 4769 13300
rect 4803 13266 4841 13300
rect 4875 13266 4881 13300
rect 4763 13227 4881 13266
rect 4763 13193 4769 13227
rect 4803 13193 4841 13227
rect 4875 13193 4881 13227
rect 4763 13154 4881 13193
rect 4763 12714 4769 13154
rect 4875 12714 4881 13154
rect 4763 12645 4769 12662
rect 4875 12645 4881 12662
rect 4763 12576 4769 12593
rect 4875 12576 4881 12593
rect 4763 12507 4769 12524
rect 4875 12507 4881 12524
rect 4763 12438 4769 12455
rect 4875 12438 4881 12455
rect 4763 12368 4769 12386
rect 4875 12368 4881 12386
rect 4763 12298 4769 12316
rect 4875 12298 4881 12316
rect 4763 12228 4769 12246
rect 4875 12228 4881 12246
rect 4763 12158 4769 12176
rect 4875 12158 4881 12176
rect 4815 12106 4829 12112
rect 4763 12100 4881 12106
rect 5040 13452 5158 13458
rect 5092 13400 5106 13452
rect 5040 13383 5158 13400
rect 5092 13331 5106 13383
rect 5040 13314 5158 13331
rect 5092 13262 5106 13314
rect 5040 13245 5158 13262
rect 5092 13193 5106 13245
rect 5040 13176 5158 13193
rect 5092 13154 5106 13176
rect 5040 13107 5046 13124
rect 5152 13107 5158 13124
rect 5040 13038 5046 13055
rect 5152 13038 5158 13055
rect 5040 12968 5046 12986
rect 5152 12968 5158 12986
rect 5040 12898 5046 12916
rect 5152 12898 5158 12916
rect 5040 12112 5046 12846
rect 5152 12112 5158 12846
rect 5040 12100 5158 12112
rect 5317 13446 5435 13458
rect 5317 13412 5323 13446
rect 5357 13412 5395 13446
rect 5429 13412 5435 13446
rect 5317 13373 5435 13412
rect 5317 13339 5323 13373
rect 5357 13339 5395 13373
rect 5429 13339 5435 13373
rect 5317 13300 5435 13339
rect 5317 13266 5323 13300
rect 5357 13266 5395 13300
rect 5429 13266 5435 13300
rect 5317 13227 5435 13266
rect 5317 13193 5323 13227
rect 5357 13193 5395 13227
rect 5429 13193 5435 13227
rect 5317 13154 5435 13193
rect 5317 12714 5323 13154
rect 5429 12714 5435 13154
rect 5317 12645 5323 12662
rect 5429 12645 5435 12662
rect 5317 12576 5323 12593
rect 5429 12576 5435 12593
rect 5317 12507 5323 12524
rect 5429 12507 5435 12524
rect 5317 12438 5323 12455
rect 5429 12438 5435 12455
rect 5317 12368 5323 12386
rect 5429 12368 5435 12386
rect 5317 12298 5323 12316
rect 5429 12298 5435 12316
rect 5317 12228 5323 12246
rect 5429 12228 5435 12246
rect 5317 12158 5323 12176
rect 5429 12158 5435 12176
rect 5369 12106 5383 12112
rect 5317 12100 5435 12106
rect 5594 13452 5712 13458
rect 5646 13400 5660 13452
rect 5594 13383 5712 13400
rect 5646 13331 5660 13383
rect 5594 13314 5712 13331
rect 5646 13262 5660 13314
rect 5594 13245 5712 13262
rect 5646 13193 5660 13245
rect 5594 13176 5712 13193
rect 5646 13154 5660 13176
rect 5594 13107 5600 13124
rect 5706 13107 5712 13124
rect 5594 13038 5600 13055
rect 5706 13038 5712 13055
rect 5594 12968 5600 12986
rect 5706 12968 5712 12986
rect 5594 12898 5600 12916
rect 5706 12898 5712 12916
rect 5594 12112 5600 12846
rect 5706 12112 5712 12846
rect 5594 12100 5712 12112
rect 5871 13446 5989 13458
rect 5871 13412 5877 13446
rect 5911 13412 5949 13446
rect 5983 13412 5989 13446
rect 5871 13373 5989 13412
rect 5871 13339 5877 13373
rect 5911 13339 5949 13373
rect 5983 13339 5989 13373
rect 5871 13300 5989 13339
rect 5871 13266 5877 13300
rect 5911 13266 5949 13300
rect 5983 13266 5989 13300
rect 5871 13227 5989 13266
rect 5871 13193 5877 13227
rect 5911 13193 5949 13227
rect 5983 13193 5989 13227
rect 5871 13154 5989 13193
rect 5871 12714 5877 13154
rect 5983 12714 5989 13154
rect 5871 12645 5877 12662
rect 5983 12645 5989 12662
rect 5871 12576 5877 12593
rect 5983 12576 5989 12593
rect 5871 12507 5877 12524
rect 5983 12507 5989 12524
rect 5871 12438 5877 12455
rect 5983 12438 5989 12455
rect 5871 12368 5877 12386
rect 5983 12368 5989 12386
rect 5871 12298 5877 12316
rect 5983 12298 5989 12316
rect 5871 12228 5877 12246
rect 5983 12228 5989 12246
rect 5871 12158 5877 12176
rect 5983 12158 5989 12176
rect 5923 12106 5937 12112
rect 5871 12100 5989 12106
rect 6148 13452 6266 13458
rect 6200 13400 6214 13452
rect 6148 13383 6266 13400
rect 6200 13331 6214 13383
rect 6148 13314 6266 13331
rect 6200 13262 6214 13314
rect 6148 13245 6266 13262
rect 6200 13193 6214 13245
rect 6148 13176 6266 13193
rect 6200 13154 6214 13176
rect 6148 13107 6154 13124
rect 6260 13107 6266 13124
rect 6148 13038 6154 13055
rect 6260 13038 6266 13055
rect 6148 12968 6154 12986
rect 6260 12968 6266 12986
rect 6148 12898 6154 12916
rect 6260 12898 6266 12916
rect 6148 12112 6154 12846
rect 6260 12112 6266 12846
rect 6148 12100 6266 12112
rect 6425 13446 6543 13458
rect 6425 13412 6431 13446
rect 6465 13412 6503 13446
rect 6537 13412 6543 13446
rect 6425 13373 6543 13412
rect 6425 13339 6431 13373
rect 6465 13339 6503 13373
rect 6537 13339 6543 13373
rect 6425 13300 6543 13339
rect 6425 13266 6431 13300
rect 6465 13266 6503 13300
rect 6537 13266 6543 13300
rect 6425 13227 6543 13266
rect 6425 13193 6431 13227
rect 6465 13193 6503 13227
rect 6537 13193 6543 13227
rect 6425 13154 6543 13193
rect 6425 12714 6431 13154
rect 6537 12714 6543 13154
rect 6425 12645 6431 12662
rect 6537 12645 6543 12662
rect 6425 12576 6431 12593
rect 6537 12576 6543 12593
rect 6425 12507 6431 12524
rect 6537 12507 6543 12524
rect 6425 12438 6431 12455
rect 6537 12438 6543 12455
rect 6425 12368 6431 12386
rect 6537 12368 6543 12386
rect 6425 12298 6431 12316
rect 6537 12298 6543 12316
rect 6425 12228 6431 12246
rect 6537 12228 6543 12246
rect 6425 12158 6431 12176
rect 6537 12158 6543 12176
rect 6477 12106 6491 12112
rect 6425 12100 6543 12106
rect 6702 13452 6820 13458
rect 6754 13400 6768 13452
rect 6702 13383 6820 13400
rect 6754 13331 6768 13383
rect 6702 13314 6820 13331
rect 6754 13262 6768 13314
rect 6702 13245 6820 13262
rect 6754 13193 6768 13245
rect 6702 13176 6820 13193
rect 6754 13154 6768 13176
rect 6702 13107 6708 13124
rect 6814 13107 6820 13124
rect 6702 13038 6708 13055
rect 6814 13038 6820 13055
rect 6702 12968 6708 12986
rect 6814 12968 6820 12986
rect 6702 12898 6708 12916
rect 6814 12898 6820 12916
rect 6702 12112 6708 12846
rect 6814 12112 6820 12846
rect 6702 12100 6820 12112
rect 6979 13446 7097 13458
rect 6979 13412 6985 13446
rect 7019 13412 7057 13446
rect 7091 13412 7097 13446
rect 6979 13373 7097 13412
rect 6979 13339 6985 13373
rect 7019 13339 7057 13373
rect 7091 13339 7097 13373
rect 6979 13300 7097 13339
rect 6979 13266 6985 13300
rect 7019 13266 7057 13300
rect 7091 13266 7097 13300
rect 6979 13227 7097 13266
rect 6979 13193 6985 13227
rect 7019 13193 7057 13227
rect 7091 13193 7097 13227
rect 6979 13154 7097 13193
rect 6979 12714 6985 13154
rect 7091 12714 7097 13154
rect 6979 12645 6985 12662
rect 7091 12645 7097 12662
rect 6979 12576 6985 12593
rect 7091 12576 7097 12593
rect 6979 12507 6985 12524
rect 7091 12507 7097 12524
rect 6979 12438 6985 12455
rect 7091 12438 7097 12455
rect 6979 12368 6985 12386
rect 7091 12368 7097 12386
rect 6979 12298 6985 12316
rect 7091 12298 7097 12316
rect 6979 12228 6985 12246
rect 7091 12228 7097 12246
rect 6979 12158 6985 12176
rect 7091 12158 7097 12176
rect 7031 12106 7045 12112
rect 6979 12100 7097 12106
rect 7256 13452 7374 13458
rect 7308 13400 7322 13452
rect 7256 13383 7374 13400
rect 7308 13331 7322 13383
rect 7256 13314 7374 13331
rect 7308 13262 7322 13314
rect 7256 13245 7374 13262
rect 7308 13193 7322 13245
rect 7256 13176 7374 13193
rect 7308 13154 7322 13176
rect 7256 13107 7262 13124
rect 7368 13107 7374 13124
rect 7256 13038 7262 13055
rect 7368 13038 7374 13055
rect 7256 12968 7262 12986
rect 7368 12968 7374 12986
rect 7256 12898 7262 12916
rect 7368 12898 7374 12916
rect 7256 12112 7262 12846
rect 7368 12112 7374 12846
rect 7256 12100 7374 12112
rect 7533 13446 7651 13458
rect 7533 13412 7539 13446
rect 7573 13412 7611 13446
rect 7645 13412 7651 13446
rect 7533 13373 7651 13412
rect 7533 13339 7539 13373
rect 7573 13339 7611 13373
rect 7645 13339 7651 13373
rect 7533 13300 7651 13339
rect 7533 13266 7539 13300
rect 7573 13266 7611 13300
rect 7645 13266 7651 13300
rect 7533 13227 7651 13266
rect 7533 13193 7539 13227
rect 7573 13193 7611 13227
rect 7645 13193 7651 13227
rect 7533 13154 7651 13193
rect 7533 12714 7539 13154
rect 7645 12714 7651 13154
rect 7533 12645 7539 12662
rect 7645 12645 7651 12662
rect 7533 12576 7539 12593
rect 7645 12576 7651 12593
rect 7533 12507 7539 12524
rect 7645 12507 7651 12524
rect 7533 12438 7539 12455
rect 7645 12438 7651 12455
rect 7533 12368 7539 12386
rect 7645 12368 7651 12386
rect 7533 12298 7539 12316
rect 7645 12298 7651 12316
rect 7533 12228 7539 12246
rect 7645 12228 7651 12246
rect 7533 12158 7539 12176
rect 7645 12158 7651 12176
rect 7585 12106 7599 12112
rect 7533 12100 7651 12106
rect 7810 13452 7928 13458
rect 7862 13400 7876 13452
rect 7810 13383 7928 13400
rect 7862 13331 7876 13383
rect 7810 13314 7928 13331
rect 7862 13262 7876 13314
rect 7810 13245 7928 13262
rect 7862 13193 7876 13245
rect 7810 13176 7928 13193
rect 7862 13154 7876 13176
rect 7810 13107 7816 13124
rect 7922 13107 7928 13124
rect 7810 13038 7816 13055
rect 7922 13038 7928 13055
rect 7810 12968 7816 12986
rect 7922 12968 7928 12986
rect 7810 12898 7816 12916
rect 7922 12898 7928 12916
rect 7810 12112 7816 12846
rect 7922 12112 7928 12846
rect 7810 12100 7928 12112
rect 8044 13456 8224 13475
rect 8044 13404 8047 13456
rect 8099 13404 8169 13456
rect 8221 13404 8224 13456
rect 8044 13403 8184 13404
rect 8218 13403 8224 13404
rect 8044 13387 8224 13403
rect 8044 13335 8047 13387
rect 8099 13335 8169 13387
rect 8221 13335 8224 13387
rect 8044 13331 8184 13335
rect 8218 13331 8224 13335
rect 8044 13318 8224 13331
rect 8044 13266 8047 13318
rect 8099 13266 8169 13318
rect 8221 13266 8224 13318
rect 8044 13259 8184 13266
rect 8218 13259 8224 13266
rect 8044 13249 8224 13259
rect 8044 13197 8047 13249
rect 8099 13197 8169 13249
rect 8221 13197 8224 13249
rect 8044 13187 8184 13197
rect 8218 13187 8224 13197
rect 8044 13180 8224 13187
rect 8044 13128 8047 13180
rect 8099 13128 8169 13180
rect 8221 13128 8224 13180
rect 8044 13125 8050 13128
rect 8084 13125 8184 13128
rect 8044 13115 8184 13125
rect 8218 13115 8224 13128
rect 8044 13110 8224 13115
rect 8044 13058 8047 13110
rect 8099 13058 8169 13110
rect 8221 13058 8224 13110
rect 8044 13053 8050 13058
rect 8084 13053 8184 13058
rect 8044 13043 8184 13053
rect 8218 13043 8224 13058
rect 8044 13040 8224 13043
rect 8044 12988 8047 13040
rect 8099 12988 8169 13040
rect 8221 12988 8224 13040
rect 8044 12981 8050 12988
rect 8084 12981 8184 12988
rect 8044 12971 8184 12981
rect 8218 12971 8224 12988
rect 8044 12970 8224 12971
rect 8044 12918 8047 12970
rect 8099 12918 8169 12970
rect 8221 12918 8224 12970
rect 8044 12908 8050 12918
rect 8084 12908 8184 12918
rect 8044 12900 8184 12908
rect 8218 12900 8224 12918
rect 8044 12848 8047 12900
rect 8099 12848 8169 12900
rect 8221 12848 8224 12900
rect 8044 12835 8050 12848
rect 8084 12835 8184 12848
rect 8044 12827 8184 12835
rect 8218 12827 8224 12848
rect 8044 12796 8224 12827
rect 8044 12762 8050 12796
rect 8084 12789 8224 12796
rect 8084 12762 8184 12789
rect 8044 12755 8184 12762
rect 8218 12755 8224 12789
rect 8044 12723 8224 12755
rect 8044 12689 8050 12723
rect 8084 12717 8224 12723
rect 8084 12689 8184 12717
rect 8044 12683 8184 12689
rect 8218 12683 8224 12717
rect 8044 12650 8224 12683
rect 8044 12616 8050 12650
rect 8084 12645 8224 12650
rect 8084 12616 8184 12645
rect 8044 12611 8184 12616
rect 8218 12611 8224 12645
rect 8044 12577 8224 12611
rect 8044 12543 8050 12577
rect 8084 12573 8224 12577
rect 8084 12543 8184 12573
rect 8044 12539 8184 12543
rect 8218 12539 8224 12573
rect 8044 12504 8224 12539
rect 8044 12470 8050 12504
rect 8084 12501 8224 12504
rect 8084 12470 8184 12501
rect 8044 12467 8184 12470
rect 8218 12467 8224 12501
rect 8044 12431 8224 12467
rect 8044 12397 8050 12431
rect 8084 12429 8224 12431
rect 8084 12397 8184 12429
rect 8044 12395 8184 12397
rect 8218 12395 8224 12429
rect 8044 12358 8224 12395
rect 8044 12324 8050 12358
rect 8084 12357 8224 12358
rect 8084 12324 8184 12357
rect 8044 12323 8184 12324
rect 8218 12323 8224 12357
rect 8044 12285 8224 12323
rect 8044 12251 8050 12285
rect 8084 12251 8184 12285
rect 8218 12251 8224 12285
rect 8044 12212 8224 12251
rect 8044 12178 8050 12212
rect 8084 12178 8184 12212
rect 8218 12178 8224 12212
rect 8044 12139 8224 12178
rect 8044 12105 8050 12139
rect 8084 12105 8184 12139
rect 8218 12105 8224 12139
rect 8044 12066 8224 12105
rect 8044 12032 8050 12066
rect 8084 12032 8184 12066
rect 8218 12032 8224 12066
rect 8044 11993 8224 12032
tri 2712 11959 2736 11983 sw
rect 8044 11959 8050 11993
rect 8084 11959 8184 11993
rect 8218 11959 8224 11993
rect 2580 11936 2736 11959
tri 2736 11936 2759 11959 sw
rect 2580 11920 2759 11936
tri 2759 11920 2775 11936 sw
rect 8044 11920 8224 11959
rect 2580 11895 2775 11920
tri 2775 11895 2800 11920 sw
rect 2580 11818 7748 11895
rect 2580 11784 3035 11818
rect 3069 11784 3108 11818
rect 3142 11784 3181 11818
rect 3215 11784 3254 11818
rect 3288 11784 3327 11818
rect 3361 11784 3400 11818
rect 3434 11784 3473 11818
rect 3507 11784 3546 11818
rect 3580 11784 3619 11818
rect 3653 11784 3692 11818
rect 3726 11784 3765 11818
rect 3799 11784 3838 11818
rect 3872 11784 3911 11818
rect 3945 11784 3984 11818
rect 4018 11784 4057 11818
rect 4091 11784 4130 11818
rect 4164 11784 4203 11818
rect 4237 11784 4276 11818
rect 4310 11784 4349 11818
rect 4383 11784 4422 11818
rect 4456 11784 4495 11818
rect 4529 11784 4568 11818
rect 4602 11784 4641 11818
rect 4675 11784 4714 11818
rect 4748 11784 4787 11818
rect 4821 11784 4860 11818
rect 4894 11784 4933 11818
rect 4967 11784 5006 11818
rect 5040 11784 5079 11818
rect 5113 11784 5152 11818
rect 5186 11784 5225 11818
rect 5259 11784 5298 11818
rect 5332 11784 5371 11818
rect 5405 11784 5444 11818
rect 5478 11784 5517 11818
rect 5551 11784 5590 11818
rect 5624 11784 5663 11818
rect 5697 11784 5736 11818
rect 5770 11784 5809 11818
rect 5843 11784 5881 11818
rect 5915 11784 5953 11818
rect 5987 11784 6025 11818
rect 6059 11784 6097 11818
rect 6131 11784 6169 11818
rect 6203 11784 6241 11818
rect 6275 11784 6313 11818
rect 6347 11784 6385 11818
rect 6419 11784 6457 11818
rect 6491 11784 6529 11818
rect 6563 11784 6601 11818
rect 6635 11784 6673 11818
rect 6707 11784 6745 11818
rect 6779 11784 6817 11818
rect 6851 11784 6889 11818
rect 6923 11784 6961 11818
rect 6995 11784 7033 11818
rect 7067 11784 7105 11818
rect 7139 11784 7177 11818
rect 7211 11784 7249 11818
rect 7283 11784 7321 11818
rect 7355 11784 7393 11818
rect 7427 11784 7465 11818
rect 7499 11784 7537 11818
rect 7571 11784 7609 11818
rect 7643 11784 7681 11818
rect 7715 11784 7748 11818
rect 2580 11752 7748 11784
rect 8044 11886 8050 11920
rect 8084 11886 8184 11920
rect 8218 11886 8224 11920
rect 8044 11847 8224 11886
rect 8044 11813 8050 11847
rect 8084 11813 8184 11847
rect 8218 11813 8224 11847
rect 8044 11774 8224 11813
rect 2580 11740 2797 11752
tri 2797 11740 2809 11752 nw
rect 8044 11740 8050 11774
rect 8084 11740 8184 11774
rect 8218 11740 8224 11774
rect 2580 11717 2774 11740
tri 2774 11717 2797 11740 nw
rect 2580 11701 2758 11717
tri 2758 11701 2774 11717 nw
rect 8044 11701 8224 11740
rect 2580 11667 2724 11701
tri 2724 11667 2758 11701 nw
rect 8044 11667 8050 11701
rect 8084 11667 8184 11701
rect 8218 11667 8224 11701
rect 2580 10522 2712 11667
tri 2712 11655 2724 11667 nw
rect 8044 11628 8224 11667
rect 8044 11594 8050 11628
rect 8084 11594 8184 11628
rect 8218 11594 8224 11628
rect 8044 11555 8224 11594
rect 8044 11521 8050 11555
rect 8084 11521 8184 11555
rect 8218 11521 8224 11555
rect 8044 11482 8224 11521
rect 2632 10470 2660 10522
rect 2580 10456 2712 10470
rect 2632 10404 2660 10456
rect 2580 10390 2712 10404
rect 2632 10338 2660 10390
rect 2580 10324 2712 10338
rect 2632 10272 2660 10324
rect 2580 10258 2712 10272
rect 2632 10206 2660 10258
rect 2580 10192 2712 10206
rect 2632 10140 2660 10192
rect 2580 10126 2712 10140
rect 2632 10074 2660 10126
rect 2824 11452 2942 11458
rect 2876 11400 2890 11452
rect 2824 11383 2942 11400
rect 2876 11331 2890 11383
rect 2824 11314 2942 11331
rect 2876 11262 2890 11314
rect 2824 11245 2942 11262
rect 2876 11193 2890 11245
rect 2824 11176 2942 11193
rect 2876 11154 2890 11176
rect 2824 11107 2830 11124
rect 2936 11107 2942 11124
rect 2824 11038 2830 11055
rect 2936 11038 2942 11055
rect 2824 10968 2830 10986
rect 2936 10968 2942 10986
rect 2824 10898 2830 10916
rect 2936 10898 2942 10916
rect 2824 10112 2830 10846
rect 2936 10112 2942 10846
rect 2824 10100 2942 10112
rect 3101 11446 3219 11458
rect 3101 11412 3107 11446
rect 3141 11412 3179 11446
rect 3213 11412 3219 11446
rect 3101 11373 3219 11412
rect 3101 11339 3107 11373
rect 3141 11339 3179 11373
rect 3213 11339 3219 11373
rect 3101 11300 3219 11339
rect 3101 11266 3107 11300
rect 3141 11266 3179 11300
rect 3213 11266 3219 11300
rect 3101 11227 3219 11266
rect 3101 11193 3107 11227
rect 3141 11193 3179 11227
rect 3213 11193 3219 11227
rect 3101 11154 3219 11193
rect 3101 10714 3107 11154
rect 3213 10714 3219 11154
rect 3101 10645 3107 10662
rect 3213 10645 3219 10662
rect 3101 10576 3107 10593
rect 3213 10576 3219 10593
rect 3101 10507 3107 10524
rect 3213 10507 3219 10524
rect 3101 10438 3107 10455
rect 3213 10438 3219 10455
rect 3101 10368 3107 10386
rect 3213 10368 3219 10386
rect 3101 10298 3107 10316
rect 3213 10298 3219 10316
rect 3101 10228 3107 10246
rect 3213 10228 3219 10246
rect 3101 10158 3107 10176
rect 3213 10158 3219 10176
rect 3153 10106 3167 10112
rect 3101 10100 3219 10106
rect 3378 11452 3496 11458
rect 3430 11400 3444 11452
rect 3378 11383 3496 11400
rect 3430 11331 3444 11383
rect 3378 11314 3496 11331
rect 3430 11262 3444 11314
rect 3378 11245 3496 11262
rect 3430 11193 3444 11245
rect 3378 11176 3496 11193
rect 3430 11154 3444 11176
rect 3378 11107 3384 11124
rect 3490 11107 3496 11124
rect 3378 11038 3384 11055
rect 3490 11038 3496 11055
rect 3378 10968 3384 10986
rect 3490 10968 3496 10986
rect 3378 10898 3384 10916
rect 3490 10898 3496 10916
rect 3378 10112 3384 10846
rect 3490 10112 3496 10846
rect 3378 10100 3496 10112
rect 3655 11446 3773 11458
rect 3655 11412 3661 11446
rect 3695 11412 3733 11446
rect 3767 11412 3773 11446
rect 3655 11373 3773 11412
rect 3655 11339 3661 11373
rect 3695 11339 3733 11373
rect 3767 11339 3773 11373
rect 3655 11300 3773 11339
rect 3655 11266 3661 11300
rect 3695 11266 3733 11300
rect 3767 11266 3773 11300
rect 3655 11227 3773 11266
rect 3655 11193 3661 11227
rect 3695 11193 3733 11227
rect 3767 11193 3773 11227
rect 3655 11154 3773 11193
rect 3655 10714 3661 11154
rect 3767 10714 3773 11154
rect 3655 10645 3661 10662
rect 3767 10645 3773 10662
rect 3655 10576 3661 10593
rect 3767 10576 3773 10593
rect 3655 10507 3661 10524
rect 3767 10507 3773 10524
rect 3655 10438 3661 10455
rect 3767 10438 3773 10455
rect 3655 10368 3661 10386
rect 3767 10368 3773 10386
rect 3655 10298 3661 10316
rect 3767 10298 3773 10316
rect 3655 10228 3661 10246
rect 3767 10228 3773 10246
rect 3655 10158 3661 10176
rect 3767 10158 3773 10176
rect 3707 10106 3721 10112
rect 3655 10100 3773 10106
rect 3932 11452 4050 11458
rect 3984 11400 3998 11452
rect 3932 11383 4050 11400
rect 3984 11331 3998 11383
rect 3932 11314 4050 11331
rect 3984 11262 3998 11314
rect 3932 11245 4050 11262
rect 3984 11193 3998 11245
rect 3932 11176 4050 11193
rect 3984 11154 3998 11176
rect 3932 11107 3938 11124
rect 4044 11107 4050 11124
rect 3932 11038 3938 11055
rect 4044 11038 4050 11055
rect 3932 10968 3938 10986
rect 4044 10968 4050 10986
rect 3932 10898 3938 10916
rect 4044 10898 4050 10916
rect 3932 10112 3938 10846
rect 4044 10112 4050 10846
rect 3932 10100 4050 10112
rect 4209 11446 4327 11458
rect 4209 11412 4215 11446
rect 4249 11412 4287 11446
rect 4321 11412 4327 11446
rect 4209 11373 4327 11412
rect 4209 11339 4215 11373
rect 4249 11339 4287 11373
rect 4321 11339 4327 11373
rect 4209 11300 4327 11339
rect 4209 11266 4215 11300
rect 4249 11266 4287 11300
rect 4321 11266 4327 11300
rect 4209 11227 4327 11266
rect 4209 11193 4215 11227
rect 4249 11193 4287 11227
rect 4321 11193 4327 11227
rect 4209 11154 4327 11193
rect 4209 10714 4215 11154
rect 4321 10714 4327 11154
rect 4209 10645 4215 10662
rect 4321 10645 4327 10662
rect 4209 10576 4215 10593
rect 4321 10576 4327 10593
rect 4209 10507 4215 10524
rect 4321 10507 4327 10524
rect 4209 10438 4215 10455
rect 4321 10438 4327 10455
rect 4209 10368 4215 10386
rect 4321 10368 4327 10386
rect 4209 10298 4215 10316
rect 4321 10298 4327 10316
rect 4209 10228 4215 10246
rect 4321 10228 4327 10246
rect 4209 10158 4215 10176
rect 4321 10158 4327 10176
rect 4261 10106 4275 10112
rect 4209 10100 4327 10106
rect 4486 11452 4604 11458
rect 4538 11400 4552 11452
rect 4486 11383 4604 11400
rect 4538 11331 4552 11383
rect 4486 11314 4604 11331
rect 4538 11262 4552 11314
rect 4486 11245 4604 11262
rect 4538 11193 4552 11245
rect 4486 11176 4604 11193
rect 4538 11154 4552 11176
rect 4486 11107 4492 11124
rect 4598 11107 4604 11124
rect 4486 11038 4492 11055
rect 4598 11038 4604 11055
rect 4486 10968 4492 10986
rect 4598 10968 4604 10986
rect 4486 10898 4492 10916
rect 4598 10898 4604 10916
rect 4486 10112 4492 10846
rect 4598 10112 4604 10846
rect 4486 10100 4604 10112
rect 4763 11446 4881 11458
rect 4763 11412 4769 11446
rect 4803 11412 4841 11446
rect 4875 11412 4881 11446
rect 4763 11373 4881 11412
rect 4763 11339 4769 11373
rect 4803 11339 4841 11373
rect 4875 11339 4881 11373
rect 4763 11300 4881 11339
rect 4763 11266 4769 11300
rect 4803 11266 4841 11300
rect 4875 11266 4881 11300
rect 4763 11227 4881 11266
rect 4763 11193 4769 11227
rect 4803 11193 4841 11227
rect 4875 11193 4881 11227
rect 4763 11154 4881 11193
rect 4763 10714 4769 11154
rect 4875 10714 4881 11154
rect 4763 10645 4769 10662
rect 4875 10645 4881 10662
rect 4763 10576 4769 10593
rect 4875 10576 4881 10593
rect 4763 10507 4769 10524
rect 4875 10507 4881 10524
rect 4763 10438 4769 10455
rect 4875 10438 4881 10455
rect 4763 10368 4769 10386
rect 4875 10368 4881 10386
rect 4763 10298 4769 10316
rect 4875 10298 4881 10316
rect 4763 10228 4769 10246
rect 4875 10228 4881 10246
rect 4763 10158 4769 10176
rect 4875 10158 4881 10176
rect 4815 10106 4829 10112
rect 4763 10100 4881 10106
rect 5040 11452 5158 11458
rect 5092 11400 5106 11452
rect 5040 11383 5158 11400
rect 5092 11331 5106 11383
rect 5040 11314 5158 11331
rect 5092 11262 5106 11314
rect 5040 11245 5158 11262
rect 5092 11193 5106 11245
rect 5040 11176 5158 11193
rect 5092 11154 5106 11176
rect 5040 11107 5046 11124
rect 5152 11107 5158 11124
rect 5040 11038 5046 11055
rect 5152 11038 5158 11055
rect 5040 10968 5046 10986
rect 5152 10968 5158 10986
rect 5040 10898 5046 10916
rect 5152 10898 5158 10916
rect 5040 10112 5046 10846
rect 5152 10112 5158 10846
rect 5040 10100 5158 10112
rect 5317 11446 5435 11458
rect 5317 11412 5323 11446
rect 5357 11412 5395 11446
rect 5429 11412 5435 11446
rect 5317 11373 5435 11412
rect 5317 11339 5323 11373
rect 5357 11339 5395 11373
rect 5429 11339 5435 11373
rect 5317 11300 5435 11339
rect 5317 11266 5323 11300
rect 5357 11266 5395 11300
rect 5429 11266 5435 11300
rect 5317 11227 5435 11266
rect 5317 11193 5323 11227
rect 5357 11193 5395 11227
rect 5429 11193 5435 11227
rect 5317 11154 5435 11193
rect 5317 10714 5323 11154
rect 5429 10714 5435 11154
rect 5317 10645 5323 10662
rect 5429 10645 5435 10662
rect 5317 10576 5323 10593
rect 5429 10576 5435 10593
rect 5317 10507 5323 10524
rect 5429 10507 5435 10524
rect 5317 10438 5323 10455
rect 5429 10438 5435 10455
rect 5317 10368 5323 10386
rect 5429 10368 5435 10386
rect 5317 10298 5323 10316
rect 5429 10298 5435 10316
rect 5317 10228 5323 10246
rect 5429 10228 5435 10246
rect 5317 10158 5323 10176
rect 5429 10158 5435 10176
rect 5369 10106 5383 10112
rect 5317 10100 5435 10106
rect 5594 11452 5712 11458
rect 5646 11400 5660 11452
rect 5594 11383 5712 11400
rect 5646 11331 5660 11383
rect 5594 11314 5712 11331
rect 5646 11262 5660 11314
rect 5594 11245 5712 11262
rect 5646 11193 5660 11245
rect 5594 11176 5712 11193
rect 5646 11154 5660 11176
rect 5594 11107 5600 11124
rect 5706 11107 5712 11124
rect 5594 11038 5600 11055
rect 5706 11038 5712 11055
rect 5594 10968 5600 10986
rect 5706 10968 5712 10986
rect 5594 10898 5600 10916
rect 5706 10898 5712 10916
rect 5594 10112 5600 10846
rect 5706 10112 5712 10846
rect 5594 10100 5712 10112
rect 5871 11446 5989 11458
rect 5871 11412 5877 11446
rect 5911 11412 5949 11446
rect 5983 11412 5989 11446
rect 5871 11373 5989 11412
rect 5871 11339 5877 11373
rect 5911 11339 5949 11373
rect 5983 11339 5989 11373
rect 5871 11300 5989 11339
rect 5871 11266 5877 11300
rect 5911 11266 5949 11300
rect 5983 11266 5989 11300
rect 5871 11227 5989 11266
rect 5871 11193 5877 11227
rect 5911 11193 5949 11227
rect 5983 11193 5989 11227
rect 5871 11154 5989 11193
rect 5871 10714 5877 11154
rect 5983 10714 5989 11154
rect 5871 10645 5877 10662
rect 5983 10645 5989 10662
rect 5871 10576 5877 10593
rect 5983 10576 5989 10593
rect 5871 10507 5877 10524
rect 5983 10507 5989 10524
rect 5871 10438 5877 10455
rect 5983 10438 5989 10455
rect 5871 10368 5877 10386
rect 5983 10368 5989 10386
rect 5871 10298 5877 10316
rect 5983 10298 5989 10316
rect 5871 10228 5877 10246
rect 5983 10228 5989 10246
rect 5871 10158 5877 10176
rect 5983 10158 5989 10176
rect 5923 10106 5937 10112
rect 5871 10100 5989 10106
rect 6148 11452 6266 11458
rect 6200 11400 6214 11452
rect 6148 11383 6266 11400
rect 6200 11331 6214 11383
rect 6148 11314 6266 11331
rect 6200 11262 6214 11314
rect 6148 11245 6266 11262
rect 6200 11193 6214 11245
rect 6148 11176 6266 11193
rect 6200 11154 6214 11176
rect 6148 11107 6154 11124
rect 6260 11107 6266 11124
rect 6148 11038 6154 11055
rect 6260 11038 6266 11055
rect 6148 10968 6154 10986
rect 6260 10968 6266 10986
rect 6148 10898 6154 10916
rect 6260 10898 6266 10916
rect 6148 10112 6154 10846
rect 6260 10112 6266 10846
rect 6148 10100 6266 10112
rect 6425 11446 6543 11458
rect 6425 11412 6431 11446
rect 6465 11412 6503 11446
rect 6537 11412 6543 11446
rect 6425 11373 6543 11412
rect 6425 11339 6431 11373
rect 6465 11339 6503 11373
rect 6537 11339 6543 11373
rect 6425 11300 6543 11339
rect 6425 11266 6431 11300
rect 6465 11266 6503 11300
rect 6537 11266 6543 11300
rect 6425 11227 6543 11266
rect 6425 11193 6431 11227
rect 6465 11193 6503 11227
rect 6537 11193 6543 11227
rect 6425 11154 6543 11193
rect 6425 10714 6431 11154
rect 6537 10714 6543 11154
rect 6425 10645 6431 10662
rect 6537 10645 6543 10662
rect 6425 10576 6431 10593
rect 6537 10576 6543 10593
rect 6425 10507 6431 10524
rect 6537 10507 6543 10524
rect 6425 10438 6431 10455
rect 6537 10438 6543 10455
rect 6425 10368 6431 10386
rect 6537 10368 6543 10386
rect 6425 10298 6431 10316
rect 6537 10298 6543 10316
rect 6425 10228 6431 10246
rect 6537 10228 6543 10246
rect 6425 10158 6431 10176
rect 6537 10158 6543 10176
rect 6477 10106 6491 10112
rect 6425 10100 6543 10106
rect 6702 11452 6820 11458
rect 6754 11400 6768 11452
rect 6702 11383 6820 11400
rect 6754 11331 6768 11383
rect 6702 11314 6820 11331
rect 6754 11262 6768 11314
rect 6702 11245 6820 11262
rect 6754 11193 6768 11245
rect 6702 11176 6820 11193
rect 6754 11154 6768 11176
rect 6702 11107 6708 11124
rect 6814 11107 6820 11124
rect 6702 11038 6708 11055
rect 6814 11038 6820 11055
rect 6702 10968 6708 10986
rect 6814 10968 6820 10986
rect 6702 10898 6708 10916
rect 6814 10898 6820 10916
rect 6702 10112 6708 10846
rect 6814 10112 6820 10846
rect 6702 10100 6820 10112
rect 6979 11446 7097 11458
rect 6979 11412 6985 11446
rect 7019 11412 7057 11446
rect 7091 11412 7097 11446
rect 6979 11373 7097 11412
rect 6979 11339 6985 11373
rect 7019 11339 7057 11373
rect 7091 11339 7097 11373
rect 6979 11300 7097 11339
rect 6979 11266 6985 11300
rect 7019 11266 7057 11300
rect 7091 11266 7097 11300
rect 6979 11227 7097 11266
rect 6979 11193 6985 11227
rect 7019 11193 7057 11227
rect 7091 11193 7097 11227
rect 6979 11154 7097 11193
rect 6979 10714 6985 11154
rect 7091 10714 7097 11154
rect 6979 10645 6985 10662
rect 7091 10645 7097 10662
rect 6979 10576 6985 10593
rect 7091 10576 7097 10593
rect 6979 10507 6985 10524
rect 7091 10507 7097 10524
rect 6979 10438 6985 10455
rect 7091 10438 7097 10455
rect 6979 10368 6985 10386
rect 7091 10368 7097 10386
rect 6979 10298 6985 10316
rect 7091 10298 7097 10316
rect 6979 10228 6985 10246
rect 7091 10228 7097 10246
rect 6979 10158 6985 10176
rect 7091 10158 7097 10176
rect 7031 10106 7045 10112
rect 6979 10100 7097 10106
rect 7256 11452 7374 11458
rect 7308 11400 7322 11452
rect 7256 11383 7374 11400
rect 7308 11331 7322 11383
rect 7256 11314 7374 11331
rect 7308 11262 7322 11314
rect 7256 11245 7374 11262
rect 7308 11193 7322 11245
rect 7256 11176 7374 11193
rect 7308 11154 7322 11176
rect 7256 11107 7262 11124
rect 7368 11107 7374 11124
rect 7256 11038 7262 11055
rect 7368 11038 7374 11055
rect 7256 10968 7262 10986
rect 7368 10968 7374 10986
rect 7256 10898 7262 10916
rect 7368 10898 7374 10916
rect 7256 10112 7262 10846
rect 7368 10112 7374 10846
rect 7256 10100 7374 10112
rect 7533 11446 7651 11458
rect 7533 11412 7539 11446
rect 7573 11412 7611 11446
rect 7645 11412 7651 11446
rect 7533 11373 7651 11412
rect 7533 11339 7539 11373
rect 7573 11339 7611 11373
rect 7645 11339 7651 11373
rect 7533 11300 7651 11339
rect 7533 11266 7539 11300
rect 7573 11266 7611 11300
rect 7645 11266 7651 11300
rect 7533 11227 7651 11266
rect 7533 11193 7539 11227
rect 7573 11193 7611 11227
rect 7645 11193 7651 11227
rect 7533 11154 7651 11193
rect 7533 10714 7539 11154
rect 7645 10714 7651 11154
rect 7533 10645 7539 10662
rect 7645 10645 7651 10662
rect 7533 10576 7539 10593
rect 7645 10576 7651 10593
rect 7533 10507 7539 10524
rect 7645 10507 7651 10524
rect 7533 10438 7539 10455
rect 7645 10438 7651 10455
rect 7533 10368 7539 10386
rect 7645 10368 7651 10386
rect 7533 10298 7539 10316
rect 7645 10298 7651 10316
rect 7533 10228 7539 10246
rect 7645 10228 7651 10246
rect 7533 10158 7539 10176
rect 7645 10158 7651 10176
rect 7585 10106 7599 10112
rect 7533 10100 7651 10106
rect 7810 11452 7928 11458
rect 7862 11400 7876 11452
rect 7810 11383 7928 11400
rect 7862 11331 7876 11383
rect 7810 11314 7928 11331
rect 7862 11262 7876 11314
rect 7810 11245 7928 11262
rect 7862 11193 7876 11245
rect 7810 11176 7928 11193
rect 7862 11154 7876 11176
rect 7810 11107 7816 11124
rect 7922 11107 7928 11124
rect 7810 11038 7816 11055
rect 7922 11038 7928 11055
rect 7810 10968 7816 10986
rect 7922 10968 7928 10986
rect 7810 10898 7816 10916
rect 7922 10898 7928 10916
rect 7810 10112 7816 10846
rect 7922 10112 7928 10846
rect 7810 10100 7928 10112
rect 8044 11456 8050 11482
rect 8084 11456 8184 11482
rect 8218 11456 8224 11482
rect 8044 11404 8047 11456
rect 8099 11404 8169 11456
rect 8221 11404 8224 11456
rect 8044 11387 8050 11404
rect 8084 11387 8184 11404
rect 8218 11387 8224 11404
rect 8044 11335 8047 11387
rect 8099 11335 8169 11387
rect 8221 11335 8224 11387
rect 8044 11318 8050 11335
rect 8084 11318 8184 11335
rect 8218 11318 8224 11335
rect 8044 11266 8047 11318
rect 8099 11266 8169 11318
rect 8221 11266 8224 11318
rect 8044 11263 8224 11266
rect 8044 11249 8050 11263
rect 8084 11249 8184 11263
rect 8218 11249 8224 11263
rect 8044 11197 8047 11249
rect 8099 11197 8169 11249
rect 8221 11197 8224 11249
rect 8044 11190 8224 11197
rect 8044 11180 8050 11190
rect 8084 11180 8184 11190
rect 8218 11180 8224 11190
rect 8044 11128 8047 11180
rect 8099 11128 8169 11180
rect 8221 11128 8224 11180
rect 8044 11117 8224 11128
rect 8044 11110 8050 11117
rect 8084 11110 8184 11117
rect 8218 11110 8224 11117
rect 8044 11058 8047 11110
rect 8099 11058 8169 11110
rect 8221 11058 8224 11110
rect 8044 11044 8224 11058
rect 8044 11040 8050 11044
rect 8084 11040 8184 11044
rect 8218 11040 8224 11044
rect 8044 10988 8047 11040
rect 8099 10988 8169 11040
rect 8221 10988 8224 11040
rect 8044 10971 8224 10988
rect 8044 10970 8050 10971
rect 8084 10970 8184 10971
rect 8218 10970 8224 10971
rect 8044 10918 8047 10970
rect 8099 10918 8169 10970
rect 8221 10918 8224 10970
rect 8044 10900 8224 10918
rect 8044 10848 8047 10900
rect 8099 10848 8169 10900
rect 8221 10848 8224 10900
rect 8044 10825 8224 10848
rect 8044 10791 8050 10825
rect 8084 10791 8184 10825
rect 8218 10791 8224 10825
rect 8044 10752 8224 10791
rect 8044 10718 8050 10752
rect 8084 10718 8184 10752
rect 8218 10718 8224 10752
rect 8044 10679 8224 10718
rect 8044 10645 8050 10679
rect 8084 10645 8184 10679
rect 8218 10645 8224 10679
rect 8044 10606 8224 10645
rect 8044 10572 8050 10606
rect 8084 10572 8184 10606
rect 8218 10572 8224 10606
rect 8044 10533 8224 10572
rect 8044 10499 8050 10533
rect 8084 10499 8184 10533
rect 8218 10499 8224 10533
rect 8044 10460 8224 10499
rect 8044 10426 8050 10460
rect 8084 10426 8184 10460
rect 8218 10426 8224 10460
rect 8044 10387 8224 10426
rect 8044 10353 8050 10387
rect 8084 10353 8184 10387
rect 8218 10353 8224 10387
rect 8044 10314 8224 10353
rect 8044 10280 8050 10314
rect 8084 10280 8184 10314
rect 8218 10280 8224 10314
rect 8044 10241 8224 10280
rect 8044 10207 8050 10241
rect 8084 10207 8184 10241
rect 8218 10207 8224 10241
rect 8044 10168 8224 10207
rect 8044 10134 8050 10168
rect 8084 10134 8184 10168
rect 8218 10134 8224 10168
rect 8044 10095 8224 10134
rect 2580 10061 2712 10074
tri 2712 10061 2739 10088 sw
rect 8044 10061 8050 10095
rect 8084 10061 8184 10095
rect 8218 10061 8224 10095
rect 2580 10060 2739 10061
rect 2632 10008 2660 10060
rect 2712 10056 2739 10060
tri 2739 10056 2744 10061 sw
rect 2712 10050 7729 10056
rect 2712 10016 3035 10050
rect 3069 10016 3108 10050
rect 3142 10016 3181 10050
rect 3215 10016 3254 10050
rect 3288 10016 3327 10050
rect 3361 10016 3400 10050
rect 3434 10016 3473 10050
rect 3507 10016 3546 10050
rect 3580 10016 3619 10050
rect 3653 10016 3692 10050
rect 3726 10016 3765 10050
rect 3799 10016 3838 10050
rect 3872 10016 3911 10050
rect 3945 10016 3984 10050
rect 4018 10016 4057 10050
rect 4091 10016 4130 10050
rect 4164 10016 4203 10050
rect 4237 10016 4276 10050
rect 4310 10016 4349 10050
rect 4383 10016 4422 10050
rect 4456 10016 4495 10050
rect 4529 10016 4568 10050
rect 4602 10016 4641 10050
rect 4675 10016 4714 10050
rect 4748 10016 4787 10050
rect 4821 10016 4860 10050
rect 4894 10016 4933 10050
rect 4967 10016 5006 10050
rect 5040 10016 5079 10050
rect 5113 10016 5152 10050
rect 5186 10016 5225 10050
rect 5259 10016 5298 10050
rect 5332 10016 5371 10050
rect 5405 10016 5444 10050
rect 5478 10016 5517 10050
rect 5551 10016 5590 10050
rect 5624 10016 5663 10050
rect 5697 10016 5736 10050
rect 5770 10016 5809 10050
rect 5843 10016 5882 10050
rect 5916 10016 5955 10050
rect 5989 10016 6027 10050
rect 6061 10016 6099 10050
rect 6133 10016 6171 10050
rect 6205 10016 6243 10050
rect 6277 10016 6315 10050
rect 6349 10016 6387 10050
rect 6421 10016 6459 10050
rect 6493 10016 6531 10050
rect 6565 10016 6603 10050
rect 6637 10016 6675 10050
rect 6709 10016 6747 10050
rect 6781 10016 6819 10050
rect 6853 10016 6891 10050
rect 6925 10016 6963 10050
rect 6997 10016 7035 10050
rect 7069 10016 7107 10050
rect 7141 10016 7179 10050
rect 7213 10016 7251 10050
rect 7285 10016 7323 10050
rect 7357 10016 7395 10050
rect 7429 10016 7467 10050
rect 7501 10016 7539 10050
rect 7573 10016 7611 10050
rect 7645 10016 7683 10050
rect 7717 10016 7729 10050
rect 2712 10008 7729 10016
rect 2580 10002 7729 10008
rect 8044 10022 8224 10061
rect 2270 9948 2450 9986
rect 2270 9914 2276 9948
rect 2310 9914 2410 9948
rect 2444 9914 2450 9948
rect 2270 9892 2450 9914
rect 8044 9988 8050 10022
rect 8084 9988 8184 10022
rect 8218 9988 8224 10022
rect 8044 9949 8224 9988
rect 8044 9915 8050 9949
rect 8084 9915 8184 9949
rect 8218 9915 8224 9949
tri 8039 9904 8044 9909 se
rect 8044 9904 8224 9915
tri 2450 9892 2462 9904 sw
tri 8027 9892 8039 9904 se
rect 8039 9892 8224 9904
rect 2270 9876 2462 9892
tri 2462 9876 2478 9892 sw
tri 8011 9876 8027 9892 se
rect 8027 9876 8224 9892
rect 2270 9842 2276 9876
rect 2310 9842 2410 9876
rect 2444 9870 8050 9876
rect 2444 9842 2482 9870
rect 2270 9836 2482 9842
rect 2516 9836 2555 9870
rect 2589 9836 2628 9870
rect 2662 9836 2701 9870
rect 2735 9836 2774 9870
rect 2808 9836 2847 9870
rect 2881 9836 2920 9870
rect 2954 9836 2993 9870
rect 3027 9836 3066 9870
rect 3100 9836 3139 9870
rect 3173 9836 3212 9870
rect 3246 9836 3285 9870
rect 3319 9836 3358 9870
rect 3392 9836 3431 9870
rect 3465 9836 3504 9870
rect 3538 9836 3577 9870
rect 3611 9836 3650 9870
rect 3684 9836 3723 9870
rect 3757 9836 3796 9870
rect 3830 9836 3869 9870
rect 3903 9836 3942 9870
rect 3976 9836 4015 9870
rect 4049 9836 4088 9870
rect 4122 9836 4161 9870
rect 4195 9836 4234 9870
rect 4268 9836 4306 9870
rect 4340 9836 4378 9870
rect 4412 9836 4450 9870
rect 4484 9836 4522 9870
rect 4556 9836 4594 9870
rect 4628 9836 4666 9870
rect 4700 9836 4738 9870
rect 4772 9836 4810 9870
rect 4844 9836 4882 9870
rect 4916 9836 4954 9870
rect 4988 9836 5026 9870
rect 5060 9836 5098 9870
rect 5132 9836 5170 9870
rect 5204 9836 5242 9870
rect 5276 9836 5314 9870
rect 5348 9836 5386 9870
rect 5420 9836 5458 9870
rect 5492 9836 5530 9870
rect 5564 9836 5602 9870
rect 5636 9836 5674 9870
rect 5708 9836 5746 9870
rect 5780 9836 5818 9870
rect 5852 9836 5890 9870
rect 5924 9836 5962 9870
rect 5996 9836 6034 9870
rect 6068 9836 6106 9870
rect 6140 9836 6178 9870
rect 6212 9836 6250 9870
rect 6284 9836 6322 9870
rect 6356 9836 6394 9870
rect 6428 9836 6466 9870
rect 6500 9836 6538 9870
rect 6572 9836 6610 9870
rect 6644 9836 6682 9870
rect 6716 9836 6754 9870
rect 6788 9836 6826 9870
rect 6860 9836 6898 9870
rect 6932 9836 6970 9870
rect 7004 9836 7042 9870
rect 7076 9836 7114 9870
rect 7148 9836 7186 9870
rect 7220 9836 7258 9870
rect 7292 9836 7330 9870
rect 7364 9836 7402 9870
rect 7436 9836 7474 9870
rect 7508 9836 7546 9870
rect 7580 9836 7618 9870
rect 7652 9836 7690 9870
rect 7724 9836 7762 9870
rect 7796 9836 7834 9870
rect 7868 9836 7906 9870
rect 7940 9836 7978 9870
rect 8012 9842 8050 9870
rect 8084 9842 8184 9876
rect 8218 9842 8224 9876
rect 8012 9836 8224 9842
rect 2270 9830 8224 9836
rect 8423 14530 8429 39330
rect 8535 27019 8573 39404
rect 8567 26967 8573 27019
rect 8535 26951 8573 26967
rect 8567 26899 8573 26951
rect 8535 14530 8573 26899
rect 8423 14491 8573 14530
rect 8423 14457 8429 14491
rect 8463 14457 8501 14491
rect 8535 14457 8573 14491
rect 8423 14418 8573 14457
rect 8423 14384 8429 14418
rect 8463 14384 8501 14418
rect 8535 14384 8573 14418
rect 8423 14345 8573 14384
rect 8423 14311 8429 14345
rect 8463 14311 8501 14345
rect 8535 14311 8573 14345
rect 8423 14272 8573 14311
rect 8423 14238 8429 14272
rect 8463 14238 8501 14272
rect 8535 14238 8573 14272
rect 8423 14199 8573 14238
rect 8423 14165 8429 14199
rect 8463 14165 8501 14199
rect 8535 14165 8573 14199
rect 8423 14126 8573 14165
rect 8423 14092 8429 14126
rect 8463 14092 8501 14126
rect 8535 14092 8573 14126
rect 8423 14053 8573 14092
rect 8423 14019 8429 14053
rect 8463 14019 8501 14053
rect 8535 14019 8573 14053
rect 8423 13980 8573 14019
rect 8423 13946 8429 13980
rect 8463 13946 8501 13980
rect 8535 13946 8573 13980
rect 8423 13907 8573 13946
rect 8423 13873 8429 13907
rect 8463 13873 8501 13907
rect 8535 13873 8573 13907
rect 8423 13834 8573 13873
rect 8423 13800 8429 13834
rect 8463 13800 8501 13834
rect 8535 13800 8573 13834
rect 8423 13761 8573 13800
rect 8423 13727 8429 13761
rect 8463 13727 8501 13761
rect 8535 13727 8573 13761
rect 8423 13688 8573 13727
rect 8423 13654 8429 13688
rect 8463 13654 8501 13688
rect 8535 13654 8573 13688
rect 8423 13615 8573 13654
rect 8423 13581 8429 13615
rect 8463 13581 8501 13615
rect 8535 13581 8573 13615
rect 8423 13542 8573 13581
rect 8423 13508 8429 13542
rect 8463 13508 8501 13542
rect 8535 13508 8573 13542
rect 8423 13469 8573 13508
rect 8423 13435 8429 13469
rect 8463 13435 8501 13469
rect 8535 13435 8573 13469
rect 8423 13396 8573 13435
rect 8423 13362 8429 13396
rect 8463 13362 8501 13396
rect 8535 13362 8573 13396
rect 8423 13323 8573 13362
rect 8423 13289 8429 13323
rect 8463 13289 8501 13323
rect 8535 13289 8573 13323
rect 8423 13250 8573 13289
rect 8423 13216 8429 13250
rect 8463 13216 8501 13250
rect 8535 13216 8573 13250
rect 8423 13177 8573 13216
rect 8423 13143 8429 13177
rect 8463 13143 8501 13177
rect 8535 13143 8573 13177
rect 8423 13104 8573 13143
rect 8423 13070 8429 13104
rect 8463 13070 8501 13104
rect 8535 13070 8573 13104
rect 8423 13031 8573 13070
rect 8423 12997 8429 13031
rect 8463 12997 8501 13031
rect 8535 12997 8573 13031
rect 8423 12958 8573 12997
rect 8423 12924 8429 12958
rect 8463 12924 8501 12958
rect 8535 12924 8573 12958
rect 8423 12885 8573 12924
rect 8423 12851 8429 12885
rect 8463 12851 8501 12885
rect 8535 12851 8573 12885
rect 8423 12812 8573 12851
rect 8423 12778 8429 12812
rect 8463 12778 8501 12812
rect 8535 12778 8573 12812
rect 8423 12739 8573 12778
rect 8423 12705 8429 12739
rect 8463 12705 8501 12739
rect 8535 12705 8573 12739
rect 8423 12666 8573 12705
rect 8423 12632 8429 12666
rect 8463 12632 8501 12666
rect 8535 12632 8573 12666
rect 8423 12593 8573 12632
rect 8423 12559 8429 12593
rect 8463 12559 8501 12593
rect 8535 12559 8573 12593
rect 8423 12520 8573 12559
rect 8423 12486 8429 12520
rect 8463 12486 8501 12520
rect 8535 12486 8573 12520
rect 8423 12447 8573 12486
rect 8423 12413 8429 12447
rect 8463 12413 8501 12447
rect 8535 12413 8573 12447
rect 8423 12374 8573 12413
rect 8423 12340 8429 12374
rect 8463 12340 8501 12374
rect 8535 12340 8573 12374
rect 8423 12301 8573 12340
rect 8423 12267 8429 12301
rect 8463 12267 8501 12301
rect 8535 12267 8573 12301
rect 8423 12228 8573 12267
rect 8423 12194 8429 12228
rect 8463 12194 8501 12228
rect 8535 12194 8573 12228
rect 8423 12155 8573 12194
rect 8423 12121 8429 12155
rect 8463 12121 8501 12155
rect 8535 12121 8573 12155
rect 8423 12082 8573 12121
rect 8423 12048 8429 12082
rect 8463 12048 8501 12082
rect 8535 12048 8573 12082
rect 8423 12009 8573 12048
rect 8423 11975 8429 12009
rect 8463 11975 8501 12009
rect 8535 11975 8573 12009
rect 8423 11936 8573 11975
rect 8423 11902 8429 11936
rect 8463 11902 8501 11936
rect 8535 11902 8573 11936
rect 8423 11863 8573 11902
rect 8423 11829 8429 11863
rect 8463 11829 8501 11863
rect 8535 11829 8573 11863
rect 8423 11790 8573 11829
rect 8423 11756 8429 11790
rect 8463 11756 8501 11790
rect 8535 11756 8573 11790
rect 8423 11717 8573 11756
rect 8423 11683 8429 11717
rect 8463 11683 8501 11717
rect 8535 11683 8573 11717
rect 8423 11644 8573 11683
rect 8423 11610 8429 11644
rect 8463 11610 8501 11644
rect 8535 11610 8573 11644
rect 8423 11571 8573 11610
rect 8423 11537 8429 11571
rect 8463 11537 8501 11571
rect 8535 11537 8573 11571
rect 8423 11498 8573 11537
rect 8423 11464 8429 11498
rect 8463 11464 8501 11498
rect 8535 11464 8573 11498
rect 8423 11425 8573 11464
rect 8423 11391 8429 11425
rect 8463 11391 8501 11425
rect 8535 11391 8573 11425
rect 8423 11352 8573 11391
rect 8423 11318 8429 11352
rect 8463 11318 8501 11352
rect 8535 11318 8573 11352
rect 8423 11279 8573 11318
rect 8423 11245 8429 11279
rect 8463 11245 8501 11279
rect 8535 11245 8573 11279
rect 8423 11206 8573 11245
rect 8423 11172 8429 11206
rect 8463 11172 8501 11206
rect 8535 11172 8573 11206
rect 8423 11133 8573 11172
rect 8423 11099 8429 11133
rect 8463 11099 8501 11133
rect 8535 11099 8573 11133
rect 8423 11060 8573 11099
rect 8423 11026 8429 11060
rect 8463 11026 8501 11060
rect 8535 11026 8573 11060
rect 8423 10987 8573 11026
rect 8423 10953 8429 10987
rect 8463 10953 8501 10987
rect 8535 10953 8573 10987
rect 8423 10914 8573 10953
rect 8423 10880 8429 10914
rect 8463 10880 8501 10914
rect 8535 10880 8573 10914
rect 8423 10841 8573 10880
rect 8423 10807 8429 10841
rect 8463 10807 8501 10841
rect 8535 10807 8573 10841
rect 8423 10768 8573 10807
rect 8423 10734 8429 10768
rect 8463 10734 8501 10768
rect 8535 10734 8573 10768
rect 8423 10695 8573 10734
rect 8423 10661 8429 10695
rect 8463 10661 8501 10695
rect 8535 10661 8573 10695
rect 8423 10622 8573 10661
rect 8423 10588 8429 10622
rect 8463 10588 8501 10622
rect 8535 10588 8573 10622
rect 8423 10549 8573 10588
rect 8423 10515 8429 10549
rect 8463 10515 8501 10549
rect 8535 10515 8573 10549
rect 8423 10476 8573 10515
rect 8423 10442 8429 10476
rect 8463 10442 8501 10476
rect 8535 10442 8573 10476
rect 8423 10403 8573 10442
rect 8423 10369 8429 10403
rect 8463 10369 8501 10403
rect 8535 10369 8573 10403
rect 8423 10330 8573 10369
rect 8423 10296 8429 10330
rect 8463 10296 8501 10330
rect 8535 10296 8573 10330
rect 8423 10257 8573 10296
rect 8423 10223 8429 10257
rect 8463 10223 8501 10257
rect 8535 10223 8573 10257
rect 8423 10184 8573 10223
rect 8423 10150 8429 10184
rect 8463 10150 8501 10184
rect 8535 10150 8573 10184
rect 8423 10111 8573 10150
rect 8423 10077 8429 10111
rect 8463 10077 8501 10111
rect 8535 10077 8573 10111
rect 8423 10038 8573 10077
rect 8423 10004 8429 10038
rect 8463 10004 8501 10038
rect 8535 10004 8573 10038
rect 8423 9965 8573 10004
rect 8423 9931 8429 9965
rect 8463 9931 8501 9965
rect 8535 9931 8573 9965
rect 8423 9892 8573 9931
rect 8423 9858 8429 9892
rect 8463 9858 8501 9892
rect 8535 9858 8573 9892
tri 8421 9819 8423 9821 se
rect 8423 9819 8573 9858
tri 8407 9805 8421 9819 se
rect 8421 9805 8429 9819
tri 2056 9785 2076 9805 sw
tri 8387 9785 8407 9805 se
rect 8407 9785 8429 9805
rect 8463 9785 8501 9819
rect 8535 9785 8573 9819
rect 2050 9752 2076 9785
tri 2076 9752 2109 9785 sw
tri 8354 9752 8387 9785 se
rect 8387 9752 8573 9785
rect 2050 9746 8573 9752
rect 2050 9712 7805 9746
rect 7839 9712 7883 9746
rect 7917 9712 7961 9746
rect 7995 9712 8039 9746
rect 8073 9712 8116 9746
rect 8150 9712 8193 9746
rect 8227 9712 8270 9746
rect 8304 9712 8347 9746
rect 8381 9712 8429 9746
rect 8463 9712 8501 9746
rect 8535 9712 8573 9746
rect 2050 9699 8573 9712
rect 2122 9665 2161 9699
rect 2195 9665 2234 9699
rect 2268 9665 2307 9699
rect 2341 9665 2380 9699
rect 2414 9665 2453 9699
rect 2487 9665 2526 9699
rect 2560 9665 2599 9699
rect 2633 9665 2672 9699
rect 2706 9665 2745 9699
rect 2779 9665 2818 9699
rect 2852 9665 2891 9699
rect 2925 9665 2964 9699
rect 2998 9665 3037 9699
rect 3071 9665 3110 9699
rect 3144 9665 3183 9699
rect 3217 9665 3256 9699
rect 3290 9665 3329 9699
rect 3363 9665 3402 9699
rect 3436 9665 3475 9699
rect 3509 9665 3548 9699
rect 3582 9665 3621 9699
rect 3655 9665 3694 9699
rect 3728 9665 3767 9699
rect 3801 9665 3840 9699
rect 3874 9665 3913 9699
rect 3947 9665 3986 9699
rect 4020 9665 4059 9699
rect 4093 9665 4132 9699
rect 4166 9665 4205 9699
rect 7695 9674 8573 9699
rect 2122 9627 4205 9665
rect 2122 9593 2161 9627
rect 2195 9593 2234 9627
rect 2268 9593 2307 9627
rect 2341 9593 2380 9627
rect 2414 9593 2453 9627
rect 2487 9593 2526 9627
rect 2560 9593 2599 9627
rect 2633 9593 2672 9627
rect 2706 9593 2745 9627
rect 2779 9593 2818 9627
rect 2852 9593 2891 9627
rect 2925 9593 2964 9627
rect 2998 9593 3037 9627
rect 3071 9593 3110 9627
rect 3144 9593 3183 9627
rect 3217 9593 3256 9627
rect 3290 9593 3329 9627
rect 3363 9593 3402 9627
rect 3436 9593 3475 9627
rect 3509 9593 3548 9627
rect 3582 9593 3621 9627
rect 3655 9593 3694 9627
rect 3728 9593 3767 9627
rect 3801 9593 3840 9627
rect 3874 9593 3913 9627
rect 3947 9593 3986 9627
rect 4020 9593 4059 9627
rect 4093 9593 4132 9627
rect 4166 9593 4205 9627
rect 7839 9640 7883 9674
rect 7917 9640 7961 9674
rect 7995 9640 8039 9674
rect 8073 9640 8116 9674
rect 8150 9640 8193 9674
rect 8227 9640 8270 9674
rect 8304 9640 8347 9674
rect 8381 9640 8424 9674
rect 8458 9640 8573 9674
rect 2050 9540 7733 9593
rect 2050 8938 2056 9540
tri 2056 9487 2109 9540 nw
tri 7694 9507 7727 9540 ne
tri 5195 9455 5198 9458 se
rect 5198 9455 5204 9458
rect 1938 8874 2056 8938
rect 1938 8840 1944 8874
rect 1978 8840 2016 8874
rect 2050 8840 2056 8874
rect 1938 8801 2056 8840
rect 1938 8767 1944 8801
rect 1978 8767 2016 8801
rect 2050 8767 2056 8801
rect 1938 8728 2056 8767
rect 1938 8694 1944 8728
rect 1978 8694 2016 8728
rect 2050 8694 2056 8728
rect 1938 8655 2056 8694
rect 1938 8621 1944 8655
rect 1978 8621 2016 8655
rect 2050 8621 2056 8655
rect 1938 8582 2056 8621
rect 1938 8548 1944 8582
rect 1978 8548 2016 8582
rect 2050 8548 2056 8582
rect 1938 8509 2056 8548
rect 1938 8475 1944 8509
rect 1978 8475 2016 8509
rect 2050 8475 2056 8509
rect 1938 8436 2056 8475
rect 1938 8402 1944 8436
rect 1978 8402 2016 8436
rect 2050 8402 2056 8436
rect 1938 8363 2056 8402
rect 1938 8329 1944 8363
rect 1978 8329 2016 8363
rect 2050 8329 2056 8363
rect 1938 8290 2056 8329
rect 1938 8256 1944 8290
rect 1978 8256 2016 8290
rect 2050 8256 2056 8290
rect 1938 8217 2056 8256
rect 1938 8183 1944 8217
rect 1978 8183 2016 8217
rect 2050 8183 2056 8217
rect 1938 8144 2056 8183
rect 1938 8110 1944 8144
rect 1978 8110 2016 8144
rect 2050 8110 2056 8144
rect 1938 8071 2056 8110
rect 1938 8037 1944 8071
rect 1978 8037 2016 8071
rect 2050 8037 2056 8071
rect 1938 7998 2056 8037
rect 1938 7964 1944 7998
rect 1978 7964 2016 7998
rect 2050 7964 2056 7998
rect 1938 7925 2056 7964
rect 1938 7891 1944 7925
rect 1978 7891 2016 7925
rect 2050 7891 2056 7925
rect 1938 7852 2056 7891
rect 1938 7818 1944 7852
rect 1978 7818 2016 7852
rect 2050 7818 2056 7852
rect 1938 7779 2056 7818
rect 1938 7745 1944 7779
rect 1978 7745 2016 7779
rect 2050 7745 2056 7779
rect 1938 7706 2056 7745
rect 1938 7672 1944 7706
rect 1978 7672 2016 7706
rect 2050 7672 2056 7706
rect 1938 7633 2056 7672
rect 1938 7599 1944 7633
rect 1978 7599 2016 7633
rect 2050 7599 2056 7633
rect 1938 7560 2056 7599
rect 1938 7526 1944 7560
rect 1978 7526 2016 7560
rect 2050 7526 2056 7560
rect 1938 7487 2056 7526
rect 1938 7453 1944 7487
rect 1978 7453 2016 7487
rect 2050 7453 2056 7487
rect 1938 7414 2056 7453
rect 1938 7380 1944 7414
rect 1978 7380 2016 7414
rect 2050 7380 2056 7414
rect 1938 7341 2056 7380
rect 1938 3491 1944 7341
rect 2050 3491 2056 7341
rect 2135 9449 5204 9455
rect 2135 9443 2359 9449
rect 2135 5305 2141 9443
rect 2319 9415 2359 9443
rect 2393 9415 2432 9449
rect 2466 9415 2505 9449
rect 2539 9415 2578 9449
rect 2612 9415 2651 9449
rect 2685 9415 2724 9449
rect 2758 9415 2797 9449
rect 2831 9415 2870 9449
rect 2904 9415 2943 9449
rect 2977 9415 3016 9449
rect 3050 9415 3089 9449
rect 3123 9415 3162 9449
rect 3196 9415 3235 9449
rect 3269 9415 3308 9449
rect 3342 9415 3381 9449
rect 3415 9415 3454 9449
rect 3488 9415 3527 9449
rect 3561 9415 3600 9449
rect 3634 9415 3673 9449
rect 3707 9415 3746 9449
rect 3780 9415 3819 9449
rect 3853 9415 3892 9449
rect 3926 9415 3965 9449
rect 3999 9415 4038 9449
rect 4072 9415 4111 9449
rect 4145 9415 4184 9449
rect 4218 9415 4257 9449
rect 4291 9415 4330 9449
rect 4364 9415 4403 9449
rect 4437 9415 4476 9449
rect 4510 9415 4549 9449
rect 4583 9415 4622 9449
rect 4656 9415 4694 9449
rect 4728 9415 4766 9449
rect 4800 9415 4838 9449
rect 4872 9415 4910 9449
rect 4944 9415 4982 9449
rect 5016 9415 5054 9449
rect 5088 9415 5126 9449
rect 5160 9415 5198 9449
rect 2319 9409 5204 9415
rect 2319 9403 2349 9409
tri 2349 9403 2355 9409 nw
tri 5195 9406 5198 9409 ne
rect 5198 9406 5204 9409
rect 5256 9406 5268 9458
rect 5320 9406 5332 9458
rect 5384 9406 5396 9458
rect 5448 9406 5460 9458
rect 5512 9449 5524 9458
rect 5576 9449 5588 9458
rect 5640 9449 5652 9458
rect 5704 9449 5716 9458
rect 5768 9449 5780 9458
rect 5520 9415 5524 9449
rect 5768 9415 5774 9449
rect 5512 9406 5524 9415
rect 5576 9406 5588 9415
rect 5640 9406 5652 9415
rect 5704 9406 5716 9415
rect 5768 9406 5780 9415
rect 5832 9406 5844 9458
rect 5896 9406 5908 9458
rect 5960 9406 5972 9458
rect 6024 9406 6036 9458
rect 6088 9449 6100 9458
rect 6152 9449 6164 9458
rect 6216 9449 6228 9458
rect 6280 9449 6292 9458
rect 6344 9449 6356 9458
rect 6096 9415 6100 9449
rect 6344 9415 6350 9449
rect 6088 9406 6100 9415
rect 6152 9406 6164 9415
rect 6216 9406 6228 9415
rect 6280 9406 6292 9415
rect 6344 9406 6356 9415
rect 6408 9406 6420 9458
rect 6472 9406 6484 9458
rect 6536 9406 6548 9458
rect 6600 9406 6612 9458
rect 6664 9449 6676 9458
rect 6728 9449 6740 9458
rect 6792 9449 6804 9458
rect 6856 9449 6868 9458
rect 6920 9449 6932 9458
rect 6672 9415 6676 9449
rect 6920 9415 6926 9449
rect 6664 9406 6676 9415
rect 6728 9406 6740 9415
rect 6792 9406 6804 9415
rect 6856 9406 6868 9415
rect 6920 9406 6932 9415
rect 6984 9406 6996 9458
rect 7048 9406 7060 9458
rect 7112 9406 7124 9458
rect 7176 9406 7188 9458
rect 7240 9449 7252 9458
rect 7304 9449 7316 9458
rect 7368 9455 7374 9458
tri 7374 9455 7377 9458 sw
rect 7368 9449 7619 9455
rect 7248 9415 7252 9449
rect 7392 9437 7619 9449
rect 7392 9415 7493 9437
rect 7240 9406 7252 9415
rect 7304 9406 7316 9415
rect 7368 9409 7493 9415
rect 7368 9406 7374 9409
tri 7374 9406 7377 9409 nw
tri 7415 9406 7418 9409 ne
rect 7418 9406 7493 9409
tri 7418 9403 7421 9406 ne
rect 7421 9403 7493 9406
rect 7527 9403 7579 9437
rect 7613 9403 7619 9437
rect 2319 7709 2325 9403
tri 2325 9379 2349 9403 nw
tri 7421 9379 7445 9403 ne
rect 7445 9379 7619 9403
tri 7445 9365 7459 9379 ne
rect 7459 9365 7619 9379
tri 7459 9350 7474 9365 ne
rect 7474 9350 7493 9365
rect 2468 9298 2474 9350
rect 2526 9298 2539 9350
rect 2591 9298 2604 9350
rect 2656 9341 7380 9350
rect 2660 9307 2699 9341
rect 2733 9307 2772 9341
rect 2806 9307 2845 9341
rect 2879 9307 2918 9341
rect 2952 9307 2991 9341
rect 3025 9307 3064 9341
rect 3098 9307 3137 9341
rect 3171 9307 3210 9341
rect 3244 9307 3283 9341
rect 3317 9307 3356 9341
rect 3390 9307 3429 9341
rect 3463 9307 3502 9341
rect 3536 9307 3575 9341
rect 3609 9307 3648 9341
rect 3682 9307 3721 9341
rect 3755 9307 3794 9341
rect 3828 9307 3867 9341
rect 3901 9307 3940 9341
rect 3974 9307 4013 9341
rect 4047 9307 4086 9341
rect 4120 9307 4159 9341
rect 4193 9307 4232 9341
rect 4266 9307 4305 9341
rect 4339 9307 4378 9341
rect 4412 9307 4451 9341
rect 4485 9307 4524 9341
rect 4558 9307 4597 9341
rect 4631 9307 4670 9341
rect 4704 9307 4742 9341
rect 4776 9307 4814 9341
rect 4848 9307 4886 9341
rect 4920 9307 4958 9341
rect 4992 9307 5030 9341
rect 5064 9307 5102 9341
rect 5136 9307 5174 9341
rect 5208 9307 5246 9341
rect 5280 9307 5318 9341
rect 5352 9307 5390 9341
rect 5424 9307 5462 9341
rect 5496 9307 5534 9341
rect 5568 9307 5606 9341
rect 5640 9307 5678 9341
rect 5712 9307 5750 9341
rect 5784 9307 5822 9341
rect 5856 9307 5894 9341
rect 5928 9307 5966 9341
rect 6000 9307 6038 9341
rect 6072 9307 6110 9341
rect 6144 9307 6182 9341
rect 6216 9307 6254 9341
rect 6288 9307 6326 9341
rect 6360 9307 6398 9341
rect 6432 9307 6470 9341
rect 6504 9307 6542 9341
rect 6576 9307 6614 9341
rect 6648 9307 6686 9341
rect 6720 9307 6758 9341
rect 6792 9307 6830 9341
rect 6864 9307 6902 9341
rect 6936 9307 6974 9341
rect 7008 9307 7046 9341
rect 7080 9307 7118 9341
rect 7152 9307 7190 9341
rect 7224 9307 7262 9341
rect 7296 9307 7334 9341
rect 7368 9307 7380 9341
tri 7474 9337 7487 9350 ne
rect 2656 9298 7380 9307
rect 7487 9331 7493 9350
rect 7527 9331 7579 9365
rect 7613 9331 7619 9365
rect 7487 9293 7619 9331
rect 7487 9259 7493 9293
rect 7527 9259 7579 9293
rect 7613 9259 7619 9293
rect 2411 9212 2467 9224
rect 2411 9178 2422 9212
rect 2456 9178 2467 9212
rect 2411 9139 2467 9178
rect 2411 9105 2422 9139
rect 2456 9105 2467 9139
rect 2411 9066 2467 9105
rect 2411 9032 2422 9066
rect 2456 9032 2467 9066
rect 2411 8993 2467 9032
rect 2411 8959 2422 8993
rect 2456 8959 2467 8993
rect 2411 8920 2467 8959
rect 2411 8886 2422 8920
rect 2456 8886 2467 8920
rect 2411 8847 2467 8886
rect 2411 8813 2422 8847
rect 2456 8813 2467 8847
rect 2411 8774 2467 8813
rect 2411 8740 2422 8774
rect 2456 8740 2467 8774
rect 4068 9212 4124 9224
rect 4068 9178 4079 9212
rect 4113 9178 4124 9212
rect 4068 9139 4124 9178
rect 4068 9105 4079 9139
rect 4113 9105 4124 9139
rect 4068 9066 4124 9105
rect 4068 9032 4079 9066
rect 4113 9032 4124 9066
rect 4068 8993 4124 9032
rect 4068 8959 4079 8993
rect 4113 8959 4124 8993
rect 4068 8920 4124 8959
rect 4068 8886 4079 8920
rect 4113 8886 4124 8920
rect 4068 8847 4124 8886
rect 4068 8813 4079 8847
rect 4113 8813 4124 8847
rect 4068 8774 4124 8813
tri 4067 8757 4068 8758 se
rect 4068 8757 4079 8774
tri 2467 8740 2484 8757 sw
tri 4050 8740 4067 8757 se
rect 4067 8740 4079 8757
rect 4113 8740 4124 8774
rect 5726 9212 5782 9224
rect 5726 9178 5737 9212
rect 5771 9178 5782 9212
rect 5726 9139 5782 9178
rect 5726 9105 5737 9139
rect 5771 9105 5782 9139
rect 5726 9066 5782 9105
rect 5726 9032 5737 9066
rect 5771 9032 5782 9066
rect 5726 8993 5782 9032
rect 5726 8959 5737 8993
rect 5771 8959 5782 8993
rect 5726 8920 5782 8959
rect 5726 8886 5737 8920
rect 5771 8886 5782 8920
rect 5726 8847 5782 8886
rect 5726 8813 5737 8847
rect 5771 8813 5782 8847
rect 5726 8774 5782 8813
tri 4124 8740 4142 8758 sw
tri 5708 8740 5726 8758 se
rect 5726 8740 5737 8774
rect 5771 8740 5782 8774
rect 7375 9212 7431 9224
rect 7375 9178 7386 9212
rect 7420 9178 7431 9212
rect 7375 9139 7431 9178
rect 7375 9105 7386 9139
rect 7420 9105 7431 9139
rect 7375 9066 7431 9105
rect 7375 9032 7386 9066
rect 7420 9032 7431 9066
rect 7375 8993 7431 9032
rect 7375 8959 7386 8993
rect 7420 8959 7431 8993
rect 7375 8920 7431 8959
rect 7375 8886 7386 8920
rect 7420 8886 7431 8920
rect 7375 8847 7431 8886
rect 7375 8813 7386 8847
rect 7420 8813 7431 8847
rect 7375 8774 7431 8813
tri 5782 8740 5800 8758 sw
tri 7357 8740 7375 8758 se
rect 7375 8740 7386 8774
rect 7420 8740 7431 8774
rect 2411 8729 2484 8740
tri 2484 8729 2495 8740 sw
tri 4039 8729 4050 8740 se
rect 4050 8729 4142 8740
tri 4142 8729 4153 8740 sw
tri 5697 8729 5708 8740 se
rect 5708 8729 5800 8740
tri 5800 8729 5811 8740 sw
tri 7346 8729 7357 8740 se
rect 7357 8729 7431 8740
rect 2411 8727 7431 8729
rect 2411 8701 5204 8727
rect 7368 8701 7431 8727
rect 2411 8667 2422 8701
rect 2456 8667 4079 8701
rect 4113 8667 5204 8701
rect 7368 8667 7386 8701
rect 7420 8667 7431 8701
rect 2411 8628 5204 8667
rect 7368 8628 7431 8667
rect 2411 8594 2422 8628
rect 2456 8594 4079 8628
rect 4113 8594 5204 8628
rect 7368 8594 7386 8628
rect 7420 8594 7431 8628
rect 2411 8554 5204 8594
rect 7368 8554 7431 8594
rect 2411 8520 2422 8554
rect 2456 8520 4079 8554
rect 4113 8520 5204 8554
rect 7368 8520 7386 8554
rect 7420 8520 7431 8554
rect 2411 8480 5204 8520
rect 7368 8480 7431 8520
rect 2411 8446 2422 8480
rect 2456 8446 4079 8480
rect 4113 8446 5204 8480
rect 7368 8446 7386 8480
rect 7420 8446 7431 8480
rect 2411 8406 5204 8446
rect 7368 8406 7431 8446
rect 2411 8372 2422 8406
rect 2456 8372 4079 8406
rect 4113 8372 5204 8406
rect 7368 8372 7386 8406
rect 7420 8372 7431 8406
rect 2411 8332 5204 8372
rect 7368 8332 7431 8372
rect 2411 8298 2422 8332
rect 2456 8298 4079 8332
rect 4113 8298 5204 8332
rect 7368 8298 7386 8332
rect 7420 8298 7431 8332
rect 2411 8258 5204 8298
rect 7368 8258 7431 8298
rect 2411 8224 2422 8258
rect 2456 8224 4079 8258
rect 4113 8224 5204 8258
rect 7368 8224 7386 8258
rect 7420 8224 7431 8258
rect 2411 8184 5204 8224
rect 7368 8184 7431 8224
rect 2411 8150 2422 8184
rect 2456 8150 4079 8184
rect 4113 8150 5204 8184
rect 7368 8150 7386 8184
rect 7420 8150 7431 8184
rect 2411 8110 5204 8150
rect 7368 8110 7431 8150
rect 2411 8076 2422 8110
rect 2456 8076 4079 8110
rect 4113 8076 5204 8110
rect 7368 8076 7386 8110
rect 7420 8076 7431 8110
rect 2411 8036 5204 8076
rect 7368 8036 7431 8076
rect 2411 8002 2422 8036
rect 2456 8002 4079 8036
rect 4113 8002 5204 8036
rect 7368 8002 7386 8036
rect 7420 8002 7431 8036
rect 2411 7962 5204 8002
rect 7368 7962 7431 8002
rect 2411 7928 2422 7962
rect 2456 7928 4079 7962
rect 4113 7928 5204 7962
rect 7368 7928 7386 7962
rect 7420 7928 7431 7962
rect 2411 7888 5204 7928
rect 7368 7888 7431 7928
rect 2411 7854 2422 7888
rect 2456 7854 4079 7888
rect 4113 7854 5204 7888
rect 7368 7854 7386 7888
rect 7420 7854 7431 7888
rect 2411 7843 5204 7854
rect 7368 7843 7431 7854
rect 2411 7842 7431 7843
rect 7487 9221 7619 9259
rect 7487 9187 7493 9221
rect 7527 9187 7579 9221
rect 7613 9187 7619 9221
rect 7487 9149 7619 9187
rect 7487 9115 7493 9149
rect 7527 9115 7579 9149
rect 7613 9115 7619 9149
rect 7487 9077 7619 9115
rect 7487 9043 7493 9077
rect 7527 9043 7579 9077
rect 7613 9043 7619 9077
rect 7487 9005 7619 9043
rect 7487 8971 7493 9005
rect 7527 8971 7579 9005
rect 7613 8971 7619 9005
rect 7487 8933 7619 8971
rect 7487 8899 7493 8933
rect 7527 8899 7579 8933
rect 7613 8899 7619 8933
rect 7487 8861 7619 8899
rect 7487 8827 7493 8861
rect 7527 8827 7579 8861
rect 7613 8827 7619 8861
rect 7487 8789 7619 8827
rect 7487 8755 7493 8789
rect 7527 8755 7579 8789
rect 7613 8755 7619 8789
rect 7487 8717 7619 8755
rect 7487 8683 7493 8717
rect 7527 8683 7579 8717
rect 7613 8683 7619 8717
rect 7487 8645 7619 8683
rect 7487 8611 7493 8645
rect 7527 8611 7579 8645
rect 7613 8611 7619 8645
rect 7487 8573 7619 8611
rect 7487 8539 7493 8573
rect 7527 8539 7579 8573
rect 7613 8539 7619 8573
rect 7487 8501 7619 8539
rect 7487 8467 7493 8501
rect 7527 8467 7579 8501
rect 7613 8467 7619 8501
rect 7487 8429 7619 8467
rect 7487 8395 7493 8429
rect 7527 8395 7579 8429
rect 7613 8395 7619 8429
rect 7487 8357 7619 8395
rect 7487 8323 7493 8357
rect 7527 8323 7579 8357
rect 7613 8323 7619 8357
rect 7487 8285 7619 8323
rect 7487 8251 7493 8285
rect 7527 8251 7579 8285
rect 7613 8251 7619 8285
rect 7487 8213 7619 8251
rect 7487 8179 7493 8213
rect 7527 8179 7579 8213
rect 7613 8179 7619 8213
rect 7487 8141 7619 8179
rect 7487 8107 7493 8141
rect 7527 8107 7579 8141
rect 7613 8107 7619 8141
rect 7487 8069 7619 8107
rect 7487 8035 7493 8069
rect 7527 8035 7579 8069
rect 7613 8035 7619 8069
rect 7487 7997 7619 8035
rect 7487 7963 7493 7997
rect 7527 7963 7579 7997
rect 7613 7963 7619 7997
rect 7487 7925 7619 7963
rect 7487 7891 7493 7925
rect 7527 7891 7579 7925
rect 7613 7891 7619 7925
rect 7487 7853 7619 7891
rect 7487 7819 7493 7853
rect 7527 7819 7579 7853
rect 7613 7819 7619 7853
rect 7487 7781 7619 7819
rect 7487 7747 7493 7781
rect 7527 7747 7579 7781
rect 7613 7747 7619 7781
tri 2325 7709 2337 7721 sw
tri 7475 7709 7487 7721 se
rect 7487 7709 7619 7747
rect 2319 7687 2337 7709
tri 2337 7687 2359 7709 sw
tri 7456 7690 7475 7709 se
rect 7475 7690 7493 7709
tri 5195 7687 5198 7690 se
rect 5198 7687 5204 7690
rect 2319 7681 5204 7687
rect 5256 7681 5268 7690
rect 5320 7681 5332 7690
rect 5384 7681 5396 7690
rect 5448 7681 5460 7690
rect 2319 7647 2357 7681
rect 2391 7647 2429 7681
rect 2463 7647 2501 7681
rect 2535 7647 2573 7681
rect 2607 7647 2645 7681
rect 2679 7647 2717 7681
rect 2751 7647 2789 7681
rect 2823 7647 2861 7681
rect 2895 7647 2933 7681
rect 2967 7647 3005 7681
rect 3039 7647 3077 7681
rect 3111 7647 3149 7681
rect 3183 7647 3221 7681
rect 3255 7647 3293 7681
rect 3327 7647 3365 7681
rect 3399 7647 3437 7681
rect 3471 7647 3509 7681
rect 3543 7647 3581 7681
rect 3615 7647 3653 7681
rect 3687 7647 3725 7681
rect 3759 7647 3797 7681
rect 3831 7647 3869 7681
rect 3903 7647 3941 7681
rect 3975 7647 4013 7681
rect 4047 7647 4085 7681
rect 4119 7647 4157 7681
rect 4191 7647 4229 7681
rect 4263 7647 4301 7681
rect 4335 7647 4373 7681
rect 4407 7647 4445 7681
rect 4479 7647 4517 7681
rect 4551 7647 4589 7681
rect 4623 7647 4661 7681
rect 4695 7647 4733 7681
rect 4767 7647 4805 7681
rect 4839 7647 4877 7681
rect 4911 7647 4949 7681
rect 4983 7647 5021 7681
rect 5055 7647 5093 7681
rect 5127 7647 5165 7681
rect 5199 7647 5204 7681
rect 5448 7647 5453 7681
rect 2319 7641 5204 7647
rect 2319 7637 2355 7641
tri 2355 7637 2359 7641 nw
tri 5195 7638 5198 7641 ne
rect 5198 7638 5204 7641
rect 5256 7638 5268 7647
rect 5320 7638 5332 7647
rect 5384 7638 5396 7647
rect 5448 7638 5460 7647
rect 5512 7638 5524 7690
rect 5576 7638 5588 7690
rect 5640 7638 5652 7690
rect 5704 7638 5716 7690
rect 5768 7681 5780 7690
rect 5832 7681 5844 7690
rect 5896 7681 5908 7690
rect 5960 7681 5972 7690
rect 6024 7681 6036 7690
rect 5775 7647 5780 7681
rect 6024 7647 6029 7681
rect 5768 7638 5780 7647
rect 5832 7638 5844 7647
rect 5896 7638 5908 7647
rect 5960 7638 5972 7647
rect 6024 7638 6036 7647
rect 6088 7638 6100 7690
rect 6152 7638 6164 7690
rect 6216 7638 6228 7690
rect 6280 7638 6292 7690
rect 6344 7681 6356 7690
rect 6408 7681 6420 7690
rect 6472 7681 6484 7690
rect 6536 7681 6548 7690
rect 6600 7681 6612 7690
rect 6351 7647 6356 7681
rect 6600 7647 6605 7681
rect 6344 7638 6356 7647
rect 6408 7638 6420 7647
rect 6472 7638 6484 7647
rect 6536 7638 6548 7647
rect 6600 7638 6612 7647
rect 6664 7638 6676 7690
rect 6728 7638 6740 7690
rect 6792 7638 6804 7690
rect 6856 7638 6868 7690
rect 6920 7681 6932 7690
rect 6984 7681 6996 7690
rect 7048 7681 7060 7690
rect 7112 7681 7124 7690
rect 7176 7681 7188 7690
rect 6927 7647 6932 7681
rect 7176 7647 7181 7681
rect 6920 7638 6932 7647
rect 6984 7638 6996 7647
rect 7048 7638 7060 7647
rect 7112 7638 7124 7647
rect 7176 7638 7188 7647
rect 7240 7638 7252 7690
rect 7304 7638 7316 7690
rect 7368 7687 7374 7690
tri 7374 7687 7377 7690 sw
tri 7453 7687 7456 7690 se
rect 7456 7687 7493 7690
rect 7368 7681 7493 7687
rect 7368 7647 7397 7681
rect 7431 7675 7493 7681
rect 7527 7675 7579 7709
rect 7613 7675 7619 7709
rect 7431 7647 7619 7675
rect 7368 7641 7619 7647
rect 7368 7638 7374 7641
tri 7374 7638 7377 7641 nw
tri 7453 7638 7456 7641 ne
rect 7456 7638 7619 7641
tri 7456 7637 7457 7638 ne
rect 7457 7637 7619 7638
rect 2319 5875 2325 7637
tri 2325 7607 2355 7637 nw
tri 7457 7607 7487 7637 ne
rect 7487 7603 7493 7637
rect 7527 7603 7579 7637
rect 7613 7603 7619 7637
rect 7487 7565 7619 7603
rect 2468 7497 2474 7549
rect 2526 7497 2539 7549
rect 2591 7497 2604 7549
rect 2656 7540 7380 7549
rect 2660 7506 2699 7540
rect 2733 7506 2772 7540
rect 2806 7506 2845 7540
rect 2879 7506 2918 7540
rect 2952 7506 2991 7540
rect 3025 7506 3064 7540
rect 3098 7506 3137 7540
rect 3171 7506 3210 7540
rect 3244 7506 3283 7540
rect 3317 7506 3356 7540
rect 3390 7506 3429 7540
rect 3463 7506 3502 7540
rect 3536 7506 3575 7540
rect 3609 7506 3648 7540
rect 3682 7506 3721 7540
rect 3755 7506 3794 7540
rect 3828 7506 3867 7540
rect 3901 7506 3940 7540
rect 3974 7506 4013 7540
rect 4047 7506 4086 7540
rect 4120 7506 4159 7540
rect 4193 7506 4232 7540
rect 4266 7506 4305 7540
rect 4339 7506 4378 7540
rect 4412 7506 4451 7540
rect 4485 7506 4524 7540
rect 4558 7506 4597 7540
rect 4631 7506 4670 7540
rect 4704 7506 4742 7540
rect 4776 7506 4814 7540
rect 4848 7506 4886 7540
rect 4920 7506 4958 7540
rect 4992 7506 5030 7540
rect 5064 7506 5102 7540
rect 5136 7506 5174 7540
rect 5208 7506 5246 7540
rect 5280 7506 5318 7540
rect 5352 7506 5390 7540
rect 5424 7506 5462 7540
rect 5496 7506 5534 7540
rect 5568 7506 5606 7540
rect 5640 7506 5678 7540
rect 5712 7506 5750 7540
rect 5784 7506 5822 7540
rect 5856 7506 5894 7540
rect 5928 7506 5966 7540
rect 6000 7506 6038 7540
rect 6072 7506 6110 7540
rect 6144 7506 6182 7540
rect 6216 7506 6254 7540
rect 6288 7506 6326 7540
rect 6360 7506 6398 7540
rect 6432 7506 6470 7540
rect 6504 7506 6542 7540
rect 6576 7506 6614 7540
rect 6648 7506 6686 7540
rect 6720 7506 6758 7540
rect 6792 7506 6830 7540
rect 6864 7506 6902 7540
rect 6936 7506 6974 7540
rect 7008 7506 7046 7540
rect 7080 7506 7118 7540
rect 7152 7506 7190 7540
rect 7224 7506 7262 7540
rect 7296 7506 7334 7540
rect 7368 7506 7380 7540
rect 2656 7497 7380 7506
rect 7487 7531 7493 7565
rect 7527 7531 7579 7565
rect 7613 7531 7619 7565
rect 7487 7493 7619 7531
rect 7487 7459 7493 7493
rect 7527 7459 7579 7493
rect 7613 7459 7619 7493
rect 2411 7412 2467 7424
rect 2411 7378 2422 7412
rect 2456 7378 2467 7412
rect 2411 7339 2467 7378
rect 2411 7305 2422 7339
rect 2456 7305 2467 7339
rect 2411 7266 2467 7305
rect 2411 7232 2422 7266
rect 2456 7232 2467 7266
rect 2411 7193 2467 7232
rect 2411 7159 2422 7193
rect 2456 7159 2467 7193
rect 2411 7120 2467 7159
rect 2411 7086 2422 7120
rect 2456 7086 2467 7120
rect 2411 7047 2467 7086
rect 2411 7013 2422 7047
rect 2456 7013 2467 7047
rect 2411 6974 2467 7013
rect 2411 6940 2422 6974
rect 2456 6940 2467 6974
rect 4068 7412 4124 7424
rect 4068 7378 4079 7412
rect 4113 7378 4124 7412
rect 4068 7339 4124 7378
rect 4068 7305 4079 7339
rect 4113 7305 4124 7339
rect 4068 7266 4124 7305
rect 4068 7232 4079 7266
rect 4113 7232 4124 7266
rect 4068 7193 4124 7232
rect 4068 7159 4079 7193
rect 4113 7159 4124 7193
rect 4068 7120 4124 7159
rect 4068 7086 4079 7120
rect 4113 7086 4124 7120
rect 4068 7047 4124 7086
rect 4068 7013 4079 7047
rect 4113 7013 4124 7047
rect 4068 6974 4124 7013
tri 2467 6940 2492 6965 sw
tri 4050 6940 4068 6958 se
rect 4068 6940 4079 6974
rect 4113 6940 4124 6974
rect 5726 7412 5782 7424
rect 5726 7378 5737 7412
rect 5771 7378 5782 7412
rect 5726 7339 5782 7378
rect 5726 7305 5737 7339
rect 5771 7305 5782 7339
rect 5726 7266 5782 7305
rect 5726 7232 5737 7266
rect 5771 7232 5782 7266
rect 5726 7193 5782 7232
rect 5726 7159 5737 7193
rect 5771 7159 5782 7193
rect 5726 7120 5782 7159
rect 5726 7086 5737 7120
rect 5771 7086 5782 7120
rect 5726 7047 5782 7086
rect 5726 7013 5737 7047
rect 5771 7013 5782 7047
rect 5726 6974 5782 7013
tri 4124 6940 4142 6958 sw
tri 5708 6940 5726 6958 se
rect 5726 6940 5737 6974
rect 5771 6940 5782 6974
rect 7375 7412 7431 7424
rect 7375 7378 7386 7412
rect 7420 7378 7431 7412
rect 7375 7339 7431 7378
rect 7375 7305 7386 7339
rect 7420 7305 7431 7339
rect 7375 7266 7431 7305
rect 7375 7232 7386 7266
rect 7420 7232 7431 7266
rect 7375 7193 7431 7232
rect 7375 7159 7386 7193
rect 7420 7159 7431 7193
rect 7375 7120 7431 7159
rect 7375 7086 7386 7120
rect 7420 7086 7431 7120
rect 7375 7047 7431 7086
rect 7375 7013 7386 7047
rect 7420 7013 7431 7047
rect 7375 6974 7431 7013
tri 7367 6958 7375 6966 se
rect 7375 6958 7386 6974
tri 5782 6940 5800 6958 sw
tri 7349 6940 7367 6958 se
rect 7367 6940 7386 6958
rect 7420 6940 7431 6974
rect 2411 6929 2492 6940
tri 2492 6929 2503 6940 sw
tri 4039 6929 4050 6940 se
rect 4050 6929 4142 6940
tri 4142 6929 4153 6940 sw
tri 5697 6929 5708 6940 se
rect 5708 6929 5800 6940
tri 5800 6929 5811 6940 sw
tri 7338 6929 7349 6940 se
rect 7349 6929 7431 6940
rect 2411 6927 7431 6929
rect 2411 6901 5204 6927
rect 7368 6901 7431 6927
rect 2411 6867 2422 6901
rect 2456 6867 4079 6901
rect 4113 6867 5204 6901
rect 7368 6867 7386 6901
rect 7420 6867 7431 6901
rect 2411 6828 5204 6867
rect 7368 6828 7431 6867
rect 2411 6794 2422 6828
rect 2456 6794 4079 6828
rect 4113 6794 5204 6828
rect 7368 6794 7386 6828
rect 7420 6794 7431 6828
rect 2411 6754 5204 6794
rect 7368 6754 7431 6794
rect 2411 6720 2422 6754
rect 2456 6720 4079 6754
rect 4113 6720 5204 6754
rect 7368 6720 7386 6754
rect 7420 6720 7431 6754
rect 2411 6680 5204 6720
rect 7368 6680 7431 6720
rect 2411 6646 2422 6680
rect 2456 6646 4079 6680
rect 4113 6646 5204 6680
rect 7368 6646 7386 6680
rect 7420 6646 7431 6680
rect 2411 6606 5204 6646
rect 7368 6606 7431 6646
rect 2411 6572 2422 6606
rect 2456 6572 4079 6606
rect 4113 6572 5204 6606
rect 7368 6572 7386 6606
rect 7420 6572 7431 6606
rect 2411 6532 5204 6572
rect 7368 6532 7431 6572
rect 2411 6498 2422 6532
rect 2456 6498 4079 6532
rect 4113 6498 5204 6532
rect 7368 6498 7386 6532
rect 7420 6498 7431 6532
rect 2411 6458 5204 6498
rect 7368 6458 7431 6498
rect 2411 6424 2422 6458
rect 2456 6424 4079 6458
rect 4113 6424 5204 6458
rect 7368 6424 7386 6458
rect 7420 6424 7431 6458
rect 2411 6384 5204 6424
rect 7368 6384 7431 6424
rect 2411 6350 2422 6384
rect 2456 6350 4079 6384
rect 4113 6350 5204 6384
rect 7368 6350 7386 6384
rect 7420 6350 7431 6384
rect 2411 6310 5204 6350
rect 7368 6310 7431 6350
rect 2411 6276 2422 6310
rect 2456 6276 4079 6310
rect 4113 6276 5204 6310
rect 7368 6276 7386 6310
rect 7420 6276 7431 6310
rect 2411 6236 5204 6276
rect 7368 6236 7431 6276
rect 2411 6202 2422 6236
rect 2456 6202 4079 6236
rect 4113 6202 5204 6236
rect 7368 6202 7386 6236
rect 7420 6202 7431 6236
rect 2411 6162 5204 6202
rect 7368 6162 7431 6202
rect 2411 6128 2422 6162
rect 2456 6128 4079 6162
rect 4113 6128 5204 6162
rect 7368 6128 7386 6162
rect 7420 6128 7431 6162
rect 2411 6088 5204 6128
rect 7368 6088 7431 6128
rect 2411 6054 2422 6088
rect 2456 6054 4079 6088
rect 4113 6054 5204 6088
rect 7368 6054 7386 6088
rect 7420 6054 7431 6088
rect 2411 6043 5204 6054
rect 7368 6043 7431 6054
rect 2411 6042 7431 6043
rect 7487 7421 7619 7459
rect 7487 7387 7493 7421
rect 7527 7387 7579 7421
rect 7613 7387 7619 7421
rect 7487 7349 7619 7387
rect 7487 7315 7493 7349
rect 7527 7315 7579 7349
rect 7613 7315 7619 7349
rect 7487 7277 7619 7315
rect 7487 7243 7493 7277
rect 7527 7243 7579 7277
rect 7613 7243 7619 7277
rect 7487 7205 7619 7243
rect 7487 7171 7493 7205
rect 7527 7171 7579 7205
rect 7613 7171 7619 7205
rect 7487 7133 7619 7171
rect 7487 7099 7493 7133
rect 7527 7099 7579 7133
rect 7613 7099 7619 7133
rect 7487 7061 7619 7099
rect 7487 7027 7493 7061
rect 7527 7027 7579 7061
rect 7613 7027 7619 7061
rect 7487 6989 7619 7027
rect 7487 6955 7493 6989
rect 7527 6955 7579 6989
rect 7613 6955 7619 6989
rect 7487 6917 7619 6955
rect 7487 6883 7493 6917
rect 7527 6883 7579 6917
rect 7613 6883 7619 6917
rect 7487 6845 7619 6883
rect 7487 6811 7493 6845
rect 7527 6811 7579 6845
rect 7613 6811 7619 6845
rect 7487 6773 7619 6811
rect 7487 6739 7493 6773
rect 7527 6739 7579 6773
rect 7613 6739 7619 6773
rect 7487 6701 7619 6739
rect 7487 6667 7493 6701
rect 7527 6667 7579 6701
rect 7613 6667 7619 6701
rect 7487 6629 7619 6667
rect 7487 6595 7493 6629
rect 7527 6595 7579 6629
rect 7613 6595 7619 6629
rect 7487 6557 7619 6595
rect 7487 6523 7493 6557
rect 7527 6523 7579 6557
rect 7613 6523 7619 6557
rect 7487 6485 7619 6523
rect 7487 6451 7493 6485
rect 7527 6451 7579 6485
rect 7613 6451 7619 6485
rect 7487 6413 7619 6451
rect 7487 6379 7493 6413
rect 7527 6379 7579 6413
rect 7613 6379 7619 6413
rect 7487 6341 7619 6379
rect 7487 6307 7493 6341
rect 7527 6307 7579 6341
rect 7613 6307 7619 6341
rect 7487 6269 7619 6307
rect 7487 6235 7493 6269
rect 7527 6235 7579 6269
rect 7613 6235 7619 6269
rect 7487 6197 7619 6235
rect 7487 6163 7493 6197
rect 7527 6163 7579 6197
rect 7613 6163 7619 6197
rect 7487 6125 7619 6163
rect 7487 6091 7493 6125
rect 7527 6091 7579 6125
rect 7613 6091 7619 6125
rect 7487 6053 7619 6091
rect 7487 6019 7493 6053
rect 7527 6019 7579 6053
rect 7613 6019 7619 6053
rect 7487 5981 7619 6019
rect 7487 5947 7493 5981
rect 7527 5947 7579 5981
rect 7613 5947 7619 5981
rect 7487 5909 7619 5947
tri 2325 5875 2331 5881 sw
tri 7481 5875 7487 5881 se
rect 7487 5875 7493 5909
rect 7527 5875 7579 5909
rect 7613 5875 7619 5909
rect 2319 5847 2331 5875
tri 2331 5847 2359 5875 sw
tri 7456 5850 7481 5875 se
rect 7481 5850 7619 5875
tri 5195 5847 5198 5850 se
rect 5198 5847 5204 5850
rect 2319 5841 5204 5847
rect 2319 5807 2363 5841
rect 2397 5807 2436 5841
rect 2470 5807 2509 5841
rect 2543 5807 2582 5841
rect 2616 5807 2655 5841
rect 2689 5807 2728 5841
rect 2762 5807 2801 5841
rect 2835 5807 2874 5841
rect 2908 5807 2947 5841
rect 2981 5807 3020 5841
rect 3054 5807 3093 5841
rect 3127 5807 3166 5841
rect 3200 5807 3239 5841
rect 3273 5807 3312 5841
rect 3346 5807 3385 5841
rect 3419 5807 3458 5841
rect 3492 5807 3531 5841
rect 3565 5807 3604 5841
rect 3638 5807 3677 5841
rect 3711 5807 3750 5841
rect 3784 5807 3823 5841
rect 3857 5807 3896 5841
rect 3930 5807 3969 5841
rect 4003 5807 4042 5841
rect 4076 5807 4115 5841
rect 4149 5807 4188 5841
rect 4222 5807 4261 5841
rect 4295 5807 4334 5841
rect 4368 5807 4407 5841
rect 4441 5807 4480 5841
rect 4514 5807 4553 5841
rect 4587 5807 4626 5841
rect 4660 5807 4699 5841
rect 4733 5807 4772 5841
rect 4806 5807 4845 5841
rect 4879 5807 4918 5841
rect 4952 5807 4991 5841
rect 5025 5807 5064 5841
rect 5098 5807 5137 5841
rect 5171 5807 5204 5841
rect 2319 5801 5204 5807
rect 2319 5305 2325 5801
tri 2325 5767 2359 5801 nw
tri 5195 5798 5198 5801 ne
rect 5198 5798 5204 5801
rect 5256 5798 5268 5850
rect 5320 5798 5332 5850
rect 5384 5841 5396 5850
rect 5448 5841 5460 5850
rect 5512 5841 5524 5850
rect 5576 5841 5588 5850
rect 5640 5841 5652 5850
rect 5390 5807 5396 5841
rect 5640 5807 5648 5841
rect 5384 5798 5396 5807
rect 5448 5798 5460 5807
rect 5512 5798 5524 5807
rect 5576 5798 5588 5807
rect 5640 5798 5652 5807
rect 5704 5798 5716 5850
rect 5768 5798 5780 5850
rect 5832 5798 5844 5850
rect 5896 5841 5908 5850
rect 5960 5841 5972 5850
rect 6024 5841 6036 5850
rect 6088 5841 6100 5850
rect 6152 5841 6164 5850
rect 5901 5807 5908 5841
rect 6152 5807 6159 5841
rect 5896 5798 5908 5807
rect 5960 5798 5972 5807
rect 6024 5798 6036 5807
rect 6088 5798 6100 5807
rect 6152 5798 6164 5807
rect 6216 5798 6228 5850
rect 6280 5798 6292 5850
rect 6344 5798 6356 5850
rect 6408 5841 6420 5850
rect 6472 5841 6484 5850
rect 6536 5841 6548 5850
rect 6600 5841 6612 5850
rect 6664 5841 6676 5850
rect 6412 5807 6420 5841
rect 6664 5807 6670 5841
rect 6408 5798 6420 5807
rect 6472 5798 6484 5807
rect 6536 5798 6548 5807
rect 6600 5798 6612 5807
rect 6664 5798 6676 5807
rect 6728 5798 6740 5850
rect 6792 5798 6804 5850
rect 6856 5798 6868 5850
rect 6920 5841 6932 5850
rect 6984 5841 6996 5850
rect 7048 5841 7060 5850
rect 7112 5841 7124 5850
rect 7176 5841 7188 5850
rect 6923 5807 6932 5841
rect 7176 5807 7181 5841
rect 6920 5798 6932 5807
rect 6984 5798 6996 5807
rect 7048 5798 7060 5807
rect 7112 5798 7124 5807
rect 7176 5798 7188 5807
rect 7240 5798 7252 5850
rect 7304 5798 7316 5850
rect 7368 5847 7374 5850
tri 7374 5847 7377 5850 sw
tri 7453 5847 7456 5850 se
rect 7456 5847 7619 5850
rect 7368 5841 7619 5847
rect 7368 5807 7397 5841
rect 7431 5837 7619 5841
rect 7431 5807 7493 5837
rect 7368 5803 7493 5807
rect 7527 5803 7579 5837
rect 7613 5803 7619 5837
rect 7368 5801 7619 5803
rect 7368 5798 7374 5801
tri 7374 5798 7377 5801 nw
tri 7453 5798 7456 5801 ne
rect 7456 5798 7619 5801
tri 7456 5767 7487 5798 ne
rect 7487 5765 7619 5798
rect 7487 5731 7493 5765
rect 7527 5731 7579 5765
rect 7613 5731 7619 5765
rect 7487 5693 7619 5731
rect 7487 5659 7493 5693
rect 7527 5659 7579 5693
rect 7613 5659 7619 5693
rect 2468 5602 2474 5654
rect 2526 5602 2539 5654
rect 2591 5602 2604 5654
rect 2656 5645 7380 5654
rect 2674 5611 2713 5645
rect 2747 5611 2786 5645
rect 2820 5611 2859 5645
rect 2893 5611 2932 5645
rect 2966 5611 3005 5645
rect 3039 5611 3078 5645
rect 3112 5611 3151 5645
rect 3185 5611 3224 5645
rect 3258 5611 3297 5645
rect 3331 5611 3370 5645
rect 3404 5611 3443 5645
rect 3477 5611 3516 5645
rect 3550 5611 3589 5645
rect 3623 5611 3662 5645
rect 3696 5611 3735 5645
rect 3769 5611 3808 5645
rect 3842 5611 3881 5645
rect 3915 5611 3954 5645
rect 3988 5611 4027 5645
rect 4061 5611 4100 5645
rect 4134 5611 4173 5645
rect 4207 5611 4246 5645
rect 4280 5611 4319 5645
rect 4353 5611 4392 5645
rect 4426 5611 4465 5645
rect 4499 5611 4538 5645
rect 4572 5611 4611 5645
rect 4645 5611 4684 5645
rect 4718 5611 4757 5645
rect 4791 5611 4830 5645
rect 4864 5611 4903 5645
rect 4937 5611 4976 5645
rect 5010 5611 5049 5645
rect 5083 5611 5122 5645
rect 5156 5611 5195 5645
rect 5229 5611 5268 5645
rect 5302 5611 5341 5645
rect 5375 5611 5414 5645
rect 5448 5611 5487 5645
rect 5521 5611 5560 5645
rect 5594 5611 5633 5645
rect 5667 5611 5706 5645
rect 5740 5611 5778 5645
rect 5812 5611 5850 5645
rect 5884 5611 5922 5645
rect 5956 5611 5994 5645
rect 6028 5611 6066 5645
rect 6100 5611 6138 5645
rect 6172 5611 6210 5645
rect 6244 5611 6282 5645
rect 6316 5611 6354 5645
rect 6388 5611 6426 5645
rect 6460 5611 6498 5645
rect 6532 5611 6570 5645
rect 6604 5611 6642 5645
rect 6676 5611 6714 5645
rect 6748 5611 6786 5645
rect 6820 5611 6858 5645
rect 6892 5611 6930 5645
rect 6964 5611 7002 5645
rect 7036 5611 7380 5645
rect 2656 5602 7380 5611
rect 7487 5621 7619 5659
rect 7487 5587 7493 5621
rect 7527 5587 7579 5621
rect 7613 5587 7619 5621
rect 2681 5557 3041 5558
rect 2681 5546 2798 5557
rect 2681 5512 2687 5546
rect 2721 5512 2798 5546
rect 2681 5505 2798 5512
rect 2850 5505 2891 5557
rect 2943 5505 2983 5557
rect 3035 5505 3041 5557
rect 2681 5479 3041 5505
rect 2681 5472 2798 5479
rect 2681 5438 2687 5472
rect 2721 5438 2798 5472
rect 2681 5427 2798 5438
rect 2850 5427 2891 5479
rect 2943 5427 2983 5479
rect 3035 5427 3041 5479
rect 7487 5549 7619 5587
rect 7487 5515 7493 5549
rect 7527 5515 7579 5549
rect 7613 5515 7619 5549
rect 7487 5477 7619 5515
rect 7487 5443 7493 5477
rect 7527 5443 7579 5477
rect 7613 5443 7619 5477
rect 2681 5405 2738 5427
tri 2738 5405 2760 5427 nw
rect 7487 5405 7619 5443
rect 2681 5398 2727 5405
rect 2681 5364 2687 5398
rect 2721 5364 2727 5398
tri 2727 5394 2738 5405 nw
rect 2135 5266 2325 5305
rect 2135 5232 2141 5266
rect 2175 5232 2213 5266
rect 2247 5232 2285 5266
rect 2319 5232 2325 5266
rect 2135 5193 2325 5232
rect 2135 5159 2141 5193
rect 2175 5159 2213 5193
rect 2247 5159 2285 5193
rect 2319 5159 2325 5193
rect 2135 5120 2325 5159
rect 2135 5086 2141 5120
rect 2175 5086 2213 5120
rect 2247 5086 2285 5120
rect 2319 5086 2325 5120
rect 2135 5047 2325 5086
rect 2135 5013 2141 5047
rect 2175 5013 2213 5047
rect 2247 5013 2285 5047
rect 2319 5013 2325 5047
rect 2135 4974 2325 5013
rect 2135 4940 2141 4974
rect 2175 4940 2213 4974
rect 2247 4940 2285 4974
rect 2319 4940 2325 4974
rect 2135 4901 2325 4940
rect 2135 4867 2141 4901
rect 2175 4867 2213 4901
rect 2247 4867 2285 4901
rect 2319 4867 2325 4901
rect 2135 4828 2325 4867
rect 2135 4794 2141 4828
rect 2175 4794 2213 4828
rect 2247 4794 2285 4828
rect 2319 4794 2325 4828
rect 2135 4755 2325 4794
rect 2135 4721 2141 4755
rect 2175 4721 2213 4755
rect 2247 4721 2285 4755
rect 2319 4721 2325 4755
rect 2135 4682 2325 4721
rect 2135 4648 2141 4682
rect 2175 4648 2213 4682
rect 2247 4648 2285 4682
rect 2319 4648 2325 4682
rect 2135 4609 2325 4648
rect 2135 4575 2141 4609
rect 2175 4575 2213 4609
rect 2247 4575 2285 4609
rect 2319 4575 2325 4609
rect 2135 4536 2325 4575
rect 2135 4502 2141 4536
rect 2175 4502 2213 4536
rect 2247 4502 2285 4536
rect 2319 4502 2325 4536
rect 2135 4463 2325 4502
rect 2135 4429 2141 4463
rect 2175 4429 2213 4463
rect 2247 4429 2285 4463
rect 2319 4429 2325 4463
rect 2135 4390 2325 4429
rect 2135 4356 2141 4390
rect 2175 4356 2213 4390
rect 2247 4356 2285 4390
rect 2319 4356 2325 4390
rect 2135 4317 2325 4356
rect 2135 4283 2141 4317
rect 2175 4283 2213 4317
rect 2247 4283 2285 4317
rect 2319 4283 2325 4317
rect 2135 4244 2325 4283
rect 2135 4210 2141 4244
rect 2175 4210 2213 4244
rect 2247 4210 2285 4244
rect 2319 4210 2325 4244
rect 2135 4171 2325 4210
rect 2135 4137 2141 4171
rect 2175 4137 2213 4171
rect 2247 4137 2285 4171
rect 2319 4137 2325 4171
rect 2135 4098 2325 4137
rect 2135 4064 2141 4098
rect 2175 4064 2213 4098
rect 2247 4064 2285 4098
rect 2319 4064 2325 4098
rect 2589 5319 2635 5331
rect 2589 5285 2595 5319
rect 2629 5285 2635 5319
rect 2589 5245 2635 5285
rect 2589 5211 2595 5245
rect 2629 5211 2635 5245
rect 2589 5171 2635 5211
rect 2589 5137 2595 5171
rect 2629 5137 2635 5171
rect 2589 5097 2635 5137
rect 2589 5063 2595 5097
rect 2629 5063 2635 5097
rect 2589 5023 2635 5063
rect 2589 4989 2595 5023
rect 2629 4989 2635 5023
rect 2589 4949 2635 4989
rect 2589 4915 2595 4949
rect 2629 4915 2635 4949
rect 2589 4875 2635 4915
rect 2589 4841 2595 4875
rect 2629 4841 2635 4875
rect 2589 4801 2635 4841
rect 2589 4767 2595 4801
rect 2629 4767 2635 4801
rect 2589 4727 2635 4767
rect 2589 4693 2595 4727
rect 2629 4693 2635 4727
rect 2589 4653 2635 4693
rect 2589 4619 2595 4653
rect 2629 4619 2635 4653
rect 2589 4579 2635 4619
rect 2589 4545 2595 4579
rect 2629 4545 2635 4579
rect 2589 4504 2635 4545
rect 2589 4470 2595 4504
rect 2629 4470 2635 4504
rect 2589 4429 2635 4470
rect 2589 4395 2595 4429
rect 2629 4395 2635 4429
rect 2589 4354 2635 4395
rect 2589 4320 2595 4354
rect 2629 4320 2635 4354
rect 2589 4279 2635 4320
rect 2589 4245 2595 4279
rect 2629 4245 2635 4279
rect 2589 4204 2635 4245
rect 2589 4170 2595 4204
rect 2629 4170 2635 4204
rect 2589 4141 2635 4170
rect 2681 5324 2727 5364
rect 7487 5371 7493 5405
rect 7527 5371 7579 5405
rect 7613 5371 7619 5405
rect 7487 5333 7619 5371
rect 2681 5290 2687 5324
rect 2721 5290 2727 5324
rect 2681 5250 2727 5290
rect 2681 5216 2687 5250
rect 2721 5216 2727 5250
rect 2681 5176 2727 5216
rect 2681 5142 2687 5176
rect 2721 5142 2727 5176
rect 2681 5102 2727 5142
rect 2681 5068 2687 5102
rect 2721 5068 2727 5102
rect 2681 5028 2727 5068
rect 2681 4994 2687 5028
rect 2721 4994 2727 5028
rect 2681 4954 2727 4994
rect 2681 4920 2687 4954
rect 2721 4920 2727 4954
rect 2681 4879 2727 4920
rect 2681 4845 2687 4879
rect 2721 4845 2727 4879
rect 2681 4804 2727 4845
rect 2681 4770 2687 4804
rect 2721 4770 2727 4804
rect 2681 4729 2727 4770
rect 2681 4695 2687 4729
rect 2721 4695 2727 4729
rect 2681 4654 2727 4695
rect 2681 4620 2687 4654
rect 2721 4620 2727 4654
rect 2681 4579 2727 4620
rect 2681 4545 2687 4579
rect 2721 4545 2727 4579
rect 2681 4504 2727 4545
rect 2681 4470 2687 4504
rect 2721 4470 2727 4504
rect 2681 4429 2727 4470
rect 2681 4395 2687 4429
rect 2721 4395 2727 4429
rect 2681 4354 2727 4395
rect 2681 4320 2687 4354
rect 2721 4320 2727 4354
rect 2681 4279 2727 4320
rect 2681 4245 2687 4279
rect 2721 4245 2727 4279
rect 2681 4204 2727 4245
rect 2681 4170 2687 4204
rect 2721 4170 2727 4204
rect 2681 4158 2727 4170
rect 2773 5319 2819 5331
rect 2773 5285 2779 5319
rect 2813 5285 2819 5319
rect 2773 5245 2819 5285
rect 2773 5211 2779 5245
rect 2813 5211 2819 5245
rect 2773 5171 2819 5211
rect 2773 5137 2779 5171
rect 2813 5137 2819 5171
rect 2773 5097 2819 5137
rect 2773 5063 2779 5097
rect 2813 5063 2819 5097
rect 2773 5023 2819 5063
rect 2773 4989 2779 5023
rect 2813 4989 2819 5023
rect 2773 4949 2819 4989
rect 2773 4915 2779 4949
rect 2813 4915 2819 4949
rect 2773 4875 2819 4915
rect 2773 4841 2779 4875
rect 2813 4841 2819 4875
rect 2773 4801 2819 4841
rect 2773 4767 2779 4801
rect 2813 4767 2819 4801
rect 3621 5319 3677 5331
rect 3621 5285 3632 5319
rect 3666 5285 3677 5319
rect 3621 5244 3677 5285
rect 3621 5210 3632 5244
rect 3666 5210 3677 5244
rect 3621 5169 3677 5210
rect 3621 5135 3632 5169
rect 3666 5135 3677 5169
rect 3621 5094 3677 5135
rect 3621 5060 3632 5094
rect 3666 5060 3677 5094
rect 3621 5019 3677 5060
rect 3621 4985 3632 5019
rect 3666 4985 3677 5019
rect 3621 4944 3677 4985
rect 3621 4910 3632 4944
rect 3666 4910 3677 4944
rect 3621 4869 3677 4910
rect 3621 4835 3632 4869
rect 3666 4835 3677 4869
rect 3621 4794 3677 4835
rect 2773 4760 2819 4767
tri 2819 4760 2849 4790 sw
tri 3609 4760 3621 4772 se
rect 3621 4760 3632 4794
rect 3666 4760 3677 4794
rect 4480 5319 4536 5331
rect 4480 5285 4491 5319
rect 4525 5285 4536 5319
rect 4480 5244 4536 5285
rect 4480 5210 4491 5244
rect 4525 5210 4536 5244
rect 4480 5169 4536 5210
rect 4480 5135 4491 5169
rect 4525 5135 4536 5169
rect 4480 5094 4536 5135
rect 4480 5060 4491 5094
rect 4525 5060 4536 5094
rect 4480 5019 4536 5060
rect 4480 4985 4491 5019
rect 4525 4985 4536 5019
rect 4480 4944 4536 4985
rect 4480 4910 4491 4944
rect 4525 4910 4536 4944
rect 4480 4869 4536 4910
rect 4480 4835 4491 4869
rect 4525 4835 4536 4869
rect 4480 4794 4536 4835
tri 3677 4760 3689 4772 sw
tri 4468 4760 4480 4772 se
rect 4480 4760 4491 4794
rect 4525 4760 4536 4794
rect 5336 5319 5392 5331
rect 5336 5285 5347 5319
rect 5381 5285 5392 5319
rect 5336 5244 5392 5285
rect 5336 5210 5347 5244
rect 5381 5210 5392 5244
rect 5336 5169 5392 5210
rect 5336 5135 5347 5169
rect 5381 5135 5392 5169
rect 5336 5094 5392 5135
rect 5336 5060 5347 5094
rect 5381 5060 5392 5094
rect 5336 5019 5392 5060
rect 5336 4985 5347 5019
rect 5381 4985 5392 5019
rect 5336 4944 5392 4985
rect 5336 4910 5347 4944
rect 5381 4910 5392 4944
rect 5336 4869 5392 4910
rect 5336 4835 5347 4869
rect 5381 4835 5392 4869
rect 5336 4794 5392 4835
tri 4536 4760 4548 4772 sw
tri 5324 4760 5336 4772 se
rect 5336 4760 5347 4794
rect 5381 4760 5392 4794
rect 6195 5319 6251 5331
rect 6195 5285 6206 5319
rect 6240 5285 6251 5319
rect 6195 5244 6251 5285
rect 6195 5210 6206 5244
rect 6240 5210 6251 5244
rect 6195 5169 6251 5210
rect 6195 5135 6206 5169
rect 6240 5135 6251 5169
rect 6195 5094 6251 5135
rect 6195 5060 6206 5094
rect 6240 5060 6251 5094
rect 6195 5019 6251 5060
rect 6195 4985 6206 5019
rect 6240 4985 6251 5019
rect 6195 4944 6251 4985
rect 6195 4910 6206 4944
rect 6240 4910 6251 4944
rect 6195 4869 6251 4910
rect 6195 4835 6206 4869
rect 6240 4835 6251 4869
rect 6195 4794 6251 4835
tri 5392 4760 5404 4772 sw
tri 6183 4760 6195 4772 se
rect 6195 4760 6206 4794
rect 6240 4760 6251 4794
rect 7048 5319 7104 5331
rect 7048 5285 7059 5319
rect 7093 5285 7104 5319
rect 7048 5244 7104 5285
rect 7048 5210 7059 5244
rect 7093 5210 7104 5244
rect 7048 5169 7104 5210
rect 7048 5135 7059 5169
rect 7093 5135 7104 5169
rect 7048 5094 7104 5135
rect 7048 5060 7059 5094
rect 7093 5060 7104 5094
rect 7048 5019 7104 5060
rect 7048 4985 7059 5019
rect 7093 4985 7104 5019
rect 7048 4944 7104 4985
rect 7048 4910 7059 4944
rect 7093 4910 7104 4944
rect 7048 4869 7104 4910
rect 7048 4835 7059 4869
rect 7093 4835 7104 4869
rect 7048 4794 7104 4835
tri 6251 4760 6263 4772 sw
tri 7036 4760 7048 4772 se
rect 7048 4760 7059 4794
rect 7093 4760 7104 4794
rect 7487 5299 7493 5333
rect 7527 5299 7579 5333
rect 7613 5299 7619 5333
rect 7487 5261 7619 5299
rect 7487 5227 7493 5261
rect 7527 5227 7579 5261
rect 7613 5227 7619 5261
rect 7487 5189 7619 5227
rect 7487 5155 7493 5189
rect 7527 5155 7579 5189
rect 7613 5155 7619 5189
rect 7487 5117 7619 5155
rect 7487 5083 7493 5117
rect 7527 5083 7579 5117
rect 7613 5083 7619 5117
rect 7487 5045 7619 5083
rect 7487 5011 7493 5045
rect 7527 5011 7579 5045
rect 7613 5011 7619 5045
rect 7487 4973 7619 5011
rect 7487 4939 7493 4973
rect 7527 4939 7579 4973
rect 7613 4939 7619 4973
rect 7487 4901 7619 4939
rect 7487 4867 7493 4901
rect 7527 4867 7579 4901
rect 7613 4867 7619 4901
rect 7487 4829 7619 4867
rect 7487 4795 7493 4829
rect 7527 4795 7579 4829
rect 7613 4795 7619 4829
rect 2773 4757 2849 4760
tri 2849 4757 2852 4760 sw
tri 3606 4757 3609 4760 se
rect 3609 4757 3689 4760
tri 3689 4757 3692 4760 sw
tri 4465 4757 4468 4760 se
rect 4468 4757 4548 4760
tri 4548 4757 4551 4760 sw
tri 5321 4757 5324 4760 se
rect 5324 4757 5404 4760
tri 5404 4757 5407 4760 sw
tri 6180 4757 6183 4760 se
rect 6183 4757 6263 4760
tri 6263 4757 6266 4760 sw
tri 7033 4757 7036 4760 se
rect 7036 4757 7104 4760
tri 7104 4757 7119 4772 sw
rect 7487 4757 7619 4795
rect 2773 4747 2852 4757
tri 2852 4747 2862 4757 sw
tri 3596 4747 3606 4757 se
rect 3606 4747 3692 4757
tri 3692 4747 3702 4757 sw
tri 4455 4747 4465 4757 se
rect 4465 4747 4551 4757
tri 4551 4747 4561 4757 sw
tri 5311 4747 5321 4757 se
rect 5321 4747 5407 4757
tri 5407 4747 5417 4757 sw
tri 6170 4747 6180 4757 se
rect 6180 4747 6266 4757
tri 6266 4747 6276 4757 sw
tri 7023 4747 7033 4757 se
rect 7033 4747 7119 4757
tri 7119 4747 7129 4757 sw
rect 2773 4743 7374 4747
rect 2773 4727 5204 4743
rect 2773 4693 2779 4727
rect 2813 4719 5204 4727
rect 2813 4693 3632 4719
rect 2773 4685 3632 4693
rect 3666 4685 4491 4719
rect 4525 4691 5204 4719
rect 5256 4691 5336 4743
rect 5388 4691 5468 4743
rect 5520 4691 5600 4743
rect 5652 4691 5732 4743
rect 5784 4691 5864 4743
rect 5916 4691 5996 4743
rect 6048 4691 6128 4743
rect 6180 4719 6260 4743
rect 6180 4691 6206 4719
rect 4525 4685 5347 4691
rect 5381 4685 6206 4691
rect 6240 4691 6260 4719
rect 6312 4691 6392 4743
rect 6444 4691 6524 4743
rect 6576 4691 6656 4743
rect 6708 4691 6788 4743
rect 6840 4691 6920 4743
rect 6972 4691 7052 4743
rect 7104 4691 7184 4743
rect 7236 4691 7316 4743
rect 7368 4691 7374 4743
rect 6240 4685 7059 4691
rect 7093 4685 7374 4691
rect 2773 4653 7374 4685
rect 2773 4619 2779 4653
rect 2813 4644 7374 4653
rect 2813 4619 3632 4644
rect 2773 4610 3632 4619
rect 3666 4610 4491 4644
rect 4525 4635 5347 4644
rect 5381 4635 6206 4644
rect 4525 4610 5204 4635
rect 2773 4583 5204 4610
rect 5256 4583 5336 4635
rect 5388 4583 5468 4635
rect 5520 4583 5600 4635
rect 5652 4583 5732 4635
rect 5784 4583 5864 4635
rect 5916 4583 5996 4635
rect 6048 4583 6128 4635
rect 6180 4610 6206 4635
rect 6240 4635 7059 4644
rect 7093 4635 7374 4644
rect 6240 4610 6260 4635
rect 6180 4583 6260 4610
rect 6312 4583 6392 4635
rect 6444 4583 6524 4635
rect 6576 4583 6656 4635
rect 6708 4583 6788 4635
rect 6840 4583 6920 4635
rect 6972 4583 7052 4635
rect 7104 4583 7184 4635
rect 7236 4583 7316 4635
rect 7368 4583 7374 4635
rect 2773 4579 7374 4583
rect 2773 4545 2779 4579
rect 2813 4569 7374 4579
rect 2813 4545 3632 4569
rect 2773 4535 3632 4545
rect 3666 4535 4491 4569
rect 4525 4535 5347 4569
rect 5381 4535 6206 4569
rect 6240 4535 7059 4569
rect 7093 4535 7374 4569
rect 2773 4527 7374 4535
rect 2773 4504 5204 4527
rect 2773 4470 2779 4504
rect 2813 4494 5204 4504
rect 2813 4470 3632 4494
rect 2773 4460 3632 4470
rect 3666 4460 4491 4494
rect 4525 4475 5204 4494
rect 5256 4475 5336 4527
rect 5388 4475 5468 4527
rect 5520 4475 5600 4527
rect 5652 4475 5732 4527
rect 5784 4475 5864 4527
rect 5916 4475 5996 4527
rect 6048 4475 6128 4527
rect 6180 4494 6260 4527
rect 6180 4475 6206 4494
rect 4525 4460 5347 4475
rect 5381 4460 6206 4475
rect 6240 4475 6260 4494
rect 6312 4475 6392 4527
rect 6444 4475 6524 4527
rect 6576 4475 6656 4527
rect 6708 4475 6788 4527
rect 6840 4475 6920 4527
rect 6972 4475 7052 4527
rect 7104 4475 7184 4527
rect 7236 4475 7316 4527
rect 7368 4475 7374 4527
rect 6240 4460 7059 4475
rect 7093 4460 7374 4475
rect 2773 4429 7374 4460
rect 2773 4395 2779 4429
rect 2813 4419 7374 4429
rect 2813 4395 3632 4419
rect 2773 4385 3632 4395
rect 3666 4385 4491 4419
rect 4525 4385 5204 4419
rect 2773 4367 5204 4385
rect 5256 4367 5336 4419
rect 5388 4367 5468 4419
rect 5520 4367 5600 4419
rect 5652 4367 5732 4419
rect 5784 4367 5864 4419
rect 5916 4367 5996 4419
rect 6048 4367 6128 4419
rect 6180 4385 6206 4419
rect 6240 4385 6260 4419
rect 6180 4367 6260 4385
rect 6312 4367 6392 4419
rect 6444 4367 6524 4419
rect 6576 4367 6656 4419
rect 6708 4367 6788 4419
rect 6840 4367 6920 4419
rect 6972 4367 7052 4419
rect 7104 4367 7184 4419
rect 7236 4367 7316 4419
rect 7368 4367 7374 4419
rect 2773 4354 7374 4367
rect 2773 4320 2779 4354
rect 2813 4344 7374 4354
rect 2813 4320 3632 4344
rect 2773 4310 3632 4320
rect 3666 4310 4491 4344
rect 4525 4311 5347 4344
rect 5381 4311 6206 4344
rect 4525 4310 5204 4311
rect 2773 4279 5204 4310
rect 2773 4245 2779 4279
rect 2813 4269 5204 4279
rect 2813 4245 3632 4269
rect 2773 4235 3632 4245
rect 3666 4235 4491 4269
rect 4525 4259 5204 4269
rect 5256 4259 5336 4311
rect 5388 4259 5468 4311
rect 5520 4259 5600 4311
rect 5652 4259 5732 4311
rect 5784 4259 5864 4311
rect 5916 4259 5996 4311
rect 6048 4259 6128 4311
rect 6180 4310 6206 4311
rect 6240 4311 7059 4344
rect 7093 4311 7374 4344
rect 6240 4310 6260 4311
rect 6180 4269 6260 4310
rect 6180 4259 6206 4269
rect 4525 4235 5347 4259
rect 5381 4235 6206 4259
rect 6240 4259 6260 4269
rect 6312 4259 6392 4311
rect 6444 4259 6524 4311
rect 6576 4259 6656 4311
rect 6708 4259 6788 4311
rect 6840 4259 6920 4311
rect 6972 4259 7052 4311
rect 7104 4259 7184 4311
rect 7236 4259 7316 4311
rect 7368 4259 7374 4311
rect 6240 4235 7059 4259
rect 7093 4235 7374 4259
rect 2773 4204 7374 4235
rect 2773 4170 2779 4204
rect 2813 4203 7374 4204
rect 2813 4193 5204 4203
rect 2813 4170 3632 4193
rect 2773 4159 3632 4170
rect 3666 4159 4491 4193
rect 4525 4159 5204 4193
rect 2773 4151 5204 4159
rect 5256 4151 5336 4203
rect 5388 4151 5468 4203
rect 5520 4151 5600 4203
rect 5652 4151 5732 4203
rect 5784 4151 5864 4203
rect 5916 4151 5996 4203
rect 6048 4151 6128 4203
rect 6180 4193 6260 4203
rect 6180 4159 6206 4193
rect 6240 4159 6260 4193
rect 6180 4151 6260 4159
rect 6312 4151 6392 4203
rect 6444 4151 6524 4203
rect 6576 4151 6656 4203
rect 6708 4151 6788 4203
rect 6840 4151 6920 4203
rect 6972 4151 7052 4203
rect 7104 4151 7184 4203
rect 7236 4151 7316 4203
rect 7368 4151 7374 4203
rect 2773 4147 7374 4151
rect 7487 4723 7493 4757
rect 7527 4723 7579 4757
rect 7613 4723 7619 4757
rect 7487 4685 7619 4723
rect 7487 4651 7493 4685
rect 7527 4651 7579 4685
rect 7613 4651 7619 4685
rect 7487 4613 7619 4651
rect 7487 4579 7493 4613
rect 7527 4579 7579 4613
rect 7613 4579 7619 4613
rect 7487 4540 7619 4579
rect 7487 4506 7493 4540
rect 7527 4506 7579 4540
rect 7613 4506 7619 4540
rect 7487 4467 7619 4506
rect 7487 4433 7493 4467
rect 7527 4433 7579 4467
rect 7613 4433 7619 4467
rect 7487 4394 7619 4433
rect 7487 4360 7493 4394
rect 7527 4360 7579 4394
rect 7613 4360 7619 4394
rect 7487 4321 7619 4360
rect 7487 4287 7493 4321
rect 7527 4287 7579 4321
rect 7613 4287 7619 4321
rect 7487 4248 7619 4287
rect 7487 4214 7493 4248
rect 7527 4214 7579 4248
rect 7613 4214 7619 4248
rect 7487 4175 7619 4214
tri 2635 4141 2640 4146 sw
tri 2772 4141 2773 4142 se
rect 2773 4141 2839 4147
tri 2839 4141 2845 4147 nw
rect 7487 4141 7493 4175
rect 7527 4141 7579 4175
rect 7613 4141 7619 4175
rect 2589 4124 2640 4141
tri 2640 4124 2657 4141 sw
tri 2755 4124 2772 4141 se
rect 2772 4124 2822 4141
tri 2822 4124 2839 4141 nw
rect 2589 4116 2657 4124
tri 2657 4116 2665 4124 sw
tri 2747 4116 2755 4124 se
rect 2755 4116 2816 4124
tri 2816 4118 2822 4124 nw
rect 2589 4070 2816 4116
rect 7487 4102 7619 4141
rect 2135 4025 2325 4064
rect 2135 3991 2141 4025
rect 2175 3991 2213 4025
rect 2247 3991 2285 4025
rect 2319 3991 2325 4025
rect 7487 4068 7493 4102
rect 7527 4068 7579 4102
rect 7613 4068 7619 4102
rect 7487 4029 7619 4068
tri 7470 3995 7487 4012 se
rect 7487 3995 7493 4029
rect 7527 3995 7579 4029
rect 7613 3995 7619 4029
rect 2135 3978 2325 3991
tri 7458 3983 7470 3995 se
rect 7470 3983 7619 3995
tri 2325 3978 2330 3983 sw
tri 7453 3978 7458 3983 se
rect 7458 3978 7619 3983
rect 2135 3949 2330 3978
tri 2330 3949 2359 3978 sw
tri 7424 3949 7453 3978 se
rect 7453 3949 7619 3978
rect 2135 3943 5204 3949
rect 5256 3943 5339 3949
rect 5391 3943 5474 3949
rect 5526 3943 5609 3949
rect 5661 3943 5744 3949
rect 5796 3943 5879 3949
rect 5931 3943 6014 3949
rect 6066 3943 6149 3949
rect 6201 3943 6284 3949
rect 6336 3943 6419 3949
rect 6471 3943 6553 3949
rect 6605 3943 6687 3949
rect 6739 3943 6821 3949
rect 6873 3943 6955 3949
rect 7007 3943 7089 3949
rect 7141 3943 7223 3949
rect 7275 3943 7619 3949
rect 2135 3909 2147 3943
rect 2181 3909 2220 3943
rect 2254 3909 2293 3943
rect 2327 3909 2366 3943
rect 2400 3909 2439 3943
rect 2473 3909 2512 3943
rect 2546 3909 2585 3943
rect 2619 3909 2658 3943
rect 2692 3909 2731 3943
rect 2765 3909 2804 3943
rect 2838 3909 2877 3943
rect 2911 3909 2950 3943
rect 2984 3909 3023 3943
rect 2135 3871 3023 3909
rect 2135 3837 2147 3871
rect 2181 3837 2220 3871
rect 2254 3837 2293 3871
rect 2327 3837 2366 3871
rect 2400 3837 2439 3871
rect 2473 3837 2512 3871
rect 2546 3837 2585 3871
rect 2619 3837 2658 3871
rect 2692 3837 2731 3871
rect 2765 3837 2804 3871
rect 2838 3837 2877 3871
rect 2911 3837 2950 3871
rect 2984 3837 3023 3871
rect 7593 3837 7619 3943
rect 2135 3831 5204 3837
rect 5256 3831 5339 3837
rect 5391 3831 5474 3837
rect 5526 3831 5609 3837
rect 5661 3831 5744 3837
rect 5796 3831 5879 3837
rect 5931 3831 6014 3837
rect 6066 3831 6149 3837
rect 6201 3831 6284 3837
rect 6336 3831 6419 3837
rect 6471 3831 6553 3837
rect 6605 3831 6687 3837
rect 6739 3831 6821 3837
rect 6873 3831 6955 3837
rect 7007 3831 7089 3837
rect 7141 3831 7223 3837
rect 7275 3831 7619 3837
rect 7727 4528 7733 9540
rect 7839 9540 8573 9640
rect 7839 4528 7877 9540
tri 7877 9506 7911 9540 nw
rect 7727 4489 7877 4528
rect 7727 4455 7733 4489
rect 7767 4455 7805 4489
rect 7839 4455 7877 4489
rect 7727 4416 7877 4455
rect 7727 4382 7733 4416
rect 7767 4382 7805 4416
rect 7839 4382 7877 4416
rect 7727 4343 7877 4382
rect 7727 4309 7733 4343
rect 7767 4309 7805 4343
rect 7839 4309 7877 4343
rect 7727 4270 7877 4309
rect 7727 4236 7733 4270
rect 7767 4236 7805 4270
rect 7839 4236 7877 4270
rect 7727 4197 7877 4236
rect 7727 4163 7733 4197
rect 7767 4163 7805 4197
rect 7839 4163 7877 4197
rect 7727 4124 7877 4163
rect 7727 4090 7733 4124
rect 7767 4090 7805 4124
rect 7839 4090 7877 4124
rect 7727 4051 7877 4090
rect 7727 4017 7733 4051
rect 7767 4017 7805 4051
rect 7839 4017 7877 4051
rect 7727 3978 7877 4017
rect 7727 3944 7733 3978
rect 7767 3944 7805 3978
rect 7839 3944 7877 3978
rect 7727 3905 7877 3944
rect 7727 3871 7733 3905
rect 7767 3871 7805 3905
rect 7839 3871 7877 3905
rect 7727 3832 7877 3871
rect 7727 3798 7733 3832
rect 7767 3798 7805 3832
rect 7839 3798 7877 3832
rect 7727 3759 7877 3798
rect 7727 3725 7733 3759
rect 7767 3725 7805 3759
rect 7839 3725 7877 3759
rect 7727 3686 7877 3725
rect 7727 3652 7733 3686
rect 7767 3652 7805 3686
rect 7839 3652 7877 3686
rect 7727 3613 7877 3652
rect 7727 3579 7733 3613
rect 7767 3579 7805 3613
rect 7839 3579 7877 3613
rect 7727 3540 7877 3579
rect 7727 3506 7733 3540
rect 7767 3506 7805 3540
rect 7839 3506 7877 3540
rect 1938 3467 2056 3491
tri 7719 3484 7727 3492 se
rect 7727 3484 7877 3506
tri 2056 3467 2073 3484 sw
tri 7702 3467 7719 3484 se
rect 7719 3467 7877 3484
rect 1938 3459 2073 3467
tri 2073 3459 2081 3467 sw
tri 7694 3459 7702 3467 se
rect 7702 3459 7733 3467
rect 1938 3453 7733 3459
rect 1938 3419 1950 3453
rect 1984 3419 2023 3453
rect 2057 3419 2096 3453
rect 2130 3419 2169 3453
rect 2203 3419 2242 3453
rect 2276 3419 2315 3453
rect 2349 3419 2388 3453
rect 2422 3419 2461 3453
rect 2495 3419 2534 3453
rect 2568 3419 2607 3453
rect 2641 3419 2680 3453
rect 2714 3419 2753 3453
rect 2787 3419 2826 3453
rect 2860 3419 2899 3453
rect 2933 3419 2972 3453
rect 3006 3419 3045 3453
rect 3079 3419 3118 3453
rect 3152 3419 3191 3453
rect 3225 3419 3264 3453
rect 3298 3419 3337 3453
rect 3371 3419 3410 3453
rect 3444 3419 3483 3453
rect 3517 3419 3556 3453
rect 3590 3419 3629 3453
rect 3663 3419 3702 3453
rect 3736 3419 3775 3453
rect 3809 3419 3848 3453
rect 3882 3419 3921 3453
rect 3955 3419 3994 3453
rect 4028 3419 4067 3453
rect 4101 3419 4140 3453
rect 4174 3419 4213 3453
rect 4247 3419 4286 3453
rect 4320 3419 4359 3453
rect 4393 3419 4432 3453
rect 4466 3419 4505 3453
rect 4539 3419 4578 3453
rect 4612 3419 4651 3453
rect 4685 3419 4724 3453
rect 4758 3419 4797 3453
rect 4831 3419 4870 3453
rect 4904 3419 4943 3453
rect 4977 3419 5016 3453
rect 5050 3419 5089 3453
rect 5123 3419 5162 3453
rect 5196 3419 5235 3453
rect 5269 3419 5308 3453
rect 5342 3419 5381 3453
rect 5415 3419 5454 3453
rect 5488 3419 5527 3453
rect 5561 3419 5600 3453
rect 5634 3419 5673 3453
rect 5707 3419 5746 3453
rect 5780 3419 5819 3453
rect 5853 3419 5892 3453
rect 5926 3419 5965 3453
rect 5999 3419 6038 3453
rect 6072 3419 6111 3453
rect 6145 3419 6184 3453
rect 6218 3419 6257 3453
rect 6291 3419 6330 3453
rect 1938 3381 6330 3419
rect 1938 3347 1950 3381
rect 1984 3347 2023 3381
rect 2057 3347 2096 3381
rect 2130 3347 2169 3381
rect 2203 3347 2242 3381
rect 2276 3347 2315 3381
rect 2349 3347 2388 3381
rect 2422 3347 2461 3381
rect 2495 3347 2534 3381
rect 2568 3347 2607 3381
rect 2641 3347 2680 3381
rect 2714 3347 2753 3381
rect 2787 3347 2826 3381
rect 2860 3347 2899 3381
rect 2933 3347 2972 3381
rect 3006 3347 3045 3381
rect 3079 3347 3118 3381
rect 3152 3347 3191 3381
rect 3225 3347 3264 3381
rect 3298 3347 3337 3381
rect 3371 3347 3410 3381
rect 3444 3347 3483 3381
rect 3517 3347 3556 3381
rect 3590 3347 3629 3381
rect 3663 3347 3702 3381
rect 3736 3347 3775 3381
rect 3809 3347 3848 3381
rect 3882 3347 3921 3381
rect 3955 3347 3994 3381
rect 4028 3347 4067 3381
rect 4101 3347 4140 3381
rect 4174 3347 4213 3381
rect 4247 3347 4286 3381
rect 4320 3347 4359 3381
rect 4393 3347 4432 3381
rect 4466 3347 4505 3381
rect 4539 3347 4578 3381
rect 4612 3347 4651 3381
rect 4685 3347 4724 3381
rect 4758 3347 4797 3381
rect 4831 3347 4870 3381
rect 4904 3347 4943 3381
rect 4977 3347 5016 3381
rect 5050 3347 5089 3381
rect 5123 3347 5162 3381
rect 5196 3347 5235 3381
rect 5269 3347 5308 3381
rect 5342 3347 5381 3381
rect 5415 3347 5454 3381
rect 5488 3347 5527 3381
rect 5561 3347 5600 3381
rect 5634 3347 5673 3381
rect 5707 3347 5746 3381
rect 5780 3347 5819 3381
rect 5853 3347 5892 3381
rect 5926 3347 5965 3381
rect 5999 3347 6038 3381
rect 6072 3347 6111 3381
rect 6145 3347 6184 3381
rect 6218 3347 6257 3381
rect 6291 3347 6330 3381
rect 7660 3433 7733 3453
rect 7767 3433 7805 3467
rect 7839 3433 7877 3467
rect 7660 3394 7877 3433
rect 7660 3360 7733 3394
rect 7767 3360 7805 3394
rect 7839 3360 7877 3394
rect 7660 3347 7877 3360
rect 1938 3341 7877 3347
tri 7701 3315 7727 3341 ne
rect 1923 3057 7573 3058
rect 1923 3049 5204 3057
rect 1923 3015 1935 3049
rect 1969 3015 2008 3049
rect 2042 3015 2081 3049
rect 2115 3015 2154 3049
rect 2188 3015 2227 3049
rect 2261 3015 2300 3049
rect 2334 3015 2373 3049
rect 2407 3015 2446 3049
rect 2480 3015 2519 3049
rect 2553 3015 2592 3049
rect 2626 3015 2665 3049
rect 2699 3015 2738 3049
rect 2772 3015 2811 3049
rect 2845 3015 2884 3049
rect 2918 3015 2957 3049
rect 2991 3015 3030 3049
rect 3064 3015 3103 3049
rect 3137 3015 3176 3049
rect 3210 3015 3249 3049
rect 3283 3015 3322 3049
rect 3356 3015 3395 3049
rect 3429 3015 3468 3049
rect 3502 3015 3541 3049
rect 3575 3015 3614 3049
rect 3648 3015 3687 3049
rect 3721 3015 3760 3049
rect 3794 3015 3833 3049
rect 3867 3015 3906 3049
rect 3940 3015 3979 3049
rect 4013 3015 4052 3049
rect 4086 3015 4125 3049
rect 4159 3015 4198 3049
rect 4232 3015 4271 3049
rect 4305 3015 4344 3049
rect 4378 3015 4417 3049
rect 4451 3015 4490 3049
rect 4524 3015 4563 3049
rect 4597 3015 4636 3049
rect 4670 3015 4709 3049
rect 4743 3015 4782 3049
rect 4816 3015 4855 3049
rect 4889 3015 4928 3049
rect 4962 3015 5001 3049
rect 5035 3015 5074 3049
rect 5108 3015 5147 3049
rect 5181 3015 5204 3049
rect 1923 3005 5204 3015
rect 5256 3005 5270 3057
rect 5322 3049 5336 3057
rect 5388 3049 5402 3057
rect 5454 3049 5468 3057
rect 5520 3049 5534 3057
rect 5586 3049 5599 3057
rect 5651 3049 5664 3057
rect 5716 3049 5729 3057
rect 5327 3015 5336 3049
rect 5400 3015 5402 3049
rect 5651 3015 5655 3049
rect 5716 3015 5727 3049
rect 5322 3005 5336 3015
rect 5388 3005 5402 3015
rect 5454 3005 5468 3015
rect 5520 3005 5534 3015
rect 5586 3005 5599 3015
rect 5651 3005 5664 3015
rect 5716 3005 5729 3015
rect 5781 3005 5794 3057
rect 5846 3005 5859 3057
rect 5911 3005 5924 3057
rect 5976 3049 5989 3057
rect 6041 3049 6054 3057
rect 6106 3049 6119 3057
rect 6171 3049 6184 3057
rect 6236 3049 6249 3057
rect 6301 3049 6314 3057
rect 6366 3049 6379 3057
rect 5977 3015 5989 3049
rect 6049 3015 6054 3049
rect 6301 3015 6303 3049
rect 6366 3015 6375 3049
rect 5976 3005 5989 3015
rect 6041 3005 6054 3015
rect 6106 3005 6119 3015
rect 6171 3005 6184 3015
rect 6236 3005 6249 3015
rect 6301 3005 6314 3015
rect 6366 3005 6379 3015
rect 6431 3005 6444 3057
rect 6496 3005 6509 3057
rect 6561 3005 6574 3057
rect 6626 3005 6639 3057
rect 6691 3049 6704 3057
rect 6756 3049 6769 3057
rect 6821 3049 6834 3057
rect 6886 3049 6899 3057
rect 6951 3049 6964 3057
rect 7016 3049 7029 3057
rect 6697 3015 6704 3049
rect 7016 3015 7023 3049
rect 6691 3005 6704 3015
rect 6756 3005 6769 3015
rect 6821 3005 6834 3015
rect 6886 3005 6899 3015
rect 6951 3005 6964 3015
rect 7016 3005 7029 3015
rect 7081 3005 7094 3057
rect 7146 3005 7159 3057
rect 7211 3005 7224 3057
rect 7276 3005 7289 3057
rect 7341 3049 7354 3057
rect 7406 3049 7419 3057
rect 7471 3049 7484 3057
rect 7536 3049 7573 3057
rect 7345 3015 7354 3049
rect 7417 3015 7419 3049
rect 7561 3015 7573 3049
rect 7341 3005 7354 3015
rect 7406 3005 7419 3015
rect 7471 3005 7484 3015
rect 7536 3005 7573 3015
rect 1923 2989 7573 3005
rect 1923 2971 5204 2989
rect 1923 2937 1935 2971
rect 1969 2937 2008 2971
rect 2042 2937 2081 2971
rect 2115 2937 2154 2971
rect 2188 2937 2227 2971
rect 2261 2937 2300 2971
rect 2334 2937 2373 2971
rect 2407 2937 2446 2971
rect 2480 2937 2519 2971
rect 2553 2937 2592 2971
rect 2626 2937 2665 2971
rect 2699 2937 2738 2971
rect 2772 2937 2811 2971
rect 2845 2937 2884 2971
rect 2918 2937 2957 2971
rect 2991 2937 3030 2971
rect 3064 2937 3103 2971
rect 3137 2937 3176 2971
rect 3210 2937 3249 2971
rect 3283 2937 3322 2971
rect 3356 2937 3395 2971
rect 3429 2937 3468 2971
rect 3502 2937 3541 2971
rect 3575 2937 3614 2971
rect 3648 2937 3687 2971
rect 3721 2937 3760 2971
rect 3794 2937 3833 2971
rect 3867 2937 3906 2971
rect 3940 2937 3979 2971
rect 4013 2937 4052 2971
rect 4086 2937 4125 2971
rect 4159 2937 4198 2971
rect 4232 2937 4271 2971
rect 4305 2937 4344 2971
rect 4378 2937 4417 2971
rect 4451 2937 4490 2971
rect 4524 2937 4563 2971
rect 4597 2937 4636 2971
rect 4670 2937 4709 2971
rect 4743 2937 4782 2971
rect 4816 2937 4855 2971
rect 4889 2937 4928 2971
rect 4962 2937 5001 2971
rect 5035 2937 5074 2971
rect 5108 2937 5147 2971
rect 5181 2937 5204 2971
rect 5256 2937 5270 2989
rect 5322 2971 5336 2989
rect 5388 2971 5402 2989
rect 5454 2971 5468 2989
rect 5520 2971 5534 2989
rect 5586 2971 5599 2989
rect 5651 2971 5664 2989
rect 5716 2971 5729 2989
rect 5327 2937 5336 2971
rect 5400 2937 5402 2971
rect 5651 2937 5655 2971
rect 5716 2937 5727 2971
rect 5781 2937 5794 2989
rect 5846 2937 5859 2989
rect 5911 2937 5924 2989
rect 5976 2971 5989 2989
rect 6041 2971 6054 2989
rect 6106 2971 6119 2989
rect 6171 2971 6184 2989
rect 6236 2971 6249 2989
rect 6301 2971 6314 2989
rect 6366 2971 6379 2989
rect 5977 2937 5989 2971
rect 6049 2937 6054 2971
rect 6301 2937 6303 2971
rect 6366 2937 6375 2971
rect 6431 2937 6444 2989
rect 6496 2937 6509 2989
rect 6561 2937 6574 2989
rect 6626 2937 6639 2989
rect 6691 2971 6704 2989
rect 6756 2971 6769 2989
rect 6821 2971 6834 2989
rect 6886 2971 6899 2989
rect 6951 2971 6964 2989
rect 7016 2971 7029 2989
rect 6697 2937 6704 2971
rect 7016 2937 7023 2971
rect 7081 2937 7094 2989
rect 7146 2937 7159 2989
rect 7211 2937 7224 2989
rect 7276 2937 7289 2989
rect 7341 2971 7354 2989
rect 7406 2971 7419 2989
rect 7471 2971 7484 2989
rect 7536 2971 7573 2989
rect 7345 2937 7354 2971
rect 7417 2937 7419 2971
rect 7561 2937 7573 2971
rect 1923 2921 7573 2937
rect 1923 2893 5204 2921
rect 1923 2859 1935 2893
rect 1969 2859 2008 2893
rect 2042 2859 2081 2893
rect 2115 2859 2154 2893
rect 2188 2859 2227 2893
rect 2261 2859 2300 2893
rect 2334 2859 2373 2893
rect 2407 2859 2446 2893
rect 2480 2859 2519 2893
rect 2553 2859 2592 2893
rect 2626 2859 2665 2893
rect 2699 2859 2738 2893
rect 2772 2859 2811 2893
rect 2845 2859 2884 2893
rect 2918 2859 2957 2893
rect 2991 2859 3030 2893
rect 3064 2859 3103 2893
rect 3137 2859 3176 2893
rect 3210 2859 3249 2893
rect 3283 2859 3322 2893
rect 3356 2859 3395 2893
rect 3429 2859 3468 2893
rect 3502 2859 3541 2893
rect 3575 2859 3614 2893
rect 3648 2859 3687 2893
rect 3721 2859 3760 2893
rect 3794 2859 3833 2893
rect 3867 2859 3906 2893
rect 3940 2859 3979 2893
rect 4013 2859 4052 2893
rect 4086 2859 4125 2893
rect 4159 2859 4198 2893
rect 4232 2859 4271 2893
rect 4305 2859 4344 2893
rect 4378 2859 4417 2893
rect 4451 2859 4490 2893
rect 4524 2859 4563 2893
rect 4597 2859 4636 2893
rect 4670 2859 4709 2893
rect 4743 2859 4782 2893
rect 4816 2859 4855 2893
rect 4889 2859 4928 2893
rect 4962 2859 5001 2893
rect 5035 2859 5074 2893
rect 5108 2859 5147 2893
rect 5181 2869 5204 2893
rect 5256 2869 5270 2921
rect 5322 2893 5336 2921
rect 5388 2893 5402 2921
rect 5454 2893 5468 2921
rect 5520 2893 5534 2921
rect 5586 2893 5599 2921
rect 5651 2893 5664 2921
rect 5716 2893 5729 2921
rect 5327 2869 5336 2893
rect 5400 2869 5402 2893
rect 5651 2869 5655 2893
rect 5716 2869 5727 2893
rect 5781 2869 5794 2921
rect 5846 2869 5859 2921
rect 5911 2869 5924 2921
rect 5976 2893 5989 2921
rect 6041 2893 6054 2921
rect 6106 2893 6119 2921
rect 6171 2893 6184 2921
rect 6236 2893 6249 2921
rect 6301 2893 6314 2921
rect 6366 2893 6379 2921
rect 5977 2869 5989 2893
rect 6049 2869 6054 2893
rect 6301 2869 6303 2893
rect 6366 2869 6375 2893
rect 6431 2869 6444 2921
rect 6496 2869 6509 2921
rect 6561 2869 6574 2921
rect 6626 2869 6639 2921
rect 6691 2893 6704 2921
rect 6756 2893 6769 2921
rect 6821 2893 6834 2921
rect 6886 2893 6899 2921
rect 6951 2893 6964 2921
rect 7016 2893 7029 2921
rect 6697 2869 6704 2893
rect 7016 2869 7023 2893
rect 7081 2869 7094 2921
rect 7146 2869 7159 2921
rect 7211 2869 7224 2921
rect 7276 2869 7289 2921
rect 7341 2893 7354 2921
rect 7406 2893 7419 2921
rect 7471 2893 7484 2921
rect 7536 2893 7573 2921
rect 7345 2869 7354 2893
rect 7417 2869 7419 2893
rect 5181 2859 5220 2869
rect 5254 2859 5293 2869
rect 5327 2859 5366 2869
rect 5400 2859 5439 2869
rect 5473 2859 5511 2869
rect 5545 2859 5583 2869
rect 5617 2859 5655 2869
rect 5689 2859 5727 2869
rect 5761 2859 5799 2869
rect 5833 2859 5871 2869
rect 5905 2859 5943 2869
rect 5977 2859 6015 2869
rect 6049 2859 6087 2869
rect 6121 2859 6159 2869
rect 6193 2859 6231 2869
rect 6265 2859 6303 2869
rect 6337 2859 6375 2869
rect 6409 2859 6447 2869
rect 6481 2859 6519 2869
rect 6553 2859 6591 2869
rect 6625 2859 6663 2869
rect 6697 2859 6735 2869
rect 6769 2859 6807 2869
rect 6841 2859 6879 2869
rect 6913 2859 6951 2869
rect 6985 2859 7023 2869
rect 7057 2859 7095 2869
rect 7129 2859 7167 2869
rect 7201 2859 7239 2869
rect 7273 2859 7311 2869
rect 7345 2859 7383 2869
rect 7417 2859 7455 2869
rect 7489 2859 7527 2869
rect 7561 2859 7573 2893
rect 1923 2853 7573 2859
rect 1923 2815 5204 2853
rect 1923 2781 1935 2815
rect 1969 2781 2008 2815
rect 2042 2781 2081 2815
rect 2115 2781 2154 2815
rect 2188 2781 2227 2815
rect 2261 2781 2300 2815
rect 2334 2781 2373 2815
rect 2407 2781 2446 2815
rect 2480 2781 2519 2815
rect 2553 2781 2592 2815
rect 2626 2781 2665 2815
rect 2699 2781 2738 2815
rect 2772 2781 2811 2815
rect 2845 2781 2884 2815
rect 2918 2781 2957 2815
rect 2991 2781 3030 2815
rect 3064 2781 3103 2815
rect 3137 2781 3176 2815
rect 3210 2781 3249 2815
rect 3283 2781 3322 2815
rect 3356 2781 3395 2815
rect 3429 2781 3468 2815
rect 3502 2781 3541 2815
rect 3575 2781 3614 2815
rect 3648 2781 3687 2815
rect 3721 2781 3760 2815
rect 3794 2781 3833 2815
rect 3867 2781 3906 2815
rect 3940 2781 3979 2815
rect 4013 2781 4052 2815
rect 4086 2781 4125 2815
rect 4159 2781 4198 2815
rect 4232 2781 4271 2815
rect 4305 2781 4344 2815
rect 4378 2781 4417 2815
rect 4451 2781 4490 2815
rect 4524 2781 4563 2815
rect 4597 2781 4636 2815
rect 4670 2781 4709 2815
rect 4743 2781 4782 2815
rect 4816 2781 4855 2815
rect 4889 2781 4928 2815
rect 4962 2781 5001 2815
rect 5035 2781 5074 2815
rect 5108 2781 5147 2815
rect 5181 2801 5204 2815
rect 5256 2801 5270 2853
rect 5322 2815 5336 2853
rect 5388 2815 5402 2853
rect 5454 2815 5468 2853
rect 5520 2815 5534 2853
rect 5586 2815 5599 2853
rect 5651 2815 5664 2853
rect 5716 2815 5729 2853
rect 5327 2801 5336 2815
rect 5400 2801 5402 2815
rect 5651 2801 5655 2815
rect 5716 2801 5727 2815
rect 5781 2801 5794 2853
rect 5846 2801 5859 2853
rect 5911 2801 5924 2853
rect 5976 2815 5989 2853
rect 6041 2815 6054 2853
rect 6106 2815 6119 2853
rect 6171 2815 6184 2853
rect 6236 2815 6249 2853
rect 6301 2815 6314 2853
rect 6366 2815 6379 2853
rect 5977 2801 5989 2815
rect 6049 2801 6054 2815
rect 6301 2801 6303 2815
rect 6366 2801 6375 2815
rect 6431 2801 6444 2853
rect 6496 2801 6509 2853
rect 6561 2801 6574 2853
rect 6626 2801 6639 2853
rect 6691 2815 6704 2853
rect 6756 2815 6769 2853
rect 6821 2815 6834 2853
rect 6886 2815 6899 2853
rect 6951 2815 6964 2853
rect 7016 2815 7029 2853
rect 6697 2801 6704 2815
rect 7016 2801 7023 2815
rect 7081 2801 7094 2853
rect 7146 2801 7159 2853
rect 7211 2801 7224 2853
rect 7276 2801 7289 2853
rect 7341 2815 7354 2853
rect 7406 2815 7419 2853
rect 7471 2815 7484 2853
rect 7536 2815 7573 2853
rect 7345 2801 7354 2815
rect 7417 2801 7419 2815
rect 5181 2785 5220 2801
rect 5254 2785 5293 2801
rect 5327 2785 5366 2801
rect 5400 2785 5439 2801
rect 5473 2785 5511 2801
rect 5545 2785 5583 2801
rect 5617 2785 5655 2801
rect 5689 2785 5727 2801
rect 5761 2785 5799 2801
rect 5833 2785 5871 2801
rect 5905 2785 5943 2801
rect 5977 2785 6015 2801
rect 6049 2785 6087 2801
rect 6121 2785 6159 2801
rect 6193 2785 6231 2801
rect 6265 2785 6303 2801
rect 6337 2785 6375 2801
rect 6409 2785 6447 2801
rect 6481 2785 6519 2801
rect 6553 2785 6591 2801
rect 6625 2785 6663 2801
rect 6697 2785 6735 2801
rect 6769 2785 6807 2801
rect 6841 2785 6879 2801
rect 6913 2785 6951 2801
rect 6985 2785 7023 2801
rect 7057 2785 7095 2801
rect 7129 2785 7167 2801
rect 7201 2785 7239 2801
rect 7273 2785 7311 2801
rect 7345 2785 7383 2801
rect 7417 2785 7455 2801
rect 7489 2785 7527 2801
rect 5181 2781 5204 2785
rect 1923 2737 5204 2781
rect 1923 2703 1935 2737
rect 1969 2703 2008 2737
rect 2042 2703 2081 2737
rect 2115 2703 2154 2737
rect 2188 2703 2227 2737
rect 2261 2703 2300 2737
rect 2334 2703 2373 2737
rect 2407 2703 2446 2737
rect 2480 2703 2519 2737
rect 2553 2703 2592 2737
rect 2626 2703 2665 2737
rect 2699 2703 2738 2737
rect 2772 2703 2811 2737
rect 2845 2703 2884 2737
rect 2918 2703 2957 2737
rect 2991 2703 3030 2737
rect 3064 2703 3103 2737
rect 3137 2703 3176 2737
rect 3210 2703 3249 2737
rect 3283 2703 3322 2737
rect 3356 2703 3395 2737
rect 3429 2703 3468 2737
rect 3502 2703 3541 2737
rect 3575 2703 3614 2737
rect 3648 2703 3687 2737
rect 3721 2703 3760 2737
rect 3794 2703 3833 2737
rect 3867 2703 3906 2737
rect 3940 2703 3979 2737
rect 4013 2703 4052 2737
rect 4086 2703 4125 2737
rect 4159 2703 4198 2737
rect 4232 2703 4271 2737
rect 4305 2703 4344 2737
rect 4378 2703 4417 2737
rect 4451 2703 4490 2737
rect 4524 2703 4563 2737
rect 4597 2703 4636 2737
rect 4670 2703 4709 2737
rect 4743 2703 4782 2737
rect 4816 2703 4855 2737
rect 4889 2703 4928 2737
rect 4962 2703 5001 2737
rect 5035 2703 5074 2737
rect 5108 2703 5147 2737
rect 5181 2733 5204 2737
rect 5256 2733 5270 2785
rect 5327 2781 5336 2785
rect 5400 2781 5402 2785
rect 5651 2781 5655 2785
rect 5716 2781 5727 2785
rect 5322 2737 5336 2781
rect 5388 2737 5402 2781
rect 5454 2737 5468 2781
rect 5520 2737 5534 2781
rect 5586 2737 5599 2781
rect 5651 2737 5664 2781
rect 5716 2737 5729 2781
rect 5327 2733 5336 2737
rect 5400 2733 5402 2737
rect 5651 2733 5655 2737
rect 5716 2733 5727 2737
rect 5781 2733 5794 2785
rect 5846 2733 5859 2785
rect 5911 2733 5924 2785
rect 5977 2781 5989 2785
rect 6049 2781 6054 2785
rect 6301 2781 6303 2785
rect 6366 2781 6375 2785
rect 5976 2737 5989 2781
rect 6041 2737 6054 2781
rect 6106 2737 6119 2781
rect 6171 2737 6184 2781
rect 6236 2737 6249 2781
rect 6301 2737 6314 2781
rect 6366 2737 6379 2781
rect 5977 2733 5989 2737
rect 6049 2733 6054 2737
rect 6301 2733 6303 2737
rect 6366 2733 6375 2737
rect 6431 2733 6444 2785
rect 6496 2733 6509 2785
rect 6561 2733 6574 2785
rect 6626 2733 6639 2785
rect 6697 2781 6704 2785
rect 7016 2781 7023 2785
rect 6691 2737 6704 2781
rect 6756 2737 6769 2781
rect 6821 2737 6834 2781
rect 6886 2737 6899 2781
rect 6951 2737 6964 2781
rect 7016 2737 7029 2781
rect 6697 2733 6704 2737
rect 7016 2733 7023 2737
rect 7081 2733 7094 2785
rect 7146 2733 7159 2785
rect 7211 2733 7224 2785
rect 7276 2733 7289 2785
rect 7345 2781 7354 2785
rect 7417 2781 7419 2785
rect 7561 2781 7573 2815
rect 7341 2737 7354 2781
rect 7406 2737 7419 2781
rect 7471 2737 7484 2781
rect 7536 2737 7573 2781
rect 7345 2733 7354 2737
rect 7417 2733 7419 2737
rect 5181 2717 5220 2733
rect 5254 2717 5293 2733
rect 5327 2717 5366 2733
rect 5400 2717 5439 2733
rect 5473 2717 5511 2733
rect 5545 2717 5583 2733
rect 5617 2717 5655 2733
rect 5689 2717 5727 2733
rect 5761 2717 5799 2733
rect 5833 2717 5871 2733
rect 5905 2717 5943 2733
rect 5977 2717 6015 2733
rect 6049 2717 6087 2733
rect 6121 2717 6159 2733
rect 6193 2717 6231 2733
rect 6265 2717 6303 2733
rect 6337 2717 6375 2733
rect 6409 2717 6447 2733
rect 6481 2717 6519 2733
rect 6553 2717 6591 2733
rect 6625 2717 6663 2733
rect 6697 2717 6735 2733
rect 6769 2717 6807 2733
rect 6841 2717 6879 2733
rect 6913 2717 6951 2733
rect 6985 2717 7023 2733
rect 7057 2717 7095 2733
rect 7129 2717 7167 2733
rect 7201 2717 7239 2733
rect 7273 2717 7311 2733
rect 7345 2717 7383 2733
rect 7417 2717 7455 2733
rect 7489 2717 7527 2733
rect 5181 2703 5204 2717
rect 1923 2665 5204 2703
rect 5256 2665 5270 2717
rect 5327 2703 5336 2717
rect 5400 2703 5402 2717
rect 5651 2703 5655 2717
rect 5716 2703 5727 2717
rect 5322 2665 5336 2703
rect 5388 2665 5402 2703
rect 5454 2665 5468 2703
rect 5520 2665 5534 2703
rect 5586 2665 5599 2703
rect 5651 2665 5664 2703
rect 5716 2665 5729 2703
rect 5781 2665 5794 2717
rect 5846 2665 5859 2717
rect 5911 2665 5924 2717
rect 5977 2703 5989 2717
rect 6049 2703 6054 2717
rect 6301 2703 6303 2717
rect 6366 2703 6375 2717
rect 5976 2665 5989 2703
rect 6041 2665 6054 2703
rect 6106 2665 6119 2703
rect 6171 2665 6184 2703
rect 6236 2665 6249 2703
rect 6301 2665 6314 2703
rect 6366 2665 6379 2703
rect 6431 2665 6444 2717
rect 6496 2665 6509 2717
rect 6561 2665 6574 2717
rect 6626 2665 6639 2717
rect 6697 2703 6704 2717
rect 7016 2703 7023 2717
rect 6691 2665 6704 2703
rect 6756 2665 6769 2703
rect 6821 2665 6834 2703
rect 6886 2665 6899 2703
rect 6951 2665 6964 2703
rect 7016 2665 7029 2703
rect 7081 2665 7094 2717
rect 7146 2665 7159 2717
rect 7211 2665 7224 2717
rect 7276 2665 7289 2717
rect 7345 2703 7354 2717
rect 7417 2703 7419 2717
rect 7561 2703 7573 2737
rect 7341 2665 7354 2703
rect 7406 2665 7419 2703
rect 7471 2665 7484 2703
rect 7536 2665 7573 2703
rect 1923 2659 7573 2665
rect 1923 2625 1935 2659
rect 1969 2625 2008 2659
rect 2042 2625 2081 2659
rect 2115 2625 2154 2659
rect 2188 2625 2227 2659
rect 2261 2625 2300 2659
rect 2334 2625 2373 2659
rect 2407 2625 2446 2659
rect 2480 2625 2519 2659
rect 2553 2625 2592 2659
rect 2626 2625 2665 2659
rect 2699 2625 2738 2659
rect 2772 2625 2811 2659
rect 2845 2625 2884 2659
rect 2918 2625 2957 2659
rect 2991 2625 3030 2659
rect 3064 2625 3103 2659
rect 3137 2625 3176 2659
rect 3210 2625 3249 2659
rect 3283 2625 3322 2659
rect 3356 2625 3395 2659
rect 3429 2625 3468 2659
rect 3502 2625 3541 2659
rect 3575 2625 3614 2659
rect 3648 2625 3687 2659
rect 3721 2625 3760 2659
rect 3794 2625 3833 2659
rect 3867 2625 3906 2659
rect 3940 2625 3979 2659
rect 4013 2625 4052 2659
rect 4086 2625 4125 2659
rect 4159 2625 4198 2659
rect 4232 2625 4271 2659
rect 4305 2625 4344 2659
rect 4378 2625 4417 2659
rect 4451 2625 4490 2659
rect 4524 2625 4563 2659
rect 4597 2625 4636 2659
rect 4670 2625 4709 2659
rect 4743 2625 4782 2659
rect 4816 2625 4855 2659
rect 4889 2625 4928 2659
rect 4962 2625 5001 2659
rect 5035 2625 5074 2659
rect 5108 2625 5147 2659
rect 5181 2649 5220 2659
rect 5254 2649 5293 2659
rect 5327 2649 5366 2659
rect 5400 2649 5439 2659
rect 5473 2649 5511 2659
rect 5545 2649 5583 2659
rect 5617 2649 5655 2659
rect 5689 2649 5727 2659
rect 5761 2649 5799 2659
rect 5833 2649 5871 2659
rect 5905 2649 5943 2659
rect 5977 2649 6015 2659
rect 6049 2649 6087 2659
rect 6121 2649 6159 2659
rect 6193 2649 6231 2659
rect 6265 2649 6303 2659
rect 6337 2649 6375 2659
rect 6409 2649 6447 2659
rect 6481 2649 6519 2659
rect 6553 2649 6591 2659
rect 6625 2649 6663 2659
rect 6697 2649 6735 2659
rect 6769 2649 6807 2659
rect 6841 2649 6879 2659
rect 6913 2649 6951 2659
rect 6985 2649 7023 2659
rect 7057 2649 7095 2659
rect 7129 2649 7167 2659
rect 7201 2649 7239 2659
rect 7273 2649 7311 2659
rect 7345 2649 7383 2659
rect 7417 2649 7455 2659
rect 7489 2649 7527 2659
rect 5181 2625 5204 2649
rect 1923 2597 5204 2625
rect 5256 2597 5270 2649
rect 5327 2625 5336 2649
rect 5400 2625 5402 2649
rect 5651 2625 5655 2649
rect 5716 2625 5727 2649
rect 5322 2597 5336 2625
rect 5388 2597 5402 2625
rect 5454 2597 5468 2625
rect 5520 2597 5534 2625
rect 5586 2597 5599 2625
rect 5651 2597 5664 2625
rect 5716 2597 5729 2625
rect 5781 2597 5794 2649
rect 5846 2597 5859 2649
rect 5911 2597 5924 2649
rect 5977 2625 5989 2649
rect 6049 2625 6054 2649
rect 6301 2625 6303 2649
rect 6366 2625 6375 2649
rect 5976 2597 5989 2625
rect 6041 2597 6054 2625
rect 6106 2597 6119 2625
rect 6171 2597 6184 2625
rect 6236 2597 6249 2625
rect 6301 2597 6314 2625
rect 6366 2597 6379 2625
rect 6431 2597 6444 2649
rect 6496 2597 6509 2649
rect 6561 2597 6574 2649
rect 6626 2597 6639 2649
rect 6697 2625 6704 2649
rect 7016 2625 7023 2649
rect 6691 2597 6704 2625
rect 6756 2597 6769 2625
rect 6821 2597 6834 2625
rect 6886 2597 6899 2625
rect 6951 2597 6964 2625
rect 7016 2597 7029 2625
rect 7081 2597 7094 2649
rect 7146 2597 7159 2649
rect 7211 2597 7224 2649
rect 7276 2597 7289 2649
rect 7345 2625 7354 2649
rect 7417 2625 7419 2649
rect 7561 2625 7573 2659
rect 7341 2597 7354 2625
rect 7406 2597 7419 2625
rect 7471 2597 7484 2625
rect 7536 2597 7573 2625
rect 1923 2581 7573 2597
rect 1923 2547 1935 2581
rect 1969 2547 2008 2581
rect 2042 2547 2081 2581
rect 2115 2547 2154 2581
rect 2188 2547 2227 2581
rect 2261 2547 2300 2581
rect 2334 2547 2373 2581
rect 2407 2547 2446 2581
rect 2480 2547 2519 2581
rect 2553 2547 2592 2581
rect 2626 2547 2665 2581
rect 2699 2547 2738 2581
rect 2772 2547 2811 2581
rect 2845 2547 2884 2581
rect 2918 2547 2957 2581
rect 2991 2547 3030 2581
rect 3064 2547 3103 2581
rect 3137 2547 3176 2581
rect 3210 2547 3249 2581
rect 3283 2547 3322 2581
rect 3356 2547 3395 2581
rect 3429 2547 3468 2581
rect 3502 2547 3541 2581
rect 3575 2547 3614 2581
rect 3648 2547 3687 2581
rect 3721 2547 3760 2581
rect 3794 2547 3833 2581
rect 3867 2547 3906 2581
rect 3940 2547 3979 2581
rect 4013 2547 4052 2581
rect 4086 2547 4125 2581
rect 4159 2547 4198 2581
rect 4232 2547 4271 2581
rect 4305 2547 4344 2581
rect 4378 2547 4417 2581
rect 4451 2547 4490 2581
rect 4524 2547 4563 2581
rect 4597 2547 4636 2581
rect 4670 2547 4709 2581
rect 4743 2547 4782 2581
rect 4816 2547 4855 2581
rect 4889 2547 4928 2581
rect 4962 2547 5001 2581
rect 5035 2547 5074 2581
rect 5108 2547 5147 2581
rect 5181 2547 5204 2581
rect 1923 2529 5204 2547
rect 5256 2529 5270 2581
rect 5327 2547 5336 2581
rect 5400 2547 5402 2581
rect 5651 2547 5655 2581
rect 5716 2547 5727 2581
rect 5322 2529 5336 2547
rect 5388 2529 5402 2547
rect 5454 2529 5468 2547
rect 5520 2529 5534 2547
rect 5586 2529 5599 2547
rect 5651 2529 5664 2547
rect 5716 2529 5729 2547
rect 5781 2529 5794 2581
rect 5846 2529 5859 2581
rect 5911 2529 5924 2581
rect 5977 2547 5989 2581
rect 6049 2547 6054 2581
rect 6301 2547 6303 2581
rect 6366 2547 6375 2581
rect 5976 2529 5989 2547
rect 6041 2529 6054 2547
rect 6106 2529 6119 2547
rect 6171 2529 6184 2547
rect 6236 2529 6249 2547
rect 6301 2529 6314 2547
rect 6366 2529 6379 2547
rect 6431 2529 6444 2581
rect 6496 2529 6509 2581
rect 6561 2529 6574 2581
rect 6626 2529 6639 2581
rect 6697 2547 6704 2581
rect 7016 2547 7023 2581
rect 6691 2529 6704 2547
rect 6756 2529 6769 2547
rect 6821 2529 6834 2547
rect 6886 2529 6899 2547
rect 6951 2529 6964 2547
rect 7016 2529 7029 2547
rect 7081 2529 7094 2581
rect 7146 2529 7159 2581
rect 7211 2529 7224 2581
rect 7276 2529 7289 2581
rect 7345 2547 7354 2581
rect 7417 2547 7419 2581
rect 7561 2547 7573 2581
rect 7341 2529 7354 2547
rect 7406 2529 7419 2547
rect 7471 2529 7484 2547
rect 7536 2529 7573 2547
rect 1923 2513 7573 2529
rect 1923 2503 5204 2513
rect 1923 2469 1935 2503
rect 1969 2469 2008 2503
rect 2042 2469 2081 2503
rect 2115 2469 2154 2503
rect 2188 2469 2227 2503
rect 2261 2469 2300 2503
rect 2334 2469 2373 2503
rect 2407 2469 2446 2503
rect 2480 2469 2519 2503
rect 2553 2469 2592 2503
rect 2626 2469 2665 2503
rect 2699 2469 2738 2503
rect 2772 2469 2811 2503
rect 2845 2469 2884 2503
rect 2918 2469 2957 2503
rect 2991 2469 3030 2503
rect 3064 2469 3103 2503
rect 3137 2469 3176 2503
rect 3210 2469 3249 2503
rect 3283 2469 3322 2503
rect 3356 2469 3395 2503
rect 3429 2469 3468 2503
rect 3502 2469 3541 2503
rect 3575 2469 3614 2503
rect 3648 2469 3687 2503
rect 3721 2469 3760 2503
rect 3794 2469 3833 2503
rect 3867 2469 3906 2503
rect 3940 2469 3979 2503
rect 4013 2469 4052 2503
rect 4086 2469 4125 2503
rect 4159 2469 4198 2503
rect 4232 2469 4271 2503
rect 4305 2469 4344 2503
rect 4378 2469 4417 2503
rect 4451 2469 4490 2503
rect 4524 2469 4563 2503
rect 4597 2469 4636 2503
rect 4670 2469 4709 2503
rect 4743 2469 4782 2503
rect 4816 2469 4855 2503
rect 4889 2469 4928 2503
rect 4962 2469 5001 2503
rect 5035 2469 5074 2503
rect 5108 2469 5147 2503
rect 5181 2469 5204 2503
rect 1923 2461 5204 2469
rect 5256 2461 5270 2513
rect 5322 2503 5336 2513
rect 5388 2503 5402 2513
rect 5454 2503 5468 2513
rect 5520 2503 5534 2513
rect 5586 2503 5599 2513
rect 5651 2503 5664 2513
rect 5716 2503 5729 2513
rect 5327 2469 5336 2503
rect 5400 2469 5402 2503
rect 5651 2469 5655 2503
rect 5716 2469 5727 2503
rect 5322 2461 5336 2469
rect 5388 2461 5402 2469
rect 5454 2461 5468 2469
rect 5520 2461 5534 2469
rect 5586 2461 5599 2469
rect 5651 2461 5664 2469
rect 5716 2461 5729 2469
rect 5781 2461 5794 2513
rect 5846 2461 5859 2513
rect 5911 2461 5924 2513
rect 5976 2503 5989 2513
rect 6041 2503 6054 2513
rect 6106 2503 6119 2513
rect 6171 2503 6184 2513
rect 6236 2503 6249 2513
rect 6301 2503 6314 2513
rect 6366 2503 6379 2513
rect 5977 2469 5989 2503
rect 6049 2469 6054 2503
rect 6301 2469 6303 2503
rect 6366 2469 6375 2503
rect 5976 2461 5989 2469
rect 6041 2461 6054 2469
rect 6106 2461 6119 2469
rect 6171 2461 6184 2469
rect 6236 2461 6249 2469
rect 6301 2461 6314 2469
rect 6366 2461 6379 2469
rect 6431 2461 6444 2513
rect 6496 2461 6509 2513
rect 6561 2461 6574 2513
rect 6626 2461 6639 2513
rect 6691 2503 6704 2513
rect 6756 2503 6769 2513
rect 6821 2503 6834 2513
rect 6886 2503 6899 2513
rect 6951 2503 6964 2513
rect 7016 2503 7029 2513
rect 6697 2469 6704 2503
rect 7016 2469 7023 2503
rect 6691 2461 6704 2469
rect 6756 2461 6769 2469
rect 6821 2461 6834 2469
rect 6886 2461 6899 2469
rect 6951 2461 6964 2469
rect 7016 2461 7029 2469
rect 7081 2461 7094 2513
rect 7146 2461 7159 2513
rect 7211 2461 7224 2513
rect 7276 2461 7289 2513
rect 7341 2503 7354 2513
rect 7406 2503 7419 2513
rect 7471 2503 7484 2513
rect 7536 2503 7573 2513
rect 7345 2469 7354 2503
rect 7417 2469 7419 2503
rect 7561 2469 7573 2503
rect 7341 2461 7354 2469
rect 7406 2461 7419 2469
rect 7471 2461 7484 2469
rect 7536 2461 7573 2469
rect 1923 2460 7573 2461
tri 5230 2284 5406 2460 ne
rect 5406 2269 7573 2460
rect 2241 2263 5172 2267
rect 2241 2211 3192 2263
rect 3244 2211 3258 2263
rect 3310 2211 3324 2263
rect 3376 2211 3390 2263
rect 3442 2211 3456 2263
rect 3508 2211 3522 2263
rect 3574 2211 3588 2263
rect 3640 2211 3654 2263
rect 3706 2211 3720 2263
rect 3772 2211 3786 2263
rect 3838 2211 3852 2263
rect 3904 2211 3918 2263
rect 3970 2211 3984 2263
rect 4036 2211 4050 2263
rect 4102 2211 4116 2263
rect 4168 2211 4182 2263
rect 4234 2211 4248 2263
rect 4300 2211 4314 2263
rect 4366 2211 4380 2263
rect 4432 2211 4446 2263
rect 4498 2211 4512 2263
rect 4564 2211 4578 2263
rect 4630 2211 4644 2263
rect 4696 2211 4710 2263
rect 4762 2211 4776 2263
rect 4828 2211 4841 2263
rect 4893 2211 5172 2263
rect 2241 2197 5172 2211
tri 1942 2121 1971 2150 se
rect 1971 2121 1977 2150
tri 1908 2087 1942 2121 se
rect 1942 2098 1977 2121
rect 2029 2098 2042 2150
rect 2094 2098 2107 2150
rect 2159 2098 2165 2150
rect 1942 2087 2165 2098
tri 1878 2057 1908 2087 se
rect 1908 2067 2165 2087
rect 2241 2145 3192 2197
rect 3244 2145 3258 2197
rect 3310 2145 3324 2197
rect 3376 2145 3390 2197
rect 3442 2145 3456 2197
rect 3508 2145 3522 2197
rect 3574 2145 3588 2197
rect 3640 2145 3654 2197
rect 3706 2145 3720 2197
rect 3772 2145 3786 2197
rect 3838 2145 3852 2197
rect 3904 2145 3918 2197
rect 3970 2145 3984 2197
rect 4036 2145 4050 2197
rect 4102 2145 4116 2197
rect 4168 2145 4182 2197
rect 4234 2145 4248 2197
rect 4300 2145 4314 2197
rect 4366 2145 4380 2197
rect 4432 2145 4446 2197
rect 4498 2145 4512 2197
rect 4564 2145 4578 2197
rect 4630 2145 4644 2197
rect 4696 2145 4710 2197
rect 4762 2145 4776 2197
rect 4828 2145 4841 2197
rect 4893 2145 5172 2197
rect 2241 2131 5172 2145
rect 2241 2079 3192 2131
rect 3244 2079 3258 2131
rect 3310 2079 3324 2131
rect 3376 2079 3390 2131
rect 3442 2079 3456 2131
rect 3508 2079 3522 2131
rect 3574 2079 3588 2131
rect 3640 2079 3654 2131
rect 3706 2079 3720 2131
rect 3772 2079 3786 2131
rect 3838 2079 3852 2131
rect 3904 2079 3918 2131
rect 3970 2079 3984 2131
rect 4036 2079 4050 2131
rect 4102 2079 4116 2131
rect 4168 2079 4182 2131
rect 4234 2079 4248 2131
rect 4300 2079 4314 2131
rect 4366 2079 4380 2131
rect 4432 2079 4446 2131
rect 4498 2079 4512 2131
rect 4564 2079 4578 2131
rect 4630 2079 4644 2131
rect 4696 2079 4710 2131
rect 4762 2079 4776 2131
rect 4828 2079 4841 2131
rect 4893 2079 5172 2131
rect 1908 2057 1992 2067
tri 1992 2057 2002 2067 nw
rect 2241 2065 5172 2079
rect 1878 2047 1982 2057
tri 1982 2047 1992 2057 nw
rect 1878 1860 1959 2047
tri 1959 2024 1982 2047 nw
rect 2241 2016 3192 2065
rect 2241 1982 2253 2016
rect 2287 1982 2326 2016
rect 2360 1982 2399 2016
rect 2433 1982 2472 2016
rect 2506 1982 2545 2016
rect 2579 1982 2618 2016
rect 2652 1982 2691 2016
rect 2725 1982 2764 2016
rect 2798 1982 2837 2016
rect 2871 1982 2910 2016
rect 2944 1982 2983 2016
rect 3017 1982 3056 2016
rect 3090 1982 3129 2016
rect 3163 2013 3192 2016
rect 3244 2013 3258 2065
rect 3310 2013 3324 2065
rect 3376 2016 3390 2065
rect 3442 2016 3456 2065
rect 3508 2016 3522 2065
rect 3574 2016 3588 2065
rect 3640 2016 3654 2065
rect 3706 2016 3720 2065
rect 3772 2016 3786 2065
rect 3382 2013 3390 2016
rect 3455 2013 3456 2016
rect 3706 2013 3709 2016
rect 3772 2013 3781 2016
rect 3838 2013 3852 2065
rect 3904 2013 3918 2065
rect 3970 2013 3984 2065
rect 4036 2013 4050 2065
rect 4102 2016 4116 2065
rect 4168 2016 4182 2065
rect 4234 2016 4248 2065
rect 4300 2016 4314 2065
rect 4366 2016 4380 2065
rect 4432 2016 4446 2065
rect 4498 2016 4512 2065
rect 4564 2016 4578 2065
rect 4103 2013 4116 2016
rect 4175 2013 4182 2016
rect 4247 2013 4248 2016
rect 4498 2013 4501 2016
rect 4564 2013 4573 2016
rect 4630 2013 4644 2065
rect 4696 2013 4710 2065
rect 4762 2013 4776 2065
rect 4828 2013 4841 2065
rect 4893 2016 5172 2065
rect 3163 1999 3202 2013
rect 3236 1999 3275 2013
rect 3309 1999 3348 2013
rect 3382 1999 3421 2013
rect 3455 1999 3493 2013
rect 3527 1999 3565 2013
rect 3599 1999 3637 2013
rect 3671 1999 3709 2013
rect 3743 1999 3781 2013
rect 3815 1999 3853 2013
rect 3887 1999 3925 2013
rect 3959 1999 3997 2013
rect 4031 1999 4069 2013
rect 4103 1999 4141 2013
rect 4175 1999 4213 2013
rect 4247 1999 4285 2013
rect 4319 1999 4357 2013
rect 4391 1999 4429 2013
rect 4463 1999 4501 2013
rect 4535 1999 4573 2013
rect 4607 1999 4645 2013
rect 4679 1999 4717 2013
rect 4751 1999 4789 2013
rect 4823 1999 4861 2013
rect 3163 1982 3192 1999
tri 2228 1944 2241 1957 se
rect 2241 1947 3192 1982
rect 3244 1947 3258 1999
rect 3310 1947 3324 1999
rect 3382 1982 3390 1999
rect 3455 1982 3456 1999
rect 3706 1982 3709 1999
rect 3772 1982 3781 1999
rect 3376 1947 3390 1982
rect 3442 1947 3456 1982
rect 3508 1947 3522 1982
rect 3574 1947 3588 1982
rect 3640 1947 3654 1982
rect 3706 1947 3720 1982
rect 3772 1947 3786 1982
rect 3838 1947 3852 1999
rect 3904 1947 3918 1999
rect 3970 1947 3984 1999
rect 4036 1947 4050 1999
rect 4103 1982 4116 1999
rect 4175 1982 4182 1999
rect 4247 1982 4248 1999
rect 4498 1982 4501 1999
rect 4564 1982 4573 1999
rect 4102 1947 4116 1982
rect 4168 1947 4182 1982
rect 4234 1947 4248 1982
rect 4300 1947 4314 1982
rect 4366 1947 4380 1982
rect 4432 1947 4446 1982
rect 4498 1947 4512 1982
rect 4564 1947 4578 1982
rect 4630 1947 4644 1999
rect 4696 1947 4710 1999
rect 4762 1947 4776 1999
rect 4828 1947 4841 1999
rect 4895 1982 4933 2016
rect 4967 1982 5172 2016
rect 4893 1947 5172 1982
rect 2241 1944 5172 1947
tri 2207 1923 2228 1944 se
rect 2228 1933 5005 1944
rect 2228 1923 3192 1933
rect 1997 1917 3192 1923
rect 1997 1883 2009 1917
rect 2043 1883 2084 1917
rect 2118 1883 2159 1917
rect 2193 1883 2234 1917
rect 2268 1883 2309 1917
rect 2343 1883 2384 1917
rect 2418 1883 2459 1917
rect 2493 1883 2534 1917
rect 2568 1883 2609 1917
rect 2643 1883 2684 1917
rect 2718 1883 2759 1917
rect 2793 1883 2834 1917
rect 2868 1883 2909 1917
rect 2943 1883 2984 1917
rect 3018 1883 3059 1917
rect 3093 1883 3133 1917
rect 3167 1883 3192 1917
rect 1997 1881 3192 1883
rect 3244 1881 3258 1933
rect 3310 1917 3324 1933
rect 3376 1917 3390 1933
rect 3315 1883 3324 1917
rect 3389 1883 3390 1917
rect 3310 1881 3324 1883
rect 3376 1881 3390 1883
rect 3442 1881 3456 1933
rect 3508 1881 3522 1933
rect 3574 1881 3588 1933
rect 3640 1917 3654 1933
rect 3706 1917 3720 1933
rect 3772 1917 3786 1933
rect 3838 1917 3852 1933
rect 3904 1917 3918 1933
rect 3648 1883 3654 1917
rect 3838 1883 3839 1917
rect 3904 1883 3914 1917
rect 3640 1881 3654 1883
rect 3706 1881 3720 1883
rect 3772 1881 3786 1883
rect 3838 1881 3852 1883
rect 3904 1881 3918 1883
rect 3970 1881 3984 1933
rect 4036 1881 4050 1933
rect 4102 1881 4116 1933
rect 4168 1917 4182 1933
rect 4234 1917 4248 1933
rect 4300 1917 4314 1933
rect 4366 1917 4380 1933
rect 4432 1917 4446 1933
rect 4173 1883 4182 1917
rect 4432 1883 4439 1917
rect 4168 1881 4182 1883
rect 4234 1881 4248 1883
rect 4300 1881 4314 1883
rect 4366 1881 4380 1883
rect 4432 1881 4446 1883
rect 4498 1881 4512 1933
rect 4564 1881 4578 1933
rect 4630 1881 4644 1933
rect 4696 1917 4710 1933
rect 4762 1917 4776 1933
rect 4828 1917 4841 1933
rect 4893 1917 5005 1933
rect 4697 1883 4710 1917
rect 4771 1883 4776 1917
rect 4919 1910 5005 1917
rect 5039 1910 5172 1944
rect 4919 1883 5172 1910
rect 4696 1881 4710 1883
rect 4762 1881 4776 1883
rect 4828 1881 4841 1883
rect 4893 1881 5172 1883
rect 1997 1877 5172 1881
tri 4727 1869 4735 1877 ne
rect 4735 1869 5172 1877
rect 1878 1826 1919 1860
rect 1953 1826 1959 1860
tri 4735 1843 4761 1869 ne
rect 4761 1835 5005 1869
rect 5039 1835 5172 1869
rect 1878 1787 1959 1826
rect 1878 1753 1919 1787
rect 1953 1753 1959 1787
rect 2083 1825 2798 1834
rect 2850 1825 2891 1834
rect 2943 1825 2983 1834
rect 3035 1825 4697 1834
rect 2083 1791 2095 1825
rect 2129 1791 2170 1825
rect 2204 1791 2245 1825
rect 2279 1791 2319 1825
rect 2353 1791 2393 1825
rect 2427 1791 2467 1825
rect 2501 1791 2541 1825
rect 2575 1791 2615 1825
rect 2649 1791 2689 1825
rect 2723 1791 2763 1825
rect 2797 1791 2798 1825
rect 2871 1791 2891 1825
rect 2945 1791 2983 1825
rect 3035 1791 3059 1825
rect 3093 1791 3133 1825
rect 3167 1791 3207 1825
rect 3241 1791 3281 1825
rect 3315 1791 3355 1825
rect 3389 1791 3625 1825
rect 3659 1791 3699 1825
rect 3733 1791 3773 1825
rect 3807 1791 3847 1825
rect 3881 1791 3921 1825
rect 3955 1791 3994 1825
rect 4028 1791 4067 1825
rect 4101 1791 4140 1825
rect 4174 1791 4213 1825
rect 4247 1791 4286 1825
rect 4320 1791 4359 1825
rect 4393 1791 4432 1825
rect 4466 1791 4505 1825
rect 4539 1791 4578 1825
rect 4612 1791 4651 1825
rect 4685 1791 4697 1825
rect 2083 1782 2798 1791
rect 2850 1782 2891 1791
rect 2943 1782 2983 1791
rect 3035 1782 4697 1791
rect 4761 1794 5172 1835
tri 4748 1760 4761 1773 se
rect 4761 1760 5005 1794
rect 5039 1760 5172 1794
rect 1878 1714 1959 1753
tri 4739 1751 4748 1760 se
rect 4748 1751 5172 1760
tri 4727 1739 4739 1751 se
rect 4739 1739 5172 1751
rect 1878 1680 1919 1714
rect 1953 1680 1959 1714
rect 2229 1733 5172 1739
rect 2229 1699 2241 1733
rect 2275 1699 2316 1733
rect 2350 1699 2391 1733
rect 2425 1699 2466 1733
rect 2500 1699 2541 1733
rect 2575 1699 2615 1733
rect 2649 1699 2689 1733
rect 2723 1699 2763 1733
rect 2797 1699 2837 1733
rect 2871 1699 2911 1733
rect 2945 1699 2985 1733
rect 3019 1699 3059 1733
rect 3093 1699 3133 1733
rect 3167 1699 3207 1733
rect 3241 1699 3281 1733
rect 3315 1699 3355 1733
rect 3389 1699 3539 1733
rect 3573 1699 3614 1733
rect 3648 1699 3689 1733
rect 3723 1699 3764 1733
rect 3798 1699 3839 1733
rect 3873 1699 3914 1733
rect 3948 1699 3989 1733
rect 4023 1699 4064 1733
rect 4098 1699 4139 1733
rect 4173 1699 4214 1733
rect 4248 1699 4289 1733
rect 4323 1699 4364 1733
rect 4398 1699 4439 1733
rect 4473 1699 4514 1733
rect 4548 1699 4589 1733
rect 4623 1699 4663 1733
rect 4697 1699 4737 1733
rect 4771 1699 4811 1733
rect 4845 1699 4885 1733
rect 4919 1719 5172 1733
rect 4919 1699 5005 1719
rect 2229 1693 5005 1699
tri 4727 1685 4735 1693 ne
rect 4735 1685 5005 1693
rect 5039 1685 5172 1719
rect 1878 1641 1959 1680
tri 4735 1676 4744 1685 ne
rect 4744 1676 5172 1685
tri 4744 1659 4761 1676 ne
rect 1878 1607 1919 1641
rect 1953 1607 1959 1641
rect 1878 1568 1959 1607
rect 2083 1641 2798 1650
rect 2850 1641 2891 1650
rect 2943 1641 2983 1650
rect 3035 1641 4697 1650
rect 2083 1607 2095 1641
rect 2129 1607 2170 1641
rect 2204 1607 2245 1641
rect 2279 1607 2319 1641
rect 2353 1607 2393 1641
rect 2427 1607 2467 1641
rect 2501 1607 2541 1641
rect 2575 1607 2615 1641
rect 2649 1607 2689 1641
rect 2723 1607 2763 1641
rect 2797 1607 2798 1641
rect 2871 1607 2891 1641
rect 2945 1607 2983 1641
rect 3035 1607 3059 1641
rect 3093 1607 3133 1641
rect 3167 1607 3207 1641
rect 3241 1607 3281 1641
rect 3315 1607 3355 1641
rect 3389 1607 3625 1641
rect 3659 1607 3699 1641
rect 3733 1607 3773 1641
rect 3807 1607 3847 1641
rect 3881 1607 3921 1641
rect 3955 1607 3994 1641
rect 4028 1607 4067 1641
rect 4101 1607 4140 1641
rect 4174 1607 4213 1641
rect 4247 1607 4286 1641
rect 4320 1607 4359 1641
rect 4393 1607 4432 1641
rect 4466 1607 4505 1641
rect 4539 1607 4578 1641
rect 4612 1607 4651 1641
rect 4685 1607 4697 1641
rect 2083 1598 2798 1607
rect 2850 1598 2891 1607
rect 2943 1598 2983 1607
rect 3035 1598 4697 1607
rect 4761 1644 5172 1676
rect 4761 1610 5005 1644
rect 5039 1610 5172 1644
tri 4741 1569 4761 1589 se
rect 4761 1569 5172 1610
rect 1878 1534 1919 1568
rect 1953 1534 1959 1568
tri 4727 1555 4741 1569 se
rect 4741 1555 5005 1569
rect 1878 1495 1959 1534
rect 2229 1549 5005 1555
rect 2229 1515 2241 1549
rect 2275 1515 2316 1549
rect 2350 1515 2391 1549
rect 2425 1515 2466 1549
rect 2500 1515 2541 1549
rect 2575 1515 2615 1549
rect 2649 1515 2689 1549
rect 2723 1515 2763 1549
rect 2797 1515 2837 1549
rect 2871 1515 2911 1549
rect 2945 1515 2985 1549
rect 3019 1515 3059 1549
rect 3093 1515 3133 1549
rect 3167 1515 3207 1549
rect 3241 1515 3281 1549
rect 3315 1515 3355 1549
rect 3389 1515 3539 1549
rect 3573 1515 3614 1549
rect 3648 1515 3689 1549
rect 3723 1515 3764 1549
rect 3798 1515 3839 1549
rect 3873 1515 3914 1549
rect 3948 1515 3989 1549
rect 4023 1515 4064 1549
rect 4098 1515 4139 1549
rect 4173 1515 4214 1549
rect 4248 1515 4289 1549
rect 4323 1515 4364 1549
rect 4398 1515 4439 1549
rect 4473 1515 4514 1549
rect 4548 1515 4589 1549
rect 4623 1515 4663 1549
rect 4697 1515 4737 1549
rect 4771 1515 4811 1549
rect 4845 1515 4885 1549
rect 4919 1535 5005 1549
rect 5039 1535 5172 1569
rect 4919 1515 5172 1535
rect 2229 1509 5172 1515
rect 1878 1461 1919 1495
rect 1953 1461 1959 1495
tri 4727 1494 4742 1509 ne
rect 4742 1494 5172 1509
tri 4742 1475 4761 1494 ne
rect 1878 1422 1959 1461
rect 1878 1388 1919 1422
rect 1953 1388 1959 1422
rect 2083 1457 2798 1467
rect 2850 1457 2891 1467
rect 2943 1457 2983 1467
rect 3035 1457 4697 1467
rect 2083 1423 2095 1457
rect 2129 1423 2170 1457
rect 2204 1423 2245 1457
rect 2279 1423 2319 1457
rect 2353 1423 2393 1457
rect 2427 1423 2467 1457
rect 2501 1423 2541 1457
rect 2575 1423 2615 1457
rect 2649 1423 2689 1457
rect 2723 1423 2763 1457
rect 2797 1423 2798 1457
rect 2871 1423 2891 1457
rect 2945 1423 2983 1457
rect 3035 1423 3059 1457
rect 3093 1423 3133 1457
rect 3167 1423 3207 1457
rect 3241 1423 3281 1457
rect 3315 1423 3355 1457
rect 3389 1423 3625 1457
rect 3659 1423 3699 1457
rect 3733 1423 3773 1457
rect 3807 1423 3847 1457
rect 3881 1423 3921 1457
rect 3955 1423 3994 1457
rect 4028 1423 4067 1457
rect 4101 1423 4140 1457
rect 4174 1423 4213 1457
rect 4247 1423 4286 1457
rect 4320 1423 4359 1457
rect 4393 1423 4432 1457
rect 4466 1423 4505 1457
rect 4539 1423 4578 1457
rect 4612 1423 4651 1457
rect 4685 1423 4697 1457
rect 2083 1415 2798 1423
rect 2850 1415 2891 1423
rect 2943 1415 2983 1423
rect 3035 1415 4697 1423
rect 4761 1460 5005 1494
rect 5039 1460 5172 1494
rect 4761 1419 5172 1460
rect 1878 1349 1959 1388
tri 4741 1385 4761 1405 se
rect 4761 1385 5005 1419
rect 5039 1385 5172 1419
tri 4732 1376 4741 1385 se
rect 4741 1376 5172 1385
tri 4727 1371 4732 1376 se
rect 4732 1371 5172 1376
rect 1878 1315 1919 1349
rect 1953 1315 1959 1349
rect 2229 1365 5172 1371
rect 2229 1331 2241 1365
rect 2275 1331 2316 1365
rect 2350 1331 2391 1365
rect 2425 1331 2466 1365
rect 2500 1331 2541 1365
rect 2575 1331 2615 1365
rect 2649 1331 2689 1365
rect 2723 1331 2763 1365
rect 2797 1331 2837 1365
rect 2871 1331 2911 1365
rect 2945 1331 2985 1365
rect 3019 1331 3059 1365
rect 3093 1331 3133 1365
rect 3167 1331 3207 1365
rect 3241 1331 3281 1365
rect 3315 1331 3355 1365
rect 3389 1331 3539 1365
rect 3573 1331 3614 1365
rect 3648 1331 3689 1365
rect 3723 1331 3764 1365
rect 3798 1331 3839 1365
rect 3873 1331 3914 1365
rect 3948 1331 3989 1365
rect 4023 1331 4064 1365
rect 4098 1331 4139 1365
rect 4173 1331 4214 1365
rect 4248 1331 4289 1365
rect 4323 1331 4364 1365
rect 4398 1331 4439 1365
rect 4473 1331 4514 1365
rect 4548 1331 4589 1365
rect 4623 1331 4663 1365
rect 4697 1331 4737 1365
rect 4771 1331 4811 1365
rect 4845 1331 4885 1365
rect 4919 1344 5172 1365
rect 4919 1331 5005 1344
rect 2229 1325 5005 1331
rect 1878 1276 1959 1315
tri 4727 1310 4742 1325 ne
rect 4742 1310 5005 1325
rect 5039 1310 5172 1344
tri 4742 1301 4751 1310 ne
rect 4751 1301 5172 1310
tri 4751 1291 4761 1301 ne
rect 1878 1242 1919 1276
rect 1953 1242 1959 1276
rect 1878 1202 1959 1242
rect 2083 1273 2798 1282
rect 2850 1273 2891 1282
rect 2943 1273 2983 1282
rect 3035 1273 4697 1282
rect 2083 1239 2095 1273
rect 2129 1239 2170 1273
rect 2204 1239 2245 1273
rect 2279 1239 2319 1273
rect 2353 1239 2393 1273
rect 2427 1239 2467 1273
rect 2501 1239 2541 1273
rect 2575 1239 2615 1273
rect 2649 1239 2689 1273
rect 2723 1239 2763 1273
rect 2797 1239 2798 1273
rect 2871 1239 2891 1273
rect 2945 1239 2983 1273
rect 3035 1239 3059 1273
rect 3093 1239 3133 1273
rect 3167 1239 3207 1273
rect 3241 1239 3281 1273
rect 3315 1239 3355 1273
rect 3389 1239 3625 1273
rect 3659 1239 3699 1273
rect 3733 1239 3773 1273
rect 3807 1239 3847 1273
rect 3881 1239 3921 1273
rect 3955 1239 3994 1273
rect 4028 1239 4067 1273
rect 4101 1239 4140 1273
rect 4174 1239 4213 1273
rect 4247 1239 4286 1273
rect 4320 1239 4359 1273
rect 4393 1239 4432 1273
rect 4466 1239 4505 1273
rect 4539 1239 4578 1273
rect 4612 1239 4651 1273
rect 4685 1239 4697 1273
rect 2083 1230 2798 1239
rect 2850 1230 2891 1239
rect 2943 1230 2983 1239
rect 3035 1230 4697 1239
rect 4761 1270 5172 1301
rect 4761 1236 5005 1270
rect 5039 1236 5172 1270
rect 1878 1168 1919 1202
rect 1953 1168 1959 1202
tri 4736 1196 4761 1221 se
rect 4761 1196 5172 1236
tri 4727 1187 4736 1196 se
rect 4736 1187 5005 1196
rect 1878 1128 1959 1168
rect 2229 1181 5005 1187
rect 2229 1147 2241 1181
rect 2275 1147 2316 1181
rect 2350 1147 2391 1181
rect 2425 1147 2466 1181
rect 2500 1147 2541 1181
rect 2575 1147 2615 1181
rect 2649 1147 2689 1181
rect 2723 1147 2763 1181
rect 2797 1147 2837 1181
rect 2871 1147 2911 1181
rect 2945 1147 2985 1181
rect 3019 1147 3059 1181
rect 3093 1147 3133 1181
rect 3167 1147 3207 1181
rect 3241 1147 3281 1181
rect 3315 1147 3355 1181
rect 3389 1147 3539 1181
rect 3573 1147 3614 1181
rect 3648 1147 3689 1181
rect 3723 1147 3764 1181
rect 3798 1147 3839 1181
rect 3873 1147 3914 1181
rect 3948 1147 3989 1181
rect 4023 1147 4064 1181
rect 4098 1147 4139 1181
rect 4173 1147 4214 1181
rect 4248 1147 4289 1181
rect 4323 1147 4364 1181
rect 4398 1147 4439 1181
rect 4473 1147 4514 1181
rect 4548 1147 4589 1181
rect 4623 1147 4663 1181
rect 4697 1147 4737 1181
rect 4771 1147 4811 1181
rect 4845 1147 4885 1181
rect 4919 1162 5005 1181
rect 5039 1162 5172 1196
rect 4919 1147 5172 1162
rect 2229 1141 5172 1147
rect 1878 1094 1919 1128
rect 1953 1094 1959 1128
tri 4727 1122 4746 1141 ne
rect 4746 1122 5172 1141
tri 4746 1107 4761 1122 ne
rect 1878 1054 1959 1094
rect 1878 1020 1919 1054
rect 1953 1020 1959 1054
rect 2083 1089 2798 1098
rect 2850 1089 2891 1098
rect 2943 1089 2983 1098
rect 3035 1089 4697 1098
rect 2083 1055 2095 1089
rect 2129 1055 2170 1089
rect 2204 1055 2245 1089
rect 2279 1055 2319 1089
rect 2353 1055 2393 1089
rect 2427 1055 2467 1089
rect 2501 1055 2541 1089
rect 2575 1055 2615 1089
rect 2649 1055 2689 1089
rect 2723 1055 2763 1089
rect 2797 1055 2798 1089
rect 2871 1055 2891 1089
rect 2945 1055 2983 1089
rect 3035 1055 3059 1089
rect 3093 1055 3133 1089
rect 3167 1055 3207 1089
rect 3241 1055 3281 1089
rect 3315 1055 3355 1089
rect 3389 1055 3625 1089
rect 3659 1055 3699 1089
rect 3733 1055 3773 1089
rect 3807 1055 3847 1089
rect 3881 1055 3921 1089
rect 3955 1055 3994 1089
rect 4028 1055 4067 1089
rect 4101 1055 4140 1089
rect 4174 1055 4213 1089
rect 4247 1055 4286 1089
rect 4320 1055 4359 1089
rect 4393 1055 4432 1089
rect 4466 1055 4505 1089
rect 4539 1055 4578 1089
rect 4612 1055 4651 1089
rect 4685 1055 4697 1089
rect 2083 1046 2798 1055
rect 2850 1046 2891 1055
rect 2943 1046 2983 1055
rect 3035 1046 4697 1055
rect 4761 1088 5005 1122
rect 5039 1088 5172 1122
tri 1852 517 1878 543 se
rect 1878 517 1959 1020
tri 4727 1003 4761 1037 se
rect 4761 1003 5172 1088
rect 2229 998 5172 1003
rect 2229 997 5005 998
rect 2229 963 2241 997
rect 2275 963 2316 997
rect 2350 963 2391 997
rect 2425 963 2466 997
rect 2500 963 2541 997
rect 2575 963 2615 997
rect 2649 963 2689 997
rect 2723 963 2763 997
rect 2797 963 2837 997
rect 2871 963 2911 997
rect 2945 963 2985 997
rect 3019 963 3059 997
rect 3093 963 3133 997
rect 3167 963 3207 997
rect 3241 963 3281 997
rect 3315 963 3355 997
rect 3389 963 3539 997
rect 3573 963 3614 997
rect 3648 963 3689 997
rect 3723 963 3764 997
rect 3798 963 3839 997
rect 3873 963 3914 997
rect 3948 963 3989 997
rect 4023 963 4064 997
rect 4098 963 4139 997
rect 4173 963 4214 997
rect 4248 963 4289 997
rect 4323 963 4364 997
rect 4398 963 4439 997
rect 4473 963 4514 997
rect 4548 963 4589 997
rect 4623 963 4663 997
rect 4697 963 4737 997
rect 4771 963 4811 997
rect 4845 963 4885 997
rect 4919 964 5005 997
rect 5039 964 5172 998
rect 4919 963 5172 964
tri 2198 926 2229 957 se
rect 2229 926 5172 963
tri 2170 898 2198 926 se
rect 2198 898 5172 926
tri 2136 864 2170 898 se
rect 2170 864 2471 898
rect 2505 864 2543 898
rect 2577 864 2615 898
rect 2649 864 2687 898
rect 2721 864 2759 898
rect 2793 864 2831 898
rect 2865 864 2903 898
rect 2937 864 2975 898
rect 3009 864 3047 898
rect 3081 864 3119 898
rect 3153 864 3191 898
rect 3225 864 3263 898
rect 3297 864 3335 898
rect 3369 864 3407 898
rect 3441 864 3479 898
rect 3513 864 3551 898
rect 3585 864 3623 898
rect 3657 864 3695 898
rect 3729 864 3767 898
rect 3801 864 3839 898
rect 3873 864 3911 898
rect 3945 864 3984 898
rect 4018 864 4057 898
rect 4091 864 4130 898
rect 4164 864 4203 898
rect 4237 864 4276 898
rect 4310 864 4349 898
rect 4383 864 4422 898
rect 4456 864 4495 898
rect 4529 864 4568 898
rect 4602 864 4641 898
rect 4675 864 4714 898
rect 4748 864 4787 898
rect 4821 864 4860 898
rect 4894 864 4933 898
rect 4967 864 5172 898
tri 2123 851 2136 864 se
rect 2136 858 5172 864
rect 5406 2235 5414 2269
rect 5448 2235 5486 2269
rect 5520 2235 5558 2269
rect 5592 2235 5630 2269
rect 5664 2235 5702 2269
rect 5736 2235 5774 2269
rect 5808 2235 5846 2269
rect 5880 2235 5918 2269
rect 5952 2235 5990 2269
rect 6024 2235 6062 2269
rect 6096 2235 6134 2269
rect 6168 2235 6206 2269
rect 6240 2235 6278 2269
rect 6312 2235 6350 2269
rect 6384 2235 6595 2269
rect 6629 2242 6667 2269
rect 6663 2235 6667 2242
rect 6701 2242 6739 2269
rect 6701 2235 6711 2242
rect 6773 2235 6811 2269
rect 6845 2242 6883 2269
rect 6917 2242 6955 2269
rect 6989 2242 7027 2269
rect 7061 2242 7099 2269
rect 7133 2242 7171 2269
rect 6863 2235 6883 2242
rect 6989 2235 7011 2242
rect 7063 2235 7099 2242
rect 7163 2235 7171 2242
rect 7205 2242 7243 2269
rect 7277 2242 7315 2269
rect 7349 2242 7387 2269
rect 7205 2235 7211 2242
rect 7277 2235 7311 2242
rect 7363 2235 7387 2242
rect 7421 2235 7459 2269
rect 7493 2235 7531 2269
rect 7565 2235 7573 2269
rect 5406 2228 6611 2235
rect 5406 2195 5628 2228
rect 6320 2195 6611 2228
rect 6663 2195 6711 2235
rect 6763 2195 6811 2235
rect 6863 2195 6911 2235
rect 6963 2195 7011 2235
rect 7063 2195 7111 2235
rect 7163 2195 7211 2235
rect 7263 2195 7311 2235
rect 7363 2195 7573 2235
rect 5406 2161 5414 2195
rect 5448 2161 5486 2195
rect 5520 2161 5558 2195
rect 5592 2161 5628 2195
rect 6320 2161 6350 2195
rect 6384 2161 6595 2195
rect 6663 2190 6667 2195
rect 6629 2161 6667 2190
rect 6701 2190 6711 2195
rect 6701 2161 6739 2190
rect 6773 2161 6811 2195
rect 6863 2190 6883 2195
rect 6989 2190 7011 2195
rect 7063 2190 7099 2195
rect 7163 2190 7171 2195
rect 6845 2161 6883 2190
rect 6917 2161 6955 2190
rect 6989 2161 7027 2190
rect 7061 2161 7099 2190
rect 7133 2161 7171 2190
rect 7205 2190 7211 2195
rect 7277 2190 7311 2195
rect 7363 2190 7387 2195
rect 7205 2161 7243 2190
rect 7277 2161 7315 2190
rect 7349 2161 7387 2190
rect 7421 2161 7459 2195
rect 7493 2161 7531 2195
rect 7565 2161 7573 2195
rect 5406 2121 5628 2161
rect 6320 2121 7573 2161
rect 5406 2087 5414 2121
rect 5448 2087 5486 2121
rect 5520 2087 5558 2121
rect 5592 2087 5628 2121
rect 6320 2087 6350 2121
rect 6384 2087 6595 2121
rect 6629 2108 6667 2121
rect 6663 2087 6667 2108
rect 6701 2108 6739 2121
rect 6701 2087 6711 2108
rect 6773 2087 6811 2121
rect 6845 2108 6883 2121
rect 6917 2108 6955 2121
rect 6989 2108 7027 2121
rect 7061 2108 7099 2121
rect 7133 2108 7171 2121
rect 6863 2087 6883 2108
rect 6989 2087 7011 2108
rect 7063 2087 7099 2108
rect 7163 2087 7171 2108
rect 7205 2108 7243 2121
rect 7277 2108 7315 2121
rect 7349 2108 7387 2121
rect 7205 2087 7211 2108
rect 7277 2087 7311 2108
rect 7363 2087 7387 2108
rect 7421 2087 7459 2121
rect 7493 2087 7531 2121
rect 7565 2087 7573 2121
rect 5406 2047 5628 2087
rect 6320 2056 6611 2087
rect 6663 2056 6711 2087
rect 6763 2056 6811 2087
rect 6863 2056 6911 2087
rect 6963 2056 7011 2087
rect 7063 2056 7111 2087
rect 7163 2056 7211 2087
rect 7263 2056 7311 2087
rect 7363 2056 7573 2087
rect 6320 2047 7573 2056
rect 5406 2013 5414 2047
rect 5448 2013 5486 2047
rect 5520 2013 5558 2047
rect 5592 2013 5628 2047
rect 6320 2013 6350 2047
rect 6384 2013 6595 2047
rect 6629 2013 6667 2047
rect 6701 2013 6739 2047
rect 6773 2013 6811 2047
rect 6845 2013 6883 2047
rect 6917 2013 6955 2047
rect 6989 2013 7027 2047
rect 7061 2013 7099 2047
rect 7133 2013 7171 2047
rect 7205 2013 7243 2047
rect 7277 2013 7315 2047
rect 7349 2013 7387 2047
rect 7421 2013 7459 2047
rect 7493 2013 7531 2047
rect 7565 2013 7573 2047
rect 5406 1973 5628 2013
rect 6320 1973 7573 2013
rect 5406 1939 5414 1973
rect 5448 1939 5486 1973
rect 5520 1939 5558 1973
rect 5592 1939 5628 1973
rect 6320 1939 6350 1973
rect 6384 1939 6595 1973
rect 6663 1939 6667 1973
rect 6701 1939 6711 1973
rect 6773 1939 6811 1973
rect 6863 1939 6883 1973
rect 6989 1939 7011 1973
rect 7063 1939 7099 1973
rect 7163 1939 7171 1973
rect 7205 1939 7211 1973
rect 7277 1939 7311 1973
rect 7363 1939 7387 1973
rect 7421 1939 7459 1973
rect 7493 1939 7531 1973
rect 7565 1939 7573 1973
rect 5406 1899 5628 1939
rect 6320 1921 6611 1939
rect 6663 1921 6711 1939
rect 6763 1921 6811 1939
rect 6863 1921 6911 1939
rect 6963 1921 7011 1939
rect 7063 1921 7111 1939
rect 7163 1921 7211 1939
rect 7263 1921 7311 1939
rect 7363 1921 7573 1939
rect 6320 1899 7573 1921
rect 5406 1865 5414 1899
rect 5448 1865 5486 1899
rect 5520 1865 5558 1899
rect 5592 1865 5628 1899
rect 6320 1865 6350 1899
rect 6384 1865 6595 1899
rect 6629 1865 6667 1899
rect 6701 1865 6739 1899
rect 6773 1865 6811 1899
rect 6845 1865 6883 1899
rect 6917 1865 6955 1899
rect 6989 1865 7027 1899
rect 7061 1865 7099 1899
rect 7133 1865 7171 1899
rect 7205 1865 7243 1899
rect 7277 1865 7315 1899
rect 7349 1865 7387 1899
rect 7421 1865 7459 1899
rect 7493 1865 7531 1899
rect 7565 1865 7573 1899
rect 5406 1825 5628 1865
rect 6320 1838 7573 1865
rect 6320 1825 6611 1838
rect 6663 1825 6711 1838
rect 6763 1825 6811 1838
rect 6863 1825 6911 1838
rect 6963 1825 7011 1838
rect 7063 1825 7111 1838
rect 7163 1825 7211 1838
rect 7263 1825 7311 1838
rect 7363 1825 7573 1838
rect 5406 1791 5414 1825
rect 5448 1791 5486 1825
rect 5520 1791 5558 1825
rect 5592 1791 5628 1825
rect 6320 1791 6350 1825
rect 6384 1791 6595 1825
rect 6663 1791 6667 1825
rect 6701 1791 6711 1825
rect 6773 1791 6811 1825
rect 6863 1791 6883 1825
rect 6989 1791 7011 1825
rect 7063 1791 7099 1825
rect 7163 1791 7171 1825
rect 7205 1791 7211 1825
rect 7277 1791 7311 1825
rect 7363 1791 7387 1825
rect 7421 1791 7459 1825
rect 7493 1791 7531 1825
rect 7565 1791 7573 1825
rect 5406 1751 5628 1791
rect 6320 1786 6611 1791
rect 6663 1786 6711 1791
rect 6763 1786 6811 1791
rect 6863 1786 6911 1791
rect 6963 1786 7011 1791
rect 7063 1786 7111 1791
rect 7163 1786 7211 1791
rect 7263 1786 7311 1791
rect 7363 1786 7573 1791
rect 6320 1751 7573 1786
rect 5406 1717 5414 1751
rect 5448 1717 5486 1751
rect 5520 1717 5558 1751
rect 5592 1717 5628 1751
rect 6320 1717 6350 1751
rect 6384 1717 6595 1751
rect 6629 1717 6667 1751
rect 6701 1717 6739 1751
rect 6773 1717 6811 1751
rect 6845 1717 6883 1751
rect 6917 1717 6955 1751
rect 6989 1717 7027 1751
rect 7061 1717 7099 1751
rect 7133 1717 7171 1751
rect 7205 1717 7243 1751
rect 7277 1717 7315 1751
rect 7349 1717 7387 1751
rect 7421 1717 7459 1751
rect 7493 1717 7531 1751
rect 7565 1717 7573 1751
rect 5406 1676 5628 1717
rect 6320 1703 7573 1717
rect 6320 1676 6611 1703
rect 6663 1676 6711 1703
rect 6763 1676 6811 1703
rect 6863 1676 6911 1703
rect 6963 1676 7011 1703
rect 7063 1676 7111 1703
rect 7163 1676 7211 1703
rect 7263 1676 7311 1703
rect 7363 1676 7573 1703
rect 5406 1642 5414 1676
rect 5448 1642 5486 1676
rect 5520 1642 5558 1676
rect 5592 1642 5628 1676
rect 6320 1642 6350 1676
rect 6384 1642 6595 1676
rect 6663 1651 6667 1676
rect 6629 1642 6667 1651
rect 6701 1651 6711 1676
rect 6701 1642 6739 1651
rect 6773 1642 6811 1676
rect 6863 1651 6883 1676
rect 6989 1651 7011 1676
rect 7063 1651 7099 1676
rect 7163 1651 7171 1676
rect 6845 1642 6883 1651
rect 6917 1642 6955 1651
rect 6989 1642 7027 1651
rect 7061 1642 7099 1651
rect 7133 1642 7171 1651
rect 7205 1651 7211 1676
rect 7277 1651 7311 1676
rect 7363 1651 7387 1676
rect 7205 1642 7243 1651
rect 7277 1642 7315 1651
rect 7349 1642 7387 1651
rect 7421 1642 7459 1676
rect 7493 1642 7531 1676
rect 7565 1642 7573 1676
rect 5406 1601 5628 1642
rect 6320 1601 7573 1642
rect 5406 1567 5414 1601
rect 5448 1567 5486 1601
rect 5520 1567 5558 1601
rect 5592 1567 5628 1601
rect 6320 1567 6350 1601
rect 6384 1567 6595 1601
rect 6629 1568 6667 1601
rect 6663 1567 6667 1568
rect 6701 1568 6739 1601
rect 6701 1567 6711 1568
rect 6773 1567 6811 1601
rect 6845 1568 6883 1601
rect 6917 1568 6955 1601
rect 6989 1568 7027 1601
rect 7061 1568 7099 1601
rect 7133 1568 7171 1601
rect 6863 1567 6883 1568
rect 6989 1567 7011 1568
rect 7063 1567 7099 1568
rect 7163 1567 7171 1568
rect 7205 1568 7243 1601
rect 7277 1568 7315 1601
rect 7349 1568 7387 1601
rect 7205 1567 7211 1568
rect 7277 1567 7311 1568
rect 7363 1567 7387 1568
rect 7421 1567 7459 1601
rect 7493 1567 7531 1601
rect 7565 1567 7573 1601
rect 5406 1526 5628 1567
rect 6320 1526 6611 1567
rect 6663 1526 6711 1567
rect 6763 1526 6811 1567
rect 6863 1526 6911 1567
rect 6963 1526 7011 1567
rect 7063 1526 7111 1567
rect 7163 1526 7211 1567
rect 7263 1526 7311 1567
rect 7363 1526 7573 1567
rect 5406 1492 5414 1526
rect 5448 1492 5486 1526
rect 5520 1492 5558 1526
rect 5592 1492 5628 1526
rect 6320 1492 6350 1526
rect 6384 1492 6595 1526
rect 6663 1516 6667 1526
rect 6629 1492 6667 1516
rect 6701 1516 6711 1526
rect 6701 1492 6739 1516
rect 6773 1492 6811 1526
rect 6863 1516 6883 1526
rect 6989 1516 7011 1526
rect 7063 1516 7099 1526
rect 7163 1516 7171 1526
rect 6845 1492 6883 1516
rect 6917 1492 6955 1516
rect 6989 1492 7027 1516
rect 7061 1492 7099 1516
rect 7133 1492 7171 1516
rect 7205 1516 7211 1526
rect 7277 1516 7311 1526
rect 7363 1516 7387 1526
rect 7205 1492 7243 1516
rect 7277 1492 7315 1516
rect 7349 1492 7387 1516
rect 7421 1492 7459 1526
rect 7493 1492 7531 1526
rect 7565 1492 7573 1526
rect 5406 1451 5628 1492
rect 6320 1451 7573 1492
rect 5406 1417 5414 1451
rect 5448 1417 5486 1451
rect 5520 1417 5558 1451
rect 5592 1417 5628 1451
rect 6320 1417 6350 1451
rect 6384 1417 6595 1451
rect 6629 1433 6667 1451
rect 6663 1417 6667 1433
rect 6701 1433 6739 1451
rect 6701 1417 6711 1433
rect 6773 1417 6811 1451
rect 6845 1433 6883 1451
rect 6917 1433 6955 1451
rect 6989 1433 7027 1451
rect 7061 1433 7099 1451
rect 7133 1433 7171 1451
rect 6863 1417 6883 1433
rect 6989 1417 7011 1433
rect 7063 1417 7099 1433
rect 7163 1417 7171 1433
rect 7205 1433 7243 1451
rect 7277 1433 7315 1451
rect 7349 1433 7387 1451
rect 7205 1417 7211 1433
rect 7277 1417 7311 1433
rect 7363 1417 7387 1433
rect 7421 1417 7459 1451
rect 7493 1417 7531 1451
rect 7565 1417 7573 1451
rect 5406 1376 5628 1417
rect 6320 1381 6611 1417
rect 6663 1381 6711 1417
rect 6763 1381 6811 1417
rect 6863 1381 6911 1417
rect 6963 1381 7011 1417
rect 7063 1381 7111 1417
rect 7163 1381 7211 1417
rect 7263 1381 7311 1417
rect 7363 1381 7573 1417
rect 6320 1376 7573 1381
rect 5406 1342 5414 1376
rect 5448 1342 5486 1376
rect 5520 1342 5558 1376
rect 5592 1342 5628 1376
rect 6320 1342 6350 1376
rect 6384 1342 6595 1376
rect 6629 1342 6667 1376
rect 6701 1342 6739 1376
rect 6773 1342 6811 1376
rect 6845 1342 6883 1376
rect 6917 1342 6955 1376
rect 6989 1342 7027 1376
rect 7061 1342 7099 1376
rect 7133 1342 7171 1376
rect 7205 1342 7243 1376
rect 7277 1342 7315 1376
rect 7349 1342 7387 1376
rect 7421 1342 7459 1376
rect 7493 1342 7531 1376
rect 7565 1342 7573 1376
rect 5406 1301 5628 1342
rect 6320 1301 7573 1342
rect 5406 1267 5414 1301
rect 5448 1267 5486 1301
rect 5520 1267 5558 1301
rect 5592 1267 5628 1301
rect 6320 1267 6350 1301
rect 6384 1267 6595 1301
rect 6629 1298 6667 1301
rect 6663 1267 6667 1298
rect 6701 1298 6739 1301
rect 6701 1267 6711 1298
rect 6773 1267 6811 1301
rect 6845 1298 6883 1301
rect 6917 1298 6955 1301
rect 6989 1298 7027 1301
rect 7061 1298 7099 1301
rect 7133 1298 7171 1301
rect 6863 1267 6883 1298
rect 6989 1267 7011 1298
rect 7063 1267 7099 1298
rect 7163 1267 7171 1298
rect 7205 1298 7243 1301
rect 7277 1298 7315 1301
rect 7349 1298 7387 1301
rect 7205 1267 7211 1298
rect 7277 1267 7311 1298
rect 7363 1267 7387 1298
rect 7421 1267 7459 1301
rect 7493 1267 7531 1301
rect 7565 1267 7573 1301
rect 5406 1226 5628 1267
rect 6320 1246 6611 1267
rect 6663 1246 6711 1267
rect 6763 1246 6811 1267
rect 6863 1246 6911 1267
rect 6963 1246 7011 1267
rect 7063 1246 7111 1267
rect 7163 1246 7211 1267
rect 7263 1246 7311 1267
rect 7363 1246 7573 1267
rect 6320 1226 7573 1246
rect 5406 1192 5414 1226
rect 5448 1192 5486 1226
rect 5520 1192 5558 1226
rect 5592 1192 5628 1226
rect 6320 1192 6350 1226
rect 6384 1192 6595 1226
rect 6629 1192 6667 1226
rect 6701 1192 6739 1226
rect 6773 1192 6811 1226
rect 6845 1192 6883 1226
rect 6917 1192 6955 1226
rect 6989 1192 7027 1226
rect 7061 1192 7099 1226
rect 7133 1192 7171 1226
rect 7205 1192 7243 1226
rect 7277 1192 7315 1226
rect 7349 1192 7387 1226
rect 7421 1192 7459 1226
rect 7493 1192 7531 1226
rect 7565 1192 7573 1226
rect 5406 1152 5628 1192
rect 6320 1163 7573 1192
rect 6320 1152 6611 1163
rect 5406 1151 6611 1152
rect 6663 1151 6711 1163
rect 6763 1151 6811 1163
rect 6863 1151 6911 1163
rect 6963 1151 7011 1163
rect 7063 1151 7111 1163
rect 7163 1151 7211 1163
rect 7263 1151 7311 1163
rect 7363 1151 7573 1163
rect 5406 1117 5414 1151
rect 5448 1117 5486 1151
rect 5520 1117 5558 1151
rect 5592 1139 5630 1151
rect 5664 1139 5702 1151
rect 5736 1139 5774 1151
rect 5808 1139 5846 1151
rect 5880 1139 5918 1151
rect 5952 1139 5990 1151
rect 6024 1139 6062 1151
rect 6096 1139 6134 1151
rect 6168 1139 6206 1151
rect 6240 1139 6278 1151
rect 6312 1139 6350 1151
rect 5592 1117 5628 1139
rect 5406 1087 5628 1117
rect 5680 1087 5692 1139
rect 5744 1087 5756 1139
rect 5808 1087 5820 1139
rect 5880 1117 5884 1139
rect 6128 1117 6134 1139
rect 5872 1087 5884 1117
rect 5936 1087 5948 1117
rect 6000 1087 6012 1117
rect 6064 1087 6076 1117
rect 6128 1087 6140 1117
rect 6192 1087 6204 1139
rect 6256 1087 6268 1139
rect 6320 1117 6350 1139
rect 6384 1117 6595 1151
rect 6663 1117 6667 1151
rect 6701 1117 6711 1151
rect 6773 1117 6811 1151
rect 6863 1117 6883 1151
rect 6989 1117 7011 1151
rect 7063 1117 7099 1151
rect 7163 1117 7171 1151
rect 7205 1117 7211 1151
rect 7277 1117 7311 1151
rect 7363 1117 7387 1151
rect 7421 1117 7459 1151
rect 7493 1117 7531 1151
rect 7565 1117 7573 1151
rect 6320 1111 6611 1117
rect 6663 1111 6711 1117
rect 6763 1111 6811 1117
rect 6863 1111 6911 1117
rect 6963 1111 7011 1117
rect 7063 1111 7111 1117
rect 7163 1111 7211 1117
rect 7263 1111 7311 1117
rect 7363 1111 7573 1117
rect 6320 1087 7573 1111
rect 5406 1076 7573 1087
rect 5406 1042 5414 1076
rect 5448 1042 5486 1076
rect 5520 1042 5558 1076
rect 5592 1074 5630 1076
rect 5664 1074 5702 1076
rect 5736 1074 5774 1076
rect 5808 1074 5846 1076
rect 5880 1074 5918 1076
rect 5952 1074 5990 1076
rect 6024 1074 6062 1076
rect 6096 1074 6134 1076
rect 6168 1074 6206 1076
rect 6240 1074 6278 1076
rect 6312 1074 6350 1076
rect 5592 1042 5628 1074
rect 5406 1022 5628 1042
rect 5680 1022 5692 1074
rect 5744 1022 5756 1074
rect 5808 1022 5820 1074
rect 5880 1042 5884 1074
rect 6128 1042 6134 1074
rect 5872 1022 5884 1042
rect 5936 1022 5948 1042
rect 6000 1022 6012 1042
rect 6064 1022 6076 1042
rect 6128 1022 6140 1042
rect 6192 1022 6204 1074
rect 6256 1022 6268 1074
rect 6320 1042 6350 1074
rect 6384 1042 6595 1076
rect 6629 1042 6667 1076
rect 6701 1042 6739 1076
rect 6773 1042 6811 1076
rect 6845 1042 6883 1076
rect 6917 1042 6955 1076
rect 6989 1042 7027 1076
rect 7061 1042 7099 1076
rect 7133 1042 7171 1076
rect 7205 1042 7243 1076
rect 7277 1042 7315 1076
rect 7349 1042 7387 1076
rect 7421 1042 7459 1076
rect 7493 1042 7531 1076
rect 7565 1042 7573 1076
rect 6320 1028 7573 1042
rect 6320 1022 6611 1028
rect 5406 1009 6611 1022
rect 5406 1001 5628 1009
rect 5406 967 5414 1001
rect 5448 967 5486 1001
rect 5520 967 5558 1001
rect 5592 967 5628 1001
rect 5406 957 5628 967
rect 5680 957 5692 1009
rect 5744 957 5756 1009
rect 5808 957 5820 1009
rect 5872 1001 5884 1009
rect 5936 1001 5948 1009
rect 6000 1001 6012 1009
rect 6064 1001 6076 1009
rect 6128 1001 6140 1009
rect 5880 967 5884 1001
rect 6128 967 6134 1001
rect 5872 957 5884 967
rect 5936 957 5948 967
rect 6000 957 6012 967
rect 6064 957 6076 967
rect 6128 957 6140 967
rect 6192 957 6204 1009
rect 6256 957 6268 1009
rect 6320 1001 6611 1009
rect 6663 1001 6711 1028
rect 6763 1001 6811 1028
rect 6863 1001 6911 1028
rect 6963 1001 7011 1028
rect 7063 1001 7111 1028
rect 7163 1001 7211 1028
rect 7263 1001 7311 1028
rect 7363 1001 7573 1028
rect 6320 967 6350 1001
rect 6384 967 6595 1001
rect 6663 976 6667 1001
rect 6629 967 6667 976
rect 6701 976 6711 1001
rect 6701 967 6739 976
rect 6773 967 6811 1001
rect 6863 976 6883 1001
rect 6989 976 7011 1001
rect 7063 976 7099 1001
rect 7163 976 7171 1001
rect 6845 967 6883 976
rect 6917 967 6955 976
rect 6989 967 7027 976
rect 7061 967 7099 976
rect 7133 967 7171 976
rect 7205 976 7211 1001
rect 7277 976 7311 1001
rect 7363 976 7387 1001
rect 7205 967 7243 976
rect 7277 967 7315 976
rect 7349 967 7387 976
rect 7421 967 7459 1001
rect 7493 967 7531 1001
rect 7565 967 7573 1001
rect 6320 957 7573 967
rect 5406 944 7573 957
rect 5406 926 5628 944
rect 5406 892 5414 926
rect 5448 892 5486 926
rect 5520 892 5558 926
rect 5592 892 5628 926
rect 5680 892 5692 944
rect 5744 892 5756 944
rect 5808 892 5820 944
rect 5872 926 5884 944
rect 5936 926 5948 944
rect 6000 926 6012 944
rect 6064 926 6076 944
rect 6128 926 6140 944
rect 5880 892 5884 926
rect 6128 892 6134 926
rect 6192 892 6204 944
rect 6256 892 6268 944
rect 6320 926 7573 944
rect 6320 892 6350 926
rect 6384 892 6595 926
rect 6629 893 6667 926
rect 6663 892 6667 893
rect 6701 893 6739 926
rect 6701 892 6711 893
rect 6773 892 6811 926
rect 6845 893 6883 926
rect 6917 893 6955 926
rect 6989 893 7027 926
rect 7061 893 7099 926
rect 7133 893 7171 926
rect 6863 892 6883 893
rect 6989 892 7011 893
rect 7063 892 7099 893
rect 7163 892 7171 893
rect 7205 893 7243 926
rect 7277 893 7315 926
rect 7349 893 7387 926
rect 7205 892 7211 893
rect 7277 892 7311 893
rect 7363 892 7387 893
rect 7421 892 7459 926
rect 7493 892 7531 926
rect 7565 892 7573 926
rect 5406 879 6611 892
rect 2136 851 2263 858
tri 2263 851 2270 858 nw
rect 5406 851 5628 879
tri 2089 817 2123 851 se
rect 2123 817 2229 851
tri 2229 817 2263 851 nw
rect 5406 817 5414 851
rect 5448 817 5486 851
rect 5520 817 5558 851
rect 5592 827 5628 851
rect 5680 827 5692 879
rect 5744 827 5756 879
rect 5808 827 5820 879
rect 5872 851 5884 879
rect 5936 851 5948 879
rect 6000 851 6012 879
rect 6064 851 6076 879
rect 6128 851 6140 879
rect 5880 827 5884 851
rect 6128 827 6134 851
rect 6192 827 6204 879
rect 6256 827 6268 879
rect 6320 851 6611 879
rect 6663 851 6711 892
rect 6763 851 6811 892
rect 6863 851 6911 892
rect 6963 851 7011 892
rect 7063 851 7111 892
rect 7163 851 7211 892
rect 7263 851 7311 892
rect 7363 851 7573 892
rect 6320 827 6350 851
rect 5592 817 5630 827
rect 5664 817 5702 827
rect 5736 817 5774 827
rect 5808 817 5846 827
rect 5880 817 5918 827
rect 5952 817 5990 827
rect 6024 817 6062 827
rect 6096 817 6134 827
rect 6168 817 6206 827
rect 6240 817 6278 827
rect 6312 817 6350 827
rect 6384 817 6595 851
rect 6663 841 6667 851
rect 6629 817 6667 841
rect 6701 841 6711 851
rect 6701 817 6739 841
rect 6773 817 6811 851
rect 6863 841 6883 851
rect 6989 841 7011 851
rect 7063 841 7099 851
rect 7163 841 7171 851
rect 6845 817 6883 841
rect 6917 817 6955 841
rect 6989 817 7027 841
rect 7061 817 7099 841
rect 7133 817 7171 841
rect 7205 841 7211 851
rect 7277 841 7311 851
rect 7363 841 7387 851
rect 7205 817 7243 841
rect 7277 817 7315 841
rect 7349 817 7387 841
rect 7421 817 7459 851
rect 7493 817 7531 851
rect 7565 817 7573 851
tri 1811 476 1852 517 se
rect 1852 508 1959 517
rect 1852 476 1927 508
tri 1927 476 1959 508 nw
tri 2081 809 2089 817 se
rect 2089 809 2188 817
rect 2081 776 2188 809
tri 2188 776 2229 817 nw
rect 5406 814 7573 817
rect 5406 776 5628 814
tri 1777 442 1811 476 se
rect 1811 442 1893 476
tri 1893 442 1927 476 nw
tri 1762 427 1777 442 se
rect 1777 427 1878 442
tri 1878 427 1893 442 nw
tri 1682 347 1762 427 se
rect 1762 347 1798 427
tri 1798 347 1878 427 nw
rect 1346 341 1681 347
rect 75 296 215 308
rect 75 262 81 296
rect 115 262 175 296
rect 209 262 215 296
rect 75 213 215 262
rect 1346 307 1358 341
rect 1392 307 1451 341
rect 1485 307 1543 341
rect 1577 307 1635 341
rect 1669 307 1681 341
rect 1346 269 1681 307
rect 1346 235 1358 269
rect 1392 235 1451 269
rect 1485 235 1543 269
rect 1577 235 1635 269
rect 1669 235 1681 269
rect 1346 229 1681 235
tri 1681 230 1798 347 nw
rect 75 179 81 213
rect 115 179 175 213
rect 209 179 215 213
rect 75 158 215 179
tri 215 158 278 221 sw
tri 2031 158 2081 208 se
rect 2081 158 2180 776
tri 2180 768 2188 776 nw
rect 5406 742 5414 776
rect 5448 742 5486 776
rect 5520 742 5558 776
rect 5592 762 5628 776
rect 5680 762 5692 814
rect 5744 762 5756 814
rect 5808 762 5820 814
rect 5872 776 5884 814
rect 5936 776 5948 814
rect 6000 776 6012 814
rect 6064 776 6076 814
rect 6128 776 6140 814
rect 5880 762 5884 776
rect 6128 762 6134 776
rect 6192 762 6204 814
rect 6256 762 6268 814
rect 6320 776 7573 814
rect 6320 762 6350 776
rect 5592 749 5630 762
rect 5664 749 5702 762
rect 5736 749 5774 762
rect 5808 749 5846 762
rect 5880 749 5918 762
rect 5952 749 5990 762
rect 6024 749 6062 762
rect 6096 749 6134 762
rect 6168 749 6206 762
rect 6240 749 6278 762
rect 6312 749 6350 762
rect 5592 742 5628 749
rect 5406 701 5628 742
rect 5406 667 5414 701
rect 5448 667 5486 701
rect 5520 667 5558 701
rect 5592 697 5628 701
rect 5680 697 5692 749
rect 5744 697 5756 749
rect 5808 697 5820 749
rect 5880 742 5884 749
rect 6128 742 6134 749
rect 5872 701 5884 742
rect 5936 701 5948 742
rect 6000 701 6012 742
rect 6064 701 6076 742
rect 6128 701 6140 742
rect 5880 697 5884 701
rect 6128 697 6134 701
rect 6192 697 6204 749
rect 6256 697 6268 749
rect 6320 742 6350 749
rect 6384 742 6595 776
rect 6629 758 6667 776
rect 6663 742 6667 758
rect 6701 758 6739 776
rect 6701 742 6711 758
rect 6773 742 6811 776
rect 6845 758 6883 776
rect 6917 758 6955 776
rect 6989 758 7027 776
rect 7061 758 7099 776
rect 7133 758 7171 776
rect 6863 742 6883 758
rect 6989 742 7011 758
rect 7063 742 7099 758
rect 7163 742 7171 758
rect 7205 758 7243 776
rect 7277 758 7315 776
rect 7349 758 7387 776
rect 7205 742 7211 758
rect 7277 742 7311 758
rect 7363 742 7387 758
rect 7421 742 7459 776
rect 7493 742 7531 776
rect 7565 742 7573 776
rect 6320 706 6611 742
rect 6663 706 6711 742
rect 6763 706 6811 742
rect 6863 706 6911 742
rect 6963 706 7011 742
rect 7063 706 7111 742
rect 7163 706 7211 742
rect 7263 706 7311 742
rect 7363 706 7573 742
rect 6320 701 7573 706
rect 6320 697 6350 701
rect 5592 684 5630 697
rect 5664 684 5702 697
rect 5736 684 5774 697
rect 5808 684 5846 697
rect 5880 684 5918 697
rect 5952 684 5990 697
rect 6024 684 6062 697
rect 6096 684 6134 697
rect 6168 684 6206 697
rect 6240 684 6278 697
rect 6312 684 6350 697
rect 5592 667 5628 684
rect 5406 632 5628 667
rect 5680 632 5692 684
rect 5744 632 5756 684
rect 5808 632 5820 684
rect 5880 667 5884 684
rect 6128 667 6134 684
rect 5872 632 5884 667
rect 5936 632 5948 667
rect 6000 632 6012 667
rect 6064 632 6076 667
rect 6128 632 6140 667
rect 6192 632 6204 684
rect 6256 632 6268 684
rect 6320 667 6350 684
rect 6384 667 6595 701
rect 6629 667 6667 701
rect 6701 667 6739 701
rect 6773 667 6811 701
rect 6845 667 6883 701
rect 6917 667 6955 701
rect 6989 667 7027 701
rect 7061 667 7099 701
rect 7133 667 7171 701
rect 7205 667 7243 701
rect 7277 667 7315 701
rect 7349 667 7387 701
rect 7421 667 7459 701
rect 7493 667 7531 701
rect 7565 667 7573 701
rect 6320 632 7573 667
rect 5406 626 7573 632
rect 5406 592 5414 626
rect 5448 592 5486 626
rect 5520 592 5558 626
rect 5592 619 5630 626
rect 5664 619 5702 626
rect 5736 619 5774 626
rect 5808 619 5846 626
rect 5880 619 5918 626
rect 5952 619 5990 626
rect 6024 619 6062 626
rect 6096 619 6134 626
rect 6168 619 6206 626
rect 6240 619 6278 626
rect 6312 619 6350 626
rect 5592 592 5628 619
rect 5406 567 5628 592
rect 5680 567 5692 619
rect 5744 567 5756 619
rect 5808 567 5820 619
rect 5880 592 5884 619
rect 6128 592 6134 619
rect 5872 567 5884 592
rect 5936 567 5948 592
rect 6000 567 6012 592
rect 6064 567 6076 592
rect 6128 567 6140 592
rect 6192 567 6204 619
rect 6256 567 6268 619
rect 6320 592 6350 619
rect 6384 592 6595 626
rect 6629 623 6667 626
rect 6663 592 6667 623
rect 6701 623 6739 626
rect 6701 592 6711 623
rect 6773 592 6811 626
rect 6845 623 6883 626
rect 6917 623 6955 626
rect 6989 623 7027 626
rect 7061 623 7099 626
rect 7133 623 7171 626
rect 6863 592 6883 623
rect 6989 592 7011 623
rect 7063 592 7099 623
rect 7163 592 7171 623
rect 7205 623 7243 626
rect 7277 623 7315 626
rect 7349 623 7387 626
rect 7205 592 7211 623
rect 7277 592 7311 623
rect 7363 592 7387 623
rect 7421 592 7459 626
rect 7493 592 7531 626
rect 7565 592 7573 626
rect 6320 571 6611 592
rect 6663 571 6711 592
rect 6763 571 6811 592
rect 6863 571 6911 592
rect 6963 571 7011 592
rect 7063 571 7111 592
rect 7163 571 7211 592
rect 7263 571 7311 592
rect 7363 571 7573 592
rect 6320 567 7573 571
rect 5406 554 7573 567
rect 5406 551 5628 554
rect 5406 517 5414 551
rect 5448 517 5486 551
rect 5520 517 5558 551
rect 5592 517 5628 551
rect 5406 502 5628 517
rect 5680 502 5692 554
rect 5744 502 5756 554
rect 5808 502 5820 554
rect 5872 551 5884 554
rect 5936 551 5948 554
rect 6000 551 6012 554
rect 6064 551 6076 554
rect 6128 551 6140 554
rect 5880 517 5884 551
rect 6128 517 6134 551
rect 5872 502 5884 517
rect 5936 502 5948 517
rect 6000 502 6012 517
rect 6064 502 6076 517
rect 6128 502 6140 517
rect 6192 502 6204 554
rect 6256 502 6268 554
rect 6320 551 7573 554
rect 6320 517 6350 551
rect 6384 517 6595 551
rect 6629 517 6667 551
rect 6701 517 6739 551
rect 6773 517 6811 551
rect 6845 517 6883 551
rect 6917 517 6955 551
rect 6989 517 7027 551
rect 7061 517 7099 551
rect 7133 517 7171 551
rect 7205 517 7243 551
rect 7277 517 7315 551
rect 7349 517 7387 551
rect 7421 517 7459 551
rect 7493 517 7531 551
rect 7565 517 7573 551
rect 6320 502 7573 517
rect 5406 489 7573 502
rect 5406 476 5628 489
rect 5406 442 5414 476
rect 5448 442 5486 476
rect 5520 442 5558 476
rect 5592 442 5628 476
rect 5406 437 5628 442
rect 5680 437 5692 489
rect 5744 437 5756 489
rect 5808 437 5820 489
rect 5872 476 5884 489
rect 5936 476 5948 489
rect 6000 476 6012 489
rect 6064 476 6076 489
rect 6128 476 6140 489
rect 5880 442 5884 476
rect 6128 442 6134 476
rect 5872 437 5884 442
rect 5936 437 5948 442
rect 6000 437 6012 442
rect 6064 437 6076 442
rect 6128 437 6140 442
rect 6192 437 6204 489
rect 6256 437 6268 489
rect 6320 488 7573 489
rect 6320 476 6611 488
rect 6663 476 6711 488
rect 6763 476 6811 488
rect 6863 476 6911 488
rect 6963 476 7011 488
rect 7063 476 7111 488
rect 7163 476 7211 488
rect 7263 476 7311 488
rect 7363 476 7573 488
rect 6320 442 6350 476
rect 6384 442 6595 476
rect 6663 442 6667 476
rect 6701 442 6711 476
rect 6773 442 6811 476
rect 6863 442 6883 476
rect 6989 442 7011 476
rect 7063 442 7099 476
rect 7163 442 7171 476
rect 7205 442 7211 476
rect 7277 442 7311 476
rect 7363 442 7387 476
rect 7421 442 7459 476
rect 7493 442 7531 476
rect 7565 442 7573 476
rect 6320 437 6611 442
rect 5406 436 6611 437
rect 6663 436 6711 442
rect 6763 436 6811 442
rect 6863 436 6911 442
rect 6963 436 7011 442
rect 7063 436 7111 442
rect 7163 436 7211 442
rect 7263 436 7311 442
rect 7363 436 7573 442
rect 5406 430 7573 436
rect 75 143 2180 158
rect 75 130 2099 143
rect 75 96 81 130
rect 115 96 175 130
rect 209 96 2099 130
rect 75 62 2099 96
tri 2099 62 2180 143 nw
rect 7727 0 7877 3341
<< via1 >>
rect 1938 26968 1944 27020
rect 1944 26968 1990 27020
rect 2004 26968 2050 27020
rect 2050 26968 2056 27020
rect 1938 26904 1944 26956
rect 1944 26904 1990 26956
rect 2004 26904 2050 26956
rect 2050 26904 2056 26956
rect 2270 38704 2322 38724
rect 2270 38672 2276 38704
rect 2276 38672 2310 38704
rect 2310 38672 2322 38704
rect 2392 38715 2444 38724
rect 2392 38681 2410 38715
rect 2410 38681 2444 38715
rect 2392 38672 2444 38681
rect 2270 38631 2322 38655
rect 2270 38603 2276 38631
rect 2276 38603 2310 38631
rect 2310 38603 2322 38631
rect 2392 38642 2444 38655
rect 2392 38608 2410 38642
rect 2410 38608 2444 38642
rect 2392 38603 2444 38608
rect 2270 38558 2322 38586
rect 2270 38534 2276 38558
rect 2276 38534 2310 38558
rect 2310 38534 2322 38558
rect 2392 38569 2444 38586
rect 2392 38535 2410 38569
rect 2410 38535 2444 38569
rect 2392 38534 2444 38535
rect 2270 38485 2322 38517
rect 2270 38465 2276 38485
rect 2276 38465 2310 38485
rect 2310 38465 2322 38485
rect 2392 38496 2444 38517
rect 2392 38465 2410 38496
rect 2410 38465 2444 38496
rect 2270 38412 2322 38448
rect 2270 38396 2276 38412
rect 2276 38396 2310 38412
rect 2310 38396 2322 38412
rect 2392 38423 2444 38448
rect 2392 38396 2410 38423
rect 2410 38396 2444 38423
rect 2270 38339 2322 38378
rect 2270 38326 2276 38339
rect 2276 38326 2310 38339
rect 2310 38326 2322 38339
rect 2392 38350 2444 38378
rect 2392 38326 2410 38350
rect 2410 38326 2444 38350
rect 2270 38305 2276 38308
rect 2276 38305 2310 38308
rect 2310 38305 2322 38308
rect 2270 38266 2322 38305
rect 2270 38256 2276 38266
rect 2276 38256 2310 38266
rect 2310 38256 2322 38266
rect 2392 38277 2444 38308
rect 2392 38256 2410 38277
rect 2410 38256 2444 38277
rect 2270 38232 2276 38238
rect 2276 38232 2310 38238
rect 2310 38232 2322 38238
rect 2270 38193 2322 38232
rect 2270 38186 2276 38193
rect 2276 38186 2310 38193
rect 2310 38186 2322 38193
rect 2392 38204 2444 38238
rect 2392 38186 2410 38204
rect 2410 38186 2444 38204
rect 2270 38159 2276 38168
rect 2276 38159 2310 38168
rect 2310 38159 2322 38168
rect 2270 38120 2322 38159
rect 2270 38116 2276 38120
rect 2276 38116 2310 38120
rect 2310 38116 2322 38120
rect 2392 38131 2444 38168
rect 2392 38116 2410 38131
rect 2410 38116 2444 38131
rect 2270 36699 2276 36724
rect 2276 36699 2310 36724
rect 2310 36699 2322 36724
rect 2270 36672 2322 36699
rect 2392 36710 2410 36724
rect 2410 36710 2444 36724
rect 2392 36672 2444 36710
rect 2270 36626 2276 36655
rect 2276 36626 2310 36655
rect 2310 36626 2322 36655
rect 2270 36603 2322 36626
rect 2392 36637 2410 36655
rect 2410 36637 2444 36655
rect 2392 36603 2444 36637
rect 2270 36554 2276 36586
rect 2276 36554 2310 36586
rect 2310 36554 2322 36586
rect 2270 36534 2322 36554
rect 2392 36564 2410 36586
rect 2410 36564 2444 36586
rect 2392 36534 2444 36564
rect 2270 36516 2322 36517
rect 2270 36482 2276 36516
rect 2276 36482 2310 36516
rect 2310 36482 2322 36516
rect 2270 36465 2322 36482
rect 2392 36491 2410 36517
rect 2410 36491 2444 36517
rect 2392 36465 2444 36491
rect 2270 36444 2322 36448
rect 2270 36410 2276 36444
rect 2276 36410 2310 36444
rect 2310 36410 2322 36444
rect 2270 36396 2322 36410
rect 2392 36418 2410 36448
rect 2410 36418 2444 36448
rect 2392 36396 2444 36418
rect 2270 36372 2322 36378
rect 2270 36338 2276 36372
rect 2276 36338 2310 36372
rect 2310 36338 2322 36372
rect 2270 36326 2322 36338
rect 2392 36345 2410 36378
rect 2410 36345 2444 36378
rect 2392 36326 2444 36345
rect 2270 36300 2322 36308
rect 2270 36266 2276 36300
rect 2276 36266 2310 36300
rect 2310 36266 2322 36300
rect 2270 36256 2322 36266
rect 2392 36306 2444 36308
rect 2392 36272 2410 36306
rect 2410 36272 2444 36306
rect 2392 36256 2444 36272
rect 2270 36228 2322 36238
rect 2270 36194 2276 36228
rect 2276 36194 2310 36228
rect 2310 36194 2322 36228
rect 2270 36186 2322 36194
rect 2392 36233 2444 36238
rect 2392 36199 2410 36233
rect 2410 36199 2444 36233
rect 2392 36186 2444 36199
rect 2270 36156 2322 36168
rect 2270 36122 2276 36156
rect 2276 36122 2310 36156
rect 2310 36122 2322 36156
rect 2270 36116 2322 36122
rect 2392 36160 2444 36168
rect 2392 36126 2410 36160
rect 2410 36126 2444 36160
rect 2392 36116 2444 36126
rect 2270 34716 2322 34724
rect 2270 34682 2276 34716
rect 2276 34682 2310 34716
rect 2310 34682 2322 34716
rect 2270 34672 2322 34682
rect 2392 34716 2444 34724
rect 2392 34682 2410 34716
rect 2410 34682 2444 34716
rect 2392 34672 2444 34682
rect 2270 34644 2322 34655
rect 2270 34610 2276 34644
rect 2276 34610 2310 34644
rect 2310 34610 2322 34644
rect 2270 34603 2322 34610
rect 2392 34644 2444 34655
rect 2392 34610 2410 34644
rect 2410 34610 2444 34644
rect 2392 34603 2444 34610
rect 2270 34572 2322 34586
rect 2270 34538 2276 34572
rect 2276 34538 2310 34572
rect 2310 34538 2322 34572
rect 2270 34534 2322 34538
rect 2392 34572 2444 34586
rect 2392 34538 2410 34572
rect 2410 34538 2444 34572
rect 2392 34534 2444 34538
rect 2270 34500 2322 34517
rect 2270 34466 2276 34500
rect 2276 34466 2310 34500
rect 2310 34466 2322 34500
rect 2270 34465 2322 34466
rect 2392 34500 2444 34517
rect 2392 34466 2410 34500
rect 2410 34466 2444 34500
rect 2392 34465 2444 34466
rect 2270 34428 2322 34448
rect 2270 34396 2276 34428
rect 2276 34396 2310 34428
rect 2310 34396 2322 34428
rect 2392 34428 2444 34448
rect 2392 34396 2410 34428
rect 2410 34396 2444 34428
rect 2270 34356 2322 34378
rect 2270 34326 2276 34356
rect 2276 34326 2310 34356
rect 2310 34326 2322 34356
rect 2392 34356 2444 34378
rect 2392 34326 2410 34356
rect 2410 34326 2444 34356
rect 2270 34284 2322 34308
rect 2270 34256 2276 34284
rect 2276 34256 2310 34284
rect 2310 34256 2322 34284
rect 2392 34284 2444 34308
rect 2392 34256 2410 34284
rect 2410 34256 2444 34284
rect 2270 34212 2322 34238
rect 2270 34186 2276 34212
rect 2276 34186 2310 34212
rect 2310 34186 2322 34212
rect 2392 34212 2444 34238
rect 2392 34186 2410 34212
rect 2410 34186 2444 34212
rect 2270 34140 2322 34168
rect 2270 34116 2276 34140
rect 2276 34116 2310 34140
rect 2310 34116 2322 34140
rect 2392 34140 2444 34168
rect 2392 34116 2410 34140
rect 2410 34116 2444 34140
rect 2270 32700 2322 32724
rect 2270 32672 2276 32700
rect 2276 32672 2310 32700
rect 2310 32672 2322 32700
rect 2392 32700 2444 32724
rect 2392 32672 2410 32700
rect 2410 32672 2444 32700
rect 2270 32628 2322 32655
rect 2270 32603 2276 32628
rect 2276 32603 2310 32628
rect 2310 32603 2322 32628
rect 2392 32628 2444 32655
rect 2392 32603 2410 32628
rect 2410 32603 2444 32628
rect 2270 32556 2322 32586
rect 2270 32534 2276 32556
rect 2276 32534 2310 32556
rect 2310 32534 2322 32556
rect 2392 32556 2444 32586
rect 2392 32534 2410 32556
rect 2410 32534 2444 32556
rect 2270 32484 2322 32517
rect 2270 32465 2276 32484
rect 2276 32465 2310 32484
rect 2310 32465 2322 32484
rect 2392 32484 2444 32517
rect 2392 32465 2410 32484
rect 2410 32465 2444 32484
rect 2270 32412 2322 32448
rect 2270 32396 2276 32412
rect 2276 32396 2310 32412
rect 2310 32396 2322 32412
rect 2392 32412 2444 32448
rect 2392 32396 2410 32412
rect 2410 32396 2444 32412
rect 2270 32340 2322 32378
rect 2270 32326 2276 32340
rect 2276 32326 2310 32340
rect 2310 32326 2322 32340
rect 2392 32340 2444 32378
rect 2392 32326 2410 32340
rect 2410 32326 2444 32340
rect 2270 32306 2276 32308
rect 2276 32306 2310 32308
rect 2310 32306 2322 32308
rect 2270 32268 2322 32306
rect 2270 32256 2276 32268
rect 2276 32256 2310 32268
rect 2310 32256 2322 32268
rect 2392 32306 2410 32308
rect 2410 32306 2444 32308
rect 2392 32268 2444 32306
rect 2392 32256 2410 32268
rect 2410 32256 2444 32268
rect 2270 32234 2276 32238
rect 2276 32234 2310 32238
rect 2310 32234 2322 32238
rect 2270 32196 2322 32234
rect 2270 32186 2276 32196
rect 2276 32186 2310 32196
rect 2310 32186 2322 32196
rect 2392 32234 2410 32238
rect 2410 32234 2444 32238
rect 2392 32196 2444 32234
rect 2392 32186 2410 32196
rect 2410 32186 2444 32196
rect 2270 32162 2276 32168
rect 2276 32162 2310 32168
rect 2310 32162 2322 32168
rect 2270 32124 2322 32162
rect 2270 32116 2276 32124
rect 2276 32116 2310 32124
rect 2310 32116 2322 32124
rect 2392 32162 2410 32168
rect 2410 32162 2444 32168
rect 2392 32124 2444 32162
rect 2392 32116 2410 32124
rect 2410 32116 2444 32124
rect 2270 30722 2276 30724
rect 2276 30722 2310 30724
rect 2310 30722 2322 30724
rect 2270 30684 2322 30722
rect 2270 30672 2276 30684
rect 2276 30672 2310 30684
rect 2310 30672 2322 30684
rect 2392 30722 2410 30724
rect 2410 30722 2444 30724
rect 2392 30684 2444 30722
rect 2392 30672 2410 30684
rect 2410 30672 2444 30684
rect 2270 30650 2276 30655
rect 2276 30650 2310 30655
rect 2310 30650 2322 30655
rect 2270 30612 2322 30650
rect 2270 30603 2276 30612
rect 2276 30603 2310 30612
rect 2310 30603 2322 30612
rect 2392 30650 2410 30655
rect 2410 30650 2444 30655
rect 2392 30612 2444 30650
rect 2392 30603 2410 30612
rect 2410 30603 2444 30612
rect 2270 30578 2276 30586
rect 2276 30578 2310 30586
rect 2310 30578 2322 30586
rect 2270 30540 2322 30578
rect 2270 30534 2276 30540
rect 2276 30534 2310 30540
rect 2310 30534 2322 30540
rect 2392 30578 2410 30586
rect 2410 30578 2444 30586
rect 2392 30540 2444 30578
rect 2392 30534 2410 30540
rect 2410 30534 2444 30540
rect 2270 30506 2276 30517
rect 2276 30506 2310 30517
rect 2310 30506 2322 30517
rect 2270 30468 2322 30506
rect 2270 30465 2276 30468
rect 2276 30465 2310 30468
rect 2310 30465 2322 30468
rect 2392 30506 2410 30517
rect 2410 30506 2444 30517
rect 2392 30468 2444 30506
rect 2392 30465 2410 30468
rect 2410 30465 2444 30468
rect 2270 30434 2276 30448
rect 2276 30434 2310 30448
rect 2310 30434 2322 30448
rect 2270 30396 2322 30434
rect 2392 30434 2410 30448
rect 2410 30434 2444 30448
rect 2392 30396 2444 30434
rect 2270 30362 2276 30378
rect 2276 30362 2310 30378
rect 2310 30362 2322 30378
rect 2270 30326 2322 30362
rect 2392 30362 2410 30378
rect 2410 30362 2444 30378
rect 2392 30326 2444 30362
rect 2270 30290 2276 30308
rect 2276 30290 2310 30308
rect 2310 30290 2322 30308
rect 2270 30256 2322 30290
rect 2392 30290 2410 30308
rect 2410 30290 2444 30308
rect 2392 30256 2444 30290
rect 2270 30218 2276 30238
rect 2276 30218 2310 30238
rect 2310 30218 2322 30238
rect 2270 30186 2322 30218
rect 2392 30218 2410 30238
rect 2410 30218 2444 30238
rect 2392 30186 2444 30218
rect 2270 30146 2276 30168
rect 2276 30146 2310 30168
rect 2310 30146 2322 30168
rect 2270 30116 2322 30146
rect 2392 30146 2410 30168
rect 2410 30146 2444 30168
rect 2392 30116 2444 30146
rect 2824 38714 2876 38720
rect 2824 38680 2830 38714
rect 2830 38680 2864 38714
rect 2864 38680 2876 38714
rect 2824 38668 2876 38680
rect 2890 38714 2942 38720
rect 2890 38680 2902 38714
rect 2902 38680 2936 38714
rect 2936 38680 2942 38714
rect 2890 38668 2942 38680
rect 2824 38641 2876 38651
rect 2824 38607 2830 38641
rect 2830 38607 2864 38641
rect 2864 38607 2876 38641
rect 2824 38599 2876 38607
rect 2890 38641 2942 38651
rect 2890 38607 2902 38641
rect 2902 38607 2936 38641
rect 2936 38607 2942 38641
rect 2890 38599 2942 38607
rect 2824 38568 2876 38582
rect 2824 38534 2830 38568
rect 2830 38534 2864 38568
rect 2864 38534 2876 38568
rect 2824 38530 2876 38534
rect 2890 38568 2942 38582
rect 2890 38534 2902 38568
rect 2902 38534 2936 38568
rect 2936 38534 2942 38568
rect 2890 38530 2942 38534
rect 2824 38495 2876 38513
rect 2824 38461 2830 38495
rect 2830 38461 2864 38495
rect 2864 38461 2876 38495
rect 2890 38495 2942 38513
rect 2890 38461 2902 38495
rect 2902 38461 2936 38495
rect 2936 38461 2942 38495
rect 2824 38422 2876 38444
rect 2890 38422 2942 38444
rect 2824 38392 2830 38422
rect 2830 38392 2876 38422
rect 2890 38392 2936 38422
rect 2936 38392 2942 38422
rect 2824 38323 2830 38375
rect 2830 38323 2876 38375
rect 2890 38323 2936 38375
rect 2936 38323 2942 38375
rect 2824 38254 2830 38306
rect 2830 38254 2876 38306
rect 2890 38254 2936 38306
rect 2936 38254 2942 38306
rect 2824 38184 2830 38236
rect 2830 38184 2876 38236
rect 2890 38184 2936 38236
rect 2936 38184 2942 38236
rect 2824 38114 2830 38166
rect 2830 38114 2876 38166
rect 2890 38114 2936 38166
rect 2936 38114 2942 38166
rect 3101 37930 3107 37982
rect 3107 37930 3153 37982
rect 3167 37930 3213 37982
rect 3213 37930 3219 37982
rect 3101 37861 3107 37913
rect 3107 37861 3153 37913
rect 3167 37861 3213 37913
rect 3213 37861 3219 37913
rect 3101 37792 3107 37844
rect 3107 37792 3153 37844
rect 3167 37792 3213 37844
rect 3213 37792 3219 37844
rect 3101 37723 3107 37775
rect 3107 37723 3153 37775
rect 3167 37723 3213 37775
rect 3213 37723 3219 37775
rect 3101 37654 3107 37706
rect 3107 37654 3153 37706
rect 3167 37654 3213 37706
rect 3213 37654 3219 37706
rect 3101 37584 3107 37636
rect 3107 37584 3153 37636
rect 3167 37584 3213 37636
rect 3213 37584 3219 37636
rect 3101 37514 3107 37566
rect 3107 37514 3153 37566
rect 3167 37514 3213 37566
rect 3213 37514 3219 37566
rect 3101 37444 3107 37496
rect 3107 37444 3153 37496
rect 3167 37444 3213 37496
rect 3213 37444 3219 37496
rect 3101 37380 3107 37426
rect 3107 37380 3153 37426
rect 3167 37380 3213 37426
rect 3213 37380 3219 37426
rect 3101 37374 3153 37380
rect 3167 37374 3219 37380
rect 3378 38714 3430 38720
rect 3378 38680 3384 38714
rect 3384 38680 3418 38714
rect 3418 38680 3430 38714
rect 3378 38668 3430 38680
rect 3444 38714 3496 38720
rect 3444 38680 3456 38714
rect 3456 38680 3490 38714
rect 3490 38680 3496 38714
rect 3444 38668 3496 38680
rect 3378 38641 3430 38651
rect 3378 38607 3384 38641
rect 3384 38607 3418 38641
rect 3418 38607 3430 38641
rect 3378 38599 3430 38607
rect 3444 38641 3496 38651
rect 3444 38607 3456 38641
rect 3456 38607 3490 38641
rect 3490 38607 3496 38641
rect 3444 38599 3496 38607
rect 3378 38568 3430 38582
rect 3378 38534 3384 38568
rect 3384 38534 3418 38568
rect 3418 38534 3430 38568
rect 3378 38530 3430 38534
rect 3444 38568 3496 38582
rect 3444 38534 3456 38568
rect 3456 38534 3490 38568
rect 3490 38534 3496 38568
rect 3444 38530 3496 38534
rect 3378 38495 3430 38513
rect 3378 38461 3384 38495
rect 3384 38461 3418 38495
rect 3418 38461 3430 38495
rect 3444 38495 3496 38513
rect 3444 38461 3456 38495
rect 3456 38461 3490 38495
rect 3490 38461 3496 38495
rect 3378 38422 3430 38444
rect 3444 38422 3496 38444
rect 3378 38392 3384 38422
rect 3384 38392 3430 38422
rect 3444 38392 3490 38422
rect 3490 38392 3496 38422
rect 3378 38323 3384 38375
rect 3384 38323 3430 38375
rect 3444 38323 3490 38375
rect 3490 38323 3496 38375
rect 3378 38254 3384 38306
rect 3384 38254 3430 38306
rect 3444 38254 3490 38306
rect 3490 38254 3496 38306
rect 3378 38184 3384 38236
rect 3384 38184 3430 38236
rect 3444 38184 3490 38236
rect 3490 38184 3496 38236
rect 3378 38114 3384 38166
rect 3384 38114 3430 38166
rect 3444 38114 3490 38166
rect 3490 38114 3496 38166
rect 3655 37930 3661 37982
rect 3661 37930 3707 37982
rect 3721 37930 3767 37982
rect 3767 37930 3773 37982
rect 3655 37861 3661 37913
rect 3661 37861 3707 37913
rect 3721 37861 3767 37913
rect 3767 37861 3773 37913
rect 3655 37792 3661 37844
rect 3661 37792 3707 37844
rect 3721 37792 3767 37844
rect 3767 37792 3773 37844
rect 3655 37723 3661 37775
rect 3661 37723 3707 37775
rect 3721 37723 3767 37775
rect 3767 37723 3773 37775
rect 3655 37654 3661 37706
rect 3661 37654 3707 37706
rect 3721 37654 3767 37706
rect 3767 37654 3773 37706
rect 3655 37584 3661 37636
rect 3661 37584 3707 37636
rect 3721 37584 3767 37636
rect 3767 37584 3773 37636
rect 3655 37514 3661 37566
rect 3661 37514 3707 37566
rect 3721 37514 3767 37566
rect 3767 37514 3773 37566
rect 3655 37444 3661 37496
rect 3661 37444 3707 37496
rect 3721 37444 3767 37496
rect 3767 37444 3773 37496
rect 3655 37380 3661 37426
rect 3661 37380 3707 37426
rect 3721 37380 3767 37426
rect 3767 37380 3773 37426
rect 3655 37374 3707 37380
rect 3721 37374 3773 37380
rect 3932 38714 3984 38720
rect 3932 38680 3938 38714
rect 3938 38680 3972 38714
rect 3972 38680 3984 38714
rect 3932 38668 3984 38680
rect 3998 38714 4050 38720
rect 3998 38680 4010 38714
rect 4010 38680 4044 38714
rect 4044 38680 4050 38714
rect 3998 38668 4050 38680
rect 3932 38641 3984 38651
rect 3932 38607 3938 38641
rect 3938 38607 3972 38641
rect 3972 38607 3984 38641
rect 3932 38599 3984 38607
rect 3998 38641 4050 38651
rect 3998 38607 4010 38641
rect 4010 38607 4044 38641
rect 4044 38607 4050 38641
rect 3998 38599 4050 38607
rect 3932 38568 3984 38582
rect 3932 38534 3938 38568
rect 3938 38534 3972 38568
rect 3972 38534 3984 38568
rect 3932 38530 3984 38534
rect 3998 38568 4050 38582
rect 3998 38534 4010 38568
rect 4010 38534 4044 38568
rect 4044 38534 4050 38568
rect 3998 38530 4050 38534
rect 3932 38495 3984 38513
rect 3932 38461 3938 38495
rect 3938 38461 3972 38495
rect 3972 38461 3984 38495
rect 3998 38495 4050 38513
rect 3998 38461 4010 38495
rect 4010 38461 4044 38495
rect 4044 38461 4050 38495
rect 3932 38422 3984 38444
rect 3998 38422 4050 38444
rect 3932 38392 3938 38422
rect 3938 38392 3984 38422
rect 3998 38392 4044 38422
rect 4044 38392 4050 38422
rect 3932 38323 3938 38375
rect 3938 38323 3984 38375
rect 3998 38323 4044 38375
rect 4044 38323 4050 38375
rect 3932 38254 3938 38306
rect 3938 38254 3984 38306
rect 3998 38254 4044 38306
rect 4044 38254 4050 38306
rect 3932 38184 3938 38236
rect 3938 38184 3984 38236
rect 3998 38184 4044 38236
rect 4044 38184 4050 38236
rect 3932 38114 3938 38166
rect 3938 38114 3984 38166
rect 3998 38114 4044 38166
rect 4044 38114 4050 38166
rect 4209 37930 4215 37982
rect 4215 37930 4261 37982
rect 4275 37930 4321 37982
rect 4321 37930 4327 37982
rect 4209 37861 4215 37913
rect 4215 37861 4261 37913
rect 4275 37861 4321 37913
rect 4321 37861 4327 37913
rect 4209 37792 4215 37844
rect 4215 37792 4261 37844
rect 4275 37792 4321 37844
rect 4321 37792 4327 37844
rect 4209 37723 4215 37775
rect 4215 37723 4261 37775
rect 4275 37723 4321 37775
rect 4321 37723 4327 37775
rect 4209 37654 4215 37706
rect 4215 37654 4261 37706
rect 4275 37654 4321 37706
rect 4321 37654 4327 37706
rect 4209 37584 4215 37636
rect 4215 37584 4261 37636
rect 4275 37584 4321 37636
rect 4321 37584 4327 37636
rect 4209 37514 4215 37566
rect 4215 37514 4261 37566
rect 4275 37514 4321 37566
rect 4321 37514 4327 37566
rect 4209 37444 4215 37496
rect 4215 37444 4261 37496
rect 4275 37444 4321 37496
rect 4321 37444 4327 37496
rect 4209 37380 4215 37426
rect 4215 37380 4261 37426
rect 4275 37380 4321 37426
rect 4321 37380 4327 37426
rect 4209 37374 4261 37380
rect 4275 37374 4327 37380
rect 4486 38714 4538 38720
rect 4486 38680 4492 38714
rect 4492 38680 4526 38714
rect 4526 38680 4538 38714
rect 4486 38668 4538 38680
rect 4552 38714 4604 38720
rect 4552 38680 4564 38714
rect 4564 38680 4598 38714
rect 4598 38680 4604 38714
rect 4552 38668 4604 38680
rect 4486 38641 4538 38651
rect 4486 38607 4492 38641
rect 4492 38607 4526 38641
rect 4526 38607 4538 38641
rect 4486 38599 4538 38607
rect 4552 38641 4604 38651
rect 4552 38607 4564 38641
rect 4564 38607 4598 38641
rect 4598 38607 4604 38641
rect 4552 38599 4604 38607
rect 4486 38568 4538 38582
rect 4486 38534 4492 38568
rect 4492 38534 4526 38568
rect 4526 38534 4538 38568
rect 4486 38530 4538 38534
rect 4552 38568 4604 38582
rect 4552 38534 4564 38568
rect 4564 38534 4598 38568
rect 4598 38534 4604 38568
rect 4552 38530 4604 38534
rect 4486 38495 4538 38513
rect 4486 38461 4492 38495
rect 4492 38461 4526 38495
rect 4526 38461 4538 38495
rect 4552 38495 4604 38513
rect 4552 38461 4564 38495
rect 4564 38461 4598 38495
rect 4598 38461 4604 38495
rect 4486 38422 4538 38444
rect 4552 38422 4604 38444
rect 4486 38392 4492 38422
rect 4492 38392 4538 38422
rect 4552 38392 4598 38422
rect 4598 38392 4604 38422
rect 4486 38323 4492 38375
rect 4492 38323 4538 38375
rect 4552 38323 4598 38375
rect 4598 38323 4604 38375
rect 4486 38254 4492 38306
rect 4492 38254 4538 38306
rect 4552 38254 4598 38306
rect 4598 38254 4604 38306
rect 4486 38184 4492 38236
rect 4492 38184 4538 38236
rect 4552 38184 4598 38236
rect 4598 38184 4604 38236
rect 4486 38114 4492 38166
rect 4492 38114 4538 38166
rect 4552 38114 4598 38166
rect 4598 38114 4604 38166
rect 4763 37930 4769 37982
rect 4769 37930 4815 37982
rect 4829 37930 4875 37982
rect 4875 37930 4881 37982
rect 4763 37861 4769 37913
rect 4769 37861 4815 37913
rect 4829 37861 4875 37913
rect 4875 37861 4881 37913
rect 4763 37792 4769 37844
rect 4769 37792 4815 37844
rect 4829 37792 4875 37844
rect 4875 37792 4881 37844
rect 4763 37723 4769 37775
rect 4769 37723 4815 37775
rect 4829 37723 4875 37775
rect 4875 37723 4881 37775
rect 4763 37654 4769 37706
rect 4769 37654 4815 37706
rect 4829 37654 4875 37706
rect 4875 37654 4881 37706
rect 4763 37584 4769 37636
rect 4769 37584 4815 37636
rect 4829 37584 4875 37636
rect 4875 37584 4881 37636
rect 4763 37514 4769 37566
rect 4769 37514 4815 37566
rect 4829 37514 4875 37566
rect 4875 37514 4881 37566
rect 4763 37444 4769 37496
rect 4769 37444 4815 37496
rect 4829 37444 4875 37496
rect 4875 37444 4881 37496
rect 4763 37380 4769 37426
rect 4769 37380 4815 37426
rect 4829 37380 4875 37426
rect 4875 37380 4881 37426
rect 4763 37374 4815 37380
rect 4829 37374 4881 37380
rect 5040 38714 5092 38720
rect 5040 38680 5046 38714
rect 5046 38680 5080 38714
rect 5080 38680 5092 38714
rect 5040 38668 5092 38680
rect 5106 38714 5158 38720
rect 5106 38680 5118 38714
rect 5118 38680 5152 38714
rect 5152 38680 5158 38714
rect 5106 38668 5158 38680
rect 5040 38641 5092 38651
rect 5040 38607 5046 38641
rect 5046 38607 5080 38641
rect 5080 38607 5092 38641
rect 5040 38599 5092 38607
rect 5106 38641 5158 38651
rect 5106 38607 5118 38641
rect 5118 38607 5152 38641
rect 5152 38607 5158 38641
rect 5106 38599 5158 38607
rect 5040 38568 5092 38582
rect 5040 38534 5046 38568
rect 5046 38534 5080 38568
rect 5080 38534 5092 38568
rect 5040 38530 5092 38534
rect 5106 38568 5158 38582
rect 5106 38534 5118 38568
rect 5118 38534 5152 38568
rect 5152 38534 5158 38568
rect 5106 38530 5158 38534
rect 5040 38495 5092 38513
rect 5040 38461 5046 38495
rect 5046 38461 5080 38495
rect 5080 38461 5092 38495
rect 5106 38495 5158 38513
rect 5106 38461 5118 38495
rect 5118 38461 5152 38495
rect 5152 38461 5158 38495
rect 5040 38422 5092 38444
rect 5106 38422 5158 38444
rect 5040 38392 5046 38422
rect 5046 38392 5092 38422
rect 5106 38392 5152 38422
rect 5152 38392 5158 38422
rect 5040 38323 5046 38375
rect 5046 38323 5092 38375
rect 5106 38323 5152 38375
rect 5152 38323 5158 38375
rect 5040 38254 5046 38306
rect 5046 38254 5092 38306
rect 5106 38254 5152 38306
rect 5152 38254 5158 38306
rect 5040 38184 5046 38236
rect 5046 38184 5092 38236
rect 5106 38184 5152 38236
rect 5152 38184 5158 38236
rect 5040 38114 5046 38166
rect 5046 38114 5092 38166
rect 5106 38114 5152 38166
rect 5152 38114 5158 38166
rect 5317 37930 5323 37982
rect 5323 37930 5369 37982
rect 5383 37930 5429 37982
rect 5429 37930 5435 37982
rect 5317 37861 5323 37913
rect 5323 37861 5369 37913
rect 5383 37861 5429 37913
rect 5429 37861 5435 37913
rect 5317 37792 5323 37844
rect 5323 37792 5369 37844
rect 5383 37792 5429 37844
rect 5429 37792 5435 37844
rect 5317 37723 5323 37775
rect 5323 37723 5369 37775
rect 5383 37723 5429 37775
rect 5429 37723 5435 37775
rect 5317 37654 5323 37706
rect 5323 37654 5369 37706
rect 5383 37654 5429 37706
rect 5429 37654 5435 37706
rect 5317 37584 5323 37636
rect 5323 37584 5369 37636
rect 5383 37584 5429 37636
rect 5429 37584 5435 37636
rect 5317 37514 5323 37566
rect 5323 37514 5369 37566
rect 5383 37514 5429 37566
rect 5429 37514 5435 37566
rect 5317 37444 5323 37496
rect 5323 37444 5369 37496
rect 5383 37444 5429 37496
rect 5429 37444 5435 37496
rect 5317 37380 5323 37426
rect 5323 37380 5369 37426
rect 5383 37380 5429 37426
rect 5429 37380 5435 37426
rect 5317 37374 5369 37380
rect 5383 37374 5435 37380
rect 5594 38714 5646 38720
rect 5594 38680 5600 38714
rect 5600 38680 5634 38714
rect 5634 38680 5646 38714
rect 5594 38668 5646 38680
rect 5660 38714 5712 38720
rect 5660 38680 5672 38714
rect 5672 38680 5706 38714
rect 5706 38680 5712 38714
rect 5660 38668 5712 38680
rect 5594 38641 5646 38651
rect 5594 38607 5600 38641
rect 5600 38607 5634 38641
rect 5634 38607 5646 38641
rect 5594 38599 5646 38607
rect 5660 38641 5712 38651
rect 5660 38607 5672 38641
rect 5672 38607 5706 38641
rect 5706 38607 5712 38641
rect 5660 38599 5712 38607
rect 5594 38568 5646 38582
rect 5594 38534 5600 38568
rect 5600 38534 5634 38568
rect 5634 38534 5646 38568
rect 5594 38530 5646 38534
rect 5660 38568 5712 38582
rect 5660 38534 5672 38568
rect 5672 38534 5706 38568
rect 5706 38534 5712 38568
rect 5660 38530 5712 38534
rect 5594 38495 5646 38513
rect 5594 38461 5600 38495
rect 5600 38461 5634 38495
rect 5634 38461 5646 38495
rect 5660 38495 5712 38513
rect 5660 38461 5672 38495
rect 5672 38461 5706 38495
rect 5706 38461 5712 38495
rect 5594 38422 5646 38444
rect 5660 38422 5712 38444
rect 5594 38392 5600 38422
rect 5600 38392 5646 38422
rect 5660 38392 5706 38422
rect 5706 38392 5712 38422
rect 5594 38323 5600 38375
rect 5600 38323 5646 38375
rect 5660 38323 5706 38375
rect 5706 38323 5712 38375
rect 5594 38254 5600 38306
rect 5600 38254 5646 38306
rect 5660 38254 5706 38306
rect 5706 38254 5712 38306
rect 5594 38184 5600 38236
rect 5600 38184 5646 38236
rect 5660 38184 5706 38236
rect 5706 38184 5712 38236
rect 5594 38114 5600 38166
rect 5600 38114 5646 38166
rect 5660 38114 5706 38166
rect 5706 38114 5712 38166
rect 5871 37930 5877 37982
rect 5877 37930 5923 37982
rect 5937 37930 5983 37982
rect 5983 37930 5989 37982
rect 5871 37861 5877 37913
rect 5877 37861 5923 37913
rect 5937 37861 5983 37913
rect 5983 37861 5989 37913
rect 5871 37792 5877 37844
rect 5877 37792 5923 37844
rect 5937 37792 5983 37844
rect 5983 37792 5989 37844
rect 5871 37723 5877 37775
rect 5877 37723 5923 37775
rect 5937 37723 5983 37775
rect 5983 37723 5989 37775
rect 5871 37654 5877 37706
rect 5877 37654 5923 37706
rect 5937 37654 5983 37706
rect 5983 37654 5989 37706
rect 5871 37584 5877 37636
rect 5877 37584 5923 37636
rect 5937 37584 5983 37636
rect 5983 37584 5989 37636
rect 5871 37514 5877 37566
rect 5877 37514 5923 37566
rect 5937 37514 5983 37566
rect 5983 37514 5989 37566
rect 5871 37444 5877 37496
rect 5877 37444 5923 37496
rect 5937 37444 5983 37496
rect 5983 37444 5989 37496
rect 5871 37380 5877 37426
rect 5877 37380 5923 37426
rect 5937 37380 5983 37426
rect 5983 37380 5989 37426
rect 5871 37374 5923 37380
rect 5937 37374 5989 37380
rect 6148 38714 6200 38720
rect 6148 38680 6154 38714
rect 6154 38680 6188 38714
rect 6188 38680 6200 38714
rect 6148 38668 6200 38680
rect 6214 38714 6266 38720
rect 6214 38680 6226 38714
rect 6226 38680 6260 38714
rect 6260 38680 6266 38714
rect 6214 38668 6266 38680
rect 6148 38641 6200 38651
rect 6148 38607 6154 38641
rect 6154 38607 6188 38641
rect 6188 38607 6200 38641
rect 6148 38599 6200 38607
rect 6214 38641 6266 38651
rect 6214 38607 6226 38641
rect 6226 38607 6260 38641
rect 6260 38607 6266 38641
rect 6214 38599 6266 38607
rect 6148 38568 6200 38582
rect 6148 38534 6154 38568
rect 6154 38534 6188 38568
rect 6188 38534 6200 38568
rect 6148 38530 6200 38534
rect 6214 38568 6266 38582
rect 6214 38534 6226 38568
rect 6226 38534 6260 38568
rect 6260 38534 6266 38568
rect 6214 38530 6266 38534
rect 6148 38495 6200 38513
rect 6148 38461 6154 38495
rect 6154 38461 6188 38495
rect 6188 38461 6200 38495
rect 6214 38495 6266 38513
rect 6214 38461 6226 38495
rect 6226 38461 6260 38495
rect 6260 38461 6266 38495
rect 6148 38422 6200 38444
rect 6214 38422 6266 38444
rect 6148 38392 6154 38422
rect 6154 38392 6200 38422
rect 6214 38392 6260 38422
rect 6260 38392 6266 38422
rect 6148 38323 6154 38375
rect 6154 38323 6200 38375
rect 6214 38323 6260 38375
rect 6260 38323 6266 38375
rect 6148 38254 6154 38306
rect 6154 38254 6200 38306
rect 6214 38254 6260 38306
rect 6260 38254 6266 38306
rect 6148 38184 6154 38236
rect 6154 38184 6200 38236
rect 6214 38184 6260 38236
rect 6260 38184 6266 38236
rect 6148 38114 6154 38166
rect 6154 38114 6200 38166
rect 6214 38114 6260 38166
rect 6260 38114 6266 38166
rect 6425 37930 6431 37982
rect 6431 37930 6477 37982
rect 6491 37930 6537 37982
rect 6537 37930 6543 37982
rect 6425 37861 6431 37913
rect 6431 37861 6477 37913
rect 6491 37861 6537 37913
rect 6537 37861 6543 37913
rect 6425 37792 6431 37844
rect 6431 37792 6477 37844
rect 6491 37792 6537 37844
rect 6537 37792 6543 37844
rect 6425 37723 6431 37775
rect 6431 37723 6477 37775
rect 6491 37723 6537 37775
rect 6537 37723 6543 37775
rect 6425 37654 6431 37706
rect 6431 37654 6477 37706
rect 6491 37654 6537 37706
rect 6537 37654 6543 37706
rect 6425 37584 6431 37636
rect 6431 37584 6477 37636
rect 6491 37584 6537 37636
rect 6537 37584 6543 37636
rect 6425 37514 6431 37566
rect 6431 37514 6477 37566
rect 6491 37514 6537 37566
rect 6537 37514 6543 37566
rect 6425 37444 6431 37496
rect 6431 37444 6477 37496
rect 6491 37444 6537 37496
rect 6537 37444 6543 37496
rect 6425 37380 6431 37426
rect 6431 37380 6477 37426
rect 6491 37380 6537 37426
rect 6537 37380 6543 37426
rect 6425 37374 6477 37380
rect 6491 37374 6543 37380
rect 6702 38714 6754 38720
rect 6702 38680 6708 38714
rect 6708 38680 6742 38714
rect 6742 38680 6754 38714
rect 6702 38668 6754 38680
rect 6768 38714 6820 38720
rect 6768 38680 6780 38714
rect 6780 38680 6814 38714
rect 6814 38680 6820 38714
rect 6768 38668 6820 38680
rect 6702 38641 6754 38651
rect 6702 38607 6708 38641
rect 6708 38607 6742 38641
rect 6742 38607 6754 38641
rect 6702 38599 6754 38607
rect 6768 38641 6820 38651
rect 6768 38607 6780 38641
rect 6780 38607 6814 38641
rect 6814 38607 6820 38641
rect 6768 38599 6820 38607
rect 6702 38568 6754 38582
rect 6702 38534 6708 38568
rect 6708 38534 6742 38568
rect 6742 38534 6754 38568
rect 6702 38530 6754 38534
rect 6768 38568 6820 38582
rect 6768 38534 6780 38568
rect 6780 38534 6814 38568
rect 6814 38534 6820 38568
rect 6768 38530 6820 38534
rect 6702 38495 6754 38513
rect 6702 38461 6708 38495
rect 6708 38461 6742 38495
rect 6742 38461 6754 38495
rect 6768 38495 6820 38513
rect 6768 38461 6780 38495
rect 6780 38461 6814 38495
rect 6814 38461 6820 38495
rect 6702 38422 6754 38444
rect 6768 38422 6820 38444
rect 6702 38392 6708 38422
rect 6708 38392 6754 38422
rect 6768 38392 6814 38422
rect 6814 38392 6820 38422
rect 6702 38323 6708 38375
rect 6708 38323 6754 38375
rect 6768 38323 6814 38375
rect 6814 38323 6820 38375
rect 6702 38254 6708 38306
rect 6708 38254 6754 38306
rect 6768 38254 6814 38306
rect 6814 38254 6820 38306
rect 6702 38184 6708 38236
rect 6708 38184 6754 38236
rect 6768 38184 6814 38236
rect 6814 38184 6820 38236
rect 6702 38114 6708 38166
rect 6708 38114 6754 38166
rect 6768 38114 6814 38166
rect 6814 38114 6820 38166
rect 6979 37930 6985 37982
rect 6985 37930 7031 37982
rect 7045 37930 7091 37982
rect 7091 37930 7097 37982
rect 6979 37861 6985 37913
rect 6985 37861 7031 37913
rect 7045 37861 7091 37913
rect 7091 37861 7097 37913
rect 6979 37792 6985 37844
rect 6985 37792 7031 37844
rect 7045 37792 7091 37844
rect 7091 37792 7097 37844
rect 6979 37723 6985 37775
rect 6985 37723 7031 37775
rect 7045 37723 7091 37775
rect 7091 37723 7097 37775
rect 6979 37654 6985 37706
rect 6985 37654 7031 37706
rect 7045 37654 7091 37706
rect 7091 37654 7097 37706
rect 6979 37584 6985 37636
rect 6985 37584 7031 37636
rect 7045 37584 7091 37636
rect 7091 37584 7097 37636
rect 6979 37514 6985 37566
rect 6985 37514 7031 37566
rect 7045 37514 7091 37566
rect 7091 37514 7097 37566
rect 6979 37444 6985 37496
rect 6985 37444 7031 37496
rect 7045 37444 7091 37496
rect 7091 37444 7097 37496
rect 6979 37380 6985 37426
rect 6985 37380 7031 37426
rect 7045 37380 7091 37426
rect 7091 37380 7097 37426
rect 6979 37374 7031 37380
rect 7045 37374 7097 37380
rect 7256 38714 7308 38720
rect 7256 38680 7262 38714
rect 7262 38680 7296 38714
rect 7296 38680 7308 38714
rect 7256 38668 7308 38680
rect 7322 38714 7374 38720
rect 7322 38680 7334 38714
rect 7334 38680 7368 38714
rect 7368 38680 7374 38714
rect 7322 38668 7374 38680
rect 7256 38641 7308 38651
rect 7256 38607 7262 38641
rect 7262 38607 7296 38641
rect 7296 38607 7308 38641
rect 7256 38599 7308 38607
rect 7322 38641 7374 38651
rect 7322 38607 7334 38641
rect 7334 38607 7368 38641
rect 7368 38607 7374 38641
rect 7322 38599 7374 38607
rect 7256 38568 7308 38582
rect 7256 38534 7262 38568
rect 7262 38534 7296 38568
rect 7296 38534 7308 38568
rect 7256 38530 7308 38534
rect 7322 38568 7374 38582
rect 7322 38534 7334 38568
rect 7334 38534 7368 38568
rect 7368 38534 7374 38568
rect 7322 38530 7374 38534
rect 7256 38495 7308 38513
rect 7256 38461 7262 38495
rect 7262 38461 7296 38495
rect 7296 38461 7308 38495
rect 7322 38495 7374 38513
rect 7322 38461 7334 38495
rect 7334 38461 7368 38495
rect 7368 38461 7374 38495
rect 7256 38422 7308 38444
rect 7322 38422 7374 38444
rect 7256 38392 7262 38422
rect 7262 38392 7308 38422
rect 7322 38392 7368 38422
rect 7368 38392 7374 38422
rect 7256 38323 7262 38375
rect 7262 38323 7308 38375
rect 7322 38323 7368 38375
rect 7368 38323 7374 38375
rect 7256 38254 7262 38306
rect 7262 38254 7308 38306
rect 7322 38254 7368 38306
rect 7368 38254 7374 38306
rect 7256 38184 7262 38236
rect 7262 38184 7308 38236
rect 7322 38184 7368 38236
rect 7368 38184 7374 38236
rect 7256 38114 7262 38166
rect 7262 38114 7308 38166
rect 7322 38114 7368 38166
rect 7368 38114 7374 38166
rect 7533 37930 7539 37982
rect 7539 37930 7585 37982
rect 7599 37930 7645 37982
rect 7645 37930 7651 37982
rect 7533 37861 7539 37913
rect 7539 37861 7585 37913
rect 7599 37861 7645 37913
rect 7645 37861 7651 37913
rect 7533 37792 7539 37844
rect 7539 37792 7585 37844
rect 7599 37792 7645 37844
rect 7645 37792 7651 37844
rect 7533 37723 7539 37775
rect 7539 37723 7585 37775
rect 7599 37723 7645 37775
rect 7645 37723 7651 37775
rect 7533 37654 7539 37706
rect 7539 37654 7585 37706
rect 7599 37654 7645 37706
rect 7645 37654 7651 37706
rect 7533 37584 7539 37636
rect 7539 37584 7585 37636
rect 7599 37584 7645 37636
rect 7645 37584 7651 37636
rect 7533 37514 7539 37566
rect 7539 37514 7585 37566
rect 7599 37514 7645 37566
rect 7645 37514 7651 37566
rect 7533 37444 7539 37496
rect 7539 37444 7585 37496
rect 7599 37444 7645 37496
rect 7645 37444 7651 37496
rect 7533 37380 7539 37426
rect 7539 37380 7585 37426
rect 7599 37380 7645 37426
rect 7645 37380 7651 37426
rect 7533 37374 7585 37380
rect 7599 37374 7651 37380
rect 7810 38714 7862 38720
rect 7810 38680 7816 38714
rect 7816 38680 7850 38714
rect 7850 38680 7862 38714
rect 7810 38668 7862 38680
rect 7876 38714 7928 38720
rect 7876 38680 7888 38714
rect 7888 38680 7922 38714
rect 7922 38680 7928 38714
rect 7876 38668 7928 38680
rect 7810 38641 7862 38651
rect 7810 38607 7816 38641
rect 7816 38607 7850 38641
rect 7850 38607 7862 38641
rect 7810 38599 7862 38607
rect 7876 38641 7928 38651
rect 7876 38607 7888 38641
rect 7888 38607 7922 38641
rect 7922 38607 7928 38641
rect 7876 38599 7928 38607
rect 7810 38568 7862 38582
rect 7810 38534 7816 38568
rect 7816 38534 7850 38568
rect 7850 38534 7862 38568
rect 7810 38530 7862 38534
rect 7876 38568 7928 38582
rect 7876 38534 7888 38568
rect 7888 38534 7922 38568
rect 7922 38534 7928 38568
rect 7876 38530 7928 38534
rect 7810 38495 7862 38513
rect 7810 38461 7816 38495
rect 7816 38461 7850 38495
rect 7850 38461 7862 38495
rect 7876 38495 7928 38513
rect 7876 38461 7888 38495
rect 7888 38461 7922 38495
rect 7922 38461 7928 38495
rect 7810 38422 7862 38444
rect 7876 38422 7928 38444
rect 7810 38392 7816 38422
rect 7816 38392 7862 38422
rect 7876 38392 7922 38422
rect 7922 38392 7928 38422
rect 7810 38323 7816 38375
rect 7816 38323 7862 38375
rect 7876 38323 7922 38375
rect 7922 38323 7928 38375
rect 7810 38254 7816 38306
rect 7816 38254 7862 38306
rect 7876 38254 7922 38306
rect 7922 38254 7928 38306
rect 7810 38184 7816 38236
rect 7816 38184 7862 38236
rect 7876 38184 7922 38236
rect 7922 38184 7928 38236
rect 7810 38114 7816 38166
rect 7816 38114 7862 38166
rect 7876 38114 7922 38166
rect 7922 38114 7928 38166
rect 8047 38719 8099 38724
rect 8047 38685 8050 38719
rect 8050 38685 8084 38719
rect 8084 38685 8099 38719
rect 8047 38672 8099 38685
rect 8169 38709 8221 38724
rect 8169 38675 8184 38709
rect 8184 38675 8218 38709
rect 8218 38675 8221 38709
rect 8169 38672 8221 38675
rect 8047 38647 8099 38655
rect 8047 38613 8050 38647
rect 8050 38613 8084 38647
rect 8084 38613 8099 38647
rect 8047 38603 8099 38613
rect 8169 38637 8221 38655
rect 8169 38603 8184 38637
rect 8184 38603 8218 38637
rect 8218 38603 8221 38637
rect 8047 38575 8099 38586
rect 8047 38541 8050 38575
rect 8050 38541 8084 38575
rect 8084 38541 8099 38575
rect 8047 38534 8099 38541
rect 8169 38565 8221 38586
rect 8169 38534 8184 38565
rect 8184 38534 8218 38565
rect 8218 38534 8221 38565
rect 8047 38503 8099 38517
rect 8047 38469 8050 38503
rect 8050 38469 8084 38503
rect 8084 38469 8099 38503
rect 8047 38465 8099 38469
rect 8169 38493 8221 38517
rect 8169 38465 8184 38493
rect 8184 38465 8218 38493
rect 8218 38465 8221 38493
rect 8047 38431 8099 38448
rect 8047 38397 8050 38431
rect 8050 38397 8084 38431
rect 8084 38397 8099 38431
rect 8047 38396 8099 38397
rect 8169 38421 8221 38448
rect 8169 38396 8184 38421
rect 8184 38396 8218 38421
rect 8218 38396 8221 38421
rect 8047 38359 8099 38378
rect 8047 38326 8050 38359
rect 8050 38326 8084 38359
rect 8084 38326 8099 38359
rect 8169 38349 8221 38378
rect 8169 38326 8184 38349
rect 8184 38326 8218 38349
rect 8218 38326 8221 38349
rect 8047 38287 8099 38308
rect 8047 38256 8050 38287
rect 8050 38256 8084 38287
rect 8084 38256 8099 38287
rect 8169 38277 8221 38308
rect 8169 38256 8184 38277
rect 8184 38256 8218 38277
rect 8218 38256 8221 38277
rect 8047 38215 8099 38238
rect 8047 38186 8050 38215
rect 8050 38186 8084 38215
rect 8084 38186 8099 38215
rect 8169 38205 8221 38238
rect 8169 38186 8184 38205
rect 8184 38186 8218 38205
rect 8218 38186 8221 38205
rect 8047 38143 8099 38168
rect 8047 38116 8050 38143
rect 8050 38116 8084 38143
rect 8084 38116 8099 38143
rect 8169 38133 8221 38168
rect 8169 38116 8184 38133
rect 8184 38116 8218 38133
rect 8218 38116 8221 38133
rect 2824 36714 2876 36720
rect 2824 36680 2830 36714
rect 2830 36680 2864 36714
rect 2864 36680 2876 36714
rect 2824 36668 2876 36680
rect 2890 36714 2942 36720
rect 2890 36680 2902 36714
rect 2902 36680 2936 36714
rect 2936 36680 2942 36714
rect 2890 36668 2942 36680
rect 2824 36641 2876 36651
rect 2824 36607 2830 36641
rect 2830 36607 2864 36641
rect 2864 36607 2876 36641
rect 2824 36599 2876 36607
rect 2890 36641 2942 36651
rect 2890 36607 2902 36641
rect 2902 36607 2936 36641
rect 2936 36607 2942 36641
rect 2890 36599 2942 36607
rect 2824 36568 2876 36582
rect 2824 36534 2830 36568
rect 2830 36534 2864 36568
rect 2864 36534 2876 36568
rect 2824 36530 2876 36534
rect 2890 36568 2942 36582
rect 2890 36534 2902 36568
rect 2902 36534 2936 36568
rect 2936 36534 2942 36568
rect 2890 36530 2942 36534
rect 2824 36495 2876 36513
rect 2824 36461 2830 36495
rect 2830 36461 2864 36495
rect 2864 36461 2876 36495
rect 2890 36495 2942 36513
rect 2890 36461 2902 36495
rect 2902 36461 2936 36495
rect 2936 36461 2942 36495
rect 2824 36422 2876 36444
rect 2890 36422 2942 36444
rect 2824 36392 2830 36422
rect 2830 36392 2876 36422
rect 2890 36392 2936 36422
rect 2936 36392 2942 36422
rect 2824 36323 2830 36375
rect 2830 36323 2876 36375
rect 2890 36323 2936 36375
rect 2936 36323 2942 36375
rect 2824 36254 2830 36306
rect 2830 36254 2876 36306
rect 2890 36254 2936 36306
rect 2936 36254 2942 36306
rect 2824 36184 2830 36236
rect 2830 36184 2876 36236
rect 2890 36184 2936 36236
rect 2936 36184 2942 36236
rect 2824 36114 2830 36166
rect 2830 36114 2876 36166
rect 2890 36114 2936 36166
rect 2936 36114 2942 36166
rect 3101 35930 3107 35982
rect 3107 35930 3153 35982
rect 3167 35930 3213 35982
rect 3213 35930 3219 35982
rect 3101 35861 3107 35913
rect 3107 35861 3153 35913
rect 3167 35861 3213 35913
rect 3213 35861 3219 35913
rect 3101 35792 3107 35844
rect 3107 35792 3153 35844
rect 3167 35792 3213 35844
rect 3213 35792 3219 35844
rect 3101 35723 3107 35775
rect 3107 35723 3153 35775
rect 3167 35723 3213 35775
rect 3213 35723 3219 35775
rect 3101 35654 3107 35706
rect 3107 35654 3153 35706
rect 3167 35654 3213 35706
rect 3213 35654 3219 35706
rect 3101 35584 3107 35636
rect 3107 35584 3153 35636
rect 3167 35584 3213 35636
rect 3213 35584 3219 35636
rect 3101 35514 3107 35566
rect 3107 35514 3153 35566
rect 3167 35514 3213 35566
rect 3213 35514 3219 35566
rect 3101 35444 3107 35496
rect 3107 35444 3153 35496
rect 3167 35444 3213 35496
rect 3213 35444 3219 35496
rect 3101 35380 3107 35426
rect 3107 35380 3153 35426
rect 3167 35380 3213 35426
rect 3213 35380 3219 35426
rect 3101 35374 3153 35380
rect 3167 35374 3219 35380
rect 3378 36714 3430 36720
rect 3378 36680 3384 36714
rect 3384 36680 3418 36714
rect 3418 36680 3430 36714
rect 3378 36668 3430 36680
rect 3444 36714 3496 36720
rect 3444 36680 3456 36714
rect 3456 36680 3490 36714
rect 3490 36680 3496 36714
rect 3444 36668 3496 36680
rect 3378 36641 3430 36651
rect 3378 36607 3384 36641
rect 3384 36607 3418 36641
rect 3418 36607 3430 36641
rect 3378 36599 3430 36607
rect 3444 36641 3496 36651
rect 3444 36607 3456 36641
rect 3456 36607 3490 36641
rect 3490 36607 3496 36641
rect 3444 36599 3496 36607
rect 3378 36568 3430 36582
rect 3378 36534 3384 36568
rect 3384 36534 3418 36568
rect 3418 36534 3430 36568
rect 3378 36530 3430 36534
rect 3444 36568 3496 36582
rect 3444 36534 3456 36568
rect 3456 36534 3490 36568
rect 3490 36534 3496 36568
rect 3444 36530 3496 36534
rect 3378 36495 3430 36513
rect 3378 36461 3384 36495
rect 3384 36461 3418 36495
rect 3418 36461 3430 36495
rect 3444 36495 3496 36513
rect 3444 36461 3456 36495
rect 3456 36461 3490 36495
rect 3490 36461 3496 36495
rect 3378 36422 3430 36444
rect 3444 36422 3496 36444
rect 3378 36392 3384 36422
rect 3384 36392 3430 36422
rect 3444 36392 3490 36422
rect 3490 36392 3496 36422
rect 3378 36323 3384 36375
rect 3384 36323 3430 36375
rect 3444 36323 3490 36375
rect 3490 36323 3496 36375
rect 3378 36254 3384 36306
rect 3384 36254 3430 36306
rect 3444 36254 3490 36306
rect 3490 36254 3496 36306
rect 3378 36184 3384 36236
rect 3384 36184 3430 36236
rect 3444 36184 3490 36236
rect 3490 36184 3496 36236
rect 3378 36114 3384 36166
rect 3384 36114 3430 36166
rect 3444 36114 3490 36166
rect 3490 36114 3496 36166
rect 3655 35930 3661 35982
rect 3661 35930 3707 35982
rect 3721 35930 3767 35982
rect 3767 35930 3773 35982
rect 3655 35861 3661 35913
rect 3661 35861 3707 35913
rect 3721 35861 3767 35913
rect 3767 35861 3773 35913
rect 3655 35792 3661 35844
rect 3661 35792 3707 35844
rect 3721 35792 3767 35844
rect 3767 35792 3773 35844
rect 3655 35723 3661 35775
rect 3661 35723 3707 35775
rect 3721 35723 3767 35775
rect 3767 35723 3773 35775
rect 3655 35654 3661 35706
rect 3661 35654 3707 35706
rect 3721 35654 3767 35706
rect 3767 35654 3773 35706
rect 3655 35584 3661 35636
rect 3661 35584 3707 35636
rect 3721 35584 3767 35636
rect 3767 35584 3773 35636
rect 3655 35514 3661 35566
rect 3661 35514 3707 35566
rect 3721 35514 3767 35566
rect 3767 35514 3773 35566
rect 3655 35444 3661 35496
rect 3661 35444 3707 35496
rect 3721 35444 3767 35496
rect 3767 35444 3773 35496
rect 3655 35380 3661 35426
rect 3661 35380 3707 35426
rect 3721 35380 3767 35426
rect 3767 35380 3773 35426
rect 3655 35374 3707 35380
rect 3721 35374 3773 35380
rect 3932 36714 3984 36720
rect 3932 36680 3938 36714
rect 3938 36680 3972 36714
rect 3972 36680 3984 36714
rect 3932 36668 3984 36680
rect 3998 36714 4050 36720
rect 3998 36680 4010 36714
rect 4010 36680 4044 36714
rect 4044 36680 4050 36714
rect 3998 36668 4050 36680
rect 3932 36641 3984 36651
rect 3932 36607 3938 36641
rect 3938 36607 3972 36641
rect 3972 36607 3984 36641
rect 3932 36599 3984 36607
rect 3998 36641 4050 36651
rect 3998 36607 4010 36641
rect 4010 36607 4044 36641
rect 4044 36607 4050 36641
rect 3998 36599 4050 36607
rect 3932 36568 3984 36582
rect 3932 36534 3938 36568
rect 3938 36534 3972 36568
rect 3972 36534 3984 36568
rect 3932 36530 3984 36534
rect 3998 36568 4050 36582
rect 3998 36534 4010 36568
rect 4010 36534 4044 36568
rect 4044 36534 4050 36568
rect 3998 36530 4050 36534
rect 3932 36495 3984 36513
rect 3932 36461 3938 36495
rect 3938 36461 3972 36495
rect 3972 36461 3984 36495
rect 3998 36495 4050 36513
rect 3998 36461 4010 36495
rect 4010 36461 4044 36495
rect 4044 36461 4050 36495
rect 3932 36422 3984 36444
rect 3998 36422 4050 36444
rect 3932 36392 3938 36422
rect 3938 36392 3984 36422
rect 3998 36392 4044 36422
rect 4044 36392 4050 36422
rect 3932 36323 3938 36375
rect 3938 36323 3984 36375
rect 3998 36323 4044 36375
rect 4044 36323 4050 36375
rect 3932 36254 3938 36306
rect 3938 36254 3984 36306
rect 3998 36254 4044 36306
rect 4044 36254 4050 36306
rect 3932 36184 3938 36236
rect 3938 36184 3984 36236
rect 3998 36184 4044 36236
rect 4044 36184 4050 36236
rect 3932 36114 3938 36166
rect 3938 36114 3984 36166
rect 3998 36114 4044 36166
rect 4044 36114 4050 36166
rect 4209 35930 4215 35982
rect 4215 35930 4261 35982
rect 4275 35930 4321 35982
rect 4321 35930 4327 35982
rect 4209 35861 4215 35913
rect 4215 35861 4261 35913
rect 4275 35861 4321 35913
rect 4321 35861 4327 35913
rect 4209 35792 4215 35844
rect 4215 35792 4261 35844
rect 4275 35792 4321 35844
rect 4321 35792 4327 35844
rect 4209 35723 4215 35775
rect 4215 35723 4261 35775
rect 4275 35723 4321 35775
rect 4321 35723 4327 35775
rect 4209 35654 4215 35706
rect 4215 35654 4261 35706
rect 4275 35654 4321 35706
rect 4321 35654 4327 35706
rect 4209 35584 4215 35636
rect 4215 35584 4261 35636
rect 4275 35584 4321 35636
rect 4321 35584 4327 35636
rect 4209 35514 4215 35566
rect 4215 35514 4261 35566
rect 4275 35514 4321 35566
rect 4321 35514 4327 35566
rect 4209 35444 4215 35496
rect 4215 35444 4261 35496
rect 4275 35444 4321 35496
rect 4321 35444 4327 35496
rect 4209 35380 4215 35426
rect 4215 35380 4261 35426
rect 4275 35380 4321 35426
rect 4321 35380 4327 35426
rect 4209 35374 4261 35380
rect 4275 35374 4327 35380
rect 4486 36714 4538 36720
rect 4486 36680 4492 36714
rect 4492 36680 4526 36714
rect 4526 36680 4538 36714
rect 4486 36668 4538 36680
rect 4552 36714 4604 36720
rect 4552 36680 4564 36714
rect 4564 36680 4598 36714
rect 4598 36680 4604 36714
rect 4552 36668 4604 36680
rect 4486 36641 4538 36651
rect 4486 36607 4492 36641
rect 4492 36607 4526 36641
rect 4526 36607 4538 36641
rect 4486 36599 4538 36607
rect 4552 36641 4604 36651
rect 4552 36607 4564 36641
rect 4564 36607 4598 36641
rect 4598 36607 4604 36641
rect 4552 36599 4604 36607
rect 4486 36568 4538 36582
rect 4486 36534 4492 36568
rect 4492 36534 4526 36568
rect 4526 36534 4538 36568
rect 4486 36530 4538 36534
rect 4552 36568 4604 36582
rect 4552 36534 4564 36568
rect 4564 36534 4598 36568
rect 4598 36534 4604 36568
rect 4552 36530 4604 36534
rect 4486 36495 4538 36513
rect 4486 36461 4492 36495
rect 4492 36461 4526 36495
rect 4526 36461 4538 36495
rect 4552 36495 4604 36513
rect 4552 36461 4564 36495
rect 4564 36461 4598 36495
rect 4598 36461 4604 36495
rect 4486 36422 4538 36444
rect 4552 36422 4604 36444
rect 4486 36392 4492 36422
rect 4492 36392 4538 36422
rect 4552 36392 4598 36422
rect 4598 36392 4604 36422
rect 4486 36323 4492 36375
rect 4492 36323 4538 36375
rect 4552 36323 4598 36375
rect 4598 36323 4604 36375
rect 4486 36254 4492 36306
rect 4492 36254 4538 36306
rect 4552 36254 4598 36306
rect 4598 36254 4604 36306
rect 4486 36184 4492 36236
rect 4492 36184 4538 36236
rect 4552 36184 4598 36236
rect 4598 36184 4604 36236
rect 4486 36114 4492 36166
rect 4492 36114 4538 36166
rect 4552 36114 4598 36166
rect 4598 36114 4604 36166
rect 4763 35930 4769 35982
rect 4769 35930 4815 35982
rect 4829 35930 4875 35982
rect 4875 35930 4881 35982
rect 4763 35861 4769 35913
rect 4769 35861 4815 35913
rect 4829 35861 4875 35913
rect 4875 35861 4881 35913
rect 4763 35792 4769 35844
rect 4769 35792 4815 35844
rect 4829 35792 4875 35844
rect 4875 35792 4881 35844
rect 4763 35723 4769 35775
rect 4769 35723 4815 35775
rect 4829 35723 4875 35775
rect 4875 35723 4881 35775
rect 4763 35654 4769 35706
rect 4769 35654 4815 35706
rect 4829 35654 4875 35706
rect 4875 35654 4881 35706
rect 4763 35584 4769 35636
rect 4769 35584 4815 35636
rect 4829 35584 4875 35636
rect 4875 35584 4881 35636
rect 4763 35514 4769 35566
rect 4769 35514 4815 35566
rect 4829 35514 4875 35566
rect 4875 35514 4881 35566
rect 4763 35444 4769 35496
rect 4769 35444 4815 35496
rect 4829 35444 4875 35496
rect 4875 35444 4881 35496
rect 4763 35380 4769 35426
rect 4769 35380 4815 35426
rect 4829 35380 4875 35426
rect 4875 35380 4881 35426
rect 4763 35374 4815 35380
rect 4829 35374 4881 35380
rect 5040 36714 5092 36720
rect 5040 36680 5046 36714
rect 5046 36680 5080 36714
rect 5080 36680 5092 36714
rect 5040 36668 5092 36680
rect 5106 36714 5158 36720
rect 5106 36680 5118 36714
rect 5118 36680 5152 36714
rect 5152 36680 5158 36714
rect 5106 36668 5158 36680
rect 5040 36641 5092 36651
rect 5040 36607 5046 36641
rect 5046 36607 5080 36641
rect 5080 36607 5092 36641
rect 5040 36599 5092 36607
rect 5106 36641 5158 36651
rect 5106 36607 5118 36641
rect 5118 36607 5152 36641
rect 5152 36607 5158 36641
rect 5106 36599 5158 36607
rect 5040 36568 5092 36582
rect 5040 36534 5046 36568
rect 5046 36534 5080 36568
rect 5080 36534 5092 36568
rect 5040 36530 5092 36534
rect 5106 36568 5158 36582
rect 5106 36534 5118 36568
rect 5118 36534 5152 36568
rect 5152 36534 5158 36568
rect 5106 36530 5158 36534
rect 5040 36495 5092 36513
rect 5040 36461 5046 36495
rect 5046 36461 5080 36495
rect 5080 36461 5092 36495
rect 5106 36495 5158 36513
rect 5106 36461 5118 36495
rect 5118 36461 5152 36495
rect 5152 36461 5158 36495
rect 5040 36422 5092 36444
rect 5106 36422 5158 36444
rect 5040 36392 5046 36422
rect 5046 36392 5092 36422
rect 5106 36392 5152 36422
rect 5152 36392 5158 36422
rect 5040 36323 5046 36375
rect 5046 36323 5092 36375
rect 5106 36323 5152 36375
rect 5152 36323 5158 36375
rect 5040 36254 5046 36306
rect 5046 36254 5092 36306
rect 5106 36254 5152 36306
rect 5152 36254 5158 36306
rect 5040 36184 5046 36236
rect 5046 36184 5092 36236
rect 5106 36184 5152 36236
rect 5152 36184 5158 36236
rect 5040 36114 5046 36166
rect 5046 36114 5092 36166
rect 5106 36114 5152 36166
rect 5152 36114 5158 36166
rect 5317 35930 5323 35982
rect 5323 35930 5369 35982
rect 5383 35930 5429 35982
rect 5429 35930 5435 35982
rect 5317 35861 5323 35913
rect 5323 35861 5369 35913
rect 5383 35861 5429 35913
rect 5429 35861 5435 35913
rect 5317 35792 5323 35844
rect 5323 35792 5369 35844
rect 5383 35792 5429 35844
rect 5429 35792 5435 35844
rect 5317 35723 5323 35775
rect 5323 35723 5369 35775
rect 5383 35723 5429 35775
rect 5429 35723 5435 35775
rect 5317 35654 5323 35706
rect 5323 35654 5369 35706
rect 5383 35654 5429 35706
rect 5429 35654 5435 35706
rect 5317 35584 5323 35636
rect 5323 35584 5369 35636
rect 5383 35584 5429 35636
rect 5429 35584 5435 35636
rect 5317 35514 5323 35566
rect 5323 35514 5369 35566
rect 5383 35514 5429 35566
rect 5429 35514 5435 35566
rect 5317 35444 5323 35496
rect 5323 35444 5369 35496
rect 5383 35444 5429 35496
rect 5429 35444 5435 35496
rect 5317 35380 5323 35426
rect 5323 35380 5369 35426
rect 5383 35380 5429 35426
rect 5429 35380 5435 35426
rect 5317 35374 5369 35380
rect 5383 35374 5435 35380
rect 5594 36714 5646 36720
rect 5594 36680 5600 36714
rect 5600 36680 5634 36714
rect 5634 36680 5646 36714
rect 5594 36668 5646 36680
rect 5660 36714 5712 36720
rect 5660 36680 5672 36714
rect 5672 36680 5706 36714
rect 5706 36680 5712 36714
rect 5660 36668 5712 36680
rect 5594 36641 5646 36651
rect 5594 36607 5600 36641
rect 5600 36607 5634 36641
rect 5634 36607 5646 36641
rect 5594 36599 5646 36607
rect 5660 36641 5712 36651
rect 5660 36607 5672 36641
rect 5672 36607 5706 36641
rect 5706 36607 5712 36641
rect 5660 36599 5712 36607
rect 5594 36568 5646 36582
rect 5594 36534 5600 36568
rect 5600 36534 5634 36568
rect 5634 36534 5646 36568
rect 5594 36530 5646 36534
rect 5660 36568 5712 36582
rect 5660 36534 5672 36568
rect 5672 36534 5706 36568
rect 5706 36534 5712 36568
rect 5660 36530 5712 36534
rect 5594 36495 5646 36513
rect 5594 36461 5600 36495
rect 5600 36461 5634 36495
rect 5634 36461 5646 36495
rect 5660 36495 5712 36513
rect 5660 36461 5672 36495
rect 5672 36461 5706 36495
rect 5706 36461 5712 36495
rect 5594 36422 5646 36444
rect 5660 36422 5712 36444
rect 5594 36392 5600 36422
rect 5600 36392 5646 36422
rect 5660 36392 5706 36422
rect 5706 36392 5712 36422
rect 5594 36323 5600 36375
rect 5600 36323 5646 36375
rect 5660 36323 5706 36375
rect 5706 36323 5712 36375
rect 5594 36254 5600 36306
rect 5600 36254 5646 36306
rect 5660 36254 5706 36306
rect 5706 36254 5712 36306
rect 5594 36184 5600 36236
rect 5600 36184 5646 36236
rect 5660 36184 5706 36236
rect 5706 36184 5712 36236
rect 5594 36114 5600 36166
rect 5600 36114 5646 36166
rect 5660 36114 5706 36166
rect 5706 36114 5712 36166
rect 5871 35930 5877 35982
rect 5877 35930 5923 35982
rect 5937 35930 5983 35982
rect 5983 35930 5989 35982
rect 5871 35861 5877 35913
rect 5877 35861 5923 35913
rect 5937 35861 5983 35913
rect 5983 35861 5989 35913
rect 5871 35792 5877 35844
rect 5877 35792 5923 35844
rect 5937 35792 5983 35844
rect 5983 35792 5989 35844
rect 5871 35723 5877 35775
rect 5877 35723 5923 35775
rect 5937 35723 5983 35775
rect 5983 35723 5989 35775
rect 5871 35654 5877 35706
rect 5877 35654 5923 35706
rect 5937 35654 5983 35706
rect 5983 35654 5989 35706
rect 5871 35584 5877 35636
rect 5877 35584 5923 35636
rect 5937 35584 5983 35636
rect 5983 35584 5989 35636
rect 5871 35514 5877 35566
rect 5877 35514 5923 35566
rect 5937 35514 5983 35566
rect 5983 35514 5989 35566
rect 5871 35444 5877 35496
rect 5877 35444 5923 35496
rect 5937 35444 5983 35496
rect 5983 35444 5989 35496
rect 5871 35380 5877 35426
rect 5877 35380 5923 35426
rect 5937 35380 5983 35426
rect 5983 35380 5989 35426
rect 5871 35374 5923 35380
rect 5937 35374 5989 35380
rect 6148 36714 6200 36720
rect 6148 36680 6154 36714
rect 6154 36680 6188 36714
rect 6188 36680 6200 36714
rect 6148 36668 6200 36680
rect 6214 36714 6266 36720
rect 6214 36680 6226 36714
rect 6226 36680 6260 36714
rect 6260 36680 6266 36714
rect 6214 36668 6266 36680
rect 6148 36641 6200 36651
rect 6148 36607 6154 36641
rect 6154 36607 6188 36641
rect 6188 36607 6200 36641
rect 6148 36599 6200 36607
rect 6214 36641 6266 36651
rect 6214 36607 6226 36641
rect 6226 36607 6260 36641
rect 6260 36607 6266 36641
rect 6214 36599 6266 36607
rect 6148 36568 6200 36582
rect 6148 36534 6154 36568
rect 6154 36534 6188 36568
rect 6188 36534 6200 36568
rect 6148 36530 6200 36534
rect 6214 36568 6266 36582
rect 6214 36534 6226 36568
rect 6226 36534 6260 36568
rect 6260 36534 6266 36568
rect 6214 36530 6266 36534
rect 6148 36495 6200 36513
rect 6148 36461 6154 36495
rect 6154 36461 6188 36495
rect 6188 36461 6200 36495
rect 6214 36495 6266 36513
rect 6214 36461 6226 36495
rect 6226 36461 6260 36495
rect 6260 36461 6266 36495
rect 6148 36422 6200 36444
rect 6214 36422 6266 36444
rect 6148 36392 6154 36422
rect 6154 36392 6200 36422
rect 6214 36392 6260 36422
rect 6260 36392 6266 36422
rect 6148 36323 6154 36375
rect 6154 36323 6200 36375
rect 6214 36323 6260 36375
rect 6260 36323 6266 36375
rect 6148 36254 6154 36306
rect 6154 36254 6200 36306
rect 6214 36254 6260 36306
rect 6260 36254 6266 36306
rect 6148 36184 6154 36236
rect 6154 36184 6200 36236
rect 6214 36184 6260 36236
rect 6260 36184 6266 36236
rect 6148 36114 6154 36166
rect 6154 36114 6200 36166
rect 6214 36114 6260 36166
rect 6260 36114 6266 36166
rect 6425 35930 6431 35982
rect 6431 35930 6477 35982
rect 6491 35930 6537 35982
rect 6537 35930 6543 35982
rect 6425 35861 6431 35913
rect 6431 35861 6477 35913
rect 6491 35861 6537 35913
rect 6537 35861 6543 35913
rect 6425 35792 6431 35844
rect 6431 35792 6477 35844
rect 6491 35792 6537 35844
rect 6537 35792 6543 35844
rect 6425 35723 6431 35775
rect 6431 35723 6477 35775
rect 6491 35723 6537 35775
rect 6537 35723 6543 35775
rect 6425 35654 6431 35706
rect 6431 35654 6477 35706
rect 6491 35654 6537 35706
rect 6537 35654 6543 35706
rect 6425 35584 6431 35636
rect 6431 35584 6477 35636
rect 6491 35584 6537 35636
rect 6537 35584 6543 35636
rect 6425 35514 6431 35566
rect 6431 35514 6477 35566
rect 6491 35514 6537 35566
rect 6537 35514 6543 35566
rect 6425 35444 6431 35496
rect 6431 35444 6477 35496
rect 6491 35444 6537 35496
rect 6537 35444 6543 35496
rect 6425 35380 6431 35426
rect 6431 35380 6477 35426
rect 6491 35380 6537 35426
rect 6537 35380 6543 35426
rect 6425 35374 6477 35380
rect 6491 35374 6543 35380
rect 6702 36714 6754 36720
rect 6702 36680 6708 36714
rect 6708 36680 6742 36714
rect 6742 36680 6754 36714
rect 6702 36668 6754 36680
rect 6768 36714 6820 36720
rect 6768 36680 6780 36714
rect 6780 36680 6814 36714
rect 6814 36680 6820 36714
rect 6768 36668 6820 36680
rect 6702 36641 6754 36651
rect 6702 36607 6708 36641
rect 6708 36607 6742 36641
rect 6742 36607 6754 36641
rect 6702 36599 6754 36607
rect 6768 36641 6820 36651
rect 6768 36607 6780 36641
rect 6780 36607 6814 36641
rect 6814 36607 6820 36641
rect 6768 36599 6820 36607
rect 6702 36568 6754 36582
rect 6702 36534 6708 36568
rect 6708 36534 6742 36568
rect 6742 36534 6754 36568
rect 6702 36530 6754 36534
rect 6768 36568 6820 36582
rect 6768 36534 6780 36568
rect 6780 36534 6814 36568
rect 6814 36534 6820 36568
rect 6768 36530 6820 36534
rect 6702 36495 6754 36513
rect 6702 36461 6708 36495
rect 6708 36461 6742 36495
rect 6742 36461 6754 36495
rect 6768 36495 6820 36513
rect 6768 36461 6780 36495
rect 6780 36461 6814 36495
rect 6814 36461 6820 36495
rect 6702 36422 6754 36444
rect 6768 36422 6820 36444
rect 6702 36392 6708 36422
rect 6708 36392 6754 36422
rect 6768 36392 6814 36422
rect 6814 36392 6820 36422
rect 6702 36323 6708 36375
rect 6708 36323 6754 36375
rect 6768 36323 6814 36375
rect 6814 36323 6820 36375
rect 6702 36254 6708 36306
rect 6708 36254 6754 36306
rect 6768 36254 6814 36306
rect 6814 36254 6820 36306
rect 6702 36184 6708 36236
rect 6708 36184 6754 36236
rect 6768 36184 6814 36236
rect 6814 36184 6820 36236
rect 6702 36114 6708 36166
rect 6708 36114 6754 36166
rect 6768 36114 6814 36166
rect 6814 36114 6820 36166
rect 6979 35930 6985 35982
rect 6985 35930 7031 35982
rect 7045 35930 7091 35982
rect 7091 35930 7097 35982
rect 6979 35861 6985 35913
rect 6985 35861 7031 35913
rect 7045 35861 7091 35913
rect 7091 35861 7097 35913
rect 6979 35792 6985 35844
rect 6985 35792 7031 35844
rect 7045 35792 7091 35844
rect 7091 35792 7097 35844
rect 6979 35723 6985 35775
rect 6985 35723 7031 35775
rect 7045 35723 7091 35775
rect 7091 35723 7097 35775
rect 6979 35654 6985 35706
rect 6985 35654 7031 35706
rect 7045 35654 7091 35706
rect 7091 35654 7097 35706
rect 6979 35584 6985 35636
rect 6985 35584 7031 35636
rect 7045 35584 7091 35636
rect 7091 35584 7097 35636
rect 6979 35514 6985 35566
rect 6985 35514 7031 35566
rect 7045 35514 7091 35566
rect 7091 35514 7097 35566
rect 6979 35444 6985 35496
rect 6985 35444 7031 35496
rect 7045 35444 7091 35496
rect 7091 35444 7097 35496
rect 6979 35380 6985 35426
rect 6985 35380 7031 35426
rect 7045 35380 7091 35426
rect 7091 35380 7097 35426
rect 6979 35374 7031 35380
rect 7045 35374 7097 35380
rect 7256 36714 7308 36720
rect 7256 36680 7262 36714
rect 7262 36680 7296 36714
rect 7296 36680 7308 36714
rect 7256 36668 7308 36680
rect 7322 36714 7374 36720
rect 7322 36680 7334 36714
rect 7334 36680 7368 36714
rect 7368 36680 7374 36714
rect 7322 36668 7374 36680
rect 7256 36641 7308 36651
rect 7256 36607 7262 36641
rect 7262 36607 7296 36641
rect 7296 36607 7308 36641
rect 7256 36599 7308 36607
rect 7322 36641 7374 36651
rect 7322 36607 7334 36641
rect 7334 36607 7368 36641
rect 7368 36607 7374 36641
rect 7322 36599 7374 36607
rect 7256 36568 7308 36582
rect 7256 36534 7262 36568
rect 7262 36534 7296 36568
rect 7296 36534 7308 36568
rect 7256 36530 7308 36534
rect 7322 36568 7374 36582
rect 7322 36534 7334 36568
rect 7334 36534 7368 36568
rect 7368 36534 7374 36568
rect 7322 36530 7374 36534
rect 7256 36495 7308 36513
rect 7256 36461 7262 36495
rect 7262 36461 7296 36495
rect 7296 36461 7308 36495
rect 7322 36495 7374 36513
rect 7322 36461 7334 36495
rect 7334 36461 7368 36495
rect 7368 36461 7374 36495
rect 7256 36422 7308 36444
rect 7322 36422 7374 36444
rect 7256 36392 7262 36422
rect 7262 36392 7308 36422
rect 7322 36392 7368 36422
rect 7368 36392 7374 36422
rect 7256 36323 7262 36375
rect 7262 36323 7308 36375
rect 7322 36323 7368 36375
rect 7368 36323 7374 36375
rect 7256 36254 7262 36306
rect 7262 36254 7308 36306
rect 7322 36254 7368 36306
rect 7368 36254 7374 36306
rect 7256 36184 7262 36236
rect 7262 36184 7308 36236
rect 7322 36184 7368 36236
rect 7368 36184 7374 36236
rect 7256 36114 7262 36166
rect 7262 36114 7308 36166
rect 7322 36114 7368 36166
rect 7368 36114 7374 36166
rect 7533 35930 7539 35982
rect 7539 35930 7585 35982
rect 7599 35930 7645 35982
rect 7645 35930 7651 35982
rect 7533 35861 7539 35913
rect 7539 35861 7585 35913
rect 7599 35861 7645 35913
rect 7645 35861 7651 35913
rect 7533 35792 7539 35844
rect 7539 35792 7585 35844
rect 7599 35792 7645 35844
rect 7645 35792 7651 35844
rect 7533 35723 7539 35775
rect 7539 35723 7585 35775
rect 7599 35723 7645 35775
rect 7645 35723 7651 35775
rect 7533 35654 7539 35706
rect 7539 35654 7585 35706
rect 7599 35654 7645 35706
rect 7645 35654 7651 35706
rect 7533 35584 7539 35636
rect 7539 35584 7585 35636
rect 7599 35584 7645 35636
rect 7645 35584 7651 35636
rect 7533 35514 7539 35566
rect 7539 35514 7585 35566
rect 7599 35514 7645 35566
rect 7645 35514 7651 35566
rect 7533 35444 7539 35496
rect 7539 35444 7585 35496
rect 7599 35444 7645 35496
rect 7645 35444 7651 35496
rect 7533 35380 7539 35426
rect 7539 35380 7585 35426
rect 7599 35380 7645 35426
rect 7645 35380 7651 35426
rect 7533 35374 7585 35380
rect 7599 35374 7651 35380
rect 7810 36714 7862 36720
rect 7810 36680 7816 36714
rect 7816 36680 7850 36714
rect 7850 36680 7862 36714
rect 7810 36668 7862 36680
rect 7876 36714 7928 36720
rect 7876 36680 7888 36714
rect 7888 36680 7922 36714
rect 7922 36680 7928 36714
rect 7876 36668 7928 36680
rect 7810 36641 7862 36651
rect 7810 36607 7816 36641
rect 7816 36607 7850 36641
rect 7850 36607 7862 36641
rect 7810 36599 7862 36607
rect 7876 36641 7928 36651
rect 7876 36607 7888 36641
rect 7888 36607 7922 36641
rect 7922 36607 7928 36641
rect 7876 36599 7928 36607
rect 7810 36568 7862 36582
rect 7810 36534 7816 36568
rect 7816 36534 7850 36568
rect 7850 36534 7862 36568
rect 7810 36530 7862 36534
rect 7876 36568 7928 36582
rect 7876 36534 7888 36568
rect 7888 36534 7922 36568
rect 7922 36534 7928 36568
rect 7876 36530 7928 36534
rect 7810 36495 7862 36513
rect 7810 36461 7816 36495
rect 7816 36461 7850 36495
rect 7850 36461 7862 36495
rect 7876 36495 7928 36513
rect 7876 36461 7888 36495
rect 7888 36461 7922 36495
rect 7922 36461 7928 36495
rect 7810 36422 7862 36444
rect 7876 36422 7928 36444
rect 7810 36392 7816 36422
rect 7816 36392 7862 36422
rect 7876 36392 7922 36422
rect 7922 36392 7928 36422
rect 7810 36323 7816 36375
rect 7816 36323 7862 36375
rect 7876 36323 7922 36375
rect 7922 36323 7928 36375
rect 7810 36254 7816 36306
rect 7816 36254 7862 36306
rect 7876 36254 7922 36306
rect 7922 36254 7928 36306
rect 7810 36184 7816 36236
rect 7816 36184 7862 36236
rect 7876 36184 7922 36236
rect 7922 36184 7928 36236
rect 7810 36114 7816 36166
rect 7816 36114 7862 36166
rect 7876 36114 7922 36166
rect 7922 36114 7928 36166
rect 8047 36703 8099 36724
rect 8047 36672 8050 36703
rect 8050 36672 8084 36703
rect 8084 36672 8099 36703
rect 8169 36693 8221 36724
rect 8169 36672 8184 36693
rect 8184 36672 8218 36693
rect 8218 36672 8221 36693
rect 8047 36631 8099 36655
rect 8047 36603 8050 36631
rect 8050 36603 8084 36631
rect 8084 36603 8099 36631
rect 8169 36621 8221 36655
rect 8169 36603 8184 36621
rect 8184 36603 8218 36621
rect 8218 36603 8221 36621
rect 8047 36559 8099 36586
rect 8047 36534 8050 36559
rect 8050 36534 8084 36559
rect 8084 36534 8099 36559
rect 8169 36549 8221 36586
rect 8169 36534 8184 36549
rect 8184 36534 8218 36549
rect 8218 36534 8221 36549
rect 8047 36487 8099 36517
rect 8047 36465 8050 36487
rect 8050 36465 8084 36487
rect 8084 36465 8099 36487
rect 8169 36515 8184 36517
rect 8184 36515 8218 36517
rect 8218 36515 8221 36517
rect 8169 36477 8221 36515
rect 8169 36465 8184 36477
rect 8184 36465 8218 36477
rect 8218 36465 8221 36477
rect 8047 36415 8099 36448
rect 8047 36396 8050 36415
rect 8050 36396 8084 36415
rect 8084 36396 8099 36415
rect 8169 36443 8184 36448
rect 8184 36443 8218 36448
rect 8218 36443 8221 36448
rect 8169 36405 8221 36443
rect 8169 36396 8184 36405
rect 8184 36396 8218 36405
rect 8218 36396 8221 36405
rect 8047 36343 8099 36378
rect 8047 36326 8050 36343
rect 8050 36326 8084 36343
rect 8084 36326 8099 36343
rect 8169 36371 8184 36378
rect 8184 36371 8218 36378
rect 8218 36371 8221 36378
rect 8169 36333 8221 36371
rect 8169 36326 8184 36333
rect 8184 36326 8218 36333
rect 8218 36326 8221 36333
rect 8047 36271 8099 36308
rect 8047 36256 8050 36271
rect 8050 36256 8084 36271
rect 8084 36256 8099 36271
rect 8169 36299 8184 36308
rect 8184 36299 8218 36308
rect 8218 36299 8221 36308
rect 8169 36261 8221 36299
rect 8169 36256 8184 36261
rect 8184 36256 8218 36261
rect 8218 36256 8221 36261
rect 8047 36237 8050 36238
rect 8050 36237 8084 36238
rect 8084 36237 8099 36238
rect 8047 36199 8099 36237
rect 8047 36186 8050 36199
rect 8050 36186 8084 36199
rect 8084 36186 8099 36199
rect 8169 36227 8184 36238
rect 8184 36227 8218 36238
rect 8218 36227 8221 36238
rect 8169 36189 8221 36227
rect 8169 36186 8184 36189
rect 8184 36186 8218 36189
rect 8218 36186 8221 36189
rect 8047 36165 8050 36168
rect 8050 36165 8084 36168
rect 8084 36165 8099 36168
rect 8047 36127 8099 36165
rect 8047 36116 8050 36127
rect 8050 36116 8084 36127
rect 8084 36116 8099 36127
rect 8169 36155 8184 36168
rect 8184 36155 8218 36168
rect 8218 36155 8221 36168
rect 8169 36117 8221 36155
rect 8169 36116 8184 36117
rect 8184 36116 8218 36117
rect 8218 36116 8221 36117
rect 2824 34714 2876 34720
rect 2824 34680 2830 34714
rect 2830 34680 2864 34714
rect 2864 34680 2876 34714
rect 2824 34668 2876 34680
rect 2890 34714 2942 34720
rect 2890 34680 2902 34714
rect 2902 34680 2936 34714
rect 2936 34680 2942 34714
rect 2890 34668 2942 34680
rect 2824 34641 2876 34651
rect 2824 34607 2830 34641
rect 2830 34607 2864 34641
rect 2864 34607 2876 34641
rect 2824 34599 2876 34607
rect 2890 34641 2942 34651
rect 2890 34607 2902 34641
rect 2902 34607 2936 34641
rect 2936 34607 2942 34641
rect 2890 34599 2942 34607
rect 2824 34568 2876 34582
rect 2824 34534 2830 34568
rect 2830 34534 2864 34568
rect 2864 34534 2876 34568
rect 2824 34530 2876 34534
rect 2890 34568 2942 34582
rect 2890 34534 2902 34568
rect 2902 34534 2936 34568
rect 2936 34534 2942 34568
rect 2890 34530 2942 34534
rect 2824 34495 2876 34513
rect 2824 34461 2830 34495
rect 2830 34461 2864 34495
rect 2864 34461 2876 34495
rect 2890 34495 2942 34513
rect 2890 34461 2902 34495
rect 2902 34461 2936 34495
rect 2936 34461 2942 34495
rect 2824 34422 2876 34444
rect 2890 34422 2942 34444
rect 2824 34392 2830 34422
rect 2830 34392 2876 34422
rect 2890 34392 2936 34422
rect 2936 34392 2942 34422
rect 2824 34323 2830 34375
rect 2830 34323 2876 34375
rect 2890 34323 2936 34375
rect 2936 34323 2942 34375
rect 2824 34254 2830 34306
rect 2830 34254 2876 34306
rect 2890 34254 2936 34306
rect 2936 34254 2942 34306
rect 2824 34184 2830 34236
rect 2830 34184 2876 34236
rect 2890 34184 2936 34236
rect 2936 34184 2942 34236
rect 2824 34114 2830 34166
rect 2830 34114 2876 34166
rect 2890 34114 2936 34166
rect 2936 34114 2942 34166
rect 3101 33930 3107 33982
rect 3107 33930 3153 33982
rect 3167 33930 3213 33982
rect 3213 33930 3219 33982
rect 3101 33861 3107 33913
rect 3107 33861 3153 33913
rect 3167 33861 3213 33913
rect 3213 33861 3219 33913
rect 3101 33792 3107 33844
rect 3107 33792 3153 33844
rect 3167 33792 3213 33844
rect 3213 33792 3219 33844
rect 3101 33723 3107 33775
rect 3107 33723 3153 33775
rect 3167 33723 3213 33775
rect 3213 33723 3219 33775
rect 3101 33654 3107 33706
rect 3107 33654 3153 33706
rect 3167 33654 3213 33706
rect 3213 33654 3219 33706
rect 3101 33584 3107 33636
rect 3107 33584 3153 33636
rect 3167 33584 3213 33636
rect 3213 33584 3219 33636
rect 3101 33514 3107 33566
rect 3107 33514 3153 33566
rect 3167 33514 3213 33566
rect 3213 33514 3219 33566
rect 3101 33444 3107 33496
rect 3107 33444 3153 33496
rect 3167 33444 3213 33496
rect 3213 33444 3219 33496
rect 3101 33380 3107 33426
rect 3107 33380 3153 33426
rect 3167 33380 3213 33426
rect 3213 33380 3219 33426
rect 3101 33374 3153 33380
rect 3167 33374 3219 33380
rect 3378 34714 3430 34720
rect 3378 34680 3384 34714
rect 3384 34680 3418 34714
rect 3418 34680 3430 34714
rect 3378 34668 3430 34680
rect 3444 34714 3496 34720
rect 3444 34680 3456 34714
rect 3456 34680 3490 34714
rect 3490 34680 3496 34714
rect 3444 34668 3496 34680
rect 3378 34641 3430 34651
rect 3378 34607 3384 34641
rect 3384 34607 3418 34641
rect 3418 34607 3430 34641
rect 3378 34599 3430 34607
rect 3444 34641 3496 34651
rect 3444 34607 3456 34641
rect 3456 34607 3490 34641
rect 3490 34607 3496 34641
rect 3444 34599 3496 34607
rect 3378 34568 3430 34582
rect 3378 34534 3384 34568
rect 3384 34534 3418 34568
rect 3418 34534 3430 34568
rect 3378 34530 3430 34534
rect 3444 34568 3496 34582
rect 3444 34534 3456 34568
rect 3456 34534 3490 34568
rect 3490 34534 3496 34568
rect 3444 34530 3496 34534
rect 3378 34495 3430 34513
rect 3378 34461 3384 34495
rect 3384 34461 3418 34495
rect 3418 34461 3430 34495
rect 3444 34495 3496 34513
rect 3444 34461 3456 34495
rect 3456 34461 3490 34495
rect 3490 34461 3496 34495
rect 3378 34422 3430 34444
rect 3444 34422 3496 34444
rect 3378 34392 3384 34422
rect 3384 34392 3430 34422
rect 3444 34392 3490 34422
rect 3490 34392 3496 34422
rect 3378 34323 3384 34375
rect 3384 34323 3430 34375
rect 3444 34323 3490 34375
rect 3490 34323 3496 34375
rect 3378 34254 3384 34306
rect 3384 34254 3430 34306
rect 3444 34254 3490 34306
rect 3490 34254 3496 34306
rect 3378 34184 3384 34236
rect 3384 34184 3430 34236
rect 3444 34184 3490 34236
rect 3490 34184 3496 34236
rect 3378 34114 3384 34166
rect 3384 34114 3430 34166
rect 3444 34114 3490 34166
rect 3490 34114 3496 34166
rect 3655 33930 3661 33982
rect 3661 33930 3707 33982
rect 3721 33930 3767 33982
rect 3767 33930 3773 33982
rect 3655 33861 3661 33913
rect 3661 33861 3707 33913
rect 3721 33861 3767 33913
rect 3767 33861 3773 33913
rect 3655 33792 3661 33844
rect 3661 33792 3707 33844
rect 3721 33792 3767 33844
rect 3767 33792 3773 33844
rect 3655 33723 3661 33775
rect 3661 33723 3707 33775
rect 3721 33723 3767 33775
rect 3767 33723 3773 33775
rect 3655 33654 3661 33706
rect 3661 33654 3707 33706
rect 3721 33654 3767 33706
rect 3767 33654 3773 33706
rect 3655 33584 3661 33636
rect 3661 33584 3707 33636
rect 3721 33584 3767 33636
rect 3767 33584 3773 33636
rect 3655 33514 3661 33566
rect 3661 33514 3707 33566
rect 3721 33514 3767 33566
rect 3767 33514 3773 33566
rect 3655 33444 3661 33496
rect 3661 33444 3707 33496
rect 3721 33444 3767 33496
rect 3767 33444 3773 33496
rect 3655 33380 3661 33426
rect 3661 33380 3707 33426
rect 3721 33380 3767 33426
rect 3767 33380 3773 33426
rect 3655 33374 3707 33380
rect 3721 33374 3773 33380
rect 3932 34714 3984 34720
rect 3932 34680 3938 34714
rect 3938 34680 3972 34714
rect 3972 34680 3984 34714
rect 3932 34668 3984 34680
rect 3998 34714 4050 34720
rect 3998 34680 4010 34714
rect 4010 34680 4044 34714
rect 4044 34680 4050 34714
rect 3998 34668 4050 34680
rect 3932 34641 3984 34651
rect 3932 34607 3938 34641
rect 3938 34607 3972 34641
rect 3972 34607 3984 34641
rect 3932 34599 3984 34607
rect 3998 34641 4050 34651
rect 3998 34607 4010 34641
rect 4010 34607 4044 34641
rect 4044 34607 4050 34641
rect 3998 34599 4050 34607
rect 3932 34568 3984 34582
rect 3932 34534 3938 34568
rect 3938 34534 3972 34568
rect 3972 34534 3984 34568
rect 3932 34530 3984 34534
rect 3998 34568 4050 34582
rect 3998 34534 4010 34568
rect 4010 34534 4044 34568
rect 4044 34534 4050 34568
rect 3998 34530 4050 34534
rect 3932 34495 3984 34513
rect 3932 34461 3938 34495
rect 3938 34461 3972 34495
rect 3972 34461 3984 34495
rect 3998 34495 4050 34513
rect 3998 34461 4010 34495
rect 4010 34461 4044 34495
rect 4044 34461 4050 34495
rect 3932 34422 3984 34444
rect 3998 34422 4050 34444
rect 3932 34392 3938 34422
rect 3938 34392 3984 34422
rect 3998 34392 4044 34422
rect 4044 34392 4050 34422
rect 3932 34323 3938 34375
rect 3938 34323 3984 34375
rect 3998 34323 4044 34375
rect 4044 34323 4050 34375
rect 3932 34254 3938 34306
rect 3938 34254 3984 34306
rect 3998 34254 4044 34306
rect 4044 34254 4050 34306
rect 3932 34184 3938 34236
rect 3938 34184 3984 34236
rect 3998 34184 4044 34236
rect 4044 34184 4050 34236
rect 3932 34114 3938 34166
rect 3938 34114 3984 34166
rect 3998 34114 4044 34166
rect 4044 34114 4050 34166
rect 4209 33930 4215 33982
rect 4215 33930 4261 33982
rect 4275 33930 4321 33982
rect 4321 33930 4327 33982
rect 4209 33861 4215 33913
rect 4215 33861 4261 33913
rect 4275 33861 4321 33913
rect 4321 33861 4327 33913
rect 4209 33792 4215 33844
rect 4215 33792 4261 33844
rect 4275 33792 4321 33844
rect 4321 33792 4327 33844
rect 4209 33723 4215 33775
rect 4215 33723 4261 33775
rect 4275 33723 4321 33775
rect 4321 33723 4327 33775
rect 4209 33654 4215 33706
rect 4215 33654 4261 33706
rect 4275 33654 4321 33706
rect 4321 33654 4327 33706
rect 4209 33584 4215 33636
rect 4215 33584 4261 33636
rect 4275 33584 4321 33636
rect 4321 33584 4327 33636
rect 4209 33514 4215 33566
rect 4215 33514 4261 33566
rect 4275 33514 4321 33566
rect 4321 33514 4327 33566
rect 4209 33444 4215 33496
rect 4215 33444 4261 33496
rect 4275 33444 4321 33496
rect 4321 33444 4327 33496
rect 4209 33380 4215 33426
rect 4215 33380 4261 33426
rect 4275 33380 4321 33426
rect 4321 33380 4327 33426
rect 4209 33374 4261 33380
rect 4275 33374 4327 33380
rect 4486 34714 4538 34720
rect 4486 34680 4492 34714
rect 4492 34680 4526 34714
rect 4526 34680 4538 34714
rect 4486 34668 4538 34680
rect 4552 34714 4604 34720
rect 4552 34680 4564 34714
rect 4564 34680 4598 34714
rect 4598 34680 4604 34714
rect 4552 34668 4604 34680
rect 4486 34641 4538 34651
rect 4486 34607 4492 34641
rect 4492 34607 4526 34641
rect 4526 34607 4538 34641
rect 4486 34599 4538 34607
rect 4552 34641 4604 34651
rect 4552 34607 4564 34641
rect 4564 34607 4598 34641
rect 4598 34607 4604 34641
rect 4552 34599 4604 34607
rect 4486 34568 4538 34582
rect 4486 34534 4492 34568
rect 4492 34534 4526 34568
rect 4526 34534 4538 34568
rect 4486 34530 4538 34534
rect 4552 34568 4604 34582
rect 4552 34534 4564 34568
rect 4564 34534 4598 34568
rect 4598 34534 4604 34568
rect 4552 34530 4604 34534
rect 4486 34495 4538 34513
rect 4486 34461 4492 34495
rect 4492 34461 4526 34495
rect 4526 34461 4538 34495
rect 4552 34495 4604 34513
rect 4552 34461 4564 34495
rect 4564 34461 4598 34495
rect 4598 34461 4604 34495
rect 4486 34422 4538 34444
rect 4552 34422 4604 34444
rect 4486 34392 4492 34422
rect 4492 34392 4538 34422
rect 4552 34392 4598 34422
rect 4598 34392 4604 34422
rect 4486 34323 4492 34375
rect 4492 34323 4538 34375
rect 4552 34323 4598 34375
rect 4598 34323 4604 34375
rect 4486 34254 4492 34306
rect 4492 34254 4538 34306
rect 4552 34254 4598 34306
rect 4598 34254 4604 34306
rect 4486 34184 4492 34236
rect 4492 34184 4538 34236
rect 4552 34184 4598 34236
rect 4598 34184 4604 34236
rect 4486 34114 4492 34166
rect 4492 34114 4538 34166
rect 4552 34114 4598 34166
rect 4598 34114 4604 34166
rect 4763 33930 4769 33982
rect 4769 33930 4815 33982
rect 4829 33930 4875 33982
rect 4875 33930 4881 33982
rect 4763 33861 4769 33913
rect 4769 33861 4815 33913
rect 4829 33861 4875 33913
rect 4875 33861 4881 33913
rect 4763 33792 4769 33844
rect 4769 33792 4815 33844
rect 4829 33792 4875 33844
rect 4875 33792 4881 33844
rect 4763 33723 4769 33775
rect 4769 33723 4815 33775
rect 4829 33723 4875 33775
rect 4875 33723 4881 33775
rect 4763 33654 4769 33706
rect 4769 33654 4815 33706
rect 4829 33654 4875 33706
rect 4875 33654 4881 33706
rect 4763 33584 4769 33636
rect 4769 33584 4815 33636
rect 4829 33584 4875 33636
rect 4875 33584 4881 33636
rect 4763 33514 4769 33566
rect 4769 33514 4815 33566
rect 4829 33514 4875 33566
rect 4875 33514 4881 33566
rect 4763 33444 4769 33496
rect 4769 33444 4815 33496
rect 4829 33444 4875 33496
rect 4875 33444 4881 33496
rect 4763 33380 4769 33426
rect 4769 33380 4815 33426
rect 4829 33380 4875 33426
rect 4875 33380 4881 33426
rect 4763 33374 4815 33380
rect 4829 33374 4881 33380
rect 5040 34714 5092 34720
rect 5040 34680 5046 34714
rect 5046 34680 5080 34714
rect 5080 34680 5092 34714
rect 5040 34668 5092 34680
rect 5106 34714 5158 34720
rect 5106 34680 5118 34714
rect 5118 34680 5152 34714
rect 5152 34680 5158 34714
rect 5106 34668 5158 34680
rect 5040 34641 5092 34651
rect 5040 34607 5046 34641
rect 5046 34607 5080 34641
rect 5080 34607 5092 34641
rect 5040 34599 5092 34607
rect 5106 34641 5158 34651
rect 5106 34607 5118 34641
rect 5118 34607 5152 34641
rect 5152 34607 5158 34641
rect 5106 34599 5158 34607
rect 5040 34568 5092 34582
rect 5040 34534 5046 34568
rect 5046 34534 5080 34568
rect 5080 34534 5092 34568
rect 5040 34530 5092 34534
rect 5106 34568 5158 34582
rect 5106 34534 5118 34568
rect 5118 34534 5152 34568
rect 5152 34534 5158 34568
rect 5106 34530 5158 34534
rect 5040 34495 5092 34513
rect 5040 34461 5046 34495
rect 5046 34461 5080 34495
rect 5080 34461 5092 34495
rect 5106 34495 5158 34513
rect 5106 34461 5118 34495
rect 5118 34461 5152 34495
rect 5152 34461 5158 34495
rect 5040 34422 5092 34444
rect 5106 34422 5158 34444
rect 5040 34392 5046 34422
rect 5046 34392 5092 34422
rect 5106 34392 5152 34422
rect 5152 34392 5158 34422
rect 5040 34323 5046 34375
rect 5046 34323 5092 34375
rect 5106 34323 5152 34375
rect 5152 34323 5158 34375
rect 5040 34254 5046 34306
rect 5046 34254 5092 34306
rect 5106 34254 5152 34306
rect 5152 34254 5158 34306
rect 5040 34184 5046 34236
rect 5046 34184 5092 34236
rect 5106 34184 5152 34236
rect 5152 34184 5158 34236
rect 5040 34114 5046 34166
rect 5046 34114 5092 34166
rect 5106 34114 5152 34166
rect 5152 34114 5158 34166
rect 5317 33930 5323 33982
rect 5323 33930 5369 33982
rect 5383 33930 5429 33982
rect 5429 33930 5435 33982
rect 5317 33861 5323 33913
rect 5323 33861 5369 33913
rect 5383 33861 5429 33913
rect 5429 33861 5435 33913
rect 5317 33792 5323 33844
rect 5323 33792 5369 33844
rect 5383 33792 5429 33844
rect 5429 33792 5435 33844
rect 5317 33723 5323 33775
rect 5323 33723 5369 33775
rect 5383 33723 5429 33775
rect 5429 33723 5435 33775
rect 5317 33654 5323 33706
rect 5323 33654 5369 33706
rect 5383 33654 5429 33706
rect 5429 33654 5435 33706
rect 5317 33584 5323 33636
rect 5323 33584 5369 33636
rect 5383 33584 5429 33636
rect 5429 33584 5435 33636
rect 5317 33514 5323 33566
rect 5323 33514 5369 33566
rect 5383 33514 5429 33566
rect 5429 33514 5435 33566
rect 5317 33444 5323 33496
rect 5323 33444 5369 33496
rect 5383 33444 5429 33496
rect 5429 33444 5435 33496
rect 5317 33380 5323 33426
rect 5323 33380 5369 33426
rect 5383 33380 5429 33426
rect 5429 33380 5435 33426
rect 5317 33374 5369 33380
rect 5383 33374 5435 33380
rect 5594 34714 5646 34720
rect 5594 34680 5600 34714
rect 5600 34680 5634 34714
rect 5634 34680 5646 34714
rect 5594 34668 5646 34680
rect 5660 34714 5712 34720
rect 5660 34680 5672 34714
rect 5672 34680 5706 34714
rect 5706 34680 5712 34714
rect 5660 34668 5712 34680
rect 5594 34641 5646 34651
rect 5594 34607 5600 34641
rect 5600 34607 5634 34641
rect 5634 34607 5646 34641
rect 5594 34599 5646 34607
rect 5660 34641 5712 34651
rect 5660 34607 5672 34641
rect 5672 34607 5706 34641
rect 5706 34607 5712 34641
rect 5660 34599 5712 34607
rect 5594 34568 5646 34582
rect 5594 34534 5600 34568
rect 5600 34534 5634 34568
rect 5634 34534 5646 34568
rect 5594 34530 5646 34534
rect 5660 34568 5712 34582
rect 5660 34534 5672 34568
rect 5672 34534 5706 34568
rect 5706 34534 5712 34568
rect 5660 34530 5712 34534
rect 5594 34495 5646 34513
rect 5594 34461 5600 34495
rect 5600 34461 5634 34495
rect 5634 34461 5646 34495
rect 5660 34495 5712 34513
rect 5660 34461 5672 34495
rect 5672 34461 5706 34495
rect 5706 34461 5712 34495
rect 5594 34422 5646 34444
rect 5660 34422 5712 34444
rect 5594 34392 5600 34422
rect 5600 34392 5646 34422
rect 5660 34392 5706 34422
rect 5706 34392 5712 34422
rect 5594 34323 5600 34375
rect 5600 34323 5646 34375
rect 5660 34323 5706 34375
rect 5706 34323 5712 34375
rect 5594 34254 5600 34306
rect 5600 34254 5646 34306
rect 5660 34254 5706 34306
rect 5706 34254 5712 34306
rect 5594 34184 5600 34236
rect 5600 34184 5646 34236
rect 5660 34184 5706 34236
rect 5706 34184 5712 34236
rect 5594 34114 5600 34166
rect 5600 34114 5646 34166
rect 5660 34114 5706 34166
rect 5706 34114 5712 34166
rect 5871 33930 5877 33982
rect 5877 33930 5923 33982
rect 5937 33930 5983 33982
rect 5983 33930 5989 33982
rect 5871 33861 5877 33913
rect 5877 33861 5923 33913
rect 5937 33861 5983 33913
rect 5983 33861 5989 33913
rect 5871 33792 5877 33844
rect 5877 33792 5923 33844
rect 5937 33792 5983 33844
rect 5983 33792 5989 33844
rect 5871 33723 5877 33775
rect 5877 33723 5923 33775
rect 5937 33723 5983 33775
rect 5983 33723 5989 33775
rect 5871 33654 5877 33706
rect 5877 33654 5923 33706
rect 5937 33654 5983 33706
rect 5983 33654 5989 33706
rect 5871 33584 5877 33636
rect 5877 33584 5923 33636
rect 5937 33584 5983 33636
rect 5983 33584 5989 33636
rect 5871 33514 5877 33566
rect 5877 33514 5923 33566
rect 5937 33514 5983 33566
rect 5983 33514 5989 33566
rect 5871 33444 5877 33496
rect 5877 33444 5923 33496
rect 5937 33444 5983 33496
rect 5983 33444 5989 33496
rect 5871 33380 5877 33426
rect 5877 33380 5923 33426
rect 5937 33380 5983 33426
rect 5983 33380 5989 33426
rect 5871 33374 5923 33380
rect 5937 33374 5989 33380
rect 6148 34714 6200 34720
rect 6148 34680 6154 34714
rect 6154 34680 6188 34714
rect 6188 34680 6200 34714
rect 6148 34668 6200 34680
rect 6214 34714 6266 34720
rect 6214 34680 6226 34714
rect 6226 34680 6260 34714
rect 6260 34680 6266 34714
rect 6214 34668 6266 34680
rect 6148 34641 6200 34651
rect 6148 34607 6154 34641
rect 6154 34607 6188 34641
rect 6188 34607 6200 34641
rect 6148 34599 6200 34607
rect 6214 34641 6266 34651
rect 6214 34607 6226 34641
rect 6226 34607 6260 34641
rect 6260 34607 6266 34641
rect 6214 34599 6266 34607
rect 6148 34568 6200 34582
rect 6148 34534 6154 34568
rect 6154 34534 6188 34568
rect 6188 34534 6200 34568
rect 6148 34530 6200 34534
rect 6214 34568 6266 34582
rect 6214 34534 6226 34568
rect 6226 34534 6260 34568
rect 6260 34534 6266 34568
rect 6214 34530 6266 34534
rect 6148 34495 6200 34513
rect 6148 34461 6154 34495
rect 6154 34461 6188 34495
rect 6188 34461 6200 34495
rect 6214 34495 6266 34513
rect 6214 34461 6226 34495
rect 6226 34461 6260 34495
rect 6260 34461 6266 34495
rect 6148 34422 6200 34444
rect 6214 34422 6266 34444
rect 6148 34392 6154 34422
rect 6154 34392 6200 34422
rect 6214 34392 6260 34422
rect 6260 34392 6266 34422
rect 6148 34323 6154 34375
rect 6154 34323 6200 34375
rect 6214 34323 6260 34375
rect 6260 34323 6266 34375
rect 6148 34254 6154 34306
rect 6154 34254 6200 34306
rect 6214 34254 6260 34306
rect 6260 34254 6266 34306
rect 6148 34184 6154 34236
rect 6154 34184 6200 34236
rect 6214 34184 6260 34236
rect 6260 34184 6266 34236
rect 6148 34114 6154 34166
rect 6154 34114 6200 34166
rect 6214 34114 6260 34166
rect 6260 34114 6266 34166
rect 6425 33930 6431 33982
rect 6431 33930 6477 33982
rect 6491 33930 6537 33982
rect 6537 33930 6543 33982
rect 6425 33861 6431 33913
rect 6431 33861 6477 33913
rect 6491 33861 6537 33913
rect 6537 33861 6543 33913
rect 6425 33792 6431 33844
rect 6431 33792 6477 33844
rect 6491 33792 6537 33844
rect 6537 33792 6543 33844
rect 6425 33723 6431 33775
rect 6431 33723 6477 33775
rect 6491 33723 6537 33775
rect 6537 33723 6543 33775
rect 6425 33654 6431 33706
rect 6431 33654 6477 33706
rect 6491 33654 6537 33706
rect 6537 33654 6543 33706
rect 6425 33584 6431 33636
rect 6431 33584 6477 33636
rect 6491 33584 6537 33636
rect 6537 33584 6543 33636
rect 6425 33514 6431 33566
rect 6431 33514 6477 33566
rect 6491 33514 6537 33566
rect 6537 33514 6543 33566
rect 6425 33444 6431 33496
rect 6431 33444 6477 33496
rect 6491 33444 6537 33496
rect 6537 33444 6543 33496
rect 6425 33380 6431 33426
rect 6431 33380 6477 33426
rect 6491 33380 6537 33426
rect 6537 33380 6543 33426
rect 6425 33374 6477 33380
rect 6491 33374 6543 33380
rect 6702 34714 6754 34720
rect 6702 34680 6708 34714
rect 6708 34680 6742 34714
rect 6742 34680 6754 34714
rect 6702 34668 6754 34680
rect 6768 34714 6820 34720
rect 6768 34680 6780 34714
rect 6780 34680 6814 34714
rect 6814 34680 6820 34714
rect 6768 34668 6820 34680
rect 6702 34641 6754 34651
rect 6702 34607 6708 34641
rect 6708 34607 6742 34641
rect 6742 34607 6754 34641
rect 6702 34599 6754 34607
rect 6768 34641 6820 34651
rect 6768 34607 6780 34641
rect 6780 34607 6814 34641
rect 6814 34607 6820 34641
rect 6768 34599 6820 34607
rect 6702 34568 6754 34582
rect 6702 34534 6708 34568
rect 6708 34534 6742 34568
rect 6742 34534 6754 34568
rect 6702 34530 6754 34534
rect 6768 34568 6820 34582
rect 6768 34534 6780 34568
rect 6780 34534 6814 34568
rect 6814 34534 6820 34568
rect 6768 34530 6820 34534
rect 6702 34495 6754 34513
rect 6702 34461 6708 34495
rect 6708 34461 6742 34495
rect 6742 34461 6754 34495
rect 6768 34495 6820 34513
rect 6768 34461 6780 34495
rect 6780 34461 6814 34495
rect 6814 34461 6820 34495
rect 6702 34422 6754 34444
rect 6768 34422 6820 34444
rect 6702 34392 6708 34422
rect 6708 34392 6754 34422
rect 6768 34392 6814 34422
rect 6814 34392 6820 34422
rect 6702 34323 6708 34375
rect 6708 34323 6754 34375
rect 6768 34323 6814 34375
rect 6814 34323 6820 34375
rect 6702 34254 6708 34306
rect 6708 34254 6754 34306
rect 6768 34254 6814 34306
rect 6814 34254 6820 34306
rect 6702 34184 6708 34236
rect 6708 34184 6754 34236
rect 6768 34184 6814 34236
rect 6814 34184 6820 34236
rect 6702 34114 6708 34166
rect 6708 34114 6754 34166
rect 6768 34114 6814 34166
rect 6814 34114 6820 34166
rect 6979 33930 6985 33982
rect 6985 33930 7031 33982
rect 7045 33930 7091 33982
rect 7091 33930 7097 33982
rect 6979 33861 6985 33913
rect 6985 33861 7031 33913
rect 7045 33861 7091 33913
rect 7091 33861 7097 33913
rect 6979 33792 6985 33844
rect 6985 33792 7031 33844
rect 7045 33792 7091 33844
rect 7091 33792 7097 33844
rect 6979 33723 6985 33775
rect 6985 33723 7031 33775
rect 7045 33723 7091 33775
rect 7091 33723 7097 33775
rect 6979 33654 6985 33706
rect 6985 33654 7031 33706
rect 7045 33654 7091 33706
rect 7091 33654 7097 33706
rect 6979 33584 6985 33636
rect 6985 33584 7031 33636
rect 7045 33584 7091 33636
rect 7091 33584 7097 33636
rect 6979 33514 6985 33566
rect 6985 33514 7031 33566
rect 7045 33514 7091 33566
rect 7091 33514 7097 33566
rect 6979 33444 6985 33496
rect 6985 33444 7031 33496
rect 7045 33444 7091 33496
rect 7091 33444 7097 33496
rect 6979 33380 6985 33426
rect 6985 33380 7031 33426
rect 7045 33380 7091 33426
rect 7091 33380 7097 33426
rect 6979 33374 7031 33380
rect 7045 33374 7097 33380
rect 7256 34714 7308 34720
rect 7256 34680 7262 34714
rect 7262 34680 7296 34714
rect 7296 34680 7308 34714
rect 7256 34668 7308 34680
rect 7322 34714 7374 34720
rect 7322 34680 7334 34714
rect 7334 34680 7368 34714
rect 7368 34680 7374 34714
rect 7322 34668 7374 34680
rect 7256 34641 7308 34651
rect 7256 34607 7262 34641
rect 7262 34607 7296 34641
rect 7296 34607 7308 34641
rect 7256 34599 7308 34607
rect 7322 34641 7374 34651
rect 7322 34607 7334 34641
rect 7334 34607 7368 34641
rect 7368 34607 7374 34641
rect 7322 34599 7374 34607
rect 7256 34568 7308 34582
rect 7256 34534 7262 34568
rect 7262 34534 7296 34568
rect 7296 34534 7308 34568
rect 7256 34530 7308 34534
rect 7322 34568 7374 34582
rect 7322 34534 7334 34568
rect 7334 34534 7368 34568
rect 7368 34534 7374 34568
rect 7322 34530 7374 34534
rect 7256 34495 7308 34513
rect 7256 34461 7262 34495
rect 7262 34461 7296 34495
rect 7296 34461 7308 34495
rect 7322 34495 7374 34513
rect 7322 34461 7334 34495
rect 7334 34461 7368 34495
rect 7368 34461 7374 34495
rect 7256 34422 7308 34444
rect 7322 34422 7374 34444
rect 7256 34392 7262 34422
rect 7262 34392 7308 34422
rect 7322 34392 7368 34422
rect 7368 34392 7374 34422
rect 7256 34323 7262 34375
rect 7262 34323 7308 34375
rect 7322 34323 7368 34375
rect 7368 34323 7374 34375
rect 7256 34254 7262 34306
rect 7262 34254 7308 34306
rect 7322 34254 7368 34306
rect 7368 34254 7374 34306
rect 7256 34184 7262 34236
rect 7262 34184 7308 34236
rect 7322 34184 7368 34236
rect 7368 34184 7374 34236
rect 7256 34114 7262 34166
rect 7262 34114 7308 34166
rect 7322 34114 7368 34166
rect 7368 34114 7374 34166
rect 7533 33930 7539 33982
rect 7539 33930 7585 33982
rect 7599 33930 7645 33982
rect 7645 33930 7651 33982
rect 7533 33861 7539 33913
rect 7539 33861 7585 33913
rect 7599 33861 7645 33913
rect 7645 33861 7651 33913
rect 7533 33792 7539 33844
rect 7539 33792 7585 33844
rect 7599 33792 7645 33844
rect 7645 33792 7651 33844
rect 7533 33723 7539 33775
rect 7539 33723 7585 33775
rect 7599 33723 7645 33775
rect 7645 33723 7651 33775
rect 7533 33654 7539 33706
rect 7539 33654 7585 33706
rect 7599 33654 7645 33706
rect 7645 33654 7651 33706
rect 7533 33584 7539 33636
rect 7539 33584 7585 33636
rect 7599 33584 7645 33636
rect 7645 33584 7651 33636
rect 7533 33514 7539 33566
rect 7539 33514 7585 33566
rect 7599 33514 7645 33566
rect 7645 33514 7651 33566
rect 7533 33444 7539 33496
rect 7539 33444 7585 33496
rect 7599 33444 7645 33496
rect 7645 33444 7651 33496
rect 7533 33380 7539 33426
rect 7539 33380 7585 33426
rect 7599 33380 7645 33426
rect 7645 33380 7651 33426
rect 7533 33374 7585 33380
rect 7599 33374 7651 33380
rect 7810 34714 7862 34720
rect 7810 34680 7816 34714
rect 7816 34680 7850 34714
rect 7850 34680 7862 34714
rect 7810 34668 7862 34680
rect 7876 34714 7928 34720
rect 7876 34680 7888 34714
rect 7888 34680 7922 34714
rect 7922 34680 7928 34714
rect 7876 34668 7928 34680
rect 7810 34641 7862 34651
rect 7810 34607 7816 34641
rect 7816 34607 7850 34641
rect 7850 34607 7862 34641
rect 7810 34599 7862 34607
rect 7876 34641 7928 34651
rect 7876 34607 7888 34641
rect 7888 34607 7922 34641
rect 7922 34607 7928 34641
rect 7876 34599 7928 34607
rect 7810 34568 7862 34582
rect 7810 34534 7816 34568
rect 7816 34534 7850 34568
rect 7850 34534 7862 34568
rect 7810 34530 7862 34534
rect 7876 34568 7928 34582
rect 7876 34534 7888 34568
rect 7888 34534 7922 34568
rect 7922 34534 7928 34568
rect 7876 34530 7928 34534
rect 7810 34495 7862 34513
rect 7810 34461 7816 34495
rect 7816 34461 7850 34495
rect 7850 34461 7862 34495
rect 7876 34495 7928 34513
rect 7876 34461 7888 34495
rect 7888 34461 7922 34495
rect 7922 34461 7928 34495
rect 7810 34422 7862 34444
rect 7876 34422 7928 34444
rect 7810 34392 7816 34422
rect 7816 34392 7862 34422
rect 7876 34392 7922 34422
rect 7922 34392 7928 34422
rect 7810 34323 7816 34375
rect 7816 34323 7862 34375
rect 7876 34323 7922 34375
rect 7922 34323 7928 34375
rect 7810 34254 7816 34306
rect 7816 34254 7862 34306
rect 7876 34254 7922 34306
rect 7922 34254 7928 34306
rect 7810 34184 7816 34236
rect 7816 34184 7862 34236
rect 7876 34184 7922 34236
rect 7922 34184 7928 34236
rect 7810 34114 7816 34166
rect 7816 34114 7862 34166
rect 7876 34114 7922 34166
rect 7922 34114 7928 34166
rect 8047 34687 8099 34724
rect 8047 34672 8050 34687
rect 8050 34672 8084 34687
rect 8084 34672 8099 34687
rect 8169 34715 8184 34724
rect 8184 34715 8218 34724
rect 8218 34715 8221 34724
rect 8169 34677 8221 34715
rect 8169 34672 8184 34677
rect 8184 34672 8218 34677
rect 8218 34672 8221 34677
rect 8047 34653 8050 34655
rect 8050 34653 8084 34655
rect 8084 34653 8099 34655
rect 8047 34615 8099 34653
rect 8047 34603 8050 34615
rect 8050 34603 8084 34615
rect 8084 34603 8099 34615
rect 8169 34643 8184 34655
rect 8184 34643 8218 34655
rect 8218 34643 8221 34655
rect 8169 34605 8221 34643
rect 8169 34603 8184 34605
rect 8184 34603 8218 34605
rect 8218 34603 8221 34605
rect 8047 34581 8050 34586
rect 8050 34581 8084 34586
rect 8084 34581 8099 34586
rect 8047 34543 8099 34581
rect 8047 34534 8050 34543
rect 8050 34534 8084 34543
rect 8084 34534 8099 34543
rect 8169 34571 8184 34586
rect 8184 34571 8218 34586
rect 8218 34571 8221 34586
rect 8169 34534 8221 34571
rect 8047 34509 8050 34517
rect 8050 34509 8084 34517
rect 8084 34509 8099 34517
rect 8047 34471 8099 34509
rect 8047 34465 8050 34471
rect 8050 34465 8084 34471
rect 8084 34465 8099 34471
rect 8169 34499 8184 34517
rect 8184 34499 8218 34517
rect 8218 34499 8221 34517
rect 8169 34465 8221 34499
rect 8047 34437 8050 34448
rect 8050 34437 8084 34448
rect 8084 34437 8099 34448
rect 8047 34399 8099 34437
rect 8047 34396 8050 34399
rect 8050 34396 8084 34399
rect 8084 34396 8099 34399
rect 8169 34427 8184 34448
rect 8184 34427 8218 34448
rect 8218 34427 8221 34448
rect 8169 34396 8221 34427
rect 8047 34365 8050 34378
rect 8050 34365 8084 34378
rect 8084 34365 8099 34378
rect 8047 34327 8099 34365
rect 8047 34326 8050 34327
rect 8050 34326 8084 34327
rect 8084 34326 8099 34327
rect 8169 34355 8184 34378
rect 8184 34355 8218 34378
rect 8218 34355 8221 34378
rect 8169 34326 8221 34355
rect 8047 34293 8050 34308
rect 8050 34293 8084 34308
rect 8084 34293 8099 34308
rect 8047 34256 8099 34293
rect 8169 34283 8184 34308
rect 8184 34283 8218 34308
rect 8218 34283 8221 34308
rect 8169 34256 8221 34283
rect 8047 34221 8050 34238
rect 8050 34221 8084 34238
rect 8084 34221 8099 34238
rect 8047 34186 8099 34221
rect 8169 34211 8184 34238
rect 8184 34211 8218 34238
rect 8218 34211 8221 34238
rect 8169 34186 8221 34211
rect 8047 34149 8050 34168
rect 8050 34149 8084 34168
rect 8084 34149 8099 34168
rect 8047 34116 8099 34149
rect 8169 34139 8184 34168
rect 8184 34139 8218 34168
rect 8218 34139 8221 34168
rect 8169 34116 8221 34139
rect 2824 32714 2876 32720
rect 2824 32680 2830 32714
rect 2830 32680 2864 32714
rect 2864 32680 2876 32714
rect 2824 32668 2876 32680
rect 2890 32714 2942 32720
rect 2890 32680 2902 32714
rect 2902 32680 2936 32714
rect 2936 32680 2942 32714
rect 2890 32668 2942 32680
rect 2824 32641 2876 32651
rect 2824 32607 2830 32641
rect 2830 32607 2864 32641
rect 2864 32607 2876 32641
rect 2824 32599 2876 32607
rect 2890 32641 2942 32651
rect 2890 32607 2902 32641
rect 2902 32607 2936 32641
rect 2936 32607 2942 32641
rect 2890 32599 2942 32607
rect 2824 32568 2876 32582
rect 2824 32534 2830 32568
rect 2830 32534 2864 32568
rect 2864 32534 2876 32568
rect 2824 32530 2876 32534
rect 2890 32568 2942 32582
rect 2890 32534 2902 32568
rect 2902 32534 2936 32568
rect 2936 32534 2942 32568
rect 2890 32530 2942 32534
rect 2824 32495 2876 32513
rect 2824 32461 2830 32495
rect 2830 32461 2864 32495
rect 2864 32461 2876 32495
rect 2890 32495 2942 32513
rect 2890 32461 2902 32495
rect 2902 32461 2936 32495
rect 2936 32461 2942 32495
rect 2824 32422 2876 32444
rect 2890 32422 2942 32444
rect 2824 32392 2830 32422
rect 2830 32392 2876 32422
rect 2890 32392 2936 32422
rect 2936 32392 2942 32422
rect 2824 32323 2830 32375
rect 2830 32323 2876 32375
rect 2890 32323 2936 32375
rect 2936 32323 2942 32375
rect 2824 32254 2830 32306
rect 2830 32254 2876 32306
rect 2890 32254 2936 32306
rect 2936 32254 2942 32306
rect 2824 32184 2830 32236
rect 2830 32184 2876 32236
rect 2890 32184 2936 32236
rect 2936 32184 2942 32236
rect 2824 32114 2830 32166
rect 2830 32114 2876 32166
rect 2890 32114 2936 32166
rect 2936 32114 2942 32166
rect 3101 31930 3107 31982
rect 3107 31930 3153 31982
rect 3167 31930 3213 31982
rect 3213 31930 3219 31982
rect 3101 31861 3107 31913
rect 3107 31861 3153 31913
rect 3167 31861 3213 31913
rect 3213 31861 3219 31913
rect 3101 31792 3107 31844
rect 3107 31792 3153 31844
rect 3167 31792 3213 31844
rect 3213 31792 3219 31844
rect 3101 31723 3107 31775
rect 3107 31723 3153 31775
rect 3167 31723 3213 31775
rect 3213 31723 3219 31775
rect 3101 31654 3107 31706
rect 3107 31654 3153 31706
rect 3167 31654 3213 31706
rect 3213 31654 3219 31706
rect 3101 31584 3107 31636
rect 3107 31584 3153 31636
rect 3167 31584 3213 31636
rect 3213 31584 3219 31636
rect 3101 31514 3107 31566
rect 3107 31514 3153 31566
rect 3167 31514 3213 31566
rect 3213 31514 3219 31566
rect 3101 31444 3107 31496
rect 3107 31444 3153 31496
rect 3167 31444 3213 31496
rect 3213 31444 3219 31496
rect 3101 31380 3107 31426
rect 3107 31380 3153 31426
rect 3167 31380 3213 31426
rect 3213 31380 3219 31426
rect 3101 31374 3153 31380
rect 3167 31374 3219 31380
rect 3378 32714 3430 32720
rect 3378 32680 3384 32714
rect 3384 32680 3418 32714
rect 3418 32680 3430 32714
rect 3378 32668 3430 32680
rect 3444 32714 3496 32720
rect 3444 32680 3456 32714
rect 3456 32680 3490 32714
rect 3490 32680 3496 32714
rect 3444 32668 3496 32680
rect 3378 32641 3430 32651
rect 3378 32607 3384 32641
rect 3384 32607 3418 32641
rect 3418 32607 3430 32641
rect 3378 32599 3430 32607
rect 3444 32641 3496 32651
rect 3444 32607 3456 32641
rect 3456 32607 3490 32641
rect 3490 32607 3496 32641
rect 3444 32599 3496 32607
rect 3378 32568 3430 32582
rect 3378 32534 3384 32568
rect 3384 32534 3418 32568
rect 3418 32534 3430 32568
rect 3378 32530 3430 32534
rect 3444 32568 3496 32582
rect 3444 32534 3456 32568
rect 3456 32534 3490 32568
rect 3490 32534 3496 32568
rect 3444 32530 3496 32534
rect 3378 32495 3430 32513
rect 3378 32461 3384 32495
rect 3384 32461 3418 32495
rect 3418 32461 3430 32495
rect 3444 32495 3496 32513
rect 3444 32461 3456 32495
rect 3456 32461 3490 32495
rect 3490 32461 3496 32495
rect 3378 32422 3430 32444
rect 3444 32422 3496 32444
rect 3378 32392 3384 32422
rect 3384 32392 3430 32422
rect 3444 32392 3490 32422
rect 3490 32392 3496 32422
rect 3378 32323 3384 32375
rect 3384 32323 3430 32375
rect 3444 32323 3490 32375
rect 3490 32323 3496 32375
rect 3378 32254 3384 32306
rect 3384 32254 3430 32306
rect 3444 32254 3490 32306
rect 3490 32254 3496 32306
rect 3378 32184 3384 32236
rect 3384 32184 3430 32236
rect 3444 32184 3490 32236
rect 3490 32184 3496 32236
rect 3378 32114 3384 32166
rect 3384 32114 3430 32166
rect 3444 32114 3490 32166
rect 3490 32114 3496 32166
rect 3655 31930 3661 31982
rect 3661 31930 3707 31982
rect 3721 31930 3767 31982
rect 3767 31930 3773 31982
rect 3655 31861 3661 31913
rect 3661 31861 3707 31913
rect 3721 31861 3767 31913
rect 3767 31861 3773 31913
rect 3655 31792 3661 31844
rect 3661 31792 3707 31844
rect 3721 31792 3767 31844
rect 3767 31792 3773 31844
rect 3655 31723 3661 31775
rect 3661 31723 3707 31775
rect 3721 31723 3767 31775
rect 3767 31723 3773 31775
rect 3655 31654 3661 31706
rect 3661 31654 3707 31706
rect 3721 31654 3767 31706
rect 3767 31654 3773 31706
rect 3655 31584 3661 31636
rect 3661 31584 3707 31636
rect 3721 31584 3767 31636
rect 3767 31584 3773 31636
rect 3655 31514 3661 31566
rect 3661 31514 3707 31566
rect 3721 31514 3767 31566
rect 3767 31514 3773 31566
rect 3655 31444 3661 31496
rect 3661 31444 3707 31496
rect 3721 31444 3767 31496
rect 3767 31444 3773 31496
rect 3655 31380 3661 31426
rect 3661 31380 3707 31426
rect 3721 31380 3767 31426
rect 3767 31380 3773 31426
rect 3655 31374 3707 31380
rect 3721 31374 3773 31380
rect 3932 32714 3984 32720
rect 3932 32680 3938 32714
rect 3938 32680 3972 32714
rect 3972 32680 3984 32714
rect 3932 32668 3984 32680
rect 3998 32714 4050 32720
rect 3998 32680 4010 32714
rect 4010 32680 4044 32714
rect 4044 32680 4050 32714
rect 3998 32668 4050 32680
rect 3932 32641 3984 32651
rect 3932 32607 3938 32641
rect 3938 32607 3972 32641
rect 3972 32607 3984 32641
rect 3932 32599 3984 32607
rect 3998 32641 4050 32651
rect 3998 32607 4010 32641
rect 4010 32607 4044 32641
rect 4044 32607 4050 32641
rect 3998 32599 4050 32607
rect 3932 32568 3984 32582
rect 3932 32534 3938 32568
rect 3938 32534 3972 32568
rect 3972 32534 3984 32568
rect 3932 32530 3984 32534
rect 3998 32568 4050 32582
rect 3998 32534 4010 32568
rect 4010 32534 4044 32568
rect 4044 32534 4050 32568
rect 3998 32530 4050 32534
rect 3932 32495 3984 32513
rect 3932 32461 3938 32495
rect 3938 32461 3972 32495
rect 3972 32461 3984 32495
rect 3998 32495 4050 32513
rect 3998 32461 4010 32495
rect 4010 32461 4044 32495
rect 4044 32461 4050 32495
rect 3932 32422 3984 32444
rect 3998 32422 4050 32444
rect 3932 32392 3938 32422
rect 3938 32392 3984 32422
rect 3998 32392 4044 32422
rect 4044 32392 4050 32422
rect 3932 32323 3938 32375
rect 3938 32323 3984 32375
rect 3998 32323 4044 32375
rect 4044 32323 4050 32375
rect 3932 32254 3938 32306
rect 3938 32254 3984 32306
rect 3998 32254 4044 32306
rect 4044 32254 4050 32306
rect 3932 32184 3938 32236
rect 3938 32184 3984 32236
rect 3998 32184 4044 32236
rect 4044 32184 4050 32236
rect 3932 32114 3938 32166
rect 3938 32114 3984 32166
rect 3998 32114 4044 32166
rect 4044 32114 4050 32166
rect 4209 31930 4215 31982
rect 4215 31930 4261 31982
rect 4275 31930 4321 31982
rect 4321 31930 4327 31982
rect 4209 31861 4215 31913
rect 4215 31861 4261 31913
rect 4275 31861 4321 31913
rect 4321 31861 4327 31913
rect 4209 31792 4215 31844
rect 4215 31792 4261 31844
rect 4275 31792 4321 31844
rect 4321 31792 4327 31844
rect 4209 31723 4215 31775
rect 4215 31723 4261 31775
rect 4275 31723 4321 31775
rect 4321 31723 4327 31775
rect 4209 31654 4215 31706
rect 4215 31654 4261 31706
rect 4275 31654 4321 31706
rect 4321 31654 4327 31706
rect 4209 31584 4215 31636
rect 4215 31584 4261 31636
rect 4275 31584 4321 31636
rect 4321 31584 4327 31636
rect 4209 31514 4215 31566
rect 4215 31514 4261 31566
rect 4275 31514 4321 31566
rect 4321 31514 4327 31566
rect 4209 31444 4215 31496
rect 4215 31444 4261 31496
rect 4275 31444 4321 31496
rect 4321 31444 4327 31496
rect 4209 31380 4215 31426
rect 4215 31380 4261 31426
rect 4275 31380 4321 31426
rect 4321 31380 4327 31426
rect 4209 31374 4261 31380
rect 4275 31374 4327 31380
rect 4486 32714 4538 32720
rect 4486 32680 4492 32714
rect 4492 32680 4526 32714
rect 4526 32680 4538 32714
rect 4486 32668 4538 32680
rect 4552 32714 4604 32720
rect 4552 32680 4564 32714
rect 4564 32680 4598 32714
rect 4598 32680 4604 32714
rect 4552 32668 4604 32680
rect 4486 32641 4538 32651
rect 4486 32607 4492 32641
rect 4492 32607 4526 32641
rect 4526 32607 4538 32641
rect 4486 32599 4538 32607
rect 4552 32641 4604 32651
rect 4552 32607 4564 32641
rect 4564 32607 4598 32641
rect 4598 32607 4604 32641
rect 4552 32599 4604 32607
rect 4486 32568 4538 32582
rect 4486 32534 4492 32568
rect 4492 32534 4526 32568
rect 4526 32534 4538 32568
rect 4486 32530 4538 32534
rect 4552 32568 4604 32582
rect 4552 32534 4564 32568
rect 4564 32534 4598 32568
rect 4598 32534 4604 32568
rect 4552 32530 4604 32534
rect 4486 32495 4538 32513
rect 4486 32461 4492 32495
rect 4492 32461 4526 32495
rect 4526 32461 4538 32495
rect 4552 32495 4604 32513
rect 4552 32461 4564 32495
rect 4564 32461 4598 32495
rect 4598 32461 4604 32495
rect 4486 32422 4538 32444
rect 4552 32422 4604 32444
rect 4486 32392 4492 32422
rect 4492 32392 4538 32422
rect 4552 32392 4598 32422
rect 4598 32392 4604 32422
rect 4486 32323 4492 32375
rect 4492 32323 4538 32375
rect 4552 32323 4598 32375
rect 4598 32323 4604 32375
rect 4486 32254 4492 32306
rect 4492 32254 4538 32306
rect 4552 32254 4598 32306
rect 4598 32254 4604 32306
rect 4486 32184 4492 32236
rect 4492 32184 4538 32236
rect 4552 32184 4598 32236
rect 4598 32184 4604 32236
rect 4486 32114 4492 32166
rect 4492 32114 4538 32166
rect 4552 32114 4598 32166
rect 4598 32114 4604 32166
rect 4763 31930 4769 31982
rect 4769 31930 4815 31982
rect 4829 31930 4875 31982
rect 4875 31930 4881 31982
rect 4763 31861 4769 31913
rect 4769 31861 4815 31913
rect 4829 31861 4875 31913
rect 4875 31861 4881 31913
rect 4763 31792 4769 31844
rect 4769 31792 4815 31844
rect 4829 31792 4875 31844
rect 4875 31792 4881 31844
rect 4763 31723 4769 31775
rect 4769 31723 4815 31775
rect 4829 31723 4875 31775
rect 4875 31723 4881 31775
rect 4763 31654 4769 31706
rect 4769 31654 4815 31706
rect 4829 31654 4875 31706
rect 4875 31654 4881 31706
rect 4763 31584 4769 31636
rect 4769 31584 4815 31636
rect 4829 31584 4875 31636
rect 4875 31584 4881 31636
rect 4763 31514 4769 31566
rect 4769 31514 4815 31566
rect 4829 31514 4875 31566
rect 4875 31514 4881 31566
rect 4763 31444 4769 31496
rect 4769 31444 4815 31496
rect 4829 31444 4875 31496
rect 4875 31444 4881 31496
rect 4763 31380 4769 31426
rect 4769 31380 4815 31426
rect 4829 31380 4875 31426
rect 4875 31380 4881 31426
rect 4763 31374 4815 31380
rect 4829 31374 4881 31380
rect 5040 32714 5092 32720
rect 5040 32680 5046 32714
rect 5046 32680 5080 32714
rect 5080 32680 5092 32714
rect 5040 32668 5092 32680
rect 5106 32714 5158 32720
rect 5106 32680 5118 32714
rect 5118 32680 5152 32714
rect 5152 32680 5158 32714
rect 5106 32668 5158 32680
rect 5040 32641 5092 32651
rect 5040 32607 5046 32641
rect 5046 32607 5080 32641
rect 5080 32607 5092 32641
rect 5040 32599 5092 32607
rect 5106 32641 5158 32651
rect 5106 32607 5118 32641
rect 5118 32607 5152 32641
rect 5152 32607 5158 32641
rect 5106 32599 5158 32607
rect 5040 32568 5092 32582
rect 5040 32534 5046 32568
rect 5046 32534 5080 32568
rect 5080 32534 5092 32568
rect 5040 32530 5092 32534
rect 5106 32568 5158 32582
rect 5106 32534 5118 32568
rect 5118 32534 5152 32568
rect 5152 32534 5158 32568
rect 5106 32530 5158 32534
rect 5040 32495 5092 32513
rect 5040 32461 5046 32495
rect 5046 32461 5080 32495
rect 5080 32461 5092 32495
rect 5106 32495 5158 32513
rect 5106 32461 5118 32495
rect 5118 32461 5152 32495
rect 5152 32461 5158 32495
rect 5040 32422 5092 32444
rect 5106 32422 5158 32444
rect 5040 32392 5046 32422
rect 5046 32392 5092 32422
rect 5106 32392 5152 32422
rect 5152 32392 5158 32422
rect 5040 32323 5046 32375
rect 5046 32323 5092 32375
rect 5106 32323 5152 32375
rect 5152 32323 5158 32375
rect 5040 32254 5046 32306
rect 5046 32254 5092 32306
rect 5106 32254 5152 32306
rect 5152 32254 5158 32306
rect 5040 32184 5046 32236
rect 5046 32184 5092 32236
rect 5106 32184 5152 32236
rect 5152 32184 5158 32236
rect 5040 32114 5046 32166
rect 5046 32114 5092 32166
rect 5106 32114 5152 32166
rect 5152 32114 5158 32166
rect 5317 31930 5323 31982
rect 5323 31930 5369 31982
rect 5383 31930 5429 31982
rect 5429 31930 5435 31982
rect 5317 31861 5323 31913
rect 5323 31861 5369 31913
rect 5383 31861 5429 31913
rect 5429 31861 5435 31913
rect 5317 31792 5323 31844
rect 5323 31792 5369 31844
rect 5383 31792 5429 31844
rect 5429 31792 5435 31844
rect 5317 31723 5323 31775
rect 5323 31723 5369 31775
rect 5383 31723 5429 31775
rect 5429 31723 5435 31775
rect 5317 31654 5323 31706
rect 5323 31654 5369 31706
rect 5383 31654 5429 31706
rect 5429 31654 5435 31706
rect 5317 31584 5323 31636
rect 5323 31584 5369 31636
rect 5383 31584 5429 31636
rect 5429 31584 5435 31636
rect 5317 31514 5323 31566
rect 5323 31514 5369 31566
rect 5383 31514 5429 31566
rect 5429 31514 5435 31566
rect 5317 31444 5323 31496
rect 5323 31444 5369 31496
rect 5383 31444 5429 31496
rect 5429 31444 5435 31496
rect 5317 31380 5323 31426
rect 5323 31380 5369 31426
rect 5383 31380 5429 31426
rect 5429 31380 5435 31426
rect 5317 31374 5369 31380
rect 5383 31374 5435 31380
rect 5594 32714 5646 32720
rect 5594 32680 5600 32714
rect 5600 32680 5634 32714
rect 5634 32680 5646 32714
rect 5594 32668 5646 32680
rect 5660 32714 5712 32720
rect 5660 32680 5672 32714
rect 5672 32680 5706 32714
rect 5706 32680 5712 32714
rect 5660 32668 5712 32680
rect 5594 32641 5646 32651
rect 5594 32607 5600 32641
rect 5600 32607 5634 32641
rect 5634 32607 5646 32641
rect 5594 32599 5646 32607
rect 5660 32641 5712 32651
rect 5660 32607 5672 32641
rect 5672 32607 5706 32641
rect 5706 32607 5712 32641
rect 5660 32599 5712 32607
rect 5594 32568 5646 32582
rect 5594 32534 5600 32568
rect 5600 32534 5634 32568
rect 5634 32534 5646 32568
rect 5594 32530 5646 32534
rect 5660 32568 5712 32582
rect 5660 32534 5672 32568
rect 5672 32534 5706 32568
rect 5706 32534 5712 32568
rect 5660 32530 5712 32534
rect 5594 32495 5646 32513
rect 5594 32461 5600 32495
rect 5600 32461 5634 32495
rect 5634 32461 5646 32495
rect 5660 32495 5712 32513
rect 5660 32461 5672 32495
rect 5672 32461 5706 32495
rect 5706 32461 5712 32495
rect 5594 32422 5646 32444
rect 5660 32422 5712 32444
rect 5594 32392 5600 32422
rect 5600 32392 5646 32422
rect 5660 32392 5706 32422
rect 5706 32392 5712 32422
rect 5594 32323 5600 32375
rect 5600 32323 5646 32375
rect 5660 32323 5706 32375
rect 5706 32323 5712 32375
rect 5594 32254 5600 32306
rect 5600 32254 5646 32306
rect 5660 32254 5706 32306
rect 5706 32254 5712 32306
rect 5594 32184 5600 32236
rect 5600 32184 5646 32236
rect 5660 32184 5706 32236
rect 5706 32184 5712 32236
rect 5594 32114 5600 32166
rect 5600 32114 5646 32166
rect 5660 32114 5706 32166
rect 5706 32114 5712 32166
rect 5871 31930 5877 31982
rect 5877 31930 5923 31982
rect 5937 31930 5983 31982
rect 5983 31930 5989 31982
rect 5871 31861 5877 31913
rect 5877 31861 5923 31913
rect 5937 31861 5983 31913
rect 5983 31861 5989 31913
rect 5871 31792 5877 31844
rect 5877 31792 5923 31844
rect 5937 31792 5983 31844
rect 5983 31792 5989 31844
rect 5871 31723 5877 31775
rect 5877 31723 5923 31775
rect 5937 31723 5983 31775
rect 5983 31723 5989 31775
rect 5871 31654 5877 31706
rect 5877 31654 5923 31706
rect 5937 31654 5983 31706
rect 5983 31654 5989 31706
rect 5871 31584 5877 31636
rect 5877 31584 5923 31636
rect 5937 31584 5983 31636
rect 5983 31584 5989 31636
rect 5871 31514 5877 31566
rect 5877 31514 5923 31566
rect 5937 31514 5983 31566
rect 5983 31514 5989 31566
rect 5871 31444 5877 31496
rect 5877 31444 5923 31496
rect 5937 31444 5983 31496
rect 5983 31444 5989 31496
rect 5871 31380 5877 31426
rect 5877 31380 5923 31426
rect 5937 31380 5983 31426
rect 5983 31380 5989 31426
rect 5871 31374 5923 31380
rect 5937 31374 5989 31380
rect 6148 32714 6200 32720
rect 6148 32680 6154 32714
rect 6154 32680 6188 32714
rect 6188 32680 6200 32714
rect 6148 32668 6200 32680
rect 6214 32714 6266 32720
rect 6214 32680 6226 32714
rect 6226 32680 6260 32714
rect 6260 32680 6266 32714
rect 6214 32668 6266 32680
rect 6148 32641 6200 32651
rect 6148 32607 6154 32641
rect 6154 32607 6188 32641
rect 6188 32607 6200 32641
rect 6148 32599 6200 32607
rect 6214 32641 6266 32651
rect 6214 32607 6226 32641
rect 6226 32607 6260 32641
rect 6260 32607 6266 32641
rect 6214 32599 6266 32607
rect 6148 32568 6200 32582
rect 6148 32534 6154 32568
rect 6154 32534 6188 32568
rect 6188 32534 6200 32568
rect 6148 32530 6200 32534
rect 6214 32568 6266 32582
rect 6214 32534 6226 32568
rect 6226 32534 6260 32568
rect 6260 32534 6266 32568
rect 6214 32530 6266 32534
rect 6148 32495 6200 32513
rect 6148 32461 6154 32495
rect 6154 32461 6188 32495
rect 6188 32461 6200 32495
rect 6214 32495 6266 32513
rect 6214 32461 6226 32495
rect 6226 32461 6260 32495
rect 6260 32461 6266 32495
rect 6148 32422 6200 32444
rect 6214 32422 6266 32444
rect 6148 32392 6154 32422
rect 6154 32392 6200 32422
rect 6214 32392 6260 32422
rect 6260 32392 6266 32422
rect 6148 32323 6154 32375
rect 6154 32323 6200 32375
rect 6214 32323 6260 32375
rect 6260 32323 6266 32375
rect 6148 32254 6154 32306
rect 6154 32254 6200 32306
rect 6214 32254 6260 32306
rect 6260 32254 6266 32306
rect 6148 32184 6154 32236
rect 6154 32184 6200 32236
rect 6214 32184 6260 32236
rect 6260 32184 6266 32236
rect 6148 32114 6154 32166
rect 6154 32114 6200 32166
rect 6214 32114 6260 32166
rect 6260 32114 6266 32166
rect 6425 31930 6431 31982
rect 6431 31930 6477 31982
rect 6491 31930 6537 31982
rect 6537 31930 6543 31982
rect 6425 31861 6431 31913
rect 6431 31861 6477 31913
rect 6491 31861 6537 31913
rect 6537 31861 6543 31913
rect 6425 31792 6431 31844
rect 6431 31792 6477 31844
rect 6491 31792 6537 31844
rect 6537 31792 6543 31844
rect 6425 31723 6431 31775
rect 6431 31723 6477 31775
rect 6491 31723 6537 31775
rect 6537 31723 6543 31775
rect 6425 31654 6431 31706
rect 6431 31654 6477 31706
rect 6491 31654 6537 31706
rect 6537 31654 6543 31706
rect 6425 31584 6431 31636
rect 6431 31584 6477 31636
rect 6491 31584 6537 31636
rect 6537 31584 6543 31636
rect 6425 31514 6431 31566
rect 6431 31514 6477 31566
rect 6491 31514 6537 31566
rect 6537 31514 6543 31566
rect 6425 31444 6431 31496
rect 6431 31444 6477 31496
rect 6491 31444 6537 31496
rect 6537 31444 6543 31496
rect 6425 31380 6431 31426
rect 6431 31380 6477 31426
rect 6491 31380 6537 31426
rect 6537 31380 6543 31426
rect 6425 31374 6477 31380
rect 6491 31374 6543 31380
rect 6702 32714 6754 32720
rect 6702 32680 6708 32714
rect 6708 32680 6742 32714
rect 6742 32680 6754 32714
rect 6702 32668 6754 32680
rect 6768 32714 6820 32720
rect 6768 32680 6780 32714
rect 6780 32680 6814 32714
rect 6814 32680 6820 32714
rect 6768 32668 6820 32680
rect 6702 32641 6754 32651
rect 6702 32607 6708 32641
rect 6708 32607 6742 32641
rect 6742 32607 6754 32641
rect 6702 32599 6754 32607
rect 6768 32641 6820 32651
rect 6768 32607 6780 32641
rect 6780 32607 6814 32641
rect 6814 32607 6820 32641
rect 6768 32599 6820 32607
rect 6702 32568 6754 32582
rect 6702 32534 6708 32568
rect 6708 32534 6742 32568
rect 6742 32534 6754 32568
rect 6702 32530 6754 32534
rect 6768 32568 6820 32582
rect 6768 32534 6780 32568
rect 6780 32534 6814 32568
rect 6814 32534 6820 32568
rect 6768 32530 6820 32534
rect 6702 32495 6754 32513
rect 6702 32461 6708 32495
rect 6708 32461 6742 32495
rect 6742 32461 6754 32495
rect 6768 32495 6820 32513
rect 6768 32461 6780 32495
rect 6780 32461 6814 32495
rect 6814 32461 6820 32495
rect 6702 32422 6754 32444
rect 6768 32422 6820 32444
rect 6702 32392 6708 32422
rect 6708 32392 6754 32422
rect 6768 32392 6814 32422
rect 6814 32392 6820 32422
rect 6702 32323 6708 32375
rect 6708 32323 6754 32375
rect 6768 32323 6814 32375
rect 6814 32323 6820 32375
rect 6702 32254 6708 32306
rect 6708 32254 6754 32306
rect 6768 32254 6814 32306
rect 6814 32254 6820 32306
rect 6702 32184 6708 32236
rect 6708 32184 6754 32236
rect 6768 32184 6814 32236
rect 6814 32184 6820 32236
rect 6702 32114 6708 32166
rect 6708 32114 6754 32166
rect 6768 32114 6814 32166
rect 6814 32114 6820 32166
rect 6979 31930 6985 31982
rect 6985 31930 7031 31982
rect 7045 31930 7091 31982
rect 7091 31930 7097 31982
rect 6979 31861 6985 31913
rect 6985 31861 7031 31913
rect 7045 31861 7091 31913
rect 7091 31861 7097 31913
rect 6979 31792 6985 31844
rect 6985 31792 7031 31844
rect 7045 31792 7091 31844
rect 7091 31792 7097 31844
rect 6979 31723 6985 31775
rect 6985 31723 7031 31775
rect 7045 31723 7091 31775
rect 7091 31723 7097 31775
rect 6979 31654 6985 31706
rect 6985 31654 7031 31706
rect 7045 31654 7091 31706
rect 7091 31654 7097 31706
rect 6979 31584 6985 31636
rect 6985 31584 7031 31636
rect 7045 31584 7091 31636
rect 7091 31584 7097 31636
rect 6979 31514 6985 31566
rect 6985 31514 7031 31566
rect 7045 31514 7091 31566
rect 7091 31514 7097 31566
rect 6979 31444 6985 31496
rect 6985 31444 7031 31496
rect 7045 31444 7091 31496
rect 7091 31444 7097 31496
rect 6979 31380 6985 31426
rect 6985 31380 7031 31426
rect 7045 31380 7091 31426
rect 7091 31380 7097 31426
rect 6979 31374 7031 31380
rect 7045 31374 7097 31380
rect 7256 32714 7308 32720
rect 7256 32680 7262 32714
rect 7262 32680 7296 32714
rect 7296 32680 7308 32714
rect 7256 32668 7308 32680
rect 7322 32714 7374 32720
rect 7322 32680 7334 32714
rect 7334 32680 7368 32714
rect 7368 32680 7374 32714
rect 7322 32668 7374 32680
rect 7256 32641 7308 32651
rect 7256 32607 7262 32641
rect 7262 32607 7296 32641
rect 7296 32607 7308 32641
rect 7256 32599 7308 32607
rect 7322 32641 7374 32651
rect 7322 32607 7334 32641
rect 7334 32607 7368 32641
rect 7368 32607 7374 32641
rect 7322 32599 7374 32607
rect 7256 32568 7308 32582
rect 7256 32534 7262 32568
rect 7262 32534 7296 32568
rect 7296 32534 7308 32568
rect 7256 32530 7308 32534
rect 7322 32568 7374 32582
rect 7322 32534 7334 32568
rect 7334 32534 7368 32568
rect 7368 32534 7374 32568
rect 7322 32530 7374 32534
rect 7256 32495 7308 32513
rect 7256 32461 7262 32495
rect 7262 32461 7296 32495
rect 7296 32461 7308 32495
rect 7322 32495 7374 32513
rect 7322 32461 7334 32495
rect 7334 32461 7368 32495
rect 7368 32461 7374 32495
rect 7256 32422 7308 32444
rect 7322 32422 7374 32444
rect 7256 32392 7262 32422
rect 7262 32392 7308 32422
rect 7322 32392 7368 32422
rect 7368 32392 7374 32422
rect 7256 32323 7262 32375
rect 7262 32323 7308 32375
rect 7322 32323 7368 32375
rect 7368 32323 7374 32375
rect 7256 32254 7262 32306
rect 7262 32254 7308 32306
rect 7322 32254 7368 32306
rect 7368 32254 7374 32306
rect 7256 32184 7262 32236
rect 7262 32184 7308 32236
rect 7322 32184 7368 32236
rect 7368 32184 7374 32236
rect 7256 32114 7262 32166
rect 7262 32114 7308 32166
rect 7322 32114 7368 32166
rect 7368 32114 7374 32166
rect 7533 31930 7539 31982
rect 7539 31930 7585 31982
rect 7599 31930 7645 31982
rect 7645 31930 7651 31982
rect 7533 31861 7539 31913
rect 7539 31861 7585 31913
rect 7599 31861 7645 31913
rect 7645 31861 7651 31913
rect 7533 31792 7539 31844
rect 7539 31792 7585 31844
rect 7599 31792 7645 31844
rect 7645 31792 7651 31844
rect 7533 31723 7539 31775
rect 7539 31723 7585 31775
rect 7599 31723 7645 31775
rect 7645 31723 7651 31775
rect 7533 31654 7539 31706
rect 7539 31654 7585 31706
rect 7599 31654 7645 31706
rect 7645 31654 7651 31706
rect 7533 31584 7539 31636
rect 7539 31584 7585 31636
rect 7599 31584 7645 31636
rect 7645 31584 7651 31636
rect 7533 31514 7539 31566
rect 7539 31514 7585 31566
rect 7599 31514 7645 31566
rect 7645 31514 7651 31566
rect 7533 31444 7539 31496
rect 7539 31444 7585 31496
rect 7599 31444 7645 31496
rect 7645 31444 7651 31496
rect 7533 31380 7539 31426
rect 7539 31380 7585 31426
rect 7599 31380 7645 31426
rect 7645 31380 7651 31426
rect 7533 31374 7585 31380
rect 7599 31374 7651 31380
rect 7810 32714 7862 32720
rect 7810 32680 7816 32714
rect 7816 32680 7850 32714
rect 7850 32680 7862 32714
rect 7810 32668 7862 32680
rect 7876 32714 7928 32720
rect 7876 32680 7888 32714
rect 7888 32680 7922 32714
rect 7922 32680 7928 32714
rect 7876 32668 7928 32680
rect 7810 32641 7862 32651
rect 7810 32607 7816 32641
rect 7816 32607 7850 32641
rect 7850 32607 7862 32641
rect 7810 32599 7862 32607
rect 7876 32641 7928 32651
rect 7876 32607 7888 32641
rect 7888 32607 7922 32641
rect 7922 32607 7928 32641
rect 7876 32599 7928 32607
rect 7810 32568 7862 32582
rect 7810 32534 7816 32568
rect 7816 32534 7850 32568
rect 7850 32534 7862 32568
rect 7810 32530 7862 32534
rect 7876 32568 7928 32582
rect 7876 32534 7888 32568
rect 7888 32534 7922 32568
rect 7922 32534 7928 32568
rect 7876 32530 7928 32534
rect 7810 32495 7862 32513
rect 7810 32461 7816 32495
rect 7816 32461 7850 32495
rect 7850 32461 7862 32495
rect 7876 32495 7928 32513
rect 7876 32461 7888 32495
rect 7888 32461 7922 32495
rect 7922 32461 7928 32495
rect 7810 32422 7862 32444
rect 7876 32422 7928 32444
rect 7810 32392 7816 32422
rect 7816 32392 7862 32422
rect 7876 32392 7922 32422
rect 7922 32392 7928 32422
rect 7810 32323 7816 32375
rect 7816 32323 7862 32375
rect 7876 32323 7922 32375
rect 7922 32323 7928 32375
rect 7810 32254 7816 32306
rect 7816 32254 7862 32306
rect 7876 32254 7922 32306
rect 7922 32254 7928 32306
rect 7810 32184 7816 32236
rect 7816 32184 7862 32236
rect 7876 32184 7922 32236
rect 7922 32184 7928 32236
rect 7810 32114 7816 32166
rect 7816 32114 7862 32166
rect 7876 32114 7922 32166
rect 7922 32114 7928 32166
rect 8047 32709 8050 32724
rect 8050 32709 8084 32724
rect 8084 32709 8099 32724
rect 8047 32672 8099 32709
rect 8169 32699 8184 32724
rect 8184 32699 8218 32724
rect 8218 32699 8221 32724
rect 8169 32672 8221 32699
rect 8047 32637 8050 32655
rect 8050 32637 8084 32655
rect 8084 32637 8099 32655
rect 8047 32603 8099 32637
rect 8169 32627 8184 32655
rect 8184 32627 8218 32655
rect 8218 32627 8221 32655
rect 8169 32603 8221 32627
rect 8047 32565 8050 32586
rect 8050 32565 8084 32586
rect 8084 32565 8099 32586
rect 8047 32534 8099 32565
rect 8169 32555 8184 32586
rect 8184 32555 8218 32586
rect 8218 32555 8221 32586
rect 8169 32534 8221 32555
rect 8047 32493 8050 32517
rect 8050 32493 8084 32517
rect 8084 32493 8099 32517
rect 8047 32465 8099 32493
rect 8169 32483 8184 32517
rect 8184 32483 8218 32517
rect 8218 32483 8221 32517
rect 8169 32465 8221 32483
rect 8047 32421 8050 32448
rect 8050 32421 8084 32448
rect 8084 32421 8099 32448
rect 8047 32396 8099 32421
rect 8169 32445 8221 32448
rect 8169 32411 8184 32445
rect 8184 32411 8218 32445
rect 8218 32411 8221 32445
rect 8169 32396 8221 32411
rect 8047 32349 8050 32378
rect 8050 32349 8084 32378
rect 8084 32349 8099 32378
rect 8047 32326 8099 32349
rect 8169 32373 8221 32378
rect 8169 32339 8184 32373
rect 8184 32339 8218 32373
rect 8218 32339 8221 32373
rect 8169 32326 8221 32339
rect 8047 32277 8050 32308
rect 8050 32277 8084 32308
rect 8084 32277 8099 32308
rect 8047 32256 8099 32277
rect 8169 32301 8221 32308
rect 8169 32267 8184 32301
rect 8184 32267 8218 32301
rect 8218 32267 8221 32301
rect 8169 32256 8221 32267
rect 8047 32205 8050 32238
rect 8050 32205 8084 32238
rect 8084 32205 8099 32238
rect 8047 32186 8099 32205
rect 8169 32229 8221 32238
rect 8169 32195 8184 32229
rect 8184 32195 8218 32229
rect 8218 32195 8221 32229
rect 8169 32186 8221 32195
rect 8047 32167 8099 32168
rect 8047 32133 8050 32167
rect 8050 32133 8084 32167
rect 8084 32133 8099 32167
rect 8047 32116 8099 32133
rect 8169 32157 8221 32168
rect 8169 32123 8184 32157
rect 8184 32123 8218 32157
rect 8218 32123 8221 32157
rect 8169 32116 8221 32123
rect 2824 30714 2876 30720
rect 2824 30680 2830 30714
rect 2830 30680 2864 30714
rect 2864 30680 2876 30714
rect 2824 30668 2876 30680
rect 2890 30714 2942 30720
rect 2890 30680 2902 30714
rect 2902 30680 2936 30714
rect 2936 30680 2942 30714
rect 2890 30668 2942 30680
rect 2824 30641 2876 30651
rect 2824 30607 2830 30641
rect 2830 30607 2864 30641
rect 2864 30607 2876 30641
rect 2824 30599 2876 30607
rect 2890 30641 2942 30651
rect 2890 30607 2902 30641
rect 2902 30607 2936 30641
rect 2936 30607 2942 30641
rect 2890 30599 2942 30607
rect 2824 30568 2876 30582
rect 2824 30534 2830 30568
rect 2830 30534 2864 30568
rect 2864 30534 2876 30568
rect 2824 30530 2876 30534
rect 2890 30568 2942 30582
rect 2890 30534 2902 30568
rect 2902 30534 2936 30568
rect 2936 30534 2942 30568
rect 2890 30530 2942 30534
rect 2824 30495 2876 30513
rect 2824 30461 2830 30495
rect 2830 30461 2864 30495
rect 2864 30461 2876 30495
rect 2890 30495 2942 30513
rect 2890 30461 2902 30495
rect 2902 30461 2936 30495
rect 2936 30461 2942 30495
rect 2824 30422 2876 30444
rect 2890 30422 2942 30444
rect 2824 30392 2830 30422
rect 2830 30392 2876 30422
rect 2890 30392 2936 30422
rect 2936 30392 2942 30422
rect 2824 30323 2830 30375
rect 2830 30323 2876 30375
rect 2890 30323 2936 30375
rect 2936 30323 2942 30375
rect 2824 30254 2830 30306
rect 2830 30254 2876 30306
rect 2890 30254 2936 30306
rect 2936 30254 2942 30306
rect 2824 30184 2830 30236
rect 2830 30184 2876 30236
rect 2890 30184 2936 30236
rect 2936 30184 2942 30236
rect 2824 30114 2830 30166
rect 2830 30114 2876 30166
rect 2890 30114 2936 30166
rect 2936 30114 2942 30166
rect 3101 29930 3107 29982
rect 3107 29930 3153 29982
rect 3167 29930 3213 29982
rect 3213 29930 3219 29982
rect 3101 29861 3107 29913
rect 3107 29861 3153 29913
rect 3167 29861 3213 29913
rect 3213 29861 3219 29913
rect 3101 29792 3107 29844
rect 3107 29792 3153 29844
rect 3167 29792 3213 29844
rect 3213 29792 3219 29844
rect 3101 29723 3107 29775
rect 3107 29723 3153 29775
rect 3167 29723 3213 29775
rect 3213 29723 3219 29775
rect 3101 29654 3107 29706
rect 3107 29654 3153 29706
rect 3167 29654 3213 29706
rect 3213 29654 3219 29706
rect 3101 29584 3107 29636
rect 3107 29584 3153 29636
rect 3167 29584 3213 29636
rect 3213 29584 3219 29636
rect 3101 29514 3107 29566
rect 3107 29514 3153 29566
rect 3167 29514 3213 29566
rect 3213 29514 3219 29566
rect 3101 29444 3107 29496
rect 3107 29444 3153 29496
rect 3167 29444 3213 29496
rect 3213 29444 3219 29496
rect 3101 29380 3107 29426
rect 3107 29380 3153 29426
rect 3167 29380 3213 29426
rect 3213 29380 3219 29426
rect 3101 29374 3153 29380
rect 3167 29374 3219 29380
rect 3378 30714 3430 30720
rect 3378 30680 3384 30714
rect 3384 30680 3418 30714
rect 3418 30680 3430 30714
rect 3378 30668 3430 30680
rect 3444 30714 3496 30720
rect 3444 30680 3456 30714
rect 3456 30680 3490 30714
rect 3490 30680 3496 30714
rect 3444 30668 3496 30680
rect 3378 30641 3430 30651
rect 3378 30607 3384 30641
rect 3384 30607 3418 30641
rect 3418 30607 3430 30641
rect 3378 30599 3430 30607
rect 3444 30641 3496 30651
rect 3444 30607 3456 30641
rect 3456 30607 3490 30641
rect 3490 30607 3496 30641
rect 3444 30599 3496 30607
rect 3378 30568 3430 30582
rect 3378 30534 3384 30568
rect 3384 30534 3418 30568
rect 3418 30534 3430 30568
rect 3378 30530 3430 30534
rect 3444 30568 3496 30582
rect 3444 30534 3456 30568
rect 3456 30534 3490 30568
rect 3490 30534 3496 30568
rect 3444 30530 3496 30534
rect 3378 30495 3430 30513
rect 3378 30461 3384 30495
rect 3384 30461 3418 30495
rect 3418 30461 3430 30495
rect 3444 30495 3496 30513
rect 3444 30461 3456 30495
rect 3456 30461 3490 30495
rect 3490 30461 3496 30495
rect 3378 30422 3430 30444
rect 3444 30422 3496 30444
rect 3378 30392 3384 30422
rect 3384 30392 3430 30422
rect 3444 30392 3490 30422
rect 3490 30392 3496 30422
rect 3378 30323 3384 30375
rect 3384 30323 3430 30375
rect 3444 30323 3490 30375
rect 3490 30323 3496 30375
rect 3378 30254 3384 30306
rect 3384 30254 3430 30306
rect 3444 30254 3490 30306
rect 3490 30254 3496 30306
rect 3378 30184 3384 30236
rect 3384 30184 3430 30236
rect 3444 30184 3490 30236
rect 3490 30184 3496 30236
rect 3378 30114 3384 30166
rect 3384 30114 3430 30166
rect 3444 30114 3490 30166
rect 3490 30114 3496 30166
rect 3655 29930 3661 29982
rect 3661 29930 3707 29982
rect 3721 29930 3767 29982
rect 3767 29930 3773 29982
rect 3655 29861 3661 29913
rect 3661 29861 3707 29913
rect 3721 29861 3767 29913
rect 3767 29861 3773 29913
rect 3655 29792 3661 29844
rect 3661 29792 3707 29844
rect 3721 29792 3767 29844
rect 3767 29792 3773 29844
rect 3655 29723 3661 29775
rect 3661 29723 3707 29775
rect 3721 29723 3767 29775
rect 3767 29723 3773 29775
rect 3655 29654 3661 29706
rect 3661 29654 3707 29706
rect 3721 29654 3767 29706
rect 3767 29654 3773 29706
rect 3655 29584 3661 29636
rect 3661 29584 3707 29636
rect 3721 29584 3767 29636
rect 3767 29584 3773 29636
rect 3655 29514 3661 29566
rect 3661 29514 3707 29566
rect 3721 29514 3767 29566
rect 3767 29514 3773 29566
rect 3655 29444 3661 29496
rect 3661 29444 3707 29496
rect 3721 29444 3767 29496
rect 3767 29444 3773 29496
rect 3655 29380 3661 29426
rect 3661 29380 3707 29426
rect 3721 29380 3767 29426
rect 3767 29380 3773 29426
rect 3655 29374 3707 29380
rect 3721 29374 3773 29380
rect 3932 30714 3984 30720
rect 3932 30680 3938 30714
rect 3938 30680 3972 30714
rect 3972 30680 3984 30714
rect 3932 30668 3984 30680
rect 3998 30714 4050 30720
rect 3998 30680 4010 30714
rect 4010 30680 4044 30714
rect 4044 30680 4050 30714
rect 3998 30668 4050 30680
rect 3932 30641 3984 30651
rect 3932 30607 3938 30641
rect 3938 30607 3972 30641
rect 3972 30607 3984 30641
rect 3932 30599 3984 30607
rect 3998 30641 4050 30651
rect 3998 30607 4010 30641
rect 4010 30607 4044 30641
rect 4044 30607 4050 30641
rect 3998 30599 4050 30607
rect 3932 30568 3984 30582
rect 3932 30534 3938 30568
rect 3938 30534 3972 30568
rect 3972 30534 3984 30568
rect 3932 30530 3984 30534
rect 3998 30568 4050 30582
rect 3998 30534 4010 30568
rect 4010 30534 4044 30568
rect 4044 30534 4050 30568
rect 3998 30530 4050 30534
rect 3932 30495 3984 30513
rect 3932 30461 3938 30495
rect 3938 30461 3972 30495
rect 3972 30461 3984 30495
rect 3998 30495 4050 30513
rect 3998 30461 4010 30495
rect 4010 30461 4044 30495
rect 4044 30461 4050 30495
rect 3932 30422 3984 30444
rect 3998 30422 4050 30444
rect 3932 30392 3938 30422
rect 3938 30392 3984 30422
rect 3998 30392 4044 30422
rect 4044 30392 4050 30422
rect 3932 30323 3938 30375
rect 3938 30323 3984 30375
rect 3998 30323 4044 30375
rect 4044 30323 4050 30375
rect 3932 30254 3938 30306
rect 3938 30254 3984 30306
rect 3998 30254 4044 30306
rect 4044 30254 4050 30306
rect 3932 30184 3938 30236
rect 3938 30184 3984 30236
rect 3998 30184 4044 30236
rect 4044 30184 4050 30236
rect 3932 30114 3938 30166
rect 3938 30114 3984 30166
rect 3998 30114 4044 30166
rect 4044 30114 4050 30166
rect 4209 29930 4215 29982
rect 4215 29930 4261 29982
rect 4275 29930 4321 29982
rect 4321 29930 4327 29982
rect 4209 29861 4215 29913
rect 4215 29861 4261 29913
rect 4275 29861 4321 29913
rect 4321 29861 4327 29913
rect 4209 29792 4215 29844
rect 4215 29792 4261 29844
rect 4275 29792 4321 29844
rect 4321 29792 4327 29844
rect 4209 29723 4215 29775
rect 4215 29723 4261 29775
rect 4275 29723 4321 29775
rect 4321 29723 4327 29775
rect 4209 29654 4215 29706
rect 4215 29654 4261 29706
rect 4275 29654 4321 29706
rect 4321 29654 4327 29706
rect 4209 29584 4215 29636
rect 4215 29584 4261 29636
rect 4275 29584 4321 29636
rect 4321 29584 4327 29636
rect 4209 29514 4215 29566
rect 4215 29514 4261 29566
rect 4275 29514 4321 29566
rect 4321 29514 4327 29566
rect 4209 29444 4215 29496
rect 4215 29444 4261 29496
rect 4275 29444 4321 29496
rect 4321 29444 4327 29496
rect 4209 29380 4215 29426
rect 4215 29380 4261 29426
rect 4275 29380 4321 29426
rect 4321 29380 4327 29426
rect 4209 29374 4261 29380
rect 4275 29374 4327 29380
rect 4486 30714 4538 30720
rect 4486 30680 4492 30714
rect 4492 30680 4526 30714
rect 4526 30680 4538 30714
rect 4486 30668 4538 30680
rect 4552 30714 4604 30720
rect 4552 30680 4564 30714
rect 4564 30680 4598 30714
rect 4598 30680 4604 30714
rect 4552 30668 4604 30680
rect 4486 30641 4538 30651
rect 4486 30607 4492 30641
rect 4492 30607 4526 30641
rect 4526 30607 4538 30641
rect 4486 30599 4538 30607
rect 4552 30641 4604 30651
rect 4552 30607 4564 30641
rect 4564 30607 4598 30641
rect 4598 30607 4604 30641
rect 4552 30599 4604 30607
rect 4486 30568 4538 30582
rect 4486 30534 4492 30568
rect 4492 30534 4526 30568
rect 4526 30534 4538 30568
rect 4486 30530 4538 30534
rect 4552 30568 4604 30582
rect 4552 30534 4564 30568
rect 4564 30534 4598 30568
rect 4598 30534 4604 30568
rect 4552 30530 4604 30534
rect 4486 30495 4538 30513
rect 4486 30461 4492 30495
rect 4492 30461 4526 30495
rect 4526 30461 4538 30495
rect 4552 30495 4604 30513
rect 4552 30461 4564 30495
rect 4564 30461 4598 30495
rect 4598 30461 4604 30495
rect 4486 30422 4538 30444
rect 4552 30422 4604 30444
rect 4486 30392 4492 30422
rect 4492 30392 4538 30422
rect 4552 30392 4598 30422
rect 4598 30392 4604 30422
rect 4486 30323 4492 30375
rect 4492 30323 4538 30375
rect 4552 30323 4598 30375
rect 4598 30323 4604 30375
rect 4486 30254 4492 30306
rect 4492 30254 4538 30306
rect 4552 30254 4598 30306
rect 4598 30254 4604 30306
rect 4486 30184 4492 30236
rect 4492 30184 4538 30236
rect 4552 30184 4598 30236
rect 4598 30184 4604 30236
rect 4486 30114 4492 30166
rect 4492 30114 4538 30166
rect 4552 30114 4598 30166
rect 4598 30114 4604 30166
rect 4763 29930 4769 29982
rect 4769 29930 4815 29982
rect 4829 29930 4875 29982
rect 4875 29930 4881 29982
rect 4763 29861 4769 29913
rect 4769 29861 4815 29913
rect 4829 29861 4875 29913
rect 4875 29861 4881 29913
rect 4763 29792 4769 29844
rect 4769 29792 4815 29844
rect 4829 29792 4875 29844
rect 4875 29792 4881 29844
rect 4763 29723 4769 29775
rect 4769 29723 4815 29775
rect 4829 29723 4875 29775
rect 4875 29723 4881 29775
rect 4763 29654 4769 29706
rect 4769 29654 4815 29706
rect 4829 29654 4875 29706
rect 4875 29654 4881 29706
rect 4763 29584 4769 29636
rect 4769 29584 4815 29636
rect 4829 29584 4875 29636
rect 4875 29584 4881 29636
rect 4763 29514 4769 29566
rect 4769 29514 4815 29566
rect 4829 29514 4875 29566
rect 4875 29514 4881 29566
rect 4763 29444 4769 29496
rect 4769 29444 4815 29496
rect 4829 29444 4875 29496
rect 4875 29444 4881 29496
rect 4763 29380 4769 29426
rect 4769 29380 4815 29426
rect 4829 29380 4875 29426
rect 4875 29380 4881 29426
rect 4763 29374 4815 29380
rect 4829 29374 4881 29380
rect 5040 30714 5092 30720
rect 5040 30680 5046 30714
rect 5046 30680 5080 30714
rect 5080 30680 5092 30714
rect 5040 30668 5092 30680
rect 5106 30714 5158 30720
rect 5106 30680 5118 30714
rect 5118 30680 5152 30714
rect 5152 30680 5158 30714
rect 5106 30668 5158 30680
rect 5040 30641 5092 30651
rect 5040 30607 5046 30641
rect 5046 30607 5080 30641
rect 5080 30607 5092 30641
rect 5040 30599 5092 30607
rect 5106 30641 5158 30651
rect 5106 30607 5118 30641
rect 5118 30607 5152 30641
rect 5152 30607 5158 30641
rect 5106 30599 5158 30607
rect 5040 30568 5092 30582
rect 5040 30534 5046 30568
rect 5046 30534 5080 30568
rect 5080 30534 5092 30568
rect 5040 30530 5092 30534
rect 5106 30568 5158 30582
rect 5106 30534 5118 30568
rect 5118 30534 5152 30568
rect 5152 30534 5158 30568
rect 5106 30530 5158 30534
rect 5040 30495 5092 30513
rect 5040 30461 5046 30495
rect 5046 30461 5080 30495
rect 5080 30461 5092 30495
rect 5106 30495 5158 30513
rect 5106 30461 5118 30495
rect 5118 30461 5152 30495
rect 5152 30461 5158 30495
rect 5040 30422 5092 30444
rect 5106 30422 5158 30444
rect 5040 30392 5046 30422
rect 5046 30392 5092 30422
rect 5106 30392 5152 30422
rect 5152 30392 5158 30422
rect 5040 30323 5046 30375
rect 5046 30323 5092 30375
rect 5106 30323 5152 30375
rect 5152 30323 5158 30375
rect 5040 30254 5046 30306
rect 5046 30254 5092 30306
rect 5106 30254 5152 30306
rect 5152 30254 5158 30306
rect 5040 30184 5046 30236
rect 5046 30184 5092 30236
rect 5106 30184 5152 30236
rect 5152 30184 5158 30236
rect 5040 30114 5046 30166
rect 5046 30114 5092 30166
rect 5106 30114 5152 30166
rect 5152 30114 5158 30166
rect 5317 29930 5323 29982
rect 5323 29930 5369 29982
rect 5383 29930 5429 29982
rect 5429 29930 5435 29982
rect 5317 29861 5323 29913
rect 5323 29861 5369 29913
rect 5383 29861 5429 29913
rect 5429 29861 5435 29913
rect 5317 29792 5323 29844
rect 5323 29792 5369 29844
rect 5383 29792 5429 29844
rect 5429 29792 5435 29844
rect 5317 29723 5323 29775
rect 5323 29723 5369 29775
rect 5383 29723 5429 29775
rect 5429 29723 5435 29775
rect 5317 29654 5323 29706
rect 5323 29654 5369 29706
rect 5383 29654 5429 29706
rect 5429 29654 5435 29706
rect 5317 29584 5323 29636
rect 5323 29584 5369 29636
rect 5383 29584 5429 29636
rect 5429 29584 5435 29636
rect 5317 29514 5323 29566
rect 5323 29514 5369 29566
rect 5383 29514 5429 29566
rect 5429 29514 5435 29566
rect 5317 29444 5323 29496
rect 5323 29444 5369 29496
rect 5383 29444 5429 29496
rect 5429 29444 5435 29496
rect 5317 29380 5323 29426
rect 5323 29380 5369 29426
rect 5383 29380 5429 29426
rect 5429 29380 5435 29426
rect 5317 29374 5369 29380
rect 5383 29374 5435 29380
rect 5594 30714 5646 30720
rect 5594 30680 5600 30714
rect 5600 30680 5634 30714
rect 5634 30680 5646 30714
rect 5594 30668 5646 30680
rect 5660 30714 5712 30720
rect 5660 30680 5672 30714
rect 5672 30680 5706 30714
rect 5706 30680 5712 30714
rect 5660 30668 5712 30680
rect 5594 30641 5646 30651
rect 5594 30607 5600 30641
rect 5600 30607 5634 30641
rect 5634 30607 5646 30641
rect 5594 30599 5646 30607
rect 5660 30641 5712 30651
rect 5660 30607 5672 30641
rect 5672 30607 5706 30641
rect 5706 30607 5712 30641
rect 5660 30599 5712 30607
rect 5594 30568 5646 30582
rect 5594 30534 5600 30568
rect 5600 30534 5634 30568
rect 5634 30534 5646 30568
rect 5594 30530 5646 30534
rect 5660 30568 5712 30582
rect 5660 30534 5672 30568
rect 5672 30534 5706 30568
rect 5706 30534 5712 30568
rect 5660 30530 5712 30534
rect 5594 30495 5646 30513
rect 5594 30461 5600 30495
rect 5600 30461 5634 30495
rect 5634 30461 5646 30495
rect 5660 30495 5712 30513
rect 5660 30461 5672 30495
rect 5672 30461 5706 30495
rect 5706 30461 5712 30495
rect 5594 30422 5646 30444
rect 5660 30422 5712 30444
rect 5594 30392 5600 30422
rect 5600 30392 5646 30422
rect 5660 30392 5706 30422
rect 5706 30392 5712 30422
rect 5594 30323 5600 30375
rect 5600 30323 5646 30375
rect 5660 30323 5706 30375
rect 5706 30323 5712 30375
rect 5594 30254 5600 30306
rect 5600 30254 5646 30306
rect 5660 30254 5706 30306
rect 5706 30254 5712 30306
rect 5594 30184 5600 30236
rect 5600 30184 5646 30236
rect 5660 30184 5706 30236
rect 5706 30184 5712 30236
rect 5594 30114 5600 30166
rect 5600 30114 5646 30166
rect 5660 30114 5706 30166
rect 5706 30114 5712 30166
rect 5871 29930 5877 29982
rect 5877 29930 5923 29982
rect 5937 29930 5983 29982
rect 5983 29930 5989 29982
rect 5871 29861 5877 29913
rect 5877 29861 5923 29913
rect 5937 29861 5983 29913
rect 5983 29861 5989 29913
rect 5871 29792 5877 29844
rect 5877 29792 5923 29844
rect 5937 29792 5983 29844
rect 5983 29792 5989 29844
rect 5871 29723 5877 29775
rect 5877 29723 5923 29775
rect 5937 29723 5983 29775
rect 5983 29723 5989 29775
rect 5871 29654 5877 29706
rect 5877 29654 5923 29706
rect 5937 29654 5983 29706
rect 5983 29654 5989 29706
rect 5871 29584 5877 29636
rect 5877 29584 5923 29636
rect 5937 29584 5983 29636
rect 5983 29584 5989 29636
rect 5871 29514 5877 29566
rect 5877 29514 5923 29566
rect 5937 29514 5983 29566
rect 5983 29514 5989 29566
rect 5871 29444 5877 29496
rect 5877 29444 5923 29496
rect 5937 29444 5983 29496
rect 5983 29444 5989 29496
rect 5871 29380 5877 29426
rect 5877 29380 5923 29426
rect 5937 29380 5983 29426
rect 5983 29380 5989 29426
rect 5871 29374 5923 29380
rect 5937 29374 5989 29380
rect 6148 30714 6200 30720
rect 6148 30680 6154 30714
rect 6154 30680 6188 30714
rect 6188 30680 6200 30714
rect 6148 30668 6200 30680
rect 6214 30714 6266 30720
rect 6214 30680 6226 30714
rect 6226 30680 6260 30714
rect 6260 30680 6266 30714
rect 6214 30668 6266 30680
rect 6148 30641 6200 30651
rect 6148 30607 6154 30641
rect 6154 30607 6188 30641
rect 6188 30607 6200 30641
rect 6148 30599 6200 30607
rect 6214 30641 6266 30651
rect 6214 30607 6226 30641
rect 6226 30607 6260 30641
rect 6260 30607 6266 30641
rect 6214 30599 6266 30607
rect 6148 30568 6200 30582
rect 6148 30534 6154 30568
rect 6154 30534 6188 30568
rect 6188 30534 6200 30568
rect 6148 30530 6200 30534
rect 6214 30568 6266 30582
rect 6214 30534 6226 30568
rect 6226 30534 6260 30568
rect 6260 30534 6266 30568
rect 6214 30530 6266 30534
rect 6148 30495 6200 30513
rect 6148 30461 6154 30495
rect 6154 30461 6188 30495
rect 6188 30461 6200 30495
rect 6214 30495 6266 30513
rect 6214 30461 6226 30495
rect 6226 30461 6260 30495
rect 6260 30461 6266 30495
rect 6148 30422 6200 30444
rect 6214 30422 6266 30444
rect 6148 30392 6154 30422
rect 6154 30392 6200 30422
rect 6214 30392 6260 30422
rect 6260 30392 6266 30422
rect 6148 30323 6154 30375
rect 6154 30323 6200 30375
rect 6214 30323 6260 30375
rect 6260 30323 6266 30375
rect 6148 30254 6154 30306
rect 6154 30254 6200 30306
rect 6214 30254 6260 30306
rect 6260 30254 6266 30306
rect 6148 30184 6154 30236
rect 6154 30184 6200 30236
rect 6214 30184 6260 30236
rect 6260 30184 6266 30236
rect 6148 30114 6154 30166
rect 6154 30114 6200 30166
rect 6214 30114 6260 30166
rect 6260 30114 6266 30166
rect 6425 29930 6431 29982
rect 6431 29930 6477 29982
rect 6491 29930 6537 29982
rect 6537 29930 6543 29982
rect 6425 29861 6431 29913
rect 6431 29861 6477 29913
rect 6491 29861 6537 29913
rect 6537 29861 6543 29913
rect 6425 29792 6431 29844
rect 6431 29792 6477 29844
rect 6491 29792 6537 29844
rect 6537 29792 6543 29844
rect 6425 29723 6431 29775
rect 6431 29723 6477 29775
rect 6491 29723 6537 29775
rect 6537 29723 6543 29775
rect 6425 29654 6431 29706
rect 6431 29654 6477 29706
rect 6491 29654 6537 29706
rect 6537 29654 6543 29706
rect 6425 29584 6431 29636
rect 6431 29584 6477 29636
rect 6491 29584 6537 29636
rect 6537 29584 6543 29636
rect 6425 29514 6431 29566
rect 6431 29514 6477 29566
rect 6491 29514 6537 29566
rect 6537 29514 6543 29566
rect 6425 29444 6431 29496
rect 6431 29444 6477 29496
rect 6491 29444 6537 29496
rect 6537 29444 6543 29496
rect 6425 29380 6431 29426
rect 6431 29380 6477 29426
rect 6491 29380 6537 29426
rect 6537 29380 6543 29426
rect 6425 29374 6477 29380
rect 6491 29374 6543 29380
rect 6702 30714 6754 30720
rect 6702 30680 6708 30714
rect 6708 30680 6742 30714
rect 6742 30680 6754 30714
rect 6702 30668 6754 30680
rect 6768 30714 6820 30720
rect 6768 30680 6780 30714
rect 6780 30680 6814 30714
rect 6814 30680 6820 30714
rect 6768 30668 6820 30680
rect 6702 30641 6754 30651
rect 6702 30607 6708 30641
rect 6708 30607 6742 30641
rect 6742 30607 6754 30641
rect 6702 30599 6754 30607
rect 6768 30641 6820 30651
rect 6768 30607 6780 30641
rect 6780 30607 6814 30641
rect 6814 30607 6820 30641
rect 6768 30599 6820 30607
rect 6702 30568 6754 30582
rect 6702 30534 6708 30568
rect 6708 30534 6742 30568
rect 6742 30534 6754 30568
rect 6702 30530 6754 30534
rect 6768 30568 6820 30582
rect 6768 30534 6780 30568
rect 6780 30534 6814 30568
rect 6814 30534 6820 30568
rect 6768 30530 6820 30534
rect 6702 30495 6754 30513
rect 6702 30461 6708 30495
rect 6708 30461 6742 30495
rect 6742 30461 6754 30495
rect 6768 30495 6820 30513
rect 6768 30461 6780 30495
rect 6780 30461 6814 30495
rect 6814 30461 6820 30495
rect 6702 30422 6754 30444
rect 6768 30422 6820 30444
rect 6702 30392 6708 30422
rect 6708 30392 6754 30422
rect 6768 30392 6814 30422
rect 6814 30392 6820 30422
rect 6702 30323 6708 30375
rect 6708 30323 6754 30375
rect 6768 30323 6814 30375
rect 6814 30323 6820 30375
rect 6702 30254 6708 30306
rect 6708 30254 6754 30306
rect 6768 30254 6814 30306
rect 6814 30254 6820 30306
rect 6702 30184 6708 30236
rect 6708 30184 6754 30236
rect 6768 30184 6814 30236
rect 6814 30184 6820 30236
rect 6702 30114 6708 30166
rect 6708 30114 6754 30166
rect 6768 30114 6814 30166
rect 6814 30114 6820 30166
rect 6979 29930 6985 29982
rect 6985 29930 7031 29982
rect 7045 29930 7091 29982
rect 7091 29930 7097 29982
rect 6979 29861 6985 29913
rect 6985 29861 7031 29913
rect 7045 29861 7091 29913
rect 7091 29861 7097 29913
rect 6979 29792 6985 29844
rect 6985 29792 7031 29844
rect 7045 29792 7091 29844
rect 7091 29792 7097 29844
rect 6979 29723 6985 29775
rect 6985 29723 7031 29775
rect 7045 29723 7091 29775
rect 7091 29723 7097 29775
rect 6979 29654 6985 29706
rect 6985 29654 7031 29706
rect 7045 29654 7091 29706
rect 7091 29654 7097 29706
rect 6979 29584 6985 29636
rect 6985 29584 7031 29636
rect 7045 29584 7091 29636
rect 7091 29584 7097 29636
rect 6979 29514 6985 29566
rect 6985 29514 7031 29566
rect 7045 29514 7091 29566
rect 7091 29514 7097 29566
rect 6979 29444 6985 29496
rect 6985 29444 7031 29496
rect 7045 29444 7091 29496
rect 7091 29444 7097 29496
rect 6979 29380 6985 29426
rect 6985 29380 7031 29426
rect 7045 29380 7091 29426
rect 7091 29380 7097 29426
rect 6979 29374 7031 29380
rect 7045 29374 7097 29380
rect 7256 30714 7308 30720
rect 7256 30680 7262 30714
rect 7262 30680 7296 30714
rect 7296 30680 7308 30714
rect 7256 30668 7308 30680
rect 7322 30714 7374 30720
rect 7322 30680 7334 30714
rect 7334 30680 7368 30714
rect 7368 30680 7374 30714
rect 7322 30668 7374 30680
rect 7256 30641 7308 30651
rect 7256 30607 7262 30641
rect 7262 30607 7296 30641
rect 7296 30607 7308 30641
rect 7256 30599 7308 30607
rect 7322 30641 7374 30651
rect 7322 30607 7334 30641
rect 7334 30607 7368 30641
rect 7368 30607 7374 30641
rect 7322 30599 7374 30607
rect 7256 30568 7308 30582
rect 7256 30534 7262 30568
rect 7262 30534 7296 30568
rect 7296 30534 7308 30568
rect 7256 30530 7308 30534
rect 7322 30568 7374 30582
rect 7322 30534 7334 30568
rect 7334 30534 7368 30568
rect 7368 30534 7374 30568
rect 7322 30530 7374 30534
rect 7256 30495 7308 30513
rect 7256 30461 7262 30495
rect 7262 30461 7296 30495
rect 7296 30461 7308 30495
rect 7322 30495 7374 30513
rect 7322 30461 7334 30495
rect 7334 30461 7368 30495
rect 7368 30461 7374 30495
rect 7256 30422 7308 30444
rect 7322 30422 7374 30444
rect 7256 30392 7262 30422
rect 7262 30392 7308 30422
rect 7322 30392 7368 30422
rect 7368 30392 7374 30422
rect 7256 30323 7262 30375
rect 7262 30323 7308 30375
rect 7322 30323 7368 30375
rect 7368 30323 7374 30375
rect 7256 30254 7262 30306
rect 7262 30254 7308 30306
rect 7322 30254 7368 30306
rect 7368 30254 7374 30306
rect 7256 30184 7262 30236
rect 7262 30184 7308 30236
rect 7322 30184 7368 30236
rect 7368 30184 7374 30236
rect 7256 30114 7262 30166
rect 7262 30114 7308 30166
rect 7322 30114 7368 30166
rect 7368 30114 7374 30166
rect 7533 29930 7539 29982
rect 7539 29930 7585 29982
rect 7599 29930 7645 29982
rect 7645 29930 7651 29982
rect 7533 29861 7539 29913
rect 7539 29861 7585 29913
rect 7599 29861 7645 29913
rect 7645 29861 7651 29913
rect 7533 29792 7539 29844
rect 7539 29792 7585 29844
rect 7599 29792 7645 29844
rect 7645 29792 7651 29844
rect 7533 29723 7539 29775
rect 7539 29723 7585 29775
rect 7599 29723 7645 29775
rect 7645 29723 7651 29775
rect 7533 29654 7539 29706
rect 7539 29654 7585 29706
rect 7599 29654 7645 29706
rect 7645 29654 7651 29706
rect 7533 29584 7539 29636
rect 7539 29584 7585 29636
rect 7599 29584 7645 29636
rect 7645 29584 7651 29636
rect 7533 29514 7539 29566
rect 7539 29514 7585 29566
rect 7599 29514 7645 29566
rect 7645 29514 7651 29566
rect 7533 29444 7539 29496
rect 7539 29444 7585 29496
rect 7599 29444 7645 29496
rect 7645 29444 7651 29496
rect 7533 29380 7539 29426
rect 7539 29380 7585 29426
rect 7599 29380 7645 29426
rect 7645 29380 7651 29426
rect 7533 29374 7585 29380
rect 7599 29374 7651 29380
rect 7810 30714 7862 30720
rect 7810 30680 7816 30714
rect 7816 30680 7850 30714
rect 7850 30680 7862 30714
rect 7810 30668 7862 30680
rect 7876 30714 7928 30720
rect 7876 30680 7888 30714
rect 7888 30680 7922 30714
rect 7922 30680 7928 30714
rect 7876 30668 7928 30680
rect 7810 30641 7862 30651
rect 7810 30607 7816 30641
rect 7816 30607 7850 30641
rect 7850 30607 7862 30641
rect 7810 30599 7862 30607
rect 7876 30641 7928 30651
rect 7876 30607 7888 30641
rect 7888 30607 7922 30641
rect 7922 30607 7928 30641
rect 7876 30599 7928 30607
rect 7810 30568 7862 30582
rect 7810 30534 7816 30568
rect 7816 30534 7850 30568
rect 7850 30534 7862 30568
rect 7810 30530 7862 30534
rect 7876 30568 7928 30582
rect 7876 30534 7888 30568
rect 7888 30534 7922 30568
rect 7922 30534 7928 30568
rect 7876 30530 7928 30534
rect 7810 30495 7862 30513
rect 7810 30461 7816 30495
rect 7816 30461 7850 30495
rect 7850 30461 7862 30495
rect 7876 30495 7928 30513
rect 7876 30461 7888 30495
rect 7888 30461 7922 30495
rect 7922 30461 7928 30495
rect 7810 30422 7862 30444
rect 7876 30422 7928 30444
rect 7810 30392 7816 30422
rect 7816 30392 7862 30422
rect 7876 30392 7922 30422
rect 7922 30392 7928 30422
rect 7810 30323 7816 30375
rect 7816 30323 7862 30375
rect 7876 30323 7922 30375
rect 7922 30323 7928 30375
rect 7810 30254 7816 30306
rect 7816 30254 7862 30306
rect 7876 30254 7922 30306
rect 7922 30254 7928 30306
rect 7810 30184 7816 30236
rect 7816 30184 7862 30236
rect 7876 30184 7922 30236
rect 7922 30184 7928 30236
rect 7810 30114 7816 30166
rect 7816 30114 7862 30166
rect 7876 30114 7922 30166
rect 7922 30114 7928 30166
rect 8047 30693 8050 30724
rect 8050 30693 8084 30724
rect 8084 30693 8099 30724
rect 8047 30672 8099 30693
rect 8169 30717 8221 30724
rect 8169 30683 8184 30717
rect 8184 30683 8218 30717
rect 8218 30683 8221 30717
rect 8169 30672 8221 30683
rect 8047 30621 8050 30655
rect 8050 30621 8084 30655
rect 8084 30621 8099 30655
rect 8047 30603 8099 30621
rect 8169 30645 8221 30655
rect 8169 30611 8184 30645
rect 8184 30611 8218 30645
rect 8218 30611 8221 30645
rect 8169 30603 8221 30611
rect 8047 30583 8099 30586
rect 8047 30549 8050 30583
rect 8050 30549 8084 30583
rect 8084 30549 8099 30583
rect 8047 30534 8099 30549
rect 8169 30573 8221 30586
rect 8169 30539 8184 30573
rect 8184 30539 8218 30573
rect 8218 30539 8221 30573
rect 8169 30534 8221 30539
rect 8047 30511 8099 30517
rect 8047 30477 8050 30511
rect 8050 30477 8084 30511
rect 8084 30477 8099 30511
rect 8047 30465 8099 30477
rect 8169 30501 8221 30517
rect 8169 30467 8184 30501
rect 8184 30467 8218 30501
rect 8218 30467 8221 30501
rect 8169 30465 8221 30467
rect 8047 30439 8099 30448
rect 8047 30405 8050 30439
rect 8050 30405 8084 30439
rect 8084 30405 8099 30439
rect 8047 30396 8099 30405
rect 8169 30429 8221 30448
rect 8169 30396 8184 30429
rect 8184 30396 8218 30429
rect 8218 30396 8221 30429
rect 8047 30367 8099 30378
rect 8047 30333 8050 30367
rect 8050 30333 8084 30367
rect 8084 30333 8099 30367
rect 8047 30326 8099 30333
rect 8169 30357 8221 30378
rect 8169 30326 8184 30357
rect 8184 30326 8218 30357
rect 8218 30326 8221 30357
rect 8047 30295 8099 30308
rect 8047 30261 8050 30295
rect 8050 30261 8084 30295
rect 8084 30261 8099 30295
rect 8047 30256 8099 30261
rect 8169 30285 8221 30308
rect 8169 30256 8184 30285
rect 8184 30256 8218 30285
rect 8218 30256 8221 30285
rect 8047 30223 8099 30238
rect 8047 30189 8050 30223
rect 8050 30189 8084 30223
rect 8084 30189 8099 30223
rect 8047 30186 8099 30189
rect 8169 30213 8221 30238
rect 8169 30186 8184 30213
rect 8184 30186 8218 30213
rect 8218 30186 8221 30213
rect 8047 30151 8099 30168
rect 8047 30117 8050 30151
rect 8050 30117 8084 30151
rect 8084 30117 8099 30151
rect 8047 30116 8099 30117
rect 8169 30141 8221 30168
rect 8169 30116 8184 30141
rect 8184 30116 8218 30141
rect 8218 30116 8221 30141
rect 2270 28706 2276 28724
rect 2276 28706 2310 28724
rect 2310 28706 2322 28724
rect 2270 28672 2322 28706
rect 2392 28706 2410 28724
rect 2410 28706 2444 28724
rect 2392 28672 2444 28706
rect 2270 28634 2276 28655
rect 2276 28634 2310 28655
rect 2310 28634 2322 28655
rect 2270 28603 2322 28634
rect 2392 28634 2410 28655
rect 2410 28634 2444 28655
rect 2392 28603 2444 28634
rect 2270 28562 2276 28586
rect 2276 28562 2310 28586
rect 2310 28562 2322 28586
rect 2270 28534 2322 28562
rect 2392 28562 2410 28586
rect 2410 28562 2444 28586
rect 2392 28534 2444 28562
rect 2270 28490 2276 28517
rect 2276 28490 2310 28517
rect 2310 28490 2322 28517
rect 2270 28465 2322 28490
rect 2392 28490 2410 28517
rect 2410 28490 2444 28517
rect 2392 28465 2444 28490
rect 2270 28418 2276 28448
rect 2276 28418 2310 28448
rect 2310 28418 2322 28448
rect 2270 28396 2322 28418
rect 2392 28418 2410 28448
rect 2410 28418 2444 28448
rect 2392 28396 2444 28418
rect 2270 28346 2276 28378
rect 2276 28346 2310 28378
rect 2310 28346 2322 28378
rect 2270 28326 2322 28346
rect 2392 28346 2410 28378
rect 2410 28346 2444 28378
rect 2392 28326 2444 28346
rect 2270 28274 2276 28308
rect 2276 28274 2310 28308
rect 2310 28274 2322 28308
rect 2270 28256 2322 28274
rect 2392 28274 2410 28308
rect 2410 28274 2444 28308
rect 2392 28256 2444 28274
rect 2270 28236 2322 28238
rect 2270 28202 2276 28236
rect 2276 28202 2310 28236
rect 2310 28202 2322 28236
rect 2270 28186 2322 28202
rect 2392 28236 2444 28238
rect 2392 28202 2410 28236
rect 2410 28202 2444 28236
rect 2392 28186 2444 28202
rect 2270 28164 2322 28168
rect 2270 28130 2276 28164
rect 2276 28130 2310 28164
rect 2310 28130 2322 28164
rect 2270 28116 2322 28130
rect 2392 28164 2444 28168
rect 2392 28130 2410 28164
rect 2410 28130 2444 28164
rect 2392 28116 2444 28130
rect 2270 26690 2276 26724
rect 2276 26690 2310 26724
rect 2310 26690 2322 26724
rect 2270 26672 2322 26690
rect 2392 26690 2410 26724
rect 2410 26690 2444 26724
rect 2392 26672 2444 26690
rect 2270 26652 2322 26655
rect 2270 26618 2276 26652
rect 2276 26618 2310 26652
rect 2310 26618 2322 26652
rect 2270 26603 2322 26618
rect 2392 26652 2444 26655
rect 2392 26618 2410 26652
rect 2410 26618 2444 26652
rect 2392 26603 2444 26618
rect 2270 26580 2322 26586
rect 2270 26546 2276 26580
rect 2276 26546 2310 26580
rect 2310 26546 2322 26580
rect 2270 26534 2322 26546
rect 2392 26580 2444 26586
rect 2392 26546 2410 26580
rect 2410 26546 2444 26580
rect 2392 26534 2444 26546
rect 2270 26508 2322 26517
rect 2270 26474 2276 26508
rect 2276 26474 2310 26508
rect 2310 26474 2322 26508
rect 2270 26465 2322 26474
rect 2392 26508 2444 26517
rect 2392 26474 2410 26508
rect 2410 26474 2444 26508
rect 2392 26465 2444 26474
rect 2270 26436 2322 26448
rect 2270 26402 2276 26436
rect 2276 26402 2310 26436
rect 2310 26402 2322 26436
rect 2270 26396 2322 26402
rect 2392 26436 2444 26448
rect 2392 26402 2410 26436
rect 2410 26402 2444 26436
rect 2392 26396 2444 26402
rect 2270 26364 2322 26378
rect 2270 26330 2276 26364
rect 2276 26330 2310 26364
rect 2310 26330 2322 26364
rect 2270 26326 2322 26330
rect 2392 26364 2444 26378
rect 2392 26330 2410 26364
rect 2410 26330 2444 26364
rect 2392 26326 2444 26330
rect 2270 26292 2322 26308
rect 2270 26258 2276 26292
rect 2276 26258 2310 26292
rect 2310 26258 2322 26292
rect 2270 26256 2322 26258
rect 2392 26292 2444 26308
rect 2392 26258 2410 26292
rect 2410 26258 2444 26292
rect 2392 26256 2444 26258
rect 2270 26220 2322 26238
rect 2270 26186 2276 26220
rect 2276 26186 2310 26220
rect 2310 26186 2322 26220
rect 2392 26220 2444 26238
rect 2392 26186 2410 26220
rect 2410 26186 2444 26220
rect 2270 26148 2322 26168
rect 2270 26116 2276 26148
rect 2276 26116 2310 26148
rect 2310 26116 2322 26148
rect 2392 26148 2444 26168
rect 2392 26116 2410 26148
rect 2410 26116 2444 26148
rect 2270 24708 2322 24724
rect 2270 24674 2276 24708
rect 2276 24674 2310 24708
rect 2310 24674 2322 24708
rect 2270 24672 2322 24674
rect 2392 24708 2444 24724
rect 2392 24674 2410 24708
rect 2410 24674 2444 24708
rect 2392 24672 2444 24674
rect 2270 24636 2322 24655
rect 2270 24603 2276 24636
rect 2276 24603 2310 24636
rect 2310 24603 2322 24636
rect 2392 24636 2444 24655
rect 2392 24603 2410 24636
rect 2410 24603 2444 24636
rect 2270 24564 2322 24586
rect 2270 24534 2276 24564
rect 2276 24534 2310 24564
rect 2310 24534 2322 24564
rect 2392 24564 2444 24586
rect 2392 24534 2410 24564
rect 2410 24534 2444 24564
rect 2270 24492 2322 24517
rect 2270 24465 2276 24492
rect 2276 24465 2310 24492
rect 2310 24465 2322 24492
rect 2392 24492 2444 24517
rect 2392 24465 2410 24492
rect 2410 24465 2444 24492
rect 2270 24420 2322 24448
rect 2270 24396 2276 24420
rect 2276 24396 2310 24420
rect 2310 24396 2322 24420
rect 2392 24420 2444 24448
rect 2392 24396 2410 24420
rect 2410 24396 2444 24420
rect 2270 24348 2322 24378
rect 2270 24326 2276 24348
rect 2276 24326 2310 24348
rect 2310 24326 2322 24348
rect 2392 24348 2444 24378
rect 2392 24326 2410 24348
rect 2410 24326 2444 24348
rect 2270 24276 2322 24308
rect 2270 24256 2276 24276
rect 2276 24256 2310 24276
rect 2310 24256 2322 24276
rect 2392 24276 2444 24308
rect 2392 24256 2410 24276
rect 2410 24256 2444 24276
rect 2270 24204 2322 24238
rect 2270 24186 2276 24204
rect 2276 24186 2310 24204
rect 2310 24186 2322 24204
rect 2392 24204 2444 24238
rect 2392 24186 2410 24204
rect 2410 24186 2444 24204
rect 2270 24132 2322 24168
rect 2270 24116 2276 24132
rect 2276 24116 2310 24132
rect 2310 24116 2322 24132
rect 2392 24132 2444 24168
rect 2392 24116 2410 24132
rect 2410 24116 2444 24132
rect 2270 22692 2322 22724
rect 2270 22672 2276 22692
rect 2276 22672 2310 22692
rect 2310 22672 2322 22692
rect 2392 22692 2444 22724
rect 2392 22672 2410 22692
rect 2410 22672 2444 22692
rect 2270 22620 2322 22655
rect 2270 22603 2276 22620
rect 2276 22603 2310 22620
rect 2310 22603 2322 22620
rect 2392 22620 2444 22655
rect 2392 22603 2410 22620
rect 2410 22603 2444 22620
rect 2270 22548 2322 22586
rect 2270 22534 2276 22548
rect 2276 22534 2310 22548
rect 2310 22534 2322 22548
rect 2392 22548 2444 22586
rect 2392 22534 2410 22548
rect 2410 22534 2444 22548
rect 2270 22514 2276 22517
rect 2276 22514 2310 22517
rect 2310 22514 2322 22517
rect 2270 22476 2322 22514
rect 2270 22465 2276 22476
rect 2276 22465 2310 22476
rect 2310 22465 2322 22476
rect 2392 22514 2410 22517
rect 2410 22514 2444 22517
rect 2392 22476 2444 22514
rect 2392 22465 2410 22476
rect 2410 22465 2444 22476
rect 2270 22442 2276 22448
rect 2276 22442 2310 22448
rect 2310 22442 2322 22448
rect 2270 22404 2322 22442
rect 2270 22396 2276 22404
rect 2276 22396 2310 22404
rect 2310 22396 2322 22404
rect 2392 22442 2410 22448
rect 2410 22442 2444 22448
rect 2392 22404 2444 22442
rect 2392 22396 2410 22404
rect 2410 22396 2444 22404
rect 2270 22370 2276 22378
rect 2276 22370 2310 22378
rect 2310 22370 2322 22378
rect 2270 22332 2322 22370
rect 2270 22326 2276 22332
rect 2276 22326 2310 22332
rect 2310 22326 2322 22332
rect 2392 22370 2410 22378
rect 2410 22370 2444 22378
rect 2392 22332 2444 22370
rect 2392 22326 2410 22332
rect 2410 22326 2444 22332
rect 2270 22298 2276 22308
rect 2276 22298 2310 22308
rect 2310 22298 2322 22308
rect 2270 22260 2322 22298
rect 2270 22256 2276 22260
rect 2276 22256 2310 22260
rect 2310 22256 2322 22260
rect 2392 22298 2410 22308
rect 2410 22298 2444 22308
rect 2392 22260 2444 22298
rect 2392 22256 2410 22260
rect 2410 22256 2444 22260
rect 2270 22226 2276 22238
rect 2276 22226 2310 22238
rect 2310 22226 2322 22238
rect 2270 22188 2322 22226
rect 2270 22186 2276 22188
rect 2276 22186 2310 22188
rect 2310 22186 2322 22188
rect 2392 22226 2410 22238
rect 2410 22226 2444 22238
rect 2392 22188 2444 22226
rect 2392 22186 2410 22188
rect 2410 22186 2444 22188
rect 2270 22154 2276 22168
rect 2276 22154 2310 22168
rect 2310 22154 2322 22168
rect 2270 22116 2322 22154
rect 2392 22154 2410 22168
rect 2410 22154 2444 22168
rect 2392 22116 2444 22154
rect 2270 20714 2276 20724
rect 2276 20714 2310 20724
rect 2310 20714 2322 20724
rect 2270 20676 2322 20714
rect 2270 20672 2276 20676
rect 2276 20672 2310 20676
rect 2310 20672 2322 20676
rect 2392 20714 2410 20724
rect 2410 20714 2444 20724
rect 2392 20676 2444 20714
rect 2392 20672 2410 20676
rect 2410 20672 2444 20676
rect 2270 20642 2276 20655
rect 2276 20642 2310 20655
rect 2310 20642 2322 20655
rect 2270 20604 2322 20642
rect 2270 20603 2276 20604
rect 2276 20603 2310 20604
rect 2310 20603 2322 20604
rect 2392 20642 2410 20655
rect 2410 20642 2444 20655
rect 2392 20604 2444 20642
rect 2392 20603 2410 20604
rect 2410 20603 2444 20604
rect 2270 20570 2276 20586
rect 2276 20570 2310 20586
rect 2310 20570 2322 20586
rect 2270 20534 2322 20570
rect 2392 20570 2410 20586
rect 2410 20570 2444 20586
rect 2392 20534 2444 20570
rect 2270 20498 2276 20517
rect 2276 20498 2310 20517
rect 2310 20498 2322 20517
rect 2270 20465 2322 20498
rect 2392 20498 2410 20517
rect 2410 20498 2444 20517
rect 2392 20465 2444 20498
rect 2270 20426 2276 20448
rect 2276 20426 2310 20448
rect 2310 20426 2322 20448
rect 2270 20396 2322 20426
rect 2392 20426 2410 20448
rect 2410 20426 2444 20448
rect 2392 20396 2444 20426
rect 2270 20354 2276 20378
rect 2276 20354 2310 20378
rect 2310 20354 2322 20378
rect 2270 20326 2322 20354
rect 2392 20354 2410 20378
rect 2410 20354 2444 20378
rect 2392 20326 2444 20354
rect 2270 20282 2276 20308
rect 2276 20282 2310 20308
rect 2310 20282 2322 20308
rect 2270 20256 2322 20282
rect 2392 20282 2410 20308
rect 2410 20282 2444 20308
rect 2392 20256 2444 20282
rect 2270 20210 2276 20238
rect 2276 20210 2310 20238
rect 2310 20210 2322 20238
rect 2270 20186 2322 20210
rect 2392 20210 2410 20238
rect 2410 20210 2444 20238
rect 2392 20186 2444 20210
rect 2270 20138 2276 20168
rect 2276 20138 2310 20168
rect 2310 20138 2322 20168
rect 2270 20116 2322 20138
rect 2392 20138 2410 20168
rect 2410 20138 2444 20168
rect 2392 20116 2444 20138
rect 2270 18698 2276 18724
rect 2276 18698 2310 18724
rect 2310 18698 2322 18724
rect 2270 18672 2322 18698
rect 2392 18698 2410 18724
rect 2410 18698 2444 18724
rect 2392 18672 2444 18698
rect 2270 18626 2276 18655
rect 2276 18626 2310 18655
rect 2310 18626 2322 18655
rect 2270 18603 2322 18626
rect 2392 18626 2410 18655
rect 2410 18626 2444 18655
rect 2392 18603 2444 18626
rect 2270 18554 2276 18586
rect 2276 18554 2310 18586
rect 2310 18554 2322 18586
rect 2270 18534 2322 18554
rect 2392 18554 2410 18586
rect 2410 18554 2444 18586
rect 2392 18534 2444 18554
rect 2270 18516 2322 18517
rect 2270 18482 2276 18516
rect 2276 18482 2310 18516
rect 2310 18482 2322 18516
rect 2270 18465 2322 18482
rect 2392 18516 2444 18517
rect 2392 18482 2410 18516
rect 2410 18482 2444 18516
rect 2392 18465 2444 18482
rect 2270 18444 2322 18448
rect 2270 18410 2276 18444
rect 2276 18410 2310 18444
rect 2310 18410 2322 18444
rect 2270 18396 2322 18410
rect 2392 18444 2444 18448
rect 2392 18410 2410 18444
rect 2410 18410 2444 18444
rect 2392 18396 2444 18410
rect 2270 18372 2322 18378
rect 2270 18338 2276 18372
rect 2276 18338 2310 18372
rect 2310 18338 2322 18372
rect 2270 18326 2322 18338
rect 2392 18372 2444 18378
rect 2392 18338 2410 18372
rect 2410 18338 2444 18372
rect 2392 18326 2444 18338
rect 2270 18300 2322 18308
rect 2270 18266 2276 18300
rect 2276 18266 2310 18300
rect 2310 18266 2322 18300
rect 2270 18256 2322 18266
rect 2392 18300 2444 18308
rect 2392 18266 2410 18300
rect 2410 18266 2444 18300
rect 2392 18256 2444 18266
rect 2270 18228 2322 18238
rect 2270 18194 2276 18228
rect 2276 18194 2310 18228
rect 2310 18194 2322 18228
rect 2270 18186 2322 18194
rect 2392 18228 2444 18238
rect 2392 18194 2410 18228
rect 2410 18194 2444 18228
rect 2392 18186 2444 18194
rect 2270 18156 2322 18168
rect 2270 18122 2276 18156
rect 2276 18122 2310 18156
rect 2310 18122 2322 18156
rect 2270 18116 2322 18122
rect 2392 18156 2444 18168
rect 2392 18122 2410 18156
rect 2410 18122 2444 18156
rect 2392 18116 2444 18122
rect 2270 16970 2276 16973
rect 2276 16970 2310 16973
rect 2310 16970 2322 16973
rect 2270 16932 2322 16970
rect 2270 16921 2276 16932
rect 2276 16921 2310 16932
rect 2310 16921 2322 16932
rect 2392 16970 2410 16973
rect 2410 16970 2444 16973
rect 2392 16932 2444 16970
rect 2392 16921 2410 16932
rect 2410 16921 2444 16932
rect 2270 16898 2276 16907
rect 2276 16898 2310 16907
rect 2310 16898 2322 16907
rect 2270 16860 2322 16898
rect 2270 16855 2276 16860
rect 2276 16855 2310 16860
rect 2310 16855 2322 16860
rect 2392 16898 2410 16907
rect 2410 16898 2444 16907
rect 2392 16860 2444 16898
rect 2392 16855 2410 16860
rect 2410 16855 2444 16860
rect 2270 16826 2276 16841
rect 2276 16826 2310 16841
rect 2310 16826 2322 16841
rect 2270 16789 2322 16826
rect 2392 16826 2410 16841
rect 2410 16826 2444 16841
rect 2392 16789 2444 16826
rect 2270 16754 2276 16775
rect 2276 16754 2310 16775
rect 2310 16754 2322 16775
rect 2270 16723 2322 16754
rect 2392 16754 2410 16775
rect 2410 16754 2444 16775
rect 2392 16723 2444 16754
rect 2270 16682 2276 16709
rect 2276 16682 2310 16709
rect 2310 16682 2322 16709
rect 2270 16657 2322 16682
rect 2392 16682 2410 16709
rect 2410 16682 2444 16709
rect 2392 16657 2444 16682
rect 2270 16610 2276 16643
rect 2276 16610 2310 16643
rect 2310 16610 2322 16643
rect 2270 16591 2322 16610
rect 2392 16610 2410 16643
rect 2410 16610 2444 16643
rect 2392 16591 2444 16610
rect 2270 16572 2322 16577
rect 2270 16538 2276 16572
rect 2276 16538 2310 16572
rect 2310 16538 2322 16572
rect 2270 16525 2322 16538
rect 2392 16572 2444 16577
rect 2392 16538 2410 16572
rect 2410 16538 2444 16572
rect 2392 16525 2444 16538
rect 2270 16500 2322 16511
rect 2270 16466 2276 16500
rect 2276 16466 2310 16500
rect 2310 16466 2322 16500
rect 2270 16459 2322 16466
rect 2392 16500 2444 16511
rect 2392 16466 2410 16500
rect 2410 16466 2444 16500
rect 2392 16459 2444 16466
rect 2270 16428 2322 16445
rect 2270 16394 2276 16428
rect 2276 16394 2310 16428
rect 2310 16394 2322 16428
rect 2270 16393 2322 16394
rect 2392 16428 2444 16445
rect 2392 16394 2410 16428
rect 2410 16394 2444 16428
rect 2392 16393 2444 16394
rect 2270 16356 2322 16378
rect 2270 16326 2276 16356
rect 2276 16326 2310 16356
rect 2310 16326 2322 16356
rect 2392 16356 2444 16378
rect 2392 16326 2410 16356
rect 2410 16326 2444 16356
rect 2270 16284 2322 16311
rect 2270 16259 2276 16284
rect 2276 16259 2310 16284
rect 2310 16259 2322 16284
rect 2392 16284 2444 16311
rect 2392 16259 2410 16284
rect 2410 16259 2444 16284
rect 2270 16212 2322 16244
rect 2270 16192 2276 16212
rect 2276 16192 2310 16212
rect 2310 16192 2322 16212
rect 2392 16212 2444 16244
rect 2392 16192 2410 16212
rect 2410 16192 2444 16212
rect 2270 16140 2322 16177
rect 2270 16125 2276 16140
rect 2276 16125 2310 16140
rect 2310 16125 2322 16140
rect 2392 16140 2444 16177
rect 2392 16125 2410 16140
rect 2410 16125 2444 16140
rect 2270 16106 2276 16110
rect 2276 16106 2310 16110
rect 2310 16106 2322 16110
rect 2270 16068 2322 16106
rect 2270 16058 2276 16068
rect 2276 16058 2310 16068
rect 2310 16058 2322 16068
rect 2392 16106 2410 16110
rect 2410 16106 2444 16110
rect 2392 16068 2444 16106
rect 2392 16058 2410 16068
rect 2410 16058 2444 16068
rect 2270 16034 2276 16043
rect 2276 16034 2310 16043
rect 2310 16034 2322 16043
rect 2270 15996 2322 16034
rect 2270 15991 2276 15996
rect 2276 15991 2310 15996
rect 2310 15991 2322 15996
rect 2392 16034 2410 16043
rect 2410 16034 2444 16043
rect 2392 15996 2444 16034
rect 2392 15991 2410 15996
rect 2410 15991 2444 15996
rect 2648 26676 2663 26728
rect 2663 26676 2700 26728
rect 2713 26676 2765 26728
rect 2778 26676 2830 26728
rect 2843 26676 2895 26728
rect 2908 26676 2960 26728
rect 2973 26676 3025 26728
rect 3038 26676 3090 26728
rect 3103 26676 3155 26728
rect 3168 26676 3220 26728
rect 3233 26676 3285 26728
rect 3298 26676 3350 26728
rect 3363 26676 3415 26728
rect 3428 26676 3480 26728
rect 3493 26676 3545 26728
rect 3558 26676 3610 26728
rect 3623 26676 3675 26728
rect 3688 26676 3740 26728
rect 3753 26676 3805 26728
rect 3818 26676 3870 26728
rect 3883 26676 3935 26728
rect 3948 26676 4000 26728
rect 4013 26676 4065 26728
rect 4078 26676 4130 26728
rect 4143 26676 4195 26728
rect 4208 26676 4260 26728
rect 4273 26676 4325 26728
rect 4338 26676 4390 26728
rect 4403 26676 4455 26728
rect 4468 26676 4520 26728
rect 4532 26676 4569 26728
rect 4569 26676 4584 26728
rect 2648 26608 2663 26660
rect 2663 26608 2700 26660
rect 2713 26608 2765 26660
rect 2778 26608 2830 26660
rect 2843 26608 2895 26660
rect 2908 26608 2960 26660
rect 2973 26608 3025 26660
rect 3038 26608 3090 26660
rect 3103 26608 3155 26660
rect 3168 26608 3220 26660
rect 3233 26608 3285 26660
rect 3298 26608 3350 26660
rect 3363 26608 3415 26660
rect 3428 26608 3480 26660
rect 3493 26608 3545 26660
rect 3558 26608 3610 26660
rect 3623 26608 3675 26660
rect 3688 26608 3740 26660
rect 3753 26608 3805 26660
rect 3818 26608 3870 26660
rect 3883 26608 3935 26660
rect 3948 26608 4000 26660
rect 4013 26608 4065 26660
rect 4078 26608 4130 26660
rect 4143 26608 4195 26660
rect 4208 26608 4260 26660
rect 4273 26608 4325 26660
rect 4338 26608 4390 26660
rect 4403 26608 4455 26660
rect 4468 26608 4520 26660
rect 4532 26608 4569 26660
rect 4569 26608 4584 26660
rect 2648 26540 2663 26592
rect 2663 26540 2700 26592
rect 2713 26540 2765 26592
rect 2778 26540 2830 26592
rect 2843 26540 2895 26592
rect 2908 26540 2960 26592
rect 2973 26540 3025 26592
rect 3038 26540 3090 26592
rect 3103 26540 3155 26592
rect 3168 26540 3220 26592
rect 3233 26540 3285 26592
rect 3298 26540 3350 26592
rect 3363 26540 3415 26592
rect 3428 26540 3480 26592
rect 3493 26540 3545 26592
rect 3558 26540 3610 26592
rect 3623 26540 3675 26592
rect 3688 26540 3740 26592
rect 3753 26540 3805 26592
rect 3818 26540 3870 26592
rect 3883 26540 3935 26592
rect 3948 26540 4000 26592
rect 4013 26540 4065 26592
rect 4078 26540 4130 26592
rect 4143 26540 4195 26592
rect 4208 26540 4260 26592
rect 4273 26540 4325 26592
rect 4338 26540 4390 26592
rect 4403 26540 4455 26592
rect 4468 26540 4520 26592
rect 4532 26540 4569 26592
rect 4569 26540 4584 26592
rect 2648 26472 2663 26524
rect 2663 26472 2700 26524
rect 2713 26472 2765 26524
rect 2778 26472 2830 26524
rect 2843 26472 2895 26524
rect 2908 26472 2960 26524
rect 2973 26472 3025 26524
rect 3038 26472 3090 26524
rect 3103 26472 3155 26524
rect 3168 26472 3220 26524
rect 3233 26472 3285 26524
rect 3298 26472 3350 26524
rect 3363 26472 3415 26524
rect 3428 26472 3480 26524
rect 3493 26472 3545 26524
rect 3558 26472 3610 26524
rect 3623 26472 3675 26524
rect 3688 26472 3740 26524
rect 3753 26472 3805 26524
rect 3818 26472 3870 26524
rect 3883 26472 3935 26524
rect 3948 26472 4000 26524
rect 4013 26472 4065 26524
rect 4078 26472 4130 26524
rect 4143 26472 4195 26524
rect 4208 26472 4260 26524
rect 4273 26472 4325 26524
rect 4338 26472 4390 26524
rect 4403 26472 4455 26524
rect 4468 26472 4520 26524
rect 4532 26472 4569 26524
rect 4569 26472 4584 26524
rect 2648 26404 2663 26456
rect 2663 26404 2700 26456
rect 2713 26404 2765 26456
rect 2778 26404 2830 26456
rect 2843 26404 2895 26456
rect 2908 26404 2960 26456
rect 2973 26404 3025 26456
rect 3038 26404 3090 26456
rect 3103 26404 3155 26456
rect 3168 26404 3220 26456
rect 3233 26404 3285 26456
rect 3298 26404 3350 26456
rect 3363 26404 3415 26456
rect 3428 26404 3480 26456
rect 3493 26404 3545 26456
rect 3558 26404 3610 26456
rect 3623 26404 3675 26456
rect 3688 26404 3740 26456
rect 3753 26404 3805 26456
rect 3818 26404 3870 26456
rect 3883 26404 3935 26456
rect 3948 26404 4000 26456
rect 4013 26404 4065 26456
rect 4078 26404 4130 26456
rect 4143 26404 4195 26456
rect 4208 26404 4260 26456
rect 4273 26404 4325 26456
rect 4338 26404 4390 26456
rect 4403 26404 4455 26456
rect 4468 26404 4520 26456
rect 4532 26404 4569 26456
rect 4569 26404 4584 26456
rect 2648 26336 2663 26388
rect 2663 26336 2700 26388
rect 2713 26336 2765 26388
rect 2778 26336 2830 26388
rect 2843 26336 2895 26388
rect 2908 26336 2960 26388
rect 2973 26336 3025 26388
rect 3038 26336 3090 26388
rect 3103 26336 3155 26388
rect 3168 26336 3220 26388
rect 3233 26336 3285 26388
rect 3298 26336 3350 26388
rect 3363 26336 3415 26388
rect 3428 26336 3480 26388
rect 3493 26336 3545 26388
rect 3558 26336 3610 26388
rect 3623 26336 3675 26388
rect 3688 26336 3740 26388
rect 3753 26336 3805 26388
rect 3818 26336 3870 26388
rect 3883 26336 3935 26388
rect 3948 26336 4000 26388
rect 4013 26336 4065 26388
rect 4078 26336 4130 26388
rect 4143 26336 4195 26388
rect 4208 26336 4260 26388
rect 4273 26336 4325 26388
rect 4338 26336 4390 26388
rect 4403 26336 4455 26388
rect 4468 26336 4520 26388
rect 4532 26336 4569 26388
rect 4569 26336 4584 26388
rect 2648 26268 2663 26320
rect 2663 26268 2700 26320
rect 2713 26268 2765 26320
rect 2778 26268 2830 26320
rect 2843 26268 2895 26320
rect 2908 26268 2960 26320
rect 2973 26268 3025 26320
rect 3038 26268 3090 26320
rect 3103 26268 3155 26320
rect 3168 26268 3220 26320
rect 3233 26268 3285 26320
rect 3298 26268 3350 26320
rect 3363 26268 3415 26320
rect 3428 26268 3480 26320
rect 3493 26268 3545 26320
rect 3558 26268 3610 26320
rect 3623 26268 3675 26320
rect 3688 26268 3740 26320
rect 3753 26268 3805 26320
rect 3818 26268 3870 26320
rect 3883 26268 3935 26320
rect 3948 26268 4000 26320
rect 4013 26268 4065 26320
rect 4078 26268 4130 26320
rect 4143 26268 4195 26320
rect 4208 26268 4260 26320
rect 4273 26268 4325 26320
rect 4338 26268 4390 26320
rect 4403 26268 4455 26320
rect 4468 26268 4520 26320
rect 4532 26268 4569 26320
rect 4569 26268 4584 26320
rect 2648 26200 2663 26252
rect 2663 26200 2700 26252
rect 2713 26200 2765 26252
rect 2778 26200 2830 26252
rect 2843 26200 2895 26252
rect 2908 26200 2960 26252
rect 2973 26200 3025 26252
rect 3038 26200 3090 26252
rect 3103 26200 3155 26252
rect 3168 26200 3220 26252
rect 3233 26200 3285 26252
rect 3298 26200 3350 26252
rect 3363 26200 3415 26252
rect 3428 26200 3480 26252
rect 3493 26200 3545 26252
rect 3558 26200 3610 26252
rect 3623 26200 3675 26252
rect 3688 26200 3740 26252
rect 3753 26200 3805 26252
rect 3818 26200 3870 26252
rect 3883 26200 3935 26252
rect 3948 26200 4000 26252
rect 4013 26200 4065 26252
rect 4078 26200 4130 26252
rect 4143 26200 4195 26252
rect 4208 26200 4260 26252
rect 4273 26200 4325 26252
rect 4338 26200 4390 26252
rect 4403 26200 4455 26252
rect 4468 26200 4520 26252
rect 4532 26200 4569 26252
rect 4569 26200 4584 26252
rect 2648 24676 2663 24728
rect 2663 24676 2700 24728
rect 2713 24676 2765 24728
rect 2778 24676 2830 24728
rect 2843 24676 2895 24728
rect 2908 24676 2960 24728
rect 2973 24676 3025 24728
rect 3038 24676 3090 24728
rect 3103 24676 3155 24728
rect 3168 24676 3220 24728
rect 3233 24676 3285 24728
rect 3298 24676 3350 24728
rect 3363 24676 3415 24728
rect 3428 24676 3480 24728
rect 3493 24676 3545 24728
rect 3558 24676 3610 24728
rect 3623 24676 3675 24728
rect 3688 24676 3740 24728
rect 3753 24676 3805 24728
rect 3818 24676 3870 24728
rect 3883 24676 3935 24728
rect 3948 24676 4000 24728
rect 4013 24676 4065 24728
rect 4078 24676 4130 24728
rect 4143 24676 4195 24728
rect 4208 24676 4260 24728
rect 4273 24676 4325 24728
rect 4338 24676 4390 24728
rect 4403 24676 4455 24728
rect 4468 24676 4520 24728
rect 4532 24676 4569 24728
rect 4569 24676 4584 24728
rect 2648 24608 2663 24660
rect 2663 24608 2700 24660
rect 2713 24608 2765 24660
rect 2778 24608 2830 24660
rect 2843 24608 2895 24660
rect 2908 24608 2960 24660
rect 2973 24608 3025 24660
rect 3038 24608 3090 24660
rect 3103 24608 3155 24660
rect 3168 24608 3220 24660
rect 3233 24608 3285 24660
rect 3298 24608 3350 24660
rect 3363 24608 3415 24660
rect 3428 24608 3480 24660
rect 3493 24608 3545 24660
rect 3558 24608 3610 24660
rect 3623 24608 3675 24660
rect 3688 24608 3740 24660
rect 3753 24608 3805 24660
rect 3818 24608 3870 24660
rect 3883 24608 3935 24660
rect 3948 24608 4000 24660
rect 4013 24608 4065 24660
rect 4078 24608 4130 24660
rect 4143 24608 4195 24660
rect 4208 24608 4260 24660
rect 4273 24608 4325 24660
rect 4338 24608 4390 24660
rect 4403 24608 4455 24660
rect 4468 24608 4520 24660
rect 4532 24608 4569 24660
rect 4569 24608 4584 24660
rect 2648 24540 2663 24592
rect 2663 24540 2700 24592
rect 2713 24540 2765 24592
rect 2778 24540 2830 24592
rect 2843 24540 2895 24592
rect 2908 24540 2960 24592
rect 2973 24540 3025 24592
rect 3038 24540 3090 24592
rect 3103 24540 3155 24592
rect 3168 24540 3220 24592
rect 3233 24540 3285 24592
rect 3298 24540 3350 24592
rect 3363 24540 3415 24592
rect 3428 24540 3480 24592
rect 3493 24540 3545 24592
rect 3558 24540 3610 24592
rect 3623 24540 3675 24592
rect 3688 24540 3740 24592
rect 3753 24540 3805 24592
rect 3818 24540 3870 24592
rect 3883 24540 3935 24592
rect 3948 24540 4000 24592
rect 4013 24540 4065 24592
rect 4078 24540 4130 24592
rect 4143 24540 4195 24592
rect 4208 24540 4260 24592
rect 4273 24540 4325 24592
rect 4338 24540 4390 24592
rect 4403 24540 4455 24592
rect 4468 24540 4520 24592
rect 4532 24540 4569 24592
rect 4569 24540 4584 24592
rect 2648 24472 2663 24524
rect 2663 24472 2700 24524
rect 2713 24472 2765 24524
rect 2778 24472 2830 24524
rect 2843 24472 2895 24524
rect 2908 24472 2960 24524
rect 2973 24472 3025 24524
rect 3038 24472 3090 24524
rect 3103 24472 3155 24524
rect 3168 24472 3220 24524
rect 3233 24472 3285 24524
rect 3298 24472 3350 24524
rect 3363 24472 3415 24524
rect 3428 24472 3480 24524
rect 3493 24472 3545 24524
rect 3558 24472 3610 24524
rect 3623 24472 3675 24524
rect 3688 24472 3740 24524
rect 3753 24472 3805 24524
rect 3818 24472 3870 24524
rect 3883 24472 3935 24524
rect 3948 24472 4000 24524
rect 4013 24472 4065 24524
rect 4078 24472 4130 24524
rect 4143 24472 4195 24524
rect 4208 24472 4260 24524
rect 4273 24472 4325 24524
rect 4338 24472 4390 24524
rect 4403 24472 4455 24524
rect 4468 24472 4520 24524
rect 4532 24472 4569 24524
rect 4569 24472 4584 24524
rect 2648 24404 2663 24456
rect 2663 24404 2700 24456
rect 2713 24404 2765 24456
rect 2778 24404 2830 24456
rect 2843 24404 2895 24456
rect 2908 24404 2960 24456
rect 2973 24404 3025 24456
rect 3038 24404 3090 24456
rect 3103 24404 3155 24456
rect 3168 24404 3220 24456
rect 3233 24404 3285 24456
rect 3298 24404 3350 24456
rect 3363 24404 3415 24456
rect 3428 24404 3480 24456
rect 3493 24404 3545 24456
rect 3558 24404 3610 24456
rect 3623 24404 3675 24456
rect 3688 24404 3740 24456
rect 3753 24404 3805 24456
rect 3818 24404 3870 24456
rect 3883 24404 3935 24456
rect 3948 24404 4000 24456
rect 4013 24404 4065 24456
rect 4078 24404 4130 24456
rect 4143 24404 4195 24456
rect 4208 24404 4260 24456
rect 4273 24404 4325 24456
rect 4338 24404 4390 24456
rect 4403 24404 4455 24456
rect 4468 24404 4520 24456
rect 4532 24404 4569 24456
rect 4569 24404 4584 24456
rect 2648 24336 2663 24388
rect 2663 24336 2700 24388
rect 2713 24336 2765 24388
rect 2778 24336 2830 24388
rect 2843 24336 2895 24388
rect 2908 24336 2960 24388
rect 2973 24336 3025 24388
rect 3038 24336 3090 24388
rect 3103 24336 3155 24388
rect 3168 24336 3220 24388
rect 3233 24336 3285 24388
rect 3298 24336 3350 24388
rect 3363 24336 3415 24388
rect 3428 24336 3480 24388
rect 3493 24336 3545 24388
rect 3558 24336 3610 24388
rect 3623 24336 3675 24388
rect 3688 24336 3740 24388
rect 3753 24336 3805 24388
rect 3818 24336 3870 24388
rect 3883 24336 3935 24388
rect 3948 24336 4000 24388
rect 4013 24336 4065 24388
rect 4078 24336 4130 24388
rect 4143 24336 4195 24388
rect 4208 24336 4260 24388
rect 4273 24336 4325 24388
rect 4338 24336 4390 24388
rect 4403 24336 4455 24388
rect 4468 24336 4520 24388
rect 4532 24336 4569 24388
rect 4569 24336 4584 24388
rect 2648 24268 2663 24320
rect 2663 24268 2700 24320
rect 2713 24268 2765 24320
rect 2778 24268 2830 24320
rect 2843 24268 2895 24320
rect 2908 24268 2960 24320
rect 2973 24268 3025 24320
rect 3038 24268 3090 24320
rect 3103 24268 3155 24320
rect 3168 24268 3220 24320
rect 3233 24268 3285 24320
rect 3298 24268 3350 24320
rect 3363 24268 3415 24320
rect 3428 24268 3480 24320
rect 3493 24268 3545 24320
rect 3558 24268 3610 24320
rect 3623 24268 3675 24320
rect 3688 24268 3740 24320
rect 3753 24268 3805 24320
rect 3818 24268 3870 24320
rect 3883 24268 3935 24320
rect 3948 24268 4000 24320
rect 4013 24268 4065 24320
rect 4078 24268 4130 24320
rect 4143 24268 4195 24320
rect 4208 24268 4260 24320
rect 4273 24268 4325 24320
rect 4338 24268 4390 24320
rect 4403 24268 4455 24320
rect 4468 24268 4520 24320
rect 4532 24268 4569 24320
rect 4569 24268 4584 24320
rect 2648 24200 2663 24252
rect 2663 24200 2700 24252
rect 2713 24200 2765 24252
rect 2778 24200 2830 24252
rect 2843 24200 2895 24252
rect 2908 24200 2960 24252
rect 2973 24200 3025 24252
rect 3038 24200 3090 24252
rect 3103 24200 3155 24252
rect 3168 24200 3220 24252
rect 3233 24200 3285 24252
rect 3298 24200 3350 24252
rect 3363 24200 3415 24252
rect 3428 24200 3480 24252
rect 3493 24200 3545 24252
rect 3558 24200 3610 24252
rect 3623 24200 3675 24252
rect 3688 24200 3740 24252
rect 3753 24200 3805 24252
rect 3818 24200 3870 24252
rect 3883 24200 3935 24252
rect 3948 24200 4000 24252
rect 4013 24200 4065 24252
rect 4078 24200 4130 24252
rect 4143 24200 4195 24252
rect 4208 24200 4260 24252
rect 4273 24200 4325 24252
rect 4338 24200 4390 24252
rect 4403 24200 4455 24252
rect 4468 24200 4520 24252
rect 4532 24200 4569 24252
rect 4569 24200 4584 24252
rect 2648 22676 2663 22728
rect 2663 22676 2700 22728
rect 2713 22676 2765 22728
rect 2778 22676 2830 22728
rect 2843 22676 2895 22728
rect 2908 22676 2960 22728
rect 2973 22676 3025 22728
rect 3038 22676 3090 22728
rect 3103 22676 3155 22728
rect 3168 22676 3220 22728
rect 3233 22676 3285 22728
rect 3298 22676 3350 22728
rect 3363 22676 3415 22728
rect 3428 22676 3480 22728
rect 3493 22676 3545 22728
rect 3558 22676 3610 22728
rect 3623 22676 3675 22728
rect 3688 22676 3740 22728
rect 3753 22676 3805 22728
rect 3818 22676 3870 22728
rect 3883 22676 3935 22728
rect 3948 22676 4000 22728
rect 4013 22676 4065 22728
rect 4078 22676 4130 22728
rect 4143 22676 4195 22728
rect 4208 22676 4260 22728
rect 4273 22676 4325 22728
rect 4338 22676 4390 22728
rect 4403 22676 4455 22728
rect 4468 22676 4520 22728
rect 4532 22676 4569 22728
rect 4569 22676 4584 22728
rect 2648 22608 2663 22660
rect 2663 22608 2700 22660
rect 2713 22608 2765 22660
rect 2778 22608 2830 22660
rect 2843 22608 2895 22660
rect 2908 22608 2960 22660
rect 2973 22608 3025 22660
rect 3038 22608 3090 22660
rect 3103 22608 3155 22660
rect 3168 22608 3220 22660
rect 3233 22608 3285 22660
rect 3298 22608 3350 22660
rect 3363 22608 3415 22660
rect 3428 22608 3480 22660
rect 3493 22608 3545 22660
rect 3558 22608 3610 22660
rect 3623 22608 3675 22660
rect 3688 22608 3740 22660
rect 3753 22608 3805 22660
rect 3818 22608 3870 22660
rect 3883 22608 3935 22660
rect 3948 22608 4000 22660
rect 4013 22608 4065 22660
rect 4078 22608 4130 22660
rect 4143 22608 4195 22660
rect 4208 22608 4260 22660
rect 4273 22608 4325 22660
rect 4338 22608 4390 22660
rect 4403 22608 4455 22660
rect 4468 22608 4520 22660
rect 4532 22608 4569 22660
rect 4569 22608 4584 22660
rect 2648 22540 2663 22592
rect 2663 22540 2700 22592
rect 2713 22540 2765 22592
rect 2778 22540 2830 22592
rect 2843 22540 2895 22592
rect 2908 22540 2960 22592
rect 2973 22540 3025 22592
rect 3038 22540 3090 22592
rect 3103 22540 3155 22592
rect 3168 22540 3220 22592
rect 3233 22540 3285 22592
rect 3298 22540 3350 22592
rect 3363 22540 3415 22592
rect 3428 22540 3480 22592
rect 3493 22540 3545 22592
rect 3558 22540 3610 22592
rect 3623 22540 3675 22592
rect 3688 22540 3740 22592
rect 3753 22540 3805 22592
rect 3818 22540 3870 22592
rect 3883 22540 3935 22592
rect 3948 22540 4000 22592
rect 4013 22540 4065 22592
rect 4078 22540 4130 22592
rect 4143 22540 4195 22592
rect 4208 22540 4260 22592
rect 4273 22540 4325 22592
rect 4338 22540 4390 22592
rect 4403 22540 4455 22592
rect 4468 22540 4520 22592
rect 4532 22540 4569 22592
rect 4569 22540 4584 22592
rect 2648 22472 2663 22524
rect 2663 22472 2700 22524
rect 2713 22472 2765 22524
rect 2778 22472 2830 22524
rect 2843 22472 2895 22524
rect 2908 22472 2960 22524
rect 2973 22472 3025 22524
rect 3038 22472 3090 22524
rect 3103 22472 3155 22524
rect 3168 22472 3220 22524
rect 3233 22472 3285 22524
rect 3298 22472 3350 22524
rect 3363 22472 3415 22524
rect 3428 22472 3480 22524
rect 3493 22472 3545 22524
rect 3558 22472 3610 22524
rect 3623 22472 3675 22524
rect 3688 22472 3740 22524
rect 3753 22472 3805 22524
rect 3818 22472 3870 22524
rect 3883 22472 3935 22524
rect 3948 22472 4000 22524
rect 4013 22472 4065 22524
rect 4078 22472 4130 22524
rect 4143 22472 4195 22524
rect 4208 22472 4260 22524
rect 4273 22472 4325 22524
rect 4338 22472 4390 22524
rect 4403 22472 4455 22524
rect 4468 22472 4520 22524
rect 4532 22472 4569 22524
rect 4569 22472 4584 22524
rect 2648 22404 2663 22456
rect 2663 22404 2700 22456
rect 2713 22404 2765 22456
rect 2778 22404 2830 22456
rect 2843 22404 2895 22456
rect 2908 22404 2960 22456
rect 2973 22404 3025 22456
rect 3038 22404 3090 22456
rect 3103 22404 3155 22456
rect 3168 22404 3220 22456
rect 3233 22404 3285 22456
rect 3298 22404 3350 22456
rect 3363 22404 3415 22456
rect 3428 22404 3480 22456
rect 3493 22404 3545 22456
rect 3558 22404 3610 22456
rect 3623 22404 3675 22456
rect 3688 22404 3740 22456
rect 3753 22404 3805 22456
rect 3818 22404 3870 22456
rect 3883 22404 3935 22456
rect 3948 22404 4000 22456
rect 4013 22404 4065 22456
rect 4078 22404 4130 22456
rect 4143 22404 4195 22456
rect 4208 22404 4260 22456
rect 4273 22404 4325 22456
rect 4338 22404 4390 22456
rect 4403 22404 4455 22456
rect 4468 22404 4520 22456
rect 4532 22404 4569 22456
rect 4569 22404 4584 22456
rect 2648 22336 2663 22388
rect 2663 22336 2700 22388
rect 2713 22336 2765 22388
rect 2778 22336 2830 22388
rect 2843 22336 2895 22388
rect 2908 22336 2960 22388
rect 2973 22336 3025 22388
rect 3038 22336 3090 22388
rect 3103 22336 3155 22388
rect 3168 22336 3220 22388
rect 3233 22336 3285 22388
rect 3298 22336 3350 22388
rect 3363 22336 3415 22388
rect 3428 22336 3480 22388
rect 3493 22336 3545 22388
rect 3558 22336 3610 22388
rect 3623 22336 3675 22388
rect 3688 22336 3740 22388
rect 3753 22336 3805 22388
rect 3818 22336 3870 22388
rect 3883 22336 3935 22388
rect 3948 22336 4000 22388
rect 4013 22336 4065 22388
rect 4078 22336 4130 22388
rect 4143 22336 4195 22388
rect 4208 22336 4260 22388
rect 4273 22336 4325 22388
rect 4338 22336 4390 22388
rect 4403 22336 4455 22388
rect 4468 22336 4520 22388
rect 4532 22336 4569 22388
rect 4569 22336 4584 22388
rect 2648 22268 2663 22320
rect 2663 22268 2700 22320
rect 2713 22268 2765 22320
rect 2778 22268 2830 22320
rect 2843 22268 2895 22320
rect 2908 22268 2960 22320
rect 2973 22268 3025 22320
rect 3038 22268 3090 22320
rect 3103 22268 3155 22320
rect 3168 22268 3220 22320
rect 3233 22268 3285 22320
rect 3298 22268 3350 22320
rect 3363 22268 3415 22320
rect 3428 22268 3480 22320
rect 3493 22268 3545 22320
rect 3558 22268 3610 22320
rect 3623 22268 3675 22320
rect 3688 22268 3740 22320
rect 3753 22268 3805 22320
rect 3818 22268 3870 22320
rect 3883 22268 3935 22320
rect 3948 22268 4000 22320
rect 4013 22268 4065 22320
rect 4078 22268 4130 22320
rect 4143 22268 4195 22320
rect 4208 22268 4260 22320
rect 4273 22268 4325 22320
rect 4338 22268 4390 22320
rect 4403 22268 4455 22320
rect 4468 22268 4520 22320
rect 4532 22268 4569 22320
rect 4569 22268 4584 22320
rect 2648 22200 2663 22252
rect 2663 22200 2700 22252
rect 2713 22200 2765 22252
rect 2778 22200 2830 22252
rect 2843 22200 2895 22252
rect 2908 22200 2960 22252
rect 2973 22200 3025 22252
rect 3038 22200 3090 22252
rect 3103 22200 3155 22252
rect 3168 22200 3220 22252
rect 3233 22200 3285 22252
rect 3298 22200 3350 22252
rect 3363 22200 3415 22252
rect 3428 22200 3480 22252
rect 3493 22200 3545 22252
rect 3558 22200 3610 22252
rect 3623 22200 3675 22252
rect 3688 22200 3740 22252
rect 3753 22200 3805 22252
rect 3818 22200 3870 22252
rect 3883 22200 3935 22252
rect 3948 22200 4000 22252
rect 4013 22200 4065 22252
rect 4078 22200 4130 22252
rect 4143 22200 4195 22252
rect 4208 22200 4260 22252
rect 4273 22200 4325 22252
rect 4338 22200 4390 22252
rect 4403 22200 4455 22252
rect 4468 22200 4520 22252
rect 4532 22200 4569 22252
rect 4569 22200 4584 22252
rect 2648 20676 2663 20728
rect 2663 20676 2700 20728
rect 2713 20676 2765 20728
rect 2778 20676 2830 20728
rect 2843 20676 2895 20728
rect 2908 20676 2960 20728
rect 2973 20676 3025 20728
rect 3038 20676 3090 20728
rect 3103 20676 3155 20728
rect 3168 20676 3220 20728
rect 3233 20676 3285 20728
rect 3298 20676 3350 20728
rect 3363 20676 3415 20728
rect 3428 20676 3480 20728
rect 3493 20676 3545 20728
rect 3558 20676 3610 20728
rect 3623 20676 3675 20728
rect 3688 20676 3740 20728
rect 3753 20676 3805 20728
rect 3818 20676 3870 20728
rect 3883 20676 3935 20728
rect 3948 20676 4000 20728
rect 4013 20676 4065 20728
rect 4078 20676 4130 20728
rect 4143 20676 4195 20728
rect 4208 20676 4260 20728
rect 4273 20676 4325 20728
rect 4338 20676 4390 20728
rect 4403 20676 4455 20728
rect 4468 20676 4520 20728
rect 4532 20676 4569 20728
rect 4569 20676 4584 20728
rect 2648 20608 2663 20660
rect 2663 20608 2700 20660
rect 2713 20608 2765 20660
rect 2778 20608 2830 20660
rect 2843 20608 2895 20660
rect 2908 20608 2960 20660
rect 2973 20608 3025 20660
rect 3038 20608 3090 20660
rect 3103 20608 3155 20660
rect 3168 20608 3220 20660
rect 3233 20608 3285 20660
rect 3298 20608 3350 20660
rect 3363 20608 3415 20660
rect 3428 20608 3480 20660
rect 3493 20608 3545 20660
rect 3558 20608 3610 20660
rect 3623 20608 3675 20660
rect 3688 20608 3740 20660
rect 3753 20608 3805 20660
rect 3818 20608 3870 20660
rect 3883 20608 3935 20660
rect 3948 20608 4000 20660
rect 4013 20608 4065 20660
rect 4078 20608 4130 20660
rect 4143 20608 4195 20660
rect 4208 20608 4260 20660
rect 4273 20608 4325 20660
rect 4338 20608 4390 20660
rect 4403 20608 4455 20660
rect 4468 20608 4520 20660
rect 4532 20608 4569 20660
rect 4569 20608 4584 20660
rect 2648 20540 2663 20592
rect 2663 20540 2700 20592
rect 2713 20540 2765 20592
rect 2778 20540 2830 20592
rect 2843 20540 2895 20592
rect 2908 20540 2960 20592
rect 2973 20540 3025 20592
rect 3038 20540 3090 20592
rect 3103 20540 3155 20592
rect 3168 20540 3220 20592
rect 3233 20540 3285 20592
rect 3298 20540 3350 20592
rect 3363 20540 3415 20592
rect 3428 20540 3480 20592
rect 3493 20540 3545 20592
rect 3558 20540 3610 20592
rect 3623 20540 3675 20592
rect 3688 20540 3740 20592
rect 3753 20540 3805 20592
rect 3818 20540 3870 20592
rect 3883 20540 3935 20592
rect 3948 20540 4000 20592
rect 4013 20540 4065 20592
rect 4078 20540 4130 20592
rect 4143 20540 4195 20592
rect 4208 20540 4260 20592
rect 4273 20540 4325 20592
rect 4338 20540 4390 20592
rect 4403 20540 4455 20592
rect 4468 20540 4520 20592
rect 4532 20540 4569 20592
rect 4569 20540 4584 20592
rect 2648 20472 2663 20524
rect 2663 20472 2700 20524
rect 2713 20472 2765 20524
rect 2778 20472 2830 20524
rect 2843 20472 2895 20524
rect 2908 20472 2960 20524
rect 2973 20472 3025 20524
rect 3038 20472 3090 20524
rect 3103 20472 3155 20524
rect 3168 20472 3220 20524
rect 3233 20472 3285 20524
rect 3298 20472 3350 20524
rect 3363 20472 3415 20524
rect 3428 20472 3480 20524
rect 3493 20472 3545 20524
rect 3558 20472 3610 20524
rect 3623 20472 3675 20524
rect 3688 20472 3740 20524
rect 3753 20472 3805 20524
rect 3818 20472 3870 20524
rect 3883 20472 3935 20524
rect 3948 20472 4000 20524
rect 4013 20472 4065 20524
rect 4078 20472 4130 20524
rect 4143 20472 4195 20524
rect 4208 20472 4260 20524
rect 4273 20472 4325 20524
rect 4338 20472 4390 20524
rect 4403 20472 4455 20524
rect 4468 20472 4520 20524
rect 4532 20472 4569 20524
rect 4569 20472 4584 20524
rect 2648 20404 2663 20456
rect 2663 20404 2700 20456
rect 2713 20404 2765 20456
rect 2778 20404 2830 20456
rect 2843 20404 2895 20456
rect 2908 20404 2960 20456
rect 2973 20404 3025 20456
rect 3038 20404 3090 20456
rect 3103 20404 3155 20456
rect 3168 20404 3220 20456
rect 3233 20404 3285 20456
rect 3298 20404 3350 20456
rect 3363 20404 3415 20456
rect 3428 20404 3480 20456
rect 3493 20404 3545 20456
rect 3558 20404 3610 20456
rect 3623 20404 3675 20456
rect 3688 20404 3740 20456
rect 3753 20404 3805 20456
rect 3818 20404 3870 20456
rect 3883 20404 3935 20456
rect 3948 20404 4000 20456
rect 4013 20404 4065 20456
rect 4078 20404 4130 20456
rect 4143 20404 4195 20456
rect 4208 20404 4260 20456
rect 4273 20404 4325 20456
rect 4338 20404 4390 20456
rect 4403 20404 4455 20456
rect 4468 20404 4520 20456
rect 4532 20404 4569 20456
rect 4569 20404 4584 20456
rect 2648 20336 2663 20388
rect 2663 20336 2700 20388
rect 2713 20336 2765 20388
rect 2778 20336 2830 20388
rect 2843 20336 2895 20388
rect 2908 20336 2960 20388
rect 2973 20336 3025 20388
rect 3038 20336 3090 20388
rect 3103 20336 3155 20388
rect 3168 20336 3220 20388
rect 3233 20336 3285 20388
rect 3298 20336 3350 20388
rect 3363 20336 3415 20388
rect 3428 20336 3480 20388
rect 3493 20336 3545 20388
rect 3558 20336 3610 20388
rect 3623 20336 3675 20388
rect 3688 20336 3740 20388
rect 3753 20336 3805 20388
rect 3818 20336 3870 20388
rect 3883 20336 3935 20388
rect 3948 20336 4000 20388
rect 4013 20336 4065 20388
rect 4078 20336 4130 20388
rect 4143 20336 4195 20388
rect 4208 20336 4260 20388
rect 4273 20336 4325 20388
rect 4338 20336 4390 20388
rect 4403 20336 4455 20388
rect 4468 20336 4520 20388
rect 4532 20336 4569 20388
rect 4569 20336 4584 20388
rect 2648 20268 2663 20320
rect 2663 20268 2700 20320
rect 2713 20268 2765 20320
rect 2778 20268 2830 20320
rect 2843 20268 2895 20320
rect 2908 20268 2960 20320
rect 2973 20268 3025 20320
rect 3038 20268 3090 20320
rect 3103 20268 3155 20320
rect 3168 20268 3220 20320
rect 3233 20268 3285 20320
rect 3298 20268 3350 20320
rect 3363 20268 3415 20320
rect 3428 20268 3480 20320
rect 3493 20268 3545 20320
rect 3558 20268 3610 20320
rect 3623 20268 3675 20320
rect 3688 20268 3740 20320
rect 3753 20268 3805 20320
rect 3818 20268 3870 20320
rect 3883 20268 3935 20320
rect 3948 20268 4000 20320
rect 4013 20268 4065 20320
rect 4078 20268 4130 20320
rect 4143 20268 4195 20320
rect 4208 20268 4260 20320
rect 4273 20268 4325 20320
rect 4338 20268 4390 20320
rect 4403 20268 4455 20320
rect 4468 20268 4520 20320
rect 4532 20268 4569 20320
rect 4569 20268 4584 20320
rect 2648 20200 2663 20252
rect 2663 20200 2700 20252
rect 2713 20200 2765 20252
rect 2778 20200 2830 20252
rect 2843 20200 2895 20252
rect 2908 20200 2960 20252
rect 2973 20200 3025 20252
rect 3038 20200 3090 20252
rect 3103 20200 3155 20252
rect 3168 20200 3220 20252
rect 3233 20200 3285 20252
rect 3298 20200 3350 20252
rect 3363 20200 3415 20252
rect 3428 20200 3480 20252
rect 3493 20200 3545 20252
rect 3558 20200 3610 20252
rect 3623 20200 3675 20252
rect 3688 20200 3740 20252
rect 3753 20200 3805 20252
rect 3818 20200 3870 20252
rect 3883 20200 3935 20252
rect 3948 20200 4000 20252
rect 4013 20200 4065 20252
rect 4078 20200 4130 20252
rect 4143 20200 4195 20252
rect 4208 20200 4260 20252
rect 4273 20200 4325 20252
rect 4338 20200 4390 20252
rect 4403 20200 4455 20252
rect 4468 20200 4520 20252
rect 4532 20200 4569 20252
rect 4569 20200 4584 20252
rect 2648 18676 2663 18728
rect 2663 18676 2700 18728
rect 2713 18676 2765 18728
rect 2778 18676 2830 18728
rect 2843 18676 2895 18728
rect 2908 18676 2960 18728
rect 2973 18676 3025 18728
rect 3038 18676 3090 18728
rect 3103 18676 3155 18728
rect 3168 18676 3220 18728
rect 3233 18676 3285 18728
rect 3298 18676 3350 18728
rect 3363 18676 3415 18728
rect 3428 18676 3480 18728
rect 3493 18676 3545 18728
rect 3558 18676 3610 18728
rect 3623 18676 3675 18728
rect 3688 18676 3740 18728
rect 3753 18676 3805 18728
rect 3818 18676 3870 18728
rect 3883 18676 3935 18728
rect 3948 18676 4000 18728
rect 4013 18676 4065 18728
rect 4078 18676 4130 18728
rect 4143 18676 4195 18728
rect 4208 18676 4260 18728
rect 4273 18676 4325 18728
rect 4338 18676 4390 18728
rect 4403 18676 4455 18728
rect 4468 18676 4520 18728
rect 4532 18676 4569 18728
rect 4569 18676 4584 18728
rect 2648 18608 2663 18660
rect 2663 18608 2700 18660
rect 2713 18608 2765 18660
rect 2778 18608 2830 18660
rect 2843 18608 2895 18660
rect 2908 18608 2960 18660
rect 2973 18608 3025 18660
rect 3038 18608 3090 18660
rect 3103 18608 3155 18660
rect 3168 18608 3220 18660
rect 3233 18608 3285 18660
rect 3298 18608 3350 18660
rect 3363 18608 3415 18660
rect 3428 18608 3480 18660
rect 3493 18608 3545 18660
rect 3558 18608 3610 18660
rect 3623 18608 3675 18660
rect 3688 18608 3740 18660
rect 3753 18608 3805 18660
rect 3818 18608 3870 18660
rect 3883 18608 3935 18660
rect 3948 18608 4000 18660
rect 4013 18608 4065 18660
rect 4078 18608 4130 18660
rect 4143 18608 4195 18660
rect 4208 18608 4260 18660
rect 4273 18608 4325 18660
rect 4338 18608 4390 18660
rect 4403 18608 4455 18660
rect 4468 18608 4520 18660
rect 4532 18608 4569 18660
rect 4569 18608 4584 18660
rect 2648 18563 2663 18592
rect 2663 18563 2700 18592
rect 2713 18563 2765 18592
rect 2778 18563 2830 18592
rect 2843 18563 2895 18592
rect 2908 18563 2960 18592
rect 2973 18563 3025 18592
rect 3038 18563 3090 18592
rect 3103 18563 3155 18592
rect 3168 18563 3220 18592
rect 3233 18563 3285 18592
rect 3298 18563 3350 18592
rect 3363 18563 3415 18592
rect 3428 18563 3480 18592
rect 3493 18563 3545 18592
rect 3558 18563 3610 18592
rect 3623 18563 3675 18592
rect 3688 18563 3740 18592
rect 3753 18563 3805 18592
rect 3818 18563 3870 18592
rect 3883 18563 3935 18592
rect 3948 18563 4000 18592
rect 4013 18563 4065 18592
rect 4078 18563 4130 18592
rect 4143 18563 4195 18592
rect 4208 18563 4260 18592
rect 4273 18563 4325 18592
rect 4338 18563 4390 18592
rect 4403 18563 4455 18592
rect 4468 18563 4520 18592
rect 4532 18563 4569 18592
rect 4569 18563 4584 18592
rect 2648 18540 2700 18563
rect 2713 18540 2765 18563
rect 2778 18540 2830 18563
rect 2843 18540 2895 18563
rect 2908 18540 2960 18563
rect 2973 18540 3025 18563
rect 3038 18540 3090 18563
rect 3103 18540 3155 18563
rect 3168 18540 3220 18563
rect 3233 18540 3285 18563
rect 3298 18540 3350 18563
rect 3363 18540 3415 18563
rect 3428 18540 3480 18563
rect 3493 18540 3545 18563
rect 3558 18540 3610 18563
rect 3623 18540 3675 18563
rect 3688 18540 3740 18563
rect 3753 18540 3805 18563
rect 3818 18540 3870 18563
rect 3883 18540 3935 18563
rect 3948 18540 4000 18563
rect 4013 18540 4065 18563
rect 4078 18540 4130 18563
rect 4143 18540 4195 18563
rect 4208 18540 4260 18563
rect 4273 18540 4325 18563
rect 4338 18540 4390 18563
rect 4403 18540 4455 18563
rect 4468 18540 4520 18563
rect 4532 18540 4584 18563
rect 2648 18490 2663 18524
rect 2663 18490 2697 18524
rect 2697 18490 2700 18524
rect 2648 18472 2700 18490
rect 2713 18490 2735 18524
rect 2735 18490 2765 18524
rect 2778 18490 2807 18524
rect 2807 18490 2830 18524
rect 2843 18490 2879 18524
rect 2879 18490 2895 18524
rect 2908 18490 2913 18524
rect 2913 18490 2951 18524
rect 2951 18490 2960 18524
rect 2973 18490 2985 18524
rect 2985 18490 3023 18524
rect 3023 18490 3025 18524
rect 3038 18490 3057 18524
rect 3057 18490 3090 18524
rect 3103 18490 3129 18524
rect 3129 18490 3155 18524
rect 3168 18490 3201 18524
rect 3201 18490 3220 18524
rect 2713 18472 2765 18490
rect 2778 18472 2830 18490
rect 2843 18472 2895 18490
rect 2908 18472 2960 18490
rect 2973 18472 3025 18490
rect 3038 18472 3090 18490
rect 3103 18472 3155 18490
rect 3168 18472 3220 18490
rect 3233 18490 3239 18524
rect 3239 18490 3273 18524
rect 3273 18490 3285 18524
rect 3233 18472 3285 18490
rect 3298 18490 3311 18524
rect 3311 18490 3345 18524
rect 3345 18490 3350 18524
rect 3298 18472 3350 18490
rect 3363 18490 3383 18524
rect 3383 18490 3415 18524
rect 3428 18490 3455 18524
rect 3455 18490 3480 18524
rect 3493 18490 3527 18524
rect 3527 18490 3545 18524
rect 3558 18490 3561 18524
rect 3561 18490 3599 18524
rect 3599 18490 3610 18524
rect 3623 18490 3633 18524
rect 3633 18490 3671 18524
rect 3671 18490 3675 18524
rect 3688 18490 3705 18524
rect 3705 18490 3740 18524
rect 3753 18490 3777 18524
rect 3777 18490 3805 18524
rect 3818 18490 3849 18524
rect 3849 18490 3870 18524
rect 3363 18472 3415 18490
rect 3428 18472 3480 18490
rect 3493 18472 3545 18490
rect 3558 18472 3610 18490
rect 3623 18472 3675 18490
rect 3688 18472 3740 18490
rect 3753 18472 3805 18490
rect 3818 18472 3870 18490
rect 3883 18490 3887 18524
rect 3887 18490 3921 18524
rect 3921 18490 3935 18524
rect 3883 18472 3935 18490
rect 3948 18490 3959 18524
rect 3959 18490 3993 18524
rect 3993 18490 4000 18524
rect 3948 18472 4000 18490
rect 4013 18490 4031 18524
rect 4031 18490 4065 18524
rect 4013 18472 4065 18490
rect 4078 18490 4103 18524
rect 4103 18490 4130 18524
rect 4143 18490 4175 18524
rect 4175 18490 4195 18524
rect 4208 18490 4209 18524
rect 4209 18490 4247 18524
rect 4247 18490 4260 18524
rect 4273 18490 4281 18524
rect 4281 18490 4319 18524
rect 4319 18490 4325 18524
rect 4338 18490 4353 18524
rect 4353 18490 4390 18524
rect 4403 18490 4425 18524
rect 4425 18490 4455 18524
rect 4468 18490 4497 18524
rect 4497 18490 4520 18524
rect 4078 18472 4130 18490
rect 4143 18472 4195 18490
rect 4208 18472 4260 18490
rect 4273 18472 4325 18490
rect 4338 18472 4390 18490
rect 4403 18472 4455 18490
rect 4468 18472 4520 18490
rect 4532 18490 4535 18524
rect 4535 18490 4569 18524
rect 4569 18490 4584 18524
rect 4532 18472 4584 18490
rect 2648 18451 2700 18456
rect 2648 18417 2663 18451
rect 2663 18417 2697 18451
rect 2697 18417 2700 18451
rect 2648 18404 2700 18417
rect 2713 18451 2765 18456
rect 2778 18451 2830 18456
rect 2843 18451 2895 18456
rect 2908 18451 2960 18456
rect 2973 18451 3025 18456
rect 3038 18451 3090 18456
rect 3103 18451 3155 18456
rect 3168 18451 3220 18456
rect 2713 18417 2735 18451
rect 2735 18417 2765 18451
rect 2778 18417 2807 18451
rect 2807 18417 2830 18451
rect 2843 18417 2879 18451
rect 2879 18417 2895 18451
rect 2908 18417 2913 18451
rect 2913 18417 2951 18451
rect 2951 18417 2960 18451
rect 2973 18417 2985 18451
rect 2985 18417 3023 18451
rect 3023 18417 3025 18451
rect 3038 18417 3057 18451
rect 3057 18417 3090 18451
rect 3103 18417 3129 18451
rect 3129 18417 3155 18451
rect 3168 18417 3201 18451
rect 3201 18417 3220 18451
rect 2713 18404 2765 18417
rect 2778 18404 2830 18417
rect 2843 18404 2895 18417
rect 2908 18404 2960 18417
rect 2973 18404 3025 18417
rect 3038 18404 3090 18417
rect 3103 18404 3155 18417
rect 3168 18404 3220 18417
rect 3233 18451 3285 18456
rect 3233 18417 3239 18451
rect 3239 18417 3273 18451
rect 3273 18417 3285 18451
rect 3233 18404 3285 18417
rect 3298 18451 3350 18456
rect 3298 18417 3311 18451
rect 3311 18417 3345 18451
rect 3345 18417 3350 18451
rect 3298 18404 3350 18417
rect 3363 18451 3415 18456
rect 3428 18451 3480 18456
rect 3493 18451 3545 18456
rect 3558 18451 3610 18456
rect 3623 18451 3675 18456
rect 3688 18451 3740 18456
rect 3753 18451 3805 18456
rect 3818 18451 3870 18456
rect 3363 18417 3383 18451
rect 3383 18417 3415 18451
rect 3428 18417 3455 18451
rect 3455 18417 3480 18451
rect 3493 18417 3527 18451
rect 3527 18417 3545 18451
rect 3558 18417 3561 18451
rect 3561 18417 3599 18451
rect 3599 18417 3610 18451
rect 3623 18417 3633 18451
rect 3633 18417 3671 18451
rect 3671 18417 3675 18451
rect 3688 18417 3705 18451
rect 3705 18417 3740 18451
rect 3753 18417 3777 18451
rect 3777 18417 3805 18451
rect 3818 18417 3849 18451
rect 3849 18417 3870 18451
rect 3363 18404 3415 18417
rect 3428 18404 3480 18417
rect 3493 18404 3545 18417
rect 3558 18404 3610 18417
rect 3623 18404 3675 18417
rect 3688 18404 3740 18417
rect 3753 18404 3805 18417
rect 3818 18404 3870 18417
rect 3883 18451 3935 18456
rect 3883 18417 3887 18451
rect 3887 18417 3921 18451
rect 3921 18417 3935 18451
rect 3883 18404 3935 18417
rect 3948 18451 4000 18456
rect 3948 18417 3959 18451
rect 3959 18417 3993 18451
rect 3993 18417 4000 18451
rect 3948 18404 4000 18417
rect 4013 18451 4065 18456
rect 4013 18417 4031 18451
rect 4031 18417 4065 18451
rect 4013 18404 4065 18417
rect 4078 18451 4130 18456
rect 4143 18451 4195 18456
rect 4208 18451 4260 18456
rect 4273 18451 4325 18456
rect 4338 18451 4390 18456
rect 4403 18451 4455 18456
rect 4468 18451 4520 18456
rect 4078 18417 4103 18451
rect 4103 18417 4130 18451
rect 4143 18417 4175 18451
rect 4175 18417 4195 18451
rect 4208 18417 4209 18451
rect 4209 18417 4247 18451
rect 4247 18417 4260 18451
rect 4273 18417 4281 18451
rect 4281 18417 4319 18451
rect 4319 18417 4325 18451
rect 4338 18417 4353 18451
rect 4353 18417 4390 18451
rect 4403 18417 4425 18451
rect 4425 18417 4455 18451
rect 4468 18417 4497 18451
rect 4497 18417 4520 18451
rect 4078 18404 4130 18417
rect 4143 18404 4195 18417
rect 4208 18404 4260 18417
rect 4273 18404 4325 18417
rect 4338 18404 4390 18417
rect 4403 18404 4455 18417
rect 4468 18404 4520 18417
rect 4532 18451 4584 18456
rect 4532 18417 4535 18451
rect 4535 18417 4569 18451
rect 4569 18417 4584 18451
rect 4532 18404 4584 18417
rect 2648 18378 2700 18388
rect 2648 18344 2663 18378
rect 2663 18344 2697 18378
rect 2697 18344 2700 18378
rect 2648 18336 2700 18344
rect 2713 18378 2765 18388
rect 2778 18378 2830 18388
rect 2843 18378 2895 18388
rect 2908 18378 2960 18388
rect 2973 18378 3025 18388
rect 3038 18378 3090 18388
rect 3103 18378 3155 18388
rect 3168 18378 3220 18388
rect 2713 18344 2735 18378
rect 2735 18344 2765 18378
rect 2778 18344 2807 18378
rect 2807 18344 2830 18378
rect 2843 18344 2879 18378
rect 2879 18344 2895 18378
rect 2908 18344 2913 18378
rect 2913 18344 2951 18378
rect 2951 18344 2960 18378
rect 2973 18344 2985 18378
rect 2985 18344 3023 18378
rect 3023 18344 3025 18378
rect 3038 18344 3057 18378
rect 3057 18344 3090 18378
rect 3103 18344 3129 18378
rect 3129 18344 3155 18378
rect 3168 18344 3201 18378
rect 3201 18344 3220 18378
rect 2713 18336 2765 18344
rect 2778 18336 2830 18344
rect 2843 18336 2895 18344
rect 2908 18336 2960 18344
rect 2973 18336 3025 18344
rect 3038 18336 3090 18344
rect 3103 18336 3155 18344
rect 3168 18336 3220 18344
rect 3233 18378 3285 18388
rect 3233 18344 3239 18378
rect 3239 18344 3273 18378
rect 3273 18344 3285 18378
rect 3233 18336 3285 18344
rect 3298 18378 3350 18388
rect 3298 18344 3311 18378
rect 3311 18344 3345 18378
rect 3345 18344 3350 18378
rect 3298 18336 3350 18344
rect 3363 18378 3415 18388
rect 3428 18378 3480 18388
rect 3493 18378 3545 18388
rect 3558 18378 3610 18388
rect 3623 18378 3675 18388
rect 3688 18378 3740 18388
rect 3753 18378 3805 18388
rect 3818 18378 3870 18388
rect 3363 18344 3383 18378
rect 3383 18344 3415 18378
rect 3428 18344 3455 18378
rect 3455 18344 3480 18378
rect 3493 18344 3527 18378
rect 3527 18344 3545 18378
rect 3558 18344 3561 18378
rect 3561 18344 3599 18378
rect 3599 18344 3610 18378
rect 3623 18344 3633 18378
rect 3633 18344 3671 18378
rect 3671 18344 3675 18378
rect 3688 18344 3705 18378
rect 3705 18344 3740 18378
rect 3753 18344 3777 18378
rect 3777 18344 3805 18378
rect 3818 18344 3849 18378
rect 3849 18344 3870 18378
rect 3363 18336 3415 18344
rect 3428 18336 3480 18344
rect 3493 18336 3545 18344
rect 3558 18336 3610 18344
rect 3623 18336 3675 18344
rect 3688 18336 3740 18344
rect 3753 18336 3805 18344
rect 3818 18336 3870 18344
rect 3883 18378 3935 18388
rect 3883 18344 3887 18378
rect 3887 18344 3921 18378
rect 3921 18344 3935 18378
rect 3883 18336 3935 18344
rect 3948 18378 4000 18388
rect 3948 18344 3959 18378
rect 3959 18344 3993 18378
rect 3993 18344 4000 18378
rect 3948 18336 4000 18344
rect 4013 18378 4065 18388
rect 4013 18344 4031 18378
rect 4031 18344 4065 18378
rect 4013 18336 4065 18344
rect 4078 18378 4130 18388
rect 4143 18378 4195 18388
rect 4208 18378 4260 18388
rect 4273 18378 4325 18388
rect 4338 18378 4390 18388
rect 4403 18378 4455 18388
rect 4468 18378 4520 18388
rect 4078 18344 4103 18378
rect 4103 18344 4130 18378
rect 4143 18344 4175 18378
rect 4175 18344 4195 18378
rect 4208 18344 4209 18378
rect 4209 18344 4247 18378
rect 4247 18344 4260 18378
rect 4273 18344 4281 18378
rect 4281 18344 4319 18378
rect 4319 18344 4325 18378
rect 4338 18344 4353 18378
rect 4353 18344 4390 18378
rect 4403 18344 4425 18378
rect 4425 18344 4455 18378
rect 4468 18344 4497 18378
rect 4497 18344 4520 18378
rect 4078 18336 4130 18344
rect 4143 18336 4195 18344
rect 4208 18336 4260 18344
rect 4273 18336 4325 18344
rect 4338 18336 4390 18344
rect 4403 18336 4455 18344
rect 4468 18336 4520 18344
rect 4532 18378 4584 18388
rect 4532 18344 4535 18378
rect 4535 18344 4569 18378
rect 4569 18344 4584 18378
rect 4532 18336 4584 18344
rect 2648 18305 2700 18320
rect 2648 18271 2663 18305
rect 2663 18271 2697 18305
rect 2697 18271 2700 18305
rect 2648 18268 2700 18271
rect 2713 18305 2765 18320
rect 2778 18305 2830 18320
rect 2843 18305 2895 18320
rect 2908 18305 2960 18320
rect 2973 18305 3025 18320
rect 3038 18305 3090 18320
rect 3103 18305 3155 18320
rect 3168 18305 3220 18320
rect 2713 18271 2735 18305
rect 2735 18271 2765 18305
rect 2778 18271 2807 18305
rect 2807 18271 2830 18305
rect 2843 18271 2879 18305
rect 2879 18271 2895 18305
rect 2908 18271 2913 18305
rect 2913 18271 2951 18305
rect 2951 18271 2960 18305
rect 2973 18271 2985 18305
rect 2985 18271 3023 18305
rect 3023 18271 3025 18305
rect 3038 18271 3057 18305
rect 3057 18271 3090 18305
rect 3103 18271 3129 18305
rect 3129 18271 3155 18305
rect 3168 18271 3201 18305
rect 3201 18271 3220 18305
rect 2713 18268 2765 18271
rect 2778 18268 2830 18271
rect 2843 18268 2895 18271
rect 2908 18268 2960 18271
rect 2973 18268 3025 18271
rect 3038 18268 3090 18271
rect 3103 18268 3155 18271
rect 3168 18268 3220 18271
rect 3233 18305 3285 18320
rect 3233 18271 3239 18305
rect 3239 18271 3273 18305
rect 3273 18271 3285 18305
rect 3233 18268 3285 18271
rect 3298 18305 3350 18320
rect 3298 18271 3311 18305
rect 3311 18271 3345 18305
rect 3345 18271 3350 18305
rect 3298 18268 3350 18271
rect 3363 18305 3415 18320
rect 3428 18305 3480 18320
rect 3493 18305 3545 18320
rect 3558 18305 3610 18320
rect 3623 18305 3675 18320
rect 3688 18305 3740 18320
rect 3753 18305 3805 18320
rect 3818 18305 3870 18320
rect 3363 18271 3383 18305
rect 3383 18271 3415 18305
rect 3428 18271 3455 18305
rect 3455 18271 3480 18305
rect 3493 18271 3527 18305
rect 3527 18271 3545 18305
rect 3558 18271 3561 18305
rect 3561 18271 3599 18305
rect 3599 18271 3610 18305
rect 3623 18271 3633 18305
rect 3633 18271 3671 18305
rect 3671 18271 3675 18305
rect 3688 18271 3705 18305
rect 3705 18271 3740 18305
rect 3753 18271 3777 18305
rect 3777 18271 3805 18305
rect 3818 18271 3849 18305
rect 3849 18271 3870 18305
rect 3363 18268 3415 18271
rect 3428 18268 3480 18271
rect 3493 18268 3545 18271
rect 3558 18268 3610 18271
rect 3623 18268 3675 18271
rect 3688 18268 3740 18271
rect 3753 18268 3805 18271
rect 3818 18268 3870 18271
rect 3883 18305 3935 18320
rect 3883 18271 3887 18305
rect 3887 18271 3921 18305
rect 3921 18271 3935 18305
rect 3883 18268 3935 18271
rect 3948 18305 4000 18320
rect 3948 18271 3959 18305
rect 3959 18271 3993 18305
rect 3993 18271 4000 18305
rect 3948 18268 4000 18271
rect 4013 18305 4065 18320
rect 4013 18271 4031 18305
rect 4031 18271 4065 18305
rect 4013 18268 4065 18271
rect 4078 18305 4130 18320
rect 4143 18305 4195 18320
rect 4208 18305 4260 18320
rect 4273 18305 4325 18320
rect 4338 18305 4390 18320
rect 4403 18305 4455 18320
rect 4468 18305 4520 18320
rect 4078 18271 4103 18305
rect 4103 18271 4130 18305
rect 4143 18271 4175 18305
rect 4175 18271 4195 18305
rect 4208 18271 4209 18305
rect 4209 18271 4247 18305
rect 4247 18271 4260 18305
rect 4273 18271 4281 18305
rect 4281 18271 4319 18305
rect 4319 18271 4325 18305
rect 4338 18271 4353 18305
rect 4353 18271 4390 18305
rect 4403 18271 4425 18305
rect 4425 18271 4455 18305
rect 4468 18271 4497 18305
rect 4497 18271 4520 18305
rect 4078 18268 4130 18271
rect 4143 18268 4195 18271
rect 4208 18268 4260 18271
rect 4273 18268 4325 18271
rect 4338 18268 4390 18271
rect 4403 18268 4455 18271
rect 4468 18268 4520 18271
rect 4532 18305 4584 18320
rect 4532 18271 4535 18305
rect 4535 18271 4569 18305
rect 4569 18271 4584 18305
rect 4532 18268 4584 18271
rect 2648 18232 2700 18252
rect 2648 18200 2663 18232
rect 2663 18200 2697 18232
rect 2697 18200 2700 18232
rect 2713 18232 2765 18252
rect 2778 18232 2830 18252
rect 2843 18232 2895 18252
rect 2908 18232 2960 18252
rect 2973 18232 3025 18252
rect 3038 18232 3090 18252
rect 3103 18232 3155 18252
rect 3168 18232 3220 18252
rect 2713 18200 2735 18232
rect 2735 18200 2765 18232
rect 2778 18200 2807 18232
rect 2807 18200 2830 18232
rect 2843 18200 2879 18232
rect 2879 18200 2895 18232
rect 2908 18200 2913 18232
rect 2913 18200 2951 18232
rect 2951 18200 2960 18232
rect 2973 18200 2985 18232
rect 2985 18200 3023 18232
rect 3023 18200 3025 18232
rect 3038 18200 3057 18232
rect 3057 18200 3090 18232
rect 3103 18200 3129 18232
rect 3129 18200 3155 18232
rect 3168 18200 3201 18232
rect 3201 18200 3220 18232
rect 3233 18232 3285 18252
rect 3233 18200 3239 18232
rect 3239 18200 3273 18232
rect 3273 18200 3285 18232
rect 3298 18232 3350 18252
rect 3298 18200 3311 18232
rect 3311 18200 3345 18232
rect 3345 18200 3350 18232
rect 3363 18232 3415 18252
rect 3428 18232 3480 18252
rect 3493 18232 3545 18252
rect 3558 18232 3610 18252
rect 3623 18232 3675 18252
rect 3688 18232 3740 18252
rect 3753 18232 3805 18252
rect 3818 18232 3870 18252
rect 3363 18200 3383 18232
rect 3383 18200 3415 18232
rect 3428 18200 3455 18232
rect 3455 18200 3480 18232
rect 3493 18200 3527 18232
rect 3527 18200 3545 18232
rect 3558 18200 3561 18232
rect 3561 18200 3599 18232
rect 3599 18200 3610 18232
rect 3623 18200 3633 18232
rect 3633 18200 3671 18232
rect 3671 18200 3675 18232
rect 3688 18200 3705 18232
rect 3705 18200 3740 18232
rect 3753 18200 3777 18232
rect 3777 18200 3805 18232
rect 3818 18200 3849 18232
rect 3849 18200 3870 18232
rect 3883 18232 3935 18252
rect 3883 18200 3887 18232
rect 3887 18200 3921 18232
rect 3921 18200 3935 18232
rect 3948 18232 4000 18252
rect 3948 18200 3959 18232
rect 3959 18200 3993 18232
rect 3993 18200 4000 18232
rect 4013 18232 4065 18252
rect 4013 18200 4031 18232
rect 4031 18200 4065 18232
rect 4078 18232 4130 18252
rect 4143 18232 4195 18252
rect 4208 18232 4260 18252
rect 4273 18232 4325 18252
rect 4338 18232 4390 18252
rect 4403 18232 4455 18252
rect 4468 18232 4520 18252
rect 4078 18200 4103 18232
rect 4103 18200 4130 18232
rect 4143 18200 4175 18232
rect 4175 18200 4195 18232
rect 4208 18200 4209 18232
rect 4209 18200 4247 18232
rect 4247 18200 4260 18232
rect 4273 18200 4281 18232
rect 4281 18200 4319 18232
rect 4319 18200 4325 18232
rect 4338 18200 4353 18232
rect 4353 18200 4390 18232
rect 4403 18200 4425 18232
rect 4425 18200 4455 18232
rect 4468 18200 4497 18232
rect 4497 18200 4520 18232
rect 4532 18232 4584 18252
rect 4532 18200 4535 18232
rect 4535 18200 4569 18232
rect 4569 18200 4584 18232
rect 2746 16957 2769 16970
rect 2769 16957 2798 16970
rect 2813 16957 2841 16970
rect 2841 16957 2865 16970
rect 2880 16957 2913 16970
rect 2913 16957 2932 16970
rect 2746 16918 2798 16957
rect 2813 16918 2865 16957
rect 2880 16918 2932 16957
rect 2946 16957 2951 16970
rect 2951 16957 2985 16970
rect 2985 16957 2998 16970
rect 2946 16918 2998 16957
rect 3012 16957 3023 16970
rect 3023 16957 3057 16970
rect 3057 16957 3064 16970
rect 3012 16918 3064 16957
rect 3078 16957 3095 16970
rect 3095 16957 3129 16970
rect 3129 16957 3130 16970
rect 3078 16918 3130 16957
rect 3144 16957 3167 16970
rect 3167 16957 3196 16970
rect 3210 16957 3239 16970
rect 3239 16957 3262 16970
rect 3276 16957 3311 16970
rect 3311 16957 3328 16970
rect 3342 16957 3345 16970
rect 3345 16957 3383 16970
rect 3383 16957 3394 16970
rect 3408 16957 3417 16970
rect 3417 16957 3455 16970
rect 3455 16957 3460 16970
rect 3474 16957 3489 16970
rect 3489 16957 3526 16970
rect 3540 16957 3561 16970
rect 3561 16957 3592 16970
rect 3606 16957 3633 16970
rect 3633 16957 3658 16970
rect 3672 16957 3705 16970
rect 3705 16957 3724 16970
rect 3144 16918 3196 16957
rect 3210 16918 3262 16957
rect 3276 16918 3328 16957
rect 3342 16918 3394 16957
rect 3408 16918 3460 16957
rect 3474 16918 3526 16957
rect 3540 16918 3592 16957
rect 3606 16918 3658 16957
rect 3672 16918 3724 16957
rect 3738 16957 3743 16970
rect 3743 16957 3777 16970
rect 3777 16957 3790 16970
rect 3738 16918 3790 16957
rect 3804 16957 3815 16970
rect 3815 16957 3849 16970
rect 3849 16957 3856 16970
rect 3804 16918 3856 16957
rect 3870 16957 3887 16970
rect 3887 16957 3921 16970
rect 3921 16957 3922 16970
rect 3870 16918 3922 16957
rect 3936 16957 3959 16970
rect 3959 16957 3988 16970
rect 4002 16957 4031 16970
rect 4031 16957 4054 16970
rect 4068 16957 4103 16970
rect 4103 16957 4120 16970
rect 4134 16957 4137 16970
rect 4137 16957 4175 16970
rect 4175 16957 4186 16970
rect 4200 16957 4209 16970
rect 4209 16957 4247 16970
rect 4247 16957 4252 16970
rect 4266 16957 4281 16970
rect 4281 16957 4318 16970
rect 4332 16957 4353 16970
rect 4353 16957 4384 16970
rect 4398 16957 4425 16970
rect 4425 16957 4450 16970
rect 4464 16957 4497 16970
rect 4497 16957 4516 16970
rect 3936 16918 3988 16957
rect 4002 16918 4054 16957
rect 4068 16918 4120 16957
rect 4134 16918 4186 16957
rect 4200 16918 4252 16957
rect 4266 16918 4318 16957
rect 4332 16918 4384 16957
rect 4398 16918 4450 16957
rect 4464 16918 4516 16957
rect 2746 16884 2769 16904
rect 2769 16884 2798 16904
rect 2813 16884 2841 16904
rect 2841 16884 2865 16904
rect 2880 16884 2913 16904
rect 2913 16884 2932 16904
rect 2746 16852 2798 16884
rect 2813 16852 2865 16884
rect 2880 16852 2932 16884
rect 2946 16884 2951 16904
rect 2951 16884 2985 16904
rect 2985 16884 2998 16904
rect 2946 16852 2998 16884
rect 3012 16884 3023 16904
rect 3023 16884 3057 16904
rect 3057 16884 3064 16904
rect 3012 16852 3064 16884
rect 3078 16884 3095 16904
rect 3095 16884 3129 16904
rect 3129 16884 3130 16904
rect 3078 16852 3130 16884
rect 3144 16884 3167 16904
rect 3167 16884 3196 16904
rect 3210 16884 3239 16904
rect 3239 16884 3262 16904
rect 3276 16884 3311 16904
rect 3311 16884 3328 16904
rect 3342 16884 3345 16904
rect 3345 16884 3383 16904
rect 3383 16884 3394 16904
rect 3408 16884 3417 16904
rect 3417 16884 3455 16904
rect 3455 16884 3460 16904
rect 3474 16884 3489 16904
rect 3489 16884 3526 16904
rect 3540 16884 3561 16904
rect 3561 16884 3592 16904
rect 3606 16884 3633 16904
rect 3633 16884 3658 16904
rect 3672 16884 3705 16904
rect 3705 16884 3724 16904
rect 3144 16852 3196 16884
rect 3210 16852 3262 16884
rect 3276 16852 3328 16884
rect 3342 16852 3394 16884
rect 3408 16852 3460 16884
rect 3474 16852 3526 16884
rect 3540 16852 3592 16884
rect 3606 16852 3658 16884
rect 3672 16852 3724 16884
rect 3738 16884 3743 16904
rect 3743 16884 3777 16904
rect 3777 16884 3790 16904
rect 3738 16852 3790 16884
rect 3804 16884 3815 16904
rect 3815 16884 3849 16904
rect 3849 16884 3856 16904
rect 3804 16852 3856 16884
rect 3870 16884 3887 16904
rect 3887 16884 3921 16904
rect 3921 16884 3922 16904
rect 3870 16852 3922 16884
rect 3936 16884 3959 16904
rect 3959 16884 3988 16904
rect 4002 16884 4031 16904
rect 4031 16884 4054 16904
rect 4068 16884 4103 16904
rect 4103 16884 4120 16904
rect 4134 16884 4137 16904
rect 4137 16884 4175 16904
rect 4175 16884 4186 16904
rect 4200 16884 4209 16904
rect 4209 16884 4247 16904
rect 4247 16884 4252 16904
rect 4266 16884 4281 16904
rect 4281 16884 4318 16904
rect 4332 16884 4353 16904
rect 4353 16884 4384 16904
rect 4398 16884 4425 16904
rect 4425 16884 4450 16904
rect 4464 16884 4497 16904
rect 4497 16884 4516 16904
rect 3936 16852 3988 16884
rect 4002 16852 4054 16884
rect 4068 16852 4120 16884
rect 4134 16852 4186 16884
rect 4200 16852 4252 16884
rect 4266 16852 4318 16884
rect 4332 16852 4384 16884
rect 4398 16852 4450 16884
rect 4464 16852 4516 16884
rect 2746 16811 2769 16838
rect 2769 16811 2798 16838
rect 2813 16811 2841 16838
rect 2841 16811 2865 16838
rect 2880 16811 2913 16838
rect 2913 16811 2932 16838
rect 2746 16786 2798 16811
rect 2813 16786 2865 16811
rect 2880 16786 2932 16811
rect 2946 16811 2951 16838
rect 2951 16811 2985 16838
rect 2985 16811 2998 16838
rect 2946 16786 2998 16811
rect 3012 16811 3023 16838
rect 3023 16811 3057 16838
rect 3057 16811 3064 16838
rect 3012 16786 3064 16811
rect 3078 16811 3095 16838
rect 3095 16811 3129 16838
rect 3129 16811 3130 16838
rect 3078 16786 3130 16811
rect 3144 16811 3167 16838
rect 3167 16811 3196 16838
rect 3210 16811 3239 16838
rect 3239 16811 3262 16838
rect 3276 16811 3311 16838
rect 3311 16811 3328 16838
rect 3342 16811 3345 16838
rect 3345 16811 3383 16838
rect 3383 16811 3394 16838
rect 3408 16811 3417 16838
rect 3417 16811 3455 16838
rect 3455 16811 3460 16838
rect 3474 16811 3489 16838
rect 3489 16811 3526 16838
rect 3540 16811 3561 16838
rect 3561 16811 3592 16838
rect 3606 16811 3633 16838
rect 3633 16811 3658 16838
rect 3672 16811 3705 16838
rect 3705 16811 3724 16838
rect 3144 16786 3196 16811
rect 3210 16786 3262 16811
rect 3276 16786 3328 16811
rect 3342 16786 3394 16811
rect 3408 16786 3460 16811
rect 3474 16786 3526 16811
rect 3540 16786 3592 16811
rect 3606 16786 3658 16811
rect 3672 16786 3724 16811
rect 3738 16811 3743 16838
rect 3743 16811 3777 16838
rect 3777 16811 3790 16838
rect 3738 16786 3790 16811
rect 3804 16811 3815 16838
rect 3815 16811 3849 16838
rect 3849 16811 3856 16838
rect 3804 16786 3856 16811
rect 3870 16811 3887 16838
rect 3887 16811 3921 16838
rect 3921 16811 3922 16838
rect 3870 16786 3922 16811
rect 3936 16811 3959 16838
rect 3959 16811 3988 16838
rect 4002 16811 4031 16838
rect 4031 16811 4054 16838
rect 4068 16811 4103 16838
rect 4103 16811 4120 16838
rect 4134 16811 4137 16838
rect 4137 16811 4175 16838
rect 4175 16811 4186 16838
rect 4200 16811 4209 16838
rect 4209 16811 4247 16838
rect 4247 16811 4252 16838
rect 4266 16811 4281 16838
rect 4281 16811 4318 16838
rect 4332 16811 4353 16838
rect 4353 16811 4384 16838
rect 4398 16811 4425 16838
rect 4425 16811 4450 16838
rect 4464 16811 4497 16838
rect 4497 16811 4516 16838
rect 3936 16786 3988 16811
rect 4002 16786 4054 16811
rect 4068 16786 4120 16811
rect 4134 16786 4186 16811
rect 4200 16786 4252 16811
rect 4266 16786 4318 16811
rect 4332 16786 4384 16811
rect 4398 16786 4450 16811
rect 4464 16786 4516 16811
rect 2746 16738 2769 16772
rect 2769 16738 2798 16772
rect 2813 16738 2841 16772
rect 2841 16738 2865 16772
rect 2880 16738 2913 16772
rect 2913 16738 2932 16772
rect 2746 16720 2798 16738
rect 2813 16720 2865 16738
rect 2880 16720 2932 16738
rect 2946 16738 2951 16772
rect 2951 16738 2985 16772
rect 2985 16738 2998 16772
rect 2946 16720 2998 16738
rect 3012 16738 3023 16772
rect 3023 16738 3057 16772
rect 3057 16738 3064 16772
rect 3012 16720 3064 16738
rect 3078 16738 3095 16772
rect 3095 16738 3129 16772
rect 3129 16738 3130 16772
rect 3078 16720 3130 16738
rect 3144 16738 3167 16772
rect 3167 16738 3196 16772
rect 3210 16738 3239 16772
rect 3239 16738 3262 16772
rect 3276 16738 3311 16772
rect 3311 16738 3328 16772
rect 3342 16738 3345 16772
rect 3345 16738 3383 16772
rect 3383 16738 3394 16772
rect 3408 16738 3417 16772
rect 3417 16738 3455 16772
rect 3455 16738 3460 16772
rect 3474 16738 3489 16772
rect 3489 16738 3526 16772
rect 3540 16738 3561 16772
rect 3561 16738 3592 16772
rect 3606 16738 3633 16772
rect 3633 16738 3658 16772
rect 3672 16738 3705 16772
rect 3705 16738 3724 16772
rect 3144 16720 3196 16738
rect 3210 16720 3262 16738
rect 3276 16720 3328 16738
rect 3342 16720 3394 16738
rect 3408 16720 3460 16738
rect 3474 16720 3526 16738
rect 3540 16720 3592 16738
rect 3606 16720 3658 16738
rect 3672 16720 3724 16738
rect 3738 16738 3743 16772
rect 3743 16738 3777 16772
rect 3777 16738 3790 16772
rect 3738 16720 3790 16738
rect 3804 16738 3815 16772
rect 3815 16738 3849 16772
rect 3849 16738 3856 16772
rect 3804 16720 3856 16738
rect 3870 16738 3887 16772
rect 3887 16738 3921 16772
rect 3921 16738 3922 16772
rect 3870 16720 3922 16738
rect 3936 16738 3959 16772
rect 3959 16738 3988 16772
rect 4002 16738 4031 16772
rect 4031 16738 4054 16772
rect 4068 16738 4103 16772
rect 4103 16738 4120 16772
rect 4134 16738 4137 16772
rect 4137 16738 4175 16772
rect 4175 16738 4186 16772
rect 4200 16738 4209 16772
rect 4209 16738 4247 16772
rect 4247 16738 4252 16772
rect 4266 16738 4281 16772
rect 4281 16738 4318 16772
rect 4332 16738 4353 16772
rect 4353 16738 4384 16772
rect 4398 16738 4425 16772
rect 4425 16738 4450 16772
rect 4464 16738 4497 16772
rect 4497 16738 4516 16772
rect 3936 16720 3988 16738
rect 4002 16720 4054 16738
rect 4068 16720 4120 16738
rect 4134 16720 4186 16738
rect 4200 16720 4252 16738
rect 4266 16720 4318 16738
rect 4332 16720 4384 16738
rect 4398 16720 4450 16738
rect 4464 16720 4516 16738
rect 2746 16699 2798 16706
rect 2813 16699 2865 16706
rect 2880 16699 2932 16706
rect 2746 16665 2769 16699
rect 2769 16665 2798 16699
rect 2813 16665 2841 16699
rect 2841 16665 2865 16699
rect 2880 16665 2913 16699
rect 2913 16665 2932 16699
rect 2746 16654 2798 16665
rect 2813 16654 2865 16665
rect 2880 16654 2932 16665
rect 2946 16699 2998 16706
rect 2946 16665 2951 16699
rect 2951 16665 2985 16699
rect 2985 16665 2998 16699
rect 2946 16654 2998 16665
rect 3012 16699 3064 16706
rect 3012 16665 3023 16699
rect 3023 16665 3057 16699
rect 3057 16665 3064 16699
rect 3012 16654 3064 16665
rect 3078 16699 3130 16706
rect 3078 16665 3095 16699
rect 3095 16665 3129 16699
rect 3129 16665 3130 16699
rect 3078 16654 3130 16665
rect 3144 16699 3196 16706
rect 3210 16699 3262 16706
rect 3276 16699 3328 16706
rect 3342 16699 3394 16706
rect 3408 16699 3460 16706
rect 3474 16699 3526 16706
rect 3540 16699 3592 16706
rect 3606 16699 3658 16706
rect 3672 16699 3724 16706
rect 3144 16665 3167 16699
rect 3167 16665 3196 16699
rect 3210 16665 3239 16699
rect 3239 16665 3262 16699
rect 3276 16665 3311 16699
rect 3311 16665 3328 16699
rect 3342 16665 3345 16699
rect 3345 16665 3383 16699
rect 3383 16665 3394 16699
rect 3408 16665 3417 16699
rect 3417 16665 3455 16699
rect 3455 16665 3460 16699
rect 3474 16665 3489 16699
rect 3489 16665 3526 16699
rect 3540 16665 3561 16699
rect 3561 16665 3592 16699
rect 3606 16665 3633 16699
rect 3633 16665 3658 16699
rect 3672 16665 3705 16699
rect 3705 16665 3724 16699
rect 3144 16654 3196 16665
rect 3210 16654 3262 16665
rect 3276 16654 3328 16665
rect 3342 16654 3394 16665
rect 3408 16654 3460 16665
rect 3474 16654 3526 16665
rect 3540 16654 3592 16665
rect 3606 16654 3658 16665
rect 3672 16654 3724 16665
rect 3738 16699 3790 16706
rect 3738 16665 3743 16699
rect 3743 16665 3777 16699
rect 3777 16665 3790 16699
rect 3738 16654 3790 16665
rect 3804 16699 3856 16706
rect 3804 16665 3815 16699
rect 3815 16665 3849 16699
rect 3849 16665 3856 16699
rect 3804 16654 3856 16665
rect 3870 16699 3922 16706
rect 3870 16665 3887 16699
rect 3887 16665 3921 16699
rect 3921 16665 3922 16699
rect 3870 16654 3922 16665
rect 3936 16699 3988 16706
rect 4002 16699 4054 16706
rect 4068 16699 4120 16706
rect 4134 16699 4186 16706
rect 4200 16699 4252 16706
rect 4266 16699 4318 16706
rect 4332 16699 4384 16706
rect 4398 16699 4450 16706
rect 4464 16699 4516 16706
rect 3936 16665 3959 16699
rect 3959 16665 3988 16699
rect 4002 16665 4031 16699
rect 4031 16665 4054 16699
rect 4068 16665 4103 16699
rect 4103 16665 4120 16699
rect 4134 16665 4137 16699
rect 4137 16665 4175 16699
rect 4175 16665 4186 16699
rect 4200 16665 4209 16699
rect 4209 16665 4247 16699
rect 4247 16665 4252 16699
rect 4266 16665 4281 16699
rect 4281 16665 4318 16699
rect 4332 16665 4353 16699
rect 4353 16665 4384 16699
rect 4398 16665 4425 16699
rect 4425 16665 4450 16699
rect 4464 16665 4497 16699
rect 4497 16665 4516 16699
rect 3936 16654 3988 16665
rect 4002 16654 4054 16665
rect 4068 16654 4120 16665
rect 4134 16654 4186 16665
rect 4200 16654 4252 16665
rect 4266 16654 4318 16665
rect 4332 16654 4384 16665
rect 4398 16654 4450 16665
rect 4464 16654 4516 16665
rect 2746 16626 2798 16640
rect 2813 16626 2865 16640
rect 2880 16626 2932 16640
rect 2746 16592 2769 16626
rect 2769 16592 2798 16626
rect 2813 16592 2841 16626
rect 2841 16592 2865 16626
rect 2880 16592 2913 16626
rect 2913 16592 2932 16626
rect 2746 16588 2798 16592
rect 2813 16588 2865 16592
rect 2880 16588 2932 16592
rect 2946 16626 2998 16640
rect 2946 16592 2951 16626
rect 2951 16592 2985 16626
rect 2985 16592 2998 16626
rect 2946 16588 2998 16592
rect 3012 16626 3064 16640
rect 3012 16592 3023 16626
rect 3023 16592 3057 16626
rect 3057 16592 3064 16626
rect 3012 16588 3064 16592
rect 3078 16626 3130 16640
rect 3078 16592 3095 16626
rect 3095 16592 3129 16626
rect 3129 16592 3130 16626
rect 3078 16588 3130 16592
rect 3144 16626 3196 16640
rect 3210 16626 3262 16640
rect 3276 16626 3328 16640
rect 3342 16626 3394 16640
rect 3408 16626 3460 16640
rect 3474 16626 3526 16640
rect 3540 16626 3592 16640
rect 3606 16626 3658 16640
rect 3672 16626 3724 16640
rect 3144 16592 3167 16626
rect 3167 16592 3196 16626
rect 3210 16592 3239 16626
rect 3239 16592 3262 16626
rect 3276 16592 3311 16626
rect 3311 16592 3328 16626
rect 3342 16592 3345 16626
rect 3345 16592 3383 16626
rect 3383 16592 3394 16626
rect 3408 16592 3417 16626
rect 3417 16592 3455 16626
rect 3455 16592 3460 16626
rect 3474 16592 3489 16626
rect 3489 16592 3526 16626
rect 3540 16592 3561 16626
rect 3561 16592 3592 16626
rect 3606 16592 3633 16626
rect 3633 16592 3658 16626
rect 3672 16592 3705 16626
rect 3705 16592 3724 16626
rect 3144 16588 3196 16592
rect 3210 16588 3262 16592
rect 3276 16588 3328 16592
rect 3342 16588 3394 16592
rect 3408 16588 3460 16592
rect 3474 16588 3526 16592
rect 3540 16588 3592 16592
rect 3606 16588 3658 16592
rect 3672 16588 3724 16592
rect 3738 16626 3790 16640
rect 3738 16592 3743 16626
rect 3743 16592 3777 16626
rect 3777 16592 3790 16626
rect 3738 16588 3790 16592
rect 3804 16626 3856 16640
rect 3804 16592 3815 16626
rect 3815 16592 3849 16626
rect 3849 16592 3856 16626
rect 3804 16588 3856 16592
rect 3870 16626 3922 16640
rect 3870 16592 3887 16626
rect 3887 16592 3921 16626
rect 3921 16592 3922 16626
rect 3870 16588 3922 16592
rect 3936 16626 3988 16640
rect 4002 16626 4054 16640
rect 4068 16626 4120 16640
rect 4134 16626 4186 16640
rect 4200 16626 4252 16640
rect 4266 16626 4318 16640
rect 4332 16626 4384 16640
rect 4398 16626 4450 16640
rect 4464 16626 4516 16640
rect 3936 16592 3959 16626
rect 3959 16592 3988 16626
rect 4002 16592 4031 16626
rect 4031 16592 4054 16626
rect 4068 16592 4103 16626
rect 4103 16592 4120 16626
rect 4134 16592 4137 16626
rect 4137 16592 4175 16626
rect 4175 16592 4186 16626
rect 4200 16592 4209 16626
rect 4209 16592 4247 16626
rect 4247 16592 4252 16626
rect 4266 16592 4281 16626
rect 4281 16592 4318 16626
rect 4332 16592 4353 16626
rect 4353 16592 4384 16626
rect 4398 16592 4425 16626
rect 4425 16592 4450 16626
rect 4464 16592 4497 16626
rect 4497 16592 4516 16626
rect 3936 16588 3988 16592
rect 4002 16588 4054 16592
rect 4068 16588 4120 16592
rect 4134 16588 4186 16592
rect 4200 16588 4252 16592
rect 4266 16588 4318 16592
rect 4332 16588 4384 16592
rect 4398 16588 4450 16592
rect 4464 16588 4516 16592
rect 2746 16553 2798 16574
rect 2813 16553 2865 16574
rect 2880 16553 2932 16574
rect 2746 16522 2769 16553
rect 2769 16522 2798 16553
rect 2813 16522 2841 16553
rect 2841 16522 2865 16553
rect 2880 16522 2913 16553
rect 2913 16522 2932 16553
rect 2946 16553 2998 16574
rect 2946 16522 2951 16553
rect 2951 16522 2985 16553
rect 2985 16522 2998 16553
rect 3012 16553 3064 16574
rect 3012 16522 3023 16553
rect 3023 16522 3057 16553
rect 3057 16522 3064 16553
rect 3078 16553 3130 16574
rect 3078 16522 3095 16553
rect 3095 16522 3129 16553
rect 3129 16522 3130 16553
rect 3144 16553 3196 16574
rect 3210 16553 3262 16574
rect 3276 16553 3328 16574
rect 3342 16553 3394 16574
rect 3408 16553 3460 16574
rect 3474 16553 3526 16574
rect 3540 16553 3592 16574
rect 3606 16553 3658 16574
rect 3672 16553 3724 16574
rect 3144 16522 3167 16553
rect 3167 16522 3196 16553
rect 3210 16522 3239 16553
rect 3239 16522 3262 16553
rect 3276 16522 3311 16553
rect 3311 16522 3328 16553
rect 3342 16522 3345 16553
rect 3345 16522 3383 16553
rect 3383 16522 3394 16553
rect 3408 16522 3417 16553
rect 3417 16522 3455 16553
rect 3455 16522 3460 16553
rect 3474 16522 3489 16553
rect 3489 16522 3526 16553
rect 3540 16522 3561 16553
rect 3561 16522 3592 16553
rect 3606 16522 3633 16553
rect 3633 16522 3658 16553
rect 3672 16522 3705 16553
rect 3705 16522 3724 16553
rect 3738 16553 3790 16574
rect 3738 16522 3743 16553
rect 3743 16522 3777 16553
rect 3777 16522 3790 16553
rect 3804 16553 3856 16574
rect 3804 16522 3815 16553
rect 3815 16522 3849 16553
rect 3849 16522 3856 16553
rect 3870 16553 3922 16574
rect 3870 16522 3887 16553
rect 3887 16522 3921 16553
rect 3921 16522 3922 16553
rect 3936 16553 3988 16574
rect 4002 16553 4054 16574
rect 4068 16553 4120 16574
rect 4134 16553 4186 16574
rect 4200 16553 4252 16574
rect 4266 16553 4318 16574
rect 4332 16553 4384 16574
rect 4398 16553 4450 16574
rect 4464 16553 4516 16574
rect 3936 16522 3959 16553
rect 3959 16522 3988 16553
rect 4002 16522 4031 16553
rect 4031 16522 4054 16553
rect 4068 16522 4103 16553
rect 4103 16522 4120 16553
rect 4134 16522 4137 16553
rect 4137 16522 4175 16553
rect 4175 16522 4186 16553
rect 4200 16522 4209 16553
rect 4209 16522 4247 16553
rect 4247 16522 4252 16553
rect 4266 16522 4281 16553
rect 4281 16522 4318 16553
rect 4332 16522 4353 16553
rect 4353 16522 4384 16553
rect 4398 16522 4425 16553
rect 4425 16522 4450 16553
rect 4464 16522 4497 16553
rect 4497 16522 4516 16553
rect 2746 16480 2798 16508
rect 2813 16480 2865 16508
rect 2880 16480 2932 16508
rect 2746 16456 2769 16480
rect 2769 16456 2798 16480
rect 2813 16456 2841 16480
rect 2841 16456 2865 16480
rect 2880 16456 2913 16480
rect 2913 16456 2932 16480
rect 2946 16480 2998 16508
rect 2946 16456 2951 16480
rect 2951 16456 2985 16480
rect 2985 16456 2998 16480
rect 3012 16480 3064 16508
rect 3012 16456 3023 16480
rect 3023 16456 3057 16480
rect 3057 16456 3064 16480
rect 3078 16480 3130 16508
rect 3078 16456 3095 16480
rect 3095 16456 3129 16480
rect 3129 16456 3130 16480
rect 3144 16480 3196 16508
rect 3210 16480 3262 16508
rect 3276 16480 3328 16508
rect 3342 16480 3394 16508
rect 3408 16480 3460 16508
rect 3474 16480 3526 16508
rect 3540 16480 3592 16508
rect 3606 16480 3658 16508
rect 3672 16480 3724 16508
rect 3144 16456 3167 16480
rect 3167 16456 3196 16480
rect 3210 16456 3239 16480
rect 3239 16456 3262 16480
rect 3276 16456 3311 16480
rect 3311 16456 3328 16480
rect 3342 16456 3345 16480
rect 3345 16456 3383 16480
rect 3383 16456 3394 16480
rect 3408 16456 3417 16480
rect 3417 16456 3455 16480
rect 3455 16456 3460 16480
rect 3474 16456 3489 16480
rect 3489 16456 3526 16480
rect 3540 16456 3561 16480
rect 3561 16456 3592 16480
rect 3606 16456 3633 16480
rect 3633 16456 3658 16480
rect 3672 16456 3705 16480
rect 3705 16456 3724 16480
rect 3738 16480 3790 16508
rect 3738 16456 3743 16480
rect 3743 16456 3777 16480
rect 3777 16456 3790 16480
rect 3804 16480 3856 16508
rect 3804 16456 3815 16480
rect 3815 16456 3849 16480
rect 3849 16456 3856 16480
rect 3870 16480 3922 16508
rect 3870 16456 3887 16480
rect 3887 16456 3921 16480
rect 3921 16456 3922 16480
rect 3936 16480 3988 16508
rect 4002 16480 4054 16508
rect 4068 16480 4120 16508
rect 4134 16480 4186 16508
rect 4200 16480 4252 16508
rect 4266 16480 4318 16508
rect 4332 16480 4384 16508
rect 4398 16480 4450 16508
rect 4464 16480 4516 16508
rect 3936 16456 3959 16480
rect 3959 16456 3988 16480
rect 4002 16456 4031 16480
rect 4031 16456 4054 16480
rect 4068 16456 4103 16480
rect 4103 16456 4120 16480
rect 4134 16456 4137 16480
rect 4137 16456 4175 16480
rect 4175 16456 4186 16480
rect 4200 16456 4209 16480
rect 4209 16456 4247 16480
rect 4247 16456 4252 16480
rect 4266 16456 4281 16480
rect 4281 16456 4318 16480
rect 4332 16456 4353 16480
rect 4353 16456 4384 16480
rect 4398 16456 4425 16480
rect 4425 16456 4450 16480
rect 4464 16456 4497 16480
rect 4497 16456 4516 16480
rect 2746 16407 2798 16442
rect 2813 16407 2865 16442
rect 2880 16407 2932 16442
rect 2746 16390 2769 16407
rect 2769 16390 2798 16407
rect 2813 16390 2841 16407
rect 2841 16390 2865 16407
rect 2880 16390 2913 16407
rect 2913 16390 2932 16407
rect 2946 16407 2998 16442
rect 2946 16390 2951 16407
rect 2951 16390 2985 16407
rect 2985 16390 2998 16407
rect 3012 16407 3064 16442
rect 3012 16390 3023 16407
rect 3023 16390 3057 16407
rect 3057 16390 3064 16407
rect 3078 16407 3130 16442
rect 3078 16390 3095 16407
rect 3095 16390 3129 16407
rect 3129 16390 3130 16407
rect 3144 16407 3196 16442
rect 3210 16407 3262 16442
rect 3276 16407 3328 16442
rect 3342 16407 3394 16442
rect 3408 16407 3460 16442
rect 3474 16407 3526 16442
rect 3540 16407 3592 16442
rect 3606 16407 3658 16442
rect 3672 16407 3724 16442
rect 3144 16390 3167 16407
rect 3167 16390 3196 16407
rect 3210 16390 3239 16407
rect 3239 16390 3262 16407
rect 3276 16390 3311 16407
rect 3311 16390 3328 16407
rect 3342 16390 3345 16407
rect 3345 16390 3383 16407
rect 3383 16390 3394 16407
rect 3408 16390 3417 16407
rect 3417 16390 3455 16407
rect 3455 16390 3460 16407
rect 3474 16390 3489 16407
rect 3489 16390 3526 16407
rect 3540 16390 3561 16407
rect 3561 16390 3592 16407
rect 3606 16390 3633 16407
rect 3633 16390 3658 16407
rect 3672 16390 3705 16407
rect 3705 16390 3724 16407
rect 3738 16407 3790 16442
rect 3738 16390 3743 16407
rect 3743 16390 3777 16407
rect 3777 16390 3790 16407
rect 3804 16407 3856 16442
rect 3804 16390 3815 16407
rect 3815 16390 3849 16407
rect 3849 16390 3856 16407
rect 3870 16407 3922 16442
rect 3870 16390 3887 16407
rect 3887 16390 3921 16407
rect 3921 16390 3922 16407
rect 3936 16407 3988 16442
rect 4002 16407 4054 16442
rect 4068 16407 4120 16442
rect 4134 16407 4186 16442
rect 4200 16407 4252 16442
rect 4266 16407 4318 16442
rect 4332 16407 4384 16442
rect 4398 16407 4450 16442
rect 4464 16407 4516 16442
rect 3936 16390 3959 16407
rect 3959 16390 3988 16407
rect 4002 16390 4031 16407
rect 4031 16390 4054 16407
rect 4068 16390 4103 16407
rect 4103 16390 4120 16407
rect 4134 16390 4137 16407
rect 4137 16390 4175 16407
rect 4175 16390 4186 16407
rect 4200 16390 4209 16407
rect 4209 16390 4247 16407
rect 4247 16390 4252 16407
rect 4266 16390 4281 16407
rect 4281 16390 4318 16407
rect 4332 16390 4353 16407
rect 4353 16390 4384 16407
rect 4398 16390 4425 16407
rect 4425 16390 4450 16407
rect 4464 16390 4497 16407
rect 4497 16390 4516 16407
rect 2746 16373 2769 16376
rect 2769 16373 2798 16376
rect 2813 16373 2841 16376
rect 2841 16373 2865 16376
rect 2880 16373 2913 16376
rect 2913 16373 2932 16376
rect 2746 16334 2798 16373
rect 2813 16334 2865 16373
rect 2880 16334 2932 16373
rect 2746 16324 2769 16334
rect 2769 16324 2798 16334
rect 2813 16324 2841 16334
rect 2841 16324 2865 16334
rect 2880 16324 2913 16334
rect 2913 16324 2932 16334
rect 2946 16373 2951 16376
rect 2951 16373 2985 16376
rect 2985 16373 2998 16376
rect 2946 16334 2998 16373
rect 2946 16324 2951 16334
rect 2951 16324 2985 16334
rect 2985 16324 2998 16334
rect 3012 16373 3023 16376
rect 3023 16373 3057 16376
rect 3057 16373 3064 16376
rect 3012 16334 3064 16373
rect 3012 16324 3023 16334
rect 3023 16324 3057 16334
rect 3057 16324 3064 16334
rect 3078 16373 3095 16376
rect 3095 16373 3129 16376
rect 3129 16373 3130 16376
rect 3078 16334 3130 16373
rect 3078 16324 3095 16334
rect 3095 16324 3129 16334
rect 3129 16324 3130 16334
rect 3144 16373 3167 16376
rect 3167 16373 3196 16376
rect 3210 16373 3239 16376
rect 3239 16373 3262 16376
rect 3276 16373 3311 16376
rect 3311 16373 3328 16376
rect 3342 16373 3345 16376
rect 3345 16373 3383 16376
rect 3383 16373 3394 16376
rect 3408 16373 3417 16376
rect 3417 16373 3455 16376
rect 3455 16373 3460 16376
rect 3474 16373 3489 16376
rect 3489 16373 3526 16376
rect 3540 16373 3561 16376
rect 3561 16373 3592 16376
rect 3606 16373 3633 16376
rect 3633 16373 3658 16376
rect 3672 16373 3705 16376
rect 3705 16373 3724 16376
rect 3144 16334 3196 16373
rect 3210 16334 3262 16373
rect 3276 16334 3328 16373
rect 3342 16334 3394 16373
rect 3408 16334 3460 16373
rect 3474 16334 3526 16373
rect 3540 16334 3592 16373
rect 3606 16334 3658 16373
rect 3672 16334 3724 16373
rect 3144 16324 3167 16334
rect 3167 16324 3196 16334
rect 3210 16324 3239 16334
rect 3239 16324 3262 16334
rect 3276 16324 3311 16334
rect 3311 16324 3328 16334
rect 3342 16324 3345 16334
rect 3345 16324 3383 16334
rect 3383 16324 3394 16334
rect 3408 16324 3417 16334
rect 3417 16324 3455 16334
rect 3455 16324 3460 16334
rect 3474 16324 3489 16334
rect 3489 16324 3526 16334
rect 3540 16324 3561 16334
rect 3561 16324 3592 16334
rect 3606 16324 3633 16334
rect 3633 16324 3658 16334
rect 3672 16324 3705 16334
rect 3705 16324 3724 16334
rect 3738 16373 3743 16376
rect 3743 16373 3777 16376
rect 3777 16373 3790 16376
rect 3738 16334 3790 16373
rect 3738 16324 3743 16334
rect 3743 16324 3777 16334
rect 3777 16324 3790 16334
rect 3804 16373 3815 16376
rect 3815 16373 3849 16376
rect 3849 16373 3856 16376
rect 3804 16334 3856 16373
rect 3804 16324 3815 16334
rect 3815 16324 3849 16334
rect 3849 16324 3856 16334
rect 3870 16373 3887 16376
rect 3887 16373 3921 16376
rect 3921 16373 3922 16376
rect 3870 16334 3922 16373
rect 3870 16324 3887 16334
rect 3887 16324 3921 16334
rect 3921 16324 3922 16334
rect 3936 16373 3959 16376
rect 3959 16373 3988 16376
rect 4002 16373 4031 16376
rect 4031 16373 4054 16376
rect 4068 16373 4103 16376
rect 4103 16373 4120 16376
rect 4134 16373 4137 16376
rect 4137 16373 4175 16376
rect 4175 16373 4186 16376
rect 4200 16373 4209 16376
rect 4209 16373 4247 16376
rect 4247 16373 4252 16376
rect 4266 16373 4281 16376
rect 4281 16373 4318 16376
rect 4332 16373 4353 16376
rect 4353 16373 4384 16376
rect 4398 16373 4425 16376
rect 4425 16373 4450 16376
rect 4464 16373 4497 16376
rect 4497 16373 4516 16376
rect 3936 16334 3988 16373
rect 4002 16334 4054 16373
rect 4068 16334 4120 16373
rect 4134 16334 4186 16373
rect 4200 16334 4252 16373
rect 4266 16334 4318 16373
rect 4332 16334 4384 16373
rect 4398 16334 4450 16373
rect 4464 16334 4516 16373
rect 3936 16324 3959 16334
rect 3959 16324 3988 16334
rect 4002 16324 4031 16334
rect 4031 16324 4054 16334
rect 4068 16324 4103 16334
rect 4103 16324 4120 16334
rect 4134 16324 4137 16334
rect 4137 16324 4175 16334
rect 4175 16324 4186 16334
rect 4200 16324 4209 16334
rect 4209 16324 4247 16334
rect 4247 16324 4252 16334
rect 4266 16324 4281 16334
rect 4281 16324 4318 16334
rect 4332 16324 4353 16334
rect 4353 16324 4384 16334
rect 4398 16324 4425 16334
rect 4425 16324 4450 16334
rect 4464 16324 4497 16334
rect 4497 16324 4516 16334
rect 2746 16300 2769 16310
rect 2769 16300 2798 16310
rect 2813 16300 2841 16310
rect 2841 16300 2865 16310
rect 2880 16300 2913 16310
rect 2913 16300 2932 16310
rect 2746 16261 2798 16300
rect 2813 16261 2865 16300
rect 2880 16261 2932 16300
rect 2746 16258 2769 16261
rect 2769 16258 2798 16261
rect 2813 16258 2841 16261
rect 2841 16258 2865 16261
rect 2880 16258 2913 16261
rect 2913 16258 2932 16261
rect 2946 16300 2951 16310
rect 2951 16300 2985 16310
rect 2985 16300 2998 16310
rect 2946 16261 2998 16300
rect 2946 16258 2951 16261
rect 2951 16258 2985 16261
rect 2985 16258 2998 16261
rect 3012 16300 3023 16310
rect 3023 16300 3057 16310
rect 3057 16300 3064 16310
rect 3012 16261 3064 16300
rect 3012 16258 3023 16261
rect 3023 16258 3057 16261
rect 3057 16258 3064 16261
rect 3078 16300 3095 16310
rect 3095 16300 3129 16310
rect 3129 16300 3130 16310
rect 3078 16261 3130 16300
rect 3078 16258 3095 16261
rect 3095 16258 3129 16261
rect 3129 16258 3130 16261
rect 3144 16300 3167 16310
rect 3167 16300 3196 16310
rect 3210 16300 3239 16310
rect 3239 16300 3262 16310
rect 3276 16300 3311 16310
rect 3311 16300 3328 16310
rect 3342 16300 3345 16310
rect 3345 16300 3383 16310
rect 3383 16300 3394 16310
rect 3408 16300 3417 16310
rect 3417 16300 3455 16310
rect 3455 16300 3460 16310
rect 3474 16300 3489 16310
rect 3489 16300 3526 16310
rect 3540 16300 3561 16310
rect 3561 16300 3592 16310
rect 3606 16300 3633 16310
rect 3633 16300 3658 16310
rect 3672 16300 3705 16310
rect 3705 16300 3724 16310
rect 3144 16261 3196 16300
rect 3210 16261 3262 16300
rect 3276 16261 3328 16300
rect 3342 16261 3394 16300
rect 3408 16261 3460 16300
rect 3474 16261 3526 16300
rect 3540 16261 3592 16300
rect 3606 16261 3658 16300
rect 3672 16261 3724 16300
rect 3144 16258 3167 16261
rect 3167 16258 3196 16261
rect 3210 16258 3239 16261
rect 3239 16258 3262 16261
rect 3276 16258 3311 16261
rect 3311 16258 3328 16261
rect 3342 16258 3345 16261
rect 3345 16258 3383 16261
rect 3383 16258 3394 16261
rect 3408 16258 3417 16261
rect 3417 16258 3455 16261
rect 3455 16258 3460 16261
rect 3474 16258 3489 16261
rect 3489 16258 3526 16261
rect 3540 16258 3561 16261
rect 3561 16258 3592 16261
rect 3606 16258 3633 16261
rect 3633 16258 3658 16261
rect 3672 16258 3705 16261
rect 3705 16258 3724 16261
rect 3738 16300 3743 16310
rect 3743 16300 3777 16310
rect 3777 16300 3790 16310
rect 3738 16261 3790 16300
rect 3738 16258 3743 16261
rect 3743 16258 3777 16261
rect 3777 16258 3790 16261
rect 3804 16300 3815 16310
rect 3815 16300 3849 16310
rect 3849 16300 3856 16310
rect 3804 16261 3856 16300
rect 3804 16258 3815 16261
rect 3815 16258 3849 16261
rect 3849 16258 3856 16261
rect 3870 16300 3887 16310
rect 3887 16300 3921 16310
rect 3921 16300 3922 16310
rect 3870 16261 3922 16300
rect 3870 16258 3887 16261
rect 3887 16258 3921 16261
rect 3921 16258 3922 16261
rect 3936 16300 3959 16310
rect 3959 16300 3988 16310
rect 4002 16300 4031 16310
rect 4031 16300 4054 16310
rect 4068 16300 4103 16310
rect 4103 16300 4120 16310
rect 4134 16300 4137 16310
rect 4137 16300 4175 16310
rect 4175 16300 4186 16310
rect 4200 16300 4209 16310
rect 4209 16300 4247 16310
rect 4247 16300 4252 16310
rect 4266 16300 4281 16310
rect 4281 16300 4318 16310
rect 4332 16300 4353 16310
rect 4353 16300 4384 16310
rect 4398 16300 4425 16310
rect 4425 16300 4450 16310
rect 4464 16300 4497 16310
rect 4497 16300 4516 16310
rect 3936 16261 3988 16300
rect 4002 16261 4054 16300
rect 4068 16261 4120 16300
rect 4134 16261 4186 16300
rect 4200 16261 4252 16300
rect 4266 16261 4318 16300
rect 4332 16261 4384 16300
rect 4398 16261 4450 16300
rect 4464 16261 4516 16300
rect 3936 16258 3959 16261
rect 3959 16258 3988 16261
rect 4002 16258 4031 16261
rect 4031 16258 4054 16261
rect 4068 16258 4103 16261
rect 4103 16258 4120 16261
rect 4134 16258 4137 16261
rect 4137 16258 4175 16261
rect 4175 16258 4186 16261
rect 4200 16258 4209 16261
rect 4209 16258 4247 16261
rect 4247 16258 4252 16261
rect 4266 16258 4281 16261
rect 4281 16258 4318 16261
rect 4332 16258 4353 16261
rect 4353 16258 4384 16261
rect 4398 16258 4425 16261
rect 4425 16258 4450 16261
rect 4464 16258 4497 16261
rect 4497 16258 4516 16261
rect 2746 16227 2769 16244
rect 2769 16227 2798 16244
rect 2813 16227 2841 16244
rect 2841 16227 2865 16244
rect 2880 16227 2913 16244
rect 2913 16227 2932 16244
rect 2746 16192 2798 16227
rect 2813 16192 2865 16227
rect 2880 16192 2932 16227
rect 2946 16227 2951 16244
rect 2951 16227 2985 16244
rect 2985 16227 2998 16244
rect 2946 16192 2998 16227
rect 3012 16227 3023 16244
rect 3023 16227 3057 16244
rect 3057 16227 3064 16244
rect 3012 16192 3064 16227
rect 3078 16227 3095 16244
rect 3095 16227 3129 16244
rect 3129 16227 3130 16244
rect 3078 16192 3130 16227
rect 3144 16227 3167 16244
rect 3167 16227 3196 16244
rect 3210 16227 3239 16244
rect 3239 16227 3262 16244
rect 3276 16227 3311 16244
rect 3311 16227 3328 16244
rect 3342 16227 3345 16244
rect 3345 16227 3383 16244
rect 3383 16227 3394 16244
rect 3408 16227 3417 16244
rect 3417 16227 3455 16244
rect 3455 16227 3460 16244
rect 3474 16227 3489 16244
rect 3489 16227 3526 16244
rect 3540 16227 3561 16244
rect 3561 16227 3592 16244
rect 3606 16227 3633 16244
rect 3633 16227 3658 16244
rect 3672 16227 3705 16244
rect 3705 16227 3724 16244
rect 3144 16192 3196 16227
rect 3210 16192 3262 16227
rect 3276 16192 3328 16227
rect 3342 16192 3394 16227
rect 3408 16192 3460 16227
rect 3474 16192 3526 16227
rect 3540 16192 3592 16227
rect 3606 16192 3658 16227
rect 3672 16192 3724 16227
rect 3738 16227 3743 16244
rect 3743 16227 3777 16244
rect 3777 16227 3790 16244
rect 3738 16192 3790 16227
rect 3804 16227 3815 16244
rect 3815 16227 3849 16244
rect 3849 16227 3856 16244
rect 3804 16192 3856 16227
rect 3870 16227 3887 16244
rect 3887 16227 3921 16244
rect 3921 16227 3922 16244
rect 3870 16192 3922 16227
rect 3936 16227 3959 16244
rect 3959 16227 3988 16244
rect 4002 16227 4031 16244
rect 4031 16227 4054 16244
rect 4068 16227 4103 16244
rect 4103 16227 4120 16244
rect 4134 16227 4137 16244
rect 4137 16227 4175 16244
rect 4175 16227 4186 16244
rect 4200 16227 4209 16244
rect 4209 16227 4247 16244
rect 4247 16227 4252 16244
rect 4266 16227 4281 16244
rect 4281 16227 4318 16244
rect 4332 16227 4353 16244
rect 4353 16227 4384 16244
rect 4398 16227 4425 16244
rect 4425 16227 4450 16244
rect 4464 16227 4497 16244
rect 4497 16227 4516 16244
rect 3936 16192 3988 16227
rect 4002 16192 4054 16227
rect 4068 16192 4120 16227
rect 4134 16192 4186 16227
rect 4200 16192 4252 16227
rect 4266 16192 4318 16227
rect 4332 16192 4384 16227
rect 4398 16192 4450 16227
rect 4464 16192 4516 16227
rect 2746 16154 2769 16178
rect 2769 16154 2798 16178
rect 2813 16154 2841 16178
rect 2841 16154 2865 16178
rect 2880 16154 2913 16178
rect 2913 16154 2932 16178
rect 2746 16126 2798 16154
rect 2813 16126 2865 16154
rect 2880 16126 2932 16154
rect 2946 16154 2951 16178
rect 2951 16154 2985 16178
rect 2985 16154 2998 16178
rect 2946 16126 2998 16154
rect 3012 16154 3023 16178
rect 3023 16154 3057 16178
rect 3057 16154 3064 16178
rect 3012 16126 3064 16154
rect 3078 16154 3095 16178
rect 3095 16154 3129 16178
rect 3129 16154 3130 16178
rect 3078 16126 3130 16154
rect 3144 16154 3167 16178
rect 3167 16154 3196 16178
rect 3210 16154 3239 16178
rect 3239 16154 3262 16178
rect 3276 16154 3311 16178
rect 3311 16154 3328 16178
rect 3342 16154 3345 16178
rect 3345 16154 3383 16178
rect 3383 16154 3394 16178
rect 3408 16154 3417 16178
rect 3417 16154 3455 16178
rect 3455 16154 3460 16178
rect 3474 16154 3489 16178
rect 3489 16154 3526 16178
rect 3540 16154 3561 16178
rect 3561 16154 3592 16178
rect 3606 16154 3633 16178
rect 3633 16154 3658 16178
rect 3672 16154 3705 16178
rect 3705 16154 3724 16178
rect 3144 16126 3196 16154
rect 3210 16126 3262 16154
rect 3276 16126 3328 16154
rect 3342 16126 3394 16154
rect 3408 16126 3460 16154
rect 3474 16126 3526 16154
rect 3540 16126 3592 16154
rect 3606 16126 3658 16154
rect 3672 16126 3724 16154
rect 3738 16154 3743 16178
rect 3743 16154 3777 16178
rect 3777 16154 3790 16178
rect 3738 16126 3790 16154
rect 3804 16154 3815 16178
rect 3815 16154 3849 16178
rect 3849 16154 3856 16178
rect 3804 16126 3856 16154
rect 3870 16154 3887 16178
rect 3887 16154 3921 16178
rect 3921 16154 3922 16178
rect 3870 16126 3922 16154
rect 3936 16154 3959 16178
rect 3959 16154 3988 16178
rect 4002 16154 4031 16178
rect 4031 16154 4054 16178
rect 4068 16154 4103 16178
rect 4103 16154 4120 16178
rect 4134 16154 4137 16178
rect 4137 16154 4175 16178
rect 4175 16154 4186 16178
rect 4200 16154 4209 16178
rect 4209 16154 4247 16178
rect 4247 16154 4252 16178
rect 4266 16154 4281 16178
rect 4281 16154 4318 16178
rect 4332 16154 4353 16178
rect 4353 16154 4384 16178
rect 4398 16154 4425 16178
rect 4425 16154 4450 16178
rect 4464 16154 4497 16178
rect 4497 16154 4516 16178
rect 3936 16126 3988 16154
rect 4002 16126 4054 16154
rect 4068 16126 4120 16154
rect 4134 16126 4186 16154
rect 4200 16126 4252 16154
rect 4266 16126 4318 16154
rect 4332 16126 4384 16154
rect 4398 16126 4450 16154
rect 4464 16126 4516 16154
rect 2746 16081 2769 16112
rect 2769 16081 2798 16112
rect 2813 16081 2841 16112
rect 2841 16081 2865 16112
rect 2880 16081 2913 16112
rect 2913 16081 2932 16112
rect 2746 16060 2798 16081
rect 2813 16060 2865 16081
rect 2880 16060 2932 16081
rect 2946 16081 2951 16112
rect 2951 16081 2985 16112
rect 2985 16081 2998 16112
rect 2946 16060 2998 16081
rect 3012 16081 3023 16112
rect 3023 16081 3057 16112
rect 3057 16081 3064 16112
rect 3012 16060 3064 16081
rect 3078 16081 3095 16112
rect 3095 16081 3129 16112
rect 3129 16081 3130 16112
rect 3078 16060 3130 16081
rect 3144 16081 3167 16112
rect 3167 16081 3196 16112
rect 3210 16081 3239 16112
rect 3239 16081 3262 16112
rect 3276 16081 3311 16112
rect 3311 16081 3328 16112
rect 3342 16081 3345 16112
rect 3345 16081 3383 16112
rect 3383 16081 3394 16112
rect 3408 16081 3417 16112
rect 3417 16081 3455 16112
rect 3455 16081 3460 16112
rect 3474 16081 3489 16112
rect 3489 16081 3526 16112
rect 3540 16081 3561 16112
rect 3561 16081 3592 16112
rect 3606 16081 3633 16112
rect 3633 16081 3658 16112
rect 3672 16081 3705 16112
rect 3705 16081 3724 16112
rect 3144 16060 3196 16081
rect 3210 16060 3262 16081
rect 3276 16060 3328 16081
rect 3342 16060 3394 16081
rect 3408 16060 3460 16081
rect 3474 16060 3526 16081
rect 3540 16060 3592 16081
rect 3606 16060 3658 16081
rect 3672 16060 3724 16081
rect 3738 16081 3743 16112
rect 3743 16081 3777 16112
rect 3777 16081 3790 16112
rect 3738 16060 3790 16081
rect 3804 16081 3815 16112
rect 3815 16081 3849 16112
rect 3849 16081 3856 16112
rect 3804 16060 3856 16081
rect 3870 16081 3887 16112
rect 3887 16081 3921 16112
rect 3921 16081 3922 16112
rect 3870 16060 3922 16081
rect 3936 16081 3959 16112
rect 3959 16081 3988 16112
rect 4002 16081 4031 16112
rect 4031 16081 4054 16112
rect 4068 16081 4103 16112
rect 4103 16081 4120 16112
rect 4134 16081 4137 16112
rect 4137 16081 4175 16112
rect 4175 16081 4186 16112
rect 4200 16081 4209 16112
rect 4209 16081 4247 16112
rect 4247 16081 4252 16112
rect 4266 16081 4281 16112
rect 4281 16081 4318 16112
rect 4332 16081 4353 16112
rect 4353 16081 4384 16112
rect 4398 16081 4425 16112
rect 4425 16081 4450 16112
rect 4464 16081 4497 16112
rect 4497 16081 4516 16112
rect 3936 16060 3988 16081
rect 4002 16060 4054 16081
rect 4068 16060 4120 16081
rect 4134 16060 4186 16081
rect 4200 16060 4252 16081
rect 4266 16060 4318 16081
rect 4332 16060 4384 16081
rect 4398 16060 4450 16081
rect 4464 16060 4516 16081
rect 2746 16042 2798 16046
rect 2813 16042 2865 16046
rect 2880 16042 2932 16046
rect 2746 16008 2769 16042
rect 2769 16008 2798 16042
rect 2813 16008 2841 16042
rect 2841 16008 2865 16042
rect 2880 16008 2913 16042
rect 2913 16008 2932 16042
rect 2746 15994 2798 16008
rect 2813 15994 2865 16008
rect 2880 15994 2932 16008
rect 2946 16042 2998 16046
rect 2946 16008 2951 16042
rect 2951 16008 2985 16042
rect 2985 16008 2998 16042
rect 2946 15994 2998 16008
rect 3012 16042 3064 16046
rect 3012 16008 3023 16042
rect 3023 16008 3057 16042
rect 3057 16008 3064 16042
rect 3012 15994 3064 16008
rect 3078 16042 3130 16046
rect 3078 16008 3095 16042
rect 3095 16008 3129 16042
rect 3129 16008 3130 16042
rect 3078 15994 3130 16008
rect 3144 16042 3196 16046
rect 3210 16042 3262 16046
rect 3276 16042 3328 16046
rect 3342 16042 3394 16046
rect 3408 16042 3460 16046
rect 3474 16042 3526 16046
rect 3540 16042 3592 16046
rect 3606 16042 3658 16046
rect 3672 16042 3724 16046
rect 3144 16008 3167 16042
rect 3167 16008 3196 16042
rect 3210 16008 3239 16042
rect 3239 16008 3262 16042
rect 3276 16008 3311 16042
rect 3311 16008 3328 16042
rect 3342 16008 3345 16042
rect 3345 16008 3383 16042
rect 3383 16008 3394 16042
rect 3408 16008 3417 16042
rect 3417 16008 3455 16042
rect 3455 16008 3460 16042
rect 3474 16008 3489 16042
rect 3489 16008 3526 16042
rect 3540 16008 3561 16042
rect 3561 16008 3592 16042
rect 3606 16008 3633 16042
rect 3633 16008 3658 16042
rect 3672 16008 3705 16042
rect 3705 16008 3724 16042
rect 3144 15994 3196 16008
rect 3210 15994 3262 16008
rect 3276 15994 3328 16008
rect 3342 15994 3394 16008
rect 3408 15994 3460 16008
rect 3474 15994 3526 16008
rect 3540 15994 3592 16008
rect 3606 15994 3658 16008
rect 3672 15994 3724 16008
rect 3738 16042 3790 16046
rect 3738 16008 3743 16042
rect 3743 16008 3777 16042
rect 3777 16008 3790 16042
rect 3738 15994 3790 16008
rect 3804 16042 3856 16046
rect 3804 16008 3815 16042
rect 3815 16008 3849 16042
rect 3849 16008 3856 16042
rect 3804 15994 3856 16008
rect 3870 16042 3922 16046
rect 3870 16008 3887 16042
rect 3887 16008 3921 16042
rect 3921 16008 3922 16042
rect 3870 15994 3922 16008
rect 3936 16042 3988 16046
rect 4002 16042 4054 16046
rect 4068 16042 4120 16046
rect 4134 16042 4186 16046
rect 4200 16042 4252 16046
rect 4266 16042 4318 16046
rect 4332 16042 4384 16046
rect 4398 16042 4450 16046
rect 4464 16042 4516 16046
rect 3936 16008 3959 16042
rect 3959 16008 3988 16042
rect 4002 16008 4031 16042
rect 4031 16008 4054 16042
rect 4068 16008 4103 16042
rect 4103 16008 4120 16042
rect 4134 16008 4137 16042
rect 4137 16008 4175 16042
rect 4175 16008 4186 16042
rect 4200 16008 4209 16042
rect 4209 16008 4247 16042
rect 4247 16008 4252 16042
rect 4266 16008 4281 16042
rect 4281 16008 4318 16042
rect 4332 16008 4353 16042
rect 4353 16008 4384 16042
rect 4398 16008 4425 16042
rect 4425 16008 4450 16042
rect 4464 16008 4497 16042
rect 4497 16008 4516 16042
rect 3936 15994 3988 16008
rect 4002 15994 4054 16008
rect 4068 15994 4120 16008
rect 4134 15994 4186 16008
rect 4200 15994 4252 16008
rect 4266 15994 4318 16008
rect 4332 15994 4384 16008
rect 4398 15994 4450 16008
rect 4464 15994 4516 16008
rect 5040 28714 5092 28720
rect 5040 28680 5046 28714
rect 5046 28680 5080 28714
rect 5080 28680 5092 28714
rect 5040 28668 5092 28680
rect 5106 28714 5158 28720
rect 5106 28680 5118 28714
rect 5118 28680 5152 28714
rect 5152 28680 5158 28714
rect 5106 28668 5158 28680
rect 5040 28641 5092 28651
rect 5040 28607 5046 28641
rect 5046 28607 5080 28641
rect 5080 28607 5092 28641
rect 5040 28599 5092 28607
rect 5106 28641 5158 28651
rect 5106 28607 5118 28641
rect 5118 28607 5152 28641
rect 5152 28607 5158 28641
rect 5106 28599 5158 28607
rect 5040 28568 5092 28582
rect 5040 28534 5046 28568
rect 5046 28534 5080 28568
rect 5080 28534 5092 28568
rect 5040 28530 5092 28534
rect 5106 28568 5158 28582
rect 5106 28534 5118 28568
rect 5118 28534 5152 28568
rect 5152 28534 5158 28568
rect 5106 28530 5158 28534
rect 5040 28495 5092 28513
rect 5040 28461 5046 28495
rect 5046 28461 5080 28495
rect 5080 28461 5092 28495
rect 5106 28495 5158 28513
rect 5106 28461 5118 28495
rect 5118 28461 5152 28495
rect 5152 28461 5158 28495
rect 5040 28422 5092 28444
rect 5106 28422 5158 28444
rect 5040 28392 5046 28422
rect 5046 28392 5092 28422
rect 5106 28392 5152 28422
rect 5152 28392 5158 28422
rect 5040 28323 5046 28375
rect 5046 28323 5092 28375
rect 5106 28323 5152 28375
rect 5152 28323 5158 28375
rect 5040 28254 5046 28306
rect 5046 28254 5092 28306
rect 5106 28254 5152 28306
rect 5152 28254 5158 28306
rect 5040 28184 5046 28236
rect 5046 28184 5092 28236
rect 5106 28184 5152 28236
rect 5152 28184 5158 28236
rect 5040 28114 5046 28166
rect 5046 28114 5092 28166
rect 5106 28114 5152 28166
rect 5152 28114 5158 28166
rect 5317 27930 5323 27982
rect 5323 27930 5369 27982
rect 5383 27930 5429 27982
rect 5429 27930 5435 27982
rect 5317 27861 5323 27913
rect 5323 27861 5369 27913
rect 5383 27861 5429 27913
rect 5429 27861 5435 27913
rect 5317 27792 5323 27844
rect 5323 27792 5369 27844
rect 5383 27792 5429 27844
rect 5429 27792 5435 27844
rect 5317 27723 5323 27775
rect 5323 27723 5369 27775
rect 5383 27723 5429 27775
rect 5429 27723 5435 27775
rect 5317 27654 5323 27706
rect 5323 27654 5369 27706
rect 5383 27654 5429 27706
rect 5429 27654 5435 27706
rect 5317 27584 5323 27636
rect 5323 27584 5369 27636
rect 5383 27584 5429 27636
rect 5429 27584 5435 27636
rect 5317 27514 5323 27566
rect 5323 27514 5369 27566
rect 5383 27514 5429 27566
rect 5429 27514 5435 27566
rect 5317 27444 5323 27496
rect 5323 27444 5369 27496
rect 5383 27444 5429 27496
rect 5429 27444 5435 27496
rect 5317 27380 5323 27426
rect 5323 27380 5369 27426
rect 5383 27380 5429 27426
rect 5429 27380 5435 27426
rect 5317 27374 5369 27380
rect 5383 27374 5435 27380
rect 5594 28714 5646 28720
rect 5594 28680 5600 28714
rect 5600 28680 5634 28714
rect 5634 28680 5646 28714
rect 5594 28668 5646 28680
rect 5660 28714 5712 28720
rect 5660 28680 5672 28714
rect 5672 28680 5706 28714
rect 5706 28680 5712 28714
rect 5660 28668 5712 28680
rect 5594 28641 5646 28651
rect 5594 28607 5600 28641
rect 5600 28607 5634 28641
rect 5634 28607 5646 28641
rect 5594 28599 5646 28607
rect 5660 28641 5712 28651
rect 5660 28607 5672 28641
rect 5672 28607 5706 28641
rect 5706 28607 5712 28641
rect 5660 28599 5712 28607
rect 5594 28568 5646 28582
rect 5594 28534 5600 28568
rect 5600 28534 5634 28568
rect 5634 28534 5646 28568
rect 5594 28530 5646 28534
rect 5660 28568 5712 28582
rect 5660 28534 5672 28568
rect 5672 28534 5706 28568
rect 5706 28534 5712 28568
rect 5660 28530 5712 28534
rect 5594 28495 5646 28513
rect 5594 28461 5600 28495
rect 5600 28461 5634 28495
rect 5634 28461 5646 28495
rect 5660 28495 5712 28513
rect 5660 28461 5672 28495
rect 5672 28461 5706 28495
rect 5706 28461 5712 28495
rect 5594 28422 5646 28444
rect 5660 28422 5712 28444
rect 5594 28392 5600 28422
rect 5600 28392 5646 28422
rect 5660 28392 5706 28422
rect 5706 28392 5712 28422
rect 5594 28323 5600 28375
rect 5600 28323 5646 28375
rect 5660 28323 5706 28375
rect 5706 28323 5712 28375
rect 5594 28254 5600 28306
rect 5600 28254 5646 28306
rect 5660 28254 5706 28306
rect 5706 28254 5712 28306
rect 5594 28184 5600 28236
rect 5600 28184 5646 28236
rect 5660 28184 5706 28236
rect 5706 28184 5712 28236
rect 5594 28114 5600 28166
rect 5600 28114 5646 28166
rect 5660 28114 5706 28166
rect 5706 28114 5712 28166
rect 5871 27930 5877 27982
rect 5877 27930 5923 27982
rect 5937 27930 5983 27982
rect 5983 27930 5989 27982
rect 5871 27861 5877 27913
rect 5877 27861 5923 27913
rect 5937 27861 5983 27913
rect 5983 27861 5989 27913
rect 5871 27792 5877 27844
rect 5877 27792 5923 27844
rect 5937 27792 5983 27844
rect 5983 27792 5989 27844
rect 5871 27723 5877 27775
rect 5877 27723 5923 27775
rect 5937 27723 5983 27775
rect 5983 27723 5989 27775
rect 5871 27654 5877 27706
rect 5877 27654 5923 27706
rect 5937 27654 5983 27706
rect 5983 27654 5989 27706
rect 5871 27584 5877 27636
rect 5877 27584 5923 27636
rect 5937 27584 5983 27636
rect 5983 27584 5989 27636
rect 5871 27514 5877 27566
rect 5877 27514 5923 27566
rect 5937 27514 5983 27566
rect 5983 27514 5989 27566
rect 5871 27444 5877 27496
rect 5877 27444 5923 27496
rect 5937 27444 5983 27496
rect 5983 27444 5989 27496
rect 5871 27380 5877 27426
rect 5877 27380 5923 27426
rect 5937 27380 5983 27426
rect 5983 27380 5989 27426
rect 5871 27374 5923 27380
rect 5937 27374 5989 27380
rect 6148 28714 6200 28720
rect 6148 28680 6154 28714
rect 6154 28680 6188 28714
rect 6188 28680 6200 28714
rect 6148 28668 6200 28680
rect 6214 28714 6266 28720
rect 6214 28680 6226 28714
rect 6226 28680 6260 28714
rect 6260 28680 6266 28714
rect 6214 28668 6266 28680
rect 6148 28641 6200 28651
rect 6148 28607 6154 28641
rect 6154 28607 6188 28641
rect 6188 28607 6200 28641
rect 6148 28599 6200 28607
rect 6214 28641 6266 28651
rect 6214 28607 6226 28641
rect 6226 28607 6260 28641
rect 6260 28607 6266 28641
rect 6214 28599 6266 28607
rect 6148 28568 6200 28582
rect 6148 28534 6154 28568
rect 6154 28534 6188 28568
rect 6188 28534 6200 28568
rect 6148 28530 6200 28534
rect 6214 28568 6266 28582
rect 6214 28534 6226 28568
rect 6226 28534 6260 28568
rect 6260 28534 6266 28568
rect 6214 28530 6266 28534
rect 6148 28495 6200 28513
rect 6148 28461 6154 28495
rect 6154 28461 6188 28495
rect 6188 28461 6200 28495
rect 6214 28495 6266 28513
rect 6214 28461 6226 28495
rect 6226 28461 6260 28495
rect 6260 28461 6266 28495
rect 6148 28422 6200 28444
rect 6214 28422 6266 28444
rect 6148 28392 6154 28422
rect 6154 28392 6200 28422
rect 6214 28392 6260 28422
rect 6260 28392 6266 28422
rect 6148 28323 6154 28375
rect 6154 28323 6200 28375
rect 6214 28323 6260 28375
rect 6260 28323 6266 28375
rect 6148 28254 6154 28306
rect 6154 28254 6200 28306
rect 6214 28254 6260 28306
rect 6260 28254 6266 28306
rect 6148 28184 6154 28236
rect 6154 28184 6200 28236
rect 6214 28184 6260 28236
rect 6260 28184 6266 28236
rect 6148 28114 6154 28166
rect 6154 28114 6200 28166
rect 6214 28114 6260 28166
rect 6260 28114 6266 28166
rect 6425 27930 6431 27982
rect 6431 27930 6477 27982
rect 6491 27930 6537 27982
rect 6537 27930 6543 27982
rect 6425 27861 6431 27913
rect 6431 27861 6477 27913
rect 6491 27861 6537 27913
rect 6537 27861 6543 27913
rect 6425 27792 6431 27844
rect 6431 27792 6477 27844
rect 6491 27792 6537 27844
rect 6537 27792 6543 27844
rect 6425 27723 6431 27775
rect 6431 27723 6477 27775
rect 6491 27723 6537 27775
rect 6537 27723 6543 27775
rect 6425 27654 6431 27706
rect 6431 27654 6477 27706
rect 6491 27654 6537 27706
rect 6537 27654 6543 27706
rect 6425 27584 6431 27636
rect 6431 27584 6477 27636
rect 6491 27584 6537 27636
rect 6537 27584 6543 27636
rect 6425 27514 6431 27566
rect 6431 27514 6477 27566
rect 6491 27514 6537 27566
rect 6537 27514 6543 27566
rect 6425 27444 6431 27496
rect 6431 27444 6477 27496
rect 6491 27444 6537 27496
rect 6537 27444 6543 27496
rect 6425 27380 6431 27426
rect 6431 27380 6477 27426
rect 6491 27380 6537 27426
rect 6537 27380 6543 27426
rect 6425 27374 6477 27380
rect 6491 27374 6543 27380
rect 6702 28714 6754 28720
rect 6702 28680 6708 28714
rect 6708 28680 6742 28714
rect 6742 28680 6754 28714
rect 6702 28668 6754 28680
rect 6768 28714 6820 28720
rect 6768 28680 6780 28714
rect 6780 28680 6814 28714
rect 6814 28680 6820 28714
rect 6768 28668 6820 28680
rect 6702 28641 6754 28651
rect 6702 28607 6708 28641
rect 6708 28607 6742 28641
rect 6742 28607 6754 28641
rect 6702 28599 6754 28607
rect 6768 28641 6820 28651
rect 6768 28607 6780 28641
rect 6780 28607 6814 28641
rect 6814 28607 6820 28641
rect 6768 28599 6820 28607
rect 6702 28568 6754 28582
rect 6702 28534 6708 28568
rect 6708 28534 6742 28568
rect 6742 28534 6754 28568
rect 6702 28530 6754 28534
rect 6768 28568 6820 28582
rect 6768 28534 6780 28568
rect 6780 28534 6814 28568
rect 6814 28534 6820 28568
rect 6768 28530 6820 28534
rect 6702 28495 6754 28513
rect 6702 28461 6708 28495
rect 6708 28461 6742 28495
rect 6742 28461 6754 28495
rect 6768 28495 6820 28513
rect 6768 28461 6780 28495
rect 6780 28461 6814 28495
rect 6814 28461 6820 28495
rect 6702 28422 6754 28444
rect 6768 28422 6820 28444
rect 6702 28392 6708 28422
rect 6708 28392 6754 28422
rect 6768 28392 6814 28422
rect 6814 28392 6820 28422
rect 6702 28323 6708 28375
rect 6708 28323 6754 28375
rect 6768 28323 6814 28375
rect 6814 28323 6820 28375
rect 6702 28254 6708 28306
rect 6708 28254 6754 28306
rect 6768 28254 6814 28306
rect 6814 28254 6820 28306
rect 6702 28184 6708 28236
rect 6708 28184 6754 28236
rect 6768 28184 6814 28236
rect 6814 28184 6820 28236
rect 6702 28114 6708 28166
rect 6708 28114 6754 28166
rect 6768 28114 6814 28166
rect 6814 28114 6820 28166
rect 6979 27930 6985 27982
rect 6985 27930 7031 27982
rect 7045 27930 7091 27982
rect 7091 27930 7097 27982
rect 6979 27861 6985 27913
rect 6985 27861 7031 27913
rect 7045 27861 7091 27913
rect 7091 27861 7097 27913
rect 6979 27792 6985 27844
rect 6985 27792 7031 27844
rect 7045 27792 7091 27844
rect 7091 27792 7097 27844
rect 6979 27723 6985 27775
rect 6985 27723 7031 27775
rect 7045 27723 7091 27775
rect 7091 27723 7097 27775
rect 6979 27654 6985 27706
rect 6985 27654 7031 27706
rect 7045 27654 7091 27706
rect 7091 27654 7097 27706
rect 6979 27584 6985 27636
rect 6985 27584 7031 27636
rect 7045 27584 7091 27636
rect 7091 27584 7097 27636
rect 6979 27514 6985 27566
rect 6985 27514 7031 27566
rect 7045 27514 7091 27566
rect 7091 27514 7097 27566
rect 6979 27444 6985 27496
rect 6985 27444 7031 27496
rect 7045 27444 7091 27496
rect 7091 27444 7097 27496
rect 6979 27380 6985 27426
rect 6985 27380 7031 27426
rect 7045 27380 7091 27426
rect 7091 27380 7097 27426
rect 6979 27374 7031 27380
rect 7045 27374 7097 27380
rect 7256 28714 7308 28720
rect 7256 28680 7262 28714
rect 7262 28680 7296 28714
rect 7296 28680 7308 28714
rect 7256 28668 7308 28680
rect 7322 28714 7374 28720
rect 7322 28680 7334 28714
rect 7334 28680 7368 28714
rect 7368 28680 7374 28714
rect 7322 28668 7374 28680
rect 7256 28641 7308 28651
rect 7256 28607 7262 28641
rect 7262 28607 7296 28641
rect 7296 28607 7308 28641
rect 7256 28599 7308 28607
rect 7322 28641 7374 28651
rect 7322 28607 7334 28641
rect 7334 28607 7368 28641
rect 7368 28607 7374 28641
rect 7322 28599 7374 28607
rect 7256 28568 7308 28582
rect 7256 28534 7262 28568
rect 7262 28534 7296 28568
rect 7296 28534 7308 28568
rect 7256 28530 7308 28534
rect 7322 28568 7374 28582
rect 7322 28534 7334 28568
rect 7334 28534 7368 28568
rect 7368 28534 7374 28568
rect 7322 28530 7374 28534
rect 7256 28495 7308 28513
rect 7256 28461 7262 28495
rect 7262 28461 7296 28495
rect 7296 28461 7308 28495
rect 7322 28495 7374 28513
rect 7322 28461 7334 28495
rect 7334 28461 7368 28495
rect 7368 28461 7374 28495
rect 7256 28422 7308 28444
rect 7322 28422 7374 28444
rect 7256 28392 7262 28422
rect 7262 28392 7308 28422
rect 7322 28392 7368 28422
rect 7368 28392 7374 28422
rect 7256 28323 7262 28375
rect 7262 28323 7308 28375
rect 7322 28323 7368 28375
rect 7368 28323 7374 28375
rect 7256 28254 7262 28306
rect 7262 28254 7308 28306
rect 7322 28254 7368 28306
rect 7368 28254 7374 28306
rect 7256 28184 7262 28236
rect 7262 28184 7308 28236
rect 7322 28184 7368 28236
rect 7368 28184 7374 28236
rect 7256 28114 7262 28166
rect 7262 28114 7308 28166
rect 7322 28114 7368 28166
rect 7368 28114 7374 28166
rect 7533 27930 7539 27982
rect 7539 27930 7585 27982
rect 7599 27930 7645 27982
rect 7645 27930 7651 27982
rect 7533 27861 7539 27913
rect 7539 27861 7585 27913
rect 7599 27861 7645 27913
rect 7645 27861 7651 27913
rect 7533 27792 7539 27844
rect 7539 27792 7585 27844
rect 7599 27792 7645 27844
rect 7645 27792 7651 27844
rect 7533 27723 7539 27775
rect 7539 27723 7585 27775
rect 7599 27723 7645 27775
rect 7645 27723 7651 27775
rect 7533 27654 7539 27706
rect 7539 27654 7585 27706
rect 7599 27654 7645 27706
rect 7645 27654 7651 27706
rect 7533 27584 7539 27636
rect 7539 27584 7585 27636
rect 7599 27584 7645 27636
rect 7645 27584 7651 27636
rect 7533 27514 7539 27566
rect 7539 27514 7585 27566
rect 7599 27514 7645 27566
rect 7645 27514 7651 27566
rect 7533 27444 7539 27496
rect 7539 27444 7585 27496
rect 7599 27444 7645 27496
rect 7645 27444 7651 27496
rect 7533 27380 7539 27426
rect 7539 27380 7585 27426
rect 7599 27380 7645 27426
rect 7645 27380 7651 27426
rect 7533 27374 7585 27380
rect 7599 27374 7651 27380
rect 7810 28714 7862 28720
rect 7810 28680 7816 28714
rect 7816 28680 7850 28714
rect 7850 28680 7862 28714
rect 7810 28668 7862 28680
rect 7876 28714 7928 28720
rect 7876 28680 7888 28714
rect 7888 28680 7922 28714
rect 7922 28680 7928 28714
rect 7876 28668 7928 28680
rect 7810 28641 7862 28651
rect 7810 28607 7816 28641
rect 7816 28607 7850 28641
rect 7850 28607 7862 28641
rect 7810 28599 7862 28607
rect 7876 28641 7928 28651
rect 7876 28607 7888 28641
rect 7888 28607 7922 28641
rect 7922 28607 7928 28641
rect 7876 28599 7928 28607
rect 7810 28568 7862 28582
rect 7810 28534 7816 28568
rect 7816 28534 7850 28568
rect 7850 28534 7862 28568
rect 7810 28530 7862 28534
rect 7876 28568 7928 28582
rect 7876 28534 7888 28568
rect 7888 28534 7922 28568
rect 7922 28534 7928 28568
rect 7876 28530 7928 28534
rect 7810 28495 7862 28513
rect 7810 28461 7816 28495
rect 7816 28461 7850 28495
rect 7850 28461 7862 28495
rect 7876 28495 7928 28513
rect 7876 28461 7888 28495
rect 7888 28461 7922 28495
rect 7922 28461 7928 28495
rect 7810 28422 7862 28444
rect 7876 28422 7928 28444
rect 7810 28392 7816 28422
rect 7816 28392 7862 28422
rect 7876 28392 7922 28422
rect 7922 28392 7928 28422
rect 7810 28323 7816 28375
rect 7816 28323 7862 28375
rect 7876 28323 7922 28375
rect 7922 28323 7928 28375
rect 7810 28254 7816 28306
rect 7816 28254 7862 28306
rect 7876 28254 7922 28306
rect 7922 28254 7928 28306
rect 7810 28184 7816 28236
rect 7816 28184 7862 28236
rect 7876 28184 7922 28236
rect 7922 28184 7928 28236
rect 7810 28114 7816 28166
rect 7816 28114 7862 28166
rect 7876 28114 7922 28166
rect 7922 28114 7928 28166
rect 8047 28711 8099 28724
rect 8047 28677 8050 28711
rect 8050 28677 8084 28711
rect 8084 28677 8099 28711
rect 8047 28672 8099 28677
rect 8169 28701 8221 28724
rect 8169 28672 8184 28701
rect 8184 28672 8218 28701
rect 8218 28672 8221 28701
rect 8047 28639 8099 28655
rect 8047 28605 8050 28639
rect 8050 28605 8084 28639
rect 8084 28605 8099 28639
rect 8047 28603 8099 28605
rect 8169 28629 8221 28655
rect 8169 28603 8184 28629
rect 8184 28603 8218 28629
rect 8218 28603 8221 28629
rect 8047 28567 8099 28586
rect 8047 28534 8050 28567
rect 8050 28534 8084 28567
rect 8084 28534 8099 28567
rect 8169 28557 8221 28586
rect 8169 28534 8184 28557
rect 8184 28534 8218 28557
rect 8218 28534 8221 28557
rect 8047 28495 8099 28517
rect 8047 28465 8050 28495
rect 8050 28465 8084 28495
rect 8084 28465 8099 28495
rect 8169 28485 8221 28517
rect 8169 28465 8184 28485
rect 8184 28465 8218 28485
rect 8218 28465 8221 28485
rect 8047 28423 8099 28448
rect 8047 28396 8050 28423
rect 8050 28396 8084 28423
rect 8084 28396 8099 28423
rect 8169 28413 8221 28448
rect 8169 28396 8184 28413
rect 8184 28396 8218 28413
rect 8218 28396 8221 28413
rect 8047 28351 8099 28378
rect 8047 28326 8050 28351
rect 8050 28326 8084 28351
rect 8084 28326 8099 28351
rect 8169 28341 8221 28378
rect 8169 28326 8184 28341
rect 8184 28326 8218 28341
rect 8218 28326 8221 28341
rect 8047 28279 8099 28308
rect 8047 28256 8050 28279
rect 8050 28256 8084 28279
rect 8084 28256 8099 28279
rect 8169 28307 8184 28308
rect 8184 28307 8218 28308
rect 8218 28307 8221 28308
rect 8169 28269 8221 28307
rect 8169 28256 8184 28269
rect 8184 28256 8218 28269
rect 8218 28256 8221 28269
rect 8047 28207 8099 28238
rect 8047 28186 8050 28207
rect 8050 28186 8084 28207
rect 8084 28186 8099 28207
rect 8169 28235 8184 28238
rect 8184 28235 8218 28238
rect 8218 28235 8221 28238
rect 8169 28197 8221 28235
rect 8169 28186 8184 28197
rect 8184 28186 8218 28197
rect 8218 28186 8221 28197
rect 8047 28135 8099 28168
rect 8047 28116 8050 28135
rect 8050 28116 8084 28135
rect 8084 28116 8099 28135
rect 8169 28163 8184 28168
rect 8184 28163 8218 28168
rect 8218 28163 8221 28168
rect 8169 28125 8221 28163
rect 8169 28116 8184 28125
rect 8184 28116 8218 28125
rect 8218 28116 8221 28125
rect 5040 26714 5092 26720
rect 5040 26680 5046 26714
rect 5046 26680 5080 26714
rect 5080 26680 5092 26714
rect 5040 26668 5092 26680
rect 5106 26714 5158 26720
rect 5106 26680 5118 26714
rect 5118 26680 5152 26714
rect 5152 26680 5158 26714
rect 5106 26668 5158 26680
rect 5040 26641 5092 26651
rect 5040 26607 5046 26641
rect 5046 26607 5080 26641
rect 5080 26607 5092 26641
rect 5040 26599 5092 26607
rect 5106 26641 5158 26651
rect 5106 26607 5118 26641
rect 5118 26607 5152 26641
rect 5152 26607 5158 26641
rect 5106 26599 5158 26607
rect 5040 26568 5092 26582
rect 5040 26534 5046 26568
rect 5046 26534 5080 26568
rect 5080 26534 5092 26568
rect 5040 26530 5092 26534
rect 5106 26568 5158 26582
rect 5106 26534 5118 26568
rect 5118 26534 5152 26568
rect 5152 26534 5158 26568
rect 5106 26530 5158 26534
rect 5040 26495 5092 26513
rect 5040 26461 5046 26495
rect 5046 26461 5080 26495
rect 5080 26461 5092 26495
rect 5106 26495 5158 26513
rect 5106 26461 5118 26495
rect 5118 26461 5152 26495
rect 5152 26461 5158 26495
rect 5040 26422 5092 26444
rect 5106 26422 5158 26444
rect 5040 26392 5046 26422
rect 5046 26392 5092 26422
rect 5106 26392 5152 26422
rect 5152 26392 5158 26422
rect 5040 26323 5046 26375
rect 5046 26323 5092 26375
rect 5106 26323 5152 26375
rect 5152 26323 5158 26375
rect 5040 26254 5046 26306
rect 5046 26254 5092 26306
rect 5106 26254 5152 26306
rect 5152 26254 5158 26306
rect 5040 26184 5046 26236
rect 5046 26184 5092 26236
rect 5106 26184 5152 26236
rect 5152 26184 5158 26236
rect 5040 26114 5046 26166
rect 5046 26114 5092 26166
rect 5106 26114 5152 26166
rect 5152 26114 5158 26166
rect 5317 25930 5323 25982
rect 5323 25930 5369 25982
rect 5383 25930 5429 25982
rect 5429 25930 5435 25982
rect 5317 25861 5323 25913
rect 5323 25861 5369 25913
rect 5383 25861 5429 25913
rect 5429 25861 5435 25913
rect 5317 25792 5323 25844
rect 5323 25792 5369 25844
rect 5383 25792 5429 25844
rect 5429 25792 5435 25844
rect 5317 25723 5323 25775
rect 5323 25723 5369 25775
rect 5383 25723 5429 25775
rect 5429 25723 5435 25775
rect 5317 25654 5323 25706
rect 5323 25654 5369 25706
rect 5383 25654 5429 25706
rect 5429 25654 5435 25706
rect 5317 25584 5323 25636
rect 5323 25584 5369 25636
rect 5383 25584 5429 25636
rect 5429 25584 5435 25636
rect 5317 25514 5323 25566
rect 5323 25514 5369 25566
rect 5383 25514 5429 25566
rect 5429 25514 5435 25566
rect 5317 25444 5323 25496
rect 5323 25444 5369 25496
rect 5383 25444 5429 25496
rect 5429 25444 5435 25496
rect 5317 25380 5323 25426
rect 5323 25380 5369 25426
rect 5383 25380 5429 25426
rect 5429 25380 5435 25426
rect 5317 25374 5369 25380
rect 5383 25374 5435 25380
rect 5594 26714 5646 26720
rect 5594 26680 5600 26714
rect 5600 26680 5634 26714
rect 5634 26680 5646 26714
rect 5594 26668 5646 26680
rect 5660 26714 5712 26720
rect 5660 26680 5672 26714
rect 5672 26680 5706 26714
rect 5706 26680 5712 26714
rect 5660 26668 5712 26680
rect 5594 26641 5646 26651
rect 5594 26607 5600 26641
rect 5600 26607 5634 26641
rect 5634 26607 5646 26641
rect 5594 26599 5646 26607
rect 5660 26641 5712 26651
rect 5660 26607 5672 26641
rect 5672 26607 5706 26641
rect 5706 26607 5712 26641
rect 5660 26599 5712 26607
rect 5594 26568 5646 26582
rect 5594 26534 5600 26568
rect 5600 26534 5634 26568
rect 5634 26534 5646 26568
rect 5594 26530 5646 26534
rect 5660 26568 5712 26582
rect 5660 26534 5672 26568
rect 5672 26534 5706 26568
rect 5706 26534 5712 26568
rect 5660 26530 5712 26534
rect 5594 26495 5646 26513
rect 5594 26461 5600 26495
rect 5600 26461 5634 26495
rect 5634 26461 5646 26495
rect 5660 26495 5712 26513
rect 5660 26461 5672 26495
rect 5672 26461 5706 26495
rect 5706 26461 5712 26495
rect 5594 26422 5646 26444
rect 5660 26422 5712 26444
rect 5594 26392 5600 26422
rect 5600 26392 5646 26422
rect 5660 26392 5706 26422
rect 5706 26392 5712 26422
rect 5594 26323 5600 26375
rect 5600 26323 5646 26375
rect 5660 26323 5706 26375
rect 5706 26323 5712 26375
rect 5594 26254 5600 26306
rect 5600 26254 5646 26306
rect 5660 26254 5706 26306
rect 5706 26254 5712 26306
rect 5594 26184 5600 26236
rect 5600 26184 5646 26236
rect 5660 26184 5706 26236
rect 5706 26184 5712 26236
rect 5594 26114 5600 26166
rect 5600 26114 5646 26166
rect 5660 26114 5706 26166
rect 5706 26114 5712 26166
rect 5871 25930 5877 25982
rect 5877 25930 5923 25982
rect 5937 25930 5983 25982
rect 5983 25930 5989 25982
rect 5871 25861 5877 25913
rect 5877 25861 5923 25913
rect 5937 25861 5983 25913
rect 5983 25861 5989 25913
rect 5871 25792 5877 25844
rect 5877 25792 5923 25844
rect 5937 25792 5983 25844
rect 5983 25792 5989 25844
rect 5871 25723 5877 25775
rect 5877 25723 5923 25775
rect 5937 25723 5983 25775
rect 5983 25723 5989 25775
rect 5871 25654 5877 25706
rect 5877 25654 5923 25706
rect 5937 25654 5983 25706
rect 5983 25654 5989 25706
rect 5871 25584 5877 25636
rect 5877 25584 5923 25636
rect 5937 25584 5983 25636
rect 5983 25584 5989 25636
rect 5871 25514 5877 25566
rect 5877 25514 5923 25566
rect 5937 25514 5983 25566
rect 5983 25514 5989 25566
rect 5871 25444 5877 25496
rect 5877 25444 5923 25496
rect 5937 25444 5983 25496
rect 5983 25444 5989 25496
rect 5871 25380 5877 25426
rect 5877 25380 5923 25426
rect 5937 25380 5983 25426
rect 5983 25380 5989 25426
rect 5871 25374 5923 25380
rect 5937 25374 5989 25380
rect 6148 26714 6200 26720
rect 6148 26680 6154 26714
rect 6154 26680 6188 26714
rect 6188 26680 6200 26714
rect 6148 26668 6200 26680
rect 6214 26714 6266 26720
rect 6214 26680 6226 26714
rect 6226 26680 6260 26714
rect 6260 26680 6266 26714
rect 6214 26668 6266 26680
rect 6148 26641 6200 26651
rect 6148 26607 6154 26641
rect 6154 26607 6188 26641
rect 6188 26607 6200 26641
rect 6148 26599 6200 26607
rect 6214 26641 6266 26651
rect 6214 26607 6226 26641
rect 6226 26607 6260 26641
rect 6260 26607 6266 26641
rect 6214 26599 6266 26607
rect 6148 26568 6200 26582
rect 6148 26534 6154 26568
rect 6154 26534 6188 26568
rect 6188 26534 6200 26568
rect 6148 26530 6200 26534
rect 6214 26568 6266 26582
rect 6214 26534 6226 26568
rect 6226 26534 6260 26568
rect 6260 26534 6266 26568
rect 6214 26530 6266 26534
rect 6148 26495 6200 26513
rect 6148 26461 6154 26495
rect 6154 26461 6188 26495
rect 6188 26461 6200 26495
rect 6214 26495 6266 26513
rect 6214 26461 6226 26495
rect 6226 26461 6260 26495
rect 6260 26461 6266 26495
rect 6148 26422 6200 26444
rect 6214 26422 6266 26444
rect 6148 26392 6154 26422
rect 6154 26392 6200 26422
rect 6214 26392 6260 26422
rect 6260 26392 6266 26422
rect 6148 26323 6154 26375
rect 6154 26323 6200 26375
rect 6214 26323 6260 26375
rect 6260 26323 6266 26375
rect 6148 26254 6154 26306
rect 6154 26254 6200 26306
rect 6214 26254 6260 26306
rect 6260 26254 6266 26306
rect 6148 26184 6154 26236
rect 6154 26184 6200 26236
rect 6214 26184 6260 26236
rect 6260 26184 6266 26236
rect 6148 26114 6154 26166
rect 6154 26114 6200 26166
rect 6214 26114 6260 26166
rect 6260 26114 6266 26166
rect 6425 25930 6431 25982
rect 6431 25930 6477 25982
rect 6491 25930 6537 25982
rect 6537 25930 6543 25982
rect 6425 25861 6431 25913
rect 6431 25861 6477 25913
rect 6491 25861 6537 25913
rect 6537 25861 6543 25913
rect 6425 25792 6431 25844
rect 6431 25792 6477 25844
rect 6491 25792 6537 25844
rect 6537 25792 6543 25844
rect 6425 25723 6431 25775
rect 6431 25723 6477 25775
rect 6491 25723 6537 25775
rect 6537 25723 6543 25775
rect 6425 25654 6431 25706
rect 6431 25654 6477 25706
rect 6491 25654 6537 25706
rect 6537 25654 6543 25706
rect 6425 25584 6431 25636
rect 6431 25584 6477 25636
rect 6491 25584 6537 25636
rect 6537 25584 6543 25636
rect 6425 25514 6431 25566
rect 6431 25514 6477 25566
rect 6491 25514 6537 25566
rect 6537 25514 6543 25566
rect 6425 25444 6431 25496
rect 6431 25444 6477 25496
rect 6491 25444 6537 25496
rect 6537 25444 6543 25496
rect 6425 25380 6431 25426
rect 6431 25380 6477 25426
rect 6491 25380 6537 25426
rect 6537 25380 6543 25426
rect 6425 25374 6477 25380
rect 6491 25374 6543 25380
rect 6702 26714 6754 26720
rect 6702 26680 6708 26714
rect 6708 26680 6742 26714
rect 6742 26680 6754 26714
rect 6702 26668 6754 26680
rect 6768 26714 6820 26720
rect 6768 26680 6780 26714
rect 6780 26680 6814 26714
rect 6814 26680 6820 26714
rect 6768 26668 6820 26680
rect 6702 26641 6754 26651
rect 6702 26607 6708 26641
rect 6708 26607 6742 26641
rect 6742 26607 6754 26641
rect 6702 26599 6754 26607
rect 6768 26641 6820 26651
rect 6768 26607 6780 26641
rect 6780 26607 6814 26641
rect 6814 26607 6820 26641
rect 6768 26599 6820 26607
rect 6702 26568 6754 26582
rect 6702 26534 6708 26568
rect 6708 26534 6742 26568
rect 6742 26534 6754 26568
rect 6702 26530 6754 26534
rect 6768 26568 6820 26582
rect 6768 26534 6780 26568
rect 6780 26534 6814 26568
rect 6814 26534 6820 26568
rect 6768 26530 6820 26534
rect 6702 26495 6754 26513
rect 6702 26461 6708 26495
rect 6708 26461 6742 26495
rect 6742 26461 6754 26495
rect 6768 26495 6820 26513
rect 6768 26461 6780 26495
rect 6780 26461 6814 26495
rect 6814 26461 6820 26495
rect 6702 26422 6754 26444
rect 6768 26422 6820 26444
rect 6702 26392 6708 26422
rect 6708 26392 6754 26422
rect 6768 26392 6814 26422
rect 6814 26392 6820 26422
rect 6702 26323 6708 26375
rect 6708 26323 6754 26375
rect 6768 26323 6814 26375
rect 6814 26323 6820 26375
rect 6702 26254 6708 26306
rect 6708 26254 6754 26306
rect 6768 26254 6814 26306
rect 6814 26254 6820 26306
rect 6702 26184 6708 26236
rect 6708 26184 6754 26236
rect 6768 26184 6814 26236
rect 6814 26184 6820 26236
rect 6702 26114 6708 26166
rect 6708 26114 6754 26166
rect 6768 26114 6814 26166
rect 6814 26114 6820 26166
rect 6979 25930 6985 25982
rect 6985 25930 7031 25982
rect 7045 25930 7091 25982
rect 7091 25930 7097 25982
rect 6979 25861 6985 25913
rect 6985 25861 7031 25913
rect 7045 25861 7091 25913
rect 7091 25861 7097 25913
rect 6979 25792 6985 25844
rect 6985 25792 7031 25844
rect 7045 25792 7091 25844
rect 7091 25792 7097 25844
rect 6979 25723 6985 25775
rect 6985 25723 7031 25775
rect 7045 25723 7091 25775
rect 7091 25723 7097 25775
rect 6979 25654 6985 25706
rect 6985 25654 7031 25706
rect 7045 25654 7091 25706
rect 7091 25654 7097 25706
rect 6979 25584 6985 25636
rect 6985 25584 7031 25636
rect 7045 25584 7091 25636
rect 7091 25584 7097 25636
rect 6979 25514 6985 25566
rect 6985 25514 7031 25566
rect 7045 25514 7091 25566
rect 7091 25514 7097 25566
rect 6979 25444 6985 25496
rect 6985 25444 7031 25496
rect 7045 25444 7091 25496
rect 7091 25444 7097 25496
rect 6979 25380 6985 25426
rect 6985 25380 7031 25426
rect 7045 25380 7091 25426
rect 7091 25380 7097 25426
rect 6979 25374 7031 25380
rect 7045 25374 7097 25380
rect 7256 26714 7308 26720
rect 7256 26680 7262 26714
rect 7262 26680 7296 26714
rect 7296 26680 7308 26714
rect 7256 26668 7308 26680
rect 7322 26714 7374 26720
rect 7322 26680 7334 26714
rect 7334 26680 7368 26714
rect 7368 26680 7374 26714
rect 7322 26668 7374 26680
rect 7256 26641 7308 26651
rect 7256 26607 7262 26641
rect 7262 26607 7296 26641
rect 7296 26607 7308 26641
rect 7256 26599 7308 26607
rect 7322 26641 7374 26651
rect 7322 26607 7334 26641
rect 7334 26607 7368 26641
rect 7368 26607 7374 26641
rect 7322 26599 7374 26607
rect 7256 26568 7308 26582
rect 7256 26534 7262 26568
rect 7262 26534 7296 26568
rect 7296 26534 7308 26568
rect 7256 26530 7308 26534
rect 7322 26568 7374 26582
rect 7322 26534 7334 26568
rect 7334 26534 7368 26568
rect 7368 26534 7374 26568
rect 7322 26530 7374 26534
rect 7256 26495 7308 26513
rect 7256 26461 7262 26495
rect 7262 26461 7296 26495
rect 7296 26461 7308 26495
rect 7322 26495 7374 26513
rect 7322 26461 7334 26495
rect 7334 26461 7368 26495
rect 7368 26461 7374 26495
rect 7256 26422 7308 26444
rect 7322 26422 7374 26444
rect 7256 26392 7262 26422
rect 7262 26392 7308 26422
rect 7322 26392 7368 26422
rect 7368 26392 7374 26422
rect 7256 26323 7262 26375
rect 7262 26323 7308 26375
rect 7322 26323 7368 26375
rect 7368 26323 7374 26375
rect 7256 26254 7262 26306
rect 7262 26254 7308 26306
rect 7322 26254 7368 26306
rect 7368 26254 7374 26306
rect 7256 26184 7262 26236
rect 7262 26184 7308 26236
rect 7322 26184 7368 26236
rect 7368 26184 7374 26236
rect 7256 26114 7262 26166
rect 7262 26114 7308 26166
rect 7322 26114 7368 26166
rect 7368 26114 7374 26166
rect 7533 25930 7539 25982
rect 7539 25930 7585 25982
rect 7599 25930 7645 25982
rect 7645 25930 7651 25982
rect 7533 25861 7539 25913
rect 7539 25861 7585 25913
rect 7599 25861 7645 25913
rect 7645 25861 7651 25913
rect 7533 25792 7539 25844
rect 7539 25792 7585 25844
rect 7599 25792 7645 25844
rect 7645 25792 7651 25844
rect 7533 25723 7539 25775
rect 7539 25723 7585 25775
rect 7599 25723 7645 25775
rect 7645 25723 7651 25775
rect 7533 25654 7539 25706
rect 7539 25654 7585 25706
rect 7599 25654 7645 25706
rect 7645 25654 7651 25706
rect 7533 25584 7539 25636
rect 7539 25584 7585 25636
rect 7599 25584 7645 25636
rect 7645 25584 7651 25636
rect 7533 25514 7539 25566
rect 7539 25514 7585 25566
rect 7599 25514 7645 25566
rect 7645 25514 7651 25566
rect 7533 25444 7539 25496
rect 7539 25444 7585 25496
rect 7599 25444 7645 25496
rect 7645 25444 7651 25496
rect 7533 25380 7539 25426
rect 7539 25380 7585 25426
rect 7599 25380 7645 25426
rect 7645 25380 7651 25426
rect 7533 25374 7585 25380
rect 7599 25374 7651 25380
rect 7810 26714 7862 26720
rect 7810 26680 7816 26714
rect 7816 26680 7850 26714
rect 7850 26680 7862 26714
rect 7810 26668 7862 26680
rect 7876 26714 7928 26720
rect 7876 26680 7888 26714
rect 7888 26680 7922 26714
rect 7922 26680 7928 26714
rect 7876 26668 7928 26680
rect 7810 26641 7862 26651
rect 7810 26607 7816 26641
rect 7816 26607 7850 26641
rect 7850 26607 7862 26641
rect 7810 26599 7862 26607
rect 7876 26641 7928 26651
rect 7876 26607 7888 26641
rect 7888 26607 7922 26641
rect 7922 26607 7928 26641
rect 7876 26599 7928 26607
rect 7810 26568 7862 26582
rect 7810 26534 7816 26568
rect 7816 26534 7850 26568
rect 7850 26534 7862 26568
rect 7810 26530 7862 26534
rect 7876 26568 7928 26582
rect 7876 26534 7888 26568
rect 7888 26534 7922 26568
rect 7922 26534 7928 26568
rect 7876 26530 7928 26534
rect 7810 26495 7862 26513
rect 7810 26461 7816 26495
rect 7816 26461 7850 26495
rect 7850 26461 7862 26495
rect 7876 26495 7928 26513
rect 7876 26461 7888 26495
rect 7888 26461 7922 26495
rect 7922 26461 7928 26495
rect 7810 26422 7862 26444
rect 7876 26422 7928 26444
rect 7810 26392 7816 26422
rect 7816 26392 7862 26422
rect 7876 26392 7922 26422
rect 7922 26392 7928 26422
rect 7810 26323 7816 26375
rect 7816 26323 7862 26375
rect 7876 26323 7922 26375
rect 7922 26323 7928 26375
rect 7810 26254 7816 26306
rect 7816 26254 7862 26306
rect 7876 26254 7922 26306
rect 7922 26254 7928 26306
rect 7810 26184 7816 26236
rect 7816 26184 7862 26236
rect 7876 26184 7922 26236
rect 7922 26184 7928 26236
rect 7810 26114 7816 26166
rect 7816 26114 7862 26166
rect 7876 26114 7922 26166
rect 7922 26114 7928 26166
rect 8047 26695 8099 26724
rect 8047 26672 8050 26695
rect 8050 26672 8084 26695
rect 8084 26672 8099 26695
rect 8169 26723 8184 26724
rect 8184 26723 8218 26724
rect 8218 26723 8221 26724
rect 8169 26685 8221 26723
rect 8169 26672 8184 26685
rect 8184 26672 8218 26685
rect 8218 26672 8221 26685
rect 8047 26623 8099 26655
rect 8047 26603 8050 26623
rect 8050 26603 8084 26623
rect 8084 26603 8099 26623
rect 8169 26651 8184 26655
rect 8184 26651 8218 26655
rect 8218 26651 8221 26655
rect 8169 26613 8221 26651
rect 8169 26603 8184 26613
rect 8184 26603 8218 26613
rect 8218 26603 8221 26613
rect 8047 26551 8099 26586
rect 8047 26534 8050 26551
rect 8050 26534 8084 26551
rect 8084 26534 8099 26551
rect 8169 26579 8184 26586
rect 8184 26579 8218 26586
rect 8218 26579 8221 26586
rect 8169 26541 8221 26579
rect 8169 26534 8184 26541
rect 8184 26534 8218 26541
rect 8218 26534 8221 26541
rect 8047 26479 8099 26517
rect 8047 26465 8050 26479
rect 8050 26465 8084 26479
rect 8084 26465 8099 26479
rect 8169 26507 8184 26517
rect 8184 26507 8218 26517
rect 8218 26507 8221 26517
rect 8169 26469 8221 26507
rect 8169 26465 8184 26469
rect 8184 26465 8218 26469
rect 8218 26465 8221 26469
rect 8047 26445 8050 26448
rect 8050 26445 8084 26448
rect 8084 26445 8099 26448
rect 8047 26407 8099 26445
rect 8047 26396 8050 26407
rect 8050 26396 8084 26407
rect 8084 26396 8099 26407
rect 8169 26435 8184 26448
rect 8184 26435 8218 26448
rect 8218 26435 8221 26448
rect 8169 26397 8221 26435
rect 8169 26396 8184 26397
rect 8184 26396 8218 26397
rect 8218 26396 8221 26397
rect 8047 26373 8050 26378
rect 8050 26373 8084 26378
rect 8084 26373 8099 26378
rect 8047 26335 8099 26373
rect 8047 26326 8050 26335
rect 8050 26326 8084 26335
rect 8084 26326 8099 26335
rect 8169 26363 8184 26378
rect 8184 26363 8218 26378
rect 8218 26363 8221 26378
rect 8169 26326 8221 26363
rect 8047 26301 8050 26308
rect 8050 26301 8084 26308
rect 8084 26301 8099 26308
rect 8047 26263 8099 26301
rect 8047 26256 8050 26263
rect 8050 26256 8084 26263
rect 8084 26256 8099 26263
rect 8169 26291 8184 26308
rect 8184 26291 8218 26308
rect 8218 26291 8221 26308
rect 8169 26256 8221 26291
rect 8047 26229 8050 26238
rect 8050 26229 8084 26238
rect 8084 26229 8099 26238
rect 8047 26191 8099 26229
rect 8047 26186 8050 26191
rect 8050 26186 8084 26191
rect 8084 26186 8099 26191
rect 8169 26219 8184 26238
rect 8184 26219 8218 26238
rect 8218 26219 8221 26238
rect 8169 26186 8221 26219
rect 8047 26157 8050 26168
rect 8050 26157 8084 26168
rect 8084 26157 8099 26168
rect 8047 26119 8099 26157
rect 8047 26116 8050 26119
rect 8050 26116 8084 26119
rect 8084 26116 8099 26119
rect 8169 26147 8184 26168
rect 8184 26147 8218 26168
rect 8218 26147 8221 26168
rect 8169 26116 8221 26147
rect 5040 24714 5092 24720
rect 5040 24680 5046 24714
rect 5046 24680 5080 24714
rect 5080 24680 5092 24714
rect 5040 24668 5092 24680
rect 5106 24714 5158 24720
rect 5106 24680 5118 24714
rect 5118 24680 5152 24714
rect 5152 24680 5158 24714
rect 5106 24668 5158 24680
rect 5040 24641 5092 24651
rect 5040 24607 5046 24641
rect 5046 24607 5080 24641
rect 5080 24607 5092 24641
rect 5040 24599 5092 24607
rect 5106 24641 5158 24651
rect 5106 24607 5118 24641
rect 5118 24607 5152 24641
rect 5152 24607 5158 24641
rect 5106 24599 5158 24607
rect 5040 24568 5092 24582
rect 5040 24534 5046 24568
rect 5046 24534 5080 24568
rect 5080 24534 5092 24568
rect 5040 24530 5092 24534
rect 5106 24568 5158 24582
rect 5106 24534 5118 24568
rect 5118 24534 5152 24568
rect 5152 24534 5158 24568
rect 5106 24530 5158 24534
rect 5040 24495 5092 24513
rect 5040 24461 5046 24495
rect 5046 24461 5080 24495
rect 5080 24461 5092 24495
rect 5106 24495 5158 24513
rect 5106 24461 5118 24495
rect 5118 24461 5152 24495
rect 5152 24461 5158 24495
rect 5040 24422 5092 24444
rect 5106 24422 5158 24444
rect 5040 24392 5046 24422
rect 5046 24392 5092 24422
rect 5106 24392 5152 24422
rect 5152 24392 5158 24422
rect 5040 24323 5046 24375
rect 5046 24323 5092 24375
rect 5106 24323 5152 24375
rect 5152 24323 5158 24375
rect 5040 24254 5046 24306
rect 5046 24254 5092 24306
rect 5106 24254 5152 24306
rect 5152 24254 5158 24306
rect 5040 24184 5046 24236
rect 5046 24184 5092 24236
rect 5106 24184 5152 24236
rect 5152 24184 5158 24236
rect 5040 24114 5046 24166
rect 5046 24114 5092 24166
rect 5106 24114 5152 24166
rect 5152 24114 5158 24166
rect 5317 23930 5323 23982
rect 5323 23930 5369 23982
rect 5383 23930 5429 23982
rect 5429 23930 5435 23982
rect 5317 23861 5323 23913
rect 5323 23861 5369 23913
rect 5383 23861 5429 23913
rect 5429 23861 5435 23913
rect 5317 23792 5323 23844
rect 5323 23792 5369 23844
rect 5383 23792 5429 23844
rect 5429 23792 5435 23844
rect 5317 23723 5323 23775
rect 5323 23723 5369 23775
rect 5383 23723 5429 23775
rect 5429 23723 5435 23775
rect 5317 23654 5323 23706
rect 5323 23654 5369 23706
rect 5383 23654 5429 23706
rect 5429 23654 5435 23706
rect 5317 23584 5323 23636
rect 5323 23584 5369 23636
rect 5383 23584 5429 23636
rect 5429 23584 5435 23636
rect 5317 23514 5323 23566
rect 5323 23514 5369 23566
rect 5383 23514 5429 23566
rect 5429 23514 5435 23566
rect 5317 23444 5323 23496
rect 5323 23444 5369 23496
rect 5383 23444 5429 23496
rect 5429 23444 5435 23496
rect 5317 23380 5323 23426
rect 5323 23380 5369 23426
rect 5383 23380 5429 23426
rect 5429 23380 5435 23426
rect 5317 23374 5369 23380
rect 5383 23374 5435 23380
rect 5594 24714 5646 24720
rect 5594 24680 5600 24714
rect 5600 24680 5634 24714
rect 5634 24680 5646 24714
rect 5594 24668 5646 24680
rect 5660 24714 5712 24720
rect 5660 24680 5672 24714
rect 5672 24680 5706 24714
rect 5706 24680 5712 24714
rect 5660 24668 5712 24680
rect 5594 24641 5646 24651
rect 5594 24607 5600 24641
rect 5600 24607 5634 24641
rect 5634 24607 5646 24641
rect 5594 24599 5646 24607
rect 5660 24641 5712 24651
rect 5660 24607 5672 24641
rect 5672 24607 5706 24641
rect 5706 24607 5712 24641
rect 5660 24599 5712 24607
rect 5594 24568 5646 24582
rect 5594 24534 5600 24568
rect 5600 24534 5634 24568
rect 5634 24534 5646 24568
rect 5594 24530 5646 24534
rect 5660 24568 5712 24582
rect 5660 24534 5672 24568
rect 5672 24534 5706 24568
rect 5706 24534 5712 24568
rect 5660 24530 5712 24534
rect 5594 24495 5646 24513
rect 5594 24461 5600 24495
rect 5600 24461 5634 24495
rect 5634 24461 5646 24495
rect 5660 24495 5712 24513
rect 5660 24461 5672 24495
rect 5672 24461 5706 24495
rect 5706 24461 5712 24495
rect 5594 24422 5646 24444
rect 5660 24422 5712 24444
rect 5594 24392 5600 24422
rect 5600 24392 5646 24422
rect 5660 24392 5706 24422
rect 5706 24392 5712 24422
rect 5594 24323 5600 24375
rect 5600 24323 5646 24375
rect 5660 24323 5706 24375
rect 5706 24323 5712 24375
rect 5594 24254 5600 24306
rect 5600 24254 5646 24306
rect 5660 24254 5706 24306
rect 5706 24254 5712 24306
rect 5594 24184 5600 24236
rect 5600 24184 5646 24236
rect 5660 24184 5706 24236
rect 5706 24184 5712 24236
rect 5594 24114 5600 24166
rect 5600 24114 5646 24166
rect 5660 24114 5706 24166
rect 5706 24114 5712 24166
rect 5871 23930 5877 23982
rect 5877 23930 5923 23982
rect 5937 23930 5983 23982
rect 5983 23930 5989 23982
rect 5871 23861 5877 23913
rect 5877 23861 5923 23913
rect 5937 23861 5983 23913
rect 5983 23861 5989 23913
rect 5871 23792 5877 23844
rect 5877 23792 5923 23844
rect 5937 23792 5983 23844
rect 5983 23792 5989 23844
rect 5871 23723 5877 23775
rect 5877 23723 5923 23775
rect 5937 23723 5983 23775
rect 5983 23723 5989 23775
rect 5871 23654 5877 23706
rect 5877 23654 5923 23706
rect 5937 23654 5983 23706
rect 5983 23654 5989 23706
rect 5871 23584 5877 23636
rect 5877 23584 5923 23636
rect 5937 23584 5983 23636
rect 5983 23584 5989 23636
rect 5871 23514 5877 23566
rect 5877 23514 5923 23566
rect 5937 23514 5983 23566
rect 5983 23514 5989 23566
rect 5871 23444 5877 23496
rect 5877 23444 5923 23496
rect 5937 23444 5983 23496
rect 5983 23444 5989 23496
rect 5871 23380 5877 23426
rect 5877 23380 5923 23426
rect 5937 23380 5983 23426
rect 5983 23380 5989 23426
rect 5871 23374 5923 23380
rect 5937 23374 5989 23380
rect 6148 24714 6200 24720
rect 6148 24680 6154 24714
rect 6154 24680 6188 24714
rect 6188 24680 6200 24714
rect 6148 24668 6200 24680
rect 6214 24714 6266 24720
rect 6214 24680 6226 24714
rect 6226 24680 6260 24714
rect 6260 24680 6266 24714
rect 6214 24668 6266 24680
rect 6148 24641 6200 24651
rect 6148 24607 6154 24641
rect 6154 24607 6188 24641
rect 6188 24607 6200 24641
rect 6148 24599 6200 24607
rect 6214 24641 6266 24651
rect 6214 24607 6226 24641
rect 6226 24607 6260 24641
rect 6260 24607 6266 24641
rect 6214 24599 6266 24607
rect 6148 24568 6200 24582
rect 6148 24534 6154 24568
rect 6154 24534 6188 24568
rect 6188 24534 6200 24568
rect 6148 24530 6200 24534
rect 6214 24568 6266 24582
rect 6214 24534 6226 24568
rect 6226 24534 6260 24568
rect 6260 24534 6266 24568
rect 6214 24530 6266 24534
rect 6148 24495 6200 24513
rect 6148 24461 6154 24495
rect 6154 24461 6188 24495
rect 6188 24461 6200 24495
rect 6214 24495 6266 24513
rect 6214 24461 6226 24495
rect 6226 24461 6260 24495
rect 6260 24461 6266 24495
rect 6148 24422 6200 24444
rect 6214 24422 6266 24444
rect 6148 24392 6154 24422
rect 6154 24392 6200 24422
rect 6214 24392 6260 24422
rect 6260 24392 6266 24422
rect 6148 24323 6154 24375
rect 6154 24323 6200 24375
rect 6214 24323 6260 24375
rect 6260 24323 6266 24375
rect 6148 24254 6154 24306
rect 6154 24254 6200 24306
rect 6214 24254 6260 24306
rect 6260 24254 6266 24306
rect 6148 24184 6154 24236
rect 6154 24184 6200 24236
rect 6214 24184 6260 24236
rect 6260 24184 6266 24236
rect 6148 24114 6154 24166
rect 6154 24114 6200 24166
rect 6214 24114 6260 24166
rect 6260 24114 6266 24166
rect 6425 23930 6431 23982
rect 6431 23930 6477 23982
rect 6491 23930 6537 23982
rect 6537 23930 6543 23982
rect 6425 23861 6431 23913
rect 6431 23861 6477 23913
rect 6491 23861 6537 23913
rect 6537 23861 6543 23913
rect 6425 23792 6431 23844
rect 6431 23792 6477 23844
rect 6491 23792 6537 23844
rect 6537 23792 6543 23844
rect 6425 23723 6431 23775
rect 6431 23723 6477 23775
rect 6491 23723 6537 23775
rect 6537 23723 6543 23775
rect 6425 23654 6431 23706
rect 6431 23654 6477 23706
rect 6491 23654 6537 23706
rect 6537 23654 6543 23706
rect 6425 23584 6431 23636
rect 6431 23584 6477 23636
rect 6491 23584 6537 23636
rect 6537 23584 6543 23636
rect 6425 23514 6431 23566
rect 6431 23514 6477 23566
rect 6491 23514 6537 23566
rect 6537 23514 6543 23566
rect 6425 23444 6431 23496
rect 6431 23444 6477 23496
rect 6491 23444 6537 23496
rect 6537 23444 6543 23496
rect 6425 23380 6431 23426
rect 6431 23380 6477 23426
rect 6491 23380 6537 23426
rect 6537 23380 6543 23426
rect 6425 23374 6477 23380
rect 6491 23374 6543 23380
rect 6702 24714 6754 24720
rect 6702 24680 6708 24714
rect 6708 24680 6742 24714
rect 6742 24680 6754 24714
rect 6702 24668 6754 24680
rect 6768 24714 6820 24720
rect 6768 24680 6780 24714
rect 6780 24680 6814 24714
rect 6814 24680 6820 24714
rect 6768 24668 6820 24680
rect 6702 24641 6754 24651
rect 6702 24607 6708 24641
rect 6708 24607 6742 24641
rect 6742 24607 6754 24641
rect 6702 24599 6754 24607
rect 6768 24641 6820 24651
rect 6768 24607 6780 24641
rect 6780 24607 6814 24641
rect 6814 24607 6820 24641
rect 6768 24599 6820 24607
rect 6702 24568 6754 24582
rect 6702 24534 6708 24568
rect 6708 24534 6742 24568
rect 6742 24534 6754 24568
rect 6702 24530 6754 24534
rect 6768 24568 6820 24582
rect 6768 24534 6780 24568
rect 6780 24534 6814 24568
rect 6814 24534 6820 24568
rect 6768 24530 6820 24534
rect 6702 24495 6754 24513
rect 6702 24461 6708 24495
rect 6708 24461 6742 24495
rect 6742 24461 6754 24495
rect 6768 24495 6820 24513
rect 6768 24461 6780 24495
rect 6780 24461 6814 24495
rect 6814 24461 6820 24495
rect 6702 24422 6754 24444
rect 6768 24422 6820 24444
rect 6702 24392 6708 24422
rect 6708 24392 6754 24422
rect 6768 24392 6814 24422
rect 6814 24392 6820 24422
rect 6702 24323 6708 24375
rect 6708 24323 6754 24375
rect 6768 24323 6814 24375
rect 6814 24323 6820 24375
rect 6702 24254 6708 24306
rect 6708 24254 6754 24306
rect 6768 24254 6814 24306
rect 6814 24254 6820 24306
rect 6702 24184 6708 24236
rect 6708 24184 6754 24236
rect 6768 24184 6814 24236
rect 6814 24184 6820 24236
rect 6702 24114 6708 24166
rect 6708 24114 6754 24166
rect 6768 24114 6814 24166
rect 6814 24114 6820 24166
rect 6979 23930 6985 23982
rect 6985 23930 7031 23982
rect 7045 23930 7091 23982
rect 7091 23930 7097 23982
rect 6979 23861 6985 23913
rect 6985 23861 7031 23913
rect 7045 23861 7091 23913
rect 7091 23861 7097 23913
rect 6979 23792 6985 23844
rect 6985 23792 7031 23844
rect 7045 23792 7091 23844
rect 7091 23792 7097 23844
rect 6979 23723 6985 23775
rect 6985 23723 7031 23775
rect 7045 23723 7091 23775
rect 7091 23723 7097 23775
rect 6979 23654 6985 23706
rect 6985 23654 7031 23706
rect 7045 23654 7091 23706
rect 7091 23654 7097 23706
rect 6979 23584 6985 23636
rect 6985 23584 7031 23636
rect 7045 23584 7091 23636
rect 7091 23584 7097 23636
rect 6979 23514 6985 23566
rect 6985 23514 7031 23566
rect 7045 23514 7091 23566
rect 7091 23514 7097 23566
rect 6979 23444 6985 23496
rect 6985 23444 7031 23496
rect 7045 23444 7091 23496
rect 7091 23444 7097 23496
rect 6979 23380 6985 23426
rect 6985 23380 7031 23426
rect 7045 23380 7091 23426
rect 7091 23380 7097 23426
rect 6979 23374 7031 23380
rect 7045 23374 7097 23380
rect 7256 24714 7308 24720
rect 7256 24680 7262 24714
rect 7262 24680 7296 24714
rect 7296 24680 7308 24714
rect 7256 24668 7308 24680
rect 7322 24714 7374 24720
rect 7322 24680 7334 24714
rect 7334 24680 7368 24714
rect 7368 24680 7374 24714
rect 7322 24668 7374 24680
rect 7256 24641 7308 24651
rect 7256 24607 7262 24641
rect 7262 24607 7296 24641
rect 7296 24607 7308 24641
rect 7256 24599 7308 24607
rect 7322 24641 7374 24651
rect 7322 24607 7334 24641
rect 7334 24607 7368 24641
rect 7368 24607 7374 24641
rect 7322 24599 7374 24607
rect 7256 24568 7308 24582
rect 7256 24534 7262 24568
rect 7262 24534 7296 24568
rect 7296 24534 7308 24568
rect 7256 24530 7308 24534
rect 7322 24568 7374 24582
rect 7322 24534 7334 24568
rect 7334 24534 7368 24568
rect 7368 24534 7374 24568
rect 7322 24530 7374 24534
rect 7256 24495 7308 24513
rect 7256 24461 7262 24495
rect 7262 24461 7296 24495
rect 7296 24461 7308 24495
rect 7322 24495 7374 24513
rect 7322 24461 7334 24495
rect 7334 24461 7368 24495
rect 7368 24461 7374 24495
rect 7256 24422 7308 24444
rect 7322 24422 7374 24444
rect 7256 24392 7262 24422
rect 7262 24392 7308 24422
rect 7322 24392 7368 24422
rect 7368 24392 7374 24422
rect 7256 24323 7262 24375
rect 7262 24323 7308 24375
rect 7322 24323 7368 24375
rect 7368 24323 7374 24375
rect 7256 24254 7262 24306
rect 7262 24254 7308 24306
rect 7322 24254 7368 24306
rect 7368 24254 7374 24306
rect 7256 24184 7262 24236
rect 7262 24184 7308 24236
rect 7322 24184 7368 24236
rect 7368 24184 7374 24236
rect 7256 24114 7262 24166
rect 7262 24114 7308 24166
rect 7322 24114 7368 24166
rect 7368 24114 7374 24166
rect 7533 23930 7539 23982
rect 7539 23930 7585 23982
rect 7599 23930 7645 23982
rect 7645 23930 7651 23982
rect 7533 23861 7539 23913
rect 7539 23861 7585 23913
rect 7599 23861 7645 23913
rect 7645 23861 7651 23913
rect 7533 23792 7539 23844
rect 7539 23792 7585 23844
rect 7599 23792 7645 23844
rect 7645 23792 7651 23844
rect 7533 23723 7539 23775
rect 7539 23723 7585 23775
rect 7599 23723 7645 23775
rect 7645 23723 7651 23775
rect 7533 23654 7539 23706
rect 7539 23654 7585 23706
rect 7599 23654 7645 23706
rect 7645 23654 7651 23706
rect 7533 23584 7539 23636
rect 7539 23584 7585 23636
rect 7599 23584 7645 23636
rect 7645 23584 7651 23636
rect 7533 23514 7539 23566
rect 7539 23514 7585 23566
rect 7599 23514 7645 23566
rect 7645 23514 7651 23566
rect 7533 23444 7539 23496
rect 7539 23444 7585 23496
rect 7599 23444 7645 23496
rect 7645 23444 7651 23496
rect 7533 23380 7539 23426
rect 7539 23380 7585 23426
rect 7599 23380 7645 23426
rect 7645 23380 7651 23426
rect 7533 23374 7585 23380
rect 7599 23374 7651 23380
rect 7810 24714 7862 24720
rect 7810 24680 7816 24714
rect 7816 24680 7850 24714
rect 7850 24680 7862 24714
rect 7810 24668 7862 24680
rect 7876 24714 7928 24720
rect 7876 24680 7888 24714
rect 7888 24680 7922 24714
rect 7922 24680 7928 24714
rect 7876 24668 7928 24680
rect 7810 24641 7862 24651
rect 7810 24607 7816 24641
rect 7816 24607 7850 24641
rect 7850 24607 7862 24641
rect 7810 24599 7862 24607
rect 7876 24641 7928 24651
rect 7876 24607 7888 24641
rect 7888 24607 7922 24641
rect 7922 24607 7928 24641
rect 7876 24599 7928 24607
rect 7810 24568 7862 24582
rect 7810 24534 7816 24568
rect 7816 24534 7850 24568
rect 7850 24534 7862 24568
rect 7810 24530 7862 24534
rect 7876 24568 7928 24582
rect 7876 24534 7888 24568
rect 7888 24534 7922 24568
rect 7922 24534 7928 24568
rect 7876 24530 7928 24534
rect 7810 24495 7862 24513
rect 7810 24461 7816 24495
rect 7816 24461 7850 24495
rect 7850 24461 7862 24495
rect 7876 24495 7928 24513
rect 7876 24461 7888 24495
rect 7888 24461 7922 24495
rect 7922 24461 7928 24495
rect 7810 24422 7862 24444
rect 7876 24422 7928 24444
rect 7810 24392 7816 24422
rect 7816 24392 7862 24422
rect 7876 24392 7922 24422
rect 7922 24392 7928 24422
rect 7810 24323 7816 24375
rect 7816 24323 7862 24375
rect 7876 24323 7922 24375
rect 7922 24323 7928 24375
rect 7810 24254 7816 24306
rect 7816 24254 7862 24306
rect 7876 24254 7922 24306
rect 7922 24254 7928 24306
rect 7810 24184 7816 24236
rect 7816 24184 7862 24236
rect 7876 24184 7922 24236
rect 7922 24184 7928 24236
rect 7810 24114 7816 24166
rect 7816 24114 7862 24166
rect 7876 24114 7922 24166
rect 7922 24114 7928 24166
rect 8047 24717 8050 24724
rect 8050 24717 8084 24724
rect 8084 24717 8099 24724
rect 8047 24679 8099 24717
rect 8047 24672 8050 24679
rect 8050 24672 8084 24679
rect 8084 24672 8099 24679
rect 8169 24707 8184 24724
rect 8184 24707 8218 24724
rect 8218 24707 8221 24724
rect 8169 24672 8221 24707
rect 8047 24645 8050 24655
rect 8050 24645 8084 24655
rect 8084 24645 8099 24655
rect 8047 24607 8099 24645
rect 8047 24603 8050 24607
rect 8050 24603 8084 24607
rect 8084 24603 8099 24607
rect 8169 24635 8184 24655
rect 8184 24635 8218 24655
rect 8218 24635 8221 24655
rect 8169 24603 8221 24635
rect 8047 24573 8050 24586
rect 8050 24573 8084 24586
rect 8084 24573 8099 24586
rect 8047 24535 8099 24573
rect 8047 24534 8050 24535
rect 8050 24534 8084 24535
rect 8084 24534 8099 24535
rect 8169 24563 8184 24586
rect 8184 24563 8218 24586
rect 8218 24563 8221 24586
rect 8169 24534 8221 24563
rect 8047 24501 8050 24517
rect 8050 24501 8084 24517
rect 8084 24501 8099 24517
rect 8047 24465 8099 24501
rect 8169 24491 8184 24517
rect 8184 24491 8218 24517
rect 8218 24491 8221 24517
rect 8169 24465 8221 24491
rect 8047 24429 8050 24448
rect 8050 24429 8084 24448
rect 8084 24429 8099 24448
rect 8047 24396 8099 24429
rect 8169 24419 8184 24448
rect 8184 24419 8218 24448
rect 8218 24419 8221 24448
rect 8169 24396 8221 24419
rect 8047 24357 8050 24378
rect 8050 24357 8084 24378
rect 8084 24357 8099 24378
rect 8047 24326 8099 24357
rect 8169 24347 8184 24378
rect 8184 24347 8218 24378
rect 8218 24347 8221 24378
rect 8169 24326 8221 24347
rect 8047 24285 8050 24308
rect 8050 24285 8084 24308
rect 8084 24285 8099 24308
rect 8047 24256 8099 24285
rect 8169 24275 8184 24308
rect 8184 24275 8218 24308
rect 8218 24275 8221 24308
rect 8169 24256 8221 24275
rect 8047 24213 8050 24238
rect 8050 24213 8084 24238
rect 8084 24213 8099 24238
rect 8047 24186 8099 24213
rect 8169 24237 8221 24238
rect 8169 24203 8184 24237
rect 8184 24203 8218 24237
rect 8218 24203 8221 24237
rect 8169 24186 8221 24203
rect 8047 24141 8050 24168
rect 8050 24141 8084 24168
rect 8084 24141 8099 24168
rect 8047 24116 8099 24141
rect 8169 24165 8221 24168
rect 8169 24131 8184 24165
rect 8184 24131 8218 24165
rect 8218 24131 8221 24165
rect 8169 24116 8221 24131
rect 5040 22714 5092 22720
rect 5040 22680 5046 22714
rect 5046 22680 5080 22714
rect 5080 22680 5092 22714
rect 5040 22668 5092 22680
rect 5106 22714 5158 22720
rect 5106 22680 5118 22714
rect 5118 22680 5152 22714
rect 5152 22680 5158 22714
rect 5106 22668 5158 22680
rect 5040 22641 5092 22651
rect 5040 22607 5046 22641
rect 5046 22607 5080 22641
rect 5080 22607 5092 22641
rect 5040 22599 5092 22607
rect 5106 22641 5158 22651
rect 5106 22607 5118 22641
rect 5118 22607 5152 22641
rect 5152 22607 5158 22641
rect 5106 22599 5158 22607
rect 5040 22568 5092 22582
rect 5040 22534 5046 22568
rect 5046 22534 5080 22568
rect 5080 22534 5092 22568
rect 5040 22530 5092 22534
rect 5106 22568 5158 22582
rect 5106 22534 5118 22568
rect 5118 22534 5152 22568
rect 5152 22534 5158 22568
rect 5106 22530 5158 22534
rect 5040 22495 5092 22513
rect 5040 22461 5046 22495
rect 5046 22461 5080 22495
rect 5080 22461 5092 22495
rect 5106 22495 5158 22513
rect 5106 22461 5118 22495
rect 5118 22461 5152 22495
rect 5152 22461 5158 22495
rect 5040 22422 5092 22444
rect 5106 22422 5158 22444
rect 5040 22392 5046 22422
rect 5046 22392 5092 22422
rect 5106 22392 5152 22422
rect 5152 22392 5158 22422
rect 5040 22323 5046 22375
rect 5046 22323 5092 22375
rect 5106 22323 5152 22375
rect 5152 22323 5158 22375
rect 5040 22254 5046 22306
rect 5046 22254 5092 22306
rect 5106 22254 5152 22306
rect 5152 22254 5158 22306
rect 5040 22184 5046 22236
rect 5046 22184 5092 22236
rect 5106 22184 5152 22236
rect 5152 22184 5158 22236
rect 5040 22114 5046 22166
rect 5046 22114 5092 22166
rect 5106 22114 5152 22166
rect 5152 22114 5158 22166
rect 5317 21930 5323 21982
rect 5323 21930 5369 21982
rect 5383 21930 5429 21982
rect 5429 21930 5435 21982
rect 5317 21861 5323 21913
rect 5323 21861 5369 21913
rect 5383 21861 5429 21913
rect 5429 21861 5435 21913
rect 5317 21792 5323 21844
rect 5323 21792 5369 21844
rect 5383 21792 5429 21844
rect 5429 21792 5435 21844
rect 5317 21723 5323 21775
rect 5323 21723 5369 21775
rect 5383 21723 5429 21775
rect 5429 21723 5435 21775
rect 5317 21654 5323 21706
rect 5323 21654 5369 21706
rect 5383 21654 5429 21706
rect 5429 21654 5435 21706
rect 5317 21584 5323 21636
rect 5323 21584 5369 21636
rect 5383 21584 5429 21636
rect 5429 21584 5435 21636
rect 5317 21514 5323 21566
rect 5323 21514 5369 21566
rect 5383 21514 5429 21566
rect 5429 21514 5435 21566
rect 5317 21444 5323 21496
rect 5323 21444 5369 21496
rect 5383 21444 5429 21496
rect 5429 21444 5435 21496
rect 5317 21380 5323 21426
rect 5323 21380 5369 21426
rect 5383 21380 5429 21426
rect 5429 21380 5435 21426
rect 5317 21374 5369 21380
rect 5383 21374 5435 21380
rect 5594 22714 5646 22720
rect 5594 22680 5600 22714
rect 5600 22680 5634 22714
rect 5634 22680 5646 22714
rect 5594 22668 5646 22680
rect 5660 22714 5712 22720
rect 5660 22680 5672 22714
rect 5672 22680 5706 22714
rect 5706 22680 5712 22714
rect 5660 22668 5712 22680
rect 5594 22641 5646 22651
rect 5594 22607 5600 22641
rect 5600 22607 5634 22641
rect 5634 22607 5646 22641
rect 5594 22599 5646 22607
rect 5660 22641 5712 22651
rect 5660 22607 5672 22641
rect 5672 22607 5706 22641
rect 5706 22607 5712 22641
rect 5660 22599 5712 22607
rect 5594 22568 5646 22582
rect 5594 22534 5600 22568
rect 5600 22534 5634 22568
rect 5634 22534 5646 22568
rect 5594 22530 5646 22534
rect 5660 22568 5712 22582
rect 5660 22534 5672 22568
rect 5672 22534 5706 22568
rect 5706 22534 5712 22568
rect 5660 22530 5712 22534
rect 5594 22495 5646 22513
rect 5594 22461 5600 22495
rect 5600 22461 5634 22495
rect 5634 22461 5646 22495
rect 5660 22495 5712 22513
rect 5660 22461 5672 22495
rect 5672 22461 5706 22495
rect 5706 22461 5712 22495
rect 5594 22422 5646 22444
rect 5660 22422 5712 22444
rect 5594 22392 5600 22422
rect 5600 22392 5646 22422
rect 5660 22392 5706 22422
rect 5706 22392 5712 22422
rect 5594 22323 5600 22375
rect 5600 22323 5646 22375
rect 5660 22323 5706 22375
rect 5706 22323 5712 22375
rect 5594 22254 5600 22306
rect 5600 22254 5646 22306
rect 5660 22254 5706 22306
rect 5706 22254 5712 22306
rect 5594 22184 5600 22236
rect 5600 22184 5646 22236
rect 5660 22184 5706 22236
rect 5706 22184 5712 22236
rect 5594 22114 5600 22166
rect 5600 22114 5646 22166
rect 5660 22114 5706 22166
rect 5706 22114 5712 22166
rect 5871 21930 5877 21982
rect 5877 21930 5923 21982
rect 5937 21930 5983 21982
rect 5983 21930 5989 21982
rect 5871 21861 5877 21913
rect 5877 21861 5923 21913
rect 5937 21861 5983 21913
rect 5983 21861 5989 21913
rect 5871 21792 5877 21844
rect 5877 21792 5923 21844
rect 5937 21792 5983 21844
rect 5983 21792 5989 21844
rect 5871 21723 5877 21775
rect 5877 21723 5923 21775
rect 5937 21723 5983 21775
rect 5983 21723 5989 21775
rect 5871 21654 5877 21706
rect 5877 21654 5923 21706
rect 5937 21654 5983 21706
rect 5983 21654 5989 21706
rect 5871 21584 5877 21636
rect 5877 21584 5923 21636
rect 5937 21584 5983 21636
rect 5983 21584 5989 21636
rect 5871 21514 5877 21566
rect 5877 21514 5923 21566
rect 5937 21514 5983 21566
rect 5983 21514 5989 21566
rect 5871 21444 5877 21496
rect 5877 21444 5923 21496
rect 5937 21444 5983 21496
rect 5983 21444 5989 21496
rect 5871 21380 5877 21426
rect 5877 21380 5923 21426
rect 5937 21380 5983 21426
rect 5983 21380 5989 21426
rect 5871 21374 5923 21380
rect 5937 21374 5989 21380
rect 6148 22714 6200 22720
rect 6148 22680 6154 22714
rect 6154 22680 6188 22714
rect 6188 22680 6200 22714
rect 6148 22668 6200 22680
rect 6214 22714 6266 22720
rect 6214 22680 6226 22714
rect 6226 22680 6260 22714
rect 6260 22680 6266 22714
rect 6214 22668 6266 22680
rect 6148 22641 6200 22651
rect 6148 22607 6154 22641
rect 6154 22607 6188 22641
rect 6188 22607 6200 22641
rect 6148 22599 6200 22607
rect 6214 22641 6266 22651
rect 6214 22607 6226 22641
rect 6226 22607 6260 22641
rect 6260 22607 6266 22641
rect 6214 22599 6266 22607
rect 6148 22568 6200 22582
rect 6148 22534 6154 22568
rect 6154 22534 6188 22568
rect 6188 22534 6200 22568
rect 6148 22530 6200 22534
rect 6214 22568 6266 22582
rect 6214 22534 6226 22568
rect 6226 22534 6260 22568
rect 6260 22534 6266 22568
rect 6214 22530 6266 22534
rect 6148 22495 6200 22513
rect 6148 22461 6154 22495
rect 6154 22461 6188 22495
rect 6188 22461 6200 22495
rect 6214 22495 6266 22513
rect 6214 22461 6226 22495
rect 6226 22461 6260 22495
rect 6260 22461 6266 22495
rect 6148 22422 6200 22444
rect 6214 22422 6266 22444
rect 6148 22392 6154 22422
rect 6154 22392 6200 22422
rect 6214 22392 6260 22422
rect 6260 22392 6266 22422
rect 6148 22323 6154 22375
rect 6154 22323 6200 22375
rect 6214 22323 6260 22375
rect 6260 22323 6266 22375
rect 6148 22254 6154 22306
rect 6154 22254 6200 22306
rect 6214 22254 6260 22306
rect 6260 22254 6266 22306
rect 6148 22184 6154 22236
rect 6154 22184 6200 22236
rect 6214 22184 6260 22236
rect 6260 22184 6266 22236
rect 6148 22114 6154 22166
rect 6154 22114 6200 22166
rect 6214 22114 6260 22166
rect 6260 22114 6266 22166
rect 6425 21930 6431 21982
rect 6431 21930 6477 21982
rect 6491 21930 6537 21982
rect 6537 21930 6543 21982
rect 6425 21861 6431 21913
rect 6431 21861 6477 21913
rect 6491 21861 6537 21913
rect 6537 21861 6543 21913
rect 6425 21792 6431 21844
rect 6431 21792 6477 21844
rect 6491 21792 6537 21844
rect 6537 21792 6543 21844
rect 6425 21723 6431 21775
rect 6431 21723 6477 21775
rect 6491 21723 6537 21775
rect 6537 21723 6543 21775
rect 6425 21654 6431 21706
rect 6431 21654 6477 21706
rect 6491 21654 6537 21706
rect 6537 21654 6543 21706
rect 6425 21584 6431 21636
rect 6431 21584 6477 21636
rect 6491 21584 6537 21636
rect 6537 21584 6543 21636
rect 6425 21514 6431 21566
rect 6431 21514 6477 21566
rect 6491 21514 6537 21566
rect 6537 21514 6543 21566
rect 6425 21444 6431 21496
rect 6431 21444 6477 21496
rect 6491 21444 6537 21496
rect 6537 21444 6543 21496
rect 6425 21380 6431 21426
rect 6431 21380 6477 21426
rect 6491 21380 6537 21426
rect 6537 21380 6543 21426
rect 6425 21374 6477 21380
rect 6491 21374 6543 21380
rect 6702 22714 6754 22720
rect 6702 22680 6708 22714
rect 6708 22680 6742 22714
rect 6742 22680 6754 22714
rect 6702 22668 6754 22680
rect 6768 22714 6820 22720
rect 6768 22680 6780 22714
rect 6780 22680 6814 22714
rect 6814 22680 6820 22714
rect 6768 22668 6820 22680
rect 6702 22641 6754 22651
rect 6702 22607 6708 22641
rect 6708 22607 6742 22641
rect 6742 22607 6754 22641
rect 6702 22599 6754 22607
rect 6768 22641 6820 22651
rect 6768 22607 6780 22641
rect 6780 22607 6814 22641
rect 6814 22607 6820 22641
rect 6768 22599 6820 22607
rect 6702 22568 6754 22582
rect 6702 22534 6708 22568
rect 6708 22534 6742 22568
rect 6742 22534 6754 22568
rect 6702 22530 6754 22534
rect 6768 22568 6820 22582
rect 6768 22534 6780 22568
rect 6780 22534 6814 22568
rect 6814 22534 6820 22568
rect 6768 22530 6820 22534
rect 6702 22495 6754 22513
rect 6702 22461 6708 22495
rect 6708 22461 6742 22495
rect 6742 22461 6754 22495
rect 6768 22495 6820 22513
rect 6768 22461 6780 22495
rect 6780 22461 6814 22495
rect 6814 22461 6820 22495
rect 6702 22422 6754 22444
rect 6768 22422 6820 22444
rect 6702 22392 6708 22422
rect 6708 22392 6754 22422
rect 6768 22392 6814 22422
rect 6814 22392 6820 22422
rect 6702 22323 6708 22375
rect 6708 22323 6754 22375
rect 6768 22323 6814 22375
rect 6814 22323 6820 22375
rect 6702 22254 6708 22306
rect 6708 22254 6754 22306
rect 6768 22254 6814 22306
rect 6814 22254 6820 22306
rect 6702 22184 6708 22236
rect 6708 22184 6754 22236
rect 6768 22184 6814 22236
rect 6814 22184 6820 22236
rect 6702 22114 6708 22166
rect 6708 22114 6754 22166
rect 6768 22114 6814 22166
rect 6814 22114 6820 22166
rect 6979 21930 6985 21982
rect 6985 21930 7031 21982
rect 7045 21930 7091 21982
rect 7091 21930 7097 21982
rect 6979 21861 6985 21913
rect 6985 21861 7031 21913
rect 7045 21861 7091 21913
rect 7091 21861 7097 21913
rect 6979 21792 6985 21844
rect 6985 21792 7031 21844
rect 7045 21792 7091 21844
rect 7091 21792 7097 21844
rect 6979 21723 6985 21775
rect 6985 21723 7031 21775
rect 7045 21723 7091 21775
rect 7091 21723 7097 21775
rect 6979 21654 6985 21706
rect 6985 21654 7031 21706
rect 7045 21654 7091 21706
rect 7091 21654 7097 21706
rect 6979 21584 6985 21636
rect 6985 21584 7031 21636
rect 7045 21584 7091 21636
rect 7091 21584 7097 21636
rect 6979 21514 6985 21566
rect 6985 21514 7031 21566
rect 7045 21514 7091 21566
rect 7091 21514 7097 21566
rect 6979 21444 6985 21496
rect 6985 21444 7031 21496
rect 7045 21444 7091 21496
rect 7091 21444 7097 21496
rect 6979 21380 6985 21426
rect 6985 21380 7031 21426
rect 7045 21380 7091 21426
rect 7091 21380 7097 21426
rect 6979 21374 7031 21380
rect 7045 21374 7097 21380
rect 7256 22714 7308 22720
rect 7256 22680 7262 22714
rect 7262 22680 7296 22714
rect 7296 22680 7308 22714
rect 7256 22668 7308 22680
rect 7322 22714 7374 22720
rect 7322 22680 7334 22714
rect 7334 22680 7368 22714
rect 7368 22680 7374 22714
rect 7322 22668 7374 22680
rect 7256 22641 7308 22651
rect 7256 22607 7262 22641
rect 7262 22607 7296 22641
rect 7296 22607 7308 22641
rect 7256 22599 7308 22607
rect 7322 22641 7374 22651
rect 7322 22607 7334 22641
rect 7334 22607 7368 22641
rect 7368 22607 7374 22641
rect 7322 22599 7374 22607
rect 7256 22568 7308 22582
rect 7256 22534 7262 22568
rect 7262 22534 7296 22568
rect 7296 22534 7308 22568
rect 7256 22530 7308 22534
rect 7322 22568 7374 22582
rect 7322 22534 7334 22568
rect 7334 22534 7368 22568
rect 7368 22534 7374 22568
rect 7322 22530 7374 22534
rect 7256 22495 7308 22513
rect 7256 22461 7262 22495
rect 7262 22461 7296 22495
rect 7296 22461 7308 22495
rect 7322 22495 7374 22513
rect 7322 22461 7334 22495
rect 7334 22461 7368 22495
rect 7368 22461 7374 22495
rect 7256 22422 7308 22444
rect 7322 22422 7374 22444
rect 7256 22392 7262 22422
rect 7262 22392 7308 22422
rect 7322 22392 7368 22422
rect 7368 22392 7374 22422
rect 7256 22323 7262 22375
rect 7262 22323 7308 22375
rect 7322 22323 7368 22375
rect 7368 22323 7374 22375
rect 7256 22254 7262 22306
rect 7262 22254 7308 22306
rect 7322 22254 7368 22306
rect 7368 22254 7374 22306
rect 7256 22184 7262 22236
rect 7262 22184 7308 22236
rect 7322 22184 7368 22236
rect 7368 22184 7374 22236
rect 7256 22114 7262 22166
rect 7262 22114 7308 22166
rect 7322 22114 7368 22166
rect 7368 22114 7374 22166
rect 7533 21930 7539 21982
rect 7539 21930 7585 21982
rect 7599 21930 7645 21982
rect 7645 21930 7651 21982
rect 7533 21861 7539 21913
rect 7539 21861 7585 21913
rect 7599 21861 7645 21913
rect 7645 21861 7651 21913
rect 7533 21792 7539 21844
rect 7539 21792 7585 21844
rect 7599 21792 7645 21844
rect 7645 21792 7651 21844
rect 7533 21723 7539 21775
rect 7539 21723 7585 21775
rect 7599 21723 7645 21775
rect 7645 21723 7651 21775
rect 7533 21654 7539 21706
rect 7539 21654 7585 21706
rect 7599 21654 7645 21706
rect 7645 21654 7651 21706
rect 7533 21584 7539 21636
rect 7539 21584 7585 21636
rect 7599 21584 7645 21636
rect 7645 21584 7651 21636
rect 7533 21514 7539 21566
rect 7539 21514 7585 21566
rect 7599 21514 7645 21566
rect 7645 21514 7651 21566
rect 7533 21444 7539 21496
rect 7539 21444 7585 21496
rect 7599 21444 7645 21496
rect 7645 21444 7651 21496
rect 7533 21380 7539 21426
rect 7539 21380 7585 21426
rect 7599 21380 7645 21426
rect 7645 21380 7651 21426
rect 7533 21374 7585 21380
rect 7599 21374 7651 21380
rect 7810 22714 7862 22720
rect 7810 22680 7816 22714
rect 7816 22680 7850 22714
rect 7850 22680 7862 22714
rect 7810 22668 7862 22680
rect 7876 22714 7928 22720
rect 7876 22680 7888 22714
rect 7888 22680 7922 22714
rect 7922 22680 7928 22714
rect 7876 22668 7928 22680
rect 7810 22641 7862 22651
rect 7810 22607 7816 22641
rect 7816 22607 7850 22641
rect 7850 22607 7862 22641
rect 7810 22599 7862 22607
rect 7876 22641 7928 22651
rect 7876 22607 7888 22641
rect 7888 22607 7922 22641
rect 7922 22607 7928 22641
rect 7876 22599 7928 22607
rect 7810 22568 7862 22582
rect 7810 22534 7816 22568
rect 7816 22534 7850 22568
rect 7850 22534 7862 22568
rect 7810 22530 7862 22534
rect 7876 22568 7928 22582
rect 7876 22534 7888 22568
rect 7888 22534 7922 22568
rect 7922 22534 7928 22568
rect 7876 22530 7928 22534
rect 7810 22495 7862 22513
rect 7810 22461 7816 22495
rect 7816 22461 7850 22495
rect 7850 22461 7862 22495
rect 7876 22495 7928 22513
rect 7876 22461 7888 22495
rect 7888 22461 7922 22495
rect 7922 22461 7928 22495
rect 7810 22422 7862 22444
rect 7876 22422 7928 22444
rect 7810 22392 7816 22422
rect 7816 22392 7862 22422
rect 7876 22392 7922 22422
rect 7922 22392 7928 22422
rect 7810 22323 7816 22375
rect 7816 22323 7862 22375
rect 7876 22323 7922 22375
rect 7922 22323 7928 22375
rect 7810 22254 7816 22306
rect 7816 22254 7862 22306
rect 7876 22254 7922 22306
rect 7922 22254 7928 22306
rect 7810 22184 7816 22236
rect 7816 22184 7862 22236
rect 7876 22184 7922 22236
rect 7922 22184 7928 22236
rect 7810 22114 7816 22166
rect 7816 22114 7862 22166
rect 7876 22114 7922 22166
rect 7922 22114 7928 22166
rect 8047 22701 8050 22724
rect 8050 22701 8084 22724
rect 8084 22701 8099 22724
rect 8047 22672 8099 22701
rect 8169 22691 8184 22724
rect 8184 22691 8218 22724
rect 8218 22691 8221 22724
rect 8169 22672 8221 22691
rect 8047 22629 8050 22655
rect 8050 22629 8084 22655
rect 8084 22629 8099 22655
rect 8047 22603 8099 22629
rect 8169 22653 8221 22655
rect 8169 22619 8184 22653
rect 8184 22619 8218 22653
rect 8218 22619 8221 22653
rect 8169 22603 8221 22619
rect 8047 22557 8050 22586
rect 8050 22557 8084 22586
rect 8084 22557 8099 22586
rect 8047 22534 8099 22557
rect 8169 22581 8221 22586
rect 8169 22547 8184 22581
rect 8184 22547 8218 22581
rect 8218 22547 8221 22581
rect 8169 22534 8221 22547
rect 8047 22485 8050 22517
rect 8050 22485 8084 22517
rect 8084 22485 8099 22517
rect 8047 22465 8099 22485
rect 8169 22509 8221 22517
rect 8169 22475 8184 22509
rect 8184 22475 8218 22509
rect 8218 22475 8221 22509
rect 8169 22465 8221 22475
rect 8047 22447 8099 22448
rect 8047 22413 8050 22447
rect 8050 22413 8084 22447
rect 8084 22413 8099 22447
rect 8047 22396 8099 22413
rect 8169 22437 8221 22448
rect 8169 22403 8184 22437
rect 8184 22403 8218 22437
rect 8218 22403 8221 22437
rect 8169 22396 8221 22403
rect 8047 22375 8099 22378
rect 8047 22341 8050 22375
rect 8050 22341 8084 22375
rect 8084 22341 8099 22375
rect 8047 22326 8099 22341
rect 8169 22365 8221 22378
rect 8169 22331 8184 22365
rect 8184 22331 8218 22365
rect 8218 22331 8221 22365
rect 8169 22326 8221 22331
rect 8047 22303 8099 22308
rect 8047 22269 8050 22303
rect 8050 22269 8084 22303
rect 8084 22269 8099 22303
rect 8047 22256 8099 22269
rect 8169 22293 8221 22308
rect 8169 22259 8184 22293
rect 8184 22259 8218 22293
rect 8218 22259 8221 22293
rect 8169 22256 8221 22259
rect 8047 22231 8099 22238
rect 8047 22197 8050 22231
rect 8050 22197 8084 22231
rect 8084 22197 8099 22231
rect 8047 22186 8099 22197
rect 8169 22221 8221 22238
rect 8169 22187 8184 22221
rect 8184 22187 8218 22221
rect 8218 22187 8221 22221
rect 8169 22186 8221 22187
rect 8047 22159 8099 22168
rect 8047 22125 8050 22159
rect 8050 22125 8084 22159
rect 8084 22125 8099 22159
rect 8047 22116 8099 22125
rect 8169 22149 8221 22168
rect 8169 22116 8184 22149
rect 8184 22116 8218 22149
rect 8218 22116 8221 22149
rect 5040 20714 5092 20720
rect 5040 20680 5046 20714
rect 5046 20680 5080 20714
rect 5080 20680 5092 20714
rect 5040 20668 5092 20680
rect 5106 20714 5158 20720
rect 5106 20680 5118 20714
rect 5118 20680 5152 20714
rect 5152 20680 5158 20714
rect 5106 20668 5158 20680
rect 5040 20641 5092 20651
rect 5040 20607 5046 20641
rect 5046 20607 5080 20641
rect 5080 20607 5092 20641
rect 5040 20599 5092 20607
rect 5106 20641 5158 20651
rect 5106 20607 5118 20641
rect 5118 20607 5152 20641
rect 5152 20607 5158 20641
rect 5106 20599 5158 20607
rect 5040 20568 5092 20582
rect 5040 20534 5046 20568
rect 5046 20534 5080 20568
rect 5080 20534 5092 20568
rect 5040 20530 5092 20534
rect 5106 20568 5158 20582
rect 5106 20534 5118 20568
rect 5118 20534 5152 20568
rect 5152 20534 5158 20568
rect 5106 20530 5158 20534
rect 5040 20495 5092 20513
rect 5040 20461 5046 20495
rect 5046 20461 5080 20495
rect 5080 20461 5092 20495
rect 5106 20495 5158 20513
rect 5106 20461 5118 20495
rect 5118 20461 5152 20495
rect 5152 20461 5158 20495
rect 5040 20422 5092 20444
rect 5106 20422 5158 20444
rect 5040 20392 5046 20422
rect 5046 20392 5092 20422
rect 5106 20392 5152 20422
rect 5152 20392 5158 20422
rect 5040 20323 5046 20375
rect 5046 20323 5092 20375
rect 5106 20323 5152 20375
rect 5152 20323 5158 20375
rect 5040 20254 5046 20306
rect 5046 20254 5092 20306
rect 5106 20254 5152 20306
rect 5152 20254 5158 20306
rect 5040 20184 5046 20236
rect 5046 20184 5092 20236
rect 5106 20184 5152 20236
rect 5152 20184 5158 20236
rect 5040 20114 5046 20166
rect 5046 20114 5092 20166
rect 5106 20114 5152 20166
rect 5152 20114 5158 20166
rect 5317 19930 5323 19982
rect 5323 19930 5369 19982
rect 5383 19930 5429 19982
rect 5429 19930 5435 19982
rect 5317 19861 5323 19913
rect 5323 19861 5369 19913
rect 5383 19861 5429 19913
rect 5429 19861 5435 19913
rect 5317 19792 5323 19844
rect 5323 19792 5369 19844
rect 5383 19792 5429 19844
rect 5429 19792 5435 19844
rect 5317 19723 5323 19775
rect 5323 19723 5369 19775
rect 5383 19723 5429 19775
rect 5429 19723 5435 19775
rect 5317 19654 5323 19706
rect 5323 19654 5369 19706
rect 5383 19654 5429 19706
rect 5429 19654 5435 19706
rect 5317 19584 5323 19636
rect 5323 19584 5369 19636
rect 5383 19584 5429 19636
rect 5429 19584 5435 19636
rect 5317 19514 5323 19566
rect 5323 19514 5369 19566
rect 5383 19514 5429 19566
rect 5429 19514 5435 19566
rect 5317 19444 5323 19496
rect 5323 19444 5369 19496
rect 5383 19444 5429 19496
rect 5429 19444 5435 19496
rect 5317 19380 5323 19426
rect 5323 19380 5369 19426
rect 5383 19380 5429 19426
rect 5429 19380 5435 19426
rect 5317 19374 5369 19380
rect 5383 19374 5435 19380
rect 5594 20714 5646 20720
rect 5594 20680 5600 20714
rect 5600 20680 5634 20714
rect 5634 20680 5646 20714
rect 5594 20668 5646 20680
rect 5660 20714 5712 20720
rect 5660 20680 5672 20714
rect 5672 20680 5706 20714
rect 5706 20680 5712 20714
rect 5660 20668 5712 20680
rect 5594 20641 5646 20651
rect 5594 20607 5600 20641
rect 5600 20607 5634 20641
rect 5634 20607 5646 20641
rect 5594 20599 5646 20607
rect 5660 20641 5712 20651
rect 5660 20607 5672 20641
rect 5672 20607 5706 20641
rect 5706 20607 5712 20641
rect 5660 20599 5712 20607
rect 5594 20568 5646 20582
rect 5594 20534 5600 20568
rect 5600 20534 5634 20568
rect 5634 20534 5646 20568
rect 5594 20530 5646 20534
rect 5660 20568 5712 20582
rect 5660 20534 5672 20568
rect 5672 20534 5706 20568
rect 5706 20534 5712 20568
rect 5660 20530 5712 20534
rect 5594 20495 5646 20513
rect 5594 20461 5600 20495
rect 5600 20461 5634 20495
rect 5634 20461 5646 20495
rect 5660 20495 5712 20513
rect 5660 20461 5672 20495
rect 5672 20461 5706 20495
rect 5706 20461 5712 20495
rect 5594 20422 5646 20444
rect 5660 20422 5712 20444
rect 5594 20392 5600 20422
rect 5600 20392 5646 20422
rect 5660 20392 5706 20422
rect 5706 20392 5712 20422
rect 5594 20323 5600 20375
rect 5600 20323 5646 20375
rect 5660 20323 5706 20375
rect 5706 20323 5712 20375
rect 5594 20254 5600 20306
rect 5600 20254 5646 20306
rect 5660 20254 5706 20306
rect 5706 20254 5712 20306
rect 5594 20184 5600 20236
rect 5600 20184 5646 20236
rect 5660 20184 5706 20236
rect 5706 20184 5712 20236
rect 5594 20114 5600 20166
rect 5600 20114 5646 20166
rect 5660 20114 5706 20166
rect 5706 20114 5712 20166
rect 5871 19930 5877 19982
rect 5877 19930 5923 19982
rect 5937 19930 5983 19982
rect 5983 19930 5989 19982
rect 5871 19861 5877 19913
rect 5877 19861 5923 19913
rect 5937 19861 5983 19913
rect 5983 19861 5989 19913
rect 5871 19792 5877 19844
rect 5877 19792 5923 19844
rect 5937 19792 5983 19844
rect 5983 19792 5989 19844
rect 5871 19723 5877 19775
rect 5877 19723 5923 19775
rect 5937 19723 5983 19775
rect 5983 19723 5989 19775
rect 5871 19654 5877 19706
rect 5877 19654 5923 19706
rect 5937 19654 5983 19706
rect 5983 19654 5989 19706
rect 5871 19584 5877 19636
rect 5877 19584 5923 19636
rect 5937 19584 5983 19636
rect 5983 19584 5989 19636
rect 5871 19514 5877 19566
rect 5877 19514 5923 19566
rect 5937 19514 5983 19566
rect 5983 19514 5989 19566
rect 5871 19444 5877 19496
rect 5877 19444 5923 19496
rect 5937 19444 5983 19496
rect 5983 19444 5989 19496
rect 5871 19380 5877 19426
rect 5877 19380 5923 19426
rect 5937 19380 5983 19426
rect 5983 19380 5989 19426
rect 5871 19374 5923 19380
rect 5937 19374 5989 19380
rect 6148 20714 6200 20720
rect 6148 20680 6154 20714
rect 6154 20680 6188 20714
rect 6188 20680 6200 20714
rect 6148 20668 6200 20680
rect 6214 20714 6266 20720
rect 6214 20680 6226 20714
rect 6226 20680 6260 20714
rect 6260 20680 6266 20714
rect 6214 20668 6266 20680
rect 6148 20641 6200 20651
rect 6148 20607 6154 20641
rect 6154 20607 6188 20641
rect 6188 20607 6200 20641
rect 6148 20599 6200 20607
rect 6214 20641 6266 20651
rect 6214 20607 6226 20641
rect 6226 20607 6260 20641
rect 6260 20607 6266 20641
rect 6214 20599 6266 20607
rect 6148 20568 6200 20582
rect 6148 20534 6154 20568
rect 6154 20534 6188 20568
rect 6188 20534 6200 20568
rect 6148 20530 6200 20534
rect 6214 20568 6266 20582
rect 6214 20534 6226 20568
rect 6226 20534 6260 20568
rect 6260 20534 6266 20568
rect 6214 20530 6266 20534
rect 6148 20495 6200 20513
rect 6148 20461 6154 20495
rect 6154 20461 6188 20495
rect 6188 20461 6200 20495
rect 6214 20495 6266 20513
rect 6214 20461 6226 20495
rect 6226 20461 6260 20495
rect 6260 20461 6266 20495
rect 6148 20422 6200 20444
rect 6214 20422 6266 20444
rect 6148 20392 6154 20422
rect 6154 20392 6200 20422
rect 6214 20392 6260 20422
rect 6260 20392 6266 20422
rect 6148 20323 6154 20375
rect 6154 20323 6200 20375
rect 6214 20323 6260 20375
rect 6260 20323 6266 20375
rect 6148 20254 6154 20306
rect 6154 20254 6200 20306
rect 6214 20254 6260 20306
rect 6260 20254 6266 20306
rect 6148 20184 6154 20236
rect 6154 20184 6200 20236
rect 6214 20184 6260 20236
rect 6260 20184 6266 20236
rect 6148 20114 6154 20166
rect 6154 20114 6200 20166
rect 6214 20114 6260 20166
rect 6260 20114 6266 20166
rect 6425 19930 6431 19982
rect 6431 19930 6477 19982
rect 6491 19930 6537 19982
rect 6537 19930 6543 19982
rect 6425 19861 6431 19913
rect 6431 19861 6477 19913
rect 6491 19861 6537 19913
rect 6537 19861 6543 19913
rect 6425 19792 6431 19844
rect 6431 19792 6477 19844
rect 6491 19792 6537 19844
rect 6537 19792 6543 19844
rect 6425 19723 6431 19775
rect 6431 19723 6477 19775
rect 6491 19723 6537 19775
rect 6537 19723 6543 19775
rect 6425 19654 6431 19706
rect 6431 19654 6477 19706
rect 6491 19654 6537 19706
rect 6537 19654 6543 19706
rect 6425 19584 6431 19636
rect 6431 19584 6477 19636
rect 6491 19584 6537 19636
rect 6537 19584 6543 19636
rect 6425 19514 6431 19566
rect 6431 19514 6477 19566
rect 6491 19514 6537 19566
rect 6537 19514 6543 19566
rect 6425 19444 6431 19496
rect 6431 19444 6477 19496
rect 6491 19444 6537 19496
rect 6537 19444 6543 19496
rect 6425 19380 6431 19426
rect 6431 19380 6477 19426
rect 6491 19380 6537 19426
rect 6537 19380 6543 19426
rect 6425 19374 6477 19380
rect 6491 19374 6543 19380
rect 6702 20714 6754 20720
rect 6702 20680 6708 20714
rect 6708 20680 6742 20714
rect 6742 20680 6754 20714
rect 6702 20668 6754 20680
rect 6768 20714 6820 20720
rect 6768 20680 6780 20714
rect 6780 20680 6814 20714
rect 6814 20680 6820 20714
rect 6768 20668 6820 20680
rect 6702 20641 6754 20651
rect 6702 20607 6708 20641
rect 6708 20607 6742 20641
rect 6742 20607 6754 20641
rect 6702 20599 6754 20607
rect 6768 20641 6820 20651
rect 6768 20607 6780 20641
rect 6780 20607 6814 20641
rect 6814 20607 6820 20641
rect 6768 20599 6820 20607
rect 6702 20568 6754 20582
rect 6702 20534 6708 20568
rect 6708 20534 6742 20568
rect 6742 20534 6754 20568
rect 6702 20530 6754 20534
rect 6768 20568 6820 20582
rect 6768 20534 6780 20568
rect 6780 20534 6814 20568
rect 6814 20534 6820 20568
rect 6768 20530 6820 20534
rect 6702 20495 6754 20513
rect 6702 20461 6708 20495
rect 6708 20461 6742 20495
rect 6742 20461 6754 20495
rect 6768 20495 6820 20513
rect 6768 20461 6780 20495
rect 6780 20461 6814 20495
rect 6814 20461 6820 20495
rect 6702 20422 6754 20444
rect 6768 20422 6820 20444
rect 6702 20392 6708 20422
rect 6708 20392 6754 20422
rect 6768 20392 6814 20422
rect 6814 20392 6820 20422
rect 6702 20323 6708 20375
rect 6708 20323 6754 20375
rect 6768 20323 6814 20375
rect 6814 20323 6820 20375
rect 6702 20254 6708 20306
rect 6708 20254 6754 20306
rect 6768 20254 6814 20306
rect 6814 20254 6820 20306
rect 6702 20184 6708 20236
rect 6708 20184 6754 20236
rect 6768 20184 6814 20236
rect 6814 20184 6820 20236
rect 6702 20114 6708 20166
rect 6708 20114 6754 20166
rect 6768 20114 6814 20166
rect 6814 20114 6820 20166
rect 6979 19930 6985 19982
rect 6985 19930 7031 19982
rect 7045 19930 7091 19982
rect 7091 19930 7097 19982
rect 6979 19861 6985 19913
rect 6985 19861 7031 19913
rect 7045 19861 7091 19913
rect 7091 19861 7097 19913
rect 6979 19792 6985 19844
rect 6985 19792 7031 19844
rect 7045 19792 7091 19844
rect 7091 19792 7097 19844
rect 6979 19723 6985 19775
rect 6985 19723 7031 19775
rect 7045 19723 7091 19775
rect 7091 19723 7097 19775
rect 6979 19654 6985 19706
rect 6985 19654 7031 19706
rect 7045 19654 7091 19706
rect 7091 19654 7097 19706
rect 6979 19584 6985 19636
rect 6985 19584 7031 19636
rect 7045 19584 7091 19636
rect 7091 19584 7097 19636
rect 6979 19514 6985 19566
rect 6985 19514 7031 19566
rect 7045 19514 7091 19566
rect 7091 19514 7097 19566
rect 6979 19444 6985 19496
rect 6985 19444 7031 19496
rect 7045 19444 7091 19496
rect 7091 19444 7097 19496
rect 6979 19380 6985 19426
rect 6985 19380 7031 19426
rect 7045 19380 7091 19426
rect 7091 19380 7097 19426
rect 6979 19374 7031 19380
rect 7045 19374 7097 19380
rect 7256 20714 7308 20720
rect 7256 20680 7262 20714
rect 7262 20680 7296 20714
rect 7296 20680 7308 20714
rect 7256 20668 7308 20680
rect 7322 20714 7374 20720
rect 7322 20680 7334 20714
rect 7334 20680 7368 20714
rect 7368 20680 7374 20714
rect 7322 20668 7374 20680
rect 7256 20641 7308 20651
rect 7256 20607 7262 20641
rect 7262 20607 7296 20641
rect 7296 20607 7308 20641
rect 7256 20599 7308 20607
rect 7322 20641 7374 20651
rect 7322 20607 7334 20641
rect 7334 20607 7368 20641
rect 7368 20607 7374 20641
rect 7322 20599 7374 20607
rect 7256 20568 7308 20582
rect 7256 20534 7262 20568
rect 7262 20534 7296 20568
rect 7296 20534 7308 20568
rect 7256 20530 7308 20534
rect 7322 20568 7374 20582
rect 7322 20534 7334 20568
rect 7334 20534 7368 20568
rect 7368 20534 7374 20568
rect 7322 20530 7374 20534
rect 7256 20495 7308 20513
rect 7256 20461 7262 20495
rect 7262 20461 7296 20495
rect 7296 20461 7308 20495
rect 7322 20495 7374 20513
rect 7322 20461 7334 20495
rect 7334 20461 7368 20495
rect 7368 20461 7374 20495
rect 7256 20422 7308 20444
rect 7322 20422 7374 20444
rect 7256 20392 7262 20422
rect 7262 20392 7308 20422
rect 7322 20392 7368 20422
rect 7368 20392 7374 20422
rect 7256 20323 7262 20375
rect 7262 20323 7308 20375
rect 7322 20323 7368 20375
rect 7368 20323 7374 20375
rect 7256 20254 7262 20306
rect 7262 20254 7308 20306
rect 7322 20254 7368 20306
rect 7368 20254 7374 20306
rect 7256 20184 7262 20236
rect 7262 20184 7308 20236
rect 7322 20184 7368 20236
rect 7368 20184 7374 20236
rect 7256 20114 7262 20166
rect 7262 20114 7308 20166
rect 7322 20114 7368 20166
rect 7368 20114 7374 20166
rect 7533 19930 7539 19982
rect 7539 19930 7585 19982
rect 7599 19930 7645 19982
rect 7645 19930 7651 19982
rect 7533 19861 7539 19913
rect 7539 19861 7585 19913
rect 7599 19861 7645 19913
rect 7645 19861 7651 19913
rect 7533 19792 7539 19844
rect 7539 19792 7585 19844
rect 7599 19792 7645 19844
rect 7645 19792 7651 19844
rect 7533 19723 7539 19775
rect 7539 19723 7585 19775
rect 7599 19723 7645 19775
rect 7645 19723 7651 19775
rect 7533 19654 7539 19706
rect 7539 19654 7585 19706
rect 7599 19654 7645 19706
rect 7645 19654 7651 19706
rect 7533 19584 7539 19636
rect 7539 19584 7585 19636
rect 7599 19584 7645 19636
rect 7645 19584 7651 19636
rect 7533 19514 7539 19566
rect 7539 19514 7585 19566
rect 7599 19514 7645 19566
rect 7645 19514 7651 19566
rect 7533 19444 7539 19496
rect 7539 19444 7585 19496
rect 7599 19444 7645 19496
rect 7645 19444 7651 19496
rect 7533 19380 7539 19426
rect 7539 19380 7585 19426
rect 7599 19380 7645 19426
rect 7645 19380 7651 19426
rect 7533 19374 7585 19380
rect 7599 19374 7651 19380
rect 7810 20714 7862 20720
rect 7810 20680 7816 20714
rect 7816 20680 7850 20714
rect 7850 20680 7862 20714
rect 7810 20668 7862 20680
rect 7876 20714 7928 20720
rect 7876 20680 7888 20714
rect 7888 20680 7922 20714
rect 7922 20680 7928 20714
rect 7876 20668 7928 20680
rect 7810 20641 7862 20651
rect 7810 20607 7816 20641
rect 7816 20607 7850 20641
rect 7850 20607 7862 20641
rect 7810 20599 7862 20607
rect 7876 20641 7928 20651
rect 7876 20607 7888 20641
rect 7888 20607 7922 20641
rect 7922 20607 7928 20641
rect 7876 20599 7928 20607
rect 7810 20568 7862 20582
rect 7810 20534 7816 20568
rect 7816 20534 7850 20568
rect 7850 20534 7862 20568
rect 7810 20530 7862 20534
rect 7876 20568 7928 20582
rect 7876 20534 7888 20568
rect 7888 20534 7922 20568
rect 7922 20534 7928 20568
rect 7876 20530 7928 20534
rect 7810 20495 7862 20513
rect 7810 20461 7816 20495
rect 7816 20461 7850 20495
rect 7850 20461 7862 20495
rect 7876 20495 7928 20513
rect 7876 20461 7888 20495
rect 7888 20461 7922 20495
rect 7922 20461 7928 20495
rect 7810 20422 7862 20444
rect 7876 20422 7928 20444
rect 7810 20392 7816 20422
rect 7816 20392 7862 20422
rect 7876 20392 7922 20422
rect 7922 20392 7928 20422
rect 7810 20323 7816 20375
rect 7816 20323 7862 20375
rect 7876 20323 7922 20375
rect 7922 20323 7928 20375
rect 7810 20254 7816 20306
rect 7816 20254 7862 20306
rect 7876 20254 7922 20306
rect 7922 20254 7928 20306
rect 7810 20184 7816 20236
rect 7816 20184 7862 20236
rect 7876 20184 7922 20236
rect 7922 20184 7928 20236
rect 7810 20114 7816 20166
rect 7816 20114 7862 20166
rect 7876 20114 7922 20166
rect 7922 20114 7928 20166
rect 8047 20719 8099 20724
rect 8047 20685 8050 20719
rect 8050 20685 8084 20719
rect 8084 20685 8099 20719
rect 8047 20672 8099 20685
rect 8169 20709 8221 20724
rect 8169 20675 8184 20709
rect 8184 20675 8218 20709
rect 8218 20675 8221 20709
rect 8169 20672 8221 20675
rect 8047 20647 8099 20655
rect 8047 20613 8050 20647
rect 8050 20613 8084 20647
rect 8084 20613 8099 20647
rect 8047 20603 8099 20613
rect 8169 20637 8221 20655
rect 8169 20603 8184 20637
rect 8184 20603 8218 20637
rect 8218 20603 8221 20637
rect 8047 20575 8099 20586
rect 8047 20541 8050 20575
rect 8050 20541 8084 20575
rect 8084 20541 8099 20575
rect 8047 20534 8099 20541
rect 8169 20565 8221 20586
rect 8169 20534 8184 20565
rect 8184 20534 8218 20565
rect 8218 20534 8221 20565
rect 8047 20503 8099 20517
rect 8047 20469 8050 20503
rect 8050 20469 8084 20503
rect 8084 20469 8099 20503
rect 8047 20465 8099 20469
rect 8169 20493 8221 20517
rect 8169 20465 8184 20493
rect 8184 20465 8218 20493
rect 8218 20465 8221 20493
rect 8047 20431 8099 20448
rect 8047 20397 8050 20431
rect 8050 20397 8084 20431
rect 8084 20397 8099 20431
rect 8047 20396 8099 20397
rect 8169 20421 8221 20448
rect 8169 20396 8184 20421
rect 8184 20396 8218 20421
rect 8218 20396 8221 20421
rect 8047 20359 8099 20378
rect 8047 20326 8050 20359
rect 8050 20326 8084 20359
rect 8084 20326 8099 20359
rect 8169 20349 8221 20378
rect 8169 20326 8184 20349
rect 8184 20326 8218 20349
rect 8218 20326 8221 20349
rect 8047 20287 8099 20308
rect 8047 20256 8050 20287
rect 8050 20256 8084 20287
rect 8084 20256 8099 20287
rect 8169 20277 8221 20308
rect 8169 20256 8184 20277
rect 8184 20256 8218 20277
rect 8218 20256 8221 20277
rect 8047 20215 8099 20238
rect 8047 20186 8050 20215
rect 8050 20186 8084 20215
rect 8084 20186 8099 20215
rect 8169 20205 8221 20238
rect 8169 20186 8184 20205
rect 8184 20186 8218 20205
rect 8218 20186 8221 20205
rect 8047 20143 8099 20168
rect 8047 20116 8050 20143
rect 8050 20116 8084 20143
rect 8084 20116 8099 20143
rect 8169 20133 8221 20168
rect 8169 20116 8184 20133
rect 8184 20116 8218 20133
rect 8218 20116 8221 20133
rect 5040 18714 5092 18720
rect 5040 18680 5046 18714
rect 5046 18680 5080 18714
rect 5080 18680 5092 18714
rect 5040 18668 5092 18680
rect 5106 18714 5158 18720
rect 5106 18680 5118 18714
rect 5118 18680 5152 18714
rect 5152 18680 5158 18714
rect 5106 18668 5158 18680
rect 5040 18641 5092 18651
rect 5040 18607 5046 18641
rect 5046 18607 5080 18641
rect 5080 18607 5092 18641
rect 5040 18599 5092 18607
rect 5106 18641 5158 18651
rect 5106 18607 5118 18641
rect 5118 18607 5152 18641
rect 5152 18607 5158 18641
rect 5106 18599 5158 18607
rect 5040 18568 5092 18582
rect 5040 18534 5046 18568
rect 5046 18534 5080 18568
rect 5080 18534 5092 18568
rect 5040 18530 5092 18534
rect 5106 18568 5158 18582
rect 5106 18534 5118 18568
rect 5118 18534 5152 18568
rect 5152 18534 5158 18568
rect 5106 18530 5158 18534
rect 5040 18495 5092 18513
rect 5040 18461 5046 18495
rect 5046 18461 5080 18495
rect 5080 18461 5092 18495
rect 5106 18495 5158 18513
rect 5106 18461 5118 18495
rect 5118 18461 5152 18495
rect 5152 18461 5158 18495
rect 5040 18422 5092 18444
rect 5106 18422 5158 18444
rect 5040 18392 5046 18422
rect 5046 18392 5092 18422
rect 5106 18392 5152 18422
rect 5152 18392 5158 18422
rect 5040 18323 5046 18375
rect 5046 18323 5092 18375
rect 5106 18323 5152 18375
rect 5152 18323 5158 18375
rect 5040 18254 5046 18306
rect 5046 18254 5092 18306
rect 5106 18254 5152 18306
rect 5152 18254 5158 18306
rect 5040 18184 5046 18236
rect 5046 18184 5092 18236
rect 5106 18184 5152 18236
rect 5152 18184 5158 18236
rect 5040 18114 5046 18166
rect 5046 18114 5092 18166
rect 5106 18114 5152 18166
rect 5152 18114 5158 18166
rect 5317 17930 5323 17982
rect 5323 17930 5369 17982
rect 5383 17930 5429 17982
rect 5429 17930 5435 17982
rect 5317 17861 5323 17913
rect 5323 17861 5369 17913
rect 5383 17861 5429 17913
rect 5429 17861 5435 17913
rect 5317 17792 5323 17844
rect 5323 17792 5369 17844
rect 5383 17792 5429 17844
rect 5429 17792 5435 17844
rect 5317 17723 5323 17775
rect 5323 17723 5369 17775
rect 5383 17723 5429 17775
rect 5429 17723 5435 17775
rect 5317 17654 5323 17706
rect 5323 17654 5369 17706
rect 5383 17654 5429 17706
rect 5429 17654 5435 17706
rect 5317 17584 5323 17636
rect 5323 17584 5369 17636
rect 5383 17584 5429 17636
rect 5429 17584 5435 17636
rect 5317 17514 5323 17566
rect 5323 17514 5369 17566
rect 5383 17514 5429 17566
rect 5429 17514 5435 17566
rect 5317 17444 5323 17496
rect 5323 17444 5369 17496
rect 5383 17444 5429 17496
rect 5429 17444 5435 17496
rect 5317 17380 5323 17426
rect 5323 17380 5369 17426
rect 5383 17380 5429 17426
rect 5429 17380 5435 17426
rect 5317 17374 5369 17380
rect 5383 17374 5435 17380
rect 5594 18714 5646 18720
rect 5594 18680 5600 18714
rect 5600 18680 5634 18714
rect 5634 18680 5646 18714
rect 5594 18668 5646 18680
rect 5660 18714 5712 18720
rect 5660 18680 5672 18714
rect 5672 18680 5706 18714
rect 5706 18680 5712 18714
rect 5660 18668 5712 18680
rect 5594 18641 5646 18651
rect 5594 18607 5600 18641
rect 5600 18607 5634 18641
rect 5634 18607 5646 18641
rect 5594 18599 5646 18607
rect 5660 18641 5712 18651
rect 5660 18607 5672 18641
rect 5672 18607 5706 18641
rect 5706 18607 5712 18641
rect 5660 18599 5712 18607
rect 5594 18568 5646 18582
rect 5594 18534 5600 18568
rect 5600 18534 5634 18568
rect 5634 18534 5646 18568
rect 5594 18530 5646 18534
rect 5660 18568 5712 18582
rect 5660 18534 5672 18568
rect 5672 18534 5706 18568
rect 5706 18534 5712 18568
rect 5660 18530 5712 18534
rect 5594 18495 5646 18513
rect 5594 18461 5600 18495
rect 5600 18461 5634 18495
rect 5634 18461 5646 18495
rect 5660 18495 5712 18513
rect 5660 18461 5672 18495
rect 5672 18461 5706 18495
rect 5706 18461 5712 18495
rect 5594 18422 5646 18444
rect 5660 18422 5712 18444
rect 5594 18392 5600 18422
rect 5600 18392 5646 18422
rect 5660 18392 5706 18422
rect 5706 18392 5712 18422
rect 5594 18323 5600 18375
rect 5600 18323 5646 18375
rect 5660 18323 5706 18375
rect 5706 18323 5712 18375
rect 5594 18254 5600 18306
rect 5600 18254 5646 18306
rect 5660 18254 5706 18306
rect 5706 18254 5712 18306
rect 5594 18184 5600 18236
rect 5600 18184 5646 18236
rect 5660 18184 5706 18236
rect 5706 18184 5712 18236
rect 5594 18114 5600 18166
rect 5600 18114 5646 18166
rect 5660 18114 5706 18166
rect 5706 18114 5712 18166
rect 5871 17930 5877 17982
rect 5877 17930 5923 17982
rect 5937 17930 5983 17982
rect 5983 17930 5989 17982
rect 5871 17861 5877 17913
rect 5877 17861 5923 17913
rect 5937 17861 5983 17913
rect 5983 17861 5989 17913
rect 5871 17792 5877 17844
rect 5877 17792 5923 17844
rect 5937 17792 5983 17844
rect 5983 17792 5989 17844
rect 5871 17723 5877 17775
rect 5877 17723 5923 17775
rect 5937 17723 5983 17775
rect 5983 17723 5989 17775
rect 5871 17654 5877 17706
rect 5877 17654 5923 17706
rect 5937 17654 5983 17706
rect 5983 17654 5989 17706
rect 5871 17584 5877 17636
rect 5877 17584 5923 17636
rect 5937 17584 5983 17636
rect 5983 17584 5989 17636
rect 5871 17514 5877 17566
rect 5877 17514 5923 17566
rect 5937 17514 5983 17566
rect 5983 17514 5989 17566
rect 5871 17444 5877 17496
rect 5877 17444 5923 17496
rect 5937 17444 5983 17496
rect 5983 17444 5989 17496
rect 5871 17380 5877 17426
rect 5877 17380 5923 17426
rect 5937 17380 5983 17426
rect 5983 17380 5989 17426
rect 5871 17374 5923 17380
rect 5937 17374 5989 17380
rect 6148 18714 6200 18720
rect 6148 18680 6154 18714
rect 6154 18680 6188 18714
rect 6188 18680 6200 18714
rect 6148 18668 6200 18680
rect 6214 18714 6266 18720
rect 6214 18680 6226 18714
rect 6226 18680 6260 18714
rect 6260 18680 6266 18714
rect 6214 18668 6266 18680
rect 6148 18641 6200 18651
rect 6148 18607 6154 18641
rect 6154 18607 6188 18641
rect 6188 18607 6200 18641
rect 6148 18599 6200 18607
rect 6214 18641 6266 18651
rect 6214 18607 6226 18641
rect 6226 18607 6260 18641
rect 6260 18607 6266 18641
rect 6214 18599 6266 18607
rect 6148 18568 6200 18582
rect 6148 18534 6154 18568
rect 6154 18534 6188 18568
rect 6188 18534 6200 18568
rect 6148 18530 6200 18534
rect 6214 18568 6266 18582
rect 6214 18534 6226 18568
rect 6226 18534 6260 18568
rect 6260 18534 6266 18568
rect 6214 18530 6266 18534
rect 6148 18495 6200 18513
rect 6148 18461 6154 18495
rect 6154 18461 6188 18495
rect 6188 18461 6200 18495
rect 6214 18495 6266 18513
rect 6214 18461 6226 18495
rect 6226 18461 6260 18495
rect 6260 18461 6266 18495
rect 6148 18422 6200 18444
rect 6214 18422 6266 18444
rect 6148 18392 6154 18422
rect 6154 18392 6200 18422
rect 6214 18392 6260 18422
rect 6260 18392 6266 18422
rect 6148 18323 6154 18375
rect 6154 18323 6200 18375
rect 6214 18323 6260 18375
rect 6260 18323 6266 18375
rect 6148 18254 6154 18306
rect 6154 18254 6200 18306
rect 6214 18254 6260 18306
rect 6260 18254 6266 18306
rect 6148 18184 6154 18236
rect 6154 18184 6200 18236
rect 6214 18184 6260 18236
rect 6260 18184 6266 18236
rect 6148 18114 6154 18166
rect 6154 18114 6200 18166
rect 6214 18114 6260 18166
rect 6260 18114 6266 18166
rect 6425 17930 6431 17982
rect 6431 17930 6477 17982
rect 6491 17930 6537 17982
rect 6537 17930 6543 17982
rect 6425 17861 6431 17913
rect 6431 17861 6477 17913
rect 6491 17861 6537 17913
rect 6537 17861 6543 17913
rect 6425 17792 6431 17844
rect 6431 17792 6477 17844
rect 6491 17792 6537 17844
rect 6537 17792 6543 17844
rect 6425 17723 6431 17775
rect 6431 17723 6477 17775
rect 6491 17723 6537 17775
rect 6537 17723 6543 17775
rect 6425 17654 6431 17706
rect 6431 17654 6477 17706
rect 6491 17654 6537 17706
rect 6537 17654 6543 17706
rect 6425 17584 6431 17636
rect 6431 17584 6477 17636
rect 6491 17584 6537 17636
rect 6537 17584 6543 17636
rect 6425 17514 6431 17566
rect 6431 17514 6477 17566
rect 6491 17514 6537 17566
rect 6537 17514 6543 17566
rect 6425 17444 6431 17496
rect 6431 17444 6477 17496
rect 6491 17444 6537 17496
rect 6537 17444 6543 17496
rect 6425 17380 6431 17426
rect 6431 17380 6477 17426
rect 6491 17380 6537 17426
rect 6537 17380 6543 17426
rect 6425 17374 6477 17380
rect 6491 17374 6543 17380
rect 6702 18714 6754 18720
rect 6702 18680 6708 18714
rect 6708 18680 6742 18714
rect 6742 18680 6754 18714
rect 6702 18668 6754 18680
rect 6768 18714 6820 18720
rect 6768 18680 6780 18714
rect 6780 18680 6814 18714
rect 6814 18680 6820 18714
rect 6768 18668 6820 18680
rect 6702 18641 6754 18651
rect 6702 18607 6708 18641
rect 6708 18607 6742 18641
rect 6742 18607 6754 18641
rect 6702 18599 6754 18607
rect 6768 18641 6820 18651
rect 6768 18607 6780 18641
rect 6780 18607 6814 18641
rect 6814 18607 6820 18641
rect 6768 18599 6820 18607
rect 6702 18568 6754 18582
rect 6702 18534 6708 18568
rect 6708 18534 6742 18568
rect 6742 18534 6754 18568
rect 6702 18530 6754 18534
rect 6768 18568 6820 18582
rect 6768 18534 6780 18568
rect 6780 18534 6814 18568
rect 6814 18534 6820 18568
rect 6768 18530 6820 18534
rect 6702 18495 6754 18513
rect 6702 18461 6708 18495
rect 6708 18461 6742 18495
rect 6742 18461 6754 18495
rect 6768 18495 6820 18513
rect 6768 18461 6780 18495
rect 6780 18461 6814 18495
rect 6814 18461 6820 18495
rect 6702 18422 6754 18444
rect 6768 18422 6820 18444
rect 6702 18392 6708 18422
rect 6708 18392 6754 18422
rect 6768 18392 6814 18422
rect 6814 18392 6820 18422
rect 6702 18323 6708 18375
rect 6708 18323 6754 18375
rect 6768 18323 6814 18375
rect 6814 18323 6820 18375
rect 6702 18254 6708 18306
rect 6708 18254 6754 18306
rect 6768 18254 6814 18306
rect 6814 18254 6820 18306
rect 6702 18184 6708 18236
rect 6708 18184 6754 18236
rect 6768 18184 6814 18236
rect 6814 18184 6820 18236
rect 6702 18114 6708 18166
rect 6708 18114 6754 18166
rect 6768 18114 6814 18166
rect 6814 18114 6820 18166
rect 6979 17930 6985 17982
rect 6985 17930 7031 17982
rect 7045 17930 7091 17982
rect 7091 17930 7097 17982
rect 6979 17861 6985 17913
rect 6985 17861 7031 17913
rect 7045 17861 7091 17913
rect 7091 17861 7097 17913
rect 6979 17792 6985 17844
rect 6985 17792 7031 17844
rect 7045 17792 7091 17844
rect 7091 17792 7097 17844
rect 6979 17723 6985 17775
rect 6985 17723 7031 17775
rect 7045 17723 7091 17775
rect 7091 17723 7097 17775
rect 6979 17654 6985 17706
rect 6985 17654 7031 17706
rect 7045 17654 7091 17706
rect 7091 17654 7097 17706
rect 6979 17584 6985 17636
rect 6985 17584 7031 17636
rect 7045 17584 7091 17636
rect 7091 17584 7097 17636
rect 6979 17514 6985 17566
rect 6985 17514 7031 17566
rect 7045 17514 7091 17566
rect 7091 17514 7097 17566
rect 6979 17444 6985 17496
rect 6985 17444 7031 17496
rect 7045 17444 7091 17496
rect 7091 17444 7097 17496
rect 6979 17380 6985 17426
rect 6985 17380 7031 17426
rect 7045 17380 7091 17426
rect 7091 17380 7097 17426
rect 6979 17374 7031 17380
rect 7045 17374 7097 17380
rect 7256 18714 7308 18720
rect 7256 18680 7262 18714
rect 7262 18680 7296 18714
rect 7296 18680 7308 18714
rect 7256 18668 7308 18680
rect 7322 18714 7374 18720
rect 7322 18680 7334 18714
rect 7334 18680 7368 18714
rect 7368 18680 7374 18714
rect 7322 18668 7374 18680
rect 7256 18641 7308 18651
rect 7256 18607 7262 18641
rect 7262 18607 7296 18641
rect 7296 18607 7308 18641
rect 7256 18599 7308 18607
rect 7322 18641 7374 18651
rect 7322 18607 7334 18641
rect 7334 18607 7368 18641
rect 7368 18607 7374 18641
rect 7322 18599 7374 18607
rect 7256 18568 7308 18582
rect 7256 18534 7262 18568
rect 7262 18534 7296 18568
rect 7296 18534 7308 18568
rect 7256 18530 7308 18534
rect 7322 18568 7374 18582
rect 7322 18534 7334 18568
rect 7334 18534 7368 18568
rect 7368 18534 7374 18568
rect 7322 18530 7374 18534
rect 7256 18495 7308 18513
rect 7256 18461 7262 18495
rect 7262 18461 7296 18495
rect 7296 18461 7308 18495
rect 7322 18495 7374 18513
rect 7322 18461 7334 18495
rect 7334 18461 7368 18495
rect 7368 18461 7374 18495
rect 7256 18422 7308 18444
rect 7322 18422 7374 18444
rect 7256 18392 7262 18422
rect 7262 18392 7308 18422
rect 7322 18392 7368 18422
rect 7368 18392 7374 18422
rect 7256 18323 7262 18375
rect 7262 18323 7308 18375
rect 7322 18323 7368 18375
rect 7368 18323 7374 18375
rect 7256 18254 7262 18306
rect 7262 18254 7308 18306
rect 7322 18254 7368 18306
rect 7368 18254 7374 18306
rect 7256 18184 7262 18236
rect 7262 18184 7308 18236
rect 7322 18184 7368 18236
rect 7368 18184 7374 18236
rect 7256 18114 7262 18166
rect 7262 18114 7308 18166
rect 7322 18114 7368 18166
rect 7368 18114 7374 18166
rect 7533 17930 7539 17982
rect 7539 17930 7585 17982
rect 7599 17930 7645 17982
rect 7645 17930 7651 17982
rect 7533 17861 7539 17913
rect 7539 17861 7585 17913
rect 7599 17861 7645 17913
rect 7645 17861 7651 17913
rect 7533 17792 7539 17844
rect 7539 17792 7585 17844
rect 7599 17792 7645 17844
rect 7645 17792 7651 17844
rect 7533 17723 7539 17775
rect 7539 17723 7585 17775
rect 7599 17723 7645 17775
rect 7645 17723 7651 17775
rect 7533 17654 7539 17706
rect 7539 17654 7585 17706
rect 7599 17654 7645 17706
rect 7645 17654 7651 17706
rect 7533 17584 7539 17636
rect 7539 17584 7585 17636
rect 7599 17584 7645 17636
rect 7645 17584 7651 17636
rect 7533 17514 7539 17566
rect 7539 17514 7585 17566
rect 7599 17514 7645 17566
rect 7645 17514 7651 17566
rect 7533 17444 7539 17496
rect 7539 17444 7585 17496
rect 7599 17444 7645 17496
rect 7645 17444 7651 17496
rect 7533 17380 7539 17426
rect 7539 17380 7585 17426
rect 7599 17380 7645 17426
rect 7645 17380 7651 17426
rect 7533 17374 7585 17380
rect 7599 17374 7651 17380
rect 7810 18714 7862 18720
rect 7810 18680 7816 18714
rect 7816 18680 7850 18714
rect 7850 18680 7862 18714
rect 7810 18668 7862 18680
rect 7876 18714 7928 18720
rect 7876 18680 7888 18714
rect 7888 18680 7922 18714
rect 7922 18680 7928 18714
rect 7876 18668 7928 18680
rect 7810 18641 7862 18651
rect 7810 18607 7816 18641
rect 7816 18607 7850 18641
rect 7850 18607 7862 18641
rect 7810 18599 7862 18607
rect 7876 18641 7928 18651
rect 7876 18607 7888 18641
rect 7888 18607 7922 18641
rect 7922 18607 7928 18641
rect 7876 18599 7928 18607
rect 7810 18568 7862 18582
rect 7810 18534 7816 18568
rect 7816 18534 7850 18568
rect 7850 18534 7862 18568
rect 7810 18530 7862 18534
rect 7876 18568 7928 18582
rect 7876 18534 7888 18568
rect 7888 18534 7922 18568
rect 7922 18534 7928 18568
rect 7876 18530 7928 18534
rect 7810 18495 7862 18513
rect 7810 18461 7816 18495
rect 7816 18461 7850 18495
rect 7850 18461 7862 18495
rect 7876 18495 7928 18513
rect 7876 18461 7888 18495
rect 7888 18461 7922 18495
rect 7922 18461 7928 18495
rect 7810 18422 7862 18444
rect 7876 18422 7928 18444
rect 7810 18392 7816 18422
rect 7816 18392 7862 18422
rect 7876 18392 7922 18422
rect 7922 18392 7928 18422
rect 7810 18323 7816 18375
rect 7816 18323 7862 18375
rect 7876 18323 7922 18375
rect 7922 18323 7928 18375
rect 7810 18254 7816 18306
rect 7816 18254 7862 18306
rect 7876 18254 7922 18306
rect 7922 18254 7928 18306
rect 7810 18184 7816 18236
rect 7816 18184 7862 18236
rect 7876 18184 7922 18236
rect 7922 18184 7928 18236
rect 7810 18114 7816 18166
rect 7816 18114 7862 18166
rect 7876 18114 7922 18166
rect 7922 18114 7928 18166
rect 8047 18703 8099 18724
rect 8047 18672 8050 18703
rect 8050 18672 8084 18703
rect 8084 18672 8099 18703
rect 8169 18693 8221 18724
rect 8169 18672 8184 18693
rect 8184 18672 8218 18693
rect 8218 18672 8221 18693
rect 8047 18631 8099 18655
rect 8047 18603 8050 18631
rect 8050 18603 8084 18631
rect 8084 18603 8099 18631
rect 8169 18621 8221 18655
rect 8169 18603 8184 18621
rect 8184 18603 8218 18621
rect 8218 18603 8221 18621
rect 8047 18559 8099 18586
rect 8047 18534 8050 18559
rect 8050 18534 8084 18559
rect 8084 18534 8099 18559
rect 8169 18549 8221 18586
rect 8169 18534 8184 18549
rect 8184 18534 8218 18549
rect 8218 18534 8221 18549
rect 8047 18487 8099 18517
rect 8047 18465 8050 18487
rect 8050 18465 8084 18487
rect 8084 18465 8099 18487
rect 8169 18515 8184 18517
rect 8184 18515 8218 18517
rect 8218 18515 8221 18517
rect 8169 18477 8221 18515
rect 8169 18465 8184 18477
rect 8184 18465 8218 18477
rect 8218 18465 8221 18477
rect 8047 18415 8099 18448
rect 8047 18396 8050 18415
rect 8050 18396 8084 18415
rect 8084 18396 8099 18415
rect 8169 18443 8184 18448
rect 8184 18443 8218 18448
rect 8218 18443 8221 18448
rect 8169 18405 8221 18443
rect 8169 18396 8184 18405
rect 8184 18396 8218 18405
rect 8218 18396 8221 18405
rect 8047 18343 8099 18378
rect 8047 18326 8050 18343
rect 8050 18326 8084 18343
rect 8084 18326 8099 18343
rect 8169 18371 8184 18378
rect 8184 18371 8218 18378
rect 8218 18371 8221 18378
rect 8169 18333 8221 18371
rect 8169 18326 8184 18333
rect 8184 18326 8218 18333
rect 8218 18326 8221 18333
rect 8047 18271 8099 18308
rect 8047 18256 8050 18271
rect 8050 18256 8084 18271
rect 8084 18256 8099 18271
rect 8169 18299 8184 18308
rect 8184 18299 8218 18308
rect 8218 18299 8221 18308
rect 8169 18261 8221 18299
rect 8169 18256 8184 18261
rect 8184 18256 8218 18261
rect 8218 18256 8221 18261
rect 8047 18237 8050 18238
rect 8050 18237 8084 18238
rect 8084 18237 8099 18238
rect 8047 18199 8099 18237
rect 8047 18186 8050 18199
rect 8050 18186 8084 18199
rect 8084 18186 8099 18199
rect 8169 18227 8184 18238
rect 8184 18227 8218 18238
rect 8218 18227 8221 18238
rect 8169 18189 8221 18227
rect 8169 18186 8184 18189
rect 8184 18186 8218 18189
rect 8218 18186 8221 18189
rect 8047 18165 8050 18168
rect 8050 18165 8084 18168
rect 8084 18165 8099 18168
rect 8047 18127 8099 18165
rect 8047 18116 8050 18127
rect 8050 18116 8084 18127
rect 8084 18116 8099 18127
rect 8169 18155 8184 18168
rect 8184 18155 8218 18168
rect 8218 18155 8221 18168
rect 8169 18117 8221 18155
rect 8169 18116 8184 18117
rect 8184 18116 8218 18117
rect 8218 18116 8221 18117
rect 5116 16955 5123 16970
rect 5123 16955 5162 16970
rect 5162 16955 5168 16970
rect 5182 16955 5196 16970
rect 5196 16955 5234 16970
rect 5248 16955 5269 16970
rect 5269 16955 5300 16970
rect 5314 16955 5342 16970
rect 5342 16955 5366 16970
rect 5116 16918 5168 16955
rect 5182 16918 5234 16955
rect 5248 16918 5300 16955
rect 5314 16918 5366 16955
rect 5380 16955 5381 16970
rect 5381 16955 5415 16970
rect 5415 16955 5432 16970
rect 5380 16918 5432 16955
rect 5446 16955 5454 16970
rect 5454 16955 5488 16970
rect 5488 16955 5498 16970
rect 5446 16918 5498 16955
rect 5512 16955 5527 16970
rect 5527 16955 5561 16970
rect 5561 16955 5564 16970
rect 5512 16918 5564 16955
rect 5578 16955 5600 16970
rect 5600 16955 5630 16970
rect 5644 16955 5673 16970
rect 5673 16955 5696 16970
rect 5710 16955 5746 16970
rect 5746 16955 5762 16970
rect 5776 16955 5780 16970
rect 5780 16955 5819 16970
rect 5819 16955 5828 16970
rect 5842 16955 5853 16970
rect 5853 16955 5892 16970
rect 5892 16955 5894 16970
rect 5908 16955 5926 16970
rect 5926 16955 5960 16970
rect 5974 16955 5999 16970
rect 5999 16955 6026 16970
rect 6040 16955 6072 16970
rect 6072 16955 6092 16970
rect 5578 16918 5630 16955
rect 5644 16918 5696 16955
rect 5710 16918 5762 16955
rect 5776 16918 5828 16955
rect 5842 16918 5894 16955
rect 5908 16918 5960 16955
rect 5974 16918 6026 16955
rect 6040 16918 6092 16955
rect 6106 16955 6110 16970
rect 6110 16955 6144 16970
rect 6144 16955 6158 16970
rect 6106 16918 6158 16955
rect 6172 16955 6182 16970
rect 6182 16955 6216 16970
rect 6216 16955 6224 16970
rect 6172 16918 6224 16955
rect 6238 16955 6254 16970
rect 6254 16955 6288 16970
rect 6288 16955 6290 16970
rect 6238 16918 6290 16955
rect 6304 16955 6326 16970
rect 6326 16955 6356 16970
rect 6370 16955 6398 16970
rect 6398 16955 6422 16970
rect 6436 16955 6470 16970
rect 6470 16955 6488 16970
rect 6501 16955 6504 16970
rect 6504 16955 6542 16970
rect 6542 16955 6553 16970
rect 6566 16955 6576 16970
rect 6576 16955 6614 16970
rect 6614 16955 6618 16970
rect 6631 16955 6648 16970
rect 6648 16955 6683 16970
rect 6696 16955 6720 16970
rect 6720 16955 6748 16970
rect 6761 16955 6792 16970
rect 6792 16955 6813 16970
rect 6304 16918 6356 16955
rect 6370 16918 6422 16955
rect 6436 16918 6488 16955
rect 6501 16918 6553 16955
rect 6566 16918 6618 16955
rect 6631 16918 6683 16955
rect 6696 16918 6748 16955
rect 6761 16918 6813 16955
rect 6826 16955 6830 16970
rect 6830 16955 6864 16970
rect 6864 16955 6878 16970
rect 6826 16918 6878 16955
rect 6891 16955 6902 16970
rect 6902 16955 6936 16970
rect 6936 16955 6943 16970
rect 6891 16918 6943 16955
rect 6956 16955 6974 16970
rect 6974 16955 7008 16970
rect 6956 16918 7008 16955
rect 7021 16955 7046 16970
rect 7046 16955 7073 16970
rect 7086 16955 7118 16970
rect 7118 16955 7138 16970
rect 7151 16955 7152 16970
rect 7152 16955 7190 16970
rect 7190 16955 7203 16970
rect 7216 16955 7224 16970
rect 7224 16955 7262 16970
rect 7262 16955 7268 16970
rect 7281 16955 7296 16970
rect 7296 16955 7333 16970
rect 7346 16955 7368 16970
rect 7368 16955 7398 16970
rect 7411 16955 7440 16970
rect 7440 16955 7463 16970
rect 7021 16918 7073 16955
rect 7086 16918 7138 16955
rect 7151 16918 7203 16955
rect 7216 16918 7268 16955
rect 7281 16918 7333 16955
rect 7346 16918 7398 16955
rect 7411 16918 7463 16955
rect 7476 16955 7478 16970
rect 7478 16955 7512 16970
rect 7512 16955 7528 16970
rect 7476 16918 7528 16955
rect 7541 16955 7550 16970
rect 7550 16955 7584 16970
rect 7584 16955 7593 16970
rect 7541 16918 7593 16955
rect 7606 16955 7622 16970
rect 7622 16955 7656 16970
rect 7656 16955 7658 16970
rect 7606 16918 7658 16955
rect 7671 16955 7694 16970
rect 7694 16955 7723 16970
rect 7736 16955 7766 16970
rect 7766 16955 7788 16970
rect 7801 16955 7838 16970
rect 7838 16955 7853 16970
rect 7671 16918 7723 16955
rect 7736 16918 7788 16955
rect 7801 16918 7853 16955
rect 5116 16879 5123 16904
rect 5123 16879 5162 16904
rect 5162 16879 5168 16904
rect 5182 16879 5196 16904
rect 5196 16879 5234 16904
rect 5248 16879 5269 16904
rect 5269 16879 5300 16904
rect 5314 16879 5342 16904
rect 5342 16879 5366 16904
rect 5116 16852 5168 16879
rect 5182 16852 5234 16879
rect 5248 16852 5300 16879
rect 5314 16852 5366 16879
rect 5380 16879 5381 16904
rect 5381 16879 5415 16904
rect 5415 16879 5432 16904
rect 5380 16852 5432 16879
rect 5446 16879 5454 16904
rect 5454 16879 5488 16904
rect 5488 16879 5498 16904
rect 5446 16852 5498 16879
rect 5512 16879 5527 16904
rect 5527 16879 5561 16904
rect 5561 16879 5564 16904
rect 5512 16852 5564 16879
rect 5578 16879 5600 16904
rect 5600 16879 5630 16904
rect 5644 16879 5673 16904
rect 5673 16879 5696 16904
rect 5710 16879 5746 16904
rect 5746 16879 5762 16904
rect 5776 16879 5780 16904
rect 5780 16879 5819 16904
rect 5819 16879 5828 16904
rect 5842 16879 5853 16904
rect 5853 16879 5892 16904
rect 5892 16879 5894 16904
rect 5908 16879 5926 16904
rect 5926 16879 5960 16904
rect 5974 16879 5999 16904
rect 5999 16879 6026 16904
rect 6040 16879 6072 16904
rect 6072 16879 6092 16904
rect 5578 16852 5630 16879
rect 5644 16852 5696 16879
rect 5710 16852 5762 16879
rect 5776 16852 5828 16879
rect 5842 16852 5894 16879
rect 5908 16852 5960 16879
rect 5974 16852 6026 16879
rect 6040 16852 6092 16879
rect 6106 16879 6110 16904
rect 6110 16879 6144 16904
rect 6144 16879 6158 16904
rect 6106 16852 6158 16879
rect 6172 16879 6182 16904
rect 6182 16879 6216 16904
rect 6216 16879 6224 16904
rect 6172 16852 6224 16879
rect 6238 16879 6254 16904
rect 6254 16879 6288 16904
rect 6288 16879 6290 16904
rect 6238 16852 6290 16879
rect 6304 16879 6326 16904
rect 6326 16879 6356 16904
rect 6370 16879 6398 16904
rect 6398 16879 6422 16904
rect 6436 16879 6470 16904
rect 6470 16879 6488 16904
rect 6501 16879 6504 16904
rect 6504 16879 6542 16904
rect 6542 16879 6553 16904
rect 6566 16879 6576 16904
rect 6576 16879 6614 16904
rect 6614 16879 6618 16904
rect 6631 16879 6648 16904
rect 6648 16879 6683 16904
rect 6696 16879 6720 16904
rect 6720 16879 6748 16904
rect 6761 16879 6792 16904
rect 6792 16879 6813 16904
rect 6304 16852 6356 16879
rect 6370 16852 6422 16879
rect 6436 16852 6488 16879
rect 6501 16852 6553 16879
rect 6566 16852 6618 16879
rect 6631 16852 6683 16879
rect 6696 16852 6748 16879
rect 6761 16852 6813 16879
rect 6826 16879 6830 16904
rect 6830 16879 6864 16904
rect 6864 16879 6878 16904
rect 6826 16852 6878 16879
rect 6891 16879 6902 16904
rect 6902 16879 6936 16904
rect 6936 16879 6943 16904
rect 6891 16852 6943 16879
rect 6956 16879 6974 16904
rect 6974 16879 7008 16904
rect 6956 16852 7008 16879
rect 7021 16879 7046 16904
rect 7046 16879 7073 16904
rect 7086 16879 7118 16904
rect 7118 16879 7138 16904
rect 7151 16879 7152 16904
rect 7152 16879 7190 16904
rect 7190 16879 7203 16904
rect 7216 16879 7224 16904
rect 7224 16879 7262 16904
rect 7262 16879 7268 16904
rect 7281 16879 7296 16904
rect 7296 16879 7333 16904
rect 7346 16879 7368 16904
rect 7368 16879 7398 16904
rect 7411 16879 7440 16904
rect 7440 16879 7463 16904
rect 7021 16852 7073 16879
rect 7086 16852 7138 16879
rect 7151 16852 7203 16879
rect 7216 16852 7268 16879
rect 7281 16852 7333 16879
rect 7346 16852 7398 16879
rect 7411 16852 7463 16879
rect 7476 16879 7478 16904
rect 7478 16879 7512 16904
rect 7512 16879 7528 16904
rect 7476 16852 7528 16879
rect 7541 16879 7550 16904
rect 7550 16879 7584 16904
rect 7584 16879 7593 16904
rect 7541 16852 7593 16879
rect 7606 16879 7622 16904
rect 7622 16879 7656 16904
rect 7656 16879 7658 16904
rect 7606 16852 7658 16879
rect 7671 16879 7694 16904
rect 7694 16879 7723 16904
rect 7736 16879 7766 16904
rect 7766 16879 7788 16904
rect 7801 16879 7838 16904
rect 7838 16879 7853 16904
rect 7671 16852 7723 16879
rect 7736 16852 7788 16879
rect 7801 16852 7853 16879
rect 5116 16837 5168 16838
rect 5182 16837 5234 16838
rect 5248 16837 5300 16838
rect 5314 16837 5366 16838
rect 5116 16803 5123 16837
rect 5123 16803 5162 16837
rect 5162 16803 5168 16837
rect 5182 16803 5196 16837
rect 5196 16803 5234 16837
rect 5248 16803 5269 16837
rect 5269 16803 5300 16837
rect 5314 16803 5342 16837
rect 5342 16803 5366 16837
rect 5116 16786 5168 16803
rect 5182 16786 5234 16803
rect 5248 16786 5300 16803
rect 5314 16786 5366 16803
rect 5380 16837 5432 16838
rect 5380 16803 5381 16837
rect 5381 16803 5415 16837
rect 5415 16803 5432 16837
rect 5380 16786 5432 16803
rect 5446 16837 5498 16838
rect 5446 16803 5454 16837
rect 5454 16803 5488 16837
rect 5488 16803 5498 16837
rect 5446 16786 5498 16803
rect 5512 16837 5564 16838
rect 5512 16803 5527 16837
rect 5527 16803 5561 16837
rect 5561 16803 5564 16837
rect 5512 16786 5564 16803
rect 5578 16837 5630 16838
rect 5644 16837 5696 16838
rect 5710 16837 5762 16838
rect 5776 16837 5828 16838
rect 5842 16837 5894 16838
rect 5908 16837 5960 16838
rect 5974 16837 6026 16838
rect 6040 16837 6092 16838
rect 5578 16803 5600 16837
rect 5600 16803 5630 16837
rect 5644 16803 5673 16837
rect 5673 16803 5696 16837
rect 5710 16803 5746 16837
rect 5746 16803 5762 16837
rect 5776 16803 5780 16837
rect 5780 16803 5819 16837
rect 5819 16803 5828 16837
rect 5842 16803 5853 16837
rect 5853 16803 5892 16837
rect 5892 16803 5894 16837
rect 5908 16803 5926 16837
rect 5926 16803 5960 16837
rect 5974 16803 5999 16837
rect 5999 16803 6026 16837
rect 6040 16803 6072 16837
rect 6072 16803 6092 16837
rect 5578 16786 5630 16803
rect 5644 16786 5696 16803
rect 5710 16786 5762 16803
rect 5776 16786 5828 16803
rect 5842 16786 5894 16803
rect 5908 16786 5960 16803
rect 5974 16786 6026 16803
rect 6040 16786 6092 16803
rect 6106 16837 6158 16838
rect 6106 16803 6110 16837
rect 6110 16803 6144 16837
rect 6144 16803 6158 16837
rect 6106 16786 6158 16803
rect 6172 16837 6224 16838
rect 6172 16803 6182 16837
rect 6182 16803 6216 16837
rect 6216 16803 6224 16837
rect 6172 16786 6224 16803
rect 6238 16837 6290 16838
rect 6238 16803 6254 16837
rect 6254 16803 6288 16837
rect 6288 16803 6290 16837
rect 6238 16786 6290 16803
rect 6304 16837 6356 16838
rect 6370 16837 6422 16838
rect 6436 16837 6488 16838
rect 6501 16837 6553 16838
rect 6566 16837 6618 16838
rect 6631 16837 6683 16838
rect 6696 16837 6748 16838
rect 6761 16837 6813 16838
rect 6304 16803 6326 16837
rect 6326 16803 6356 16837
rect 6370 16803 6398 16837
rect 6398 16803 6422 16837
rect 6436 16803 6470 16837
rect 6470 16803 6488 16837
rect 6501 16803 6504 16837
rect 6504 16803 6542 16837
rect 6542 16803 6553 16837
rect 6566 16803 6576 16837
rect 6576 16803 6614 16837
rect 6614 16803 6618 16837
rect 6631 16803 6648 16837
rect 6648 16803 6683 16837
rect 6696 16803 6720 16837
rect 6720 16803 6748 16837
rect 6761 16803 6792 16837
rect 6792 16803 6813 16837
rect 6304 16786 6356 16803
rect 6370 16786 6422 16803
rect 6436 16786 6488 16803
rect 6501 16786 6553 16803
rect 6566 16786 6618 16803
rect 6631 16786 6683 16803
rect 6696 16786 6748 16803
rect 6761 16786 6813 16803
rect 6826 16837 6878 16838
rect 6826 16803 6830 16837
rect 6830 16803 6864 16837
rect 6864 16803 6878 16837
rect 6826 16786 6878 16803
rect 6891 16837 6943 16838
rect 6891 16803 6902 16837
rect 6902 16803 6936 16837
rect 6936 16803 6943 16837
rect 6891 16786 6943 16803
rect 6956 16837 7008 16838
rect 6956 16803 6974 16837
rect 6974 16803 7008 16837
rect 6956 16786 7008 16803
rect 7021 16837 7073 16838
rect 7086 16837 7138 16838
rect 7151 16837 7203 16838
rect 7216 16837 7268 16838
rect 7281 16837 7333 16838
rect 7346 16837 7398 16838
rect 7411 16837 7463 16838
rect 7021 16803 7046 16837
rect 7046 16803 7073 16837
rect 7086 16803 7118 16837
rect 7118 16803 7138 16837
rect 7151 16803 7152 16837
rect 7152 16803 7190 16837
rect 7190 16803 7203 16837
rect 7216 16803 7224 16837
rect 7224 16803 7262 16837
rect 7262 16803 7268 16837
rect 7281 16803 7296 16837
rect 7296 16803 7333 16837
rect 7346 16803 7368 16837
rect 7368 16803 7398 16837
rect 7411 16803 7440 16837
rect 7440 16803 7463 16837
rect 7021 16786 7073 16803
rect 7086 16786 7138 16803
rect 7151 16786 7203 16803
rect 7216 16786 7268 16803
rect 7281 16786 7333 16803
rect 7346 16786 7398 16803
rect 7411 16786 7463 16803
rect 7476 16837 7528 16838
rect 7476 16803 7478 16837
rect 7478 16803 7512 16837
rect 7512 16803 7528 16837
rect 7476 16786 7528 16803
rect 7541 16837 7593 16838
rect 7541 16803 7550 16837
rect 7550 16803 7584 16837
rect 7584 16803 7593 16837
rect 7541 16786 7593 16803
rect 7606 16837 7658 16838
rect 7606 16803 7622 16837
rect 7622 16803 7656 16837
rect 7656 16803 7658 16837
rect 7606 16786 7658 16803
rect 7671 16837 7723 16838
rect 7736 16837 7788 16838
rect 7801 16837 7853 16838
rect 7671 16803 7694 16837
rect 7694 16803 7723 16837
rect 7736 16803 7766 16837
rect 7766 16803 7788 16837
rect 7801 16803 7838 16837
rect 7838 16803 7853 16837
rect 7671 16786 7723 16803
rect 7736 16786 7788 16803
rect 7801 16786 7853 16803
rect 5116 16761 5168 16772
rect 5182 16761 5234 16772
rect 5248 16761 5300 16772
rect 5314 16761 5366 16772
rect 5116 16727 5123 16761
rect 5123 16727 5162 16761
rect 5162 16727 5168 16761
rect 5182 16727 5196 16761
rect 5196 16727 5234 16761
rect 5248 16727 5269 16761
rect 5269 16727 5300 16761
rect 5314 16727 5342 16761
rect 5342 16727 5366 16761
rect 5116 16720 5168 16727
rect 5182 16720 5234 16727
rect 5248 16720 5300 16727
rect 5314 16720 5366 16727
rect 5380 16761 5432 16772
rect 5380 16727 5381 16761
rect 5381 16727 5415 16761
rect 5415 16727 5432 16761
rect 5380 16720 5432 16727
rect 5446 16761 5498 16772
rect 5446 16727 5454 16761
rect 5454 16727 5488 16761
rect 5488 16727 5498 16761
rect 5446 16720 5498 16727
rect 5512 16761 5564 16772
rect 5512 16727 5527 16761
rect 5527 16727 5561 16761
rect 5561 16727 5564 16761
rect 5512 16720 5564 16727
rect 5578 16761 5630 16772
rect 5644 16761 5696 16772
rect 5710 16761 5762 16772
rect 5776 16761 5828 16772
rect 5842 16761 5894 16772
rect 5908 16761 5960 16772
rect 5974 16761 6026 16772
rect 6040 16761 6092 16772
rect 5578 16727 5600 16761
rect 5600 16727 5630 16761
rect 5644 16727 5673 16761
rect 5673 16727 5696 16761
rect 5710 16727 5746 16761
rect 5746 16727 5762 16761
rect 5776 16727 5780 16761
rect 5780 16727 5819 16761
rect 5819 16727 5828 16761
rect 5842 16727 5853 16761
rect 5853 16727 5892 16761
rect 5892 16727 5894 16761
rect 5908 16727 5926 16761
rect 5926 16727 5960 16761
rect 5974 16727 5999 16761
rect 5999 16727 6026 16761
rect 6040 16727 6072 16761
rect 6072 16727 6092 16761
rect 5578 16720 5630 16727
rect 5644 16720 5696 16727
rect 5710 16720 5762 16727
rect 5776 16720 5828 16727
rect 5842 16720 5894 16727
rect 5908 16720 5960 16727
rect 5974 16720 6026 16727
rect 6040 16720 6092 16727
rect 6106 16761 6158 16772
rect 6106 16727 6110 16761
rect 6110 16727 6144 16761
rect 6144 16727 6158 16761
rect 6106 16720 6158 16727
rect 6172 16761 6224 16772
rect 6172 16727 6182 16761
rect 6182 16727 6216 16761
rect 6216 16727 6224 16761
rect 6172 16720 6224 16727
rect 6238 16761 6290 16772
rect 6238 16727 6254 16761
rect 6254 16727 6288 16761
rect 6288 16727 6290 16761
rect 6238 16720 6290 16727
rect 6304 16761 6356 16772
rect 6370 16761 6422 16772
rect 6436 16761 6488 16772
rect 6501 16761 6553 16772
rect 6566 16761 6618 16772
rect 6631 16761 6683 16772
rect 6696 16761 6748 16772
rect 6761 16761 6813 16772
rect 6304 16727 6326 16761
rect 6326 16727 6356 16761
rect 6370 16727 6398 16761
rect 6398 16727 6422 16761
rect 6436 16727 6470 16761
rect 6470 16727 6488 16761
rect 6501 16727 6504 16761
rect 6504 16727 6542 16761
rect 6542 16727 6553 16761
rect 6566 16727 6576 16761
rect 6576 16727 6614 16761
rect 6614 16727 6618 16761
rect 6631 16727 6648 16761
rect 6648 16727 6683 16761
rect 6696 16727 6720 16761
rect 6720 16727 6748 16761
rect 6761 16727 6792 16761
rect 6792 16727 6813 16761
rect 6304 16720 6356 16727
rect 6370 16720 6422 16727
rect 6436 16720 6488 16727
rect 6501 16720 6553 16727
rect 6566 16720 6618 16727
rect 6631 16720 6683 16727
rect 6696 16720 6748 16727
rect 6761 16720 6813 16727
rect 6826 16761 6878 16772
rect 6826 16727 6830 16761
rect 6830 16727 6864 16761
rect 6864 16727 6878 16761
rect 6826 16720 6878 16727
rect 6891 16761 6943 16772
rect 6891 16727 6902 16761
rect 6902 16727 6936 16761
rect 6936 16727 6943 16761
rect 6891 16720 6943 16727
rect 6956 16761 7008 16772
rect 6956 16727 6974 16761
rect 6974 16727 7008 16761
rect 6956 16720 7008 16727
rect 7021 16761 7073 16772
rect 7086 16761 7138 16772
rect 7151 16761 7203 16772
rect 7216 16761 7268 16772
rect 7281 16761 7333 16772
rect 7346 16761 7398 16772
rect 7411 16761 7463 16772
rect 7021 16727 7046 16761
rect 7046 16727 7073 16761
rect 7086 16727 7118 16761
rect 7118 16727 7138 16761
rect 7151 16727 7152 16761
rect 7152 16727 7190 16761
rect 7190 16727 7203 16761
rect 7216 16727 7224 16761
rect 7224 16727 7262 16761
rect 7262 16727 7268 16761
rect 7281 16727 7296 16761
rect 7296 16727 7333 16761
rect 7346 16727 7368 16761
rect 7368 16727 7398 16761
rect 7411 16727 7440 16761
rect 7440 16727 7463 16761
rect 7021 16720 7073 16727
rect 7086 16720 7138 16727
rect 7151 16720 7203 16727
rect 7216 16720 7268 16727
rect 7281 16720 7333 16727
rect 7346 16720 7398 16727
rect 7411 16720 7463 16727
rect 7476 16761 7528 16772
rect 7476 16727 7478 16761
rect 7478 16727 7512 16761
rect 7512 16727 7528 16761
rect 7476 16720 7528 16727
rect 7541 16761 7593 16772
rect 7541 16727 7550 16761
rect 7550 16727 7584 16761
rect 7584 16727 7593 16761
rect 7541 16720 7593 16727
rect 7606 16761 7658 16772
rect 7606 16727 7622 16761
rect 7622 16727 7656 16761
rect 7656 16727 7658 16761
rect 7606 16720 7658 16727
rect 7671 16761 7723 16772
rect 7736 16761 7788 16772
rect 7801 16761 7853 16772
rect 7671 16727 7694 16761
rect 7694 16727 7723 16761
rect 7736 16727 7766 16761
rect 7766 16727 7788 16761
rect 7801 16727 7838 16761
rect 7838 16727 7853 16761
rect 7671 16720 7723 16727
rect 7736 16720 7788 16727
rect 7801 16720 7853 16727
rect 5116 16685 5168 16706
rect 5182 16685 5234 16706
rect 5248 16685 5300 16706
rect 5314 16685 5366 16706
rect 5116 16654 5123 16685
rect 5123 16654 5162 16685
rect 5162 16654 5168 16685
rect 5182 16654 5196 16685
rect 5196 16654 5234 16685
rect 5248 16654 5269 16685
rect 5269 16654 5300 16685
rect 5314 16654 5342 16685
rect 5342 16654 5366 16685
rect 5380 16685 5432 16706
rect 5380 16654 5381 16685
rect 5381 16654 5415 16685
rect 5415 16654 5432 16685
rect 5446 16685 5498 16706
rect 5446 16654 5454 16685
rect 5454 16654 5488 16685
rect 5488 16654 5498 16685
rect 5512 16685 5564 16706
rect 5512 16654 5527 16685
rect 5527 16654 5561 16685
rect 5561 16654 5564 16685
rect 5578 16685 5630 16706
rect 5644 16685 5696 16706
rect 5710 16685 5762 16706
rect 5776 16685 5828 16706
rect 5842 16685 5894 16706
rect 5908 16685 5960 16706
rect 5974 16685 6026 16706
rect 6040 16685 6092 16706
rect 5578 16654 5600 16685
rect 5600 16654 5630 16685
rect 5644 16654 5673 16685
rect 5673 16654 5696 16685
rect 5710 16654 5746 16685
rect 5746 16654 5762 16685
rect 5776 16654 5780 16685
rect 5780 16654 5819 16685
rect 5819 16654 5828 16685
rect 5842 16654 5853 16685
rect 5853 16654 5892 16685
rect 5892 16654 5894 16685
rect 5908 16654 5926 16685
rect 5926 16654 5960 16685
rect 5974 16654 5999 16685
rect 5999 16654 6026 16685
rect 6040 16654 6072 16685
rect 6072 16654 6092 16685
rect 6106 16685 6158 16706
rect 6106 16654 6110 16685
rect 6110 16654 6144 16685
rect 6144 16654 6158 16685
rect 6172 16685 6224 16706
rect 6172 16654 6182 16685
rect 6182 16654 6216 16685
rect 6216 16654 6224 16685
rect 6238 16685 6290 16706
rect 6238 16654 6254 16685
rect 6254 16654 6288 16685
rect 6288 16654 6290 16685
rect 6304 16685 6356 16706
rect 6370 16685 6422 16706
rect 6436 16685 6488 16706
rect 6501 16685 6553 16706
rect 6566 16685 6618 16706
rect 6631 16685 6683 16706
rect 6696 16685 6748 16706
rect 6761 16685 6813 16706
rect 6304 16654 6326 16685
rect 6326 16654 6356 16685
rect 6370 16654 6398 16685
rect 6398 16654 6422 16685
rect 6436 16654 6470 16685
rect 6470 16654 6488 16685
rect 6501 16654 6504 16685
rect 6504 16654 6542 16685
rect 6542 16654 6553 16685
rect 6566 16654 6576 16685
rect 6576 16654 6614 16685
rect 6614 16654 6618 16685
rect 6631 16654 6648 16685
rect 6648 16654 6683 16685
rect 6696 16654 6720 16685
rect 6720 16654 6748 16685
rect 6761 16654 6792 16685
rect 6792 16654 6813 16685
rect 6826 16685 6878 16706
rect 6826 16654 6830 16685
rect 6830 16654 6864 16685
rect 6864 16654 6878 16685
rect 6891 16685 6943 16706
rect 6891 16654 6902 16685
rect 6902 16654 6936 16685
rect 6936 16654 6943 16685
rect 6956 16685 7008 16706
rect 6956 16654 6974 16685
rect 6974 16654 7008 16685
rect 7021 16685 7073 16706
rect 7086 16685 7138 16706
rect 7151 16685 7203 16706
rect 7216 16685 7268 16706
rect 7281 16685 7333 16706
rect 7346 16685 7398 16706
rect 7411 16685 7463 16706
rect 7021 16654 7046 16685
rect 7046 16654 7073 16685
rect 7086 16654 7118 16685
rect 7118 16654 7138 16685
rect 7151 16654 7152 16685
rect 7152 16654 7190 16685
rect 7190 16654 7203 16685
rect 7216 16654 7224 16685
rect 7224 16654 7262 16685
rect 7262 16654 7268 16685
rect 7281 16654 7296 16685
rect 7296 16654 7333 16685
rect 7346 16654 7368 16685
rect 7368 16654 7398 16685
rect 7411 16654 7440 16685
rect 7440 16654 7463 16685
rect 7476 16685 7528 16706
rect 7476 16654 7478 16685
rect 7478 16654 7512 16685
rect 7512 16654 7528 16685
rect 7541 16685 7593 16706
rect 7541 16654 7550 16685
rect 7550 16654 7584 16685
rect 7584 16654 7593 16685
rect 7606 16685 7658 16706
rect 7606 16654 7622 16685
rect 7622 16654 7656 16685
rect 7656 16654 7658 16685
rect 7671 16685 7723 16706
rect 7736 16685 7788 16706
rect 7801 16685 7853 16706
rect 7671 16654 7694 16685
rect 7694 16654 7723 16685
rect 7736 16654 7766 16685
rect 7766 16654 7788 16685
rect 7801 16654 7838 16685
rect 7838 16654 7853 16685
rect 5116 16609 5168 16640
rect 5182 16609 5234 16640
rect 5248 16609 5300 16640
rect 5314 16609 5366 16640
rect 5116 16588 5123 16609
rect 5123 16588 5162 16609
rect 5162 16588 5168 16609
rect 5182 16588 5196 16609
rect 5196 16588 5234 16609
rect 5248 16588 5269 16609
rect 5269 16588 5300 16609
rect 5314 16588 5342 16609
rect 5342 16588 5366 16609
rect 5380 16609 5432 16640
rect 5380 16588 5381 16609
rect 5381 16588 5415 16609
rect 5415 16588 5432 16609
rect 5446 16609 5498 16640
rect 5446 16588 5454 16609
rect 5454 16588 5488 16609
rect 5488 16588 5498 16609
rect 5512 16609 5564 16640
rect 5512 16588 5527 16609
rect 5527 16588 5561 16609
rect 5561 16588 5564 16609
rect 5578 16609 5630 16640
rect 5644 16609 5696 16640
rect 5710 16609 5762 16640
rect 5776 16609 5828 16640
rect 5842 16609 5894 16640
rect 5908 16609 5960 16640
rect 5974 16609 6026 16640
rect 6040 16609 6092 16640
rect 5578 16588 5600 16609
rect 5600 16588 5630 16609
rect 5644 16588 5673 16609
rect 5673 16588 5696 16609
rect 5710 16588 5746 16609
rect 5746 16588 5762 16609
rect 5776 16588 5780 16609
rect 5780 16588 5819 16609
rect 5819 16588 5828 16609
rect 5842 16588 5853 16609
rect 5853 16588 5892 16609
rect 5892 16588 5894 16609
rect 5908 16588 5926 16609
rect 5926 16588 5960 16609
rect 5974 16588 5999 16609
rect 5999 16588 6026 16609
rect 6040 16588 6072 16609
rect 6072 16588 6092 16609
rect 6106 16609 6158 16640
rect 6106 16588 6110 16609
rect 6110 16588 6144 16609
rect 6144 16588 6158 16609
rect 6172 16609 6224 16640
rect 6172 16588 6182 16609
rect 6182 16588 6216 16609
rect 6216 16588 6224 16609
rect 6238 16609 6290 16640
rect 6238 16588 6254 16609
rect 6254 16588 6288 16609
rect 6288 16588 6290 16609
rect 6304 16609 6356 16640
rect 6370 16609 6422 16640
rect 6436 16609 6488 16640
rect 6501 16609 6553 16640
rect 6566 16609 6618 16640
rect 6631 16609 6683 16640
rect 6696 16609 6748 16640
rect 6761 16609 6813 16640
rect 6304 16588 6326 16609
rect 6326 16588 6356 16609
rect 6370 16588 6398 16609
rect 6398 16588 6422 16609
rect 6436 16588 6470 16609
rect 6470 16588 6488 16609
rect 6501 16588 6504 16609
rect 6504 16588 6542 16609
rect 6542 16588 6553 16609
rect 6566 16588 6576 16609
rect 6576 16588 6614 16609
rect 6614 16588 6618 16609
rect 6631 16588 6648 16609
rect 6648 16588 6683 16609
rect 6696 16588 6720 16609
rect 6720 16588 6748 16609
rect 6761 16588 6792 16609
rect 6792 16588 6813 16609
rect 6826 16609 6878 16640
rect 6826 16588 6830 16609
rect 6830 16588 6864 16609
rect 6864 16588 6878 16609
rect 6891 16609 6943 16640
rect 6891 16588 6902 16609
rect 6902 16588 6936 16609
rect 6936 16588 6943 16609
rect 6956 16609 7008 16640
rect 6956 16588 6974 16609
rect 6974 16588 7008 16609
rect 7021 16609 7073 16640
rect 7086 16609 7138 16640
rect 7151 16609 7203 16640
rect 7216 16609 7268 16640
rect 7281 16609 7333 16640
rect 7346 16609 7398 16640
rect 7411 16609 7463 16640
rect 7021 16588 7046 16609
rect 7046 16588 7073 16609
rect 7086 16588 7118 16609
rect 7118 16588 7138 16609
rect 7151 16588 7152 16609
rect 7152 16588 7190 16609
rect 7190 16588 7203 16609
rect 7216 16588 7224 16609
rect 7224 16588 7262 16609
rect 7262 16588 7268 16609
rect 7281 16588 7296 16609
rect 7296 16588 7333 16609
rect 7346 16588 7368 16609
rect 7368 16588 7398 16609
rect 7411 16588 7440 16609
rect 7440 16588 7463 16609
rect 7476 16609 7528 16640
rect 7476 16588 7478 16609
rect 7478 16588 7512 16609
rect 7512 16588 7528 16609
rect 7541 16609 7593 16640
rect 7541 16588 7550 16609
rect 7550 16588 7584 16609
rect 7584 16588 7593 16609
rect 7606 16609 7658 16640
rect 7606 16588 7622 16609
rect 7622 16588 7656 16609
rect 7656 16588 7658 16609
rect 7671 16609 7723 16640
rect 7736 16609 7788 16640
rect 7801 16609 7853 16640
rect 7671 16588 7694 16609
rect 7694 16588 7723 16609
rect 7736 16588 7766 16609
rect 7766 16588 7788 16609
rect 7801 16588 7838 16609
rect 7838 16588 7853 16609
rect 5116 16533 5168 16574
rect 5182 16533 5234 16574
rect 5248 16533 5300 16574
rect 5314 16533 5366 16574
rect 5116 16522 5123 16533
rect 5123 16522 5162 16533
rect 5162 16522 5168 16533
rect 5182 16522 5196 16533
rect 5196 16522 5234 16533
rect 5248 16522 5269 16533
rect 5269 16522 5300 16533
rect 5314 16522 5342 16533
rect 5342 16522 5366 16533
rect 5380 16533 5432 16574
rect 5380 16522 5381 16533
rect 5381 16522 5415 16533
rect 5415 16522 5432 16533
rect 5446 16533 5498 16574
rect 5446 16522 5454 16533
rect 5454 16522 5488 16533
rect 5488 16522 5498 16533
rect 5512 16533 5564 16574
rect 5512 16522 5527 16533
rect 5527 16522 5561 16533
rect 5561 16522 5564 16533
rect 5578 16533 5630 16574
rect 5644 16533 5696 16574
rect 5710 16533 5762 16574
rect 5776 16533 5828 16574
rect 5842 16533 5894 16574
rect 5908 16533 5960 16574
rect 5974 16533 6026 16574
rect 6040 16533 6092 16574
rect 5578 16522 5600 16533
rect 5600 16522 5630 16533
rect 5644 16522 5673 16533
rect 5673 16522 5696 16533
rect 5710 16522 5746 16533
rect 5746 16522 5762 16533
rect 5776 16522 5780 16533
rect 5780 16522 5819 16533
rect 5819 16522 5828 16533
rect 5842 16522 5853 16533
rect 5853 16522 5892 16533
rect 5892 16522 5894 16533
rect 5908 16522 5926 16533
rect 5926 16522 5960 16533
rect 5974 16522 5999 16533
rect 5999 16522 6026 16533
rect 6040 16522 6072 16533
rect 6072 16522 6092 16533
rect 6106 16533 6158 16574
rect 6106 16522 6110 16533
rect 6110 16522 6144 16533
rect 6144 16522 6158 16533
rect 6172 16533 6224 16574
rect 6172 16522 6182 16533
rect 6182 16522 6216 16533
rect 6216 16522 6224 16533
rect 6238 16533 6290 16574
rect 6238 16522 6254 16533
rect 6254 16522 6288 16533
rect 6288 16522 6290 16533
rect 6304 16533 6356 16574
rect 6370 16533 6422 16574
rect 6436 16533 6488 16574
rect 6501 16533 6553 16574
rect 6566 16533 6618 16574
rect 6631 16533 6683 16574
rect 6696 16533 6748 16574
rect 6761 16533 6813 16574
rect 6304 16522 6326 16533
rect 6326 16522 6356 16533
rect 6370 16522 6398 16533
rect 6398 16522 6422 16533
rect 6436 16522 6470 16533
rect 6470 16522 6488 16533
rect 6501 16522 6504 16533
rect 6504 16522 6542 16533
rect 6542 16522 6553 16533
rect 6566 16522 6576 16533
rect 6576 16522 6614 16533
rect 6614 16522 6618 16533
rect 6631 16522 6648 16533
rect 6648 16522 6683 16533
rect 6696 16522 6720 16533
rect 6720 16522 6748 16533
rect 6761 16522 6792 16533
rect 6792 16522 6813 16533
rect 6826 16533 6878 16574
rect 6826 16522 6830 16533
rect 6830 16522 6864 16533
rect 6864 16522 6878 16533
rect 6891 16533 6943 16574
rect 6891 16522 6902 16533
rect 6902 16522 6936 16533
rect 6936 16522 6943 16533
rect 6956 16533 7008 16574
rect 6956 16522 6974 16533
rect 6974 16522 7008 16533
rect 7021 16533 7073 16574
rect 7086 16533 7138 16574
rect 7151 16533 7203 16574
rect 7216 16533 7268 16574
rect 7281 16533 7333 16574
rect 7346 16533 7398 16574
rect 7411 16533 7463 16574
rect 7021 16522 7046 16533
rect 7046 16522 7073 16533
rect 7086 16522 7118 16533
rect 7118 16522 7138 16533
rect 7151 16522 7152 16533
rect 7152 16522 7190 16533
rect 7190 16522 7203 16533
rect 7216 16522 7224 16533
rect 7224 16522 7262 16533
rect 7262 16522 7268 16533
rect 7281 16522 7296 16533
rect 7296 16522 7333 16533
rect 7346 16522 7368 16533
rect 7368 16522 7398 16533
rect 7411 16522 7440 16533
rect 7440 16522 7463 16533
rect 7476 16533 7528 16574
rect 7476 16522 7478 16533
rect 7478 16522 7512 16533
rect 7512 16522 7528 16533
rect 7541 16533 7593 16574
rect 7541 16522 7550 16533
rect 7550 16522 7584 16533
rect 7584 16522 7593 16533
rect 7606 16533 7658 16574
rect 7606 16522 7622 16533
rect 7622 16522 7656 16533
rect 7656 16522 7658 16533
rect 7671 16533 7723 16574
rect 7736 16533 7788 16574
rect 7801 16533 7853 16574
rect 7671 16522 7694 16533
rect 7694 16522 7723 16533
rect 7736 16522 7766 16533
rect 7766 16522 7788 16533
rect 7801 16522 7838 16533
rect 7838 16522 7853 16533
rect 5116 16499 5123 16508
rect 5123 16499 5162 16508
rect 5162 16499 5168 16508
rect 5182 16499 5196 16508
rect 5196 16499 5234 16508
rect 5248 16499 5269 16508
rect 5269 16499 5300 16508
rect 5314 16499 5342 16508
rect 5342 16499 5366 16508
rect 5116 16457 5168 16499
rect 5182 16457 5234 16499
rect 5248 16457 5300 16499
rect 5314 16457 5366 16499
rect 5116 16456 5123 16457
rect 5123 16456 5162 16457
rect 5162 16456 5168 16457
rect 5182 16456 5196 16457
rect 5196 16456 5234 16457
rect 5248 16456 5269 16457
rect 5269 16456 5300 16457
rect 5314 16456 5342 16457
rect 5342 16456 5366 16457
rect 5380 16499 5381 16508
rect 5381 16499 5415 16508
rect 5415 16499 5432 16508
rect 5380 16457 5432 16499
rect 5380 16456 5381 16457
rect 5381 16456 5415 16457
rect 5415 16456 5432 16457
rect 5446 16499 5454 16508
rect 5454 16499 5488 16508
rect 5488 16499 5498 16508
rect 5446 16457 5498 16499
rect 5446 16456 5454 16457
rect 5454 16456 5488 16457
rect 5488 16456 5498 16457
rect 5512 16499 5527 16508
rect 5527 16499 5561 16508
rect 5561 16499 5564 16508
rect 5512 16457 5564 16499
rect 5512 16456 5527 16457
rect 5527 16456 5561 16457
rect 5561 16456 5564 16457
rect 5578 16499 5600 16508
rect 5600 16499 5630 16508
rect 5644 16499 5673 16508
rect 5673 16499 5696 16508
rect 5710 16499 5746 16508
rect 5746 16499 5762 16508
rect 5776 16499 5780 16508
rect 5780 16499 5819 16508
rect 5819 16499 5828 16508
rect 5842 16499 5853 16508
rect 5853 16499 5892 16508
rect 5892 16499 5894 16508
rect 5908 16499 5926 16508
rect 5926 16499 5960 16508
rect 5974 16499 5999 16508
rect 5999 16499 6026 16508
rect 6040 16499 6072 16508
rect 6072 16499 6092 16508
rect 5578 16457 5630 16499
rect 5644 16457 5696 16499
rect 5710 16457 5762 16499
rect 5776 16457 5828 16499
rect 5842 16457 5894 16499
rect 5908 16457 5960 16499
rect 5974 16457 6026 16499
rect 6040 16457 6092 16499
rect 5578 16456 5600 16457
rect 5600 16456 5630 16457
rect 5644 16456 5673 16457
rect 5673 16456 5696 16457
rect 5710 16456 5746 16457
rect 5746 16456 5762 16457
rect 5776 16456 5780 16457
rect 5780 16456 5819 16457
rect 5819 16456 5828 16457
rect 5842 16456 5853 16457
rect 5853 16456 5892 16457
rect 5892 16456 5894 16457
rect 5908 16456 5926 16457
rect 5926 16456 5960 16457
rect 5974 16456 5999 16457
rect 5999 16456 6026 16457
rect 6040 16456 6072 16457
rect 6072 16456 6092 16457
rect 6106 16499 6110 16508
rect 6110 16499 6144 16508
rect 6144 16499 6158 16508
rect 6106 16457 6158 16499
rect 6106 16456 6110 16457
rect 6110 16456 6144 16457
rect 6144 16456 6158 16457
rect 6172 16499 6182 16508
rect 6182 16499 6216 16508
rect 6216 16499 6224 16508
rect 6172 16457 6224 16499
rect 6172 16456 6182 16457
rect 6182 16456 6216 16457
rect 6216 16456 6224 16457
rect 6238 16499 6254 16508
rect 6254 16499 6288 16508
rect 6288 16499 6290 16508
rect 6238 16457 6290 16499
rect 6238 16456 6254 16457
rect 6254 16456 6288 16457
rect 6288 16456 6290 16457
rect 6304 16499 6326 16508
rect 6326 16499 6356 16508
rect 6370 16499 6398 16508
rect 6398 16499 6422 16508
rect 6436 16499 6470 16508
rect 6470 16499 6488 16508
rect 6501 16499 6504 16508
rect 6504 16499 6542 16508
rect 6542 16499 6553 16508
rect 6566 16499 6576 16508
rect 6576 16499 6614 16508
rect 6614 16499 6618 16508
rect 6631 16499 6648 16508
rect 6648 16499 6683 16508
rect 6696 16499 6720 16508
rect 6720 16499 6748 16508
rect 6761 16499 6792 16508
rect 6792 16499 6813 16508
rect 6304 16457 6356 16499
rect 6370 16457 6422 16499
rect 6436 16457 6488 16499
rect 6501 16457 6553 16499
rect 6566 16457 6618 16499
rect 6631 16457 6683 16499
rect 6696 16457 6748 16499
rect 6761 16457 6813 16499
rect 6304 16456 6326 16457
rect 6326 16456 6356 16457
rect 6370 16456 6398 16457
rect 6398 16456 6422 16457
rect 6436 16456 6470 16457
rect 6470 16456 6488 16457
rect 6501 16456 6504 16457
rect 6504 16456 6542 16457
rect 6542 16456 6553 16457
rect 6566 16456 6576 16457
rect 6576 16456 6614 16457
rect 6614 16456 6618 16457
rect 6631 16456 6648 16457
rect 6648 16456 6683 16457
rect 6696 16456 6720 16457
rect 6720 16456 6748 16457
rect 6761 16456 6792 16457
rect 6792 16456 6813 16457
rect 6826 16499 6830 16508
rect 6830 16499 6864 16508
rect 6864 16499 6878 16508
rect 6826 16457 6878 16499
rect 6826 16456 6830 16457
rect 6830 16456 6864 16457
rect 6864 16456 6878 16457
rect 6891 16499 6902 16508
rect 6902 16499 6936 16508
rect 6936 16499 6943 16508
rect 6891 16457 6943 16499
rect 6891 16456 6902 16457
rect 6902 16456 6936 16457
rect 6936 16456 6943 16457
rect 6956 16499 6974 16508
rect 6974 16499 7008 16508
rect 6956 16457 7008 16499
rect 6956 16456 6974 16457
rect 6974 16456 7008 16457
rect 7021 16499 7046 16508
rect 7046 16499 7073 16508
rect 7086 16499 7118 16508
rect 7118 16499 7138 16508
rect 7151 16499 7152 16508
rect 7152 16499 7190 16508
rect 7190 16499 7203 16508
rect 7216 16499 7224 16508
rect 7224 16499 7262 16508
rect 7262 16499 7268 16508
rect 7281 16499 7296 16508
rect 7296 16499 7333 16508
rect 7346 16499 7368 16508
rect 7368 16499 7398 16508
rect 7411 16499 7440 16508
rect 7440 16499 7463 16508
rect 7021 16457 7073 16499
rect 7086 16457 7138 16499
rect 7151 16457 7203 16499
rect 7216 16457 7268 16499
rect 7281 16457 7333 16499
rect 7346 16457 7398 16499
rect 7411 16457 7463 16499
rect 7021 16456 7046 16457
rect 7046 16456 7073 16457
rect 7086 16456 7118 16457
rect 7118 16456 7138 16457
rect 7151 16456 7152 16457
rect 7152 16456 7190 16457
rect 7190 16456 7203 16457
rect 7216 16456 7224 16457
rect 7224 16456 7262 16457
rect 7262 16456 7268 16457
rect 7281 16456 7296 16457
rect 7296 16456 7333 16457
rect 7346 16456 7368 16457
rect 7368 16456 7398 16457
rect 7411 16456 7440 16457
rect 7440 16456 7463 16457
rect 7476 16499 7478 16508
rect 7478 16499 7512 16508
rect 7512 16499 7528 16508
rect 7476 16457 7528 16499
rect 7476 16456 7478 16457
rect 7478 16456 7512 16457
rect 7512 16456 7528 16457
rect 7541 16499 7550 16508
rect 7550 16499 7584 16508
rect 7584 16499 7593 16508
rect 7541 16457 7593 16499
rect 7541 16456 7550 16457
rect 7550 16456 7584 16457
rect 7584 16456 7593 16457
rect 7606 16499 7622 16508
rect 7622 16499 7656 16508
rect 7656 16499 7658 16508
rect 7606 16457 7658 16499
rect 7606 16456 7622 16457
rect 7622 16456 7656 16457
rect 7656 16456 7658 16457
rect 7671 16499 7694 16508
rect 7694 16499 7723 16508
rect 7736 16499 7766 16508
rect 7766 16499 7788 16508
rect 7801 16499 7838 16508
rect 7838 16499 7853 16508
rect 7671 16457 7723 16499
rect 7736 16457 7788 16499
rect 7801 16457 7853 16499
rect 7671 16456 7694 16457
rect 7694 16456 7723 16457
rect 7736 16456 7766 16457
rect 7766 16456 7788 16457
rect 7801 16456 7838 16457
rect 7838 16456 7853 16457
rect 5116 16423 5123 16442
rect 5123 16423 5162 16442
rect 5162 16423 5168 16442
rect 5182 16423 5196 16442
rect 5196 16423 5234 16442
rect 5248 16423 5269 16442
rect 5269 16423 5300 16442
rect 5314 16423 5342 16442
rect 5342 16423 5366 16442
rect 5116 16390 5168 16423
rect 5182 16390 5234 16423
rect 5248 16390 5300 16423
rect 5314 16390 5366 16423
rect 5380 16423 5381 16442
rect 5381 16423 5415 16442
rect 5415 16423 5432 16442
rect 5380 16390 5432 16423
rect 5446 16423 5454 16442
rect 5454 16423 5488 16442
rect 5488 16423 5498 16442
rect 5446 16390 5498 16423
rect 5512 16423 5527 16442
rect 5527 16423 5561 16442
rect 5561 16423 5564 16442
rect 5512 16390 5564 16423
rect 5578 16423 5600 16442
rect 5600 16423 5630 16442
rect 5644 16423 5673 16442
rect 5673 16423 5696 16442
rect 5710 16423 5746 16442
rect 5746 16423 5762 16442
rect 5776 16423 5780 16442
rect 5780 16423 5819 16442
rect 5819 16423 5828 16442
rect 5842 16423 5853 16442
rect 5853 16423 5892 16442
rect 5892 16423 5894 16442
rect 5908 16423 5926 16442
rect 5926 16423 5960 16442
rect 5974 16423 5999 16442
rect 5999 16423 6026 16442
rect 6040 16423 6072 16442
rect 6072 16423 6092 16442
rect 5578 16390 5630 16423
rect 5644 16390 5696 16423
rect 5710 16390 5762 16423
rect 5776 16390 5828 16423
rect 5842 16390 5894 16423
rect 5908 16390 5960 16423
rect 5974 16390 6026 16423
rect 6040 16390 6092 16423
rect 6106 16423 6110 16442
rect 6110 16423 6144 16442
rect 6144 16423 6158 16442
rect 6106 16390 6158 16423
rect 6172 16423 6182 16442
rect 6182 16423 6216 16442
rect 6216 16423 6224 16442
rect 6172 16390 6224 16423
rect 6238 16423 6254 16442
rect 6254 16423 6288 16442
rect 6288 16423 6290 16442
rect 6238 16390 6290 16423
rect 6304 16423 6326 16442
rect 6326 16423 6356 16442
rect 6370 16423 6398 16442
rect 6398 16423 6422 16442
rect 6436 16423 6470 16442
rect 6470 16423 6488 16442
rect 6501 16423 6504 16442
rect 6504 16423 6542 16442
rect 6542 16423 6553 16442
rect 6566 16423 6576 16442
rect 6576 16423 6614 16442
rect 6614 16423 6618 16442
rect 6631 16423 6648 16442
rect 6648 16423 6683 16442
rect 6696 16423 6720 16442
rect 6720 16423 6748 16442
rect 6761 16423 6792 16442
rect 6792 16423 6813 16442
rect 6304 16390 6356 16423
rect 6370 16390 6422 16423
rect 6436 16390 6488 16423
rect 6501 16390 6553 16423
rect 6566 16390 6618 16423
rect 6631 16390 6683 16423
rect 6696 16390 6748 16423
rect 6761 16390 6813 16423
rect 6826 16423 6830 16442
rect 6830 16423 6864 16442
rect 6864 16423 6878 16442
rect 6826 16390 6878 16423
rect 6891 16423 6902 16442
rect 6902 16423 6936 16442
rect 6936 16423 6943 16442
rect 6891 16390 6943 16423
rect 6956 16423 6974 16442
rect 6974 16423 7008 16442
rect 6956 16390 7008 16423
rect 7021 16423 7046 16442
rect 7046 16423 7073 16442
rect 7086 16423 7118 16442
rect 7118 16423 7138 16442
rect 7151 16423 7152 16442
rect 7152 16423 7190 16442
rect 7190 16423 7203 16442
rect 7216 16423 7224 16442
rect 7224 16423 7262 16442
rect 7262 16423 7268 16442
rect 7281 16423 7296 16442
rect 7296 16423 7333 16442
rect 7346 16423 7368 16442
rect 7368 16423 7398 16442
rect 7411 16423 7440 16442
rect 7440 16423 7463 16442
rect 7021 16390 7073 16423
rect 7086 16390 7138 16423
rect 7151 16390 7203 16423
rect 7216 16390 7268 16423
rect 7281 16390 7333 16423
rect 7346 16390 7398 16423
rect 7411 16390 7463 16423
rect 7476 16423 7478 16442
rect 7478 16423 7512 16442
rect 7512 16423 7528 16442
rect 7476 16390 7528 16423
rect 7541 16423 7550 16442
rect 7550 16423 7584 16442
rect 7584 16423 7593 16442
rect 7541 16390 7593 16423
rect 7606 16423 7622 16442
rect 7622 16423 7656 16442
rect 7656 16423 7658 16442
rect 7606 16390 7658 16423
rect 7671 16423 7694 16442
rect 7694 16423 7723 16442
rect 7736 16423 7766 16442
rect 7766 16423 7788 16442
rect 7801 16423 7838 16442
rect 7838 16423 7853 16442
rect 7671 16390 7723 16423
rect 7736 16390 7788 16423
rect 7801 16390 7853 16423
rect 5116 16347 5123 16376
rect 5123 16347 5162 16376
rect 5162 16347 5168 16376
rect 5182 16347 5196 16376
rect 5196 16347 5234 16376
rect 5248 16347 5269 16376
rect 5269 16347 5300 16376
rect 5314 16347 5342 16376
rect 5342 16347 5366 16376
rect 5116 16324 5168 16347
rect 5182 16324 5234 16347
rect 5248 16324 5300 16347
rect 5314 16324 5366 16347
rect 5380 16347 5381 16376
rect 5381 16347 5415 16376
rect 5415 16347 5432 16376
rect 5380 16324 5432 16347
rect 5446 16347 5454 16376
rect 5454 16347 5488 16376
rect 5488 16347 5498 16376
rect 5446 16324 5498 16347
rect 5512 16347 5527 16376
rect 5527 16347 5561 16376
rect 5561 16347 5564 16376
rect 5512 16324 5564 16347
rect 5578 16347 5600 16376
rect 5600 16347 5630 16376
rect 5644 16347 5673 16376
rect 5673 16347 5696 16376
rect 5710 16347 5746 16376
rect 5746 16347 5762 16376
rect 5776 16347 5780 16376
rect 5780 16347 5819 16376
rect 5819 16347 5828 16376
rect 5842 16347 5853 16376
rect 5853 16347 5892 16376
rect 5892 16347 5894 16376
rect 5908 16347 5926 16376
rect 5926 16347 5960 16376
rect 5974 16347 5999 16376
rect 5999 16347 6026 16376
rect 6040 16347 6072 16376
rect 6072 16347 6092 16376
rect 5578 16324 5630 16347
rect 5644 16324 5696 16347
rect 5710 16324 5762 16347
rect 5776 16324 5828 16347
rect 5842 16324 5894 16347
rect 5908 16324 5960 16347
rect 5974 16324 6026 16347
rect 6040 16324 6092 16347
rect 6106 16347 6110 16376
rect 6110 16347 6144 16376
rect 6144 16347 6158 16376
rect 6106 16324 6158 16347
rect 6172 16347 6182 16376
rect 6182 16347 6216 16376
rect 6216 16347 6224 16376
rect 6172 16324 6224 16347
rect 6238 16347 6254 16376
rect 6254 16347 6288 16376
rect 6288 16347 6290 16376
rect 6238 16324 6290 16347
rect 6304 16347 6326 16376
rect 6326 16347 6356 16376
rect 6370 16347 6398 16376
rect 6398 16347 6422 16376
rect 6436 16347 6470 16376
rect 6470 16347 6488 16376
rect 6501 16347 6504 16376
rect 6504 16347 6542 16376
rect 6542 16347 6553 16376
rect 6566 16347 6576 16376
rect 6576 16347 6614 16376
rect 6614 16347 6618 16376
rect 6631 16347 6648 16376
rect 6648 16347 6683 16376
rect 6696 16347 6720 16376
rect 6720 16347 6748 16376
rect 6761 16347 6792 16376
rect 6792 16347 6813 16376
rect 6304 16324 6356 16347
rect 6370 16324 6422 16347
rect 6436 16324 6488 16347
rect 6501 16324 6553 16347
rect 6566 16324 6618 16347
rect 6631 16324 6683 16347
rect 6696 16324 6748 16347
rect 6761 16324 6813 16347
rect 6826 16347 6830 16376
rect 6830 16347 6864 16376
rect 6864 16347 6878 16376
rect 6826 16324 6878 16347
rect 6891 16347 6902 16376
rect 6902 16347 6936 16376
rect 6936 16347 6943 16376
rect 6891 16324 6943 16347
rect 6956 16347 6974 16376
rect 6974 16347 7008 16376
rect 6956 16324 7008 16347
rect 7021 16347 7046 16376
rect 7046 16347 7073 16376
rect 7086 16347 7118 16376
rect 7118 16347 7138 16376
rect 7151 16347 7152 16376
rect 7152 16347 7190 16376
rect 7190 16347 7203 16376
rect 7216 16347 7224 16376
rect 7224 16347 7262 16376
rect 7262 16347 7268 16376
rect 7281 16347 7296 16376
rect 7296 16347 7333 16376
rect 7346 16347 7368 16376
rect 7368 16347 7398 16376
rect 7411 16347 7440 16376
rect 7440 16347 7463 16376
rect 7021 16324 7073 16347
rect 7086 16324 7138 16347
rect 7151 16324 7203 16347
rect 7216 16324 7268 16347
rect 7281 16324 7333 16347
rect 7346 16324 7398 16347
rect 7411 16324 7463 16347
rect 7476 16347 7478 16376
rect 7478 16347 7512 16376
rect 7512 16347 7528 16376
rect 7476 16324 7528 16347
rect 7541 16347 7550 16376
rect 7550 16347 7584 16376
rect 7584 16347 7593 16376
rect 7541 16324 7593 16347
rect 7606 16347 7622 16376
rect 7622 16347 7656 16376
rect 7656 16347 7658 16376
rect 7606 16324 7658 16347
rect 7671 16347 7694 16376
rect 7694 16347 7723 16376
rect 7736 16347 7766 16376
rect 7766 16347 7788 16376
rect 7801 16347 7838 16376
rect 7838 16347 7853 16376
rect 7671 16324 7723 16347
rect 7736 16324 7788 16347
rect 7801 16324 7853 16347
rect 5116 16305 5168 16310
rect 5182 16305 5234 16310
rect 5248 16305 5300 16310
rect 5314 16305 5366 16310
rect 5116 16271 5123 16305
rect 5123 16271 5162 16305
rect 5162 16271 5168 16305
rect 5182 16271 5196 16305
rect 5196 16271 5234 16305
rect 5248 16271 5269 16305
rect 5269 16271 5300 16305
rect 5314 16271 5342 16305
rect 5342 16271 5366 16305
rect 5116 16258 5168 16271
rect 5182 16258 5234 16271
rect 5248 16258 5300 16271
rect 5314 16258 5366 16271
rect 5380 16305 5432 16310
rect 5380 16271 5381 16305
rect 5381 16271 5415 16305
rect 5415 16271 5432 16305
rect 5380 16258 5432 16271
rect 5446 16305 5498 16310
rect 5446 16271 5454 16305
rect 5454 16271 5488 16305
rect 5488 16271 5498 16305
rect 5446 16258 5498 16271
rect 5512 16305 5564 16310
rect 5512 16271 5527 16305
rect 5527 16271 5561 16305
rect 5561 16271 5564 16305
rect 5512 16258 5564 16271
rect 5578 16305 5630 16310
rect 5644 16305 5696 16310
rect 5710 16305 5762 16310
rect 5776 16305 5828 16310
rect 5842 16305 5894 16310
rect 5908 16305 5960 16310
rect 5974 16305 6026 16310
rect 6040 16305 6092 16310
rect 5578 16271 5600 16305
rect 5600 16271 5630 16305
rect 5644 16271 5673 16305
rect 5673 16271 5696 16305
rect 5710 16271 5746 16305
rect 5746 16271 5762 16305
rect 5776 16271 5780 16305
rect 5780 16271 5819 16305
rect 5819 16271 5828 16305
rect 5842 16271 5853 16305
rect 5853 16271 5892 16305
rect 5892 16271 5894 16305
rect 5908 16271 5926 16305
rect 5926 16271 5960 16305
rect 5974 16271 5999 16305
rect 5999 16271 6026 16305
rect 6040 16271 6072 16305
rect 6072 16271 6092 16305
rect 5578 16258 5630 16271
rect 5644 16258 5696 16271
rect 5710 16258 5762 16271
rect 5776 16258 5828 16271
rect 5842 16258 5894 16271
rect 5908 16258 5960 16271
rect 5974 16258 6026 16271
rect 6040 16258 6092 16271
rect 6106 16305 6158 16310
rect 6106 16271 6110 16305
rect 6110 16271 6144 16305
rect 6144 16271 6158 16305
rect 6106 16258 6158 16271
rect 6172 16305 6224 16310
rect 6172 16271 6182 16305
rect 6182 16271 6216 16305
rect 6216 16271 6224 16305
rect 6172 16258 6224 16271
rect 6238 16305 6290 16310
rect 6238 16271 6254 16305
rect 6254 16271 6288 16305
rect 6288 16271 6290 16305
rect 6238 16258 6290 16271
rect 6304 16305 6356 16310
rect 6370 16305 6422 16310
rect 6436 16305 6488 16310
rect 6501 16305 6553 16310
rect 6566 16305 6618 16310
rect 6631 16305 6683 16310
rect 6696 16305 6748 16310
rect 6761 16305 6813 16310
rect 6304 16271 6326 16305
rect 6326 16271 6356 16305
rect 6370 16271 6398 16305
rect 6398 16271 6422 16305
rect 6436 16271 6470 16305
rect 6470 16271 6488 16305
rect 6501 16271 6504 16305
rect 6504 16271 6542 16305
rect 6542 16271 6553 16305
rect 6566 16271 6576 16305
rect 6576 16271 6614 16305
rect 6614 16271 6618 16305
rect 6631 16271 6648 16305
rect 6648 16271 6683 16305
rect 6696 16271 6720 16305
rect 6720 16271 6748 16305
rect 6761 16271 6792 16305
rect 6792 16271 6813 16305
rect 6304 16258 6356 16271
rect 6370 16258 6422 16271
rect 6436 16258 6488 16271
rect 6501 16258 6553 16271
rect 6566 16258 6618 16271
rect 6631 16258 6683 16271
rect 6696 16258 6748 16271
rect 6761 16258 6813 16271
rect 6826 16305 6878 16310
rect 6826 16271 6830 16305
rect 6830 16271 6864 16305
rect 6864 16271 6878 16305
rect 6826 16258 6878 16271
rect 6891 16305 6943 16310
rect 6891 16271 6902 16305
rect 6902 16271 6936 16305
rect 6936 16271 6943 16305
rect 6891 16258 6943 16271
rect 6956 16305 7008 16310
rect 6956 16271 6974 16305
rect 6974 16271 7008 16305
rect 6956 16258 7008 16271
rect 7021 16305 7073 16310
rect 7086 16305 7138 16310
rect 7151 16305 7203 16310
rect 7216 16305 7268 16310
rect 7281 16305 7333 16310
rect 7346 16305 7398 16310
rect 7411 16305 7463 16310
rect 7021 16271 7046 16305
rect 7046 16271 7073 16305
rect 7086 16271 7118 16305
rect 7118 16271 7138 16305
rect 7151 16271 7152 16305
rect 7152 16271 7190 16305
rect 7190 16271 7203 16305
rect 7216 16271 7224 16305
rect 7224 16271 7262 16305
rect 7262 16271 7268 16305
rect 7281 16271 7296 16305
rect 7296 16271 7333 16305
rect 7346 16271 7368 16305
rect 7368 16271 7398 16305
rect 7411 16271 7440 16305
rect 7440 16271 7463 16305
rect 7021 16258 7073 16271
rect 7086 16258 7138 16271
rect 7151 16258 7203 16271
rect 7216 16258 7268 16271
rect 7281 16258 7333 16271
rect 7346 16258 7398 16271
rect 7411 16258 7463 16271
rect 7476 16305 7528 16310
rect 7476 16271 7478 16305
rect 7478 16271 7512 16305
rect 7512 16271 7528 16305
rect 7476 16258 7528 16271
rect 7541 16305 7593 16310
rect 7541 16271 7550 16305
rect 7550 16271 7584 16305
rect 7584 16271 7593 16305
rect 7541 16258 7593 16271
rect 7606 16305 7658 16310
rect 7606 16271 7622 16305
rect 7622 16271 7656 16305
rect 7656 16271 7658 16305
rect 7606 16258 7658 16271
rect 7671 16305 7723 16310
rect 7736 16305 7788 16310
rect 7801 16305 7853 16310
rect 7671 16271 7694 16305
rect 7694 16271 7723 16305
rect 7736 16271 7766 16305
rect 7766 16271 7788 16305
rect 7801 16271 7838 16305
rect 7838 16271 7853 16305
rect 7671 16258 7723 16271
rect 7736 16258 7788 16271
rect 7801 16258 7853 16271
rect 5116 16229 5168 16244
rect 5182 16229 5234 16244
rect 5248 16229 5300 16244
rect 5314 16229 5366 16244
rect 5116 16195 5123 16229
rect 5123 16195 5162 16229
rect 5162 16195 5168 16229
rect 5182 16195 5196 16229
rect 5196 16195 5234 16229
rect 5248 16195 5269 16229
rect 5269 16195 5300 16229
rect 5314 16195 5342 16229
rect 5342 16195 5366 16229
rect 5116 16192 5168 16195
rect 5182 16192 5234 16195
rect 5248 16192 5300 16195
rect 5314 16192 5366 16195
rect 5380 16229 5432 16244
rect 5380 16195 5381 16229
rect 5381 16195 5415 16229
rect 5415 16195 5432 16229
rect 5380 16192 5432 16195
rect 5446 16229 5498 16244
rect 5446 16195 5454 16229
rect 5454 16195 5488 16229
rect 5488 16195 5498 16229
rect 5446 16192 5498 16195
rect 5512 16229 5564 16244
rect 5512 16195 5527 16229
rect 5527 16195 5561 16229
rect 5561 16195 5564 16229
rect 5512 16192 5564 16195
rect 5578 16229 5630 16244
rect 5644 16229 5696 16244
rect 5710 16229 5762 16244
rect 5776 16229 5828 16244
rect 5842 16229 5894 16244
rect 5908 16229 5960 16244
rect 5974 16229 6026 16244
rect 6040 16229 6092 16244
rect 5578 16195 5600 16229
rect 5600 16195 5630 16229
rect 5644 16195 5673 16229
rect 5673 16195 5696 16229
rect 5710 16195 5746 16229
rect 5746 16195 5762 16229
rect 5776 16195 5780 16229
rect 5780 16195 5819 16229
rect 5819 16195 5828 16229
rect 5842 16195 5853 16229
rect 5853 16195 5892 16229
rect 5892 16195 5894 16229
rect 5908 16195 5926 16229
rect 5926 16195 5960 16229
rect 5974 16195 5999 16229
rect 5999 16195 6026 16229
rect 6040 16195 6072 16229
rect 6072 16195 6092 16229
rect 5578 16192 5630 16195
rect 5644 16192 5696 16195
rect 5710 16192 5762 16195
rect 5776 16192 5828 16195
rect 5842 16192 5894 16195
rect 5908 16192 5960 16195
rect 5974 16192 6026 16195
rect 6040 16192 6092 16195
rect 6106 16229 6158 16244
rect 6106 16195 6110 16229
rect 6110 16195 6144 16229
rect 6144 16195 6158 16229
rect 6106 16192 6158 16195
rect 6172 16229 6224 16244
rect 6172 16195 6182 16229
rect 6182 16195 6216 16229
rect 6216 16195 6224 16229
rect 6172 16192 6224 16195
rect 6238 16229 6290 16244
rect 6238 16195 6254 16229
rect 6254 16195 6288 16229
rect 6288 16195 6290 16229
rect 6238 16192 6290 16195
rect 6304 16229 6356 16244
rect 6370 16229 6422 16244
rect 6436 16229 6488 16244
rect 6501 16229 6553 16244
rect 6566 16229 6618 16244
rect 6631 16229 6683 16244
rect 6696 16229 6748 16244
rect 6761 16229 6813 16244
rect 6304 16195 6326 16229
rect 6326 16195 6356 16229
rect 6370 16195 6398 16229
rect 6398 16195 6422 16229
rect 6436 16195 6470 16229
rect 6470 16195 6488 16229
rect 6501 16195 6504 16229
rect 6504 16195 6542 16229
rect 6542 16195 6553 16229
rect 6566 16195 6576 16229
rect 6576 16195 6614 16229
rect 6614 16195 6618 16229
rect 6631 16195 6648 16229
rect 6648 16195 6683 16229
rect 6696 16195 6720 16229
rect 6720 16195 6748 16229
rect 6761 16195 6792 16229
rect 6792 16195 6813 16229
rect 6304 16192 6356 16195
rect 6370 16192 6422 16195
rect 6436 16192 6488 16195
rect 6501 16192 6553 16195
rect 6566 16192 6618 16195
rect 6631 16192 6683 16195
rect 6696 16192 6748 16195
rect 6761 16192 6813 16195
rect 6826 16229 6878 16244
rect 6826 16195 6830 16229
rect 6830 16195 6864 16229
rect 6864 16195 6878 16229
rect 6826 16192 6878 16195
rect 6891 16229 6943 16244
rect 6891 16195 6902 16229
rect 6902 16195 6936 16229
rect 6936 16195 6943 16229
rect 6891 16192 6943 16195
rect 6956 16229 7008 16244
rect 6956 16195 6974 16229
rect 6974 16195 7008 16229
rect 6956 16192 7008 16195
rect 7021 16229 7073 16244
rect 7086 16229 7138 16244
rect 7151 16229 7203 16244
rect 7216 16229 7268 16244
rect 7281 16229 7333 16244
rect 7346 16229 7398 16244
rect 7411 16229 7463 16244
rect 7021 16195 7046 16229
rect 7046 16195 7073 16229
rect 7086 16195 7118 16229
rect 7118 16195 7138 16229
rect 7151 16195 7152 16229
rect 7152 16195 7190 16229
rect 7190 16195 7203 16229
rect 7216 16195 7224 16229
rect 7224 16195 7262 16229
rect 7262 16195 7268 16229
rect 7281 16195 7296 16229
rect 7296 16195 7333 16229
rect 7346 16195 7368 16229
rect 7368 16195 7398 16229
rect 7411 16195 7440 16229
rect 7440 16195 7463 16229
rect 7021 16192 7073 16195
rect 7086 16192 7138 16195
rect 7151 16192 7203 16195
rect 7216 16192 7268 16195
rect 7281 16192 7333 16195
rect 7346 16192 7398 16195
rect 7411 16192 7463 16195
rect 7476 16229 7528 16244
rect 7476 16195 7478 16229
rect 7478 16195 7512 16229
rect 7512 16195 7528 16229
rect 7476 16192 7528 16195
rect 7541 16229 7593 16244
rect 7541 16195 7550 16229
rect 7550 16195 7584 16229
rect 7584 16195 7593 16229
rect 7541 16192 7593 16195
rect 7606 16229 7658 16244
rect 7606 16195 7622 16229
rect 7622 16195 7656 16229
rect 7656 16195 7658 16229
rect 7606 16192 7658 16195
rect 7671 16229 7723 16244
rect 7736 16229 7788 16244
rect 7801 16229 7853 16244
rect 7671 16195 7694 16229
rect 7694 16195 7723 16229
rect 7736 16195 7766 16229
rect 7766 16195 7788 16229
rect 7801 16195 7838 16229
rect 7838 16195 7853 16229
rect 7671 16192 7723 16195
rect 7736 16192 7788 16195
rect 7801 16192 7853 16195
rect 5116 16153 5168 16178
rect 5182 16153 5234 16178
rect 5248 16153 5300 16178
rect 5314 16153 5366 16178
rect 5116 16126 5123 16153
rect 5123 16126 5162 16153
rect 5162 16126 5168 16153
rect 5182 16126 5196 16153
rect 5196 16126 5234 16153
rect 5248 16126 5269 16153
rect 5269 16126 5300 16153
rect 5314 16126 5342 16153
rect 5342 16126 5366 16153
rect 5380 16153 5432 16178
rect 5380 16126 5381 16153
rect 5381 16126 5415 16153
rect 5415 16126 5432 16153
rect 5446 16153 5498 16178
rect 5446 16126 5454 16153
rect 5454 16126 5488 16153
rect 5488 16126 5498 16153
rect 5512 16153 5564 16178
rect 5512 16126 5527 16153
rect 5527 16126 5561 16153
rect 5561 16126 5564 16153
rect 5578 16153 5630 16178
rect 5644 16153 5696 16178
rect 5710 16153 5762 16178
rect 5776 16153 5828 16178
rect 5842 16153 5894 16178
rect 5908 16153 5960 16178
rect 5974 16153 6026 16178
rect 6040 16153 6092 16178
rect 5578 16126 5600 16153
rect 5600 16126 5630 16153
rect 5644 16126 5673 16153
rect 5673 16126 5696 16153
rect 5710 16126 5746 16153
rect 5746 16126 5762 16153
rect 5776 16126 5780 16153
rect 5780 16126 5819 16153
rect 5819 16126 5828 16153
rect 5842 16126 5853 16153
rect 5853 16126 5892 16153
rect 5892 16126 5894 16153
rect 5908 16126 5926 16153
rect 5926 16126 5960 16153
rect 5974 16126 5999 16153
rect 5999 16126 6026 16153
rect 6040 16126 6072 16153
rect 6072 16126 6092 16153
rect 6106 16153 6158 16178
rect 6106 16126 6110 16153
rect 6110 16126 6144 16153
rect 6144 16126 6158 16153
rect 6172 16153 6224 16178
rect 6172 16126 6182 16153
rect 6182 16126 6216 16153
rect 6216 16126 6224 16153
rect 6238 16153 6290 16178
rect 6238 16126 6254 16153
rect 6254 16126 6288 16153
rect 6288 16126 6290 16153
rect 6304 16153 6356 16178
rect 6370 16153 6422 16178
rect 6436 16153 6488 16178
rect 6501 16153 6553 16178
rect 6566 16153 6618 16178
rect 6631 16153 6683 16178
rect 6696 16153 6748 16178
rect 6761 16153 6813 16178
rect 6304 16126 6326 16153
rect 6326 16126 6356 16153
rect 6370 16126 6398 16153
rect 6398 16126 6422 16153
rect 6436 16126 6470 16153
rect 6470 16126 6488 16153
rect 6501 16126 6504 16153
rect 6504 16126 6542 16153
rect 6542 16126 6553 16153
rect 6566 16126 6576 16153
rect 6576 16126 6614 16153
rect 6614 16126 6618 16153
rect 6631 16126 6648 16153
rect 6648 16126 6683 16153
rect 6696 16126 6720 16153
rect 6720 16126 6748 16153
rect 6761 16126 6792 16153
rect 6792 16126 6813 16153
rect 6826 16153 6878 16178
rect 6826 16126 6830 16153
rect 6830 16126 6864 16153
rect 6864 16126 6878 16153
rect 6891 16153 6943 16178
rect 6891 16126 6902 16153
rect 6902 16126 6936 16153
rect 6936 16126 6943 16153
rect 6956 16153 7008 16178
rect 6956 16126 6974 16153
rect 6974 16126 7008 16153
rect 7021 16153 7073 16178
rect 7086 16153 7138 16178
rect 7151 16153 7203 16178
rect 7216 16153 7268 16178
rect 7281 16153 7333 16178
rect 7346 16153 7398 16178
rect 7411 16153 7463 16178
rect 7021 16126 7046 16153
rect 7046 16126 7073 16153
rect 7086 16126 7118 16153
rect 7118 16126 7138 16153
rect 7151 16126 7152 16153
rect 7152 16126 7190 16153
rect 7190 16126 7203 16153
rect 7216 16126 7224 16153
rect 7224 16126 7262 16153
rect 7262 16126 7268 16153
rect 7281 16126 7296 16153
rect 7296 16126 7333 16153
rect 7346 16126 7368 16153
rect 7368 16126 7398 16153
rect 7411 16126 7440 16153
rect 7440 16126 7463 16153
rect 7476 16153 7528 16178
rect 7476 16126 7478 16153
rect 7478 16126 7512 16153
rect 7512 16126 7528 16153
rect 7541 16153 7593 16178
rect 7541 16126 7550 16153
rect 7550 16126 7584 16153
rect 7584 16126 7593 16153
rect 7606 16153 7658 16178
rect 7606 16126 7622 16153
rect 7622 16126 7656 16153
rect 7656 16126 7658 16153
rect 7671 16153 7723 16178
rect 7736 16153 7788 16178
rect 7801 16153 7853 16178
rect 7671 16126 7694 16153
rect 7694 16126 7723 16153
rect 7736 16126 7766 16153
rect 7766 16126 7788 16153
rect 7801 16126 7838 16153
rect 7838 16126 7853 16153
rect 5116 16077 5168 16112
rect 5182 16077 5234 16112
rect 5248 16077 5300 16112
rect 5314 16077 5366 16112
rect 5116 16060 5123 16077
rect 5123 16060 5162 16077
rect 5162 16060 5168 16077
rect 5182 16060 5196 16077
rect 5196 16060 5234 16077
rect 5248 16060 5269 16077
rect 5269 16060 5300 16077
rect 5314 16060 5342 16077
rect 5342 16060 5366 16077
rect 5380 16077 5432 16112
rect 5380 16060 5381 16077
rect 5381 16060 5415 16077
rect 5415 16060 5432 16077
rect 5446 16077 5498 16112
rect 5446 16060 5454 16077
rect 5454 16060 5488 16077
rect 5488 16060 5498 16077
rect 5512 16077 5564 16112
rect 5512 16060 5527 16077
rect 5527 16060 5561 16077
rect 5561 16060 5564 16077
rect 5578 16077 5630 16112
rect 5644 16077 5696 16112
rect 5710 16077 5762 16112
rect 5776 16077 5828 16112
rect 5842 16077 5894 16112
rect 5908 16077 5960 16112
rect 5974 16077 6026 16112
rect 6040 16077 6092 16112
rect 5578 16060 5600 16077
rect 5600 16060 5630 16077
rect 5644 16060 5673 16077
rect 5673 16060 5696 16077
rect 5710 16060 5746 16077
rect 5746 16060 5762 16077
rect 5776 16060 5780 16077
rect 5780 16060 5819 16077
rect 5819 16060 5828 16077
rect 5842 16060 5853 16077
rect 5853 16060 5892 16077
rect 5892 16060 5894 16077
rect 5908 16060 5926 16077
rect 5926 16060 5960 16077
rect 5974 16060 5999 16077
rect 5999 16060 6026 16077
rect 6040 16060 6072 16077
rect 6072 16060 6092 16077
rect 6106 16077 6158 16112
rect 6106 16060 6110 16077
rect 6110 16060 6144 16077
rect 6144 16060 6158 16077
rect 6172 16077 6224 16112
rect 6172 16060 6182 16077
rect 6182 16060 6216 16077
rect 6216 16060 6224 16077
rect 6238 16077 6290 16112
rect 6238 16060 6254 16077
rect 6254 16060 6288 16077
rect 6288 16060 6290 16077
rect 6304 16077 6356 16112
rect 6370 16077 6422 16112
rect 6436 16077 6488 16112
rect 6501 16077 6553 16112
rect 6566 16077 6618 16112
rect 6631 16077 6683 16112
rect 6696 16077 6748 16112
rect 6761 16077 6813 16112
rect 6304 16060 6326 16077
rect 6326 16060 6356 16077
rect 6370 16060 6398 16077
rect 6398 16060 6422 16077
rect 6436 16060 6470 16077
rect 6470 16060 6488 16077
rect 6501 16060 6504 16077
rect 6504 16060 6542 16077
rect 6542 16060 6553 16077
rect 6566 16060 6576 16077
rect 6576 16060 6614 16077
rect 6614 16060 6618 16077
rect 6631 16060 6648 16077
rect 6648 16060 6683 16077
rect 6696 16060 6720 16077
rect 6720 16060 6748 16077
rect 6761 16060 6792 16077
rect 6792 16060 6813 16077
rect 6826 16077 6878 16112
rect 6826 16060 6830 16077
rect 6830 16060 6864 16077
rect 6864 16060 6878 16077
rect 6891 16077 6943 16112
rect 6891 16060 6902 16077
rect 6902 16060 6936 16077
rect 6936 16060 6943 16077
rect 6956 16077 7008 16112
rect 6956 16060 6974 16077
rect 6974 16060 7008 16077
rect 7021 16077 7073 16112
rect 7086 16077 7138 16112
rect 7151 16077 7203 16112
rect 7216 16077 7268 16112
rect 7281 16077 7333 16112
rect 7346 16077 7398 16112
rect 7411 16077 7463 16112
rect 7021 16060 7046 16077
rect 7046 16060 7073 16077
rect 7086 16060 7118 16077
rect 7118 16060 7138 16077
rect 7151 16060 7152 16077
rect 7152 16060 7190 16077
rect 7190 16060 7203 16077
rect 7216 16060 7224 16077
rect 7224 16060 7262 16077
rect 7262 16060 7268 16077
rect 7281 16060 7296 16077
rect 7296 16060 7333 16077
rect 7346 16060 7368 16077
rect 7368 16060 7398 16077
rect 7411 16060 7440 16077
rect 7440 16060 7463 16077
rect 7476 16077 7528 16112
rect 7476 16060 7478 16077
rect 7478 16060 7512 16077
rect 7512 16060 7528 16077
rect 7541 16077 7593 16112
rect 7541 16060 7550 16077
rect 7550 16060 7584 16077
rect 7584 16060 7593 16077
rect 7606 16077 7658 16112
rect 7606 16060 7622 16077
rect 7622 16060 7656 16077
rect 7656 16060 7658 16077
rect 7671 16077 7723 16112
rect 7736 16077 7788 16112
rect 7801 16077 7853 16112
rect 7671 16060 7694 16077
rect 7694 16060 7723 16077
rect 7736 16060 7766 16077
rect 7766 16060 7788 16077
rect 7801 16060 7838 16077
rect 7838 16060 7853 16077
rect 5116 16043 5123 16046
rect 5123 16043 5162 16046
rect 5162 16043 5168 16046
rect 5182 16043 5196 16046
rect 5196 16043 5234 16046
rect 5248 16043 5269 16046
rect 5269 16043 5300 16046
rect 5314 16043 5342 16046
rect 5342 16043 5366 16046
rect 5116 16001 5168 16043
rect 5182 16001 5234 16043
rect 5248 16001 5300 16043
rect 5314 16001 5366 16043
rect 5116 15994 5123 16001
rect 5123 15994 5162 16001
rect 5162 15994 5168 16001
rect 5182 15994 5196 16001
rect 5196 15994 5234 16001
rect 5248 15994 5269 16001
rect 5269 15994 5300 16001
rect 5314 15994 5342 16001
rect 5342 15994 5366 16001
rect 5380 16043 5381 16046
rect 5381 16043 5415 16046
rect 5415 16043 5432 16046
rect 5380 16001 5432 16043
rect 5380 15994 5381 16001
rect 5381 15994 5415 16001
rect 5415 15994 5432 16001
rect 5446 16043 5454 16046
rect 5454 16043 5488 16046
rect 5488 16043 5498 16046
rect 5446 16001 5498 16043
rect 5446 15994 5454 16001
rect 5454 15994 5488 16001
rect 5488 15994 5498 16001
rect 5512 16043 5527 16046
rect 5527 16043 5561 16046
rect 5561 16043 5564 16046
rect 5512 16001 5564 16043
rect 5512 15994 5527 16001
rect 5527 15994 5561 16001
rect 5561 15994 5564 16001
rect 5578 16043 5600 16046
rect 5600 16043 5630 16046
rect 5644 16043 5673 16046
rect 5673 16043 5696 16046
rect 5710 16043 5746 16046
rect 5746 16043 5762 16046
rect 5776 16043 5780 16046
rect 5780 16043 5819 16046
rect 5819 16043 5828 16046
rect 5842 16043 5853 16046
rect 5853 16043 5892 16046
rect 5892 16043 5894 16046
rect 5908 16043 5926 16046
rect 5926 16043 5960 16046
rect 5974 16043 5999 16046
rect 5999 16043 6026 16046
rect 6040 16043 6072 16046
rect 6072 16043 6092 16046
rect 5578 16001 5630 16043
rect 5644 16001 5696 16043
rect 5710 16001 5762 16043
rect 5776 16001 5828 16043
rect 5842 16001 5894 16043
rect 5908 16001 5960 16043
rect 5974 16001 6026 16043
rect 6040 16001 6092 16043
rect 5578 15994 5600 16001
rect 5600 15994 5630 16001
rect 5644 15994 5673 16001
rect 5673 15994 5696 16001
rect 5710 15994 5746 16001
rect 5746 15994 5762 16001
rect 5776 15994 5780 16001
rect 5780 15994 5819 16001
rect 5819 15994 5828 16001
rect 5842 15994 5853 16001
rect 5853 15994 5892 16001
rect 5892 15994 5894 16001
rect 5908 15994 5926 16001
rect 5926 15994 5960 16001
rect 5974 15994 5999 16001
rect 5999 15994 6026 16001
rect 6040 15994 6072 16001
rect 6072 15994 6092 16001
rect 6106 16043 6110 16046
rect 6110 16043 6144 16046
rect 6144 16043 6158 16046
rect 6106 16001 6158 16043
rect 6106 15994 6110 16001
rect 6110 15994 6144 16001
rect 6144 15994 6158 16001
rect 6172 16043 6182 16046
rect 6182 16043 6216 16046
rect 6216 16043 6224 16046
rect 6172 16001 6224 16043
rect 6172 15994 6182 16001
rect 6182 15994 6216 16001
rect 6216 15994 6224 16001
rect 6238 16043 6254 16046
rect 6254 16043 6288 16046
rect 6288 16043 6290 16046
rect 6238 16001 6290 16043
rect 6238 15994 6254 16001
rect 6254 15994 6288 16001
rect 6288 15994 6290 16001
rect 6304 16043 6326 16046
rect 6326 16043 6356 16046
rect 6370 16043 6398 16046
rect 6398 16043 6422 16046
rect 6436 16043 6470 16046
rect 6470 16043 6488 16046
rect 6501 16043 6504 16046
rect 6504 16043 6542 16046
rect 6542 16043 6553 16046
rect 6566 16043 6576 16046
rect 6576 16043 6614 16046
rect 6614 16043 6618 16046
rect 6631 16043 6648 16046
rect 6648 16043 6683 16046
rect 6696 16043 6720 16046
rect 6720 16043 6748 16046
rect 6761 16043 6792 16046
rect 6792 16043 6813 16046
rect 6304 16001 6356 16043
rect 6370 16001 6422 16043
rect 6436 16001 6488 16043
rect 6501 16001 6553 16043
rect 6566 16001 6618 16043
rect 6631 16001 6683 16043
rect 6696 16001 6748 16043
rect 6761 16001 6813 16043
rect 6304 15994 6326 16001
rect 6326 15994 6356 16001
rect 6370 15994 6398 16001
rect 6398 15994 6422 16001
rect 6436 15994 6470 16001
rect 6470 15994 6488 16001
rect 6501 15994 6504 16001
rect 6504 15994 6542 16001
rect 6542 15994 6553 16001
rect 6566 15994 6576 16001
rect 6576 15994 6614 16001
rect 6614 15994 6618 16001
rect 6631 15994 6648 16001
rect 6648 15994 6683 16001
rect 6696 15994 6720 16001
rect 6720 15994 6748 16001
rect 6761 15994 6792 16001
rect 6792 15994 6813 16001
rect 6826 16043 6830 16046
rect 6830 16043 6864 16046
rect 6864 16043 6878 16046
rect 6826 16001 6878 16043
rect 6826 15994 6830 16001
rect 6830 15994 6864 16001
rect 6864 15994 6878 16001
rect 6891 16043 6902 16046
rect 6902 16043 6936 16046
rect 6936 16043 6943 16046
rect 6891 16001 6943 16043
rect 6891 15994 6902 16001
rect 6902 15994 6936 16001
rect 6936 15994 6943 16001
rect 6956 16043 6974 16046
rect 6974 16043 7008 16046
rect 6956 16001 7008 16043
rect 6956 15994 6974 16001
rect 6974 15994 7008 16001
rect 7021 16043 7046 16046
rect 7046 16043 7073 16046
rect 7086 16043 7118 16046
rect 7118 16043 7138 16046
rect 7151 16043 7152 16046
rect 7152 16043 7190 16046
rect 7190 16043 7203 16046
rect 7216 16043 7224 16046
rect 7224 16043 7262 16046
rect 7262 16043 7268 16046
rect 7281 16043 7296 16046
rect 7296 16043 7333 16046
rect 7346 16043 7368 16046
rect 7368 16043 7398 16046
rect 7411 16043 7440 16046
rect 7440 16043 7463 16046
rect 7021 16001 7073 16043
rect 7086 16001 7138 16043
rect 7151 16001 7203 16043
rect 7216 16001 7268 16043
rect 7281 16001 7333 16043
rect 7346 16001 7398 16043
rect 7411 16001 7463 16043
rect 7021 15994 7046 16001
rect 7046 15994 7073 16001
rect 7086 15994 7118 16001
rect 7118 15994 7138 16001
rect 7151 15994 7152 16001
rect 7152 15994 7190 16001
rect 7190 15994 7203 16001
rect 7216 15994 7224 16001
rect 7224 15994 7262 16001
rect 7262 15994 7268 16001
rect 7281 15994 7296 16001
rect 7296 15994 7333 16001
rect 7346 15994 7368 16001
rect 7368 15994 7398 16001
rect 7411 15994 7440 16001
rect 7440 15994 7463 16001
rect 7476 16043 7478 16046
rect 7478 16043 7512 16046
rect 7512 16043 7528 16046
rect 7476 16001 7528 16043
rect 7476 15994 7478 16001
rect 7478 15994 7512 16001
rect 7512 15994 7528 16001
rect 7541 16043 7550 16046
rect 7550 16043 7584 16046
rect 7584 16043 7593 16046
rect 7541 16001 7593 16043
rect 7541 15994 7550 16001
rect 7550 15994 7584 16001
rect 7584 15994 7593 16001
rect 7606 16043 7622 16046
rect 7622 16043 7656 16046
rect 7656 16043 7658 16046
rect 7606 16001 7658 16043
rect 7606 15994 7622 16001
rect 7622 15994 7656 16001
rect 7656 15994 7658 16001
rect 7671 16043 7694 16046
rect 7694 16043 7723 16046
rect 7736 16043 7766 16046
rect 7766 16043 7788 16046
rect 7801 16043 7838 16046
rect 7838 16043 7853 16046
rect 7671 16001 7723 16043
rect 7736 16001 7788 16043
rect 7801 16001 7853 16043
rect 7671 15994 7694 16001
rect 7694 15994 7723 16001
rect 7736 15994 7766 16001
rect 7766 15994 7788 16001
rect 7801 15994 7838 16001
rect 7838 15994 7853 16001
rect 8047 16941 8050 16973
rect 8050 16941 8084 16973
rect 8084 16941 8099 16973
rect 8047 16921 8099 16941
rect 8169 16965 8221 16973
rect 8169 16931 8184 16965
rect 8184 16931 8218 16965
rect 8218 16931 8221 16965
rect 8169 16921 8221 16931
rect 8047 16903 8099 16907
rect 8047 16869 8050 16903
rect 8050 16869 8084 16903
rect 8084 16869 8099 16903
rect 8047 16855 8099 16869
rect 8169 16893 8221 16907
rect 8169 16859 8184 16893
rect 8184 16859 8218 16893
rect 8218 16859 8221 16893
rect 8169 16855 8221 16859
rect 8047 16831 8099 16841
rect 8047 16797 8050 16831
rect 8050 16797 8084 16831
rect 8084 16797 8099 16831
rect 8047 16789 8099 16797
rect 8169 16821 8221 16841
rect 8169 16789 8184 16821
rect 8184 16789 8218 16821
rect 8218 16789 8221 16821
rect 8047 16759 8099 16775
rect 8047 16725 8050 16759
rect 8050 16725 8084 16759
rect 8084 16725 8099 16759
rect 8047 16723 8099 16725
rect 8169 16749 8221 16775
rect 8169 16723 8184 16749
rect 8184 16723 8218 16749
rect 8218 16723 8221 16749
rect 8047 16687 8099 16709
rect 8047 16657 8050 16687
rect 8050 16657 8084 16687
rect 8084 16657 8099 16687
rect 8169 16677 8221 16709
rect 8169 16657 8184 16677
rect 8184 16657 8218 16677
rect 8218 16657 8221 16677
rect 8047 16615 8099 16643
rect 8047 16591 8050 16615
rect 8050 16591 8084 16615
rect 8084 16591 8099 16615
rect 8169 16605 8221 16643
rect 8169 16591 8184 16605
rect 8184 16591 8218 16605
rect 8218 16591 8221 16605
rect 8047 16543 8099 16577
rect 8047 16525 8050 16543
rect 8050 16525 8084 16543
rect 8084 16525 8099 16543
rect 8169 16571 8184 16577
rect 8184 16571 8218 16577
rect 8218 16571 8221 16577
rect 8169 16533 8221 16571
rect 8169 16525 8184 16533
rect 8184 16525 8218 16533
rect 8218 16525 8221 16533
rect 8047 16509 8050 16511
rect 8050 16509 8084 16511
rect 8084 16509 8099 16511
rect 8047 16471 8099 16509
rect 8047 16459 8050 16471
rect 8050 16459 8084 16471
rect 8084 16459 8099 16471
rect 8169 16499 8184 16511
rect 8184 16499 8218 16511
rect 8218 16499 8221 16511
rect 8169 16461 8221 16499
rect 8169 16459 8184 16461
rect 8184 16459 8218 16461
rect 8218 16459 8221 16461
rect 8047 16437 8050 16445
rect 8050 16437 8084 16445
rect 8084 16437 8099 16445
rect 8047 16399 8099 16437
rect 8047 16393 8050 16399
rect 8050 16393 8084 16399
rect 8084 16393 8099 16399
rect 8169 16427 8184 16445
rect 8184 16427 8218 16445
rect 8218 16427 8221 16445
rect 8169 16393 8221 16427
rect 8047 16365 8050 16378
rect 8050 16365 8084 16378
rect 8084 16365 8099 16378
rect 8047 16327 8099 16365
rect 8047 16326 8050 16327
rect 8050 16326 8084 16327
rect 8084 16326 8099 16327
rect 8169 16355 8184 16378
rect 8184 16355 8218 16378
rect 8218 16355 8221 16378
rect 8169 16326 8221 16355
rect 8047 16293 8050 16311
rect 8050 16293 8084 16311
rect 8084 16293 8099 16311
rect 8047 16259 8099 16293
rect 8169 16283 8184 16311
rect 8184 16283 8218 16311
rect 8218 16283 8221 16311
rect 8169 16259 8221 16283
rect 8047 16221 8050 16244
rect 8050 16221 8084 16244
rect 8084 16221 8099 16244
rect 8047 16192 8099 16221
rect 8169 16211 8184 16244
rect 8184 16211 8218 16244
rect 8218 16211 8221 16244
rect 8169 16192 8221 16211
rect 8047 16149 8050 16177
rect 8050 16149 8084 16177
rect 8084 16149 8099 16177
rect 8047 16125 8099 16149
rect 8169 16173 8221 16177
rect 8169 16139 8184 16173
rect 8184 16139 8218 16173
rect 8218 16139 8221 16173
rect 8169 16125 8221 16139
rect 8047 16077 8050 16110
rect 8050 16077 8084 16110
rect 8084 16077 8099 16110
rect 8047 16058 8099 16077
rect 8169 16101 8221 16110
rect 8169 16067 8184 16101
rect 8184 16067 8218 16101
rect 8218 16067 8221 16101
rect 8169 16058 8221 16067
rect 8047 16039 8099 16043
rect 8047 16005 8050 16039
rect 8050 16005 8084 16039
rect 8084 16005 8099 16039
rect 8047 15991 8099 16005
rect 8169 16029 8221 16043
rect 8169 15995 8184 16029
rect 8184 15995 8218 16029
rect 8218 15995 8221 16029
rect 8169 15991 8221 15995
rect 2270 15420 2322 15456
rect 2270 15404 2276 15420
rect 2276 15404 2310 15420
rect 2310 15404 2322 15420
rect 2392 15420 2444 15456
rect 2392 15404 2410 15420
rect 2410 15404 2444 15420
rect 2270 15386 2276 15387
rect 2276 15386 2310 15387
rect 2310 15386 2322 15387
rect 2270 15348 2322 15386
rect 2270 15335 2276 15348
rect 2276 15335 2310 15348
rect 2310 15335 2322 15348
rect 2392 15386 2410 15387
rect 2410 15386 2444 15387
rect 2392 15348 2444 15386
rect 2392 15335 2410 15348
rect 2410 15335 2444 15348
rect 2270 15314 2276 15318
rect 2276 15314 2310 15318
rect 2310 15314 2322 15318
rect 2270 15276 2322 15314
rect 2270 15266 2276 15276
rect 2276 15266 2310 15276
rect 2310 15266 2322 15276
rect 2392 15314 2410 15318
rect 2410 15314 2444 15318
rect 2392 15276 2444 15314
rect 2392 15266 2410 15276
rect 2410 15266 2444 15276
rect 2270 15242 2276 15249
rect 2276 15242 2310 15249
rect 2310 15242 2322 15249
rect 2270 15204 2322 15242
rect 2270 15197 2276 15204
rect 2276 15197 2310 15204
rect 2310 15197 2322 15204
rect 2392 15242 2410 15249
rect 2410 15242 2444 15249
rect 2392 15204 2444 15242
rect 2392 15197 2410 15204
rect 2410 15197 2444 15204
rect 2270 15170 2276 15180
rect 2276 15170 2310 15180
rect 2310 15170 2322 15180
rect 2270 15132 2322 15170
rect 2270 15128 2276 15132
rect 2276 15128 2310 15132
rect 2310 15128 2322 15132
rect 2392 15170 2410 15180
rect 2410 15170 2444 15180
rect 2392 15132 2444 15170
rect 2392 15128 2410 15132
rect 2410 15128 2444 15132
rect 2270 15098 2276 15110
rect 2276 15098 2310 15110
rect 2310 15098 2322 15110
rect 2270 15060 2322 15098
rect 2270 15058 2276 15060
rect 2276 15058 2310 15060
rect 2310 15058 2322 15060
rect 2392 15098 2410 15110
rect 2410 15098 2444 15110
rect 2392 15060 2444 15098
rect 2392 15058 2410 15060
rect 2410 15058 2444 15060
rect 2270 15026 2276 15040
rect 2276 15026 2310 15040
rect 2310 15026 2322 15040
rect 2270 14988 2322 15026
rect 2392 15026 2410 15040
rect 2410 15026 2444 15040
rect 2392 14988 2444 15026
rect 2270 14954 2276 14970
rect 2276 14954 2310 14970
rect 2310 14954 2322 14970
rect 2270 14918 2322 14954
rect 2392 14954 2410 14970
rect 2410 14954 2444 14970
rect 2392 14918 2444 14954
rect 2270 14882 2276 14900
rect 2276 14882 2310 14900
rect 2310 14882 2322 14900
rect 2270 14848 2322 14882
rect 2392 14882 2410 14900
rect 2410 14882 2444 14900
rect 2392 14848 2444 14882
rect 2270 13442 2276 13456
rect 2276 13442 2310 13456
rect 2310 13442 2322 13456
rect 2270 13404 2322 13442
rect 2392 13442 2410 13456
rect 2410 13442 2444 13456
rect 2392 13404 2444 13442
rect 2270 13370 2276 13387
rect 2276 13370 2310 13387
rect 2310 13370 2322 13387
rect 2270 13335 2322 13370
rect 2392 13370 2410 13387
rect 2410 13370 2444 13387
rect 2392 13335 2444 13370
rect 2270 13298 2276 13318
rect 2276 13298 2310 13318
rect 2310 13298 2322 13318
rect 2270 13266 2322 13298
rect 2392 13298 2410 13318
rect 2410 13298 2444 13318
rect 2392 13266 2444 13298
rect 2270 13226 2276 13249
rect 2276 13226 2310 13249
rect 2310 13226 2322 13249
rect 2270 13197 2322 13226
rect 2392 13226 2410 13249
rect 2410 13226 2444 13249
rect 2392 13197 2444 13226
rect 2270 13154 2276 13180
rect 2276 13154 2310 13180
rect 2310 13154 2322 13180
rect 2270 13128 2322 13154
rect 2392 13154 2410 13180
rect 2410 13154 2444 13180
rect 2392 13128 2444 13154
rect 2270 13082 2276 13110
rect 2276 13082 2310 13110
rect 2310 13082 2322 13110
rect 2270 13058 2322 13082
rect 2392 13082 2410 13110
rect 2410 13082 2444 13110
rect 2392 13058 2444 13082
rect 2270 13010 2276 13040
rect 2276 13010 2310 13040
rect 2310 13010 2322 13040
rect 2270 12988 2322 13010
rect 2392 13010 2410 13040
rect 2410 13010 2444 13040
rect 2392 12988 2444 13010
rect 2270 12938 2276 12970
rect 2276 12938 2310 12970
rect 2310 12938 2322 12970
rect 2270 12918 2322 12938
rect 2392 12938 2410 12970
rect 2410 12938 2444 12970
rect 2392 12918 2444 12938
rect 2270 12866 2276 12900
rect 2276 12866 2310 12900
rect 2310 12866 2322 12900
rect 2270 12848 2322 12866
rect 2392 12866 2410 12900
rect 2410 12866 2444 12900
rect 2392 12848 2444 12866
rect 2270 11426 2276 11456
rect 2276 11426 2310 11456
rect 2310 11426 2322 11456
rect 2270 11404 2322 11426
rect 2392 11426 2410 11456
rect 2410 11426 2444 11456
rect 2392 11404 2444 11426
rect 2270 11354 2276 11387
rect 2276 11354 2310 11387
rect 2310 11354 2322 11387
rect 2270 11335 2322 11354
rect 2392 11354 2410 11387
rect 2410 11354 2444 11387
rect 2392 11335 2444 11354
rect 2270 11316 2322 11318
rect 2270 11282 2276 11316
rect 2276 11282 2310 11316
rect 2310 11282 2322 11316
rect 2270 11266 2322 11282
rect 2392 11316 2444 11318
rect 2392 11282 2410 11316
rect 2410 11282 2444 11316
rect 2392 11266 2444 11282
rect 2270 11244 2322 11249
rect 2270 11210 2276 11244
rect 2276 11210 2310 11244
rect 2310 11210 2322 11244
rect 2270 11197 2322 11210
rect 2392 11244 2444 11249
rect 2392 11210 2410 11244
rect 2410 11210 2444 11244
rect 2392 11197 2444 11210
rect 2270 11172 2322 11180
rect 2270 11138 2276 11172
rect 2276 11138 2310 11172
rect 2310 11138 2322 11172
rect 2270 11128 2322 11138
rect 2392 11172 2444 11180
rect 2392 11138 2410 11172
rect 2410 11138 2444 11172
rect 2392 11128 2444 11138
rect 2270 11100 2322 11110
rect 2270 11066 2276 11100
rect 2276 11066 2310 11100
rect 2310 11066 2322 11100
rect 2270 11058 2322 11066
rect 2392 11100 2444 11110
rect 2392 11066 2410 11100
rect 2410 11066 2444 11100
rect 2392 11058 2444 11066
rect 2270 11028 2322 11040
rect 2270 10994 2276 11028
rect 2276 10994 2310 11028
rect 2310 10994 2322 11028
rect 2270 10988 2322 10994
rect 2392 11028 2444 11040
rect 2392 10994 2410 11028
rect 2410 10994 2444 11028
rect 2392 10988 2444 10994
rect 2270 10956 2322 10970
rect 2270 10922 2276 10956
rect 2276 10922 2310 10956
rect 2310 10922 2322 10956
rect 2270 10918 2322 10922
rect 2392 10956 2444 10970
rect 2392 10922 2410 10956
rect 2410 10922 2444 10956
rect 2392 10918 2444 10922
rect 2270 10884 2322 10900
rect 2270 10850 2276 10884
rect 2276 10850 2310 10884
rect 2310 10850 2322 10884
rect 2270 10848 2322 10850
rect 2392 10884 2444 10900
rect 2392 10850 2410 10884
rect 2410 10850 2444 10884
rect 2392 10848 2444 10850
rect 2824 15446 2876 15452
rect 2824 15412 2830 15446
rect 2830 15412 2864 15446
rect 2864 15412 2876 15446
rect 2824 15400 2876 15412
rect 2890 15446 2942 15452
rect 2890 15412 2902 15446
rect 2902 15412 2936 15446
rect 2936 15412 2942 15446
rect 2890 15400 2942 15412
rect 2824 15373 2876 15383
rect 2824 15339 2830 15373
rect 2830 15339 2864 15373
rect 2864 15339 2876 15373
rect 2824 15331 2876 15339
rect 2890 15373 2942 15383
rect 2890 15339 2902 15373
rect 2902 15339 2936 15373
rect 2936 15339 2942 15373
rect 2890 15331 2942 15339
rect 2824 15300 2876 15314
rect 2824 15266 2830 15300
rect 2830 15266 2864 15300
rect 2864 15266 2876 15300
rect 2824 15262 2876 15266
rect 2890 15300 2942 15314
rect 2890 15266 2902 15300
rect 2902 15266 2936 15300
rect 2936 15266 2942 15300
rect 2890 15262 2942 15266
rect 2824 15227 2876 15245
rect 2824 15193 2830 15227
rect 2830 15193 2864 15227
rect 2864 15193 2876 15227
rect 2890 15227 2942 15245
rect 2890 15193 2902 15227
rect 2902 15193 2936 15227
rect 2936 15193 2942 15227
rect 2824 15154 2876 15176
rect 2890 15154 2942 15176
rect 2824 15124 2830 15154
rect 2830 15124 2876 15154
rect 2890 15124 2936 15154
rect 2936 15124 2942 15154
rect 2824 15055 2830 15107
rect 2830 15055 2876 15107
rect 2890 15055 2936 15107
rect 2936 15055 2942 15107
rect 2824 14986 2830 15038
rect 2830 14986 2876 15038
rect 2890 14986 2936 15038
rect 2936 14986 2942 15038
rect 2824 14916 2830 14968
rect 2830 14916 2876 14968
rect 2890 14916 2936 14968
rect 2936 14916 2942 14968
rect 2824 14846 2830 14898
rect 2830 14846 2876 14898
rect 2890 14846 2936 14898
rect 2936 14846 2942 14898
rect 3101 14662 3107 14714
rect 3107 14662 3153 14714
rect 3167 14662 3213 14714
rect 3213 14662 3219 14714
rect 3101 14593 3107 14645
rect 3107 14593 3153 14645
rect 3167 14593 3213 14645
rect 3213 14593 3219 14645
rect 3101 14524 3107 14576
rect 3107 14524 3153 14576
rect 3167 14524 3213 14576
rect 3213 14524 3219 14576
rect 3101 14455 3107 14507
rect 3107 14455 3153 14507
rect 3167 14455 3213 14507
rect 3213 14455 3219 14507
rect 3101 14386 3107 14438
rect 3107 14386 3153 14438
rect 3167 14386 3213 14438
rect 3213 14386 3219 14438
rect 3101 14316 3107 14368
rect 3107 14316 3153 14368
rect 3167 14316 3213 14368
rect 3213 14316 3219 14368
rect 3101 14246 3107 14298
rect 3107 14246 3153 14298
rect 3167 14246 3213 14298
rect 3213 14246 3219 14298
rect 3101 14176 3107 14228
rect 3107 14176 3153 14228
rect 3167 14176 3213 14228
rect 3213 14176 3219 14228
rect 3101 14112 3107 14158
rect 3107 14112 3153 14158
rect 3167 14112 3213 14158
rect 3213 14112 3219 14158
rect 3101 14106 3153 14112
rect 3167 14106 3219 14112
rect 3378 15446 3430 15452
rect 3378 15412 3384 15446
rect 3384 15412 3418 15446
rect 3418 15412 3430 15446
rect 3378 15400 3430 15412
rect 3444 15446 3496 15452
rect 3444 15412 3456 15446
rect 3456 15412 3490 15446
rect 3490 15412 3496 15446
rect 3444 15400 3496 15412
rect 3378 15373 3430 15383
rect 3378 15339 3384 15373
rect 3384 15339 3418 15373
rect 3418 15339 3430 15373
rect 3378 15331 3430 15339
rect 3444 15373 3496 15383
rect 3444 15339 3456 15373
rect 3456 15339 3490 15373
rect 3490 15339 3496 15373
rect 3444 15331 3496 15339
rect 3378 15300 3430 15314
rect 3378 15266 3384 15300
rect 3384 15266 3418 15300
rect 3418 15266 3430 15300
rect 3378 15262 3430 15266
rect 3444 15300 3496 15314
rect 3444 15266 3456 15300
rect 3456 15266 3490 15300
rect 3490 15266 3496 15300
rect 3444 15262 3496 15266
rect 3378 15227 3430 15245
rect 3378 15193 3384 15227
rect 3384 15193 3418 15227
rect 3418 15193 3430 15227
rect 3444 15227 3496 15245
rect 3444 15193 3456 15227
rect 3456 15193 3490 15227
rect 3490 15193 3496 15227
rect 3378 15154 3430 15176
rect 3444 15154 3496 15176
rect 3378 15124 3384 15154
rect 3384 15124 3430 15154
rect 3444 15124 3490 15154
rect 3490 15124 3496 15154
rect 3378 15055 3384 15107
rect 3384 15055 3430 15107
rect 3444 15055 3490 15107
rect 3490 15055 3496 15107
rect 3378 14986 3384 15038
rect 3384 14986 3430 15038
rect 3444 14986 3490 15038
rect 3490 14986 3496 15038
rect 3378 14916 3384 14968
rect 3384 14916 3430 14968
rect 3444 14916 3490 14968
rect 3490 14916 3496 14968
rect 3378 14846 3384 14898
rect 3384 14846 3430 14898
rect 3444 14846 3490 14898
rect 3490 14846 3496 14898
rect 3655 14662 3661 14714
rect 3661 14662 3707 14714
rect 3721 14662 3767 14714
rect 3767 14662 3773 14714
rect 3655 14593 3661 14645
rect 3661 14593 3707 14645
rect 3721 14593 3767 14645
rect 3767 14593 3773 14645
rect 3655 14524 3661 14576
rect 3661 14524 3707 14576
rect 3721 14524 3767 14576
rect 3767 14524 3773 14576
rect 3655 14455 3661 14507
rect 3661 14455 3707 14507
rect 3721 14455 3767 14507
rect 3767 14455 3773 14507
rect 3655 14386 3661 14438
rect 3661 14386 3707 14438
rect 3721 14386 3767 14438
rect 3767 14386 3773 14438
rect 3655 14316 3661 14368
rect 3661 14316 3707 14368
rect 3721 14316 3767 14368
rect 3767 14316 3773 14368
rect 3655 14246 3661 14298
rect 3661 14246 3707 14298
rect 3721 14246 3767 14298
rect 3767 14246 3773 14298
rect 3655 14176 3661 14228
rect 3661 14176 3707 14228
rect 3721 14176 3767 14228
rect 3767 14176 3773 14228
rect 3655 14112 3661 14158
rect 3661 14112 3707 14158
rect 3721 14112 3767 14158
rect 3767 14112 3773 14158
rect 3655 14106 3707 14112
rect 3721 14106 3773 14112
rect 3932 15446 3984 15452
rect 3932 15412 3938 15446
rect 3938 15412 3972 15446
rect 3972 15412 3984 15446
rect 3932 15400 3984 15412
rect 3998 15446 4050 15452
rect 3998 15412 4010 15446
rect 4010 15412 4044 15446
rect 4044 15412 4050 15446
rect 3998 15400 4050 15412
rect 3932 15373 3984 15383
rect 3932 15339 3938 15373
rect 3938 15339 3972 15373
rect 3972 15339 3984 15373
rect 3932 15331 3984 15339
rect 3998 15373 4050 15383
rect 3998 15339 4010 15373
rect 4010 15339 4044 15373
rect 4044 15339 4050 15373
rect 3998 15331 4050 15339
rect 3932 15300 3984 15314
rect 3932 15266 3938 15300
rect 3938 15266 3972 15300
rect 3972 15266 3984 15300
rect 3932 15262 3984 15266
rect 3998 15300 4050 15314
rect 3998 15266 4010 15300
rect 4010 15266 4044 15300
rect 4044 15266 4050 15300
rect 3998 15262 4050 15266
rect 3932 15227 3984 15245
rect 3932 15193 3938 15227
rect 3938 15193 3972 15227
rect 3972 15193 3984 15227
rect 3998 15227 4050 15245
rect 3998 15193 4010 15227
rect 4010 15193 4044 15227
rect 4044 15193 4050 15227
rect 3932 15154 3984 15176
rect 3998 15154 4050 15176
rect 3932 15124 3938 15154
rect 3938 15124 3984 15154
rect 3998 15124 4044 15154
rect 4044 15124 4050 15154
rect 3932 15055 3938 15107
rect 3938 15055 3984 15107
rect 3998 15055 4044 15107
rect 4044 15055 4050 15107
rect 3932 14986 3938 15038
rect 3938 14986 3984 15038
rect 3998 14986 4044 15038
rect 4044 14986 4050 15038
rect 3932 14916 3938 14968
rect 3938 14916 3984 14968
rect 3998 14916 4044 14968
rect 4044 14916 4050 14968
rect 3932 14846 3938 14898
rect 3938 14846 3984 14898
rect 3998 14846 4044 14898
rect 4044 14846 4050 14898
rect 4209 14662 4215 14714
rect 4215 14662 4261 14714
rect 4275 14662 4321 14714
rect 4321 14662 4327 14714
rect 4209 14593 4215 14645
rect 4215 14593 4261 14645
rect 4275 14593 4321 14645
rect 4321 14593 4327 14645
rect 4209 14524 4215 14576
rect 4215 14524 4261 14576
rect 4275 14524 4321 14576
rect 4321 14524 4327 14576
rect 4209 14455 4215 14507
rect 4215 14455 4261 14507
rect 4275 14455 4321 14507
rect 4321 14455 4327 14507
rect 4209 14386 4215 14438
rect 4215 14386 4261 14438
rect 4275 14386 4321 14438
rect 4321 14386 4327 14438
rect 4209 14316 4215 14368
rect 4215 14316 4261 14368
rect 4275 14316 4321 14368
rect 4321 14316 4327 14368
rect 4209 14246 4215 14298
rect 4215 14246 4261 14298
rect 4275 14246 4321 14298
rect 4321 14246 4327 14298
rect 4209 14176 4215 14228
rect 4215 14176 4261 14228
rect 4275 14176 4321 14228
rect 4321 14176 4327 14228
rect 4209 14112 4215 14158
rect 4215 14112 4261 14158
rect 4275 14112 4321 14158
rect 4321 14112 4327 14158
rect 4209 14106 4261 14112
rect 4275 14106 4327 14112
rect 4486 15446 4538 15452
rect 4486 15412 4492 15446
rect 4492 15412 4526 15446
rect 4526 15412 4538 15446
rect 4486 15400 4538 15412
rect 4552 15446 4604 15452
rect 4552 15412 4564 15446
rect 4564 15412 4598 15446
rect 4598 15412 4604 15446
rect 4552 15400 4604 15412
rect 4486 15373 4538 15383
rect 4486 15339 4492 15373
rect 4492 15339 4526 15373
rect 4526 15339 4538 15373
rect 4486 15331 4538 15339
rect 4552 15373 4604 15383
rect 4552 15339 4564 15373
rect 4564 15339 4598 15373
rect 4598 15339 4604 15373
rect 4552 15331 4604 15339
rect 4486 15300 4538 15314
rect 4486 15266 4492 15300
rect 4492 15266 4526 15300
rect 4526 15266 4538 15300
rect 4486 15262 4538 15266
rect 4552 15300 4604 15314
rect 4552 15266 4564 15300
rect 4564 15266 4598 15300
rect 4598 15266 4604 15300
rect 4552 15262 4604 15266
rect 4486 15227 4538 15245
rect 4486 15193 4492 15227
rect 4492 15193 4526 15227
rect 4526 15193 4538 15227
rect 4552 15227 4604 15245
rect 4552 15193 4564 15227
rect 4564 15193 4598 15227
rect 4598 15193 4604 15227
rect 4486 15154 4538 15176
rect 4552 15154 4604 15176
rect 4486 15124 4492 15154
rect 4492 15124 4538 15154
rect 4552 15124 4598 15154
rect 4598 15124 4604 15154
rect 4486 15055 4492 15107
rect 4492 15055 4538 15107
rect 4552 15055 4598 15107
rect 4598 15055 4604 15107
rect 4486 14986 4492 15038
rect 4492 14986 4538 15038
rect 4552 14986 4598 15038
rect 4598 14986 4604 15038
rect 4486 14916 4492 14968
rect 4492 14916 4538 14968
rect 4552 14916 4598 14968
rect 4598 14916 4604 14968
rect 4486 14846 4492 14898
rect 4492 14846 4538 14898
rect 4552 14846 4598 14898
rect 4598 14846 4604 14898
rect 4763 14662 4769 14714
rect 4769 14662 4815 14714
rect 4829 14662 4875 14714
rect 4875 14662 4881 14714
rect 4763 14593 4769 14645
rect 4769 14593 4815 14645
rect 4829 14593 4875 14645
rect 4875 14593 4881 14645
rect 4763 14524 4769 14576
rect 4769 14524 4815 14576
rect 4829 14524 4875 14576
rect 4875 14524 4881 14576
rect 4763 14455 4769 14507
rect 4769 14455 4815 14507
rect 4829 14455 4875 14507
rect 4875 14455 4881 14507
rect 4763 14386 4769 14438
rect 4769 14386 4815 14438
rect 4829 14386 4875 14438
rect 4875 14386 4881 14438
rect 4763 14316 4769 14368
rect 4769 14316 4815 14368
rect 4829 14316 4875 14368
rect 4875 14316 4881 14368
rect 4763 14246 4769 14298
rect 4769 14246 4815 14298
rect 4829 14246 4875 14298
rect 4875 14246 4881 14298
rect 4763 14176 4769 14228
rect 4769 14176 4815 14228
rect 4829 14176 4875 14228
rect 4875 14176 4881 14228
rect 4763 14112 4769 14158
rect 4769 14112 4815 14158
rect 4829 14112 4875 14158
rect 4875 14112 4881 14158
rect 4763 14106 4815 14112
rect 4829 14106 4881 14112
rect 5040 15446 5092 15452
rect 5040 15412 5046 15446
rect 5046 15412 5080 15446
rect 5080 15412 5092 15446
rect 5040 15400 5092 15412
rect 5106 15446 5158 15452
rect 5106 15412 5118 15446
rect 5118 15412 5152 15446
rect 5152 15412 5158 15446
rect 5106 15400 5158 15412
rect 5040 15373 5092 15383
rect 5040 15339 5046 15373
rect 5046 15339 5080 15373
rect 5080 15339 5092 15373
rect 5040 15331 5092 15339
rect 5106 15373 5158 15383
rect 5106 15339 5118 15373
rect 5118 15339 5152 15373
rect 5152 15339 5158 15373
rect 5106 15331 5158 15339
rect 5040 15300 5092 15314
rect 5040 15266 5046 15300
rect 5046 15266 5080 15300
rect 5080 15266 5092 15300
rect 5040 15262 5092 15266
rect 5106 15300 5158 15314
rect 5106 15266 5118 15300
rect 5118 15266 5152 15300
rect 5152 15266 5158 15300
rect 5106 15262 5158 15266
rect 5040 15227 5092 15245
rect 5040 15193 5046 15227
rect 5046 15193 5080 15227
rect 5080 15193 5092 15227
rect 5106 15227 5158 15245
rect 5106 15193 5118 15227
rect 5118 15193 5152 15227
rect 5152 15193 5158 15227
rect 5040 15154 5092 15176
rect 5106 15154 5158 15176
rect 5040 15124 5046 15154
rect 5046 15124 5092 15154
rect 5106 15124 5152 15154
rect 5152 15124 5158 15154
rect 5040 15055 5046 15107
rect 5046 15055 5092 15107
rect 5106 15055 5152 15107
rect 5152 15055 5158 15107
rect 5040 14986 5046 15038
rect 5046 14986 5092 15038
rect 5106 14986 5152 15038
rect 5152 14986 5158 15038
rect 5040 14916 5046 14968
rect 5046 14916 5092 14968
rect 5106 14916 5152 14968
rect 5152 14916 5158 14968
rect 5040 14846 5046 14898
rect 5046 14846 5092 14898
rect 5106 14846 5152 14898
rect 5152 14846 5158 14898
rect 5317 14662 5323 14714
rect 5323 14662 5369 14714
rect 5383 14662 5429 14714
rect 5429 14662 5435 14714
rect 5317 14593 5323 14645
rect 5323 14593 5369 14645
rect 5383 14593 5429 14645
rect 5429 14593 5435 14645
rect 5317 14524 5323 14576
rect 5323 14524 5369 14576
rect 5383 14524 5429 14576
rect 5429 14524 5435 14576
rect 5317 14455 5323 14507
rect 5323 14455 5369 14507
rect 5383 14455 5429 14507
rect 5429 14455 5435 14507
rect 5317 14386 5323 14438
rect 5323 14386 5369 14438
rect 5383 14386 5429 14438
rect 5429 14386 5435 14438
rect 5317 14316 5323 14368
rect 5323 14316 5369 14368
rect 5383 14316 5429 14368
rect 5429 14316 5435 14368
rect 5317 14246 5323 14298
rect 5323 14246 5369 14298
rect 5383 14246 5429 14298
rect 5429 14246 5435 14298
rect 5317 14176 5323 14228
rect 5323 14176 5369 14228
rect 5383 14176 5429 14228
rect 5429 14176 5435 14228
rect 5317 14112 5323 14158
rect 5323 14112 5369 14158
rect 5383 14112 5429 14158
rect 5429 14112 5435 14158
rect 5317 14106 5369 14112
rect 5383 14106 5435 14112
rect 5594 15446 5646 15452
rect 5594 15412 5600 15446
rect 5600 15412 5634 15446
rect 5634 15412 5646 15446
rect 5594 15400 5646 15412
rect 5660 15446 5712 15452
rect 5660 15412 5672 15446
rect 5672 15412 5706 15446
rect 5706 15412 5712 15446
rect 5660 15400 5712 15412
rect 5594 15373 5646 15383
rect 5594 15339 5600 15373
rect 5600 15339 5634 15373
rect 5634 15339 5646 15373
rect 5594 15331 5646 15339
rect 5660 15373 5712 15383
rect 5660 15339 5672 15373
rect 5672 15339 5706 15373
rect 5706 15339 5712 15373
rect 5660 15331 5712 15339
rect 5594 15300 5646 15314
rect 5594 15266 5600 15300
rect 5600 15266 5634 15300
rect 5634 15266 5646 15300
rect 5594 15262 5646 15266
rect 5660 15300 5712 15314
rect 5660 15266 5672 15300
rect 5672 15266 5706 15300
rect 5706 15266 5712 15300
rect 5660 15262 5712 15266
rect 5594 15227 5646 15245
rect 5594 15193 5600 15227
rect 5600 15193 5634 15227
rect 5634 15193 5646 15227
rect 5660 15227 5712 15245
rect 5660 15193 5672 15227
rect 5672 15193 5706 15227
rect 5706 15193 5712 15227
rect 5594 15154 5646 15176
rect 5660 15154 5712 15176
rect 5594 15124 5600 15154
rect 5600 15124 5646 15154
rect 5660 15124 5706 15154
rect 5706 15124 5712 15154
rect 5594 15055 5600 15107
rect 5600 15055 5646 15107
rect 5660 15055 5706 15107
rect 5706 15055 5712 15107
rect 5594 14986 5600 15038
rect 5600 14986 5646 15038
rect 5660 14986 5706 15038
rect 5706 14986 5712 15038
rect 5594 14916 5600 14968
rect 5600 14916 5646 14968
rect 5660 14916 5706 14968
rect 5706 14916 5712 14968
rect 5594 14846 5600 14898
rect 5600 14846 5646 14898
rect 5660 14846 5706 14898
rect 5706 14846 5712 14898
rect 5871 14662 5877 14714
rect 5877 14662 5923 14714
rect 5937 14662 5983 14714
rect 5983 14662 5989 14714
rect 5871 14593 5877 14645
rect 5877 14593 5923 14645
rect 5937 14593 5983 14645
rect 5983 14593 5989 14645
rect 5871 14524 5877 14576
rect 5877 14524 5923 14576
rect 5937 14524 5983 14576
rect 5983 14524 5989 14576
rect 5871 14455 5877 14507
rect 5877 14455 5923 14507
rect 5937 14455 5983 14507
rect 5983 14455 5989 14507
rect 5871 14386 5877 14438
rect 5877 14386 5923 14438
rect 5937 14386 5983 14438
rect 5983 14386 5989 14438
rect 5871 14316 5877 14368
rect 5877 14316 5923 14368
rect 5937 14316 5983 14368
rect 5983 14316 5989 14368
rect 5871 14246 5877 14298
rect 5877 14246 5923 14298
rect 5937 14246 5983 14298
rect 5983 14246 5989 14298
rect 5871 14176 5877 14228
rect 5877 14176 5923 14228
rect 5937 14176 5983 14228
rect 5983 14176 5989 14228
rect 5871 14112 5877 14158
rect 5877 14112 5923 14158
rect 5937 14112 5983 14158
rect 5983 14112 5989 14158
rect 5871 14106 5923 14112
rect 5937 14106 5989 14112
rect 6148 15446 6200 15452
rect 6148 15412 6154 15446
rect 6154 15412 6188 15446
rect 6188 15412 6200 15446
rect 6148 15400 6200 15412
rect 6214 15446 6266 15452
rect 6214 15412 6226 15446
rect 6226 15412 6260 15446
rect 6260 15412 6266 15446
rect 6214 15400 6266 15412
rect 6148 15373 6200 15383
rect 6148 15339 6154 15373
rect 6154 15339 6188 15373
rect 6188 15339 6200 15373
rect 6148 15331 6200 15339
rect 6214 15373 6266 15383
rect 6214 15339 6226 15373
rect 6226 15339 6260 15373
rect 6260 15339 6266 15373
rect 6214 15331 6266 15339
rect 6148 15300 6200 15314
rect 6148 15266 6154 15300
rect 6154 15266 6188 15300
rect 6188 15266 6200 15300
rect 6148 15262 6200 15266
rect 6214 15300 6266 15314
rect 6214 15266 6226 15300
rect 6226 15266 6260 15300
rect 6260 15266 6266 15300
rect 6214 15262 6266 15266
rect 6148 15227 6200 15245
rect 6148 15193 6154 15227
rect 6154 15193 6188 15227
rect 6188 15193 6200 15227
rect 6214 15227 6266 15245
rect 6214 15193 6226 15227
rect 6226 15193 6260 15227
rect 6260 15193 6266 15227
rect 6148 15154 6200 15176
rect 6214 15154 6266 15176
rect 6148 15124 6154 15154
rect 6154 15124 6200 15154
rect 6214 15124 6260 15154
rect 6260 15124 6266 15154
rect 6148 15055 6154 15107
rect 6154 15055 6200 15107
rect 6214 15055 6260 15107
rect 6260 15055 6266 15107
rect 6148 14986 6154 15038
rect 6154 14986 6200 15038
rect 6214 14986 6260 15038
rect 6260 14986 6266 15038
rect 6148 14916 6154 14968
rect 6154 14916 6200 14968
rect 6214 14916 6260 14968
rect 6260 14916 6266 14968
rect 6148 14846 6154 14898
rect 6154 14846 6200 14898
rect 6214 14846 6260 14898
rect 6260 14846 6266 14898
rect 6425 14662 6431 14714
rect 6431 14662 6477 14714
rect 6491 14662 6537 14714
rect 6537 14662 6543 14714
rect 6425 14593 6431 14645
rect 6431 14593 6477 14645
rect 6491 14593 6537 14645
rect 6537 14593 6543 14645
rect 6425 14524 6431 14576
rect 6431 14524 6477 14576
rect 6491 14524 6537 14576
rect 6537 14524 6543 14576
rect 6425 14455 6431 14507
rect 6431 14455 6477 14507
rect 6491 14455 6537 14507
rect 6537 14455 6543 14507
rect 6425 14386 6431 14438
rect 6431 14386 6477 14438
rect 6491 14386 6537 14438
rect 6537 14386 6543 14438
rect 6425 14316 6431 14368
rect 6431 14316 6477 14368
rect 6491 14316 6537 14368
rect 6537 14316 6543 14368
rect 6425 14246 6431 14298
rect 6431 14246 6477 14298
rect 6491 14246 6537 14298
rect 6537 14246 6543 14298
rect 6425 14176 6431 14228
rect 6431 14176 6477 14228
rect 6491 14176 6537 14228
rect 6537 14176 6543 14228
rect 6425 14112 6431 14158
rect 6431 14112 6477 14158
rect 6491 14112 6537 14158
rect 6537 14112 6543 14158
rect 6425 14106 6477 14112
rect 6491 14106 6543 14112
rect 6702 15446 6754 15452
rect 6702 15412 6708 15446
rect 6708 15412 6742 15446
rect 6742 15412 6754 15446
rect 6702 15400 6754 15412
rect 6768 15446 6820 15452
rect 6768 15412 6780 15446
rect 6780 15412 6814 15446
rect 6814 15412 6820 15446
rect 6768 15400 6820 15412
rect 6702 15373 6754 15383
rect 6702 15339 6708 15373
rect 6708 15339 6742 15373
rect 6742 15339 6754 15373
rect 6702 15331 6754 15339
rect 6768 15373 6820 15383
rect 6768 15339 6780 15373
rect 6780 15339 6814 15373
rect 6814 15339 6820 15373
rect 6768 15331 6820 15339
rect 6702 15300 6754 15314
rect 6702 15266 6708 15300
rect 6708 15266 6742 15300
rect 6742 15266 6754 15300
rect 6702 15262 6754 15266
rect 6768 15300 6820 15314
rect 6768 15266 6780 15300
rect 6780 15266 6814 15300
rect 6814 15266 6820 15300
rect 6768 15262 6820 15266
rect 6702 15227 6754 15245
rect 6702 15193 6708 15227
rect 6708 15193 6742 15227
rect 6742 15193 6754 15227
rect 6768 15227 6820 15245
rect 6768 15193 6780 15227
rect 6780 15193 6814 15227
rect 6814 15193 6820 15227
rect 6702 15154 6754 15176
rect 6768 15154 6820 15176
rect 6702 15124 6708 15154
rect 6708 15124 6754 15154
rect 6768 15124 6814 15154
rect 6814 15124 6820 15154
rect 6702 15055 6708 15107
rect 6708 15055 6754 15107
rect 6768 15055 6814 15107
rect 6814 15055 6820 15107
rect 6702 14986 6708 15038
rect 6708 14986 6754 15038
rect 6768 14986 6814 15038
rect 6814 14986 6820 15038
rect 6702 14916 6708 14968
rect 6708 14916 6754 14968
rect 6768 14916 6814 14968
rect 6814 14916 6820 14968
rect 6702 14846 6708 14898
rect 6708 14846 6754 14898
rect 6768 14846 6814 14898
rect 6814 14846 6820 14898
rect 6979 14662 6985 14714
rect 6985 14662 7031 14714
rect 7045 14662 7091 14714
rect 7091 14662 7097 14714
rect 6979 14593 6985 14645
rect 6985 14593 7031 14645
rect 7045 14593 7091 14645
rect 7091 14593 7097 14645
rect 6979 14524 6985 14576
rect 6985 14524 7031 14576
rect 7045 14524 7091 14576
rect 7091 14524 7097 14576
rect 6979 14455 6985 14507
rect 6985 14455 7031 14507
rect 7045 14455 7091 14507
rect 7091 14455 7097 14507
rect 6979 14386 6985 14438
rect 6985 14386 7031 14438
rect 7045 14386 7091 14438
rect 7091 14386 7097 14438
rect 6979 14316 6985 14368
rect 6985 14316 7031 14368
rect 7045 14316 7091 14368
rect 7091 14316 7097 14368
rect 6979 14246 6985 14298
rect 6985 14246 7031 14298
rect 7045 14246 7091 14298
rect 7091 14246 7097 14298
rect 6979 14176 6985 14228
rect 6985 14176 7031 14228
rect 7045 14176 7091 14228
rect 7091 14176 7097 14228
rect 6979 14112 6985 14158
rect 6985 14112 7031 14158
rect 7045 14112 7091 14158
rect 7091 14112 7097 14158
rect 6979 14106 7031 14112
rect 7045 14106 7097 14112
rect 7256 15446 7308 15452
rect 7256 15412 7262 15446
rect 7262 15412 7296 15446
rect 7296 15412 7308 15446
rect 7256 15400 7308 15412
rect 7322 15446 7374 15452
rect 7322 15412 7334 15446
rect 7334 15412 7368 15446
rect 7368 15412 7374 15446
rect 7322 15400 7374 15412
rect 7256 15373 7308 15383
rect 7256 15339 7262 15373
rect 7262 15339 7296 15373
rect 7296 15339 7308 15373
rect 7256 15331 7308 15339
rect 7322 15373 7374 15383
rect 7322 15339 7334 15373
rect 7334 15339 7368 15373
rect 7368 15339 7374 15373
rect 7322 15331 7374 15339
rect 7256 15300 7308 15314
rect 7256 15266 7262 15300
rect 7262 15266 7296 15300
rect 7296 15266 7308 15300
rect 7256 15262 7308 15266
rect 7322 15300 7374 15314
rect 7322 15266 7334 15300
rect 7334 15266 7368 15300
rect 7368 15266 7374 15300
rect 7322 15262 7374 15266
rect 7256 15227 7308 15245
rect 7256 15193 7262 15227
rect 7262 15193 7296 15227
rect 7296 15193 7308 15227
rect 7322 15227 7374 15245
rect 7322 15193 7334 15227
rect 7334 15193 7368 15227
rect 7368 15193 7374 15227
rect 7256 15154 7308 15176
rect 7322 15154 7374 15176
rect 7256 15124 7262 15154
rect 7262 15124 7308 15154
rect 7322 15124 7368 15154
rect 7368 15124 7374 15154
rect 7256 15055 7262 15107
rect 7262 15055 7308 15107
rect 7322 15055 7368 15107
rect 7368 15055 7374 15107
rect 7256 14986 7262 15038
rect 7262 14986 7308 15038
rect 7322 14986 7368 15038
rect 7368 14986 7374 15038
rect 7256 14916 7262 14968
rect 7262 14916 7308 14968
rect 7322 14916 7368 14968
rect 7368 14916 7374 14968
rect 7256 14846 7262 14898
rect 7262 14846 7308 14898
rect 7322 14846 7368 14898
rect 7368 14846 7374 14898
rect 7533 14662 7539 14714
rect 7539 14662 7585 14714
rect 7599 14662 7645 14714
rect 7645 14662 7651 14714
rect 7533 14593 7539 14645
rect 7539 14593 7585 14645
rect 7599 14593 7645 14645
rect 7645 14593 7651 14645
rect 7533 14524 7539 14576
rect 7539 14524 7585 14576
rect 7599 14524 7645 14576
rect 7645 14524 7651 14576
rect 7533 14455 7539 14507
rect 7539 14455 7585 14507
rect 7599 14455 7645 14507
rect 7645 14455 7651 14507
rect 7533 14386 7539 14438
rect 7539 14386 7585 14438
rect 7599 14386 7645 14438
rect 7645 14386 7651 14438
rect 7533 14316 7539 14368
rect 7539 14316 7585 14368
rect 7599 14316 7645 14368
rect 7645 14316 7651 14368
rect 7533 14246 7539 14298
rect 7539 14246 7585 14298
rect 7599 14246 7645 14298
rect 7645 14246 7651 14298
rect 7533 14176 7539 14228
rect 7539 14176 7585 14228
rect 7599 14176 7645 14228
rect 7645 14176 7651 14228
rect 7533 14112 7539 14158
rect 7539 14112 7585 14158
rect 7599 14112 7645 14158
rect 7645 14112 7651 14158
rect 7533 14106 7585 14112
rect 7599 14106 7651 14112
rect 7810 15446 7862 15452
rect 7810 15412 7816 15446
rect 7816 15412 7850 15446
rect 7850 15412 7862 15446
rect 7810 15400 7862 15412
rect 7876 15446 7928 15452
rect 7876 15412 7888 15446
rect 7888 15412 7922 15446
rect 7922 15412 7928 15446
rect 7876 15400 7928 15412
rect 7810 15373 7862 15383
rect 7810 15339 7816 15373
rect 7816 15339 7850 15373
rect 7850 15339 7862 15373
rect 7810 15331 7862 15339
rect 7876 15373 7928 15383
rect 7876 15339 7888 15373
rect 7888 15339 7922 15373
rect 7922 15339 7928 15373
rect 7876 15331 7928 15339
rect 7810 15300 7862 15314
rect 7810 15266 7816 15300
rect 7816 15266 7850 15300
rect 7850 15266 7862 15300
rect 7810 15262 7862 15266
rect 7876 15300 7928 15314
rect 7876 15266 7888 15300
rect 7888 15266 7922 15300
rect 7922 15266 7928 15300
rect 7876 15262 7928 15266
rect 7810 15227 7862 15245
rect 7810 15193 7816 15227
rect 7816 15193 7850 15227
rect 7850 15193 7862 15227
rect 7876 15227 7928 15245
rect 7876 15193 7888 15227
rect 7888 15193 7922 15227
rect 7922 15193 7928 15227
rect 7810 15154 7862 15176
rect 7876 15154 7928 15176
rect 7810 15124 7816 15154
rect 7816 15124 7862 15154
rect 7876 15124 7922 15154
rect 7922 15124 7928 15154
rect 7810 15055 7816 15107
rect 7816 15055 7862 15107
rect 7876 15055 7922 15107
rect 7922 15055 7928 15107
rect 7810 14986 7816 15038
rect 7816 14986 7862 15038
rect 7876 14986 7922 15038
rect 7922 14986 7928 15038
rect 7810 14916 7816 14968
rect 7816 14916 7862 14968
rect 7876 14916 7922 14968
rect 7922 14916 7928 14968
rect 7810 14846 7816 14898
rect 7816 14846 7862 14898
rect 7876 14846 7922 14898
rect 7922 14846 7928 14898
rect 8047 15429 8050 15456
rect 8050 15429 8084 15456
rect 8084 15429 8099 15456
rect 8047 15404 8099 15429
rect 8169 15453 8221 15456
rect 8169 15419 8184 15453
rect 8184 15419 8218 15453
rect 8218 15419 8221 15453
rect 8169 15404 8221 15419
rect 8047 15357 8050 15387
rect 8050 15357 8084 15387
rect 8084 15357 8099 15387
rect 8047 15335 8099 15357
rect 8169 15381 8221 15387
rect 8169 15347 8184 15381
rect 8184 15347 8218 15381
rect 8218 15347 8221 15381
rect 8169 15335 8221 15347
rect 8047 15285 8050 15318
rect 8050 15285 8084 15318
rect 8084 15285 8099 15318
rect 8047 15266 8099 15285
rect 8169 15309 8221 15318
rect 8169 15275 8184 15309
rect 8184 15275 8218 15309
rect 8218 15275 8221 15309
rect 8169 15266 8221 15275
rect 8047 15247 8099 15249
rect 8047 15213 8050 15247
rect 8050 15213 8084 15247
rect 8084 15213 8099 15247
rect 8047 15197 8099 15213
rect 8169 15237 8221 15249
rect 8169 15203 8184 15237
rect 8184 15203 8218 15237
rect 8218 15203 8221 15237
rect 8169 15197 8221 15203
rect 8047 15175 8099 15180
rect 8047 15141 8050 15175
rect 8050 15141 8084 15175
rect 8084 15141 8099 15175
rect 8047 15128 8099 15141
rect 8169 15165 8221 15180
rect 8169 15131 8184 15165
rect 8184 15131 8218 15165
rect 8218 15131 8221 15165
rect 8169 15128 8221 15131
rect 8047 15103 8099 15110
rect 8047 15069 8050 15103
rect 8050 15069 8084 15103
rect 8084 15069 8099 15103
rect 8047 15058 8099 15069
rect 8169 15093 8221 15110
rect 8169 15059 8184 15093
rect 8184 15059 8218 15093
rect 8218 15059 8221 15093
rect 8169 15058 8221 15059
rect 8047 15031 8099 15040
rect 8047 14997 8050 15031
rect 8050 14997 8084 15031
rect 8084 14997 8099 15031
rect 8047 14988 8099 14997
rect 8169 15021 8221 15040
rect 8169 14988 8184 15021
rect 8184 14988 8218 15021
rect 8218 14988 8221 15021
rect 8047 14959 8099 14970
rect 8047 14925 8050 14959
rect 8050 14925 8084 14959
rect 8084 14925 8099 14959
rect 8047 14918 8099 14925
rect 8169 14949 8221 14970
rect 8169 14918 8184 14949
rect 8184 14918 8218 14949
rect 8218 14918 8221 14949
rect 8047 14887 8099 14900
rect 8047 14853 8050 14887
rect 8050 14853 8084 14887
rect 8084 14853 8099 14887
rect 8047 14848 8099 14853
rect 8169 14877 8221 14900
rect 8169 14848 8184 14877
rect 8184 14848 8218 14877
rect 8218 14848 8221 14877
rect 2824 13446 2876 13452
rect 2824 13412 2830 13446
rect 2830 13412 2864 13446
rect 2864 13412 2876 13446
rect 2824 13400 2876 13412
rect 2890 13446 2942 13452
rect 2890 13412 2902 13446
rect 2902 13412 2936 13446
rect 2936 13412 2942 13446
rect 2890 13400 2942 13412
rect 2824 13373 2876 13383
rect 2824 13339 2830 13373
rect 2830 13339 2864 13373
rect 2864 13339 2876 13373
rect 2824 13331 2876 13339
rect 2890 13373 2942 13383
rect 2890 13339 2902 13373
rect 2902 13339 2936 13373
rect 2936 13339 2942 13373
rect 2890 13331 2942 13339
rect 2824 13300 2876 13314
rect 2824 13266 2830 13300
rect 2830 13266 2864 13300
rect 2864 13266 2876 13300
rect 2824 13262 2876 13266
rect 2890 13300 2942 13314
rect 2890 13266 2902 13300
rect 2902 13266 2936 13300
rect 2936 13266 2942 13300
rect 2890 13262 2942 13266
rect 2824 13227 2876 13245
rect 2824 13193 2830 13227
rect 2830 13193 2864 13227
rect 2864 13193 2876 13227
rect 2890 13227 2942 13245
rect 2890 13193 2902 13227
rect 2902 13193 2936 13227
rect 2936 13193 2942 13227
rect 2824 13154 2876 13176
rect 2890 13154 2942 13176
rect 2824 13124 2830 13154
rect 2830 13124 2876 13154
rect 2890 13124 2936 13154
rect 2936 13124 2942 13154
rect 2824 13055 2830 13107
rect 2830 13055 2876 13107
rect 2890 13055 2936 13107
rect 2936 13055 2942 13107
rect 2824 12986 2830 13038
rect 2830 12986 2876 13038
rect 2890 12986 2936 13038
rect 2936 12986 2942 13038
rect 2824 12916 2830 12968
rect 2830 12916 2876 12968
rect 2890 12916 2936 12968
rect 2936 12916 2942 12968
rect 2824 12846 2830 12898
rect 2830 12846 2876 12898
rect 2890 12846 2936 12898
rect 2936 12846 2942 12898
rect 3101 12662 3107 12714
rect 3107 12662 3153 12714
rect 3167 12662 3213 12714
rect 3213 12662 3219 12714
rect 3101 12593 3107 12645
rect 3107 12593 3153 12645
rect 3167 12593 3213 12645
rect 3213 12593 3219 12645
rect 3101 12524 3107 12576
rect 3107 12524 3153 12576
rect 3167 12524 3213 12576
rect 3213 12524 3219 12576
rect 3101 12455 3107 12507
rect 3107 12455 3153 12507
rect 3167 12455 3213 12507
rect 3213 12455 3219 12507
rect 3101 12386 3107 12438
rect 3107 12386 3153 12438
rect 3167 12386 3213 12438
rect 3213 12386 3219 12438
rect 3101 12316 3107 12368
rect 3107 12316 3153 12368
rect 3167 12316 3213 12368
rect 3213 12316 3219 12368
rect 3101 12246 3107 12298
rect 3107 12246 3153 12298
rect 3167 12246 3213 12298
rect 3213 12246 3219 12298
rect 3101 12176 3107 12228
rect 3107 12176 3153 12228
rect 3167 12176 3213 12228
rect 3213 12176 3219 12228
rect 3101 12112 3107 12158
rect 3107 12112 3153 12158
rect 3167 12112 3213 12158
rect 3213 12112 3219 12158
rect 3101 12106 3153 12112
rect 3167 12106 3219 12112
rect 3378 13446 3430 13452
rect 3378 13412 3384 13446
rect 3384 13412 3418 13446
rect 3418 13412 3430 13446
rect 3378 13400 3430 13412
rect 3444 13446 3496 13452
rect 3444 13412 3456 13446
rect 3456 13412 3490 13446
rect 3490 13412 3496 13446
rect 3444 13400 3496 13412
rect 3378 13373 3430 13383
rect 3378 13339 3384 13373
rect 3384 13339 3418 13373
rect 3418 13339 3430 13373
rect 3378 13331 3430 13339
rect 3444 13373 3496 13383
rect 3444 13339 3456 13373
rect 3456 13339 3490 13373
rect 3490 13339 3496 13373
rect 3444 13331 3496 13339
rect 3378 13300 3430 13314
rect 3378 13266 3384 13300
rect 3384 13266 3418 13300
rect 3418 13266 3430 13300
rect 3378 13262 3430 13266
rect 3444 13300 3496 13314
rect 3444 13266 3456 13300
rect 3456 13266 3490 13300
rect 3490 13266 3496 13300
rect 3444 13262 3496 13266
rect 3378 13227 3430 13245
rect 3378 13193 3384 13227
rect 3384 13193 3418 13227
rect 3418 13193 3430 13227
rect 3444 13227 3496 13245
rect 3444 13193 3456 13227
rect 3456 13193 3490 13227
rect 3490 13193 3496 13227
rect 3378 13154 3430 13176
rect 3444 13154 3496 13176
rect 3378 13124 3384 13154
rect 3384 13124 3430 13154
rect 3444 13124 3490 13154
rect 3490 13124 3496 13154
rect 3378 13055 3384 13107
rect 3384 13055 3430 13107
rect 3444 13055 3490 13107
rect 3490 13055 3496 13107
rect 3378 12986 3384 13038
rect 3384 12986 3430 13038
rect 3444 12986 3490 13038
rect 3490 12986 3496 13038
rect 3378 12916 3384 12968
rect 3384 12916 3430 12968
rect 3444 12916 3490 12968
rect 3490 12916 3496 12968
rect 3378 12846 3384 12898
rect 3384 12846 3430 12898
rect 3444 12846 3490 12898
rect 3490 12846 3496 12898
rect 3655 12662 3661 12714
rect 3661 12662 3707 12714
rect 3721 12662 3767 12714
rect 3767 12662 3773 12714
rect 3655 12593 3661 12645
rect 3661 12593 3707 12645
rect 3721 12593 3767 12645
rect 3767 12593 3773 12645
rect 3655 12524 3661 12576
rect 3661 12524 3707 12576
rect 3721 12524 3767 12576
rect 3767 12524 3773 12576
rect 3655 12455 3661 12507
rect 3661 12455 3707 12507
rect 3721 12455 3767 12507
rect 3767 12455 3773 12507
rect 3655 12386 3661 12438
rect 3661 12386 3707 12438
rect 3721 12386 3767 12438
rect 3767 12386 3773 12438
rect 3655 12316 3661 12368
rect 3661 12316 3707 12368
rect 3721 12316 3767 12368
rect 3767 12316 3773 12368
rect 3655 12246 3661 12298
rect 3661 12246 3707 12298
rect 3721 12246 3767 12298
rect 3767 12246 3773 12298
rect 3655 12176 3661 12228
rect 3661 12176 3707 12228
rect 3721 12176 3767 12228
rect 3767 12176 3773 12228
rect 3655 12112 3661 12158
rect 3661 12112 3707 12158
rect 3721 12112 3767 12158
rect 3767 12112 3773 12158
rect 3655 12106 3707 12112
rect 3721 12106 3773 12112
rect 3932 13446 3984 13452
rect 3932 13412 3938 13446
rect 3938 13412 3972 13446
rect 3972 13412 3984 13446
rect 3932 13400 3984 13412
rect 3998 13446 4050 13452
rect 3998 13412 4010 13446
rect 4010 13412 4044 13446
rect 4044 13412 4050 13446
rect 3998 13400 4050 13412
rect 3932 13373 3984 13383
rect 3932 13339 3938 13373
rect 3938 13339 3972 13373
rect 3972 13339 3984 13373
rect 3932 13331 3984 13339
rect 3998 13373 4050 13383
rect 3998 13339 4010 13373
rect 4010 13339 4044 13373
rect 4044 13339 4050 13373
rect 3998 13331 4050 13339
rect 3932 13300 3984 13314
rect 3932 13266 3938 13300
rect 3938 13266 3972 13300
rect 3972 13266 3984 13300
rect 3932 13262 3984 13266
rect 3998 13300 4050 13314
rect 3998 13266 4010 13300
rect 4010 13266 4044 13300
rect 4044 13266 4050 13300
rect 3998 13262 4050 13266
rect 3932 13227 3984 13245
rect 3932 13193 3938 13227
rect 3938 13193 3972 13227
rect 3972 13193 3984 13227
rect 3998 13227 4050 13245
rect 3998 13193 4010 13227
rect 4010 13193 4044 13227
rect 4044 13193 4050 13227
rect 3932 13154 3984 13176
rect 3998 13154 4050 13176
rect 3932 13124 3938 13154
rect 3938 13124 3984 13154
rect 3998 13124 4044 13154
rect 4044 13124 4050 13154
rect 3932 13055 3938 13107
rect 3938 13055 3984 13107
rect 3998 13055 4044 13107
rect 4044 13055 4050 13107
rect 3932 12986 3938 13038
rect 3938 12986 3984 13038
rect 3998 12986 4044 13038
rect 4044 12986 4050 13038
rect 3932 12916 3938 12968
rect 3938 12916 3984 12968
rect 3998 12916 4044 12968
rect 4044 12916 4050 12968
rect 3932 12846 3938 12898
rect 3938 12846 3984 12898
rect 3998 12846 4044 12898
rect 4044 12846 4050 12898
rect 4209 12662 4215 12714
rect 4215 12662 4261 12714
rect 4275 12662 4321 12714
rect 4321 12662 4327 12714
rect 4209 12593 4215 12645
rect 4215 12593 4261 12645
rect 4275 12593 4321 12645
rect 4321 12593 4327 12645
rect 4209 12524 4215 12576
rect 4215 12524 4261 12576
rect 4275 12524 4321 12576
rect 4321 12524 4327 12576
rect 4209 12455 4215 12507
rect 4215 12455 4261 12507
rect 4275 12455 4321 12507
rect 4321 12455 4327 12507
rect 4209 12386 4215 12438
rect 4215 12386 4261 12438
rect 4275 12386 4321 12438
rect 4321 12386 4327 12438
rect 4209 12316 4215 12368
rect 4215 12316 4261 12368
rect 4275 12316 4321 12368
rect 4321 12316 4327 12368
rect 4209 12246 4215 12298
rect 4215 12246 4261 12298
rect 4275 12246 4321 12298
rect 4321 12246 4327 12298
rect 4209 12176 4215 12228
rect 4215 12176 4261 12228
rect 4275 12176 4321 12228
rect 4321 12176 4327 12228
rect 4209 12112 4215 12158
rect 4215 12112 4261 12158
rect 4275 12112 4321 12158
rect 4321 12112 4327 12158
rect 4209 12106 4261 12112
rect 4275 12106 4327 12112
rect 4486 13446 4538 13452
rect 4486 13412 4492 13446
rect 4492 13412 4526 13446
rect 4526 13412 4538 13446
rect 4486 13400 4538 13412
rect 4552 13446 4604 13452
rect 4552 13412 4564 13446
rect 4564 13412 4598 13446
rect 4598 13412 4604 13446
rect 4552 13400 4604 13412
rect 4486 13373 4538 13383
rect 4486 13339 4492 13373
rect 4492 13339 4526 13373
rect 4526 13339 4538 13373
rect 4486 13331 4538 13339
rect 4552 13373 4604 13383
rect 4552 13339 4564 13373
rect 4564 13339 4598 13373
rect 4598 13339 4604 13373
rect 4552 13331 4604 13339
rect 4486 13300 4538 13314
rect 4486 13266 4492 13300
rect 4492 13266 4526 13300
rect 4526 13266 4538 13300
rect 4486 13262 4538 13266
rect 4552 13300 4604 13314
rect 4552 13266 4564 13300
rect 4564 13266 4598 13300
rect 4598 13266 4604 13300
rect 4552 13262 4604 13266
rect 4486 13227 4538 13245
rect 4486 13193 4492 13227
rect 4492 13193 4526 13227
rect 4526 13193 4538 13227
rect 4552 13227 4604 13245
rect 4552 13193 4564 13227
rect 4564 13193 4598 13227
rect 4598 13193 4604 13227
rect 4486 13154 4538 13176
rect 4552 13154 4604 13176
rect 4486 13124 4492 13154
rect 4492 13124 4538 13154
rect 4552 13124 4598 13154
rect 4598 13124 4604 13154
rect 4486 13055 4492 13107
rect 4492 13055 4538 13107
rect 4552 13055 4598 13107
rect 4598 13055 4604 13107
rect 4486 12986 4492 13038
rect 4492 12986 4538 13038
rect 4552 12986 4598 13038
rect 4598 12986 4604 13038
rect 4486 12916 4492 12968
rect 4492 12916 4538 12968
rect 4552 12916 4598 12968
rect 4598 12916 4604 12968
rect 4486 12846 4492 12898
rect 4492 12846 4538 12898
rect 4552 12846 4598 12898
rect 4598 12846 4604 12898
rect 4763 12662 4769 12714
rect 4769 12662 4815 12714
rect 4829 12662 4875 12714
rect 4875 12662 4881 12714
rect 4763 12593 4769 12645
rect 4769 12593 4815 12645
rect 4829 12593 4875 12645
rect 4875 12593 4881 12645
rect 4763 12524 4769 12576
rect 4769 12524 4815 12576
rect 4829 12524 4875 12576
rect 4875 12524 4881 12576
rect 4763 12455 4769 12507
rect 4769 12455 4815 12507
rect 4829 12455 4875 12507
rect 4875 12455 4881 12507
rect 4763 12386 4769 12438
rect 4769 12386 4815 12438
rect 4829 12386 4875 12438
rect 4875 12386 4881 12438
rect 4763 12316 4769 12368
rect 4769 12316 4815 12368
rect 4829 12316 4875 12368
rect 4875 12316 4881 12368
rect 4763 12246 4769 12298
rect 4769 12246 4815 12298
rect 4829 12246 4875 12298
rect 4875 12246 4881 12298
rect 4763 12176 4769 12228
rect 4769 12176 4815 12228
rect 4829 12176 4875 12228
rect 4875 12176 4881 12228
rect 4763 12112 4769 12158
rect 4769 12112 4815 12158
rect 4829 12112 4875 12158
rect 4875 12112 4881 12158
rect 4763 12106 4815 12112
rect 4829 12106 4881 12112
rect 5040 13446 5092 13452
rect 5040 13412 5046 13446
rect 5046 13412 5080 13446
rect 5080 13412 5092 13446
rect 5040 13400 5092 13412
rect 5106 13446 5158 13452
rect 5106 13412 5118 13446
rect 5118 13412 5152 13446
rect 5152 13412 5158 13446
rect 5106 13400 5158 13412
rect 5040 13373 5092 13383
rect 5040 13339 5046 13373
rect 5046 13339 5080 13373
rect 5080 13339 5092 13373
rect 5040 13331 5092 13339
rect 5106 13373 5158 13383
rect 5106 13339 5118 13373
rect 5118 13339 5152 13373
rect 5152 13339 5158 13373
rect 5106 13331 5158 13339
rect 5040 13300 5092 13314
rect 5040 13266 5046 13300
rect 5046 13266 5080 13300
rect 5080 13266 5092 13300
rect 5040 13262 5092 13266
rect 5106 13300 5158 13314
rect 5106 13266 5118 13300
rect 5118 13266 5152 13300
rect 5152 13266 5158 13300
rect 5106 13262 5158 13266
rect 5040 13227 5092 13245
rect 5040 13193 5046 13227
rect 5046 13193 5080 13227
rect 5080 13193 5092 13227
rect 5106 13227 5158 13245
rect 5106 13193 5118 13227
rect 5118 13193 5152 13227
rect 5152 13193 5158 13227
rect 5040 13154 5092 13176
rect 5106 13154 5158 13176
rect 5040 13124 5046 13154
rect 5046 13124 5092 13154
rect 5106 13124 5152 13154
rect 5152 13124 5158 13154
rect 5040 13055 5046 13107
rect 5046 13055 5092 13107
rect 5106 13055 5152 13107
rect 5152 13055 5158 13107
rect 5040 12986 5046 13038
rect 5046 12986 5092 13038
rect 5106 12986 5152 13038
rect 5152 12986 5158 13038
rect 5040 12916 5046 12968
rect 5046 12916 5092 12968
rect 5106 12916 5152 12968
rect 5152 12916 5158 12968
rect 5040 12846 5046 12898
rect 5046 12846 5092 12898
rect 5106 12846 5152 12898
rect 5152 12846 5158 12898
rect 5317 12662 5323 12714
rect 5323 12662 5369 12714
rect 5383 12662 5429 12714
rect 5429 12662 5435 12714
rect 5317 12593 5323 12645
rect 5323 12593 5369 12645
rect 5383 12593 5429 12645
rect 5429 12593 5435 12645
rect 5317 12524 5323 12576
rect 5323 12524 5369 12576
rect 5383 12524 5429 12576
rect 5429 12524 5435 12576
rect 5317 12455 5323 12507
rect 5323 12455 5369 12507
rect 5383 12455 5429 12507
rect 5429 12455 5435 12507
rect 5317 12386 5323 12438
rect 5323 12386 5369 12438
rect 5383 12386 5429 12438
rect 5429 12386 5435 12438
rect 5317 12316 5323 12368
rect 5323 12316 5369 12368
rect 5383 12316 5429 12368
rect 5429 12316 5435 12368
rect 5317 12246 5323 12298
rect 5323 12246 5369 12298
rect 5383 12246 5429 12298
rect 5429 12246 5435 12298
rect 5317 12176 5323 12228
rect 5323 12176 5369 12228
rect 5383 12176 5429 12228
rect 5429 12176 5435 12228
rect 5317 12112 5323 12158
rect 5323 12112 5369 12158
rect 5383 12112 5429 12158
rect 5429 12112 5435 12158
rect 5317 12106 5369 12112
rect 5383 12106 5435 12112
rect 5594 13446 5646 13452
rect 5594 13412 5600 13446
rect 5600 13412 5634 13446
rect 5634 13412 5646 13446
rect 5594 13400 5646 13412
rect 5660 13446 5712 13452
rect 5660 13412 5672 13446
rect 5672 13412 5706 13446
rect 5706 13412 5712 13446
rect 5660 13400 5712 13412
rect 5594 13373 5646 13383
rect 5594 13339 5600 13373
rect 5600 13339 5634 13373
rect 5634 13339 5646 13373
rect 5594 13331 5646 13339
rect 5660 13373 5712 13383
rect 5660 13339 5672 13373
rect 5672 13339 5706 13373
rect 5706 13339 5712 13373
rect 5660 13331 5712 13339
rect 5594 13300 5646 13314
rect 5594 13266 5600 13300
rect 5600 13266 5634 13300
rect 5634 13266 5646 13300
rect 5594 13262 5646 13266
rect 5660 13300 5712 13314
rect 5660 13266 5672 13300
rect 5672 13266 5706 13300
rect 5706 13266 5712 13300
rect 5660 13262 5712 13266
rect 5594 13227 5646 13245
rect 5594 13193 5600 13227
rect 5600 13193 5634 13227
rect 5634 13193 5646 13227
rect 5660 13227 5712 13245
rect 5660 13193 5672 13227
rect 5672 13193 5706 13227
rect 5706 13193 5712 13227
rect 5594 13154 5646 13176
rect 5660 13154 5712 13176
rect 5594 13124 5600 13154
rect 5600 13124 5646 13154
rect 5660 13124 5706 13154
rect 5706 13124 5712 13154
rect 5594 13055 5600 13107
rect 5600 13055 5646 13107
rect 5660 13055 5706 13107
rect 5706 13055 5712 13107
rect 5594 12986 5600 13038
rect 5600 12986 5646 13038
rect 5660 12986 5706 13038
rect 5706 12986 5712 13038
rect 5594 12916 5600 12968
rect 5600 12916 5646 12968
rect 5660 12916 5706 12968
rect 5706 12916 5712 12968
rect 5594 12846 5600 12898
rect 5600 12846 5646 12898
rect 5660 12846 5706 12898
rect 5706 12846 5712 12898
rect 5871 12662 5877 12714
rect 5877 12662 5923 12714
rect 5937 12662 5983 12714
rect 5983 12662 5989 12714
rect 5871 12593 5877 12645
rect 5877 12593 5923 12645
rect 5937 12593 5983 12645
rect 5983 12593 5989 12645
rect 5871 12524 5877 12576
rect 5877 12524 5923 12576
rect 5937 12524 5983 12576
rect 5983 12524 5989 12576
rect 5871 12455 5877 12507
rect 5877 12455 5923 12507
rect 5937 12455 5983 12507
rect 5983 12455 5989 12507
rect 5871 12386 5877 12438
rect 5877 12386 5923 12438
rect 5937 12386 5983 12438
rect 5983 12386 5989 12438
rect 5871 12316 5877 12368
rect 5877 12316 5923 12368
rect 5937 12316 5983 12368
rect 5983 12316 5989 12368
rect 5871 12246 5877 12298
rect 5877 12246 5923 12298
rect 5937 12246 5983 12298
rect 5983 12246 5989 12298
rect 5871 12176 5877 12228
rect 5877 12176 5923 12228
rect 5937 12176 5983 12228
rect 5983 12176 5989 12228
rect 5871 12112 5877 12158
rect 5877 12112 5923 12158
rect 5937 12112 5983 12158
rect 5983 12112 5989 12158
rect 5871 12106 5923 12112
rect 5937 12106 5989 12112
rect 6148 13446 6200 13452
rect 6148 13412 6154 13446
rect 6154 13412 6188 13446
rect 6188 13412 6200 13446
rect 6148 13400 6200 13412
rect 6214 13446 6266 13452
rect 6214 13412 6226 13446
rect 6226 13412 6260 13446
rect 6260 13412 6266 13446
rect 6214 13400 6266 13412
rect 6148 13373 6200 13383
rect 6148 13339 6154 13373
rect 6154 13339 6188 13373
rect 6188 13339 6200 13373
rect 6148 13331 6200 13339
rect 6214 13373 6266 13383
rect 6214 13339 6226 13373
rect 6226 13339 6260 13373
rect 6260 13339 6266 13373
rect 6214 13331 6266 13339
rect 6148 13300 6200 13314
rect 6148 13266 6154 13300
rect 6154 13266 6188 13300
rect 6188 13266 6200 13300
rect 6148 13262 6200 13266
rect 6214 13300 6266 13314
rect 6214 13266 6226 13300
rect 6226 13266 6260 13300
rect 6260 13266 6266 13300
rect 6214 13262 6266 13266
rect 6148 13227 6200 13245
rect 6148 13193 6154 13227
rect 6154 13193 6188 13227
rect 6188 13193 6200 13227
rect 6214 13227 6266 13245
rect 6214 13193 6226 13227
rect 6226 13193 6260 13227
rect 6260 13193 6266 13227
rect 6148 13154 6200 13176
rect 6214 13154 6266 13176
rect 6148 13124 6154 13154
rect 6154 13124 6200 13154
rect 6214 13124 6260 13154
rect 6260 13124 6266 13154
rect 6148 13055 6154 13107
rect 6154 13055 6200 13107
rect 6214 13055 6260 13107
rect 6260 13055 6266 13107
rect 6148 12986 6154 13038
rect 6154 12986 6200 13038
rect 6214 12986 6260 13038
rect 6260 12986 6266 13038
rect 6148 12916 6154 12968
rect 6154 12916 6200 12968
rect 6214 12916 6260 12968
rect 6260 12916 6266 12968
rect 6148 12846 6154 12898
rect 6154 12846 6200 12898
rect 6214 12846 6260 12898
rect 6260 12846 6266 12898
rect 6425 12662 6431 12714
rect 6431 12662 6477 12714
rect 6491 12662 6537 12714
rect 6537 12662 6543 12714
rect 6425 12593 6431 12645
rect 6431 12593 6477 12645
rect 6491 12593 6537 12645
rect 6537 12593 6543 12645
rect 6425 12524 6431 12576
rect 6431 12524 6477 12576
rect 6491 12524 6537 12576
rect 6537 12524 6543 12576
rect 6425 12455 6431 12507
rect 6431 12455 6477 12507
rect 6491 12455 6537 12507
rect 6537 12455 6543 12507
rect 6425 12386 6431 12438
rect 6431 12386 6477 12438
rect 6491 12386 6537 12438
rect 6537 12386 6543 12438
rect 6425 12316 6431 12368
rect 6431 12316 6477 12368
rect 6491 12316 6537 12368
rect 6537 12316 6543 12368
rect 6425 12246 6431 12298
rect 6431 12246 6477 12298
rect 6491 12246 6537 12298
rect 6537 12246 6543 12298
rect 6425 12176 6431 12228
rect 6431 12176 6477 12228
rect 6491 12176 6537 12228
rect 6537 12176 6543 12228
rect 6425 12112 6431 12158
rect 6431 12112 6477 12158
rect 6491 12112 6537 12158
rect 6537 12112 6543 12158
rect 6425 12106 6477 12112
rect 6491 12106 6543 12112
rect 6702 13446 6754 13452
rect 6702 13412 6708 13446
rect 6708 13412 6742 13446
rect 6742 13412 6754 13446
rect 6702 13400 6754 13412
rect 6768 13446 6820 13452
rect 6768 13412 6780 13446
rect 6780 13412 6814 13446
rect 6814 13412 6820 13446
rect 6768 13400 6820 13412
rect 6702 13373 6754 13383
rect 6702 13339 6708 13373
rect 6708 13339 6742 13373
rect 6742 13339 6754 13373
rect 6702 13331 6754 13339
rect 6768 13373 6820 13383
rect 6768 13339 6780 13373
rect 6780 13339 6814 13373
rect 6814 13339 6820 13373
rect 6768 13331 6820 13339
rect 6702 13300 6754 13314
rect 6702 13266 6708 13300
rect 6708 13266 6742 13300
rect 6742 13266 6754 13300
rect 6702 13262 6754 13266
rect 6768 13300 6820 13314
rect 6768 13266 6780 13300
rect 6780 13266 6814 13300
rect 6814 13266 6820 13300
rect 6768 13262 6820 13266
rect 6702 13227 6754 13245
rect 6702 13193 6708 13227
rect 6708 13193 6742 13227
rect 6742 13193 6754 13227
rect 6768 13227 6820 13245
rect 6768 13193 6780 13227
rect 6780 13193 6814 13227
rect 6814 13193 6820 13227
rect 6702 13154 6754 13176
rect 6768 13154 6820 13176
rect 6702 13124 6708 13154
rect 6708 13124 6754 13154
rect 6768 13124 6814 13154
rect 6814 13124 6820 13154
rect 6702 13055 6708 13107
rect 6708 13055 6754 13107
rect 6768 13055 6814 13107
rect 6814 13055 6820 13107
rect 6702 12986 6708 13038
rect 6708 12986 6754 13038
rect 6768 12986 6814 13038
rect 6814 12986 6820 13038
rect 6702 12916 6708 12968
rect 6708 12916 6754 12968
rect 6768 12916 6814 12968
rect 6814 12916 6820 12968
rect 6702 12846 6708 12898
rect 6708 12846 6754 12898
rect 6768 12846 6814 12898
rect 6814 12846 6820 12898
rect 6979 12662 6985 12714
rect 6985 12662 7031 12714
rect 7045 12662 7091 12714
rect 7091 12662 7097 12714
rect 6979 12593 6985 12645
rect 6985 12593 7031 12645
rect 7045 12593 7091 12645
rect 7091 12593 7097 12645
rect 6979 12524 6985 12576
rect 6985 12524 7031 12576
rect 7045 12524 7091 12576
rect 7091 12524 7097 12576
rect 6979 12455 6985 12507
rect 6985 12455 7031 12507
rect 7045 12455 7091 12507
rect 7091 12455 7097 12507
rect 6979 12386 6985 12438
rect 6985 12386 7031 12438
rect 7045 12386 7091 12438
rect 7091 12386 7097 12438
rect 6979 12316 6985 12368
rect 6985 12316 7031 12368
rect 7045 12316 7091 12368
rect 7091 12316 7097 12368
rect 6979 12246 6985 12298
rect 6985 12246 7031 12298
rect 7045 12246 7091 12298
rect 7091 12246 7097 12298
rect 6979 12176 6985 12228
rect 6985 12176 7031 12228
rect 7045 12176 7091 12228
rect 7091 12176 7097 12228
rect 6979 12112 6985 12158
rect 6985 12112 7031 12158
rect 7045 12112 7091 12158
rect 7091 12112 7097 12158
rect 6979 12106 7031 12112
rect 7045 12106 7097 12112
rect 7256 13446 7308 13452
rect 7256 13412 7262 13446
rect 7262 13412 7296 13446
rect 7296 13412 7308 13446
rect 7256 13400 7308 13412
rect 7322 13446 7374 13452
rect 7322 13412 7334 13446
rect 7334 13412 7368 13446
rect 7368 13412 7374 13446
rect 7322 13400 7374 13412
rect 7256 13373 7308 13383
rect 7256 13339 7262 13373
rect 7262 13339 7296 13373
rect 7296 13339 7308 13373
rect 7256 13331 7308 13339
rect 7322 13373 7374 13383
rect 7322 13339 7334 13373
rect 7334 13339 7368 13373
rect 7368 13339 7374 13373
rect 7322 13331 7374 13339
rect 7256 13300 7308 13314
rect 7256 13266 7262 13300
rect 7262 13266 7296 13300
rect 7296 13266 7308 13300
rect 7256 13262 7308 13266
rect 7322 13300 7374 13314
rect 7322 13266 7334 13300
rect 7334 13266 7368 13300
rect 7368 13266 7374 13300
rect 7322 13262 7374 13266
rect 7256 13227 7308 13245
rect 7256 13193 7262 13227
rect 7262 13193 7296 13227
rect 7296 13193 7308 13227
rect 7322 13227 7374 13245
rect 7322 13193 7334 13227
rect 7334 13193 7368 13227
rect 7368 13193 7374 13227
rect 7256 13154 7308 13176
rect 7322 13154 7374 13176
rect 7256 13124 7262 13154
rect 7262 13124 7308 13154
rect 7322 13124 7368 13154
rect 7368 13124 7374 13154
rect 7256 13055 7262 13107
rect 7262 13055 7308 13107
rect 7322 13055 7368 13107
rect 7368 13055 7374 13107
rect 7256 12986 7262 13038
rect 7262 12986 7308 13038
rect 7322 12986 7368 13038
rect 7368 12986 7374 13038
rect 7256 12916 7262 12968
rect 7262 12916 7308 12968
rect 7322 12916 7368 12968
rect 7368 12916 7374 12968
rect 7256 12846 7262 12898
rect 7262 12846 7308 12898
rect 7322 12846 7368 12898
rect 7368 12846 7374 12898
rect 7533 12662 7539 12714
rect 7539 12662 7585 12714
rect 7599 12662 7645 12714
rect 7645 12662 7651 12714
rect 7533 12593 7539 12645
rect 7539 12593 7585 12645
rect 7599 12593 7645 12645
rect 7645 12593 7651 12645
rect 7533 12524 7539 12576
rect 7539 12524 7585 12576
rect 7599 12524 7645 12576
rect 7645 12524 7651 12576
rect 7533 12455 7539 12507
rect 7539 12455 7585 12507
rect 7599 12455 7645 12507
rect 7645 12455 7651 12507
rect 7533 12386 7539 12438
rect 7539 12386 7585 12438
rect 7599 12386 7645 12438
rect 7645 12386 7651 12438
rect 7533 12316 7539 12368
rect 7539 12316 7585 12368
rect 7599 12316 7645 12368
rect 7645 12316 7651 12368
rect 7533 12246 7539 12298
rect 7539 12246 7585 12298
rect 7599 12246 7645 12298
rect 7645 12246 7651 12298
rect 7533 12176 7539 12228
rect 7539 12176 7585 12228
rect 7599 12176 7645 12228
rect 7645 12176 7651 12228
rect 7533 12112 7539 12158
rect 7539 12112 7585 12158
rect 7599 12112 7645 12158
rect 7645 12112 7651 12158
rect 7533 12106 7585 12112
rect 7599 12106 7651 12112
rect 7810 13446 7862 13452
rect 7810 13412 7816 13446
rect 7816 13412 7850 13446
rect 7850 13412 7862 13446
rect 7810 13400 7862 13412
rect 7876 13446 7928 13452
rect 7876 13412 7888 13446
rect 7888 13412 7922 13446
rect 7922 13412 7928 13446
rect 7876 13400 7928 13412
rect 7810 13373 7862 13383
rect 7810 13339 7816 13373
rect 7816 13339 7850 13373
rect 7850 13339 7862 13373
rect 7810 13331 7862 13339
rect 7876 13373 7928 13383
rect 7876 13339 7888 13373
rect 7888 13339 7922 13373
rect 7922 13339 7928 13373
rect 7876 13331 7928 13339
rect 7810 13300 7862 13314
rect 7810 13266 7816 13300
rect 7816 13266 7850 13300
rect 7850 13266 7862 13300
rect 7810 13262 7862 13266
rect 7876 13300 7928 13314
rect 7876 13266 7888 13300
rect 7888 13266 7922 13300
rect 7922 13266 7928 13300
rect 7876 13262 7928 13266
rect 7810 13227 7862 13245
rect 7810 13193 7816 13227
rect 7816 13193 7850 13227
rect 7850 13193 7862 13227
rect 7876 13227 7928 13245
rect 7876 13193 7888 13227
rect 7888 13193 7922 13227
rect 7922 13193 7928 13227
rect 7810 13154 7862 13176
rect 7876 13154 7928 13176
rect 7810 13124 7816 13154
rect 7816 13124 7862 13154
rect 7876 13124 7922 13154
rect 7922 13124 7928 13154
rect 7810 13055 7816 13107
rect 7816 13055 7862 13107
rect 7876 13055 7922 13107
rect 7922 13055 7928 13107
rect 7810 12986 7816 13038
rect 7816 12986 7862 13038
rect 7876 12986 7922 13038
rect 7922 12986 7928 13038
rect 7810 12916 7816 12968
rect 7816 12916 7862 12968
rect 7876 12916 7922 12968
rect 7922 12916 7928 12968
rect 7810 12846 7816 12898
rect 7816 12846 7862 12898
rect 7876 12846 7922 12898
rect 7922 12846 7928 12898
rect 8047 13447 8099 13456
rect 8047 13413 8050 13447
rect 8050 13413 8084 13447
rect 8084 13413 8099 13447
rect 8047 13404 8099 13413
rect 8169 13437 8221 13456
rect 8169 13404 8184 13437
rect 8184 13404 8218 13437
rect 8218 13404 8221 13437
rect 8047 13375 8099 13387
rect 8047 13341 8050 13375
rect 8050 13341 8084 13375
rect 8084 13341 8099 13375
rect 8047 13335 8099 13341
rect 8169 13365 8221 13387
rect 8169 13335 8184 13365
rect 8184 13335 8218 13365
rect 8218 13335 8221 13365
rect 8047 13303 8099 13318
rect 8047 13269 8050 13303
rect 8050 13269 8084 13303
rect 8084 13269 8099 13303
rect 8047 13266 8099 13269
rect 8169 13293 8221 13318
rect 8169 13266 8184 13293
rect 8184 13266 8218 13293
rect 8218 13266 8221 13293
rect 8047 13231 8099 13249
rect 8047 13197 8050 13231
rect 8050 13197 8084 13231
rect 8084 13197 8099 13231
rect 8169 13221 8221 13249
rect 8169 13197 8184 13221
rect 8184 13197 8218 13221
rect 8218 13197 8221 13221
rect 8047 13159 8099 13180
rect 8047 13128 8050 13159
rect 8050 13128 8084 13159
rect 8084 13128 8099 13159
rect 8169 13149 8221 13180
rect 8169 13128 8184 13149
rect 8184 13128 8218 13149
rect 8218 13128 8221 13149
rect 8047 13087 8099 13110
rect 8047 13058 8050 13087
rect 8050 13058 8084 13087
rect 8084 13058 8099 13087
rect 8169 13077 8221 13110
rect 8169 13058 8184 13077
rect 8184 13058 8218 13077
rect 8218 13058 8221 13077
rect 8047 13015 8099 13040
rect 8047 12988 8050 13015
rect 8050 12988 8084 13015
rect 8084 12988 8099 13015
rect 8169 13005 8221 13040
rect 8169 12988 8184 13005
rect 8184 12988 8218 13005
rect 8218 12988 8221 13005
rect 8047 12942 8099 12970
rect 8047 12918 8050 12942
rect 8050 12918 8084 12942
rect 8084 12918 8099 12942
rect 8169 12933 8221 12970
rect 8169 12918 8184 12933
rect 8184 12918 8218 12933
rect 8218 12918 8221 12933
rect 8047 12869 8099 12900
rect 8047 12848 8050 12869
rect 8050 12848 8084 12869
rect 8084 12848 8099 12869
rect 8169 12899 8184 12900
rect 8184 12899 8218 12900
rect 8218 12899 8221 12900
rect 8169 12861 8221 12899
rect 8169 12848 8184 12861
rect 8184 12848 8218 12861
rect 8218 12848 8221 12861
rect 2580 10470 2632 10522
rect 2660 10470 2712 10522
rect 2580 10404 2632 10456
rect 2660 10404 2712 10456
rect 2580 10338 2632 10390
rect 2660 10338 2712 10390
rect 2580 10272 2632 10324
rect 2660 10272 2712 10324
rect 2580 10206 2632 10258
rect 2660 10206 2712 10258
rect 2580 10140 2632 10192
rect 2660 10140 2712 10192
rect 2580 10074 2632 10126
rect 2660 10074 2712 10126
rect 2824 11446 2876 11452
rect 2824 11412 2830 11446
rect 2830 11412 2864 11446
rect 2864 11412 2876 11446
rect 2824 11400 2876 11412
rect 2890 11446 2942 11452
rect 2890 11412 2902 11446
rect 2902 11412 2936 11446
rect 2936 11412 2942 11446
rect 2890 11400 2942 11412
rect 2824 11373 2876 11383
rect 2824 11339 2830 11373
rect 2830 11339 2864 11373
rect 2864 11339 2876 11373
rect 2824 11331 2876 11339
rect 2890 11373 2942 11383
rect 2890 11339 2902 11373
rect 2902 11339 2936 11373
rect 2936 11339 2942 11373
rect 2890 11331 2942 11339
rect 2824 11300 2876 11314
rect 2824 11266 2830 11300
rect 2830 11266 2864 11300
rect 2864 11266 2876 11300
rect 2824 11262 2876 11266
rect 2890 11300 2942 11314
rect 2890 11266 2902 11300
rect 2902 11266 2936 11300
rect 2936 11266 2942 11300
rect 2890 11262 2942 11266
rect 2824 11227 2876 11245
rect 2824 11193 2830 11227
rect 2830 11193 2864 11227
rect 2864 11193 2876 11227
rect 2890 11227 2942 11245
rect 2890 11193 2902 11227
rect 2902 11193 2936 11227
rect 2936 11193 2942 11227
rect 2824 11154 2876 11176
rect 2890 11154 2942 11176
rect 2824 11124 2830 11154
rect 2830 11124 2876 11154
rect 2890 11124 2936 11154
rect 2936 11124 2942 11154
rect 2824 11055 2830 11107
rect 2830 11055 2876 11107
rect 2890 11055 2936 11107
rect 2936 11055 2942 11107
rect 2824 10986 2830 11038
rect 2830 10986 2876 11038
rect 2890 10986 2936 11038
rect 2936 10986 2942 11038
rect 2824 10916 2830 10968
rect 2830 10916 2876 10968
rect 2890 10916 2936 10968
rect 2936 10916 2942 10968
rect 2824 10846 2830 10898
rect 2830 10846 2876 10898
rect 2890 10846 2936 10898
rect 2936 10846 2942 10898
rect 3101 10662 3107 10714
rect 3107 10662 3153 10714
rect 3167 10662 3213 10714
rect 3213 10662 3219 10714
rect 3101 10593 3107 10645
rect 3107 10593 3153 10645
rect 3167 10593 3213 10645
rect 3213 10593 3219 10645
rect 3101 10524 3107 10576
rect 3107 10524 3153 10576
rect 3167 10524 3213 10576
rect 3213 10524 3219 10576
rect 3101 10455 3107 10507
rect 3107 10455 3153 10507
rect 3167 10455 3213 10507
rect 3213 10455 3219 10507
rect 3101 10386 3107 10438
rect 3107 10386 3153 10438
rect 3167 10386 3213 10438
rect 3213 10386 3219 10438
rect 3101 10316 3107 10368
rect 3107 10316 3153 10368
rect 3167 10316 3213 10368
rect 3213 10316 3219 10368
rect 3101 10246 3107 10298
rect 3107 10246 3153 10298
rect 3167 10246 3213 10298
rect 3213 10246 3219 10298
rect 3101 10176 3107 10228
rect 3107 10176 3153 10228
rect 3167 10176 3213 10228
rect 3213 10176 3219 10228
rect 3101 10112 3107 10158
rect 3107 10112 3153 10158
rect 3167 10112 3213 10158
rect 3213 10112 3219 10158
rect 3101 10106 3153 10112
rect 3167 10106 3219 10112
rect 3378 11446 3430 11452
rect 3378 11412 3384 11446
rect 3384 11412 3418 11446
rect 3418 11412 3430 11446
rect 3378 11400 3430 11412
rect 3444 11446 3496 11452
rect 3444 11412 3456 11446
rect 3456 11412 3490 11446
rect 3490 11412 3496 11446
rect 3444 11400 3496 11412
rect 3378 11373 3430 11383
rect 3378 11339 3384 11373
rect 3384 11339 3418 11373
rect 3418 11339 3430 11373
rect 3378 11331 3430 11339
rect 3444 11373 3496 11383
rect 3444 11339 3456 11373
rect 3456 11339 3490 11373
rect 3490 11339 3496 11373
rect 3444 11331 3496 11339
rect 3378 11300 3430 11314
rect 3378 11266 3384 11300
rect 3384 11266 3418 11300
rect 3418 11266 3430 11300
rect 3378 11262 3430 11266
rect 3444 11300 3496 11314
rect 3444 11266 3456 11300
rect 3456 11266 3490 11300
rect 3490 11266 3496 11300
rect 3444 11262 3496 11266
rect 3378 11227 3430 11245
rect 3378 11193 3384 11227
rect 3384 11193 3418 11227
rect 3418 11193 3430 11227
rect 3444 11227 3496 11245
rect 3444 11193 3456 11227
rect 3456 11193 3490 11227
rect 3490 11193 3496 11227
rect 3378 11154 3430 11176
rect 3444 11154 3496 11176
rect 3378 11124 3384 11154
rect 3384 11124 3430 11154
rect 3444 11124 3490 11154
rect 3490 11124 3496 11154
rect 3378 11055 3384 11107
rect 3384 11055 3430 11107
rect 3444 11055 3490 11107
rect 3490 11055 3496 11107
rect 3378 10986 3384 11038
rect 3384 10986 3430 11038
rect 3444 10986 3490 11038
rect 3490 10986 3496 11038
rect 3378 10916 3384 10968
rect 3384 10916 3430 10968
rect 3444 10916 3490 10968
rect 3490 10916 3496 10968
rect 3378 10846 3384 10898
rect 3384 10846 3430 10898
rect 3444 10846 3490 10898
rect 3490 10846 3496 10898
rect 3655 10662 3661 10714
rect 3661 10662 3707 10714
rect 3721 10662 3767 10714
rect 3767 10662 3773 10714
rect 3655 10593 3661 10645
rect 3661 10593 3707 10645
rect 3721 10593 3767 10645
rect 3767 10593 3773 10645
rect 3655 10524 3661 10576
rect 3661 10524 3707 10576
rect 3721 10524 3767 10576
rect 3767 10524 3773 10576
rect 3655 10455 3661 10507
rect 3661 10455 3707 10507
rect 3721 10455 3767 10507
rect 3767 10455 3773 10507
rect 3655 10386 3661 10438
rect 3661 10386 3707 10438
rect 3721 10386 3767 10438
rect 3767 10386 3773 10438
rect 3655 10316 3661 10368
rect 3661 10316 3707 10368
rect 3721 10316 3767 10368
rect 3767 10316 3773 10368
rect 3655 10246 3661 10298
rect 3661 10246 3707 10298
rect 3721 10246 3767 10298
rect 3767 10246 3773 10298
rect 3655 10176 3661 10228
rect 3661 10176 3707 10228
rect 3721 10176 3767 10228
rect 3767 10176 3773 10228
rect 3655 10112 3661 10158
rect 3661 10112 3707 10158
rect 3721 10112 3767 10158
rect 3767 10112 3773 10158
rect 3655 10106 3707 10112
rect 3721 10106 3773 10112
rect 3932 11446 3984 11452
rect 3932 11412 3938 11446
rect 3938 11412 3972 11446
rect 3972 11412 3984 11446
rect 3932 11400 3984 11412
rect 3998 11446 4050 11452
rect 3998 11412 4010 11446
rect 4010 11412 4044 11446
rect 4044 11412 4050 11446
rect 3998 11400 4050 11412
rect 3932 11373 3984 11383
rect 3932 11339 3938 11373
rect 3938 11339 3972 11373
rect 3972 11339 3984 11373
rect 3932 11331 3984 11339
rect 3998 11373 4050 11383
rect 3998 11339 4010 11373
rect 4010 11339 4044 11373
rect 4044 11339 4050 11373
rect 3998 11331 4050 11339
rect 3932 11300 3984 11314
rect 3932 11266 3938 11300
rect 3938 11266 3972 11300
rect 3972 11266 3984 11300
rect 3932 11262 3984 11266
rect 3998 11300 4050 11314
rect 3998 11266 4010 11300
rect 4010 11266 4044 11300
rect 4044 11266 4050 11300
rect 3998 11262 4050 11266
rect 3932 11227 3984 11245
rect 3932 11193 3938 11227
rect 3938 11193 3972 11227
rect 3972 11193 3984 11227
rect 3998 11227 4050 11245
rect 3998 11193 4010 11227
rect 4010 11193 4044 11227
rect 4044 11193 4050 11227
rect 3932 11154 3984 11176
rect 3998 11154 4050 11176
rect 3932 11124 3938 11154
rect 3938 11124 3984 11154
rect 3998 11124 4044 11154
rect 4044 11124 4050 11154
rect 3932 11055 3938 11107
rect 3938 11055 3984 11107
rect 3998 11055 4044 11107
rect 4044 11055 4050 11107
rect 3932 10986 3938 11038
rect 3938 10986 3984 11038
rect 3998 10986 4044 11038
rect 4044 10986 4050 11038
rect 3932 10916 3938 10968
rect 3938 10916 3984 10968
rect 3998 10916 4044 10968
rect 4044 10916 4050 10968
rect 3932 10846 3938 10898
rect 3938 10846 3984 10898
rect 3998 10846 4044 10898
rect 4044 10846 4050 10898
rect 4209 10662 4215 10714
rect 4215 10662 4261 10714
rect 4275 10662 4321 10714
rect 4321 10662 4327 10714
rect 4209 10593 4215 10645
rect 4215 10593 4261 10645
rect 4275 10593 4321 10645
rect 4321 10593 4327 10645
rect 4209 10524 4215 10576
rect 4215 10524 4261 10576
rect 4275 10524 4321 10576
rect 4321 10524 4327 10576
rect 4209 10455 4215 10507
rect 4215 10455 4261 10507
rect 4275 10455 4321 10507
rect 4321 10455 4327 10507
rect 4209 10386 4215 10438
rect 4215 10386 4261 10438
rect 4275 10386 4321 10438
rect 4321 10386 4327 10438
rect 4209 10316 4215 10368
rect 4215 10316 4261 10368
rect 4275 10316 4321 10368
rect 4321 10316 4327 10368
rect 4209 10246 4215 10298
rect 4215 10246 4261 10298
rect 4275 10246 4321 10298
rect 4321 10246 4327 10298
rect 4209 10176 4215 10228
rect 4215 10176 4261 10228
rect 4275 10176 4321 10228
rect 4321 10176 4327 10228
rect 4209 10112 4215 10158
rect 4215 10112 4261 10158
rect 4275 10112 4321 10158
rect 4321 10112 4327 10158
rect 4209 10106 4261 10112
rect 4275 10106 4327 10112
rect 4486 11446 4538 11452
rect 4486 11412 4492 11446
rect 4492 11412 4526 11446
rect 4526 11412 4538 11446
rect 4486 11400 4538 11412
rect 4552 11446 4604 11452
rect 4552 11412 4564 11446
rect 4564 11412 4598 11446
rect 4598 11412 4604 11446
rect 4552 11400 4604 11412
rect 4486 11373 4538 11383
rect 4486 11339 4492 11373
rect 4492 11339 4526 11373
rect 4526 11339 4538 11373
rect 4486 11331 4538 11339
rect 4552 11373 4604 11383
rect 4552 11339 4564 11373
rect 4564 11339 4598 11373
rect 4598 11339 4604 11373
rect 4552 11331 4604 11339
rect 4486 11300 4538 11314
rect 4486 11266 4492 11300
rect 4492 11266 4526 11300
rect 4526 11266 4538 11300
rect 4486 11262 4538 11266
rect 4552 11300 4604 11314
rect 4552 11266 4564 11300
rect 4564 11266 4598 11300
rect 4598 11266 4604 11300
rect 4552 11262 4604 11266
rect 4486 11227 4538 11245
rect 4486 11193 4492 11227
rect 4492 11193 4526 11227
rect 4526 11193 4538 11227
rect 4552 11227 4604 11245
rect 4552 11193 4564 11227
rect 4564 11193 4598 11227
rect 4598 11193 4604 11227
rect 4486 11154 4538 11176
rect 4552 11154 4604 11176
rect 4486 11124 4492 11154
rect 4492 11124 4538 11154
rect 4552 11124 4598 11154
rect 4598 11124 4604 11154
rect 4486 11055 4492 11107
rect 4492 11055 4538 11107
rect 4552 11055 4598 11107
rect 4598 11055 4604 11107
rect 4486 10986 4492 11038
rect 4492 10986 4538 11038
rect 4552 10986 4598 11038
rect 4598 10986 4604 11038
rect 4486 10916 4492 10968
rect 4492 10916 4538 10968
rect 4552 10916 4598 10968
rect 4598 10916 4604 10968
rect 4486 10846 4492 10898
rect 4492 10846 4538 10898
rect 4552 10846 4598 10898
rect 4598 10846 4604 10898
rect 4763 10662 4769 10714
rect 4769 10662 4815 10714
rect 4829 10662 4875 10714
rect 4875 10662 4881 10714
rect 4763 10593 4769 10645
rect 4769 10593 4815 10645
rect 4829 10593 4875 10645
rect 4875 10593 4881 10645
rect 4763 10524 4769 10576
rect 4769 10524 4815 10576
rect 4829 10524 4875 10576
rect 4875 10524 4881 10576
rect 4763 10455 4769 10507
rect 4769 10455 4815 10507
rect 4829 10455 4875 10507
rect 4875 10455 4881 10507
rect 4763 10386 4769 10438
rect 4769 10386 4815 10438
rect 4829 10386 4875 10438
rect 4875 10386 4881 10438
rect 4763 10316 4769 10368
rect 4769 10316 4815 10368
rect 4829 10316 4875 10368
rect 4875 10316 4881 10368
rect 4763 10246 4769 10298
rect 4769 10246 4815 10298
rect 4829 10246 4875 10298
rect 4875 10246 4881 10298
rect 4763 10176 4769 10228
rect 4769 10176 4815 10228
rect 4829 10176 4875 10228
rect 4875 10176 4881 10228
rect 4763 10112 4769 10158
rect 4769 10112 4815 10158
rect 4829 10112 4875 10158
rect 4875 10112 4881 10158
rect 4763 10106 4815 10112
rect 4829 10106 4881 10112
rect 5040 11446 5092 11452
rect 5040 11412 5046 11446
rect 5046 11412 5080 11446
rect 5080 11412 5092 11446
rect 5040 11400 5092 11412
rect 5106 11446 5158 11452
rect 5106 11412 5118 11446
rect 5118 11412 5152 11446
rect 5152 11412 5158 11446
rect 5106 11400 5158 11412
rect 5040 11373 5092 11383
rect 5040 11339 5046 11373
rect 5046 11339 5080 11373
rect 5080 11339 5092 11373
rect 5040 11331 5092 11339
rect 5106 11373 5158 11383
rect 5106 11339 5118 11373
rect 5118 11339 5152 11373
rect 5152 11339 5158 11373
rect 5106 11331 5158 11339
rect 5040 11300 5092 11314
rect 5040 11266 5046 11300
rect 5046 11266 5080 11300
rect 5080 11266 5092 11300
rect 5040 11262 5092 11266
rect 5106 11300 5158 11314
rect 5106 11266 5118 11300
rect 5118 11266 5152 11300
rect 5152 11266 5158 11300
rect 5106 11262 5158 11266
rect 5040 11227 5092 11245
rect 5040 11193 5046 11227
rect 5046 11193 5080 11227
rect 5080 11193 5092 11227
rect 5106 11227 5158 11245
rect 5106 11193 5118 11227
rect 5118 11193 5152 11227
rect 5152 11193 5158 11227
rect 5040 11154 5092 11176
rect 5106 11154 5158 11176
rect 5040 11124 5046 11154
rect 5046 11124 5092 11154
rect 5106 11124 5152 11154
rect 5152 11124 5158 11154
rect 5040 11055 5046 11107
rect 5046 11055 5092 11107
rect 5106 11055 5152 11107
rect 5152 11055 5158 11107
rect 5040 10986 5046 11038
rect 5046 10986 5092 11038
rect 5106 10986 5152 11038
rect 5152 10986 5158 11038
rect 5040 10916 5046 10968
rect 5046 10916 5092 10968
rect 5106 10916 5152 10968
rect 5152 10916 5158 10968
rect 5040 10846 5046 10898
rect 5046 10846 5092 10898
rect 5106 10846 5152 10898
rect 5152 10846 5158 10898
rect 5317 10662 5323 10714
rect 5323 10662 5369 10714
rect 5383 10662 5429 10714
rect 5429 10662 5435 10714
rect 5317 10593 5323 10645
rect 5323 10593 5369 10645
rect 5383 10593 5429 10645
rect 5429 10593 5435 10645
rect 5317 10524 5323 10576
rect 5323 10524 5369 10576
rect 5383 10524 5429 10576
rect 5429 10524 5435 10576
rect 5317 10455 5323 10507
rect 5323 10455 5369 10507
rect 5383 10455 5429 10507
rect 5429 10455 5435 10507
rect 5317 10386 5323 10438
rect 5323 10386 5369 10438
rect 5383 10386 5429 10438
rect 5429 10386 5435 10438
rect 5317 10316 5323 10368
rect 5323 10316 5369 10368
rect 5383 10316 5429 10368
rect 5429 10316 5435 10368
rect 5317 10246 5323 10298
rect 5323 10246 5369 10298
rect 5383 10246 5429 10298
rect 5429 10246 5435 10298
rect 5317 10176 5323 10228
rect 5323 10176 5369 10228
rect 5383 10176 5429 10228
rect 5429 10176 5435 10228
rect 5317 10112 5323 10158
rect 5323 10112 5369 10158
rect 5383 10112 5429 10158
rect 5429 10112 5435 10158
rect 5317 10106 5369 10112
rect 5383 10106 5435 10112
rect 5594 11446 5646 11452
rect 5594 11412 5600 11446
rect 5600 11412 5634 11446
rect 5634 11412 5646 11446
rect 5594 11400 5646 11412
rect 5660 11446 5712 11452
rect 5660 11412 5672 11446
rect 5672 11412 5706 11446
rect 5706 11412 5712 11446
rect 5660 11400 5712 11412
rect 5594 11373 5646 11383
rect 5594 11339 5600 11373
rect 5600 11339 5634 11373
rect 5634 11339 5646 11373
rect 5594 11331 5646 11339
rect 5660 11373 5712 11383
rect 5660 11339 5672 11373
rect 5672 11339 5706 11373
rect 5706 11339 5712 11373
rect 5660 11331 5712 11339
rect 5594 11300 5646 11314
rect 5594 11266 5600 11300
rect 5600 11266 5634 11300
rect 5634 11266 5646 11300
rect 5594 11262 5646 11266
rect 5660 11300 5712 11314
rect 5660 11266 5672 11300
rect 5672 11266 5706 11300
rect 5706 11266 5712 11300
rect 5660 11262 5712 11266
rect 5594 11227 5646 11245
rect 5594 11193 5600 11227
rect 5600 11193 5634 11227
rect 5634 11193 5646 11227
rect 5660 11227 5712 11245
rect 5660 11193 5672 11227
rect 5672 11193 5706 11227
rect 5706 11193 5712 11227
rect 5594 11154 5646 11176
rect 5660 11154 5712 11176
rect 5594 11124 5600 11154
rect 5600 11124 5646 11154
rect 5660 11124 5706 11154
rect 5706 11124 5712 11154
rect 5594 11055 5600 11107
rect 5600 11055 5646 11107
rect 5660 11055 5706 11107
rect 5706 11055 5712 11107
rect 5594 10986 5600 11038
rect 5600 10986 5646 11038
rect 5660 10986 5706 11038
rect 5706 10986 5712 11038
rect 5594 10916 5600 10968
rect 5600 10916 5646 10968
rect 5660 10916 5706 10968
rect 5706 10916 5712 10968
rect 5594 10846 5600 10898
rect 5600 10846 5646 10898
rect 5660 10846 5706 10898
rect 5706 10846 5712 10898
rect 5871 10662 5877 10714
rect 5877 10662 5923 10714
rect 5937 10662 5983 10714
rect 5983 10662 5989 10714
rect 5871 10593 5877 10645
rect 5877 10593 5923 10645
rect 5937 10593 5983 10645
rect 5983 10593 5989 10645
rect 5871 10524 5877 10576
rect 5877 10524 5923 10576
rect 5937 10524 5983 10576
rect 5983 10524 5989 10576
rect 5871 10455 5877 10507
rect 5877 10455 5923 10507
rect 5937 10455 5983 10507
rect 5983 10455 5989 10507
rect 5871 10386 5877 10438
rect 5877 10386 5923 10438
rect 5937 10386 5983 10438
rect 5983 10386 5989 10438
rect 5871 10316 5877 10368
rect 5877 10316 5923 10368
rect 5937 10316 5983 10368
rect 5983 10316 5989 10368
rect 5871 10246 5877 10298
rect 5877 10246 5923 10298
rect 5937 10246 5983 10298
rect 5983 10246 5989 10298
rect 5871 10176 5877 10228
rect 5877 10176 5923 10228
rect 5937 10176 5983 10228
rect 5983 10176 5989 10228
rect 5871 10112 5877 10158
rect 5877 10112 5923 10158
rect 5937 10112 5983 10158
rect 5983 10112 5989 10158
rect 5871 10106 5923 10112
rect 5937 10106 5989 10112
rect 6148 11446 6200 11452
rect 6148 11412 6154 11446
rect 6154 11412 6188 11446
rect 6188 11412 6200 11446
rect 6148 11400 6200 11412
rect 6214 11446 6266 11452
rect 6214 11412 6226 11446
rect 6226 11412 6260 11446
rect 6260 11412 6266 11446
rect 6214 11400 6266 11412
rect 6148 11373 6200 11383
rect 6148 11339 6154 11373
rect 6154 11339 6188 11373
rect 6188 11339 6200 11373
rect 6148 11331 6200 11339
rect 6214 11373 6266 11383
rect 6214 11339 6226 11373
rect 6226 11339 6260 11373
rect 6260 11339 6266 11373
rect 6214 11331 6266 11339
rect 6148 11300 6200 11314
rect 6148 11266 6154 11300
rect 6154 11266 6188 11300
rect 6188 11266 6200 11300
rect 6148 11262 6200 11266
rect 6214 11300 6266 11314
rect 6214 11266 6226 11300
rect 6226 11266 6260 11300
rect 6260 11266 6266 11300
rect 6214 11262 6266 11266
rect 6148 11227 6200 11245
rect 6148 11193 6154 11227
rect 6154 11193 6188 11227
rect 6188 11193 6200 11227
rect 6214 11227 6266 11245
rect 6214 11193 6226 11227
rect 6226 11193 6260 11227
rect 6260 11193 6266 11227
rect 6148 11154 6200 11176
rect 6214 11154 6266 11176
rect 6148 11124 6154 11154
rect 6154 11124 6200 11154
rect 6214 11124 6260 11154
rect 6260 11124 6266 11154
rect 6148 11055 6154 11107
rect 6154 11055 6200 11107
rect 6214 11055 6260 11107
rect 6260 11055 6266 11107
rect 6148 10986 6154 11038
rect 6154 10986 6200 11038
rect 6214 10986 6260 11038
rect 6260 10986 6266 11038
rect 6148 10916 6154 10968
rect 6154 10916 6200 10968
rect 6214 10916 6260 10968
rect 6260 10916 6266 10968
rect 6148 10846 6154 10898
rect 6154 10846 6200 10898
rect 6214 10846 6260 10898
rect 6260 10846 6266 10898
rect 6425 10662 6431 10714
rect 6431 10662 6477 10714
rect 6491 10662 6537 10714
rect 6537 10662 6543 10714
rect 6425 10593 6431 10645
rect 6431 10593 6477 10645
rect 6491 10593 6537 10645
rect 6537 10593 6543 10645
rect 6425 10524 6431 10576
rect 6431 10524 6477 10576
rect 6491 10524 6537 10576
rect 6537 10524 6543 10576
rect 6425 10455 6431 10507
rect 6431 10455 6477 10507
rect 6491 10455 6537 10507
rect 6537 10455 6543 10507
rect 6425 10386 6431 10438
rect 6431 10386 6477 10438
rect 6491 10386 6537 10438
rect 6537 10386 6543 10438
rect 6425 10316 6431 10368
rect 6431 10316 6477 10368
rect 6491 10316 6537 10368
rect 6537 10316 6543 10368
rect 6425 10246 6431 10298
rect 6431 10246 6477 10298
rect 6491 10246 6537 10298
rect 6537 10246 6543 10298
rect 6425 10176 6431 10228
rect 6431 10176 6477 10228
rect 6491 10176 6537 10228
rect 6537 10176 6543 10228
rect 6425 10112 6431 10158
rect 6431 10112 6477 10158
rect 6491 10112 6537 10158
rect 6537 10112 6543 10158
rect 6425 10106 6477 10112
rect 6491 10106 6543 10112
rect 6702 11446 6754 11452
rect 6702 11412 6708 11446
rect 6708 11412 6742 11446
rect 6742 11412 6754 11446
rect 6702 11400 6754 11412
rect 6768 11446 6820 11452
rect 6768 11412 6780 11446
rect 6780 11412 6814 11446
rect 6814 11412 6820 11446
rect 6768 11400 6820 11412
rect 6702 11373 6754 11383
rect 6702 11339 6708 11373
rect 6708 11339 6742 11373
rect 6742 11339 6754 11373
rect 6702 11331 6754 11339
rect 6768 11373 6820 11383
rect 6768 11339 6780 11373
rect 6780 11339 6814 11373
rect 6814 11339 6820 11373
rect 6768 11331 6820 11339
rect 6702 11300 6754 11314
rect 6702 11266 6708 11300
rect 6708 11266 6742 11300
rect 6742 11266 6754 11300
rect 6702 11262 6754 11266
rect 6768 11300 6820 11314
rect 6768 11266 6780 11300
rect 6780 11266 6814 11300
rect 6814 11266 6820 11300
rect 6768 11262 6820 11266
rect 6702 11227 6754 11245
rect 6702 11193 6708 11227
rect 6708 11193 6742 11227
rect 6742 11193 6754 11227
rect 6768 11227 6820 11245
rect 6768 11193 6780 11227
rect 6780 11193 6814 11227
rect 6814 11193 6820 11227
rect 6702 11154 6754 11176
rect 6768 11154 6820 11176
rect 6702 11124 6708 11154
rect 6708 11124 6754 11154
rect 6768 11124 6814 11154
rect 6814 11124 6820 11154
rect 6702 11055 6708 11107
rect 6708 11055 6754 11107
rect 6768 11055 6814 11107
rect 6814 11055 6820 11107
rect 6702 10986 6708 11038
rect 6708 10986 6754 11038
rect 6768 10986 6814 11038
rect 6814 10986 6820 11038
rect 6702 10916 6708 10968
rect 6708 10916 6754 10968
rect 6768 10916 6814 10968
rect 6814 10916 6820 10968
rect 6702 10846 6708 10898
rect 6708 10846 6754 10898
rect 6768 10846 6814 10898
rect 6814 10846 6820 10898
rect 6979 10662 6985 10714
rect 6985 10662 7031 10714
rect 7045 10662 7091 10714
rect 7091 10662 7097 10714
rect 6979 10593 6985 10645
rect 6985 10593 7031 10645
rect 7045 10593 7091 10645
rect 7091 10593 7097 10645
rect 6979 10524 6985 10576
rect 6985 10524 7031 10576
rect 7045 10524 7091 10576
rect 7091 10524 7097 10576
rect 6979 10455 6985 10507
rect 6985 10455 7031 10507
rect 7045 10455 7091 10507
rect 7091 10455 7097 10507
rect 6979 10386 6985 10438
rect 6985 10386 7031 10438
rect 7045 10386 7091 10438
rect 7091 10386 7097 10438
rect 6979 10316 6985 10368
rect 6985 10316 7031 10368
rect 7045 10316 7091 10368
rect 7091 10316 7097 10368
rect 6979 10246 6985 10298
rect 6985 10246 7031 10298
rect 7045 10246 7091 10298
rect 7091 10246 7097 10298
rect 6979 10176 6985 10228
rect 6985 10176 7031 10228
rect 7045 10176 7091 10228
rect 7091 10176 7097 10228
rect 6979 10112 6985 10158
rect 6985 10112 7031 10158
rect 7045 10112 7091 10158
rect 7091 10112 7097 10158
rect 6979 10106 7031 10112
rect 7045 10106 7097 10112
rect 7256 11446 7308 11452
rect 7256 11412 7262 11446
rect 7262 11412 7296 11446
rect 7296 11412 7308 11446
rect 7256 11400 7308 11412
rect 7322 11446 7374 11452
rect 7322 11412 7334 11446
rect 7334 11412 7368 11446
rect 7368 11412 7374 11446
rect 7322 11400 7374 11412
rect 7256 11373 7308 11383
rect 7256 11339 7262 11373
rect 7262 11339 7296 11373
rect 7296 11339 7308 11373
rect 7256 11331 7308 11339
rect 7322 11373 7374 11383
rect 7322 11339 7334 11373
rect 7334 11339 7368 11373
rect 7368 11339 7374 11373
rect 7322 11331 7374 11339
rect 7256 11300 7308 11314
rect 7256 11266 7262 11300
rect 7262 11266 7296 11300
rect 7296 11266 7308 11300
rect 7256 11262 7308 11266
rect 7322 11300 7374 11314
rect 7322 11266 7334 11300
rect 7334 11266 7368 11300
rect 7368 11266 7374 11300
rect 7322 11262 7374 11266
rect 7256 11227 7308 11245
rect 7256 11193 7262 11227
rect 7262 11193 7296 11227
rect 7296 11193 7308 11227
rect 7322 11227 7374 11245
rect 7322 11193 7334 11227
rect 7334 11193 7368 11227
rect 7368 11193 7374 11227
rect 7256 11154 7308 11176
rect 7322 11154 7374 11176
rect 7256 11124 7262 11154
rect 7262 11124 7308 11154
rect 7322 11124 7368 11154
rect 7368 11124 7374 11154
rect 7256 11055 7262 11107
rect 7262 11055 7308 11107
rect 7322 11055 7368 11107
rect 7368 11055 7374 11107
rect 7256 10986 7262 11038
rect 7262 10986 7308 11038
rect 7322 10986 7368 11038
rect 7368 10986 7374 11038
rect 7256 10916 7262 10968
rect 7262 10916 7308 10968
rect 7322 10916 7368 10968
rect 7368 10916 7374 10968
rect 7256 10846 7262 10898
rect 7262 10846 7308 10898
rect 7322 10846 7368 10898
rect 7368 10846 7374 10898
rect 7533 10662 7539 10714
rect 7539 10662 7585 10714
rect 7599 10662 7645 10714
rect 7645 10662 7651 10714
rect 7533 10593 7539 10645
rect 7539 10593 7585 10645
rect 7599 10593 7645 10645
rect 7645 10593 7651 10645
rect 7533 10524 7539 10576
rect 7539 10524 7585 10576
rect 7599 10524 7645 10576
rect 7645 10524 7651 10576
rect 7533 10455 7539 10507
rect 7539 10455 7585 10507
rect 7599 10455 7645 10507
rect 7645 10455 7651 10507
rect 7533 10386 7539 10438
rect 7539 10386 7585 10438
rect 7599 10386 7645 10438
rect 7645 10386 7651 10438
rect 7533 10316 7539 10368
rect 7539 10316 7585 10368
rect 7599 10316 7645 10368
rect 7645 10316 7651 10368
rect 7533 10246 7539 10298
rect 7539 10246 7585 10298
rect 7599 10246 7645 10298
rect 7645 10246 7651 10298
rect 7533 10176 7539 10228
rect 7539 10176 7585 10228
rect 7599 10176 7645 10228
rect 7645 10176 7651 10228
rect 7533 10112 7539 10158
rect 7539 10112 7585 10158
rect 7599 10112 7645 10158
rect 7645 10112 7651 10158
rect 7533 10106 7585 10112
rect 7599 10106 7651 10112
rect 7810 11446 7862 11452
rect 7810 11412 7816 11446
rect 7816 11412 7850 11446
rect 7850 11412 7862 11446
rect 7810 11400 7862 11412
rect 7876 11446 7928 11452
rect 7876 11412 7888 11446
rect 7888 11412 7922 11446
rect 7922 11412 7928 11446
rect 7876 11400 7928 11412
rect 7810 11373 7862 11383
rect 7810 11339 7816 11373
rect 7816 11339 7850 11373
rect 7850 11339 7862 11373
rect 7810 11331 7862 11339
rect 7876 11373 7928 11383
rect 7876 11339 7888 11373
rect 7888 11339 7922 11373
rect 7922 11339 7928 11373
rect 7876 11331 7928 11339
rect 7810 11300 7862 11314
rect 7810 11266 7816 11300
rect 7816 11266 7850 11300
rect 7850 11266 7862 11300
rect 7810 11262 7862 11266
rect 7876 11300 7928 11314
rect 7876 11266 7888 11300
rect 7888 11266 7922 11300
rect 7922 11266 7928 11300
rect 7876 11262 7928 11266
rect 7810 11227 7862 11245
rect 7810 11193 7816 11227
rect 7816 11193 7850 11227
rect 7850 11193 7862 11227
rect 7876 11227 7928 11245
rect 7876 11193 7888 11227
rect 7888 11193 7922 11227
rect 7922 11193 7928 11227
rect 7810 11154 7862 11176
rect 7876 11154 7928 11176
rect 7810 11124 7816 11154
rect 7816 11124 7862 11154
rect 7876 11124 7922 11154
rect 7922 11124 7928 11154
rect 7810 11055 7816 11107
rect 7816 11055 7862 11107
rect 7876 11055 7922 11107
rect 7922 11055 7928 11107
rect 7810 10986 7816 11038
rect 7816 10986 7862 11038
rect 7876 10986 7922 11038
rect 7922 10986 7928 11038
rect 7810 10916 7816 10968
rect 7816 10916 7862 10968
rect 7876 10916 7922 10968
rect 7922 10916 7928 10968
rect 7810 10846 7816 10898
rect 7816 10846 7862 10898
rect 7876 10846 7922 10898
rect 7922 10846 7928 10898
rect 8047 11448 8050 11456
rect 8050 11448 8084 11456
rect 8084 11448 8099 11456
rect 8047 11409 8099 11448
rect 8047 11404 8050 11409
rect 8050 11404 8084 11409
rect 8084 11404 8099 11409
rect 8169 11448 8184 11456
rect 8184 11448 8218 11456
rect 8218 11448 8221 11456
rect 8169 11409 8221 11448
rect 8169 11404 8184 11409
rect 8184 11404 8218 11409
rect 8218 11404 8221 11409
rect 8047 11375 8050 11387
rect 8050 11375 8084 11387
rect 8084 11375 8099 11387
rect 8047 11336 8099 11375
rect 8047 11335 8050 11336
rect 8050 11335 8084 11336
rect 8084 11335 8099 11336
rect 8169 11375 8184 11387
rect 8184 11375 8218 11387
rect 8218 11375 8221 11387
rect 8169 11336 8221 11375
rect 8169 11335 8184 11336
rect 8184 11335 8218 11336
rect 8218 11335 8221 11336
rect 8047 11302 8050 11318
rect 8050 11302 8084 11318
rect 8084 11302 8099 11318
rect 8047 11266 8099 11302
rect 8169 11302 8184 11318
rect 8184 11302 8218 11318
rect 8218 11302 8221 11318
rect 8169 11266 8221 11302
rect 8047 11229 8050 11249
rect 8050 11229 8084 11249
rect 8084 11229 8099 11249
rect 8047 11197 8099 11229
rect 8169 11229 8184 11249
rect 8184 11229 8218 11249
rect 8218 11229 8221 11249
rect 8169 11197 8221 11229
rect 8047 11156 8050 11180
rect 8050 11156 8084 11180
rect 8084 11156 8099 11180
rect 8047 11128 8099 11156
rect 8169 11156 8184 11180
rect 8184 11156 8218 11180
rect 8218 11156 8221 11180
rect 8169 11128 8221 11156
rect 8047 11083 8050 11110
rect 8050 11083 8084 11110
rect 8084 11083 8099 11110
rect 8047 11058 8099 11083
rect 8169 11083 8184 11110
rect 8184 11083 8218 11110
rect 8218 11083 8221 11110
rect 8169 11058 8221 11083
rect 8047 11010 8050 11040
rect 8050 11010 8084 11040
rect 8084 11010 8099 11040
rect 8047 10988 8099 11010
rect 8169 11010 8184 11040
rect 8184 11010 8218 11040
rect 8218 11010 8221 11040
rect 8169 10988 8221 11010
rect 8047 10937 8050 10970
rect 8050 10937 8084 10970
rect 8084 10937 8099 10970
rect 8047 10918 8099 10937
rect 8169 10937 8184 10970
rect 8184 10937 8218 10970
rect 8218 10937 8221 10970
rect 8169 10918 8221 10937
rect 8047 10898 8099 10900
rect 8047 10864 8050 10898
rect 8050 10864 8084 10898
rect 8084 10864 8099 10898
rect 8047 10848 8099 10864
rect 8169 10898 8221 10900
rect 8169 10864 8184 10898
rect 8184 10864 8218 10898
rect 8218 10864 8221 10898
rect 8169 10848 8221 10864
rect 2580 10008 2632 10060
rect 2660 10008 2712 10060
rect 8429 26967 8481 27019
rect 8515 26967 8535 27019
rect 8535 26967 8567 27019
rect 8429 26899 8481 26951
rect 8515 26899 8535 26951
rect 8535 26899 8567 26951
rect 5204 9449 5256 9458
rect 5204 9415 5232 9449
rect 5232 9415 5256 9449
rect 5204 9406 5256 9415
rect 5268 9449 5320 9458
rect 5268 9415 5270 9449
rect 5270 9415 5304 9449
rect 5304 9415 5320 9449
rect 5268 9406 5320 9415
rect 5332 9449 5384 9458
rect 5332 9415 5342 9449
rect 5342 9415 5376 9449
rect 5376 9415 5384 9449
rect 5332 9406 5384 9415
rect 5396 9449 5448 9458
rect 5396 9415 5414 9449
rect 5414 9415 5448 9449
rect 5396 9406 5448 9415
rect 5460 9449 5512 9458
rect 5524 9449 5576 9458
rect 5588 9449 5640 9458
rect 5652 9449 5704 9458
rect 5716 9449 5768 9458
rect 5780 9449 5832 9458
rect 5460 9415 5486 9449
rect 5486 9415 5512 9449
rect 5524 9415 5558 9449
rect 5558 9415 5576 9449
rect 5588 9415 5592 9449
rect 5592 9415 5630 9449
rect 5630 9415 5640 9449
rect 5652 9415 5664 9449
rect 5664 9415 5702 9449
rect 5702 9415 5704 9449
rect 5716 9415 5736 9449
rect 5736 9415 5768 9449
rect 5780 9415 5808 9449
rect 5808 9415 5832 9449
rect 5460 9406 5512 9415
rect 5524 9406 5576 9415
rect 5588 9406 5640 9415
rect 5652 9406 5704 9415
rect 5716 9406 5768 9415
rect 5780 9406 5832 9415
rect 5844 9449 5896 9458
rect 5844 9415 5846 9449
rect 5846 9415 5880 9449
rect 5880 9415 5896 9449
rect 5844 9406 5896 9415
rect 5908 9449 5960 9458
rect 5908 9415 5918 9449
rect 5918 9415 5952 9449
rect 5952 9415 5960 9449
rect 5908 9406 5960 9415
rect 5972 9449 6024 9458
rect 5972 9415 5990 9449
rect 5990 9415 6024 9449
rect 5972 9406 6024 9415
rect 6036 9449 6088 9458
rect 6100 9449 6152 9458
rect 6164 9449 6216 9458
rect 6228 9449 6280 9458
rect 6292 9449 6344 9458
rect 6356 9449 6408 9458
rect 6036 9415 6062 9449
rect 6062 9415 6088 9449
rect 6100 9415 6134 9449
rect 6134 9415 6152 9449
rect 6164 9415 6168 9449
rect 6168 9415 6206 9449
rect 6206 9415 6216 9449
rect 6228 9415 6240 9449
rect 6240 9415 6278 9449
rect 6278 9415 6280 9449
rect 6292 9415 6312 9449
rect 6312 9415 6344 9449
rect 6356 9415 6384 9449
rect 6384 9415 6408 9449
rect 6036 9406 6088 9415
rect 6100 9406 6152 9415
rect 6164 9406 6216 9415
rect 6228 9406 6280 9415
rect 6292 9406 6344 9415
rect 6356 9406 6408 9415
rect 6420 9449 6472 9458
rect 6420 9415 6422 9449
rect 6422 9415 6456 9449
rect 6456 9415 6472 9449
rect 6420 9406 6472 9415
rect 6484 9449 6536 9458
rect 6484 9415 6494 9449
rect 6494 9415 6528 9449
rect 6528 9415 6536 9449
rect 6484 9406 6536 9415
rect 6548 9449 6600 9458
rect 6548 9415 6566 9449
rect 6566 9415 6600 9449
rect 6548 9406 6600 9415
rect 6612 9449 6664 9458
rect 6676 9449 6728 9458
rect 6740 9449 6792 9458
rect 6804 9449 6856 9458
rect 6868 9449 6920 9458
rect 6932 9449 6984 9458
rect 6612 9415 6638 9449
rect 6638 9415 6664 9449
rect 6676 9415 6710 9449
rect 6710 9415 6728 9449
rect 6740 9415 6744 9449
rect 6744 9415 6782 9449
rect 6782 9415 6792 9449
rect 6804 9415 6816 9449
rect 6816 9415 6854 9449
rect 6854 9415 6856 9449
rect 6868 9415 6888 9449
rect 6888 9415 6920 9449
rect 6932 9415 6960 9449
rect 6960 9415 6984 9449
rect 6612 9406 6664 9415
rect 6676 9406 6728 9415
rect 6740 9406 6792 9415
rect 6804 9406 6856 9415
rect 6868 9406 6920 9415
rect 6932 9406 6984 9415
rect 6996 9449 7048 9458
rect 6996 9415 6998 9449
rect 6998 9415 7032 9449
rect 7032 9415 7048 9449
rect 6996 9406 7048 9415
rect 7060 9449 7112 9458
rect 7060 9415 7070 9449
rect 7070 9415 7104 9449
rect 7104 9415 7112 9449
rect 7060 9406 7112 9415
rect 7124 9449 7176 9458
rect 7124 9415 7142 9449
rect 7142 9415 7176 9449
rect 7124 9406 7176 9415
rect 7188 9449 7240 9458
rect 7252 9449 7304 9458
rect 7316 9449 7368 9458
rect 7188 9415 7214 9449
rect 7214 9415 7240 9449
rect 7252 9415 7286 9449
rect 7286 9415 7304 9449
rect 7316 9415 7320 9449
rect 7320 9415 7358 9449
rect 7358 9415 7368 9449
rect 7188 9406 7240 9415
rect 7252 9406 7304 9415
rect 7316 9406 7368 9415
rect 2474 9341 2526 9350
rect 2474 9307 2480 9341
rect 2480 9307 2514 9341
rect 2514 9307 2526 9341
rect 2474 9298 2526 9307
rect 2539 9341 2591 9350
rect 2539 9307 2553 9341
rect 2553 9307 2587 9341
rect 2587 9307 2591 9341
rect 2539 9298 2591 9307
rect 2604 9341 2656 9350
rect 2604 9307 2626 9341
rect 2626 9307 2656 9341
rect 2604 9298 2656 9307
rect 5204 8701 7368 8727
rect 5204 8667 5737 8701
rect 5737 8667 5771 8701
rect 5771 8667 7368 8701
rect 5204 8628 7368 8667
rect 5204 8594 5737 8628
rect 5737 8594 5771 8628
rect 5771 8594 7368 8628
rect 5204 8554 7368 8594
rect 5204 8520 5737 8554
rect 5737 8520 5771 8554
rect 5771 8520 7368 8554
rect 5204 8480 7368 8520
rect 5204 8446 5737 8480
rect 5737 8446 5771 8480
rect 5771 8446 7368 8480
rect 5204 8406 7368 8446
rect 5204 8372 5737 8406
rect 5737 8372 5771 8406
rect 5771 8372 7368 8406
rect 5204 8332 7368 8372
rect 5204 8298 5737 8332
rect 5737 8298 5771 8332
rect 5771 8298 7368 8332
rect 5204 8258 7368 8298
rect 5204 8224 5737 8258
rect 5737 8224 5771 8258
rect 5771 8224 7368 8258
rect 5204 8184 7368 8224
rect 5204 8150 5737 8184
rect 5737 8150 5771 8184
rect 5771 8150 7368 8184
rect 5204 8110 7368 8150
rect 5204 8076 5737 8110
rect 5737 8076 5771 8110
rect 5771 8076 7368 8110
rect 5204 8036 7368 8076
rect 5204 8002 5737 8036
rect 5737 8002 5771 8036
rect 5771 8002 7368 8036
rect 5204 7962 7368 8002
rect 5204 7928 5737 7962
rect 5737 7928 5771 7962
rect 5771 7928 7368 7962
rect 5204 7888 7368 7928
rect 5204 7854 5737 7888
rect 5737 7854 5771 7888
rect 5771 7854 7368 7888
rect 5204 7843 7368 7854
rect 5204 7681 5256 7690
rect 5268 7681 5320 7690
rect 5332 7681 5384 7690
rect 5396 7681 5448 7690
rect 5460 7681 5512 7690
rect 5204 7647 5237 7681
rect 5237 7647 5256 7681
rect 5268 7647 5271 7681
rect 5271 7647 5309 7681
rect 5309 7647 5320 7681
rect 5332 7647 5343 7681
rect 5343 7647 5381 7681
rect 5381 7647 5384 7681
rect 5396 7647 5415 7681
rect 5415 7647 5448 7681
rect 5460 7647 5487 7681
rect 5487 7647 5512 7681
rect 5204 7638 5256 7647
rect 5268 7638 5320 7647
rect 5332 7638 5384 7647
rect 5396 7638 5448 7647
rect 5460 7638 5512 7647
rect 5524 7681 5576 7690
rect 5524 7647 5525 7681
rect 5525 7647 5559 7681
rect 5559 7647 5576 7681
rect 5524 7638 5576 7647
rect 5588 7681 5640 7690
rect 5588 7647 5597 7681
rect 5597 7647 5631 7681
rect 5631 7647 5640 7681
rect 5588 7638 5640 7647
rect 5652 7681 5704 7690
rect 5652 7647 5669 7681
rect 5669 7647 5703 7681
rect 5703 7647 5704 7681
rect 5652 7638 5704 7647
rect 5716 7681 5768 7690
rect 5780 7681 5832 7690
rect 5844 7681 5896 7690
rect 5908 7681 5960 7690
rect 5972 7681 6024 7690
rect 6036 7681 6088 7690
rect 5716 7647 5741 7681
rect 5741 7647 5768 7681
rect 5780 7647 5813 7681
rect 5813 7647 5832 7681
rect 5844 7647 5847 7681
rect 5847 7647 5885 7681
rect 5885 7647 5896 7681
rect 5908 7647 5919 7681
rect 5919 7647 5957 7681
rect 5957 7647 5960 7681
rect 5972 7647 5991 7681
rect 5991 7647 6024 7681
rect 6036 7647 6063 7681
rect 6063 7647 6088 7681
rect 5716 7638 5768 7647
rect 5780 7638 5832 7647
rect 5844 7638 5896 7647
rect 5908 7638 5960 7647
rect 5972 7638 6024 7647
rect 6036 7638 6088 7647
rect 6100 7681 6152 7690
rect 6100 7647 6101 7681
rect 6101 7647 6135 7681
rect 6135 7647 6152 7681
rect 6100 7638 6152 7647
rect 6164 7681 6216 7690
rect 6164 7647 6173 7681
rect 6173 7647 6207 7681
rect 6207 7647 6216 7681
rect 6164 7638 6216 7647
rect 6228 7681 6280 7690
rect 6228 7647 6245 7681
rect 6245 7647 6279 7681
rect 6279 7647 6280 7681
rect 6228 7638 6280 7647
rect 6292 7681 6344 7690
rect 6356 7681 6408 7690
rect 6420 7681 6472 7690
rect 6484 7681 6536 7690
rect 6548 7681 6600 7690
rect 6612 7681 6664 7690
rect 6292 7647 6317 7681
rect 6317 7647 6344 7681
rect 6356 7647 6389 7681
rect 6389 7647 6408 7681
rect 6420 7647 6423 7681
rect 6423 7647 6461 7681
rect 6461 7647 6472 7681
rect 6484 7647 6495 7681
rect 6495 7647 6533 7681
rect 6533 7647 6536 7681
rect 6548 7647 6567 7681
rect 6567 7647 6600 7681
rect 6612 7647 6639 7681
rect 6639 7647 6664 7681
rect 6292 7638 6344 7647
rect 6356 7638 6408 7647
rect 6420 7638 6472 7647
rect 6484 7638 6536 7647
rect 6548 7638 6600 7647
rect 6612 7638 6664 7647
rect 6676 7681 6728 7690
rect 6676 7647 6677 7681
rect 6677 7647 6711 7681
rect 6711 7647 6728 7681
rect 6676 7638 6728 7647
rect 6740 7681 6792 7690
rect 6740 7647 6749 7681
rect 6749 7647 6783 7681
rect 6783 7647 6792 7681
rect 6740 7638 6792 7647
rect 6804 7681 6856 7690
rect 6804 7647 6821 7681
rect 6821 7647 6855 7681
rect 6855 7647 6856 7681
rect 6804 7638 6856 7647
rect 6868 7681 6920 7690
rect 6932 7681 6984 7690
rect 6996 7681 7048 7690
rect 7060 7681 7112 7690
rect 7124 7681 7176 7690
rect 7188 7681 7240 7690
rect 6868 7647 6893 7681
rect 6893 7647 6920 7681
rect 6932 7647 6965 7681
rect 6965 7647 6984 7681
rect 6996 7647 6999 7681
rect 6999 7647 7037 7681
rect 7037 7647 7048 7681
rect 7060 7647 7071 7681
rect 7071 7647 7109 7681
rect 7109 7647 7112 7681
rect 7124 7647 7143 7681
rect 7143 7647 7176 7681
rect 7188 7647 7215 7681
rect 7215 7647 7240 7681
rect 6868 7638 6920 7647
rect 6932 7638 6984 7647
rect 6996 7638 7048 7647
rect 7060 7638 7112 7647
rect 7124 7638 7176 7647
rect 7188 7638 7240 7647
rect 7252 7681 7304 7690
rect 7252 7647 7253 7681
rect 7253 7647 7287 7681
rect 7287 7647 7304 7681
rect 7252 7638 7304 7647
rect 7316 7681 7368 7690
rect 7316 7647 7325 7681
rect 7325 7647 7359 7681
rect 7359 7647 7368 7681
rect 7316 7638 7368 7647
rect 2474 7540 2526 7549
rect 2474 7506 2480 7540
rect 2480 7506 2514 7540
rect 2514 7506 2526 7540
rect 2474 7497 2526 7506
rect 2539 7540 2591 7549
rect 2539 7506 2553 7540
rect 2553 7506 2587 7540
rect 2587 7506 2591 7540
rect 2539 7497 2591 7506
rect 2604 7540 2656 7549
rect 2604 7506 2626 7540
rect 2626 7506 2656 7540
rect 2604 7497 2656 7506
rect 5204 6901 7368 6927
rect 5204 6867 5737 6901
rect 5737 6867 5771 6901
rect 5771 6867 7368 6901
rect 5204 6828 7368 6867
rect 5204 6794 5737 6828
rect 5737 6794 5771 6828
rect 5771 6794 7368 6828
rect 5204 6754 7368 6794
rect 5204 6720 5737 6754
rect 5737 6720 5771 6754
rect 5771 6720 7368 6754
rect 5204 6680 7368 6720
rect 5204 6646 5737 6680
rect 5737 6646 5771 6680
rect 5771 6646 7368 6680
rect 5204 6606 7368 6646
rect 5204 6572 5737 6606
rect 5737 6572 5771 6606
rect 5771 6572 7368 6606
rect 5204 6532 7368 6572
rect 5204 6498 5737 6532
rect 5737 6498 5771 6532
rect 5771 6498 7368 6532
rect 5204 6458 7368 6498
rect 5204 6424 5737 6458
rect 5737 6424 5771 6458
rect 5771 6424 7368 6458
rect 5204 6384 7368 6424
rect 5204 6350 5737 6384
rect 5737 6350 5771 6384
rect 5771 6350 7368 6384
rect 5204 6310 7368 6350
rect 5204 6276 5737 6310
rect 5737 6276 5771 6310
rect 5771 6276 7368 6310
rect 5204 6236 7368 6276
rect 5204 6202 5737 6236
rect 5737 6202 5771 6236
rect 5771 6202 7368 6236
rect 5204 6162 7368 6202
rect 5204 6128 5737 6162
rect 5737 6128 5771 6162
rect 5771 6128 7368 6162
rect 5204 6088 7368 6128
rect 5204 6054 5737 6088
rect 5737 6054 5771 6088
rect 5771 6054 7368 6088
rect 5204 6043 7368 6054
rect 5204 5841 5256 5850
rect 5204 5807 5210 5841
rect 5210 5807 5244 5841
rect 5244 5807 5256 5841
rect 5204 5798 5256 5807
rect 5268 5841 5320 5850
rect 5268 5807 5283 5841
rect 5283 5807 5317 5841
rect 5317 5807 5320 5841
rect 5268 5798 5320 5807
rect 5332 5841 5384 5850
rect 5396 5841 5448 5850
rect 5460 5841 5512 5850
rect 5524 5841 5576 5850
rect 5588 5841 5640 5850
rect 5652 5841 5704 5850
rect 5332 5807 5356 5841
rect 5356 5807 5384 5841
rect 5396 5807 5429 5841
rect 5429 5807 5448 5841
rect 5460 5807 5463 5841
rect 5463 5807 5502 5841
rect 5502 5807 5512 5841
rect 5524 5807 5536 5841
rect 5536 5807 5575 5841
rect 5575 5807 5576 5841
rect 5588 5807 5609 5841
rect 5609 5807 5640 5841
rect 5652 5807 5682 5841
rect 5682 5807 5704 5841
rect 5332 5798 5384 5807
rect 5396 5798 5448 5807
rect 5460 5798 5512 5807
rect 5524 5798 5576 5807
rect 5588 5798 5640 5807
rect 5652 5798 5704 5807
rect 5716 5841 5768 5850
rect 5716 5807 5721 5841
rect 5721 5807 5755 5841
rect 5755 5807 5768 5841
rect 5716 5798 5768 5807
rect 5780 5841 5832 5850
rect 5780 5807 5794 5841
rect 5794 5807 5828 5841
rect 5828 5807 5832 5841
rect 5780 5798 5832 5807
rect 5844 5841 5896 5850
rect 5908 5841 5960 5850
rect 5972 5841 6024 5850
rect 6036 5841 6088 5850
rect 6100 5841 6152 5850
rect 6164 5841 6216 5850
rect 5844 5807 5867 5841
rect 5867 5807 5896 5841
rect 5908 5807 5940 5841
rect 5940 5807 5960 5841
rect 5972 5807 5974 5841
rect 5974 5807 6013 5841
rect 6013 5807 6024 5841
rect 6036 5807 6047 5841
rect 6047 5807 6086 5841
rect 6086 5807 6088 5841
rect 6100 5807 6120 5841
rect 6120 5807 6152 5841
rect 6164 5807 6193 5841
rect 6193 5807 6216 5841
rect 5844 5798 5896 5807
rect 5908 5798 5960 5807
rect 5972 5798 6024 5807
rect 6036 5798 6088 5807
rect 6100 5798 6152 5807
rect 6164 5798 6216 5807
rect 6228 5841 6280 5850
rect 6228 5807 6232 5841
rect 6232 5807 6266 5841
rect 6266 5807 6280 5841
rect 6228 5798 6280 5807
rect 6292 5841 6344 5850
rect 6292 5807 6305 5841
rect 6305 5807 6339 5841
rect 6339 5807 6344 5841
rect 6292 5798 6344 5807
rect 6356 5841 6408 5850
rect 6420 5841 6472 5850
rect 6484 5841 6536 5850
rect 6548 5841 6600 5850
rect 6612 5841 6664 5850
rect 6676 5841 6728 5850
rect 6356 5807 6378 5841
rect 6378 5807 6408 5841
rect 6420 5807 6451 5841
rect 6451 5807 6472 5841
rect 6484 5807 6485 5841
rect 6485 5807 6524 5841
rect 6524 5807 6536 5841
rect 6548 5807 6558 5841
rect 6558 5807 6597 5841
rect 6597 5807 6600 5841
rect 6612 5807 6631 5841
rect 6631 5807 6664 5841
rect 6676 5807 6704 5841
rect 6704 5807 6728 5841
rect 6356 5798 6408 5807
rect 6420 5798 6472 5807
rect 6484 5798 6536 5807
rect 6548 5798 6600 5807
rect 6612 5798 6664 5807
rect 6676 5798 6728 5807
rect 6740 5841 6792 5850
rect 6740 5807 6743 5841
rect 6743 5807 6777 5841
rect 6777 5807 6792 5841
rect 6740 5798 6792 5807
rect 6804 5841 6856 5850
rect 6804 5807 6816 5841
rect 6816 5807 6850 5841
rect 6850 5807 6856 5841
rect 6804 5798 6856 5807
rect 6868 5841 6920 5850
rect 6932 5841 6984 5850
rect 6996 5841 7048 5850
rect 7060 5841 7112 5850
rect 7124 5841 7176 5850
rect 7188 5841 7240 5850
rect 6868 5807 6889 5841
rect 6889 5807 6920 5841
rect 6932 5807 6962 5841
rect 6962 5807 6984 5841
rect 6996 5807 7035 5841
rect 7035 5807 7048 5841
rect 7060 5807 7069 5841
rect 7069 5807 7108 5841
rect 7108 5807 7112 5841
rect 7124 5807 7142 5841
rect 7142 5807 7176 5841
rect 7188 5807 7215 5841
rect 7215 5807 7240 5841
rect 6868 5798 6920 5807
rect 6932 5798 6984 5807
rect 6996 5798 7048 5807
rect 7060 5798 7112 5807
rect 7124 5798 7176 5807
rect 7188 5798 7240 5807
rect 7252 5841 7304 5850
rect 7252 5807 7253 5841
rect 7253 5807 7287 5841
rect 7287 5807 7304 5841
rect 7252 5798 7304 5807
rect 7316 5841 7368 5850
rect 7316 5807 7325 5841
rect 7325 5807 7359 5841
rect 7359 5807 7368 5841
rect 7316 5798 7368 5807
rect 2474 5602 2526 5654
rect 2539 5602 2591 5654
rect 2604 5645 2656 5654
rect 2604 5611 2640 5645
rect 2640 5611 2656 5645
rect 2604 5602 2656 5611
rect 2798 5505 2850 5557
rect 2891 5505 2943 5557
rect 2983 5505 3035 5557
rect 2798 5427 2850 5479
rect 2891 5427 2943 5479
rect 2983 5427 3035 5479
rect 5204 4691 5256 4743
rect 5336 4719 5388 4743
rect 5336 4691 5347 4719
rect 5347 4691 5381 4719
rect 5381 4691 5388 4719
rect 5468 4691 5520 4743
rect 5600 4691 5652 4743
rect 5732 4691 5784 4743
rect 5864 4691 5916 4743
rect 5996 4691 6048 4743
rect 6128 4691 6180 4743
rect 6260 4691 6312 4743
rect 6392 4691 6444 4743
rect 6524 4691 6576 4743
rect 6656 4691 6708 4743
rect 6788 4691 6840 4743
rect 6920 4691 6972 4743
rect 7052 4719 7104 4743
rect 7052 4691 7059 4719
rect 7059 4691 7093 4719
rect 7093 4691 7104 4719
rect 7184 4691 7236 4743
rect 7316 4691 7368 4743
rect 5204 4583 5256 4635
rect 5336 4610 5347 4635
rect 5347 4610 5381 4635
rect 5381 4610 5388 4635
rect 5336 4583 5388 4610
rect 5468 4583 5520 4635
rect 5600 4583 5652 4635
rect 5732 4583 5784 4635
rect 5864 4583 5916 4635
rect 5996 4583 6048 4635
rect 6128 4583 6180 4635
rect 6260 4583 6312 4635
rect 6392 4583 6444 4635
rect 6524 4583 6576 4635
rect 6656 4583 6708 4635
rect 6788 4583 6840 4635
rect 6920 4583 6972 4635
rect 7052 4610 7059 4635
rect 7059 4610 7093 4635
rect 7093 4610 7104 4635
rect 7052 4583 7104 4610
rect 7184 4583 7236 4635
rect 7316 4583 7368 4635
rect 5204 4475 5256 4527
rect 5336 4494 5388 4527
rect 5336 4475 5347 4494
rect 5347 4475 5381 4494
rect 5381 4475 5388 4494
rect 5468 4475 5520 4527
rect 5600 4475 5652 4527
rect 5732 4475 5784 4527
rect 5864 4475 5916 4527
rect 5996 4475 6048 4527
rect 6128 4475 6180 4527
rect 6260 4475 6312 4527
rect 6392 4475 6444 4527
rect 6524 4475 6576 4527
rect 6656 4475 6708 4527
rect 6788 4475 6840 4527
rect 6920 4475 6972 4527
rect 7052 4494 7104 4527
rect 7052 4475 7059 4494
rect 7059 4475 7093 4494
rect 7093 4475 7104 4494
rect 7184 4475 7236 4527
rect 7316 4475 7368 4527
rect 5204 4367 5256 4419
rect 5336 4385 5347 4419
rect 5347 4385 5381 4419
rect 5381 4385 5388 4419
rect 5336 4367 5388 4385
rect 5468 4367 5520 4419
rect 5600 4367 5652 4419
rect 5732 4367 5784 4419
rect 5864 4367 5916 4419
rect 5996 4367 6048 4419
rect 6128 4367 6180 4419
rect 6260 4367 6312 4419
rect 6392 4367 6444 4419
rect 6524 4367 6576 4419
rect 6656 4367 6708 4419
rect 6788 4367 6840 4419
rect 6920 4367 6972 4419
rect 7052 4385 7059 4419
rect 7059 4385 7093 4419
rect 7093 4385 7104 4419
rect 7052 4367 7104 4385
rect 7184 4367 7236 4419
rect 7316 4367 7368 4419
rect 5204 4259 5256 4311
rect 5336 4310 5347 4311
rect 5347 4310 5381 4311
rect 5381 4310 5388 4311
rect 5336 4269 5388 4310
rect 5336 4259 5347 4269
rect 5347 4259 5381 4269
rect 5381 4259 5388 4269
rect 5468 4259 5520 4311
rect 5600 4259 5652 4311
rect 5732 4259 5784 4311
rect 5864 4259 5916 4311
rect 5996 4259 6048 4311
rect 6128 4259 6180 4311
rect 6260 4259 6312 4311
rect 6392 4259 6444 4311
rect 6524 4259 6576 4311
rect 6656 4259 6708 4311
rect 6788 4259 6840 4311
rect 6920 4259 6972 4311
rect 7052 4310 7059 4311
rect 7059 4310 7093 4311
rect 7093 4310 7104 4311
rect 7052 4269 7104 4310
rect 7052 4259 7059 4269
rect 7059 4259 7093 4269
rect 7093 4259 7104 4269
rect 7184 4259 7236 4311
rect 7316 4259 7368 4311
rect 5204 4151 5256 4203
rect 5336 4193 5388 4203
rect 5336 4159 5347 4193
rect 5347 4159 5381 4193
rect 5381 4159 5388 4193
rect 5336 4151 5388 4159
rect 5468 4151 5520 4203
rect 5600 4151 5652 4203
rect 5732 4151 5784 4203
rect 5864 4151 5916 4203
rect 5996 4151 6048 4203
rect 6128 4151 6180 4203
rect 6260 4151 6312 4203
rect 6392 4151 6444 4203
rect 6524 4151 6576 4203
rect 6656 4151 6708 4203
rect 6788 4151 6840 4203
rect 6920 4151 6972 4203
rect 7052 4193 7104 4203
rect 7052 4159 7059 4193
rect 7059 4159 7093 4193
rect 7093 4159 7104 4193
rect 7052 4151 7104 4159
rect 7184 4151 7236 4203
rect 7316 4151 7368 4203
rect 5204 3943 5256 3949
rect 5339 3943 5391 3949
rect 5474 3943 5526 3949
rect 5609 3943 5661 3949
rect 5744 3943 5796 3949
rect 5879 3943 5931 3949
rect 6014 3943 6066 3949
rect 6149 3943 6201 3949
rect 6284 3943 6336 3949
rect 6419 3943 6471 3949
rect 6553 3943 6605 3949
rect 6687 3943 6739 3949
rect 6821 3943 6873 3949
rect 6955 3943 7007 3949
rect 7089 3943 7141 3949
rect 7223 3943 7275 3949
rect 5204 3897 5256 3943
rect 5339 3897 5391 3943
rect 5474 3897 5526 3943
rect 5609 3897 5661 3943
rect 5744 3897 5796 3943
rect 5879 3897 5931 3943
rect 6014 3897 6066 3943
rect 6149 3897 6201 3943
rect 6284 3897 6336 3943
rect 6419 3897 6471 3943
rect 6553 3897 6605 3943
rect 6687 3897 6739 3943
rect 6821 3897 6873 3943
rect 6955 3897 7007 3943
rect 7089 3897 7141 3943
rect 7223 3897 7275 3943
rect 5204 3837 5256 3883
rect 5339 3837 5391 3883
rect 5474 3837 5526 3883
rect 5609 3837 5661 3883
rect 5744 3837 5796 3883
rect 5879 3837 5931 3883
rect 6014 3837 6066 3883
rect 6149 3837 6201 3883
rect 6284 3837 6336 3883
rect 6419 3837 6471 3883
rect 6553 3837 6605 3883
rect 6687 3837 6739 3883
rect 6821 3837 6873 3883
rect 6955 3837 7007 3883
rect 7089 3837 7141 3883
rect 7223 3837 7275 3883
rect 5204 3831 5256 3837
rect 5339 3831 5391 3837
rect 5474 3831 5526 3837
rect 5609 3831 5661 3837
rect 5744 3831 5796 3837
rect 5879 3831 5931 3837
rect 6014 3831 6066 3837
rect 6149 3831 6201 3837
rect 6284 3831 6336 3837
rect 6419 3831 6471 3837
rect 6553 3831 6605 3837
rect 6687 3831 6739 3837
rect 6821 3831 6873 3837
rect 6955 3831 7007 3837
rect 7089 3831 7141 3837
rect 7223 3831 7275 3837
rect 5204 3049 5256 3057
rect 5204 3015 5220 3049
rect 5220 3015 5254 3049
rect 5254 3015 5256 3049
rect 5204 3005 5256 3015
rect 5270 3049 5322 3057
rect 5336 3049 5388 3057
rect 5402 3049 5454 3057
rect 5468 3049 5520 3057
rect 5534 3049 5586 3057
rect 5599 3049 5651 3057
rect 5664 3049 5716 3057
rect 5729 3049 5781 3057
rect 5270 3015 5293 3049
rect 5293 3015 5322 3049
rect 5336 3015 5366 3049
rect 5366 3015 5388 3049
rect 5402 3015 5439 3049
rect 5439 3015 5454 3049
rect 5468 3015 5473 3049
rect 5473 3015 5511 3049
rect 5511 3015 5520 3049
rect 5534 3015 5545 3049
rect 5545 3015 5583 3049
rect 5583 3015 5586 3049
rect 5599 3015 5617 3049
rect 5617 3015 5651 3049
rect 5664 3015 5689 3049
rect 5689 3015 5716 3049
rect 5729 3015 5761 3049
rect 5761 3015 5781 3049
rect 5270 3005 5322 3015
rect 5336 3005 5388 3015
rect 5402 3005 5454 3015
rect 5468 3005 5520 3015
rect 5534 3005 5586 3015
rect 5599 3005 5651 3015
rect 5664 3005 5716 3015
rect 5729 3005 5781 3015
rect 5794 3049 5846 3057
rect 5794 3015 5799 3049
rect 5799 3015 5833 3049
rect 5833 3015 5846 3049
rect 5794 3005 5846 3015
rect 5859 3049 5911 3057
rect 5859 3015 5871 3049
rect 5871 3015 5905 3049
rect 5905 3015 5911 3049
rect 5859 3005 5911 3015
rect 5924 3049 5976 3057
rect 5989 3049 6041 3057
rect 6054 3049 6106 3057
rect 6119 3049 6171 3057
rect 6184 3049 6236 3057
rect 6249 3049 6301 3057
rect 6314 3049 6366 3057
rect 6379 3049 6431 3057
rect 5924 3015 5943 3049
rect 5943 3015 5976 3049
rect 5989 3015 6015 3049
rect 6015 3015 6041 3049
rect 6054 3015 6087 3049
rect 6087 3015 6106 3049
rect 6119 3015 6121 3049
rect 6121 3015 6159 3049
rect 6159 3015 6171 3049
rect 6184 3015 6193 3049
rect 6193 3015 6231 3049
rect 6231 3015 6236 3049
rect 6249 3015 6265 3049
rect 6265 3015 6301 3049
rect 6314 3015 6337 3049
rect 6337 3015 6366 3049
rect 6379 3015 6409 3049
rect 6409 3015 6431 3049
rect 5924 3005 5976 3015
rect 5989 3005 6041 3015
rect 6054 3005 6106 3015
rect 6119 3005 6171 3015
rect 6184 3005 6236 3015
rect 6249 3005 6301 3015
rect 6314 3005 6366 3015
rect 6379 3005 6431 3015
rect 6444 3049 6496 3057
rect 6444 3015 6447 3049
rect 6447 3015 6481 3049
rect 6481 3015 6496 3049
rect 6444 3005 6496 3015
rect 6509 3049 6561 3057
rect 6509 3015 6519 3049
rect 6519 3015 6553 3049
rect 6553 3015 6561 3049
rect 6509 3005 6561 3015
rect 6574 3049 6626 3057
rect 6574 3015 6591 3049
rect 6591 3015 6625 3049
rect 6625 3015 6626 3049
rect 6574 3005 6626 3015
rect 6639 3049 6691 3057
rect 6704 3049 6756 3057
rect 6769 3049 6821 3057
rect 6834 3049 6886 3057
rect 6899 3049 6951 3057
rect 6964 3049 7016 3057
rect 7029 3049 7081 3057
rect 6639 3015 6663 3049
rect 6663 3015 6691 3049
rect 6704 3015 6735 3049
rect 6735 3015 6756 3049
rect 6769 3015 6807 3049
rect 6807 3015 6821 3049
rect 6834 3015 6841 3049
rect 6841 3015 6879 3049
rect 6879 3015 6886 3049
rect 6899 3015 6913 3049
rect 6913 3015 6951 3049
rect 6964 3015 6985 3049
rect 6985 3015 7016 3049
rect 7029 3015 7057 3049
rect 7057 3015 7081 3049
rect 6639 3005 6691 3015
rect 6704 3005 6756 3015
rect 6769 3005 6821 3015
rect 6834 3005 6886 3015
rect 6899 3005 6951 3015
rect 6964 3005 7016 3015
rect 7029 3005 7081 3015
rect 7094 3049 7146 3057
rect 7094 3015 7095 3049
rect 7095 3015 7129 3049
rect 7129 3015 7146 3049
rect 7094 3005 7146 3015
rect 7159 3049 7211 3057
rect 7159 3015 7167 3049
rect 7167 3015 7201 3049
rect 7201 3015 7211 3049
rect 7159 3005 7211 3015
rect 7224 3049 7276 3057
rect 7224 3015 7239 3049
rect 7239 3015 7273 3049
rect 7273 3015 7276 3049
rect 7224 3005 7276 3015
rect 7289 3049 7341 3057
rect 7354 3049 7406 3057
rect 7419 3049 7471 3057
rect 7484 3049 7536 3057
rect 7289 3015 7311 3049
rect 7311 3015 7341 3049
rect 7354 3015 7383 3049
rect 7383 3015 7406 3049
rect 7419 3015 7455 3049
rect 7455 3015 7471 3049
rect 7484 3015 7489 3049
rect 7489 3015 7527 3049
rect 7527 3015 7536 3049
rect 7289 3005 7341 3015
rect 7354 3005 7406 3015
rect 7419 3005 7471 3015
rect 7484 3005 7536 3015
rect 5204 2971 5256 2989
rect 5204 2937 5220 2971
rect 5220 2937 5254 2971
rect 5254 2937 5256 2971
rect 5270 2971 5322 2989
rect 5336 2971 5388 2989
rect 5402 2971 5454 2989
rect 5468 2971 5520 2989
rect 5534 2971 5586 2989
rect 5599 2971 5651 2989
rect 5664 2971 5716 2989
rect 5729 2971 5781 2989
rect 5270 2937 5293 2971
rect 5293 2937 5322 2971
rect 5336 2937 5366 2971
rect 5366 2937 5388 2971
rect 5402 2937 5439 2971
rect 5439 2937 5454 2971
rect 5468 2937 5473 2971
rect 5473 2937 5511 2971
rect 5511 2937 5520 2971
rect 5534 2937 5545 2971
rect 5545 2937 5583 2971
rect 5583 2937 5586 2971
rect 5599 2937 5617 2971
rect 5617 2937 5651 2971
rect 5664 2937 5689 2971
rect 5689 2937 5716 2971
rect 5729 2937 5761 2971
rect 5761 2937 5781 2971
rect 5794 2971 5846 2989
rect 5794 2937 5799 2971
rect 5799 2937 5833 2971
rect 5833 2937 5846 2971
rect 5859 2971 5911 2989
rect 5859 2937 5871 2971
rect 5871 2937 5905 2971
rect 5905 2937 5911 2971
rect 5924 2971 5976 2989
rect 5989 2971 6041 2989
rect 6054 2971 6106 2989
rect 6119 2971 6171 2989
rect 6184 2971 6236 2989
rect 6249 2971 6301 2989
rect 6314 2971 6366 2989
rect 6379 2971 6431 2989
rect 5924 2937 5943 2971
rect 5943 2937 5976 2971
rect 5989 2937 6015 2971
rect 6015 2937 6041 2971
rect 6054 2937 6087 2971
rect 6087 2937 6106 2971
rect 6119 2937 6121 2971
rect 6121 2937 6159 2971
rect 6159 2937 6171 2971
rect 6184 2937 6193 2971
rect 6193 2937 6231 2971
rect 6231 2937 6236 2971
rect 6249 2937 6265 2971
rect 6265 2937 6301 2971
rect 6314 2937 6337 2971
rect 6337 2937 6366 2971
rect 6379 2937 6409 2971
rect 6409 2937 6431 2971
rect 6444 2971 6496 2989
rect 6444 2937 6447 2971
rect 6447 2937 6481 2971
rect 6481 2937 6496 2971
rect 6509 2971 6561 2989
rect 6509 2937 6519 2971
rect 6519 2937 6553 2971
rect 6553 2937 6561 2971
rect 6574 2971 6626 2989
rect 6574 2937 6591 2971
rect 6591 2937 6625 2971
rect 6625 2937 6626 2971
rect 6639 2971 6691 2989
rect 6704 2971 6756 2989
rect 6769 2971 6821 2989
rect 6834 2971 6886 2989
rect 6899 2971 6951 2989
rect 6964 2971 7016 2989
rect 7029 2971 7081 2989
rect 6639 2937 6663 2971
rect 6663 2937 6691 2971
rect 6704 2937 6735 2971
rect 6735 2937 6756 2971
rect 6769 2937 6807 2971
rect 6807 2937 6821 2971
rect 6834 2937 6841 2971
rect 6841 2937 6879 2971
rect 6879 2937 6886 2971
rect 6899 2937 6913 2971
rect 6913 2937 6951 2971
rect 6964 2937 6985 2971
rect 6985 2937 7016 2971
rect 7029 2937 7057 2971
rect 7057 2937 7081 2971
rect 7094 2971 7146 2989
rect 7094 2937 7095 2971
rect 7095 2937 7129 2971
rect 7129 2937 7146 2971
rect 7159 2971 7211 2989
rect 7159 2937 7167 2971
rect 7167 2937 7201 2971
rect 7201 2937 7211 2971
rect 7224 2971 7276 2989
rect 7224 2937 7239 2971
rect 7239 2937 7273 2971
rect 7273 2937 7276 2971
rect 7289 2971 7341 2989
rect 7354 2971 7406 2989
rect 7419 2971 7471 2989
rect 7484 2971 7536 2989
rect 7289 2937 7311 2971
rect 7311 2937 7341 2971
rect 7354 2937 7383 2971
rect 7383 2937 7406 2971
rect 7419 2937 7455 2971
rect 7455 2937 7471 2971
rect 7484 2937 7489 2971
rect 7489 2937 7527 2971
rect 7527 2937 7536 2971
rect 5204 2893 5256 2921
rect 5204 2869 5220 2893
rect 5220 2869 5254 2893
rect 5254 2869 5256 2893
rect 5270 2893 5322 2921
rect 5336 2893 5388 2921
rect 5402 2893 5454 2921
rect 5468 2893 5520 2921
rect 5534 2893 5586 2921
rect 5599 2893 5651 2921
rect 5664 2893 5716 2921
rect 5729 2893 5781 2921
rect 5270 2869 5293 2893
rect 5293 2869 5322 2893
rect 5336 2869 5366 2893
rect 5366 2869 5388 2893
rect 5402 2869 5439 2893
rect 5439 2869 5454 2893
rect 5468 2869 5473 2893
rect 5473 2869 5511 2893
rect 5511 2869 5520 2893
rect 5534 2869 5545 2893
rect 5545 2869 5583 2893
rect 5583 2869 5586 2893
rect 5599 2869 5617 2893
rect 5617 2869 5651 2893
rect 5664 2869 5689 2893
rect 5689 2869 5716 2893
rect 5729 2869 5761 2893
rect 5761 2869 5781 2893
rect 5794 2893 5846 2921
rect 5794 2869 5799 2893
rect 5799 2869 5833 2893
rect 5833 2869 5846 2893
rect 5859 2893 5911 2921
rect 5859 2869 5871 2893
rect 5871 2869 5905 2893
rect 5905 2869 5911 2893
rect 5924 2893 5976 2921
rect 5989 2893 6041 2921
rect 6054 2893 6106 2921
rect 6119 2893 6171 2921
rect 6184 2893 6236 2921
rect 6249 2893 6301 2921
rect 6314 2893 6366 2921
rect 6379 2893 6431 2921
rect 5924 2869 5943 2893
rect 5943 2869 5976 2893
rect 5989 2869 6015 2893
rect 6015 2869 6041 2893
rect 6054 2869 6087 2893
rect 6087 2869 6106 2893
rect 6119 2869 6121 2893
rect 6121 2869 6159 2893
rect 6159 2869 6171 2893
rect 6184 2869 6193 2893
rect 6193 2869 6231 2893
rect 6231 2869 6236 2893
rect 6249 2869 6265 2893
rect 6265 2869 6301 2893
rect 6314 2869 6337 2893
rect 6337 2869 6366 2893
rect 6379 2869 6409 2893
rect 6409 2869 6431 2893
rect 6444 2893 6496 2921
rect 6444 2869 6447 2893
rect 6447 2869 6481 2893
rect 6481 2869 6496 2893
rect 6509 2893 6561 2921
rect 6509 2869 6519 2893
rect 6519 2869 6553 2893
rect 6553 2869 6561 2893
rect 6574 2893 6626 2921
rect 6574 2869 6591 2893
rect 6591 2869 6625 2893
rect 6625 2869 6626 2893
rect 6639 2893 6691 2921
rect 6704 2893 6756 2921
rect 6769 2893 6821 2921
rect 6834 2893 6886 2921
rect 6899 2893 6951 2921
rect 6964 2893 7016 2921
rect 7029 2893 7081 2921
rect 6639 2869 6663 2893
rect 6663 2869 6691 2893
rect 6704 2869 6735 2893
rect 6735 2869 6756 2893
rect 6769 2869 6807 2893
rect 6807 2869 6821 2893
rect 6834 2869 6841 2893
rect 6841 2869 6879 2893
rect 6879 2869 6886 2893
rect 6899 2869 6913 2893
rect 6913 2869 6951 2893
rect 6964 2869 6985 2893
rect 6985 2869 7016 2893
rect 7029 2869 7057 2893
rect 7057 2869 7081 2893
rect 7094 2893 7146 2921
rect 7094 2869 7095 2893
rect 7095 2869 7129 2893
rect 7129 2869 7146 2893
rect 7159 2893 7211 2921
rect 7159 2869 7167 2893
rect 7167 2869 7201 2893
rect 7201 2869 7211 2893
rect 7224 2893 7276 2921
rect 7224 2869 7239 2893
rect 7239 2869 7273 2893
rect 7273 2869 7276 2893
rect 7289 2893 7341 2921
rect 7354 2893 7406 2921
rect 7419 2893 7471 2921
rect 7484 2893 7536 2921
rect 7289 2869 7311 2893
rect 7311 2869 7341 2893
rect 7354 2869 7383 2893
rect 7383 2869 7406 2893
rect 7419 2869 7455 2893
rect 7455 2869 7471 2893
rect 7484 2869 7489 2893
rect 7489 2869 7527 2893
rect 7527 2869 7536 2893
rect 5204 2815 5256 2853
rect 5204 2801 5220 2815
rect 5220 2801 5254 2815
rect 5254 2801 5256 2815
rect 5270 2815 5322 2853
rect 5336 2815 5388 2853
rect 5402 2815 5454 2853
rect 5468 2815 5520 2853
rect 5534 2815 5586 2853
rect 5599 2815 5651 2853
rect 5664 2815 5716 2853
rect 5729 2815 5781 2853
rect 5270 2801 5293 2815
rect 5293 2801 5322 2815
rect 5336 2801 5366 2815
rect 5366 2801 5388 2815
rect 5402 2801 5439 2815
rect 5439 2801 5454 2815
rect 5468 2801 5473 2815
rect 5473 2801 5511 2815
rect 5511 2801 5520 2815
rect 5534 2801 5545 2815
rect 5545 2801 5583 2815
rect 5583 2801 5586 2815
rect 5599 2801 5617 2815
rect 5617 2801 5651 2815
rect 5664 2801 5689 2815
rect 5689 2801 5716 2815
rect 5729 2801 5761 2815
rect 5761 2801 5781 2815
rect 5794 2815 5846 2853
rect 5794 2801 5799 2815
rect 5799 2801 5833 2815
rect 5833 2801 5846 2815
rect 5859 2815 5911 2853
rect 5859 2801 5871 2815
rect 5871 2801 5905 2815
rect 5905 2801 5911 2815
rect 5924 2815 5976 2853
rect 5989 2815 6041 2853
rect 6054 2815 6106 2853
rect 6119 2815 6171 2853
rect 6184 2815 6236 2853
rect 6249 2815 6301 2853
rect 6314 2815 6366 2853
rect 6379 2815 6431 2853
rect 5924 2801 5943 2815
rect 5943 2801 5976 2815
rect 5989 2801 6015 2815
rect 6015 2801 6041 2815
rect 6054 2801 6087 2815
rect 6087 2801 6106 2815
rect 6119 2801 6121 2815
rect 6121 2801 6159 2815
rect 6159 2801 6171 2815
rect 6184 2801 6193 2815
rect 6193 2801 6231 2815
rect 6231 2801 6236 2815
rect 6249 2801 6265 2815
rect 6265 2801 6301 2815
rect 6314 2801 6337 2815
rect 6337 2801 6366 2815
rect 6379 2801 6409 2815
rect 6409 2801 6431 2815
rect 6444 2815 6496 2853
rect 6444 2801 6447 2815
rect 6447 2801 6481 2815
rect 6481 2801 6496 2815
rect 6509 2815 6561 2853
rect 6509 2801 6519 2815
rect 6519 2801 6553 2815
rect 6553 2801 6561 2815
rect 6574 2815 6626 2853
rect 6574 2801 6591 2815
rect 6591 2801 6625 2815
rect 6625 2801 6626 2815
rect 6639 2815 6691 2853
rect 6704 2815 6756 2853
rect 6769 2815 6821 2853
rect 6834 2815 6886 2853
rect 6899 2815 6951 2853
rect 6964 2815 7016 2853
rect 7029 2815 7081 2853
rect 6639 2801 6663 2815
rect 6663 2801 6691 2815
rect 6704 2801 6735 2815
rect 6735 2801 6756 2815
rect 6769 2801 6807 2815
rect 6807 2801 6821 2815
rect 6834 2801 6841 2815
rect 6841 2801 6879 2815
rect 6879 2801 6886 2815
rect 6899 2801 6913 2815
rect 6913 2801 6951 2815
rect 6964 2801 6985 2815
rect 6985 2801 7016 2815
rect 7029 2801 7057 2815
rect 7057 2801 7081 2815
rect 7094 2815 7146 2853
rect 7094 2801 7095 2815
rect 7095 2801 7129 2815
rect 7129 2801 7146 2815
rect 7159 2815 7211 2853
rect 7159 2801 7167 2815
rect 7167 2801 7201 2815
rect 7201 2801 7211 2815
rect 7224 2815 7276 2853
rect 7224 2801 7239 2815
rect 7239 2801 7273 2815
rect 7273 2801 7276 2815
rect 7289 2815 7341 2853
rect 7354 2815 7406 2853
rect 7419 2815 7471 2853
rect 7484 2815 7536 2853
rect 7289 2801 7311 2815
rect 7311 2801 7341 2815
rect 7354 2801 7383 2815
rect 7383 2801 7406 2815
rect 7419 2801 7455 2815
rect 7455 2801 7471 2815
rect 7484 2801 7489 2815
rect 7489 2801 7527 2815
rect 7527 2801 7536 2815
rect 5204 2781 5220 2785
rect 5220 2781 5254 2785
rect 5254 2781 5256 2785
rect 5204 2737 5256 2781
rect 5204 2733 5220 2737
rect 5220 2733 5254 2737
rect 5254 2733 5256 2737
rect 5270 2781 5293 2785
rect 5293 2781 5322 2785
rect 5336 2781 5366 2785
rect 5366 2781 5388 2785
rect 5402 2781 5439 2785
rect 5439 2781 5454 2785
rect 5468 2781 5473 2785
rect 5473 2781 5511 2785
rect 5511 2781 5520 2785
rect 5534 2781 5545 2785
rect 5545 2781 5583 2785
rect 5583 2781 5586 2785
rect 5599 2781 5617 2785
rect 5617 2781 5651 2785
rect 5664 2781 5689 2785
rect 5689 2781 5716 2785
rect 5729 2781 5761 2785
rect 5761 2781 5781 2785
rect 5270 2737 5322 2781
rect 5336 2737 5388 2781
rect 5402 2737 5454 2781
rect 5468 2737 5520 2781
rect 5534 2737 5586 2781
rect 5599 2737 5651 2781
rect 5664 2737 5716 2781
rect 5729 2737 5781 2781
rect 5270 2733 5293 2737
rect 5293 2733 5322 2737
rect 5336 2733 5366 2737
rect 5366 2733 5388 2737
rect 5402 2733 5439 2737
rect 5439 2733 5454 2737
rect 5468 2733 5473 2737
rect 5473 2733 5511 2737
rect 5511 2733 5520 2737
rect 5534 2733 5545 2737
rect 5545 2733 5583 2737
rect 5583 2733 5586 2737
rect 5599 2733 5617 2737
rect 5617 2733 5651 2737
rect 5664 2733 5689 2737
rect 5689 2733 5716 2737
rect 5729 2733 5761 2737
rect 5761 2733 5781 2737
rect 5794 2781 5799 2785
rect 5799 2781 5833 2785
rect 5833 2781 5846 2785
rect 5794 2737 5846 2781
rect 5794 2733 5799 2737
rect 5799 2733 5833 2737
rect 5833 2733 5846 2737
rect 5859 2781 5871 2785
rect 5871 2781 5905 2785
rect 5905 2781 5911 2785
rect 5859 2737 5911 2781
rect 5859 2733 5871 2737
rect 5871 2733 5905 2737
rect 5905 2733 5911 2737
rect 5924 2781 5943 2785
rect 5943 2781 5976 2785
rect 5989 2781 6015 2785
rect 6015 2781 6041 2785
rect 6054 2781 6087 2785
rect 6087 2781 6106 2785
rect 6119 2781 6121 2785
rect 6121 2781 6159 2785
rect 6159 2781 6171 2785
rect 6184 2781 6193 2785
rect 6193 2781 6231 2785
rect 6231 2781 6236 2785
rect 6249 2781 6265 2785
rect 6265 2781 6301 2785
rect 6314 2781 6337 2785
rect 6337 2781 6366 2785
rect 6379 2781 6409 2785
rect 6409 2781 6431 2785
rect 5924 2737 5976 2781
rect 5989 2737 6041 2781
rect 6054 2737 6106 2781
rect 6119 2737 6171 2781
rect 6184 2737 6236 2781
rect 6249 2737 6301 2781
rect 6314 2737 6366 2781
rect 6379 2737 6431 2781
rect 5924 2733 5943 2737
rect 5943 2733 5976 2737
rect 5989 2733 6015 2737
rect 6015 2733 6041 2737
rect 6054 2733 6087 2737
rect 6087 2733 6106 2737
rect 6119 2733 6121 2737
rect 6121 2733 6159 2737
rect 6159 2733 6171 2737
rect 6184 2733 6193 2737
rect 6193 2733 6231 2737
rect 6231 2733 6236 2737
rect 6249 2733 6265 2737
rect 6265 2733 6301 2737
rect 6314 2733 6337 2737
rect 6337 2733 6366 2737
rect 6379 2733 6409 2737
rect 6409 2733 6431 2737
rect 6444 2781 6447 2785
rect 6447 2781 6481 2785
rect 6481 2781 6496 2785
rect 6444 2737 6496 2781
rect 6444 2733 6447 2737
rect 6447 2733 6481 2737
rect 6481 2733 6496 2737
rect 6509 2781 6519 2785
rect 6519 2781 6553 2785
rect 6553 2781 6561 2785
rect 6509 2737 6561 2781
rect 6509 2733 6519 2737
rect 6519 2733 6553 2737
rect 6553 2733 6561 2737
rect 6574 2781 6591 2785
rect 6591 2781 6625 2785
rect 6625 2781 6626 2785
rect 6574 2737 6626 2781
rect 6574 2733 6591 2737
rect 6591 2733 6625 2737
rect 6625 2733 6626 2737
rect 6639 2781 6663 2785
rect 6663 2781 6691 2785
rect 6704 2781 6735 2785
rect 6735 2781 6756 2785
rect 6769 2781 6807 2785
rect 6807 2781 6821 2785
rect 6834 2781 6841 2785
rect 6841 2781 6879 2785
rect 6879 2781 6886 2785
rect 6899 2781 6913 2785
rect 6913 2781 6951 2785
rect 6964 2781 6985 2785
rect 6985 2781 7016 2785
rect 7029 2781 7057 2785
rect 7057 2781 7081 2785
rect 6639 2737 6691 2781
rect 6704 2737 6756 2781
rect 6769 2737 6821 2781
rect 6834 2737 6886 2781
rect 6899 2737 6951 2781
rect 6964 2737 7016 2781
rect 7029 2737 7081 2781
rect 6639 2733 6663 2737
rect 6663 2733 6691 2737
rect 6704 2733 6735 2737
rect 6735 2733 6756 2737
rect 6769 2733 6807 2737
rect 6807 2733 6821 2737
rect 6834 2733 6841 2737
rect 6841 2733 6879 2737
rect 6879 2733 6886 2737
rect 6899 2733 6913 2737
rect 6913 2733 6951 2737
rect 6964 2733 6985 2737
rect 6985 2733 7016 2737
rect 7029 2733 7057 2737
rect 7057 2733 7081 2737
rect 7094 2781 7095 2785
rect 7095 2781 7129 2785
rect 7129 2781 7146 2785
rect 7094 2737 7146 2781
rect 7094 2733 7095 2737
rect 7095 2733 7129 2737
rect 7129 2733 7146 2737
rect 7159 2781 7167 2785
rect 7167 2781 7201 2785
rect 7201 2781 7211 2785
rect 7159 2737 7211 2781
rect 7159 2733 7167 2737
rect 7167 2733 7201 2737
rect 7201 2733 7211 2737
rect 7224 2781 7239 2785
rect 7239 2781 7273 2785
rect 7273 2781 7276 2785
rect 7224 2737 7276 2781
rect 7224 2733 7239 2737
rect 7239 2733 7273 2737
rect 7273 2733 7276 2737
rect 7289 2781 7311 2785
rect 7311 2781 7341 2785
rect 7354 2781 7383 2785
rect 7383 2781 7406 2785
rect 7419 2781 7455 2785
rect 7455 2781 7471 2785
rect 7484 2781 7489 2785
rect 7489 2781 7527 2785
rect 7527 2781 7536 2785
rect 7289 2737 7341 2781
rect 7354 2737 7406 2781
rect 7419 2737 7471 2781
rect 7484 2737 7536 2781
rect 7289 2733 7311 2737
rect 7311 2733 7341 2737
rect 7354 2733 7383 2737
rect 7383 2733 7406 2737
rect 7419 2733 7455 2737
rect 7455 2733 7471 2737
rect 7484 2733 7489 2737
rect 7489 2733 7527 2737
rect 7527 2733 7536 2737
rect 5204 2703 5220 2717
rect 5220 2703 5254 2717
rect 5254 2703 5256 2717
rect 5204 2665 5256 2703
rect 5270 2703 5293 2717
rect 5293 2703 5322 2717
rect 5336 2703 5366 2717
rect 5366 2703 5388 2717
rect 5402 2703 5439 2717
rect 5439 2703 5454 2717
rect 5468 2703 5473 2717
rect 5473 2703 5511 2717
rect 5511 2703 5520 2717
rect 5534 2703 5545 2717
rect 5545 2703 5583 2717
rect 5583 2703 5586 2717
rect 5599 2703 5617 2717
rect 5617 2703 5651 2717
rect 5664 2703 5689 2717
rect 5689 2703 5716 2717
rect 5729 2703 5761 2717
rect 5761 2703 5781 2717
rect 5270 2665 5322 2703
rect 5336 2665 5388 2703
rect 5402 2665 5454 2703
rect 5468 2665 5520 2703
rect 5534 2665 5586 2703
rect 5599 2665 5651 2703
rect 5664 2665 5716 2703
rect 5729 2665 5781 2703
rect 5794 2703 5799 2717
rect 5799 2703 5833 2717
rect 5833 2703 5846 2717
rect 5794 2665 5846 2703
rect 5859 2703 5871 2717
rect 5871 2703 5905 2717
rect 5905 2703 5911 2717
rect 5859 2665 5911 2703
rect 5924 2703 5943 2717
rect 5943 2703 5976 2717
rect 5989 2703 6015 2717
rect 6015 2703 6041 2717
rect 6054 2703 6087 2717
rect 6087 2703 6106 2717
rect 6119 2703 6121 2717
rect 6121 2703 6159 2717
rect 6159 2703 6171 2717
rect 6184 2703 6193 2717
rect 6193 2703 6231 2717
rect 6231 2703 6236 2717
rect 6249 2703 6265 2717
rect 6265 2703 6301 2717
rect 6314 2703 6337 2717
rect 6337 2703 6366 2717
rect 6379 2703 6409 2717
rect 6409 2703 6431 2717
rect 5924 2665 5976 2703
rect 5989 2665 6041 2703
rect 6054 2665 6106 2703
rect 6119 2665 6171 2703
rect 6184 2665 6236 2703
rect 6249 2665 6301 2703
rect 6314 2665 6366 2703
rect 6379 2665 6431 2703
rect 6444 2703 6447 2717
rect 6447 2703 6481 2717
rect 6481 2703 6496 2717
rect 6444 2665 6496 2703
rect 6509 2703 6519 2717
rect 6519 2703 6553 2717
rect 6553 2703 6561 2717
rect 6509 2665 6561 2703
rect 6574 2703 6591 2717
rect 6591 2703 6625 2717
rect 6625 2703 6626 2717
rect 6574 2665 6626 2703
rect 6639 2703 6663 2717
rect 6663 2703 6691 2717
rect 6704 2703 6735 2717
rect 6735 2703 6756 2717
rect 6769 2703 6807 2717
rect 6807 2703 6821 2717
rect 6834 2703 6841 2717
rect 6841 2703 6879 2717
rect 6879 2703 6886 2717
rect 6899 2703 6913 2717
rect 6913 2703 6951 2717
rect 6964 2703 6985 2717
rect 6985 2703 7016 2717
rect 7029 2703 7057 2717
rect 7057 2703 7081 2717
rect 6639 2665 6691 2703
rect 6704 2665 6756 2703
rect 6769 2665 6821 2703
rect 6834 2665 6886 2703
rect 6899 2665 6951 2703
rect 6964 2665 7016 2703
rect 7029 2665 7081 2703
rect 7094 2703 7095 2717
rect 7095 2703 7129 2717
rect 7129 2703 7146 2717
rect 7094 2665 7146 2703
rect 7159 2703 7167 2717
rect 7167 2703 7201 2717
rect 7201 2703 7211 2717
rect 7159 2665 7211 2703
rect 7224 2703 7239 2717
rect 7239 2703 7273 2717
rect 7273 2703 7276 2717
rect 7224 2665 7276 2703
rect 7289 2703 7311 2717
rect 7311 2703 7341 2717
rect 7354 2703 7383 2717
rect 7383 2703 7406 2717
rect 7419 2703 7455 2717
rect 7455 2703 7471 2717
rect 7484 2703 7489 2717
rect 7489 2703 7527 2717
rect 7527 2703 7536 2717
rect 7289 2665 7341 2703
rect 7354 2665 7406 2703
rect 7419 2665 7471 2703
rect 7484 2665 7536 2703
rect 5204 2625 5220 2649
rect 5220 2625 5254 2649
rect 5254 2625 5256 2649
rect 5204 2597 5256 2625
rect 5270 2625 5293 2649
rect 5293 2625 5322 2649
rect 5336 2625 5366 2649
rect 5366 2625 5388 2649
rect 5402 2625 5439 2649
rect 5439 2625 5454 2649
rect 5468 2625 5473 2649
rect 5473 2625 5511 2649
rect 5511 2625 5520 2649
rect 5534 2625 5545 2649
rect 5545 2625 5583 2649
rect 5583 2625 5586 2649
rect 5599 2625 5617 2649
rect 5617 2625 5651 2649
rect 5664 2625 5689 2649
rect 5689 2625 5716 2649
rect 5729 2625 5761 2649
rect 5761 2625 5781 2649
rect 5270 2597 5322 2625
rect 5336 2597 5388 2625
rect 5402 2597 5454 2625
rect 5468 2597 5520 2625
rect 5534 2597 5586 2625
rect 5599 2597 5651 2625
rect 5664 2597 5716 2625
rect 5729 2597 5781 2625
rect 5794 2625 5799 2649
rect 5799 2625 5833 2649
rect 5833 2625 5846 2649
rect 5794 2597 5846 2625
rect 5859 2625 5871 2649
rect 5871 2625 5905 2649
rect 5905 2625 5911 2649
rect 5859 2597 5911 2625
rect 5924 2625 5943 2649
rect 5943 2625 5976 2649
rect 5989 2625 6015 2649
rect 6015 2625 6041 2649
rect 6054 2625 6087 2649
rect 6087 2625 6106 2649
rect 6119 2625 6121 2649
rect 6121 2625 6159 2649
rect 6159 2625 6171 2649
rect 6184 2625 6193 2649
rect 6193 2625 6231 2649
rect 6231 2625 6236 2649
rect 6249 2625 6265 2649
rect 6265 2625 6301 2649
rect 6314 2625 6337 2649
rect 6337 2625 6366 2649
rect 6379 2625 6409 2649
rect 6409 2625 6431 2649
rect 5924 2597 5976 2625
rect 5989 2597 6041 2625
rect 6054 2597 6106 2625
rect 6119 2597 6171 2625
rect 6184 2597 6236 2625
rect 6249 2597 6301 2625
rect 6314 2597 6366 2625
rect 6379 2597 6431 2625
rect 6444 2625 6447 2649
rect 6447 2625 6481 2649
rect 6481 2625 6496 2649
rect 6444 2597 6496 2625
rect 6509 2625 6519 2649
rect 6519 2625 6553 2649
rect 6553 2625 6561 2649
rect 6509 2597 6561 2625
rect 6574 2625 6591 2649
rect 6591 2625 6625 2649
rect 6625 2625 6626 2649
rect 6574 2597 6626 2625
rect 6639 2625 6663 2649
rect 6663 2625 6691 2649
rect 6704 2625 6735 2649
rect 6735 2625 6756 2649
rect 6769 2625 6807 2649
rect 6807 2625 6821 2649
rect 6834 2625 6841 2649
rect 6841 2625 6879 2649
rect 6879 2625 6886 2649
rect 6899 2625 6913 2649
rect 6913 2625 6951 2649
rect 6964 2625 6985 2649
rect 6985 2625 7016 2649
rect 7029 2625 7057 2649
rect 7057 2625 7081 2649
rect 6639 2597 6691 2625
rect 6704 2597 6756 2625
rect 6769 2597 6821 2625
rect 6834 2597 6886 2625
rect 6899 2597 6951 2625
rect 6964 2597 7016 2625
rect 7029 2597 7081 2625
rect 7094 2625 7095 2649
rect 7095 2625 7129 2649
rect 7129 2625 7146 2649
rect 7094 2597 7146 2625
rect 7159 2625 7167 2649
rect 7167 2625 7201 2649
rect 7201 2625 7211 2649
rect 7159 2597 7211 2625
rect 7224 2625 7239 2649
rect 7239 2625 7273 2649
rect 7273 2625 7276 2649
rect 7224 2597 7276 2625
rect 7289 2625 7311 2649
rect 7311 2625 7341 2649
rect 7354 2625 7383 2649
rect 7383 2625 7406 2649
rect 7419 2625 7455 2649
rect 7455 2625 7471 2649
rect 7484 2625 7489 2649
rect 7489 2625 7527 2649
rect 7527 2625 7536 2649
rect 7289 2597 7341 2625
rect 7354 2597 7406 2625
rect 7419 2597 7471 2625
rect 7484 2597 7536 2625
rect 5204 2547 5220 2581
rect 5220 2547 5254 2581
rect 5254 2547 5256 2581
rect 5204 2529 5256 2547
rect 5270 2547 5293 2581
rect 5293 2547 5322 2581
rect 5336 2547 5366 2581
rect 5366 2547 5388 2581
rect 5402 2547 5439 2581
rect 5439 2547 5454 2581
rect 5468 2547 5473 2581
rect 5473 2547 5511 2581
rect 5511 2547 5520 2581
rect 5534 2547 5545 2581
rect 5545 2547 5583 2581
rect 5583 2547 5586 2581
rect 5599 2547 5617 2581
rect 5617 2547 5651 2581
rect 5664 2547 5689 2581
rect 5689 2547 5716 2581
rect 5729 2547 5761 2581
rect 5761 2547 5781 2581
rect 5270 2529 5322 2547
rect 5336 2529 5388 2547
rect 5402 2529 5454 2547
rect 5468 2529 5520 2547
rect 5534 2529 5586 2547
rect 5599 2529 5651 2547
rect 5664 2529 5716 2547
rect 5729 2529 5781 2547
rect 5794 2547 5799 2581
rect 5799 2547 5833 2581
rect 5833 2547 5846 2581
rect 5794 2529 5846 2547
rect 5859 2547 5871 2581
rect 5871 2547 5905 2581
rect 5905 2547 5911 2581
rect 5859 2529 5911 2547
rect 5924 2547 5943 2581
rect 5943 2547 5976 2581
rect 5989 2547 6015 2581
rect 6015 2547 6041 2581
rect 6054 2547 6087 2581
rect 6087 2547 6106 2581
rect 6119 2547 6121 2581
rect 6121 2547 6159 2581
rect 6159 2547 6171 2581
rect 6184 2547 6193 2581
rect 6193 2547 6231 2581
rect 6231 2547 6236 2581
rect 6249 2547 6265 2581
rect 6265 2547 6301 2581
rect 6314 2547 6337 2581
rect 6337 2547 6366 2581
rect 6379 2547 6409 2581
rect 6409 2547 6431 2581
rect 5924 2529 5976 2547
rect 5989 2529 6041 2547
rect 6054 2529 6106 2547
rect 6119 2529 6171 2547
rect 6184 2529 6236 2547
rect 6249 2529 6301 2547
rect 6314 2529 6366 2547
rect 6379 2529 6431 2547
rect 6444 2547 6447 2581
rect 6447 2547 6481 2581
rect 6481 2547 6496 2581
rect 6444 2529 6496 2547
rect 6509 2547 6519 2581
rect 6519 2547 6553 2581
rect 6553 2547 6561 2581
rect 6509 2529 6561 2547
rect 6574 2547 6591 2581
rect 6591 2547 6625 2581
rect 6625 2547 6626 2581
rect 6574 2529 6626 2547
rect 6639 2547 6663 2581
rect 6663 2547 6691 2581
rect 6704 2547 6735 2581
rect 6735 2547 6756 2581
rect 6769 2547 6807 2581
rect 6807 2547 6821 2581
rect 6834 2547 6841 2581
rect 6841 2547 6879 2581
rect 6879 2547 6886 2581
rect 6899 2547 6913 2581
rect 6913 2547 6951 2581
rect 6964 2547 6985 2581
rect 6985 2547 7016 2581
rect 7029 2547 7057 2581
rect 7057 2547 7081 2581
rect 6639 2529 6691 2547
rect 6704 2529 6756 2547
rect 6769 2529 6821 2547
rect 6834 2529 6886 2547
rect 6899 2529 6951 2547
rect 6964 2529 7016 2547
rect 7029 2529 7081 2547
rect 7094 2547 7095 2581
rect 7095 2547 7129 2581
rect 7129 2547 7146 2581
rect 7094 2529 7146 2547
rect 7159 2547 7167 2581
rect 7167 2547 7201 2581
rect 7201 2547 7211 2581
rect 7159 2529 7211 2547
rect 7224 2547 7239 2581
rect 7239 2547 7273 2581
rect 7273 2547 7276 2581
rect 7224 2529 7276 2547
rect 7289 2547 7311 2581
rect 7311 2547 7341 2581
rect 7354 2547 7383 2581
rect 7383 2547 7406 2581
rect 7419 2547 7455 2581
rect 7455 2547 7471 2581
rect 7484 2547 7489 2581
rect 7489 2547 7527 2581
rect 7527 2547 7536 2581
rect 7289 2529 7341 2547
rect 7354 2529 7406 2547
rect 7419 2529 7471 2547
rect 7484 2529 7536 2547
rect 5204 2503 5256 2513
rect 5204 2469 5220 2503
rect 5220 2469 5254 2503
rect 5254 2469 5256 2503
rect 5204 2461 5256 2469
rect 5270 2503 5322 2513
rect 5336 2503 5388 2513
rect 5402 2503 5454 2513
rect 5468 2503 5520 2513
rect 5534 2503 5586 2513
rect 5599 2503 5651 2513
rect 5664 2503 5716 2513
rect 5729 2503 5781 2513
rect 5270 2469 5293 2503
rect 5293 2469 5322 2503
rect 5336 2469 5366 2503
rect 5366 2469 5388 2503
rect 5402 2469 5439 2503
rect 5439 2469 5454 2503
rect 5468 2469 5473 2503
rect 5473 2469 5511 2503
rect 5511 2469 5520 2503
rect 5534 2469 5545 2503
rect 5545 2469 5583 2503
rect 5583 2469 5586 2503
rect 5599 2469 5617 2503
rect 5617 2469 5651 2503
rect 5664 2469 5689 2503
rect 5689 2469 5716 2503
rect 5729 2469 5761 2503
rect 5761 2469 5781 2503
rect 5270 2461 5322 2469
rect 5336 2461 5388 2469
rect 5402 2461 5454 2469
rect 5468 2461 5520 2469
rect 5534 2461 5586 2469
rect 5599 2461 5651 2469
rect 5664 2461 5716 2469
rect 5729 2461 5781 2469
rect 5794 2503 5846 2513
rect 5794 2469 5799 2503
rect 5799 2469 5833 2503
rect 5833 2469 5846 2503
rect 5794 2461 5846 2469
rect 5859 2503 5911 2513
rect 5859 2469 5871 2503
rect 5871 2469 5905 2503
rect 5905 2469 5911 2503
rect 5859 2461 5911 2469
rect 5924 2503 5976 2513
rect 5989 2503 6041 2513
rect 6054 2503 6106 2513
rect 6119 2503 6171 2513
rect 6184 2503 6236 2513
rect 6249 2503 6301 2513
rect 6314 2503 6366 2513
rect 6379 2503 6431 2513
rect 5924 2469 5943 2503
rect 5943 2469 5976 2503
rect 5989 2469 6015 2503
rect 6015 2469 6041 2503
rect 6054 2469 6087 2503
rect 6087 2469 6106 2503
rect 6119 2469 6121 2503
rect 6121 2469 6159 2503
rect 6159 2469 6171 2503
rect 6184 2469 6193 2503
rect 6193 2469 6231 2503
rect 6231 2469 6236 2503
rect 6249 2469 6265 2503
rect 6265 2469 6301 2503
rect 6314 2469 6337 2503
rect 6337 2469 6366 2503
rect 6379 2469 6409 2503
rect 6409 2469 6431 2503
rect 5924 2461 5976 2469
rect 5989 2461 6041 2469
rect 6054 2461 6106 2469
rect 6119 2461 6171 2469
rect 6184 2461 6236 2469
rect 6249 2461 6301 2469
rect 6314 2461 6366 2469
rect 6379 2461 6431 2469
rect 6444 2503 6496 2513
rect 6444 2469 6447 2503
rect 6447 2469 6481 2503
rect 6481 2469 6496 2503
rect 6444 2461 6496 2469
rect 6509 2503 6561 2513
rect 6509 2469 6519 2503
rect 6519 2469 6553 2503
rect 6553 2469 6561 2503
rect 6509 2461 6561 2469
rect 6574 2503 6626 2513
rect 6574 2469 6591 2503
rect 6591 2469 6625 2503
rect 6625 2469 6626 2503
rect 6574 2461 6626 2469
rect 6639 2503 6691 2513
rect 6704 2503 6756 2513
rect 6769 2503 6821 2513
rect 6834 2503 6886 2513
rect 6899 2503 6951 2513
rect 6964 2503 7016 2513
rect 7029 2503 7081 2513
rect 6639 2469 6663 2503
rect 6663 2469 6691 2503
rect 6704 2469 6735 2503
rect 6735 2469 6756 2503
rect 6769 2469 6807 2503
rect 6807 2469 6821 2503
rect 6834 2469 6841 2503
rect 6841 2469 6879 2503
rect 6879 2469 6886 2503
rect 6899 2469 6913 2503
rect 6913 2469 6951 2503
rect 6964 2469 6985 2503
rect 6985 2469 7016 2503
rect 7029 2469 7057 2503
rect 7057 2469 7081 2503
rect 6639 2461 6691 2469
rect 6704 2461 6756 2469
rect 6769 2461 6821 2469
rect 6834 2461 6886 2469
rect 6899 2461 6951 2469
rect 6964 2461 7016 2469
rect 7029 2461 7081 2469
rect 7094 2503 7146 2513
rect 7094 2469 7095 2503
rect 7095 2469 7129 2503
rect 7129 2469 7146 2503
rect 7094 2461 7146 2469
rect 7159 2503 7211 2513
rect 7159 2469 7167 2503
rect 7167 2469 7201 2503
rect 7201 2469 7211 2503
rect 7159 2461 7211 2469
rect 7224 2503 7276 2513
rect 7224 2469 7239 2503
rect 7239 2469 7273 2503
rect 7273 2469 7276 2503
rect 7224 2461 7276 2469
rect 7289 2503 7341 2513
rect 7354 2503 7406 2513
rect 7419 2503 7471 2513
rect 7484 2503 7536 2513
rect 7289 2469 7311 2503
rect 7311 2469 7341 2503
rect 7354 2469 7383 2503
rect 7383 2469 7406 2503
rect 7419 2469 7455 2503
rect 7455 2469 7471 2503
rect 7484 2469 7489 2503
rect 7489 2469 7527 2503
rect 7527 2469 7536 2503
rect 7289 2461 7341 2469
rect 7354 2461 7406 2469
rect 7419 2461 7471 2469
rect 7484 2461 7536 2469
rect 3192 2211 3244 2263
rect 3258 2211 3310 2263
rect 3324 2211 3376 2263
rect 3390 2211 3442 2263
rect 3456 2211 3508 2263
rect 3522 2211 3574 2263
rect 3588 2211 3640 2263
rect 3654 2211 3706 2263
rect 3720 2211 3772 2263
rect 3786 2211 3838 2263
rect 3852 2211 3904 2263
rect 3918 2211 3970 2263
rect 3984 2211 4036 2263
rect 4050 2211 4102 2263
rect 4116 2211 4168 2263
rect 4182 2211 4234 2263
rect 4248 2211 4300 2263
rect 4314 2211 4366 2263
rect 4380 2211 4432 2263
rect 4446 2211 4498 2263
rect 4512 2211 4564 2263
rect 4578 2211 4630 2263
rect 4644 2211 4696 2263
rect 4710 2211 4762 2263
rect 4776 2211 4828 2263
rect 4841 2211 4893 2263
rect 1977 2098 2029 2150
rect 2042 2098 2094 2150
rect 2107 2098 2159 2150
rect 3192 2145 3244 2197
rect 3258 2145 3310 2197
rect 3324 2145 3376 2197
rect 3390 2145 3442 2197
rect 3456 2145 3508 2197
rect 3522 2145 3574 2197
rect 3588 2145 3640 2197
rect 3654 2145 3706 2197
rect 3720 2145 3772 2197
rect 3786 2145 3838 2197
rect 3852 2145 3904 2197
rect 3918 2145 3970 2197
rect 3984 2145 4036 2197
rect 4050 2145 4102 2197
rect 4116 2145 4168 2197
rect 4182 2145 4234 2197
rect 4248 2145 4300 2197
rect 4314 2145 4366 2197
rect 4380 2145 4432 2197
rect 4446 2145 4498 2197
rect 4512 2145 4564 2197
rect 4578 2145 4630 2197
rect 4644 2145 4696 2197
rect 4710 2145 4762 2197
rect 4776 2145 4828 2197
rect 4841 2145 4893 2197
rect 3192 2079 3244 2131
rect 3258 2079 3310 2131
rect 3324 2079 3376 2131
rect 3390 2079 3442 2131
rect 3456 2079 3508 2131
rect 3522 2079 3574 2131
rect 3588 2079 3640 2131
rect 3654 2079 3706 2131
rect 3720 2079 3772 2131
rect 3786 2079 3838 2131
rect 3852 2079 3904 2131
rect 3918 2079 3970 2131
rect 3984 2079 4036 2131
rect 4050 2079 4102 2131
rect 4116 2079 4168 2131
rect 4182 2079 4234 2131
rect 4248 2079 4300 2131
rect 4314 2079 4366 2131
rect 4380 2079 4432 2131
rect 4446 2079 4498 2131
rect 4512 2079 4564 2131
rect 4578 2079 4630 2131
rect 4644 2079 4696 2131
rect 4710 2079 4762 2131
rect 4776 2079 4828 2131
rect 4841 2079 4893 2131
rect 3192 2016 3244 2065
rect 3192 2013 3202 2016
rect 3202 2013 3236 2016
rect 3236 2013 3244 2016
rect 3258 2016 3310 2065
rect 3258 2013 3275 2016
rect 3275 2013 3309 2016
rect 3309 2013 3310 2016
rect 3324 2016 3376 2065
rect 3390 2016 3442 2065
rect 3456 2016 3508 2065
rect 3522 2016 3574 2065
rect 3588 2016 3640 2065
rect 3654 2016 3706 2065
rect 3720 2016 3772 2065
rect 3786 2016 3838 2065
rect 3324 2013 3348 2016
rect 3348 2013 3376 2016
rect 3390 2013 3421 2016
rect 3421 2013 3442 2016
rect 3456 2013 3493 2016
rect 3493 2013 3508 2016
rect 3522 2013 3527 2016
rect 3527 2013 3565 2016
rect 3565 2013 3574 2016
rect 3588 2013 3599 2016
rect 3599 2013 3637 2016
rect 3637 2013 3640 2016
rect 3654 2013 3671 2016
rect 3671 2013 3706 2016
rect 3720 2013 3743 2016
rect 3743 2013 3772 2016
rect 3786 2013 3815 2016
rect 3815 2013 3838 2016
rect 3852 2016 3904 2065
rect 3852 2013 3853 2016
rect 3853 2013 3887 2016
rect 3887 2013 3904 2016
rect 3918 2016 3970 2065
rect 3918 2013 3925 2016
rect 3925 2013 3959 2016
rect 3959 2013 3970 2016
rect 3984 2016 4036 2065
rect 3984 2013 3997 2016
rect 3997 2013 4031 2016
rect 4031 2013 4036 2016
rect 4050 2016 4102 2065
rect 4116 2016 4168 2065
rect 4182 2016 4234 2065
rect 4248 2016 4300 2065
rect 4314 2016 4366 2065
rect 4380 2016 4432 2065
rect 4446 2016 4498 2065
rect 4512 2016 4564 2065
rect 4578 2016 4630 2065
rect 4050 2013 4069 2016
rect 4069 2013 4102 2016
rect 4116 2013 4141 2016
rect 4141 2013 4168 2016
rect 4182 2013 4213 2016
rect 4213 2013 4234 2016
rect 4248 2013 4285 2016
rect 4285 2013 4300 2016
rect 4314 2013 4319 2016
rect 4319 2013 4357 2016
rect 4357 2013 4366 2016
rect 4380 2013 4391 2016
rect 4391 2013 4429 2016
rect 4429 2013 4432 2016
rect 4446 2013 4463 2016
rect 4463 2013 4498 2016
rect 4512 2013 4535 2016
rect 4535 2013 4564 2016
rect 4578 2013 4607 2016
rect 4607 2013 4630 2016
rect 4644 2016 4696 2065
rect 4644 2013 4645 2016
rect 4645 2013 4679 2016
rect 4679 2013 4696 2016
rect 4710 2016 4762 2065
rect 4710 2013 4717 2016
rect 4717 2013 4751 2016
rect 4751 2013 4762 2016
rect 4776 2016 4828 2065
rect 4776 2013 4789 2016
rect 4789 2013 4823 2016
rect 4823 2013 4828 2016
rect 4841 2016 4893 2065
rect 4841 2013 4861 2016
rect 4861 2013 4893 2016
rect 3192 1982 3202 1999
rect 3202 1982 3236 1999
rect 3236 1982 3244 1999
rect 3192 1947 3244 1982
rect 3258 1982 3275 1999
rect 3275 1982 3309 1999
rect 3309 1982 3310 1999
rect 3258 1947 3310 1982
rect 3324 1982 3348 1999
rect 3348 1982 3376 1999
rect 3390 1982 3421 1999
rect 3421 1982 3442 1999
rect 3456 1982 3493 1999
rect 3493 1982 3508 1999
rect 3522 1982 3527 1999
rect 3527 1982 3565 1999
rect 3565 1982 3574 1999
rect 3588 1982 3599 1999
rect 3599 1982 3637 1999
rect 3637 1982 3640 1999
rect 3654 1982 3671 1999
rect 3671 1982 3706 1999
rect 3720 1982 3743 1999
rect 3743 1982 3772 1999
rect 3786 1982 3815 1999
rect 3815 1982 3838 1999
rect 3324 1947 3376 1982
rect 3390 1947 3442 1982
rect 3456 1947 3508 1982
rect 3522 1947 3574 1982
rect 3588 1947 3640 1982
rect 3654 1947 3706 1982
rect 3720 1947 3772 1982
rect 3786 1947 3838 1982
rect 3852 1982 3853 1999
rect 3853 1982 3887 1999
rect 3887 1982 3904 1999
rect 3852 1947 3904 1982
rect 3918 1982 3925 1999
rect 3925 1982 3959 1999
rect 3959 1982 3970 1999
rect 3918 1947 3970 1982
rect 3984 1982 3997 1999
rect 3997 1982 4031 1999
rect 4031 1982 4036 1999
rect 3984 1947 4036 1982
rect 4050 1982 4069 1999
rect 4069 1982 4102 1999
rect 4116 1982 4141 1999
rect 4141 1982 4168 1999
rect 4182 1982 4213 1999
rect 4213 1982 4234 1999
rect 4248 1982 4285 1999
rect 4285 1982 4300 1999
rect 4314 1982 4319 1999
rect 4319 1982 4357 1999
rect 4357 1982 4366 1999
rect 4380 1982 4391 1999
rect 4391 1982 4429 1999
rect 4429 1982 4432 1999
rect 4446 1982 4463 1999
rect 4463 1982 4498 1999
rect 4512 1982 4535 1999
rect 4535 1982 4564 1999
rect 4578 1982 4607 1999
rect 4607 1982 4630 1999
rect 4050 1947 4102 1982
rect 4116 1947 4168 1982
rect 4182 1947 4234 1982
rect 4248 1947 4300 1982
rect 4314 1947 4366 1982
rect 4380 1947 4432 1982
rect 4446 1947 4498 1982
rect 4512 1947 4564 1982
rect 4578 1947 4630 1982
rect 4644 1982 4645 1999
rect 4645 1982 4679 1999
rect 4679 1982 4696 1999
rect 4644 1947 4696 1982
rect 4710 1982 4717 1999
rect 4717 1982 4751 1999
rect 4751 1982 4762 1999
rect 4710 1947 4762 1982
rect 4776 1982 4789 1999
rect 4789 1982 4823 1999
rect 4823 1982 4828 1999
rect 4776 1947 4828 1982
rect 4841 1982 4861 1999
rect 4861 1982 4893 1999
rect 4841 1947 4893 1982
rect 3192 1917 3244 1933
rect 3192 1883 3207 1917
rect 3207 1883 3241 1917
rect 3241 1883 3244 1917
rect 3192 1881 3244 1883
rect 3258 1917 3310 1933
rect 3324 1917 3376 1933
rect 3258 1883 3281 1917
rect 3281 1883 3310 1917
rect 3324 1883 3355 1917
rect 3355 1883 3376 1917
rect 3258 1881 3310 1883
rect 3324 1881 3376 1883
rect 3390 1881 3442 1933
rect 3456 1881 3508 1933
rect 3522 1917 3574 1933
rect 3522 1883 3539 1917
rect 3539 1883 3573 1917
rect 3573 1883 3574 1917
rect 3522 1881 3574 1883
rect 3588 1917 3640 1933
rect 3654 1917 3706 1933
rect 3720 1917 3772 1933
rect 3786 1917 3838 1933
rect 3852 1917 3904 1933
rect 3918 1917 3970 1933
rect 3588 1883 3614 1917
rect 3614 1883 3640 1917
rect 3654 1883 3689 1917
rect 3689 1883 3706 1917
rect 3720 1883 3723 1917
rect 3723 1883 3764 1917
rect 3764 1883 3772 1917
rect 3786 1883 3798 1917
rect 3798 1883 3838 1917
rect 3852 1883 3873 1917
rect 3873 1883 3904 1917
rect 3918 1883 3948 1917
rect 3948 1883 3970 1917
rect 3588 1881 3640 1883
rect 3654 1881 3706 1883
rect 3720 1881 3772 1883
rect 3786 1881 3838 1883
rect 3852 1881 3904 1883
rect 3918 1881 3970 1883
rect 3984 1917 4036 1933
rect 3984 1883 3989 1917
rect 3989 1883 4023 1917
rect 4023 1883 4036 1917
rect 3984 1881 4036 1883
rect 4050 1917 4102 1933
rect 4050 1883 4064 1917
rect 4064 1883 4098 1917
rect 4098 1883 4102 1917
rect 4050 1881 4102 1883
rect 4116 1917 4168 1933
rect 4182 1917 4234 1933
rect 4248 1917 4300 1933
rect 4314 1917 4366 1933
rect 4380 1917 4432 1933
rect 4446 1917 4498 1933
rect 4116 1883 4139 1917
rect 4139 1883 4168 1917
rect 4182 1883 4214 1917
rect 4214 1883 4234 1917
rect 4248 1883 4289 1917
rect 4289 1883 4300 1917
rect 4314 1883 4323 1917
rect 4323 1883 4364 1917
rect 4364 1883 4366 1917
rect 4380 1883 4398 1917
rect 4398 1883 4432 1917
rect 4446 1883 4473 1917
rect 4473 1883 4498 1917
rect 4116 1881 4168 1883
rect 4182 1881 4234 1883
rect 4248 1881 4300 1883
rect 4314 1881 4366 1883
rect 4380 1881 4432 1883
rect 4446 1881 4498 1883
rect 4512 1917 4564 1933
rect 4512 1883 4514 1917
rect 4514 1883 4548 1917
rect 4548 1883 4564 1917
rect 4512 1881 4564 1883
rect 4578 1917 4630 1933
rect 4578 1883 4589 1917
rect 4589 1883 4623 1917
rect 4623 1883 4630 1917
rect 4578 1881 4630 1883
rect 4644 1917 4696 1933
rect 4710 1917 4762 1933
rect 4776 1917 4828 1933
rect 4841 1917 4893 1933
rect 4644 1883 4663 1917
rect 4663 1883 4696 1917
rect 4710 1883 4737 1917
rect 4737 1883 4762 1917
rect 4776 1883 4811 1917
rect 4811 1883 4828 1917
rect 4841 1883 4845 1917
rect 4845 1883 4885 1917
rect 4885 1883 4893 1917
rect 4644 1881 4696 1883
rect 4710 1881 4762 1883
rect 4776 1881 4828 1883
rect 4841 1881 4893 1883
rect 2798 1825 2850 1834
rect 2891 1825 2943 1834
rect 2983 1825 3035 1834
rect 2798 1791 2837 1825
rect 2837 1791 2850 1825
rect 2891 1791 2911 1825
rect 2911 1791 2943 1825
rect 2983 1791 2985 1825
rect 2985 1791 3019 1825
rect 3019 1791 3035 1825
rect 2798 1782 2850 1791
rect 2891 1782 2943 1791
rect 2983 1782 3035 1791
rect 2798 1641 2850 1650
rect 2891 1641 2943 1650
rect 2983 1641 3035 1650
rect 2798 1607 2837 1641
rect 2837 1607 2850 1641
rect 2891 1607 2911 1641
rect 2911 1607 2943 1641
rect 2983 1607 2985 1641
rect 2985 1607 3019 1641
rect 3019 1607 3035 1641
rect 2798 1598 2850 1607
rect 2891 1598 2943 1607
rect 2983 1598 3035 1607
rect 2798 1457 2850 1467
rect 2891 1457 2943 1467
rect 2983 1457 3035 1467
rect 2798 1423 2837 1457
rect 2837 1423 2850 1457
rect 2891 1423 2911 1457
rect 2911 1423 2943 1457
rect 2983 1423 2985 1457
rect 2985 1423 3019 1457
rect 3019 1423 3035 1457
rect 2798 1415 2850 1423
rect 2891 1415 2943 1423
rect 2983 1415 3035 1423
rect 2798 1273 2850 1282
rect 2891 1273 2943 1282
rect 2983 1273 3035 1282
rect 2798 1239 2837 1273
rect 2837 1239 2850 1273
rect 2891 1239 2911 1273
rect 2911 1239 2943 1273
rect 2983 1239 2985 1273
rect 2985 1239 3019 1273
rect 3019 1239 3035 1273
rect 2798 1230 2850 1239
rect 2891 1230 2943 1239
rect 2983 1230 3035 1239
rect 2798 1089 2850 1098
rect 2891 1089 2943 1098
rect 2983 1089 3035 1098
rect 2798 1055 2837 1089
rect 2837 1055 2850 1089
rect 2891 1055 2911 1089
rect 2911 1055 2943 1089
rect 2983 1055 2985 1089
rect 2985 1055 3019 1089
rect 3019 1055 3035 1089
rect 2798 1046 2850 1055
rect 2891 1046 2943 1055
rect 2983 1046 3035 1055
rect 6611 2235 6629 2242
rect 6629 2235 6663 2242
rect 6711 2235 6739 2242
rect 6739 2235 6763 2242
rect 6811 2235 6845 2242
rect 6845 2235 6863 2242
rect 6911 2235 6917 2242
rect 6917 2235 6955 2242
rect 6955 2235 6963 2242
rect 7011 2235 7027 2242
rect 7027 2235 7061 2242
rect 7061 2235 7063 2242
rect 7111 2235 7133 2242
rect 7133 2235 7163 2242
rect 7211 2235 7243 2242
rect 7243 2235 7263 2242
rect 7311 2235 7315 2242
rect 7315 2235 7349 2242
rect 7349 2235 7363 2242
rect 5628 2195 6320 2228
rect 6611 2195 6663 2235
rect 6711 2195 6763 2235
rect 6811 2195 6863 2235
rect 6911 2195 6963 2235
rect 7011 2195 7063 2235
rect 7111 2195 7163 2235
rect 7211 2195 7263 2235
rect 7311 2195 7363 2235
rect 5628 2161 5630 2195
rect 5630 2161 5664 2195
rect 5664 2161 5702 2195
rect 5702 2161 5736 2195
rect 5736 2161 5774 2195
rect 5774 2161 5808 2195
rect 5808 2161 5846 2195
rect 5846 2161 5880 2195
rect 5880 2161 5918 2195
rect 5918 2161 5952 2195
rect 5952 2161 5990 2195
rect 5990 2161 6024 2195
rect 6024 2161 6062 2195
rect 6062 2161 6096 2195
rect 6096 2161 6134 2195
rect 6134 2161 6168 2195
rect 6168 2161 6206 2195
rect 6206 2161 6240 2195
rect 6240 2161 6278 2195
rect 6278 2161 6312 2195
rect 6312 2161 6320 2195
rect 6611 2190 6629 2195
rect 6629 2190 6663 2195
rect 6711 2190 6739 2195
rect 6739 2190 6763 2195
rect 6811 2190 6845 2195
rect 6845 2190 6863 2195
rect 6911 2190 6917 2195
rect 6917 2190 6955 2195
rect 6955 2190 6963 2195
rect 7011 2190 7027 2195
rect 7027 2190 7061 2195
rect 7061 2190 7063 2195
rect 7111 2190 7133 2195
rect 7133 2190 7163 2195
rect 7211 2190 7243 2195
rect 7243 2190 7263 2195
rect 7311 2190 7315 2195
rect 7315 2190 7349 2195
rect 7349 2190 7363 2195
rect 5628 2121 6320 2161
rect 5628 2087 5630 2121
rect 5630 2087 5664 2121
rect 5664 2087 5702 2121
rect 5702 2087 5736 2121
rect 5736 2087 5774 2121
rect 5774 2087 5808 2121
rect 5808 2087 5846 2121
rect 5846 2087 5880 2121
rect 5880 2087 5918 2121
rect 5918 2087 5952 2121
rect 5952 2087 5990 2121
rect 5990 2087 6024 2121
rect 6024 2087 6062 2121
rect 6062 2087 6096 2121
rect 6096 2087 6134 2121
rect 6134 2087 6168 2121
rect 6168 2087 6206 2121
rect 6206 2087 6240 2121
rect 6240 2087 6278 2121
rect 6278 2087 6312 2121
rect 6312 2087 6320 2121
rect 6611 2087 6629 2108
rect 6629 2087 6663 2108
rect 6711 2087 6739 2108
rect 6739 2087 6763 2108
rect 6811 2087 6845 2108
rect 6845 2087 6863 2108
rect 6911 2087 6917 2108
rect 6917 2087 6955 2108
rect 6955 2087 6963 2108
rect 7011 2087 7027 2108
rect 7027 2087 7061 2108
rect 7061 2087 7063 2108
rect 7111 2087 7133 2108
rect 7133 2087 7163 2108
rect 7211 2087 7243 2108
rect 7243 2087 7263 2108
rect 7311 2087 7315 2108
rect 7315 2087 7349 2108
rect 7349 2087 7363 2108
rect 5628 2047 6320 2087
rect 6611 2056 6663 2087
rect 6711 2056 6763 2087
rect 6811 2056 6863 2087
rect 6911 2056 6963 2087
rect 7011 2056 7063 2087
rect 7111 2056 7163 2087
rect 7211 2056 7263 2087
rect 7311 2056 7363 2087
rect 5628 2013 5630 2047
rect 5630 2013 5664 2047
rect 5664 2013 5702 2047
rect 5702 2013 5736 2047
rect 5736 2013 5774 2047
rect 5774 2013 5808 2047
rect 5808 2013 5846 2047
rect 5846 2013 5880 2047
rect 5880 2013 5918 2047
rect 5918 2013 5952 2047
rect 5952 2013 5990 2047
rect 5990 2013 6024 2047
rect 6024 2013 6062 2047
rect 6062 2013 6096 2047
rect 6096 2013 6134 2047
rect 6134 2013 6168 2047
rect 6168 2013 6206 2047
rect 6206 2013 6240 2047
rect 6240 2013 6278 2047
rect 6278 2013 6312 2047
rect 6312 2013 6320 2047
rect 5628 1973 6320 2013
rect 5628 1939 5630 1973
rect 5630 1939 5664 1973
rect 5664 1939 5702 1973
rect 5702 1939 5736 1973
rect 5736 1939 5774 1973
rect 5774 1939 5808 1973
rect 5808 1939 5846 1973
rect 5846 1939 5880 1973
rect 5880 1939 5918 1973
rect 5918 1939 5952 1973
rect 5952 1939 5990 1973
rect 5990 1939 6024 1973
rect 6024 1939 6062 1973
rect 6062 1939 6096 1973
rect 6096 1939 6134 1973
rect 6134 1939 6168 1973
rect 6168 1939 6206 1973
rect 6206 1939 6240 1973
rect 6240 1939 6278 1973
rect 6278 1939 6312 1973
rect 6312 1939 6320 1973
rect 6611 1939 6629 1973
rect 6629 1939 6663 1973
rect 6711 1939 6739 1973
rect 6739 1939 6763 1973
rect 6811 1939 6845 1973
rect 6845 1939 6863 1973
rect 6911 1939 6917 1973
rect 6917 1939 6955 1973
rect 6955 1939 6963 1973
rect 7011 1939 7027 1973
rect 7027 1939 7061 1973
rect 7061 1939 7063 1973
rect 7111 1939 7133 1973
rect 7133 1939 7163 1973
rect 7211 1939 7243 1973
rect 7243 1939 7263 1973
rect 7311 1939 7315 1973
rect 7315 1939 7349 1973
rect 7349 1939 7363 1973
rect 5628 1899 6320 1939
rect 6611 1921 6663 1939
rect 6711 1921 6763 1939
rect 6811 1921 6863 1939
rect 6911 1921 6963 1939
rect 7011 1921 7063 1939
rect 7111 1921 7163 1939
rect 7211 1921 7263 1939
rect 7311 1921 7363 1939
rect 5628 1865 5630 1899
rect 5630 1865 5664 1899
rect 5664 1865 5702 1899
rect 5702 1865 5736 1899
rect 5736 1865 5774 1899
rect 5774 1865 5808 1899
rect 5808 1865 5846 1899
rect 5846 1865 5880 1899
rect 5880 1865 5918 1899
rect 5918 1865 5952 1899
rect 5952 1865 5990 1899
rect 5990 1865 6024 1899
rect 6024 1865 6062 1899
rect 6062 1865 6096 1899
rect 6096 1865 6134 1899
rect 6134 1865 6168 1899
rect 6168 1865 6206 1899
rect 6206 1865 6240 1899
rect 6240 1865 6278 1899
rect 6278 1865 6312 1899
rect 6312 1865 6320 1899
rect 5628 1825 6320 1865
rect 6611 1825 6663 1838
rect 6711 1825 6763 1838
rect 6811 1825 6863 1838
rect 6911 1825 6963 1838
rect 7011 1825 7063 1838
rect 7111 1825 7163 1838
rect 7211 1825 7263 1838
rect 7311 1825 7363 1838
rect 5628 1791 5630 1825
rect 5630 1791 5664 1825
rect 5664 1791 5702 1825
rect 5702 1791 5736 1825
rect 5736 1791 5774 1825
rect 5774 1791 5808 1825
rect 5808 1791 5846 1825
rect 5846 1791 5880 1825
rect 5880 1791 5918 1825
rect 5918 1791 5952 1825
rect 5952 1791 5990 1825
rect 5990 1791 6024 1825
rect 6024 1791 6062 1825
rect 6062 1791 6096 1825
rect 6096 1791 6134 1825
rect 6134 1791 6168 1825
rect 6168 1791 6206 1825
rect 6206 1791 6240 1825
rect 6240 1791 6278 1825
rect 6278 1791 6312 1825
rect 6312 1791 6320 1825
rect 6611 1791 6629 1825
rect 6629 1791 6663 1825
rect 6711 1791 6739 1825
rect 6739 1791 6763 1825
rect 6811 1791 6845 1825
rect 6845 1791 6863 1825
rect 6911 1791 6917 1825
rect 6917 1791 6955 1825
rect 6955 1791 6963 1825
rect 7011 1791 7027 1825
rect 7027 1791 7061 1825
rect 7061 1791 7063 1825
rect 7111 1791 7133 1825
rect 7133 1791 7163 1825
rect 7211 1791 7243 1825
rect 7243 1791 7263 1825
rect 7311 1791 7315 1825
rect 7315 1791 7349 1825
rect 7349 1791 7363 1825
rect 5628 1751 6320 1791
rect 6611 1786 6663 1791
rect 6711 1786 6763 1791
rect 6811 1786 6863 1791
rect 6911 1786 6963 1791
rect 7011 1786 7063 1791
rect 7111 1786 7163 1791
rect 7211 1786 7263 1791
rect 7311 1786 7363 1791
rect 5628 1717 5630 1751
rect 5630 1717 5664 1751
rect 5664 1717 5702 1751
rect 5702 1717 5736 1751
rect 5736 1717 5774 1751
rect 5774 1717 5808 1751
rect 5808 1717 5846 1751
rect 5846 1717 5880 1751
rect 5880 1717 5918 1751
rect 5918 1717 5952 1751
rect 5952 1717 5990 1751
rect 5990 1717 6024 1751
rect 6024 1717 6062 1751
rect 6062 1717 6096 1751
rect 6096 1717 6134 1751
rect 6134 1717 6168 1751
rect 6168 1717 6206 1751
rect 6206 1717 6240 1751
rect 6240 1717 6278 1751
rect 6278 1717 6312 1751
rect 6312 1717 6320 1751
rect 5628 1676 6320 1717
rect 6611 1676 6663 1703
rect 6711 1676 6763 1703
rect 6811 1676 6863 1703
rect 6911 1676 6963 1703
rect 7011 1676 7063 1703
rect 7111 1676 7163 1703
rect 7211 1676 7263 1703
rect 7311 1676 7363 1703
rect 5628 1642 5630 1676
rect 5630 1642 5664 1676
rect 5664 1642 5702 1676
rect 5702 1642 5736 1676
rect 5736 1642 5774 1676
rect 5774 1642 5808 1676
rect 5808 1642 5846 1676
rect 5846 1642 5880 1676
rect 5880 1642 5918 1676
rect 5918 1642 5952 1676
rect 5952 1642 5990 1676
rect 5990 1642 6024 1676
rect 6024 1642 6062 1676
rect 6062 1642 6096 1676
rect 6096 1642 6134 1676
rect 6134 1642 6168 1676
rect 6168 1642 6206 1676
rect 6206 1642 6240 1676
rect 6240 1642 6278 1676
rect 6278 1642 6312 1676
rect 6312 1642 6320 1676
rect 6611 1651 6629 1676
rect 6629 1651 6663 1676
rect 6711 1651 6739 1676
rect 6739 1651 6763 1676
rect 6811 1651 6845 1676
rect 6845 1651 6863 1676
rect 6911 1651 6917 1676
rect 6917 1651 6955 1676
rect 6955 1651 6963 1676
rect 7011 1651 7027 1676
rect 7027 1651 7061 1676
rect 7061 1651 7063 1676
rect 7111 1651 7133 1676
rect 7133 1651 7163 1676
rect 7211 1651 7243 1676
rect 7243 1651 7263 1676
rect 7311 1651 7315 1676
rect 7315 1651 7349 1676
rect 7349 1651 7363 1676
rect 5628 1601 6320 1642
rect 5628 1567 5630 1601
rect 5630 1567 5664 1601
rect 5664 1567 5702 1601
rect 5702 1567 5736 1601
rect 5736 1567 5774 1601
rect 5774 1567 5808 1601
rect 5808 1567 5846 1601
rect 5846 1567 5880 1601
rect 5880 1567 5918 1601
rect 5918 1567 5952 1601
rect 5952 1567 5990 1601
rect 5990 1567 6024 1601
rect 6024 1567 6062 1601
rect 6062 1567 6096 1601
rect 6096 1567 6134 1601
rect 6134 1567 6168 1601
rect 6168 1567 6206 1601
rect 6206 1567 6240 1601
rect 6240 1567 6278 1601
rect 6278 1567 6312 1601
rect 6312 1567 6320 1601
rect 6611 1567 6629 1568
rect 6629 1567 6663 1568
rect 6711 1567 6739 1568
rect 6739 1567 6763 1568
rect 6811 1567 6845 1568
rect 6845 1567 6863 1568
rect 6911 1567 6917 1568
rect 6917 1567 6955 1568
rect 6955 1567 6963 1568
rect 7011 1567 7027 1568
rect 7027 1567 7061 1568
rect 7061 1567 7063 1568
rect 7111 1567 7133 1568
rect 7133 1567 7163 1568
rect 7211 1567 7243 1568
rect 7243 1567 7263 1568
rect 7311 1567 7315 1568
rect 7315 1567 7349 1568
rect 7349 1567 7363 1568
rect 5628 1526 6320 1567
rect 6611 1526 6663 1567
rect 6711 1526 6763 1567
rect 6811 1526 6863 1567
rect 6911 1526 6963 1567
rect 7011 1526 7063 1567
rect 7111 1526 7163 1567
rect 7211 1526 7263 1567
rect 7311 1526 7363 1567
rect 5628 1492 5630 1526
rect 5630 1492 5664 1526
rect 5664 1492 5702 1526
rect 5702 1492 5736 1526
rect 5736 1492 5774 1526
rect 5774 1492 5808 1526
rect 5808 1492 5846 1526
rect 5846 1492 5880 1526
rect 5880 1492 5918 1526
rect 5918 1492 5952 1526
rect 5952 1492 5990 1526
rect 5990 1492 6024 1526
rect 6024 1492 6062 1526
rect 6062 1492 6096 1526
rect 6096 1492 6134 1526
rect 6134 1492 6168 1526
rect 6168 1492 6206 1526
rect 6206 1492 6240 1526
rect 6240 1492 6278 1526
rect 6278 1492 6312 1526
rect 6312 1492 6320 1526
rect 6611 1516 6629 1526
rect 6629 1516 6663 1526
rect 6711 1516 6739 1526
rect 6739 1516 6763 1526
rect 6811 1516 6845 1526
rect 6845 1516 6863 1526
rect 6911 1516 6917 1526
rect 6917 1516 6955 1526
rect 6955 1516 6963 1526
rect 7011 1516 7027 1526
rect 7027 1516 7061 1526
rect 7061 1516 7063 1526
rect 7111 1516 7133 1526
rect 7133 1516 7163 1526
rect 7211 1516 7243 1526
rect 7243 1516 7263 1526
rect 7311 1516 7315 1526
rect 7315 1516 7349 1526
rect 7349 1516 7363 1526
rect 5628 1451 6320 1492
rect 5628 1417 5630 1451
rect 5630 1417 5664 1451
rect 5664 1417 5702 1451
rect 5702 1417 5736 1451
rect 5736 1417 5774 1451
rect 5774 1417 5808 1451
rect 5808 1417 5846 1451
rect 5846 1417 5880 1451
rect 5880 1417 5918 1451
rect 5918 1417 5952 1451
rect 5952 1417 5990 1451
rect 5990 1417 6024 1451
rect 6024 1417 6062 1451
rect 6062 1417 6096 1451
rect 6096 1417 6134 1451
rect 6134 1417 6168 1451
rect 6168 1417 6206 1451
rect 6206 1417 6240 1451
rect 6240 1417 6278 1451
rect 6278 1417 6312 1451
rect 6312 1417 6320 1451
rect 6611 1417 6629 1433
rect 6629 1417 6663 1433
rect 6711 1417 6739 1433
rect 6739 1417 6763 1433
rect 6811 1417 6845 1433
rect 6845 1417 6863 1433
rect 6911 1417 6917 1433
rect 6917 1417 6955 1433
rect 6955 1417 6963 1433
rect 7011 1417 7027 1433
rect 7027 1417 7061 1433
rect 7061 1417 7063 1433
rect 7111 1417 7133 1433
rect 7133 1417 7163 1433
rect 7211 1417 7243 1433
rect 7243 1417 7263 1433
rect 7311 1417 7315 1433
rect 7315 1417 7349 1433
rect 7349 1417 7363 1433
rect 5628 1376 6320 1417
rect 6611 1381 6663 1417
rect 6711 1381 6763 1417
rect 6811 1381 6863 1417
rect 6911 1381 6963 1417
rect 7011 1381 7063 1417
rect 7111 1381 7163 1417
rect 7211 1381 7263 1417
rect 7311 1381 7363 1417
rect 5628 1342 5630 1376
rect 5630 1342 5664 1376
rect 5664 1342 5702 1376
rect 5702 1342 5736 1376
rect 5736 1342 5774 1376
rect 5774 1342 5808 1376
rect 5808 1342 5846 1376
rect 5846 1342 5880 1376
rect 5880 1342 5918 1376
rect 5918 1342 5952 1376
rect 5952 1342 5990 1376
rect 5990 1342 6024 1376
rect 6024 1342 6062 1376
rect 6062 1342 6096 1376
rect 6096 1342 6134 1376
rect 6134 1342 6168 1376
rect 6168 1342 6206 1376
rect 6206 1342 6240 1376
rect 6240 1342 6278 1376
rect 6278 1342 6312 1376
rect 6312 1342 6320 1376
rect 5628 1301 6320 1342
rect 5628 1267 5630 1301
rect 5630 1267 5664 1301
rect 5664 1267 5702 1301
rect 5702 1267 5736 1301
rect 5736 1267 5774 1301
rect 5774 1267 5808 1301
rect 5808 1267 5846 1301
rect 5846 1267 5880 1301
rect 5880 1267 5918 1301
rect 5918 1267 5952 1301
rect 5952 1267 5990 1301
rect 5990 1267 6024 1301
rect 6024 1267 6062 1301
rect 6062 1267 6096 1301
rect 6096 1267 6134 1301
rect 6134 1267 6168 1301
rect 6168 1267 6206 1301
rect 6206 1267 6240 1301
rect 6240 1267 6278 1301
rect 6278 1267 6312 1301
rect 6312 1267 6320 1301
rect 6611 1267 6629 1298
rect 6629 1267 6663 1298
rect 6711 1267 6739 1298
rect 6739 1267 6763 1298
rect 6811 1267 6845 1298
rect 6845 1267 6863 1298
rect 6911 1267 6917 1298
rect 6917 1267 6955 1298
rect 6955 1267 6963 1298
rect 7011 1267 7027 1298
rect 7027 1267 7061 1298
rect 7061 1267 7063 1298
rect 7111 1267 7133 1298
rect 7133 1267 7163 1298
rect 7211 1267 7243 1298
rect 7243 1267 7263 1298
rect 7311 1267 7315 1298
rect 7315 1267 7349 1298
rect 7349 1267 7363 1298
rect 5628 1226 6320 1267
rect 6611 1246 6663 1267
rect 6711 1246 6763 1267
rect 6811 1246 6863 1267
rect 6911 1246 6963 1267
rect 7011 1246 7063 1267
rect 7111 1246 7163 1267
rect 7211 1246 7263 1267
rect 7311 1246 7363 1267
rect 5628 1192 5630 1226
rect 5630 1192 5664 1226
rect 5664 1192 5702 1226
rect 5702 1192 5736 1226
rect 5736 1192 5774 1226
rect 5774 1192 5808 1226
rect 5808 1192 5846 1226
rect 5846 1192 5880 1226
rect 5880 1192 5918 1226
rect 5918 1192 5952 1226
rect 5952 1192 5990 1226
rect 5990 1192 6024 1226
rect 6024 1192 6062 1226
rect 6062 1192 6096 1226
rect 6096 1192 6134 1226
rect 6134 1192 6168 1226
rect 6168 1192 6206 1226
rect 6206 1192 6240 1226
rect 6240 1192 6278 1226
rect 6278 1192 6312 1226
rect 6312 1192 6320 1226
rect 5628 1152 6320 1192
rect 6611 1151 6663 1163
rect 6711 1151 6763 1163
rect 6811 1151 6863 1163
rect 6911 1151 6963 1163
rect 7011 1151 7063 1163
rect 7111 1151 7163 1163
rect 7211 1151 7263 1163
rect 7311 1151 7363 1163
rect 5628 1117 5630 1139
rect 5630 1117 5664 1139
rect 5664 1117 5680 1139
rect 5628 1087 5680 1117
rect 5692 1117 5702 1139
rect 5702 1117 5736 1139
rect 5736 1117 5744 1139
rect 5692 1087 5744 1117
rect 5756 1117 5774 1139
rect 5774 1117 5808 1139
rect 5756 1087 5808 1117
rect 5820 1117 5846 1139
rect 5846 1117 5872 1139
rect 5884 1117 5918 1139
rect 5918 1117 5936 1139
rect 5948 1117 5952 1139
rect 5952 1117 5990 1139
rect 5990 1117 6000 1139
rect 6012 1117 6024 1139
rect 6024 1117 6062 1139
rect 6062 1117 6064 1139
rect 6076 1117 6096 1139
rect 6096 1117 6128 1139
rect 6140 1117 6168 1139
rect 6168 1117 6192 1139
rect 5820 1087 5872 1117
rect 5884 1087 5936 1117
rect 5948 1087 6000 1117
rect 6012 1087 6064 1117
rect 6076 1087 6128 1117
rect 6140 1087 6192 1117
rect 6204 1117 6206 1139
rect 6206 1117 6240 1139
rect 6240 1117 6256 1139
rect 6204 1087 6256 1117
rect 6268 1117 6278 1139
rect 6278 1117 6312 1139
rect 6312 1117 6320 1139
rect 6611 1117 6629 1151
rect 6629 1117 6663 1151
rect 6711 1117 6739 1151
rect 6739 1117 6763 1151
rect 6811 1117 6845 1151
rect 6845 1117 6863 1151
rect 6911 1117 6917 1151
rect 6917 1117 6955 1151
rect 6955 1117 6963 1151
rect 7011 1117 7027 1151
rect 7027 1117 7061 1151
rect 7061 1117 7063 1151
rect 7111 1117 7133 1151
rect 7133 1117 7163 1151
rect 7211 1117 7243 1151
rect 7243 1117 7263 1151
rect 7311 1117 7315 1151
rect 7315 1117 7349 1151
rect 7349 1117 7363 1151
rect 6268 1087 6320 1117
rect 6611 1111 6663 1117
rect 6711 1111 6763 1117
rect 6811 1111 6863 1117
rect 6911 1111 6963 1117
rect 7011 1111 7063 1117
rect 7111 1111 7163 1117
rect 7211 1111 7263 1117
rect 7311 1111 7363 1117
rect 5628 1042 5630 1074
rect 5630 1042 5664 1074
rect 5664 1042 5680 1074
rect 5628 1022 5680 1042
rect 5692 1042 5702 1074
rect 5702 1042 5736 1074
rect 5736 1042 5744 1074
rect 5692 1022 5744 1042
rect 5756 1042 5774 1074
rect 5774 1042 5808 1074
rect 5756 1022 5808 1042
rect 5820 1042 5846 1074
rect 5846 1042 5872 1074
rect 5884 1042 5918 1074
rect 5918 1042 5936 1074
rect 5948 1042 5952 1074
rect 5952 1042 5990 1074
rect 5990 1042 6000 1074
rect 6012 1042 6024 1074
rect 6024 1042 6062 1074
rect 6062 1042 6064 1074
rect 6076 1042 6096 1074
rect 6096 1042 6128 1074
rect 6140 1042 6168 1074
rect 6168 1042 6192 1074
rect 5820 1022 5872 1042
rect 5884 1022 5936 1042
rect 5948 1022 6000 1042
rect 6012 1022 6064 1042
rect 6076 1022 6128 1042
rect 6140 1022 6192 1042
rect 6204 1042 6206 1074
rect 6206 1042 6240 1074
rect 6240 1042 6256 1074
rect 6204 1022 6256 1042
rect 6268 1042 6278 1074
rect 6278 1042 6312 1074
rect 6312 1042 6320 1074
rect 6268 1022 6320 1042
rect 5628 1001 5680 1009
rect 5628 967 5630 1001
rect 5630 967 5664 1001
rect 5664 967 5680 1001
rect 5628 957 5680 967
rect 5692 1001 5744 1009
rect 5692 967 5702 1001
rect 5702 967 5736 1001
rect 5736 967 5744 1001
rect 5692 957 5744 967
rect 5756 1001 5808 1009
rect 5756 967 5774 1001
rect 5774 967 5808 1001
rect 5756 957 5808 967
rect 5820 1001 5872 1009
rect 5884 1001 5936 1009
rect 5948 1001 6000 1009
rect 6012 1001 6064 1009
rect 6076 1001 6128 1009
rect 6140 1001 6192 1009
rect 5820 967 5846 1001
rect 5846 967 5872 1001
rect 5884 967 5918 1001
rect 5918 967 5936 1001
rect 5948 967 5952 1001
rect 5952 967 5990 1001
rect 5990 967 6000 1001
rect 6012 967 6024 1001
rect 6024 967 6062 1001
rect 6062 967 6064 1001
rect 6076 967 6096 1001
rect 6096 967 6128 1001
rect 6140 967 6168 1001
rect 6168 967 6192 1001
rect 5820 957 5872 967
rect 5884 957 5936 967
rect 5948 957 6000 967
rect 6012 957 6064 967
rect 6076 957 6128 967
rect 6140 957 6192 967
rect 6204 1001 6256 1009
rect 6204 967 6206 1001
rect 6206 967 6240 1001
rect 6240 967 6256 1001
rect 6204 957 6256 967
rect 6268 1001 6320 1009
rect 6611 1001 6663 1028
rect 6711 1001 6763 1028
rect 6811 1001 6863 1028
rect 6911 1001 6963 1028
rect 7011 1001 7063 1028
rect 7111 1001 7163 1028
rect 7211 1001 7263 1028
rect 7311 1001 7363 1028
rect 6268 967 6278 1001
rect 6278 967 6312 1001
rect 6312 967 6320 1001
rect 6611 976 6629 1001
rect 6629 976 6663 1001
rect 6711 976 6739 1001
rect 6739 976 6763 1001
rect 6811 976 6845 1001
rect 6845 976 6863 1001
rect 6911 976 6917 1001
rect 6917 976 6955 1001
rect 6955 976 6963 1001
rect 7011 976 7027 1001
rect 7027 976 7061 1001
rect 7061 976 7063 1001
rect 7111 976 7133 1001
rect 7133 976 7163 1001
rect 7211 976 7243 1001
rect 7243 976 7263 1001
rect 7311 976 7315 1001
rect 7315 976 7349 1001
rect 7349 976 7363 1001
rect 6268 957 6320 967
rect 5628 926 5680 944
rect 5628 892 5630 926
rect 5630 892 5664 926
rect 5664 892 5680 926
rect 5692 926 5744 944
rect 5692 892 5702 926
rect 5702 892 5736 926
rect 5736 892 5744 926
rect 5756 926 5808 944
rect 5756 892 5774 926
rect 5774 892 5808 926
rect 5820 926 5872 944
rect 5884 926 5936 944
rect 5948 926 6000 944
rect 6012 926 6064 944
rect 6076 926 6128 944
rect 6140 926 6192 944
rect 5820 892 5846 926
rect 5846 892 5872 926
rect 5884 892 5918 926
rect 5918 892 5936 926
rect 5948 892 5952 926
rect 5952 892 5990 926
rect 5990 892 6000 926
rect 6012 892 6024 926
rect 6024 892 6062 926
rect 6062 892 6064 926
rect 6076 892 6096 926
rect 6096 892 6128 926
rect 6140 892 6168 926
rect 6168 892 6192 926
rect 6204 926 6256 944
rect 6204 892 6206 926
rect 6206 892 6240 926
rect 6240 892 6256 926
rect 6268 926 6320 944
rect 6268 892 6278 926
rect 6278 892 6312 926
rect 6312 892 6320 926
rect 6611 892 6629 893
rect 6629 892 6663 893
rect 6711 892 6739 893
rect 6739 892 6763 893
rect 6811 892 6845 893
rect 6845 892 6863 893
rect 6911 892 6917 893
rect 6917 892 6955 893
rect 6955 892 6963 893
rect 7011 892 7027 893
rect 7027 892 7061 893
rect 7061 892 7063 893
rect 7111 892 7133 893
rect 7133 892 7163 893
rect 7211 892 7243 893
rect 7243 892 7263 893
rect 7311 892 7315 893
rect 7315 892 7349 893
rect 7349 892 7363 893
rect 5628 851 5680 879
rect 5628 827 5630 851
rect 5630 827 5664 851
rect 5664 827 5680 851
rect 5692 851 5744 879
rect 5692 827 5702 851
rect 5702 827 5736 851
rect 5736 827 5744 851
rect 5756 851 5808 879
rect 5756 827 5774 851
rect 5774 827 5808 851
rect 5820 851 5872 879
rect 5884 851 5936 879
rect 5948 851 6000 879
rect 6012 851 6064 879
rect 6076 851 6128 879
rect 6140 851 6192 879
rect 5820 827 5846 851
rect 5846 827 5872 851
rect 5884 827 5918 851
rect 5918 827 5936 851
rect 5948 827 5952 851
rect 5952 827 5990 851
rect 5990 827 6000 851
rect 6012 827 6024 851
rect 6024 827 6062 851
rect 6062 827 6064 851
rect 6076 827 6096 851
rect 6096 827 6128 851
rect 6140 827 6168 851
rect 6168 827 6192 851
rect 6204 851 6256 879
rect 6204 827 6206 851
rect 6206 827 6240 851
rect 6240 827 6256 851
rect 6268 851 6320 879
rect 6611 851 6663 892
rect 6711 851 6763 892
rect 6811 851 6863 892
rect 6911 851 6963 892
rect 7011 851 7063 892
rect 7111 851 7163 892
rect 7211 851 7263 892
rect 7311 851 7363 892
rect 6268 827 6278 851
rect 6278 827 6312 851
rect 6312 827 6320 851
rect 6611 841 6629 851
rect 6629 841 6663 851
rect 6711 841 6739 851
rect 6739 841 6763 851
rect 6811 841 6845 851
rect 6845 841 6863 851
rect 6911 841 6917 851
rect 6917 841 6955 851
rect 6955 841 6963 851
rect 7011 841 7027 851
rect 7027 841 7061 851
rect 7061 841 7063 851
rect 7111 841 7133 851
rect 7133 841 7163 851
rect 7211 841 7243 851
rect 7243 841 7263 851
rect 7311 841 7315 851
rect 7315 841 7349 851
rect 7349 841 7363 851
rect 5628 776 5680 814
rect 5628 762 5630 776
rect 5630 762 5664 776
rect 5664 762 5680 776
rect 5692 776 5744 814
rect 5692 762 5702 776
rect 5702 762 5736 776
rect 5736 762 5744 776
rect 5756 776 5808 814
rect 5756 762 5774 776
rect 5774 762 5808 776
rect 5820 776 5872 814
rect 5884 776 5936 814
rect 5948 776 6000 814
rect 6012 776 6064 814
rect 6076 776 6128 814
rect 6140 776 6192 814
rect 5820 762 5846 776
rect 5846 762 5872 776
rect 5884 762 5918 776
rect 5918 762 5936 776
rect 5948 762 5952 776
rect 5952 762 5990 776
rect 5990 762 6000 776
rect 6012 762 6024 776
rect 6024 762 6062 776
rect 6062 762 6064 776
rect 6076 762 6096 776
rect 6096 762 6128 776
rect 6140 762 6168 776
rect 6168 762 6192 776
rect 6204 776 6256 814
rect 6204 762 6206 776
rect 6206 762 6240 776
rect 6240 762 6256 776
rect 6268 776 6320 814
rect 6268 762 6278 776
rect 6278 762 6312 776
rect 6312 762 6320 776
rect 5628 742 5630 749
rect 5630 742 5664 749
rect 5664 742 5680 749
rect 5628 701 5680 742
rect 5628 697 5630 701
rect 5630 697 5664 701
rect 5664 697 5680 701
rect 5692 742 5702 749
rect 5702 742 5736 749
rect 5736 742 5744 749
rect 5692 701 5744 742
rect 5692 697 5702 701
rect 5702 697 5736 701
rect 5736 697 5744 701
rect 5756 742 5774 749
rect 5774 742 5808 749
rect 5756 701 5808 742
rect 5756 697 5774 701
rect 5774 697 5808 701
rect 5820 742 5846 749
rect 5846 742 5872 749
rect 5884 742 5918 749
rect 5918 742 5936 749
rect 5948 742 5952 749
rect 5952 742 5990 749
rect 5990 742 6000 749
rect 6012 742 6024 749
rect 6024 742 6062 749
rect 6062 742 6064 749
rect 6076 742 6096 749
rect 6096 742 6128 749
rect 6140 742 6168 749
rect 6168 742 6192 749
rect 5820 701 5872 742
rect 5884 701 5936 742
rect 5948 701 6000 742
rect 6012 701 6064 742
rect 6076 701 6128 742
rect 6140 701 6192 742
rect 5820 697 5846 701
rect 5846 697 5872 701
rect 5884 697 5918 701
rect 5918 697 5936 701
rect 5948 697 5952 701
rect 5952 697 5990 701
rect 5990 697 6000 701
rect 6012 697 6024 701
rect 6024 697 6062 701
rect 6062 697 6064 701
rect 6076 697 6096 701
rect 6096 697 6128 701
rect 6140 697 6168 701
rect 6168 697 6192 701
rect 6204 742 6206 749
rect 6206 742 6240 749
rect 6240 742 6256 749
rect 6204 701 6256 742
rect 6204 697 6206 701
rect 6206 697 6240 701
rect 6240 697 6256 701
rect 6268 742 6278 749
rect 6278 742 6312 749
rect 6312 742 6320 749
rect 6611 742 6629 758
rect 6629 742 6663 758
rect 6711 742 6739 758
rect 6739 742 6763 758
rect 6811 742 6845 758
rect 6845 742 6863 758
rect 6911 742 6917 758
rect 6917 742 6955 758
rect 6955 742 6963 758
rect 7011 742 7027 758
rect 7027 742 7061 758
rect 7061 742 7063 758
rect 7111 742 7133 758
rect 7133 742 7163 758
rect 7211 742 7243 758
rect 7243 742 7263 758
rect 7311 742 7315 758
rect 7315 742 7349 758
rect 7349 742 7363 758
rect 6268 701 6320 742
rect 6611 706 6663 742
rect 6711 706 6763 742
rect 6811 706 6863 742
rect 6911 706 6963 742
rect 7011 706 7063 742
rect 7111 706 7163 742
rect 7211 706 7263 742
rect 7311 706 7363 742
rect 6268 697 6278 701
rect 6278 697 6312 701
rect 6312 697 6320 701
rect 5628 667 5630 684
rect 5630 667 5664 684
rect 5664 667 5680 684
rect 5628 632 5680 667
rect 5692 667 5702 684
rect 5702 667 5736 684
rect 5736 667 5744 684
rect 5692 632 5744 667
rect 5756 667 5774 684
rect 5774 667 5808 684
rect 5756 632 5808 667
rect 5820 667 5846 684
rect 5846 667 5872 684
rect 5884 667 5918 684
rect 5918 667 5936 684
rect 5948 667 5952 684
rect 5952 667 5990 684
rect 5990 667 6000 684
rect 6012 667 6024 684
rect 6024 667 6062 684
rect 6062 667 6064 684
rect 6076 667 6096 684
rect 6096 667 6128 684
rect 6140 667 6168 684
rect 6168 667 6192 684
rect 5820 632 5872 667
rect 5884 632 5936 667
rect 5948 632 6000 667
rect 6012 632 6064 667
rect 6076 632 6128 667
rect 6140 632 6192 667
rect 6204 667 6206 684
rect 6206 667 6240 684
rect 6240 667 6256 684
rect 6204 632 6256 667
rect 6268 667 6278 684
rect 6278 667 6312 684
rect 6312 667 6320 684
rect 6268 632 6320 667
rect 5628 592 5630 619
rect 5630 592 5664 619
rect 5664 592 5680 619
rect 5628 567 5680 592
rect 5692 592 5702 619
rect 5702 592 5736 619
rect 5736 592 5744 619
rect 5692 567 5744 592
rect 5756 592 5774 619
rect 5774 592 5808 619
rect 5756 567 5808 592
rect 5820 592 5846 619
rect 5846 592 5872 619
rect 5884 592 5918 619
rect 5918 592 5936 619
rect 5948 592 5952 619
rect 5952 592 5990 619
rect 5990 592 6000 619
rect 6012 592 6024 619
rect 6024 592 6062 619
rect 6062 592 6064 619
rect 6076 592 6096 619
rect 6096 592 6128 619
rect 6140 592 6168 619
rect 6168 592 6192 619
rect 5820 567 5872 592
rect 5884 567 5936 592
rect 5948 567 6000 592
rect 6012 567 6064 592
rect 6076 567 6128 592
rect 6140 567 6192 592
rect 6204 592 6206 619
rect 6206 592 6240 619
rect 6240 592 6256 619
rect 6204 567 6256 592
rect 6268 592 6278 619
rect 6278 592 6312 619
rect 6312 592 6320 619
rect 6611 592 6629 623
rect 6629 592 6663 623
rect 6711 592 6739 623
rect 6739 592 6763 623
rect 6811 592 6845 623
rect 6845 592 6863 623
rect 6911 592 6917 623
rect 6917 592 6955 623
rect 6955 592 6963 623
rect 7011 592 7027 623
rect 7027 592 7061 623
rect 7061 592 7063 623
rect 7111 592 7133 623
rect 7133 592 7163 623
rect 7211 592 7243 623
rect 7243 592 7263 623
rect 7311 592 7315 623
rect 7315 592 7349 623
rect 7349 592 7363 623
rect 6268 567 6320 592
rect 6611 571 6663 592
rect 6711 571 6763 592
rect 6811 571 6863 592
rect 6911 571 6963 592
rect 7011 571 7063 592
rect 7111 571 7163 592
rect 7211 571 7263 592
rect 7311 571 7363 592
rect 5628 551 5680 554
rect 5628 517 5630 551
rect 5630 517 5664 551
rect 5664 517 5680 551
rect 5628 502 5680 517
rect 5692 551 5744 554
rect 5692 517 5702 551
rect 5702 517 5736 551
rect 5736 517 5744 551
rect 5692 502 5744 517
rect 5756 551 5808 554
rect 5756 517 5774 551
rect 5774 517 5808 551
rect 5756 502 5808 517
rect 5820 551 5872 554
rect 5884 551 5936 554
rect 5948 551 6000 554
rect 6012 551 6064 554
rect 6076 551 6128 554
rect 6140 551 6192 554
rect 5820 517 5846 551
rect 5846 517 5872 551
rect 5884 517 5918 551
rect 5918 517 5936 551
rect 5948 517 5952 551
rect 5952 517 5990 551
rect 5990 517 6000 551
rect 6012 517 6024 551
rect 6024 517 6062 551
rect 6062 517 6064 551
rect 6076 517 6096 551
rect 6096 517 6128 551
rect 6140 517 6168 551
rect 6168 517 6192 551
rect 5820 502 5872 517
rect 5884 502 5936 517
rect 5948 502 6000 517
rect 6012 502 6064 517
rect 6076 502 6128 517
rect 6140 502 6192 517
rect 6204 551 6256 554
rect 6204 517 6206 551
rect 6206 517 6240 551
rect 6240 517 6256 551
rect 6204 502 6256 517
rect 6268 551 6320 554
rect 6268 517 6278 551
rect 6278 517 6312 551
rect 6312 517 6320 551
rect 6268 502 6320 517
rect 5628 476 5680 489
rect 5628 442 5630 476
rect 5630 442 5664 476
rect 5664 442 5680 476
rect 5628 437 5680 442
rect 5692 476 5744 489
rect 5692 442 5702 476
rect 5702 442 5736 476
rect 5736 442 5744 476
rect 5692 437 5744 442
rect 5756 476 5808 489
rect 5756 442 5774 476
rect 5774 442 5808 476
rect 5756 437 5808 442
rect 5820 476 5872 489
rect 5884 476 5936 489
rect 5948 476 6000 489
rect 6012 476 6064 489
rect 6076 476 6128 489
rect 6140 476 6192 489
rect 5820 442 5846 476
rect 5846 442 5872 476
rect 5884 442 5918 476
rect 5918 442 5936 476
rect 5948 442 5952 476
rect 5952 442 5990 476
rect 5990 442 6000 476
rect 6012 442 6024 476
rect 6024 442 6062 476
rect 6062 442 6064 476
rect 6076 442 6096 476
rect 6096 442 6128 476
rect 6140 442 6168 476
rect 6168 442 6192 476
rect 5820 437 5872 442
rect 5884 437 5936 442
rect 5948 437 6000 442
rect 6012 437 6064 442
rect 6076 437 6128 442
rect 6140 437 6192 442
rect 6204 476 6256 489
rect 6204 442 6206 476
rect 6206 442 6240 476
rect 6240 442 6256 476
rect 6204 437 6256 442
rect 6268 476 6320 489
rect 6611 476 6663 488
rect 6711 476 6763 488
rect 6811 476 6863 488
rect 6911 476 6963 488
rect 7011 476 7063 488
rect 7111 476 7163 488
rect 7211 476 7263 488
rect 7311 476 7363 488
rect 6268 442 6278 476
rect 6278 442 6312 476
rect 6312 442 6320 476
rect 6611 442 6629 476
rect 6629 442 6663 476
rect 6711 442 6739 476
rect 6739 442 6763 476
rect 6811 442 6845 476
rect 6845 442 6863 476
rect 6911 442 6917 476
rect 6917 442 6955 476
rect 6955 442 6963 476
rect 7011 442 7027 476
rect 7027 442 7061 476
rect 7061 442 7063 476
rect 7111 442 7133 476
rect 7133 442 7163 476
rect 7211 442 7243 476
rect 7243 442 7263 476
rect 7311 442 7315 476
rect 7315 442 7349 476
rect 7349 442 7363 476
rect 6268 437 6320 442
rect 6611 436 6663 442
rect 6711 436 6763 442
rect 6811 436 6863 442
rect 6911 436 6963 442
rect 7011 436 7063 442
rect 7111 436 7163 442
rect 7211 436 7263 442
rect 7311 436 7363 442
<< metal2 >>
rect 2270 38724 8222 38730
rect 2322 38672 2392 38724
rect 2444 38720 5613 38724
rect 5669 38720 5696 38724
rect 2444 38672 2824 38720
rect 2270 38668 2824 38672
rect 2876 38668 2890 38720
rect 2942 38668 3378 38720
rect 3430 38668 3444 38720
rect 3496 38668 3932 38720
rect 3984 38668 3998 38720
rect 4050 38668 4486 38720
rect 4538 38668 4552 38720
rect 4604 38668 5040 38720
rect 5092 38668 5106 38720
rect 5158 38668 5594 38720
rect 5752 38668 5779 38724
rect 5835 38668 5861 38724
rect 5917 38668 5943 38724
rect 5999 38668 6025 38724
rect 6081 38668 6107 38724
rect 6163 38720 6189 38724
rect 6245 38720 6271 38724
rect 6266 38668 6271 38720
rect 6327 38668 6353 38724
rect 6409 38668 6435 38724
rect 6491 38668 6517 38724
rect 6573 38668 6599 38724
rect 6655 38668 6681 38724
rect 6737 38720 6763 38724
rect 6819 38720 6845 38724
rect 6754 38668 6763 38720
rect 6820 38668 6845 38720
rect 6901 38668 6927 38724
rect 6983 38668 7009 38724
rect 7065 38668 7091 38724
rect 7147 38668 7173 38724
rect 7229 38668 7255 38724
rect 7311 38720 7337 38724
rect 7311 38668 7322 38720
rect 7393 38668 7419 38724
rect 7475 38668 7501 38724
rect 7557 38668 7583 38724
rect 7639 38668 7665 38724
rect 7721 38668 7747 38724
rect 7803 38720 7829 38724
rect 7885 38720 7911 38724
rect 7803 38668 7810 38720
rect 7967 38668 7993 38724
rect 8049 38668 8075 38672
rect 8131 38668 8157 38724
rect 8221 38672 8222 38724
rect 8213 38668 8222 38672
rect 2270 38655 8222 38668
rect 2322 38603 2392 38655
rect 2444 38651 8047 38655
rect 2444 38603 2824 38651
rect 2270 38599 2824 38603
rect 2876 38599 2890 38651
rect 2942 38599 3378 38651
rect 3430 38599 3444 38651
rect 3496 38599 3932 38651
rect 3984 38599 3998 38651
rect 4050 38599 4486 38651
rect 4538 38599 4552 38651
rect 4604 38599 5040 38651
rect 5092 38599 5106 38651
rect 5158 38599 5594 38651
rect 5646 38644 5660 38651
rect 5712 38644 6148 38651
rect 6200 38644 6214 38651
rect 6266 38644 6702 38651
rect 6754 38644 6768 38651
rect 6820 38644 7256 38651
rect 7308 38644 7322 38651
rect 7374 38644 7810 38651
rect 7862 38644 7876 38651
rect 7928 38644 8047 38651
rect 8099 38644 8169 38655
rect 2270 38588 5613 38599
rect 5669 38588 5696 38599
rect 5752 38588 5779 38644
rect 5835 38588 5861 38644
rect 5917 38588 5943 38644
rect 5999 38588 6025 38644
rect 6081 38588 6107 38644
rect 6266 38599 6271 38644
rect 6163 38588 6189 38599
rect 6245 38588 6271 38599
rect 6327 38588 6353 38644
rect 6409 38588 6435 38644
rect 6491 38588 6517 38644
rect 6573 38588 6599 38644
rect 6655 38588 6681 38644
rect 6754 38599 6763 38644
rect 6820 38599 6845 38644
rect 6737 38588 6763 38599
rect 6819 38588 6845 38599
rect 6901 38588 6927 38644
rect 6983 38588 7009 38644
rect 7065 38588 7091 38644
rect 7147 38588 7173 38644
rect 7229 38588 7255 38644
rect 7311 38599 7322 38644
rect 7311 38588 7337 38599
rect 7393 38588 7419 38644
rect 7475 38588 7501 38644
rect 7557 38588 7583 38644
rect 7639 38588 7665 38644
rect 7721 38588 7747 38644
rect 7803 38599 7810 38644
rect 7803 38588 7829 38599
rect 7885 38588 7911 38599
rect 7967 38588 7993 38644
rect 8049 38588 8075 38603
rect 8131 38588 8157 38644
rect 8221 38603 8222 38655
rect 8213 38588 8222 38603
rect 2270 38586 8222 38588
rect 2322 38534 2392 38586
rect 2444 38582 8047 38586
rect 2444 38534 2824 38582
rect 2270 38530 2824 38534
rect 2876 38530 2890 38582
rect 2942 38530 3378 38582
rect 3430 38530 3444 38582
rect 3496 38530 3932 38582
rect 3984 38530 3998 38582
rect 4050 38530 4486 38582
rect 4538 38530 4552 38582
rect 4604 38530 5040 38582
rect 5092 38530 5106 38582
rect 5158 38530 5594 38582
rect 5646 38564 5660 38582
rect 5712 38564 6148 38582
rect 6200 38564 6214 38582
rect 6266 38564 6702 38582
rect 6754 38564 6768 38582
rect 6820 38564 7256 38582
rect 7308 38564 7322 38582
rect 7374 38564 7810 38582
rect 7862 38564 7876 38582
rect 7928 38564 8047 38582
rect 8099 38564 8169 38586
rect 2270 38517 5613 38530
rect 2322 38465 2392 38517
rect 2444 38513 5613 38517
rect 5669 38513 5696 38530
rect 2444 38465 2824 38513
rect 2270 38461 2824 38465
rect 2876 38461 2890 38513
rect 2942 38461 3378 38513
rect 3430 38461 3444 38513
rect 3496 38461 3932 38513
rect 3984 38461 3998 38513
rect 4050 38461 4486 38513
rect 4538 38461 4552 38513
rect 4604 38461 5040 38513
rect 5092 38461 5106 38513
rect 5158 38461 5594 38513
rect 5752 38508 5779 38564
rect 5835 38508 5861 38564
rect 5917 38508 5943 38564
rect 5999 38508 6025 38564
rect 6081 38508 6107 38564
rect 6266 38530 6271 38564
rect 6163 38513 6189 38530
rect 6245 38513 6271 38530
rect 6266 38508 6271 38513
rect 6327 38508 6353 38564
rect 6409 38508 6435 38564
rect 6491 38508 6517 38564
rect 6573 38508 6599 38564
rect 6655 38508 6681 38564
rect 6754 38530 6763 38564
rect 6820 38530 6845 38564
rect 6737 38513 6763 38530
rect 6819 38513 6845 38530
rect 6754 38508 6763 38513
rect 6820 38508 6845 38513
rect 6901 38508 6927 38564
rect 6983 38508 7009 38564
rect 7065 38508 7091 38564
rect 7147 38508 7173 38564
rect 7229 38508 7255 38564
rect 7311 38530 7322 38564
rect 7311 38513 7337 38530
rect 7311 38508 7322 38513
rect 7393 38508 7419 38564
rect 7475 38508 7501 38564
rect 7557 38508 7583 38564
rect 7639 38508 7665 38564
rect 7721 38508 7747 38564
rect 7803 38530 7810 38564
rect 7803 38513 7829 38530
rect 7885 38513 7911 38530
rect 7803 38508 7810 38513
rect 7967 38508 7993 38564
rect 8049 38517 8075 38534
rect 8131 38508 8157 38564
rect 8221 38534 8222 38586
rect 8213 38517 8222 38534
rect 5646 38484 5660 38508
rect 5712 38484 6148 38508
rect 6200 38484 6214 38508
rect 6266 38484 6702 38508
rect 6754 38484 6768 38508
rect 6820 38484 7256 38508
rect 7308 38484 7322 38508
rect 7374 38484 7810 38508
rect 7862 38484 7876 38508
rect 7928 38484 8047 38508
rect 8099 38484 8169 38508
rect 2270 38448 5613 38461
rect 2322 38396 2392 38448
rect 2444 38444 5613 38448
rect 5669 38444 5696 38461
rect 2444 38396 2824 38444
rect 2270 38392 2824 38396
rect 2876 38392 2890 38444
rect 2942 38392 3378 38444
rect 3430 38392 3444 38444
rect 3496 38392 3932 38444
rect 3984 38392 3998 38444
rect 4050 38392 4486 38444
rect 4538 38392 4552 38444
rect 4604 38392 5040 38444
rect 5092 38392 5106 38444
rect 5158 38392 5594 38444
rect 5752 38428 5779 38484
rect 5835 38428 5861 38484
rect 5917 38428 5943 38484
rect 5999 38428 6025 38484
rect 6081 38428 6107 38484
rect 6266 38461 6271 38484
rect 6163 38444 6189 38461
rect 6245 38444 6271 38461
rect 6266 38428 6271 38444
rect 6327 38428 6353 38484
rect 6409 38428 6435 38484
rect 6491 38428 6517 38484
rect 6573 38428 6599 38484
rect 6655 38428 6681 38484
rect 6754 38461 6763 38484
rect 6820 38461 6845 38484
rect 6737 38444 6763 38461
rect 6819 38444 6845 38461
rect 6754 38428 6763 38444
rect 6820 38428 6845 38444
rect 6901 38428 6927 38484
rect 6983 38428 7009 38484
rect 7065 38428 7091 38484
rect 7147 38428 7173 38484
rect 7229 38428 7255 38484
rect 7311 38461 7322 38484
rect 7311 38444 7337 38461
rect 7311 38428 7322 38444
rect 7393 38428 7419 38484
rect 7475 38428 7501 38484
rect 7557 38428 7583 38484
rect 7639 38428 7665 38484
rect 7721 38428 7747 38484
rect 7803 38461 7810 38484
rect 7803 38444 7829 38461
rect 7885 38444 7911 38461
rect 7803 38428 7810 38444
rect 7967 38428 7993 38484
rect 8049 38448 8075 38465
rect 8131 38428 8157 38484
rect 8221 38465 8222 38517
rect 8213 38448 8222 38465
rect 5646 38404 5660 38428
rect 5712 38404 6148 38428
rect 6200 38404 6214 38428
rect 6266 38404 6702 38428
rect 6754 38404 6768 38428
rect 6820 38404 7256 38428
rect 7308 38404 7322 38428
rect 7374 38404 7810 38428
rect 7862 38404 7876 38428
rect 7928 38404 8047 38428
rect 8099 38404 8169 38428
rect 2270 38378 5613 38392
rect 2322 38326 2392 38378
rect 2444 38375 5613 38378
rect 5669 38375 5696 38392
rect 2444 38326 2824 38375
rect 2270 38323 2824 38326
rect 2876 38323 2890 38375
rect 2942 38323 3378 38375
rect 3430 38323 3444 38375
rect 3496 38323 3932 38375
rect 3984 38323 3998 38375
rect 4050 38323 4486 38375
rect 4538 38323 4552 38375
rect 4604 38323 5040 38375
rect 5092 38323 5106 38375
rect 5158 38323 5594 38375
rect 5752 38348 5779 38404
rect 5835 38348 5861 38404
rect 5917 38348 5943 38404
rect 5999 38348 6025 38404
rect 6081 38348 6107 38404
rect 6266 38392 6271 38404
rect 6163 38375 6189 38392
rect 6245 38375 6271 38392
rect 6266 38348 6271 38375
rect 6327 38348 6353 38404
rect 6409 38348 6435 38404
rect 6491 38348 6517 38404
rect 6573 38348 6599 38404
rect 6655 38348 6681 38404
rect 6754 38392 6763 38404
rect 6820 38392 6845 38404
rect 6737 38375 6763 38392
rect 6819 38375 6845 38392
rect 6754 38348 6763 38375
rect 6820 38348 6845 38375
rect 6901 38348 6927 38404
rect 6983 38348 7009 38404
rect 7065 38348 7091 38404
rect 7147 38348 7173 38404
rect 7229 38348 7255 38404
rect 7311 38392 7322 38404
rect 7311 38375 7337 38392
rect 7311 38348 7322 38375
rect 7393 38348 7419 38404
rect 7475 38348 7501 38404
rect 7557 38348 7583 38404
rect 7639 38348 7665 38404
rect 7721 38348 7747 38404
rect 7803 38392 7810 38404
rect 7803 38375 7829 38392
rect 7885 38375 7911 38392
rect 7803 38348 7810 38375
rect 7967 38348 7993 38404
rect 8049 38378 8075 38396
rect 8131 38348 8157 38404
rect 8221 38396 8222 38448
rect 8213 38378 8222 38396
rect 5646 38324 5660 38348
rect 5712 38324 6148 38348
rect 6200 38324 6214 38348
rect 6266 38324 6702 38348
rect 6754 38324 6768 38348
rect 6820 38324 7256 38348
rect 7308 38324 7322 38348
rect 7374 38324 7810 38348
rect 7862 38324 7876 38348
rect 7928 38326 8047 38348
rect 8099 38326 8169 38348
rect 8221 38326 8222 38378
rect 7928 38324 8222 38326
rect 2270 38308 5613 38323
rect 2322 38256 2392 38308
rect 2444 38306 5613 38308
rect 5669 38306 5696 38323
rect 2444 38256 2824 38306
rect 2270 38254 2824 38256
rect 2876 38254 2890 38306
rect 2942 38254 3378 38306
rect 3430 38254 3444 38306
rect 3496 38254 3932 38306
rect 3984 38254 3998 38306
rect 4050 38254 4486 38306
rect 4538 38254 4552 38306
rect 4604 38254 5040 38306
rect 5092 38254 5106 38306
rect 5158 38254 5594 38306
rect 5752 38268 5779 38324
rect 5835 38268 5861 38324
rect 5917 38268 5943 38324
rect 5999 38268 6025 38324
rect 6081 38268 6107 38324
rect 6266 38323 6271 38324
rect 6163 38306 6189 38323
rect 6245 38306 6271 38323
rect 6266 38268 6271 38306
rect 6327 38268 6353 38324
rect 6409 38268 6435 38324
rect 6491 38268 6517 38324
rect 6573 38268 6599 38324
rect 6655 38268 6681 38324
rect 6754 38323 6763 38324
rect 6820 38323 6845 38324
rect 6737 38306 6763 38323
rect 6819 38306 6845 38323
rect 6754 38268 6763 38306
rect 6820 38268 6845 38306
rect 6901 38268 6927 38324
rect 6983 38268 7009 38324
rect 7065 38268 7091 38324
rect 7147 38268 7173 38324
rect 7229 38268 7255 38324
rect 7311 38323 7322 38324
rect 7311 38306 7337 38323
rect 7311 38268 7322 38306
rect 7393 38268 7419 38324
rect 7475 38268 7501 38324
rect 7557 38268 7583 38324
rect 7639 38268 7665 38324
rect 7721 38268 7747 38324
rect 7803 38323 7810 38324
rect 7803 38306 7829 38323
rect 7885 38306 7911 38323
rect 7803 38268 7810 38306
rect 7967 38268 7993 38324
rect 8049 38308 8075 38324
rect 8131 38268 8157 38324
rect 8213 38308 8222 38324
rect 5646 38254 5660 38268
rect 5712 38254 6148 38268
rect 6200 38254 6214 38268
rect 6266 38254 6702 38268
rect 6754 38254 6768 38268
rect 6820 38254 7256 38268
rect 7308 38254 7322 38268
rect 7374 38254 7810 38268
rect 7862 38254 7876 38268
rect 7928 38256 8047 38268
rect 8099 38256 8169 38268
rect 8221 38256 8222 38308
rect 7928 38254 8222 38256
rect 2270 38244 8222 38254
rect 2270 38238 5613 38244
rect 2322 38186 2392 38238
rect 2444 38236 5613 38238
rect 5669 38236 5696 38244
rect 2444 38186 2824 38236
rect 2270 38184 2824 38186
rect 2876 38184 2890 38236
rect 2942 38184 3378 38236
rect 3430 38184 3444 38236
rect 3496 38184 3932 38236
rect 3984 38184 3998 38236
rect 4050 38184 4486 38236
rect 4538 38184 4552 38236
rect 4604 38184 5040 38236
rect 5092 38184 5106 38236
rect 5158 38184 5594 38236
rect 5752 38188 5779 38244
rect 5835 38188 5861 38244
rect 5917 38188 5943 38244
rect 5999 38188 6025 38244
rect 6081 38188 6107 38244
rect 6163 38236 6189 38244
rect 6245 38236 6271 38244
rect 6266 38188 6271 38236
rect 6327 38188 6353 38244
rect 6409 38188 6435 38244
rect 6491 38188 6517 38244
rect 6573 38188 6599 38244
rect 6655 38188 6681 38244
rect 6737 38236 6763 38244
rect 6819 38236 6845 38244
rect 6754 38188 6763 38236
rect 6820 38188 6845 38236
rect 6901 38188 6927 38244
rect 6983 38188 7009 38244
rect 7065 38188 7091 38244
rect 7147 38188 7173 38244
rect 7229 38188 7255 38244
rect 7311 38236 7337 38244
rect 7311 38188 7322 38236
rect 7393 38188 7419 38244
rect 7475 38188 7501 38244
rect 7557 38188 7583 38244
rect 7639 38188 7665 38244
rect 7721 38188 7747 38244
rect 7803 38236 7829 38244
rect 7885 38236 7911 38244
rect 7803 38188 7810 38236
rect 7967 38188 7993 38244
rect 8049 38238 8075 38244
rect 8131 38188 8157 38244
rect 8213 38238 8222 38244
rect 5646 38184 5660 38188
rect 5712 38184 6148 38188
rect 6200 38184 6214 38188
rect 6266 38184 6702 38188
rect 6754 38184 6768 38188
rect 6820 38184 7256 38188
rect 7308 38184 7322 38188
rect 7374 38184 7810 38188
rect 7862 38184 7876 38188
rect 7928 38186 8047 38188
rect 8099 38186 8169 38188
rect 8221 38186 8222 38238
rect 7928 38184 8222 38186
rect 2270 38168 8222 38184
rect 2322 38116 2392 38168
rect 2444 38166 8047 38168
rect 2444 38116 2824 38166
rect 2270 38114 2824 38116
rect 2876 38114 2890 38166
rect 2942 38114 3378 38166
rect 3430 38114 3444 38166
rect 3496 38114 3932 38166
rect 3984 38114 3998 38166
rect 4050 38114 4486 38166
rect 4538 38114 4552 38166
rect 4604 38114 5040 38166
rect 5092 38114 5106 38166
rect 5158 38114 5594 38166
rect 5646 38164 5660 38166
rect 5712 38164 6148 38166
rect 6200 38164 6214 38166
rect 6266 38164 6702 38166
rect 6754 38164 6768 38166
rect 6820 38164 7256 38166
rect 7308 38164 7322 38166
rect 7374 38164 7810 38166
rect 7862 38164 7876 38166
rect 7928 38164 8047 38166
rect 8099 38164 8169 38168
rect 2270 38108 5613 38114
rect 5669 38108 5696 38114
rect 5752 38108 5779 38164
rect 5835 38108 5861 38164
rect 5917 38108 5943 38164
rect 5999 38108 6025 38164
rect 6081 38108 6107 38164
rect 6266 38114 6271 38164
rect 6163 38108 6189 38114
rect 6245 38108 6271 38114
rect 6327 38108 6353 38164
rect 6409 38108 6435 38164
rect 6491 38108 6517 38164
rect 6573 38108 6599 38164
rect 6655 38108 6681 38164
rect 6754 38114 6763 38164
rect 6820 38114 6845 38164
rect 6737 38108 6763 38114
rect 6819 38108 6845 38114
rect 6901 38108 6927 38164
rect 6983 38108 7009 38164
rect 7065 38108 7091 38164
rect 7147 38108 7173 38164
rect 7229 38108 7255 38164
rect 7311 38114 7322 38164
rect 7311 38108 7337 38114
rect 7393 38108 7419 38164
rect 7475 38108 7501 38164
rect 7557 38108 7583 38164
rect 7639 38108 7665 38164
rect 7721 38108 7747 38164
rect 7803 38114 7810 38164
rect 7803 38108 7829 38114
rect 7885 38108 7911 38114
rect 7967 38108 7993 38164
rect 8049 38108 8075 38116
rect 8131 38108 8157 38164
rect 8221 38116 8222 38168
rect 8213 38108 8222 38116
rect 2729 37987 7651 37988
rect 2729 37931 2738 37987
rect 2794 37931 2819 37987
rect 2875 37931 2900 37987
rect 2956 37931 2981 37987
rect 3037 37931 3062 37987
rect 3118 37982 3143 37987
rect 3199 37982 3224 37987
rect 3219 37931 3224 37982
rect 3280 37931 3305 37987
rect 3361 37931 3386 37987
rect 3442 37931 3467 37987
rect 3523 37931 3548 37987
rect 3604 37931 3629 37987
rect 3685 37982 3710 37987
rect 3766 37982 3791 37987
rect 3707 37931 3710 37982
rect 3773 37931 3791 37982
rect 3847 37931 3872 37987
rect 3928 37931 3953 37987
rect 4009 37931 4034 37987
rect 4090 37931 4115 37987
rect 4171 37931 4196 37987
rect 4252 37982 4277 37987
rect 2729 37930 3101 37931
rect 3153 37930 3167 37931
rect 3219 37930 3655 37931
rect 3707 37930 3721 37931
rect 3773 37930 4209 37931
rect 4261 37930 4275 37982
rect 4333 37931 4358 37987
rect 4414 37931 4439 37987
rect 4495 37931 4520 37987
rect 4576 37931 4601 37987
rect 4657 37931 4682 37987
rect 4738 37931 4763 37987
rect 5299 37982 7651 37987
rect 4327 37930 4763 37931
rect 5299 37930 5317 37982
rect 5369 37930 5383 37982
rect 5435 37930 5871 37982
rect 5923 37930 5937 37982
rect 5989 37930 6425 37982
rect 6477 37930 6491 37982
rect 6543 37930 6979 37982
rect 7031 37930 7045 37982
rect 7097 37930 7533 37982
rect 7585 37930 7599 37982
rect 2729 37913 4763 37930
rect 5299 37913 7651 37930
rect 2729 37907 3101 37913
rect 3153 37907 3167 37913
rect 3219 37907 3655 37913
rect 3707 37907 3721 37913
rect 3773 37907 4209 37913
rect 2729 37851 2738 37907
rect 2794 37851 2819 37907
rect 2875 37851 2900 37907
rect 2956 37851 2981 37907
rect 3037 37851 3062 37907
rect 3219 37861 3224 37907
rect 3118 37851 3143 37861
rect 3199 37851 3224 37861
rect 3280 37851 3305 37907
rect 3361 37851 3386 37907
rect 3442 37851 3467 37907
rect 3523 37851 3548 37907
rect 3604 37851 3629 37907
rect 3707 37861 3710 37907
rect 3773 37861 3791 37907
rect 3685 37851 3710 37861
rect 3766 37851 3791 37861
rect 3847 37851 3872 37907
rect 3928 37851 3953 37907
rect 4009 37851 4034 37907
rect 4090 37851 4115 37907
rect 4171 37851 4196 37907
rect 4261 37861 4275 37913
rect 4327 37907 4763 37913
rect 4252 37851 4277 37861
rect 4333 37851 4358 37907
rect 4414 37851 4439 37907
rect 4495 37851 4520 37907
rect 4576 37851 4601 37907
rect 4657 37851 4682 37907
rect 4738 37851 4763 37907
rect 5299 37861 5317 37913
rect 5369 37861 5383 37913
rect 5435 37861 5871 37913
rect 5923 37861 5937 37913
rect 5989 37861 6425 37913
rect 6477 37861 6491 37913
rect 6543 37861 6979 37913
rect 7031 37861 7045 37913
rect 7097 37861 7533 37913
rect 7585 37861 7599 37913
rect 2729 37844 4763 37851
rect 5299 37844 7651 37861
rect 2729 37827 3101 37844
rect 3153 37827 3167 37844
rect 3219 37827 3655 37844
rect 3707 37827 3721 37844
rect 3773 37827 4209 37844
rect 2729 37771 2738 37827
rect 2794 37771 2819 37827
rect 2875 37771 2900 37827
rect 2956 37771 2981 37827
rect 3037 37771 3062 37827
rect 3219 37792 3224 37827
rect 3118 37775 3143 37792
rect 3199 37775 3224 37792
rect 3219 37771 3224 37775
rect 3280 37771 3305 37827
rect 3361 37771 3386 37827
rect 3442 37771 3467 37827
rect 3523 37771 3548 37827
rect 3604 37771 3629 37827
rect 3707 37792 3710 37827
rect 3773 37792 3791 37827
rect 3685 37775 3710 37792
rect 3766 37775 3791 37792
rect 3707 37771 3710 37775
rect 3773 37771 3791 37775
rect 3847 37771 3872 37827
rect 3928 37771 3953 37827
rect 4009 37771 4034 37827
rect 4090 37771 4115 37827
rect 4171 37771 4196 37827
rect 4261 37792 4275 37844
rect 4327 37827 4763 37844
rect 4252 37775 4277 37792
rect 2729 37747 3101 37771
rect 3153 37747 3167 37771
rect 3219 37747 3655 37771
rect 3707 37747 3721 37771
rect 3773 37747 4209 37771
rect 2729 37691 2738 37747
rect 2794 37691 2819 37747
rect 2875 37691 2900 37747
rect 2956 37691 2981 37747
rect 3037 37691 3062 37747
rect 3219 37723 3224 37747
rect 3118 37706 3143 37723
rect 3199 37706 3224 37723
rect 3219 37691 3224 37706
rect 3280 37691 3305 37747
rect 3361 37691 3386 37747
rect 3442 37691 3467 37747
rect 3523 37691 3548 37747
rect 3604 37691 3629 37747
rect 3707 37723 3710 37747
rect 3773 37723 3791 37747
rect 3685 37706 3710 37723
rect 3766 37706 3791 37723
rect 3707 37691 3710 37706
rect 3773 37691 3791 37706
rect 3847 37691 3872 37747
rect 3928 37691 3953 37747
rect 4009 37691 4034 37747
rect 4090 37691 4115 37747
rect 4171 37691 4196 37747
rect 4261 37723 4275 37775
rect 4333 37771 4358 37827
rect 4414 37771 4439 37827
rect 4495 37771 4520 37827
rect 4576 37771 4601 37827
rect 4657 37771 4682 37827
rect 4738 37771 4763 37827
rect 5299 37792 5317 37844
rect 5369 37792 5383 37844
rect 5435 37792 5871 37844
rect 5923 37792 5937 37844
rect 5989 37792 6425 37844
rect 6477 37792 6491 37844
rect 6543 37792 6979 37844
rect 7031 37792 7045 37844
rect 7097 37792 7533 37844
rect 7585 37792 7599 37844
rect 5299 37775 7651 37792
rect 4327 37747 4763 37771
rect 4252 37706 4277 37723
rect 2729 37667 3101 37691
rect 3153 37667 3167 37691
rect 3219 37667 3655 37691
rect 3707 37667 3721 37691
rect 3773 37667 4209 37691
rect 2729 37611 2738 37667
rect 2794 37611 2819 37667
rect 2875 37611 2900 37667
rect 2956 37611 2981 37667
rect 3037 37611 3062 37667
rect 3219 37654 3224 37667
rect 3118 37636 3143 37654
rect 3199 37636 3224 37654
rect 3219 37611 3224 37636
rect 3280 37611 3305 37667
rect 3361 37611 3386 37667
rect 3442 37611 3467 37667
rect 3523 37611 3548 37667
rect 3604 37611 3629 37667
rect 3707 37654 3710 37667
rect 3773 37654 3791 37667
rect 3685 37636 3710 37654
rect 3766 37636 3791 37654
rect 3707 37611 3710 37636
rect 3773 37611 3791 37636
rect 3847 37611 3872 37667
rect 3928 37611 3953 37667
rect 4009 37611 4034 37667
rect 4090 37611 4115 37667
rect 4171 37611 4196 37667
rect 4261 37654 4275 37706
rect 4333 37691 4358 37747
rect 4414 37691 4439 37747
rect 4495 37691 4520 37747
rect 4576 37691 4601 37747
rect 4657 37691 4682 37747
rect 4738 37691 4763 37747
rect 5299 37723 5317 37775
rect 5369 37723 5383 37775
rect 5435 37723 5871 37775
rect 5923 37723 5937 37775
rect 5989 37723 6425 37775
rect 6477 37723 6491 37775
rect 6543 37723 6979 37775
rect 7031 37723 7045 37775
rect 7097 37723 7533 37775
rect 7585 37723 7599 37775
rect 5299 37706 7651 37723
rect 4327 37667 4763 37691
rect 4252 37636 4277 37654
rect 2729 37587 3101 37611
rect 3153 37587 3167 37611
rect 3219 37587 3655 37611
rect 3707 37587 3721 37611
rect 3773 37587 4209 37611
rect 2729 37531 2738 37587
rect 2794 37531 2819 37587
rect 2875 37531 2900 37587
rect 2956 37531 2981 37587
rect 3037 37531 3062 37587
rect 3219 37584 3224 37587
rect 3118 37566 3143 37584
rect 3199 37566 3224 37584
rect 3219 37531 3224 37566
rect 3280 37531 3305 37587
rect 3361 37531 3386 37587
rect 3442 37531 3467 37587
rect 3523 37531 3548 37587
rect 3604 37531 3629 37587
rect 3707 37584 3710 37587
rect 3773 37584 3791 37587
rect 3685 37566 3710 37584
rect 3766 37566 3791 37584
rect 3707 37531 3710 37566
rect 3773 37531 3791 37566
rect 3847 37531 3872 37587
rect 3928 37531 3953 37587
rect 4009 37531 4034 37587
rect 4090 37531 4115 37587
rect 4171 37531 4196 37587
rect 4261 37584 4275 37636
rect 4333 37611 4358 37667
rect 4414 37611 4439 37667
rect 4495 37611 4520 37667
rect 4576 37611 4601 37667
rect 4657 37611 4682 37667
rect 4738 37611 4763 37667
rect 5299 37654 5317 37706
rect 5369 37654 5383 37706
rect 5435 37654 5871 37706
rect 5923 37654 5937 37706
rect 5989 37654 6425 37706
rect 6477 37654 6491 37706
rect 6543 37654 6979 37706
rect 7031 37654 7045 37706
rect 7097 37654 7533 37706
rect 7585 37654 7599 37706
rect 5299 37636 7651 37654
rect 4327 37587 4763 37611
rect 4252 37566 4277 37584
rect 2729 37514 3101 37531
rect 3153 37514 3167 37531
rect 3219 37514 3655 37531
rect 3707 37514 3721 37531
rect 3773 37514 4209 37531
rect 4261 37514 4275 37566
rect 4333 37531 4358 37587
rect 4414 37531 4439 37587
rect 4495 37531 4520 37587
rect 4576 37531 4601 37587
rect 4657 37531 4682 37587
rect 4738 37531 4763 37587
rect 5299 37584 5317 37636
rect 5369 37584 5383 37636
rect 5435 37584 5871 37636
rect 5923 37584 5937 37636
rect 5989 37584 6425 37636
rect 6477 37584 6491 37636
rect 6543 37584 6979 37636
rect 7031 37584 7045 37636
rect 7097 37584 7533 37636
rect 7585 37584 7599 37636
rect 5299 37566 7651 37584
rect 4327 37514 4763 37531
rect 5299 37514 5317 37566
rect 5369 37514 5383 37566
rect 5435 37514 5871 37566
rect 5923 37514 5937 37566
rect 5989 37514 6425 37566
rect 6477 37514 6491 37566
rect 6543 37514 6979 37566
rect 7031 37514 7045 37566
rect 7097 37514 7533 37566
rect 7585 37514 7599 37566
rect 2729 37507 4763 37514
rect 2729 37451 2738 37507
rect 2794 37451 2819 37507
rect 2875 37451 2900 37507
rect 2956 37451 2981 37507
rect 3037 37451 3062 37507
rect 3118 37496 3143 37507
rect 3199 37496 3224 37507
rect 3219 37451 3224 37496
rect 3280 37451 3305 37507
rect 3361 37451 3386 37507
rect 3442 37451 3467 37507
rect 3523 37451 3548 37507
rect 3604 37451 3629 37507
rect 3685 37496 3710 37507
rect 3766 37496 3791 37507
rect 3707 37451 3710 37496
rect 3773 37451 3791 37496
rect 3847 37451 3872 37507
rect 3928 37451 3953 37507
rect 4009 37451 4034 37507
rect 4090 37451 4115 37507
rect 4171 37451 4196 37507
rect 4252 37496 4277 37507
rect 2729 37444 3101 37451
rect 3153 37444 3167 37451
rect 3219 37444 3655 37451
rect 3707 37444 3721 37451
rect 3773 37444 4209 37451
rect 4261 37444 4275 37496
rect 4333 37451 4358 37507
rect 4414 37451 4439 37507
rect 4495 37451 4520 37507
rect 4576 37451 4601 37507
rect 4657 37451 4682 37507
rect 4738 37451 4763 37507
rect 5299 37496 7651 37514
rect 4327 37444 4763 37451
rect 5299 37444 5317 37496
rect 5369 37444 5383 37496
rect 5435 37444 5871 37496
rect 5923 37444 5937 37496
rect 5989 37444 6425 37496
rect 6477 37444 6491 37496
rect 6543 37444 6979 37496
rect 7031 37444 7045 37496
rect 7097 37444 7533 37496
rect 7585 37444 7599 37496
rect 2729 37427 4763 37444
rect 2729 37371 2738 37427
rect 2794 37371 2819 37427
rect 2875 37371 2900 37427
rect 2956 37371 2981 37427
rect 3037 37371 3062 37427
rect 3118 37426 3143 37427
rect 3199 37426 3224 37427
rect 3219 37374 3224 37426
rect 3118 37371 3143 37374
rect 3199 37371 3224 37374
rect 3280 37371 3305 37427
rect 3361 37371 3386 37427
rect 3442 37371 3467 37427
rect 3523 37371 3548 37427
rect 3604 37371 3629 37427
rect 3685 37426 3710 37427
rect 3766 37426 3791 37427
rect 3707 37374 3710 37426
rect 3773 37374 3791 37426
rect 3685 37371 3710 37374
rect 3766 37371 3791 37374
rect 3847 37371 3872 37427
rect 3928 37371 3953 37427
rect 4009 37371 4034 37427
rect 4090 37371 4115 37427
rect 4171 37371 4196 37427
rect 4252 37426 4277 37427
rect 4261 37374 4275 37426
rect 4252 37371 4277 37374
rect 4333 37371 4358 37427
rect 4414 37371 4439 37427
rect 4495 37371 4520 37427
rect 4576 37371 4601 37427
rect 4657 37371 4682 37427
rect 4738 37371 4763 37427
rect 5299 37426 7651 37444
rect 5299 37374 5317 37426
rect 5369 37374 5383 37426
rect 5435 37374 5871 37426
rect 5923 37374 5937 37426
rect 5989 37374 6425 37426
rect 6477 37374 6491 37426
rect 6543 37374 6979 37426
rect 7031 37374 7045 37426
rect 7097 37374 7533 37426
rect 7585 37374 7599 37426
rect 5299 37371 7651 37374
rect 2729 37368 7651 37371
rect 2270 36724 8221 36730
rect 2322 36672 2392 36724
rect 2444 36720 5613 36724
rect 5669 36720 5696 36724
rect 2444 36672 2824 36720
rect 2270 36668 2824 36672
rect 2876 36668 2890 36720
rect 2942 36668 3378 36720
rect 3430 36668 3444 36720
rect 3496 36668 3932 36720
rect 3984 36668 3998 36720
rect 4050 36668 4486 36720
rect 4538 36668 4552 36720
rect 4604 36668 5040 36720
rect 5092 36668 5106 36720
rect 5158 36668 5594 36720
rect 5752 36668 5778 36724
rect 5834 36668 5860 36724
rect 5916 36668 5942 36724
rect 5998 36668 6024 36724
rect 6080 36668 6106 36724
rect 6162 36720 6188 36724
rect 6244 36720 6270 36724
rect 6266 36668 6270 36720
rect 6326 36668 6352 36724
rect 6408 36668 6434 36724
rect 6490 36668 6516 36724
rect 6572 36668 6598 36724
rect 6654 36668 6680 36724
rect 6736 36720 6762 36724
rect 6818 36720 6844 36724
rect 6754 36668 6762 36720
rect 6820 36668 6844 36720
rect 6900 36668 6926 36724
rect 6982 36668 7008 36724
rect 7064 36668 7090 36724
rect 7146 36668 7172 36724
rect 7228 36668 7254 36724
rect 7310 36720 7336 36724
rect 7310 36668 7322 36720
rect 7392 36668 7418 36724
rect 7474 36668 7500 36724
rect 7556 36668 7582 36724
rect 7638 36668 7664 36724
rect 7720 36668 7746 36724
rect 7802 36720 7828 36724
rect 7884 36720 7910 36724
rect 7802 36668 7810 36720
rect 7966 36668 7992 36724
rect 8048 36668 8074 36672
rect 8130 36668 8156 36724
rect 8212 36668 8221 36672
rect 2270 36655 8221 36668
rect 2322 36603 2392 36655
rect 2444 36651 8047 36655
rect 2444 36603 2824 36651
rect 2270 36599 2824 36603
rect 2876 36599 2890 36651
rect 2942 36599 3378 36651
rect 3430 36599 3444 36651
rect 3496 36599 3932 36651
rect 3984 36599 3998 36651
rect 4050 36599 4486 36651
rect 4538 36599 4552 36651
rect 4604 36599 5040 36651
rect 5092 36599 5106 36651
rect 5158 36599 5594 36651
rect 5646 36644 5660 36651
rect 5712 36644 6148 36651
rect 6200 36644 6214 36651
rect 6266 36644 6702 36651
rect 6754 36644 6768 36651
rect 6820 36644 7256 36651
rect 7308 36644 7322 36651
rect 7374 36644 7810 36651
rect 7862 36644 7876 36651
rect 7928 36644 8047 36651
rect 8099 36644 8169 36655
rect 2270 36588 5613 36599
rect 5669 36588 5696 36599
rect 5752 36588 5778 36644
rect 5834 36588 5860 36644
rect 5916 36588 5942 36644
rect 5998 36588 6024 36644
rect 6080 36588 6106 36644
rect 6266 36599 6270 36644
rect 6162 36588 6188 36599
rect 6244 36588 6270 36599
rect 6326 36588 6352 36644
rect 6408 36588 6434 36644
rect 6490 36588 6516 36644
rect 6572 36588 6598 36644
rect 6654 36588 6680 36644
rect 6754 36599 6762 36644
rect 6820 36599 6844 36644
rect 6736 36588 6762 36599
rect 6818 36588 6844 36599
rect 6900 36588 6926 36644
rect 6982 36588 7008 36644
rect 7064 36588 7090 36644
rect 7146 36588 7172 36644
rect 7228 36588 7254 36644
rect 7310 36599 7322 36644
rect 7310 36588 7336 36599
rect 7392 36588 7418 36644
rect 7474 36588 7500 36644
rect 7556 36588 7582 36644
rect 7638 36588 7664 36644
rect 7720 36588 7746 36644
rect 7802 36599 7810 36644
rect 7802 36588 7828 36599
rect 7884 36588 7910 36599
rect 7966 36588 7992 36644
rect 8048 36588 8074 36603
rect 8130 36588 8156 36644
rect 8212 36588 8221 36603
rect 2270 36586 8221 36588
rect 2322 36534 2392 36586
rect 2444 36582 8047 36586
rect 2444 36534 2824 36582
rect 2270 36530 2824 36534
rect 2876 36530 2890 36582
rect 2942 36530 3378 36582
rect 3430 36530 3444 36582
rect 3496 36530 3932 36582
rect 3984 36530 3998 36582
rect 4050 36530 4486 36582
rect 4538 36530 4552 36582
rect 4604 36530 5040 36582
rect 5092 36530 5106 36582
rect 5158 36530 5594 36582
rect 5646 36564 5660 36582
rect 5712 36564 6148 36582
rect 6200 36564 6214 36582
rect 6266 36564 6702 36582
rect 6754 36564 6768 36582
rect 6820 36564 7256 36582
rect 7308 36564 7322 36582
rect 7374 36564 7810 36582
rect 7862 36564 7876 36582
rect 7928 36564 8047 36582
rect 8099 36564 8169 36586
rect 2270 36517 5613 36530
rect 2322 36465 2392 36517
rect 2444 36513 5613 36517
rect 5669 36513 5696 36530
rect 2444 36465 2824 36513
rect 2270 36461 2824 36465
rect 2876 36461 2890 36513
rect 2942 36461 3378 36513
rect 3430 36461 3444 36513
rect 3496 36461 3932 36513
rect 3984 36461 3998 36513
rect 4050 36461 4486 36513
rect 4538 36461 4552 36513
rect 4604 36461 5040 36513
rect 5092 36461 5106 36513
rect 5158 36461 5594 36513
rect 5752 36508 5778 36564
rect 5834 36508 5860 36564
rect 5916 36508 5942 36564
rect 5998 36508 6024 36564
rect 6080 36508 6106 36564
rect 6266 36530 6270 36564
rect 6162 36513 6188 36530
rect 6244 36513 6270 36530
rect 6266 36508 6270 36513
rect 6326 36508 6352 36564
rect 6408 36508 6434 36564
rect 6490 36508 6516 36564
rect 6572 36508 6598 36564
rect 6654 36508 6680 36564
rect 6754 36530 6762 36564
rect 6820 36530 6844 36564
rect 6736 36513 6762 36530
rect 6818 36513 6844 36530
rect 6754 36508 6762 36513
rect 6820 36508 6844 36513
rect 6900 36508 6926 36564
rect 6982 36508 7008 36564
rect 7064 36508 7090 36564
rect 7146 36508 7172 36564
rect 7228 36508 7254 36564
rect 7310 36530 7322 36564
rect 7310 36513 7336 36530
rect 7310 36508 7322 36513
rect 7392 36508 7418 36564
rect 7474 36508 7500 36564
rect 7556 36508 7582 36564
rect 7638 36508 7664 36564
rect 7720 36508 7746 36564
rect 7802 36530 7810 36564
rect 7802 36513 7828 36530
rect 7884 36513 7910 36530
rect 7802 36508 7810 36513
rect 7966 36508 7992 36564
rect 8048 36517 8074 36534
rect 8130 36508 8156 36564
rect 8212 36517 8221 36534
rect 5646 36484 5660 36508
rect 5712 36484 6148 36508
rect 6200 36484 6214 36508
rect 6266 36484 6702 36508
rect 6754 36484 6768 36508
rect 6820 36484 7256 36508
rect 7308 36484 7322 36508
rect 7374 36484 7810 36508
rect 7862 36484 7876 36508
rect 7928 36484 8047 36508
rect 8099 36484 8169 36508
rect 2270 36448 5613 36461
rect 2322 36396 2392 36448
rect 2444 36444 5613 36448
rect 5669 36444 5696 36461
rect 2444 36396 2824 36444
rect 2270 36392 2824 36396
rect 2876 36392 2890 36444
rect 2942 36392 3378 36444
rect 3430 36392 3444 36444
rect 3496 36392 3932 36444
rect 3984 36392 3998 36444
rect 4050 36392 4486 36444
rect 4538 36392 4552 36444
rect 4604 36392 5040 36444
rect 5092 36392 5106 36444
rect 5158 36392 5594 36444
rect 5752 36428 5778 36484
rect 5834 36428 5860 36484
rect 5916 36428 5942 36484
rect 5998 36428 6024 36484
rect 6080 36428 6106 36484
rect 6266 36461 6270 36484
rect 6162 36444 6188 36461
rect 6244 36444 6270 36461
rect 6266 36428 6270 36444
rect 6326 36428 6352 36484
rect 6408 36428 6434 36484
rect 6490 36428 6516 36484
rect 6572 36428 6598 36484
rect 6654 36428 6680 36484
rect 6754 36461 6762 36484
rect 6820 36461 6844 36484
rect 6736 36444 6762 36461
rect 6818 36444 6844 36461
rect 6754 36428 6762 36444
rect 6820 36428 6844 36444
rect 6900 36428 6926 36484
rect 6982 36428 7008 36484
rect 7064 36428 7090 36484
rect 7146 36428 7172 36484
rect 7228 36428 7254 36484
rect 7310 36461 7322 36484
rect 7310 36444 7336 36461
rect 7310 36428 7322 36444
rect 7392 36428 7418 36484
rect 7474 36428 7500 36484
rect 7556 36428 7582 36484
rect 7638 36428 7664 36484
rect 7720 36428 7746 36484
rect 7802 36461 7810 36484
rect 7802 36444 7828 36461
rect 7884 36444 7910 36461
rect 7802 36428 7810 36444
rect 7966 36428 7992 36484
rect 8048 36448 8074 36465
rect 8130 36428 8156 36484
rect 8212 36448 8221 36465
rect 5646 36404 5660 36428
rect 5712 36404 6148 36428
rect 6200 36404 6214 36428
rect 6266 36404 6702 36428
rect 6754 36404 6768 36428
rect 6820 36404 7256 36428
rect 7308 36404 7322 36428
rect 7374 36404 7810 36428
rect 7862 36404 7876 36428
rect 7928 36404 8047 36428
rect 8099 36404 8169 36428
rect 2270 36378 5613 36392
rect 2322 36326 2392 36378
rect 2444 36375 5613 36378
rect 5669 36375 5696 36392
rect 2444 36326 2824 36375
rect 2270 36323 2824 36326
rect 2876 36323 2890 36375
rect 2942 36323 3378 36375
rect 3430 36323 3444 36375
rect 3496 36323 3932 36375
rect 3984 36323 3998 36375
rect 4050 36323 4486 36375
rect 4538 36323 4552 36375
rect 4604 36323 5040 36375
rect 5092 36323 5106 36375
rect 5158 36323 5594 36375
rect 5752 36348 5778 36404
rect 5834 36348 5860 36404
rect 5916 36348 5942 36404
rect 5998 36348 6024 36404
rect 6080 36348 6106 36404
rect 6266 36392 6270 36404
rect 6162 36375 6188 36392
rect 6244 36375 6270 36392
rect 6266 36348 6270 36375
rect 6326 36348 6352 36404
rect 6408 36348 6434 36404
rect 6490 36348 6516 36404
rect 6572 36348 6598 36404
rect 6654 36348 6680 36404
rect 6754 36392 6762 36404
rect 6820 36392 6844 36404
rect 6736 36375 6762 36392
rect 6818 36375 6844 36392
rect 6754 36348 6762 36375
rect 6820 36348 6844 36375
rect 6900 36348 6926 36404
rect 6982 36348 7008 36404
rect 7064 36348 7090 36404
rect 7146 36348 7172 36404
rect 7228 36348 7254 36404
rect 7310 36392 7322 36404
rect 7310 36375 7336 36392
rect 7310 36348 7322 36375
rect 7392 36348 7418 36404
rect 7474 36348 7500 36404
rect 7556 36348 7582 36404
rect 7638 36348 7664 36404
rect 7720 36348 7746 36404
rect 7802 36392 7810 36404
rect 7802 36375 7828 36392
rect 7884 36375 7910 36392
rect 7802 36348 7810 36375
rect 7966 36348 7992 36404
rect 8048 36378 8074 36396
rect 8130 36348 8156 36404
rect 8212 36378 8221 36396
rect 5646 36324 5660 36348
rect 5712 36324 6148 36348
rect 6200 36324 6214 36348
rect 6266 36324 6702 36348
rect 6754 36324 6768 36348
rect 6820 36324 7256 36348
rect 7308 36324 7322 36348
rect 7374 36324 7810 36348
rect 7862 36324 7876 36348
rect 7928 36326 8047 36348
rect 8099 36326 8169 36348
rect 7928 36324 8221 36326
rect 2270 36308 5613 36323
rect 2322 36256 2392 36308
rect 2444 36306 5613 36308
rect 5669 36306 5696 36323
rect 2444 36256 2824 36306
rect 2270 36254 2824 36256
rect 2876 36254 2890 36306
rect 2942 36254 3378 36306
rect 3430 36254 3444 36306
rect 3496 36254 3932 36306
rect 3984 36254 3998 36306
rect 4050 36254 4486 36306
rect 4538 36254 4552 36306
rect 4604 36254 5040 36306
rect 5092 36254 5106 36306
rect 5158 36254 5594 36306
rect 5752 36268 5778 36324
rect 5834 36268 5860 36324
rect 5916 36268 5942 36324
rect 5998 36268 6024 36324
rect 6080 36268 6106 36324
rect 6266 36323 6270 36324
rect 6162 36306 6188 36323
rect 6244 36306 6270 36323
rect 6266 36268 6270 36306
rect 6326 36268 6352 36324
rect 6408 36268 6434 36324
rect 6490 36268 6516 36324
rect 6572 36268 6598 36324
rect 6654 36268 6680 36324
rect 6754 36323 6762 36324
rect 6820 36323 6844 36324
rect 6736 36306 6762 36323
rect 6818 36306 6844 36323
rect 6754 36268 6762 36306
rect 6820 36268 6844 36306
rect 6900 36268 6926 36324
rect 6982 36268 7008 36324
rect 7064 36268 7090 36324
rect 7146 36268 7172 36324
rect 7228 36268 7254 36324
rect 7310 36323 7322 36324
rect 7310 36306 7336 36323
rect 7310 36268 7322 36306
rect 7392 36268 7418 36324
rect 7474 36268 7500 36324
rect 7556 36268 7582 36324
rect 7638 36268 7664 36324
rect 7720 36268 7746 36324
rect 7802 36323 7810 36324
rect 7802 36306 7828 36323
rect 7884 36306 7910 36323
rect 7802 36268 7810 36306
rect 7966 36268 7992 36324
rect 8048 36308 8074 36324
rect 8130 36268 8156 36324
rect 8212 36308 8221 36324
rect 5646 36254 5660 36268
rect 5712 36254 6148 36268
rect 6200 36254 6214 36268
rect 6266 36254 6702 36268
rect 6754 36254 6768 36268
rect 6820 36254 7256 36268
rect 7308 36254 7322 36268
rect 7374 36254 7810 36268
rect 7862 36254 7876 36268
rect 7928 36256 8047 36268
rect 8099 36256 8169 36268
rect 7928 36254 8221 36256
rect 2270 36244 8221 36254
rect 2270 36238 5613 36244
rect 2322 36186 2392 36238
rect 2444 36236 5613 36238
rect 5669 36236 5696 36244
rect 2444 36186 2824 36236
rect 2270 36184 2824 36186
rect 2876 36184 2890 36236
rect 2942 36184 3378 36236
rect 3430 36184 3444 36236
rect 3496 36184 3932 36236
rect 3984 36184 3998 36236
rect 4050 36184 4486 36236
rect 4538 36184 4552 36236
rect 4604 36184 5040 36236
rect 5092 36184 5106 36236
rect 5158 36184 5594 36236
rect 5752 36188 5778 36244
rect 5834 36188 5860 36244
rect 5916 36188 5942 36244
rect 5998 36188 6024 36244
rect 6080 36188 6106 36244
rect 6162 36236 6188 36244
rect 6244 36236 6270 36244
rect 6266 36188 6270 36236
rect 6326 36188 6352 36244
rect 6408 36188 6434 36244
rect 6490 36188 6516 36244
rect 6572 36188 6598 36244
rect 6654 36188 6680 36244
rect 6736 36236 6762 36244
rect 6818 36236 6844 36244
rect 6754 36188 6762 36236
rect 6820 36188 6844 36236
rect 6900 36188 6926 36244
rect 6982 36188 7008 36244
rect 7064 36188 7090 36244
rect 7146 36188 7172 36244
rect 7228 36188 7254 36244
rect 7310 36236 7336 36244
rect 7310 36188 7322 36236
rect 7392 36188 7418 36244
rect 7474 36188 7500 36244
rect 7556 36188 7582 36244
rect 7638 36188 7664 36244
rect 7720 36188 7746 36244
rect 7802 36236 7828 36244
rect 7884 36236 7910 36244
rect 7802 36188 7810 36236
rect 7966 36188 7992 36244
rect 8048 36238 8074 36244
rect 8130 36188 8156 36244
rect 8212 36238 8221 36244
rect 5646 36184 5660 36188
rect 5712 36184 6148 36188
rect 6200 36184 6214 36188
rect 6266 36184 6702 36188
rect 6754 36184 6768 36188
rect 6820 36184 7256 36188
rect 7308 36184 7322 36188
rect 7374 36184 7810 36188
rect 7862 36184 7876 36188
rect 7928 36186 8047 36188
rect 8099 36186 8169 36188
rect 7928 36184 8221 36186
rect 2270 36168 8221 36184
rect 2322 36116 2392 36168
rect 2444 36166 8047 36168
rect 2444 36116 2824 36166
rect 2270 36114 2824 36116
rect 2876 36114 2890 36166
rect 2942 36114 3378 36166
rect 3430 36114 3444 36166
rect 3496 36114 3932 36166
rect 3984 36114 3998 36166
rect 4050 36114 4486 36166
rect 4538 36114 4552 36166
rect 4604 36114 5040 36166
rect 5092 36114 5106 36166
rect 5158 36114 5594 36166
rect 5646 36164 5660 36166
rect 5712 36164 6148 36166
rect 6200 36164 6214 36166
rect 6266 36164 6702 36166
rect 6754 36164 6768 36166
rect 6820 36164 7256 36166
rect 7308 36164 7322 36166
rect 7374 36164 7810 36166
rect 7862 36164 7876 36166
rect 7928 36164 8047 36166
rect 8099 36164 8169 36168
rect 2270 36108 5613 36114
rect 5669 36108 5696 36114
rect 5752 36108 5778 36164
rect 5834 36108 5860 36164
rect 5916 36108 5942 36164
rect 5998 36108 6024 36164
rect 6080 36108 6106 36164
rect 6266 36114 6270 36164
rect 6162 36108 6188 36114
rect 6244 36108 6270 36114
rect 6326 36108 6352 36164
rect 6408 36108 6434 36164
rect 6490 36108 6516 36164
rect 6572 36108 6598 36164
rect 6654 36108 6680 36164
rect 6754 36114 6762 36164
rect 6820 36114 6844 36164
rect 6736 36108 6762 36114
rect 6818 36108 6844 36114
rect 6900 36108 6926 36164
rect 6982 36108 7008 36164
rect 7064 36108 7090 36164
rect 7146 36108 7172 36164
rect 7228 36108 7254 36164
rect 7310 36114 7322 36164
rect 7310 36108 7336 36114
rect 7392 36108 7418 36164
rect 7474 36108 7500 36164
rect 7556 36108 7582 36164
rect 7638 36108 7664 36164
rect 7720 36108 7746 36164
rect 7802 36114 7810 36164
rect 7802 36108 7828 36114
rect 7884 36108 7910 36114
rect 7966 36108 7992 36164
rect 8048 36108 8074 36116
rect 8130 36108 8156 36164
rect 8212 36108 8221 36116
rect 2724 35987 7651 35988
rect 2724 35931 2733 35987
rect 2789 35931 2814 35987
rect 2870 35931 2895 35987
rect 2951 35931 2976 35987
rect 3032 35931 3057 35987
rect 3113 35982 3138 35987
rect 3194 35982 3219 35987
rect 3275 35931 3300 35987
rect 3356 35931 3381 35987
rect 3437 35931 3462 35987
rect 3518 35931 3543 35987
rect 3599 35931 3624 35987
rect 3680 35982 3705 35987
rect 3761 35982 3786 35987
rect 3773 35931 3786 35982
rect 3842 35931 3867 35987
rect 3923 35931 3948 35987
rect 4004 35931 4029 35987
rect 4085 35931 4110 35987
rect 4166 35931 4191 35987
rect 4247 35982 4272 35987
rect 4261 35931 4272 35982
rect 4328 35931 4353 35987
rect 4409 35931 4434 35987
rect 4490 35931 4515 35987
rect 4571 35931 4596 35987
rect 4652 35931 4677 35987
rect 4733 35931 4758 35987
rect 4814 35982 4839 35987
rect 2724 35930 3101 35931
rect 3153 35930 3167 35931
rect 3219 35930 3655 35931
rect 3707 35930 3721 35931
rect 3773 35930 4209 35931
rect 4261 35930 4275 35931
rect 4327 35930 4763 35931
rect 4815 35930 4829 35982
rect 4895 35931 4920 35987
rect 4976 35931 5001 35987
rect 5057 35931 5082 35987
rect 5138 35931 5163 35987
rect 4881 35930 5163 35931
rect 2724 35913 5163 35930
rect 2724 35907 3101 35913
rect 3153 35907 3167 35913
rect 3219 35907 3655 35913
rect 3707 35907 3721 35913
rect 3773 35907 4209 35913
rect 4261 35907 4275 35913
rect 4327 35907 4763 35913
rect 2724 35851 2733 35907
rect 2789 35851 2814 35907
rect 2870 35851 2895 35907
rect 2951 35851 2976 35907
rect 3032 35851 3057 35907
rect 3113 35851 3138 35861
rect 3194 35851 3219 35861
rect 3275 35851 3300 35907
rect 3356 35851 3381 35907
rect 3437 35851 3462 35907
rect 3518 35851 3543 35907
rect 3599 35851 3624 35907
rect 3773 35861 3786 35907
rect 3680 35851 3705 35861
rect 3761 35851 3786 35861
rect 3842 35851 3867 35907
rect 3923 35851 3948 35907
rect 4004 35851 4029 35907
rect 4085 35851 4110 35907
rect 4166 35851 4191 35907
rect 4261 35861 4272 35907
rect 4247 35851 4272 35861
rect 4328 35851 4353 35907
rect 4409 35851 4434 35907
rect 4490 35851 4515 35907
rect 4571 35851 4596 35907
rect 4652 35851 4677 35907
rect 4733 35851 4758 35907
rect 4815 35861 4829 35913
rect 4881 35907 5163 35913
rect 4814 35851 4839 35861
rect 4895 35851 4920 35907
rect 4976 35851 5001 35907
rect 5057 35851 5082 35907
rect 5138 35851 5163 35907
rect 2724 35844 5163 35851
rect 2724 35827 3101 35844
rect 3153 35827 3167 35844
rect 3219 35827 3655 35844
rect 3707 35827 3721 35844
rect 3773 35827 4209 35844
rect 4261 35827 4275 35844
rect 4327 35827 4763 35844
rect 2724 35771 2733 35827
rect 2789 35771 2814 35827
rect 2870 35771 2895 35827
rect 2951 35771 2976 35827
rect 3032 35771 3057 35827
rect 3113 35775 3138 35792
rect 3194 35775 3219 35792
rect 3275 35771 3300 35827
rect 3356 35771 3381 35827
rect 3437 35771 3462 35827
rect 3518 35771 3543 35827
rect 3599 35771 3624 35827
rect 3773 35792 3786 35827
rect 3680 35775 3705 35792
rect 3761 35775 3786 35792
rect 3773 35771 3786 35775
rect 3842 35771 3867 35827
rect 3923 35771 3948 35827
rect 4004 35771 4029 35827
rect 4085 35771 4110 35827
rect 4166 35771 4191 35827
rect 4261 35792 4272 35827
rect 4247 35775 4272 35792
rect 4261 35771 4272 35775
rect 4328 35771 4353 35827
rect 4409 35771 4434 35827
rect 4490 35771 4515 35827
rect 4571 35771 4596 35827
rect 4652 35771 4677 35827
rect 4733 35771 4758 35827
rect 4815 35792 4829 35844
rect 4881 35827 5163 35844
rect 4814 35775 4839 35792
rect 2724 35747 3101 35771
rect 3153 35747 3167 35771
rect 3219 35747 3655 35771
rect 3707 35747 3721 35771
rect 3773 35747 4209 35771
rect 4261 35747 4275 35771
rect 4327 35747 4763 35771
rect 2724 35691 2733 35747
rect 2789 35691 2814 35747
rect 2870 35691 2895 35747
rect 2951 35691 2976 35747
rect 3032 35691 3057 35747
rect 3113 35706 3138 35723
rect 3194 35706 3219 35723
rect 3275 35691 3300 35747
rect 3356 35691 3381 35747
rect 3437 35691 3462 35747
rect 3518 35691 3543 35747
rect 3599 35691 3624 35747
rect 3773 35723 3786 35747
rect 3680 35706 3705 35723
rect 3761 35706 3786 35723
rect 3773 35691 3786 35706
rect 3842 35691 3867 35747
rect 3923 35691 3948 35747
rect 4004 35691 4029 35747
rect 4085 35691 4110 35747
rect 4166 35691 4191 35747
rect 4261 35723 4272 35747
rect 4247 35706 4272 35723
rect 4261 35691 4272 35706
rect 4328 35691 4353 35747
rect 4409 35691 4434 35747
rect 4490 35691 4515 35747
rect 4571 35691 4596 35747
rect 4652 35691 4677 35747
rect 4733 35691 4758 35747
rect 4815 35723 4829 35775
rect 4895 35771 4920 35827
rect 4976 35771 5001 35827
rect 5057 35771 5082 35827
rect 5138 35771 5163 35827
rect 4881 35747 5163 35771
rect 4814 35706 4839 35723
rect 2724 35667 3101 35691
rect 3153 35667 3167 35691
rect 3219 35667 3655 35691
rect 3707 35667 3721 35691
rect 3773 35667 4209 35691
rect 4261 35667 4275 35691
rect 4327 35667 4763 35691
rect 2724 35611 2733 35667
rect 2789 35611 2814 35667
rect 2870 35611 2895 35667
rect 2951 35611 2976 35667
rect 3032 35611 3057 35667
rect 3113 35636 3138 35654
rect 3194 35636 3219 35654
rect 3275 35611 3300 35667
rect 3356 35611 3381 35667
rect 3437 35611 3462 35667
rect 3518 35611 3543 35667
rect 3599 35611 3624 35667
rect 3773 35654 3786 35667
rect 3680 35636 3705 35654
rect 3761 35636 3786 35654
rect 3773 35611 3786 35636
rect 3842 35611 3867 35667
rect 3923 35611 3948 35667
rect 4004 35611 4029 35667
rect 4085 35611 4110 35667
rect 4166 35611 4191 35667
rect 4261 35654 4272 35667
rect 4247 35636 4272 35654
rect 4261 35611 4272 35636
rect 4328 35611 4353 35667
rect 4409 35611 4434 35667
rect 4490 35611 4515 35667
rect 4571 35611 4596 35667
rect 4652 35611 4677 35667
rect 4733 35611 4758 35667
rect 4815 35654 4829 35706
rect 4895 35691 4920 35747
rect 4976 35691 5001 35747
rect 5057 35691 5082 35747
rect 5138 35691 5163 35747
rect 4881 35667 5163 35691
rect 4814 35636 4839 35654
rect 2724 35587 3101 35611
rect 3153 35587 3167 35611
rect 3219 35587 3655 35611
rect 3707 35587 3721 35611
rect 3773 35587 4209 35611
rect 4261 35587 4275 35611
rect 4327 35587 4763 35611
rect 2724 35531 2733 35587
rect 2789 35531 2814 35587
rect 2870 35531 2895 35587
rect 2951 35531 2976 35587
rect 3032 35531 3057 35587
rect 3113 35566 3138 35584
rect 3194 35566 3219 35584
rect 3275 35531 3300 35587
rect 3356 35531 3381 35587
rect 3437 35531 3462 35587
rect 3518 35531 3543 35587
rect 3599 35531 3624 35587
rect 3773 35584 3786 35587
rect 3680 35566 3705 35584
rect 3761 35566 3786 35584
rect 3773 35531 3786 35566
rect 3842 35531 3867 35587
rect 3923 35531 3948 35587
rect 4004 35531 4029 35587
rect 4085 35531 4110 35587
rect 4166 35531 4191 35587
rect 4261 35584 4272 35587
rect 4247 35566 4272 35584
rect 4261 35531 4272 35566
rect 4328 35531 4353 35587
rect 4409 35531 4434 35587
rect 4490 35531 4515 35587
rect 4571 35531 4596 35587
rect 4652 35531 4677 35587
rect 4733 35531 4758 35587
rect 4815 35584 4829 35636
rect 4895 35611 4920 35667
rect 4976 35611 5001 35667
rect 5057 35611 5082 35667
rect 5138 35611 5163 35667
rect 4881 35587 5163 35611
rect 4814 35566 4839 35584
rect 2724 35514 3101 35531
rect 3153 35514 3167 35531
rect 3219 35514 3655 35531
rect 3707 35514 3721 35531
rect 3773 35514 4209 35531
rect 4261 35514 4275 35531
rect 4327 35514 4763 35531
rect 4815 35514 4829 35566
rect 4895 35531 4920 35587
rect 4976 35531 5001 35587
rect 5057 35531 5082 35587
rect 5138 35531 5163 35587
rect 4881 35514 5163 35531
rect 2724 35507 5163 35514
rect 2724 35451 2733 35507
rect 2789 35451 2814 35507
rect 2870 35451 2895 35507
rect 2951 35451 2976 35507
rect 3032 35451 3057 35507
rect 3113 35496 3138 35507
rect 3194 35496 3219 35507
rect 3275 35451 3300 35507
rect 3356 35451 3381 35507
rect 3437 35451 3462 35507
rect 3518 35451 3543 35507
rect 3599 35451 3624 35507
rect 3680 35496 3705 35507
rect 3761 35496 3786 35507
rect 3773 35451 3786 35496
rect 3842 35451 3867 35507
rect 3923 35451 3948 35507
rect 4004 35451 4029 35507
rect 4085 35451 4110 35507
rect 4166 35451 4191 35507
rect 4247 35496 4272 35507
rect 4261 35451 4272 35496
rect 4328 35451 4353 35507
rect 4409 35451 4434 35507
rect 4490 35451 4515 35507
rect 4571 35451 4596 35507
rect 4652 35451 4677 35507
rect 4733 35451 4758 35507
rect 4814 35496 4839 35507
rect 2724 35444 3101 35451
rect 3153 35444 3167 35451
rect 3219 35444 3655 35451
rect 3707 35444 3721 35451
rect 3773 35444 4209 35451
rect 4261 35444 4275 35451
rect 4327 35444 4763 35451
rect 4815 35444 4829 35496
rect 4895 35451 4920 35507
rect 4976 35451 5001 35507
rect 5057 35451 5082 35507
rect 5138 35451 5163 35507
rect 4881 35444 5163 35451
rect 2724 35427 5163 35444
rect 2724 35371 2733 35427
rect 2789 35371 2814 35427
rect 2870 35371 2895 35427
rect 2951 35371 2976 35427
rect 3032 35371 3057 35427
rect 3113 35426 3138 35427
rect 3194 35426 3219 35427
rect 3113 35371 3138 35374
rect 3194 35371 3219 35374
rect 3275 35371 3300 35427
rect 3356 35371 3381 35427
rect 3437 35371 3462 35427
rect 3518 35371 3543 35427
rect 3599 35371 3624 35427
rect 3680 35426 3705 35427
rect 3761 35426 3786 35427
rect 3773 35374 3786 35426
rect 3680 35371 3705 35374
rect 3761 35371 3786 35374
rect 3842 35371 3867 35427
rect 3923 35371 3948 35427
rect 4004 35371 4029 35427
rect 4085 35371 4110 35427
rect 4166 35371 4191 35427
rect 4247 35426 4272 35427
rect 4261 35374 4272 35426
rect 4247 35371 4272 35374
rect 4328 35371 4353 35427
rect 4409 35371 4434 35427
rect 4490 35371 4515 35427
rect 4571 35371 4596 35427
rect 4652 35371 4677 35427
rect 4733 35371 4758 35427
rect 4814 35426 4839 35427
rect 4815 35374 4829 35426
rect 4814 35371 4839 35374
rect 4895 35371 4920 35427
rect 4976 35371 5001 35427
rect 5057 35371 5082 35427
rect 5138 35371 5163 35427
rect 5299 35982 7651 35987
rect 5299 35930 5317 35982
rect 5369 35930 5383 35982
rect 5435 35930 5871 35982
rect 5923 35930 5937 35982
rect 5989 35930 6425 35982
rect 6477 35930 6491 35982
rect 6543 35930 6979 35982
rect 7031 35930 7045 35982
rect 7097 35930 7533 35982
rect 7585 35930 7599 35982
rect 5299 35913 7651 35930
rect 5299 35861 5317 35913
rect 5369 35861 5383 35913
rect 5435 35861 5871 35913
rect 5923 35861 5937 35913
rect 5989 35861 6425 35913
rect 6477 35861 6491 35913
rect 6543 35861 6979 35913
rect 7031 35861 7045 35913
rect 7097 35861 7533 35913
rect 7585 35861 7599 35913
rect 5299 35844 7651 35861
rect 5299 35792 5317 35844
rect 5369 35792 5383 35844
rect 5435 35792 5871 35844
rect 5923 35792 5937 35844
rect 5989 35792 6425 35844
rect 6477 35792 6491 35844
rect 6543 35792 6979 35844
rect 7031 35792 7045 35844
rect 7097 35792 7533 35844
rect 7585 35792 7599 35844
rect 5299 35775 7651 35792
rect 5299 35723 5317 35775
rect 5369 35723 5383 35775
rect 5435 35723 5871 35775
rect 5923 35723 5937 35775
rect 5989 35723 6425 35775
rect 6477 35723 6491 35775
rect 6543 35723 6979 35775
rect 7031 35723 7045 35775
rect 7097 35723 7533 35775
rect 7585 35723 7599 35775
rect 5299 35706 7651 35723
rect 5299 35654 5317 35706
rect 5369 35654 5383 35706
rect 5435 35654 5871 35706
rect 5923 35654 5937 35706
rect 5989 35654 6425 35706
rect 6477 35654 6491 35706
rect 6543 35654 6979 35706
rect 7031 35654 7045 35706
rect 7097 35654 7533 35706
rect 7585 35654 7599 35706
rect 5299 35636 7651 35654
rect 5299 35584 5317 35636
rect 5369 35584 5383 35636
rect 5435 35584 5871 35636
rect 5923 35584 5937 35636
rect 5989 35584 6425 35636
rect 6477 35584 6491 35636
rect 6543 35584 6979 35636
rect 7031 35584 7045 35636
rect 7097 35584 7533 35636
rect 7585 35584 7599 35636
rect 5299 35566 7651 35584
rect 5299 35514 5317 35566
rect 5369 35514 5383 35566
rect 5435 35514 5871 35566
rect 5923 35514 5937 35566
rect 5989 35514 6425 35566
rect 6477 35514 6491 35566
rect 6543 35514 6979 35566
rect 7031 35514 7045 35566
rect 7097 35514 7533 35566
rect 7585 35514 7599 35566
rect 5299 35496 7651 35514
rect 5299 35444 5317 35496
rect 5369 35444 5383 35496
rect 5435 35444 5871 35496
rect 5923 35444 5937 35496
rect 5989 35444 6425 35496
rect 6477 35444 6491 35496
rect 6543 35444 6979 35496
rect 7031 35444 7045 35496
rect 7097 35444 7533 35496
rect 7585 35444 7599 35496
rect 5299 35426 7651 35444
rect 5299 35374 5317 35426
rect 5369 35374 5383 35426
rect 5435 35374 5871 35426
rect 5923 35374 5937 35426
rect 5989 35374 6425 35426
rect 6477 35374 6491 35426
rect 6543 35374 6979 35426
rect 7031 35374 7045 35426
rect 7097 35374 7533 35426
rect 7585 35374 7599 35426
rect 5299 35371 7651 35374
rect 2724 35368 7651 35371
rect 2270 34724 8222 34730
rect 2322 34672 2392 34724
rect 2444 34720 5613 34724
rect 5669 34720 5696 34724
rect 2444 34672 2824 34720
rect 2270 34668 2824 34672
rect 2876 34668 2890 34720
rect 2942 34668 3378 34720
rect 3430 34668 3444 34720
rect 3496 34668 3932 34720
rect 3984 34668 3998 34720
rect 4050 34668 4486 34720
rect 4538 34668 4552 34720
rect 4604 34668 5040 34720
rect 5092 34668 5106 34720
rect 5158 34668 5594 34720
rect 5752 34668 5779 34724
rect 5835 34668 5861 34724
rect 5917 34668 5943 34724
rect 5999 34668 6025 34724
rect 6081 34668 6107 34724
rect 6163 34720 6189 34724
rect 6245 34720 6271 34724
rect 6266 34668 6271 34720
rect 6327 34668 6353 34724
rect 6409 34668 6435 34724
rect 6491 34668 6517 34724
rect 6573 34668 6599 34724
rect 6655 34668 6681 34724
rect 6737 34720 6763 34724
rect 6819 34720 6845 34724
rect 6754 34668 6763 34720
rect 6820 34668 6845 34720
rect 6901 34668 6927 34724
rect 6983 34668 7009 34724
rect 7065 34668 7091 34724
rect 7147 34668 7173 34724
rect 7229 34668 7255 34724
rect 7311 34720 7337 34724
rect 7311 34668 7322 34720
rect 7393 34668 7419 34724
rect 7475 34668 7501 34724
rect 7557 34668 7583 34724
rect 7639 34668 7665 34724
rect 7721 34668 7747 34724
rect 7803 34720 7829 34724
rect 7885 34720 7911 34724
rect 7803 34668 7810 34720
rect 7967 34668 7993 34724
rect 8049 34668 8075 34672
rect 8131 34668 8157 34724
rect 8221 34672 8222 34724
rect 8213 34668 8222 34672
rect 2270 34655 8222 34668
rect 2322 34603 2392 34655
rect 2444 34651 8047 34655
rect 2444 34603 2824 34651
rect 2270 34599 2824 34603
rect 2876 34599 2890 34651
rect 2942 34599 3378 34651
rect 3430 34599 3444 34651
rect 3496 34599 3932 34651
rect 3984 34599 3998 34651
rect 4050 34599 4486 34651
rect 4538 34599 4552 34651
rect 4604 34599 5040 34651
rect 5092 34599 5106 34651
rect 5158 34599 5594 34651
rect 5646 34644 5660 34651
rect 5712 34644 6148 34651
rect 6200 34644 6214 34651
rect 6266 34644 6702 34651
rect 6754 34644 6768 34651
rect 6820 34644 7256 34651
rect 7308 34644 7322 34651
rect 7374 34644 7810 34651
rect 7862 34644 7876 34651
rect 7928 34644 8047 34651
rect 8099 34644 8169 34655
rect 2270 34588 5613 34599
rect 5669 34588 5696 34599
rect 5752 34588 5779 34644
rect 5835 34588 5861 34644
rect 5917 34588 5943 34644
rect 5999 34588 6025 34644
rect 6081 34588 6107 34644
rect 6266 34599 6271 34644
rect 6163 34588 6189 34599
rect 6245 34588 6271 34599
rect 6327 34588 6353 34644
rect 6409 34588 6435 34644
rect 6491 34588 6517 34644
rect 6573 34588 6599 34644
rect 6655 34588 6681 34644
rect 6754 34599 6763 34644
rect 6820 34599 6845 34644
rect 6737 34588 6763 34599
rect 6819 34588 6845 34599
rect 6901 34588 6927 34644
rect 6983 34588 7009 34644
rect 7065 34588 7091 34644
rect 7147 34588 7173 34644
rect 7229 34588 7255 34644
rect 7311 34599 7322 34644
rect 7311 34588 7337 34599
rect 7393 34588 7419 34644
rect 7475 34588 7501 34644
rect 7557 34588 7583 34644
rect 7639 34588 7665 34644
rect 7721 34588 7747 34644
rect 7803 34599 7810 34644
rect 7803 34588 7829 34599
rect 7885 34588 7911 34599
rect 7967 34588 7993 34644
rect 8049 34588 8075 34603
rect 8131 34588 8157 34644
rect 8221 34603 8222 34655
rect 8213 34588 8222 34603
rect 2270 34586 8222 34588
rect 2322 34534 2392 34586
rect 2444 34582 8047 34586
rect 2444 34534 2824 34582
rect 2270 34530 2824 34534
rect 2876 34530 2890 34582
rect 2942 34530 3378 34582
rect 3430 34530 3444 34582
rect 3496 34530 3932 34582
rect 3984 34530 3998 34582
rect 4050 34530 4486 34582
rect 4538 34530 4552 34582
rect 4604 34530 5040 34582
rect 5092 34530 5106 34582
rect 5158 34530 5594 34582
rect 5646 34564 5660 34582
rect 5712 34564 6148 34582
rect 6200 34564 6214 34582
rect 6266 34564 6702 34582
rect 6754 34564 6768 34582
rect 6820 34564 7256 34582
rect 7308 34564 7322 34582
rect 7374 34564 7810 34582
rect 7862 34564 7876 34582
rect 7928 34564 8047 34582
rect 8099 34564 8169 34586
rect 2270 34517 5613 34530
rect 2322 34465 2392 34517
rect 2444 34513 5613 34517
rect 5669 34513 5696 34530
rect 2444 34465 2824 34513
rect 2270 34461 2824 34465
rect 2876 34461 2890 34513
rect 2942 34461 3378 34513
rect 3430 34461 3444 34513
rect 3496 34461 3932 34513
rect 3984 34461 3998 34513
rect 4050 34461 4486 34513
rect 4538 34461 4552 34513
rect 4604 34461 5040 34513
rect 5092 34461 5106 34513
rect 5158 34461 5594 34513
rect 5752 34508 5779 34564
rect 5835 34508 5861 34564
rect 5917 34508 5943 34564
rect 5999 34508 6025 34564
rect 6081 34508 6107 34564
rect 6266 34530 6271 34564
rect 6163 34513 6189 34530
rect 6245 34513 6271 34530
rect 6266 34508 6271 34513
rect 6327 34508 6353 34564
rect 6409 34508 6435 34564
rect 6491 34508 6517 34564
rect 6573 34508 6599 34564
rect 6655 34508 6681 34564
rect 6754 34530 6763 34564
rect 6820 34530 6845 34564
rect 6737 34513 6763 34530
rect 6819 34513 6845 34530
rect 6754 34508 6763 34513
rect 6820 34508 6845 34513
rect 6901 34508 6927 34564
rect 6983 34508 7009 34564
rect 7065 34508 7091 34564
rect 7147 34508 7173 34564
rect 7229 34508 7255 34564
rect 7311 34530 7322 34564
rect 7311 34513 7337 34530
rect 7311 34508 7322 34513
rect 7393 34508 7419 34564
rect 7475 34508 7501 34564
rect 7557 34508 7583 34564
rect 7639 34508 7665 34564
rect 7721 34508 7747 34564
rect 7803 34530 7810 34564
rect 7803 34513 7829 34530
rect 7885 34513 7911 34530
rect 7803 34508 7810 34513
rect 7967 34508 7993 34564
rect 8049 34517 8075 34534
rect 8131 34508 8157 34564
rect 8221 34534 8222 34586
rect 8213 34517 8222 34534
rect 5646 34484 5660 34508
rect 5712 34484 6148 34508
rect 6200 34484 6214 34508
rect 6266 34484 6702 34508
rect 6754 34484 6768 34508
rect 6820 34484 7256 34508
rect 7308 34484 7322 34508
rect 7374 34484 7810 34508
rect 7862 34484 7876 34508
rect 7928 34484 8047 34508
rect 8099 34484 8169 34508
rect 2270 34448 5613 34461
rect 2322 34396 2392 34448
rect 2444 34444 5613 34448
rect 5669 34444 5696 34461
rect 2444 34396 2824 34444
rect 2270 34392 2824 34396
rect 2876 34392 2890 34444
rect 2942 34392 3378 34444
rect 3430 34392 3444 34444
rect 3496 34392 3932 34444
rect 3984 34392 3998 34444
rect 4050 34392 4486 34444
rect 4538 34392 4552 34444
rect 4604 34392 5040 34444
rect 5092 34392 5106 34444
rect 5158 34392 5594 34444
rect 5752 34428 5779 34484
rect 5835 34428 5861 34484
rect 5917 34428 5943 34484
rect 5999 34428 6025 34484
rect 6081 34428 6107 34484
rect 6266 34461 6271 34484
rect 6163 34444 6189 34461
rect 6245 34444 6271 34461
rect 6266 34428 6271 34444
rect 6327 34428 6353 34484
rect 6409 34428 6435 34484
rect 6491 34428 6517 34484
rect 6573 34428 6599 34484
rect 6655 34428 6681 34484
rect 6754 34461 6763 34484
rect 6820 34461 6845 34484
rect 6737 34444 6763 34461
rect 6819 34444 6845 34461
rect 6754 34428 6763 34444
rect 6820 34428 6845 34444
rect 6901 34428 6927 34484
rect 6983 34428 7009 34484
rect 7065 34428 7091 34484
rect 7147 34428 7173 34484
rect 7229 34428 7255 34484
rect 7311 34461 7322 34484
rect 7311 34444 7337 34461
rect 7311 34428 7322 34444
rect 7393 34428 7419 34484
rect 7475 34428 7501 34484
rect 7557 34428 7583 34484
rect 7639 34428 7665 34484
rect 7721 34428 7747 34484
rect 7803 34461 7810 34484
rect 7803 34444 7829 34461
rect 7885 34444 7911 34461
rect 7803 34428 7810 34444
rect 7967 34428 7993 34484
rect 8049 34448 8075 34465
rect 8131 34428 8157 34484
rect 8221 34465 8222 34517
rect 8213 34448 8222 34465
rect 5646 34404 5660 34428
rect 5712 34404 6148 34428
rect 6200 34404 6214 34428
rect 6266 34404 6702 34428
rect 6754 34404 6768 34428
rect 6820 34404 7256 34428
rect 7308 34404 7322 34428
rect 7374 34404 7810 34428
rect 7862 34404 7876 34428
rect 7928 34404 8047 34428
rect 8099 34404 8169 34428
rect 2270 34378 5613 34392
rect 2322 34326 2392 34378
rect 2444 34375 5613 34378
rect 5669 34375 5696 34392
rect 2444 34326 2824 34375
rect 2270 34323 2824 34326
rect 2876 34323 2890 34375
rect 2942 34323 3378 34375
rect 3430 34323 3444 34375
rect 3496 34323 3932 34375
rect 3984 34323 3998 34375
rect 4050 34323 4486 34375
rect 4538 34323 4552 34375
rect 4604 34323 5040 34375
rect 5092 34323 5106 34375
rect 5158 34323 5594 34375
rect 5752 34348 5779 34404
rect 5835 34348 5861 34404
rect 5917 34348 5943 34404
rect 5999 34348 6025 34404
rect 6081 34348 6107 34404
rect 6266 34392 6271 34404
rect 6163 34375 6189 34392
rect 6245 34375 6271 34392
rect 6266 34348 6271 34375
rect 6327 34348 6353 34404
rect 6409 34348 6435 34404
rect 6491 34348 6517 34404
rect 6573 34348 6599 34404
rect 6655 34348 6681 34404
rect 6754 34392 6763 34404
rect 6820 34392 6845 34404
rect 6737 34375 6763 34392
rect 6819 34375 6845 34392
rect 6754 34348 6763 34375
rect 6820 34348 6845 34375
rect 6901 34348 6927 34404
rect 6983 34348 7009 34404
rect 7065 34348 7091 34404
rect 7147 34348 7173 34404
rect 7229 34348 7255 34404
rect 7311 34392 7322 34404
rect 7311 34375 7337 34392
rect 7311 34348 7322 34375
rect 7393 34348 7419 34404
rect 7475 34348 7501 34404
rect 7557 34348 7583 34404
rect 7639 34348 7665 34404
rect 7721 34348 7747 34404
rect 7803 34392 7810 34404
rect 7803 34375 7829 34392
rect 7885 34375 7911 34392
rect 7803 34348 7810 34375
rect 7967 34348 7993 34404
rect 8049 34378 8075 34396
rect 8131 34348 8157 34404
rect 8221 34396 8222 34448
rect 8213 34378 8222 34396
rect 5646 34324 5660 34348
rect 5712 34324 6148 34348
rect 6200 34324 6214 34348
rect 6266 34324 6702 34348
rect 6754 34324 6768 34348
rect 6820 34324 7256 34348
rect 7308 34324 7322 34348
rect 7374 34324 7810 34348
rect 7862 34324 7876 34348
rect 7928 34326 8047 34348
rect 8099 34326 8169 34348
rect 8221 34326 8222 34378
rect 7928 34324 8222 34326
rect 2270 34308 5613 34323
rect 2322 34256 2392 34308
rect 2444 34306 5613 34308
rect 5669 34306 5696 34323
rect 2444 34256 2824 34306
rect 2270 34254 2824 34256
rect 2876 34254 2890 34306
rect 2942 34254 3378 34306
rect 3430 34254 3444 34306
rect 3496 34254 3932 34306
rect 3984 34254 3998 34306
rect 4050 34254 4486 34306
rect 4538 34254 4552 34306
rect 4604 34254 5040 34306
rect 5092 34254 5106 34306
rect 5158 34254 5594 34306
rect 5752 34268 5779 34324
rect 5835 34268 5861 34324
rect 5917 34268 5943 34324
rect 5999 34268 6025 34324
rect 6081 34268 6107 34324
rect 6266 34323 6271 34324
rect 6163 34306 6189 34323
rect 6245 34306 6271 34323
rect 6266 34268 6271 34306
rect 6327 34268 6353 34324
rect 6409 34268 6435 34324
rect 6491 34268 6517 34324
rect 6573 34268 6599 34324
rect 6655 34268 6681 34324
rect 6754 34323 6763 34324
rect 6820 34323 6845 34324
rect 6737 34306 6763 34323
rect 6819 34306 6845 34323
rect 6754 34268 6763 34306
rect 6820 34268 6845 34306
rect 6901 34268 6927 34324
rect 6983 34268 7009 34324
rect 7065 34268 7091 34324
rect 7147 34268 7173 34324
rect 7229 34268 7255 34324
rect 7311 34323 7322 34324
rect 7311 34306 7337 34323
rect 7311 34268 7322 34306
rect 7393 34268 7419 34324
rect 7475 34268 7501 34324
rect 7557 34268 7583 34324
rect 7639 34268 7665 34324
rect 7721 34268 7747 34324
rect 7803 34323 7810 34324
rect 7803 34306 7829 34323
rect 7885 34306 7911 34323
rect 7803 34268 7810 34306
rect 7967 34268 7993 34324
rect 8049 34308 8075 34324
rect 8131 34268 8157 34324
rect 8213 34308 8222 34324
rect 5646 34254 5660 34268
rect 5712 34254 6148 34268
rect 6200 34254 6214 34268
rect 6266 34254 6702 34268
rect 6754 34254 6768 34268
rect 6820 34254 7256 34268
rect 7308 34254 7322 34268
rect 7374 34254 7810 34268
rect 7862 34254 7876 34268
rect 7928 34256 8047 34268
rect 8099 34256 8169 34268
rect 8221 34256 8222 34308
rect 7928 34254 8222 34256
rect 2270 34244 8222 34254
rect 2270 34238 5613 34244
rect 2322 34186 2392 34238
rect 2444 34236 5613 34238
rect 5669 34236 5696 34244
rect 2444 34186 2824 34236
rect 2270 34184 2824 34186
rect 2876 34184 2890 34236
rect 2942 34184 3378 34236
rect 3430 34184 3444 34236
rect 3496 34184 3932 34236
rect 3984 34184 3998 34236
rect 4050 34184 4486 34236
rect 4538 34184 4552 34236
rect 4604 34184 5040 34236
rect 5092 34184 5106 34236
rect 5158 34184 5594 34236
rect 5752 34188 5779 34244
rect 5835 34188 5861 34244
rect 5917 34188 5943 34244
rect 5999 34188 6025 34244
rect 6081 34188 6107 34244
rect 6163 34236 6189 34244
rect 6245 34236 6271 34244
rect 6266 34188 6271 34236
rect 6327 34188 6353 34244
rect 6409 34188 6435 34244
rect 6491 34188 6517 34244
rect 6573 34188 6599 34244
rect 6655 34188 6681 34244
rect 6737 34236 6763 34244
rect 6819 34236 6845 34244
rect 6754 34188 6763 34236
rect 6820 34188 6845 34236
rect 6901 34188 6927 34244
rect 6983 34188 7009 34244
rect 7065 34188 7091 34244
rect 7147 34188 7173 34244
rect 7229 34188 7255 34244
rect 7311 34236 7337 34244
rect 7311 34188 7322 34236
rect 7393 34188 7419 34244
rect 7475 34188 7501 34244
rect 7557 34188 7583 34244
rect 7639 34188 7665 34244
rect 7721 34188 7747 34244
rect 7803 34236 7829 34244
rect 7885 34236 7911 34244
rect 7803 34188 7810 34236
rect 7967 34188 7993 34244
rect 8049 34238 8075 34244
rect 8131 34188 8157 34244
rect 8213 34238 8222 34244
rect 5646 34184 5660 34188
rect 5712 34184 6148 34188
rect 6200 34184 6214 34188
rect 6266 34184 6702 34188
rect 6754 34184 6768 34188
rect 6820 34184 7256 34188
rect 7308 34184 7322 34188
rect 7374 34184 7810 34188
rect 7862 34184 7876 34188
rect 7928 34186 8047 34188
rect 8099 34186 8169 34188
rect 8221 34186 8222 34238
rect 7928 34184 8222 34186
rect 2270 34168 8222 34184
rect 2322 34116 2392 34168
rect 2444 34166 8047 34168
rect 2444 34116 2824 34166
rect 2270 34114 2824 34116
rect 2876 34114 2890 34166
rect 2942 34114 3378 34166
rect 3430 34114 3444 34166
rect 3496 34114 3932 34166
rect 3984 34114 3998 34166
rect 4050 34114 4486 34166
rect 4538 34114 4552 34166
rect 4604 34114 5040 34166
rect 5092 34114 5106 34166
rect 5158 34114 5594 34166
rect 5646 34164 5660 34166
rect 5712 34164 6148 34166
rect 6200 34164 6214 34166
rect 6266 34164 6702 34166
rect 6754 34164 6768 34166
rect 6820 34164 7256 34166
rect 7308 34164 7322 34166
rect 7374 34164 7810 34166
rect 7862 34164 7876 34166
rect 7928 34164 8047 34166
rect 8099 34164 8169 34168
rect 2270 34108 5613 34114
rect 5669 34108 5696 34114
rect 5752 34108 5779 34164
rect 5835 34108 5861 34164
rect 5917 34108 5943 34164
rect 5999 34108 6025 34164
rect 6081 34108 6107 34164
rect 6266 34114 6271 34164
rect 6163 34108 6189 34114
rect 6245 34108 6271 34114
rect 6327 34108 6353 34164
rect 6409 34108 6435 34164
rect 6491 34108 6517 34164
rect 6573 34108 6599 34164
rect 6655 34108 6681 34164
rect 6754 34114 6763 34164
rect 6820 34114 6845 34164
rect 6737 34108 6763 34114
rect 6819 34108 6845 34114
rect 6901 34108 6927 34164
rect 6983 34108 7009 34164
rect 7065 34108 7091 34164
rect 7147 34108 7173 34164
rect 7229 34108 7255 34164
rect 7311 34114 7322 34164
rect 7311 34108 7337 34114
rect 7393 34108 7419 34164
rect 7475 34108 7501 34164
rect 7557 34108 7583 34164
rect 7639 34108 7665 34164
rect 7721 34108 7747 34164
rect 7803 34114 7810 34164
rect 7803 34108 7829 34114
rect 7885 34108 7911 34114
rect 7967 34108 7993 34164
rect 8049 34108 8075 34116
rect 8131 34108 8157 34164
rect 8221 34116 8222 34168
rect 8213 34108 8222 34116
rect 2724 33987 7651 33988
rect 2724 33931 2733 33987
rect 2789 33931 2814 33987
rect 2870 33931 2895 33987
rect 2951 33931 2976 33987
rect 3032 33931 3057 33987
rect 3113 33982 3138 33987
rect 3194 33982 3219 33987
rect 3275 33931 3300 33987
rect 3356 33931 3381 33987
rect 3437 33931 3462 33987
rect 3518 33931 3543 33987
rect 3599 33931 3624 33987
rect 3680 33982 3705 33987
rect 3761 33982 3786 33987
rect 3773 33931 3786 33982
rect 3842 33931 3867 33987
rect 3923 33931 3948 33987
rect 4004 33931 4029 33987
rect 4085 33931 4110 33987
rect 4166 33931 4191 33987
rect 4247 33982 4272 33987
rect 4261 33931 4272 33982
rect 4328 33931 4353 33987
rect 4409 33931 4434 33987
rect 4490 33931 4515 33987
rect 4571 33931 4596 33987
rect 4652 33931 4677 33987
rect 4733 33931 4758 33987
rect 4814 33982 4839 33987
rect 2724 33930 3101 33931
rect 3153 33930 3167 33931
rect 3219 33930 3655 33931
rect 3707 33930 3721 33931
rect 3773 33930 4209 33931
rect 4261 33930 4275 33931
rect 4327 33930 4763 33931
rect 4815 33930 4829 33982
rect 4895 33931 4920 33987
rect 4976 33931 5001 33987
rect 5057 33931 5082 33987
rect 5138 33931 5163 33987
rect 4881 33930 5163 33931
rect 2724 33913 5163 33930
rect 2724 33907 3101 33913
rect 3153 33907 3167 33913
rect 3219 33907 3655 33913
rect 3707 33907 3721 33913
rect 3773 33907 4209 33913
rect 4261 33907 4275 33913
rect 4327 33907 4763 33913
rect 2724 33851 2733 33907
rect 2789 33851 2814 33907
rect 2870 33851 2895 33907
rect 2951 33851 2976 33907
rect 3032 33851 3057 33907
rect 3113 33851 3138 33861
rect 3194 33851 3219 33861
rect 3275 33851 3300 33907
rect 3356 33851 3381 33907
rect 3437 33851 3462 33907
rect 3518 33851 3543 33907
rect 3599 33851 3624 33907
rect 3773 33861 3786 33907
rect 3680 33851 3705 33861
rect 3761 33851 3786 33861
rect 3842 33851 3867 33907
rect 3923 33851 3948 33907
rect 4004 33851 4029 33907
rect 4085 33851 4110 33907
rect 4166 33851 4191 33907
rect 4261 33861 4272 33907
rect 4247 33851 4272 33861
rect 4328 33851 4353 33907
rect 4409 33851 4434 33907
rect 4490 33851 4515 33907
rect 4571 33851 4596 33907
rect 4652 33851 4677 33907
rect 4733 33851 4758 33907
rect 4815 33861 4829 33913
rect 4881 33907 5163 33913
rect 4814 33851 4839 33861
rect 4895 33851 4920 33907
rect 4976 33851 5001 33907
rect 5057 33851 5082 33907
rect 5138 33851 5163 33907
rect 2724 33844 5163 33851
rect 2724 33827 3101 33844
rect 3153 33827 3167 33844
rect 3219 33827 3655 33844
rect 3707 33827 3721 33844
rect 3773 33827 4209 33844
rect 4261 33827 4275 33844
rect 4327 33827 4763 33844
rect 2724 33771 2733 33827
rect 2789 33771 2814 33827
rect 2870 33771 2895 33827
rect 2951 33771 2976 33827
rect 3032 33771 3057 33827
rect 3113 33775 3138 33792
rect 3194 33775 3219 33792
rect 3275 33771 3300 33827
rect 3356 33771 3381 33827
rect 3437 33771 3462 33827
rect 3518 33771 3543 33827
rect 3599 33771 3624 33827
rect 3773 33792 3786 33827
rect 3680 33775 3705 33792
rect 3761 33775 3786 33792
rect 3773 33771 3786 33775
rect 3842 33771 3867 33827
rect 3923 33771 3948 33827
rect 4004 33771 4029 33827
rect 4085 33771 4110 33827
rect 4166 33771 4191 33827
rect 4261 33792 4272 33827
rect 4247 33775 4272 33792
rect 4261 33771 4272 33775
rect 4328 33771 4353 33827
rect 4409 33771 4434 33827
rect 4490 33771 4515 33827
rect 4571 33771 4596 33827
rect 4652 33771 4677 33827
rect 4733 33771 4758 33827
rect 4815 33792 4829 33844
rect 4881 33827 5163 33844
rect 4814 33775 4839 33792
rect 2724 33747 3101 33771
rect 3153 33747 3167 33771
rect 3219 33747 3655 33771
rect 3707 33747 3721 33771
rect 3773 33747 4209 33771
rect 4261 33747 4275 33771
rect 4327 33747 4763 33771
rect 2724 33691 2733 33747
rect 2789 33691 2814 33747
rect 2870 33691 2895 33747
rect 2951 33691 2976 33747
rect 3032 33691 3057 33747
rect 3113 33706 3138 33723
rect 3194 33706 3219 33723
rect 3275 33691 3300 33747
rect 3356 33691 3381 33747
rect 3437 33691 3462 33747
rect 3518 33691 3543 33747
rect 3599 33691 3624 33747
rect 3773 33723 3786 33747
rect 3680 33706 3705 33723
rect 3761 33706 3786 33723
rect 3773 33691 3786 33706
rect 3842 33691 3867 33747
rect 3923 33691 3948 33747
rect 4004 33691 4029 33747
rect 4085 33691 4110 33747
rect 4166 33691 4191 33747
rect 4261 33723 4272 33747
rect 4247 33706 4272 33723
rect 4261 33691 4272 33706
rect 4328 33691 4353 33747
rect 4409 33691 4434 33747
rect 4490 33691 4515 33747
rect 4571 33691 4596 33747
rect 4652 33691 4677 33747
rect 4733 33691 4758 33747
rect 4815 33723 4829 33775
rect 4895 33771 4920 33827
rect 4976 33771 5001 33827
rect 5057 33771 5082 33827
rect 5138 33771 5163 33827
rect 4881 33747 5163 33771
rect 4814 33706 4839 33723
rect 2724 33667 3101 33691
rect 3153 33667 3167 33691
rect 3219 33667 3655 33691
rect 3707 33667 3721 33691
rect 3773 33667 4209 33691
rect 4261 33667 4275 33691
rect 4327 33667 4763 33691
rect 2724 33611 2733 33667
rect 2789 33611 2814 33667
rect 2870 33611 2895 33667
rect 2951 33611 2976 33667
rect 3032 33611 3057 33667
rect 3113 33636 3138 33654
rect 3194 33636 3219 33654
rect 3275 33611 3300 33667
rect 3356 33611 3381 33667
rect 3437 33611 3462 33667
rect 3518 33611 3543 33667
rect 3599 33611 3624 33667
rect 3773 33654 3786 33667
rect 3680 33636 3705 33654
rect 3761 33636 3786 33654
rect 3773 33611 3786 33636
rect 3842 33611 3867 33667
rect 3923 33611 3948 33667
rect 4004 33611 4029 33667
rect 4085 33611 4110 33667
rect 4166 33611 4191 33667
rect 4261 33654 4272 33667
rect 4247 33636 4272 33654
rect 4261 33611 4272 33636
rect 4328 33611 4353 33667
rect 4409 33611 4434 33667
rect 4490 33611 4515 33667
rect 4571 33611 4596 33667
rect 4652 33611 4677 33667
rect 4733 33611 4758 33667
rect 4815 33654 4829 33706
rect 4895 33691 4920 33747
rect 4976 33691 5001 33747
rect 5057 33691 5082 33747
rect 5138 33691 5163 33747
rect 4881 33667 5163 33691
rect 4814 33636 4839 33654
rect 2724 33587 3101 33611
rect 3153 33587 3167 33611
rect 3219 33587 3655 33611
rect 3707 33587 3721 33611
rect 3773 33587 4209 33611
rect 4261 33587 4275 33611
rect 4327 33587 4763 33611
rect 2724 33531 2733 33587
rect 2789 33531 2814 33587
rect 2870 33531 2895 33587
rect 2951 33531 2976 33587
rect 3032 33531 3057 33587
rect 3113 33566 3138 33584
rect 3194 33566 3219 33584
rect 3275 33531 3300 33587
rect 3356 33531 3381 33587
rect 3437 33531 3462 33587
rect 3518 33531 3543 33587
rect 3599 33531 3624 33587
rect 3773 33584 3786 33587
rect 3680 33566 3705 33584
rect 3761 33566 3786 33584
rect 3773 33531 3786 33566
rect 3842 33531 3867 33587
rect 3923 33531 3948 33587
rect 4004 33531 4029 33587
rect 4085 33531 4110 33587
rect 4166 33531 4191 33587
rect 4261 33584 4272 33587
rect 4247 33566 4272 33584
rect 4261 33531 4272 33566
rect 4328 33531 4353 33587
rect 4409 33531 4434 33587
rect 4490 33531 4515 33587
rect 4571 33531 4596 33587
rect 4652 33531 4677 33587
rect 4733 33531 4758 33587
rect 4815 33584 4829 33636
rect 4895 33611 4920 33667
rect 4976 33611 5001 33667
rect 5057 33611 5082 33667
rect 5138 33611 5163 33667
rect 4881 33587 5163 33611
rect 4814 33566 4839 33584
rect 2724 33514 3101 33531
rect 3153 33514 3167 33531
rect 3219 33514 3655 33531
rect 3707 33514 3721 33531
rect 3773 33514 4209 33531
rect 4261 33514 4275 33531
rect 4327 33514 4763 33531
rect 4815 33514 4829 33566
rect 4895 33531 4920 33587
rect 4976 33531 5001 33587
rect 5057 33531 5082 33587
rect 5138 33531 5163 33587
rect 4881 33514 5163 33531
rect 2724 33507 5163 33514
rect 2724 33451 2733 33507
rect 2789 33451 2814 33507
rect 2870 33451 2895 33507
rect 2951 33451 2976 33507
rect 3032 33451 3057 33507
rect 3113 33496 3138 33507
rect 3194 33496 3219 33507
rect 3275 33451 3300 33507
rect 3356 33451 3381 33507
rect 3437 33451 3462 33507
rect 3518 33451 3543 33507
rect 3599 33451 3624 33507
rect 3680 33496 3705 33507
rect 3761 33496 3786 33507
rect 3773 33451 3786 33496
rect 3842 33451 3867 33507
rect 3923 33451 3948 33507
rect 4004 33451 4029 33507
rect 4085 33451 4110 33507
rect 4166 33451 4191 33507
rect 4247 33496 4272 33507
rect 4261 33451 4272 33496
rect 4328 33451 4353 33507
rect 4409 33451 4434 33507
rect 4490 33451 4515 33507
rect 4571 33451 4596 33507
rect 4652 33451 4677 33507
rect 4733 33451 4758 33507
rect 4814 33496 4839 33507
rect 2724 33444 3101 33451
rect 3153 33444 3167 33451
rect 3219 33444 3655 33451
rect 3707 33444 3721 33451
rect 3773 33444 4209 33451
rect 4261 33444 4275 33451
rect 4327 33444 4763 33451
rect 4815 33444 4829 33496
rect 4895 33451 4920 33507
rect 4976 33451 5001 33507
rect 5057 33451 5082 33507
rect 5138 33451 5163 33507
rect 4881 33444 5163 33451
rect 2724 33427 5163 33444
rect 2724 33371 2733 33427
rect 2789 33371 2814 33427
rect 2870 33371 2895 33427
rect 2951 33371 2976 33427
rect 3032 33371 3057 33427
rect 3113 33426 3138 33427
rect 3194 33426 3219 33427
rect 3113 33371 3138 33374
rect 3194 33371 3219 33374
rect 3275 33371 3300 33427
rect 3356 33371 3381 33427
rect 3437 33371 3462 33427
rect 3518 33371 3543 33427
rect 3599 33371 3624 33427
rect 3680 33426 3705 33427
rect 3761 33426 3786 33427
rect 3773 33374 3786 33426
rect 3680 33371 3705 33374
rect 3761 33371 3786 33374
rect 3842 33371 3867 33427
rect 3923 33371 3948 33427
rect 4004 33371 4029 33427
rect 4085 33371 4110 33427
rect 4166 33371 4191 33427
rect 4247 33426 4272 33427
rect 4261 33374 4272 33426
rect 4247 33371 4272 33374
rect 4328 33371 4353 33427
rect 4409 33371 4434 33427
rect 4490 33371 4515 33427
rect 4571 33371 4596 33427
rect 4652 33371 4677 33427
rect 4733 33371 4758 33427
rect 4814 33426 4839 33427
rect 4815 33374 4829 33426
rect 4814 33371 4839 33374
rect 4895 33371 4920 33427
rect 4976 33371 5001 33427
rect 5057 33371 5082 33427
rect 5138 33371 5163 33427
rect 5299 33982 7651 33987
rect 5299 33930 5317 33982
rect 5369 33930 5383 33982
rect 5435 33930 5871 33982
rect 5923 33930 5937 33982
rect 5989 33930 6425 33982
rect 6477 33930 6491 33982
rect 6543 33930 6979 33982
rect 7031 33930 7045 33982
rect 7097 33930 7533 33982
rect 7585 33930 7599 33982
rect 5299 33913 7651 33930
rect 5299 33861 5317 33913
rect 5369 33861 5383 33913
rect 5435 33861 5871 33913
rect 5923 33861 5937 33913
rect 5989 33861 6425 33913
rect 6477 33861 6491 33913
rect 6543 33861 6979 33913
rect 7031 33861 7045 33913
rect 7097 33861 7533 33913
rect 7585 33861 7599 33913
rect 5299 33844 7651 33861
rect 5299 33792 5317 33844
rect 5369 33792 5383 33844
rect 5435 33792 5871 33844
rect 5923 33792 5937 33844
rect 5989 33792 6425 33844
rect 6477 33792 6491 33844
rect 6543 33792 6979 33844
rect 7031 33792 7045 33844
rect 7097 33792 7533 33844
rect 7585 33792 7599 33844
rect 5299 33775 7651 33792
rect 5299 33723 5317 33775
rect 5369 33723 5383 33775
rect 5435 33723 5871 33775
rect 5923 33723 5937 33775
rect 5989 33723 6425 33775
rect 6477 33723 6491 33775
rect 6543 33723 6979 33775
rect 7031 33723 7045 33775
rect 7097 33723 7533 33775
rect 7585 33723 7599 33775
rect 5299 33706 7651 33723
rect 5299 33654 5317 33706
rect 5369 33654 5383 33706
rect 5435 33654 5871 33706
rect 5923 33654 5937 33706
rect 5989 33654 6425 33706
rect 6477 33654 6491 33706
rect 6543 33654 6979 33706
rect 7031 33654 7045 33706
rect 7097 33654 7533 33706
rect 7585 33654 7599 33706
rect 5299 33636 7651 33654
rect 5299 33584 5317 33636
rect 5369 33584 5383 33636
rect 5435 33584 5871 33636
rect 5923 33584 5937 33636
rect 5989 33584 6425 33636
rect 6477 33584 6491 33636
rect 6543 33584 6979 33636
rect 7031 33584 7045 33636
rect 7097 33584 7533 33636
rect 7585 33584 7599 33636
rect 5299 33566 7651 33584
rect 5299 33514 5317 33566
rect 5369 33514 5383 33566
rect 5435 33514 5871 33566
rect 5923 33514 5937 33566
rect 5989 33514 6425 33566
rect 6477 33514 6491 33566
rect 6543 33514 6979 33566
rect 7031 33514 7045 33566
rect 7097 33514 7533 33566
rect 7585 33514 7599 33566
rect 5299 33496 7651 33514
rect 5299 33444 5317 33496
rect 5369 33444 5383 33496
rect 5435 33444 5871 33496
rect 5923 33444 5937 33496
rect 5989 33444 6425 33496
rect 6477 33444 6491 33496
rect 6543 33444 6979 33496
rect 7031 33444 7045 33496
rect 7097 33444 7533 33496
rect 7585 33444 7599 33496
rect 5299 33426 7651 33444
rect 5299 33374 5317 33426
rect 5369 33374 5383 33426
rect 5435 33374 5871 33426
rect 5923 33374 5937 33426
rect 5989 33374 6425 33426
rect 6477 33374 6491 33426
rect 6543 33374 6979 33426
rect 7031 33374 7045 33426
rect 7097 33374 7533 33426
rect 7585 33374 7599 33426
rect 5299 33371 7651 33374
rect 2724 33368 7651 33371
rect 2270 32724 8222 32730
rect 2322 32672 2392 32724
rect 2444 32720 5613 32724
rect 5669 32720 5696 32724
rect 2444 32672 2824 32720
rect 2270 32668 2824 32672
rect 2876 32668 2890 32720
rect 2942 32668 3378 32720
rect 3430 32668 3444 32720
rect 3496 32668 3932 32720
rect 3984 32668 3998 32720
rect 4050 32668 4486 32720
rect 4538 32668 4552 32720
rect 4604 32668 5040 32720
rect 5092 32668 5106 32720
rect 5158 32668 5594 32720
rect 5752 32668 5779 32724
rect 5835 32668 5861 32724
rect 5917 32668 5943 32724
rect 5999 32668 6025 32724
rect 6081 32668 6107 32724
rect 6163 32720 6189 32724
rect 6245 32720 6271 32724
rect 6266 32668 6271 32720
rect 6327 32668 6353 32724
rect 6409 32668 6435 32724
rect 6491 32668 6517 32724
rect 6573 32668 6599 32724
rect 6655 32668 6681 32724
rect 6737 32720 6763 32724
rect 6819 32720 6845 32724
rect 6754 32668 6763 32720
rect 6820 32668 6845 32720
rect 6901 32668 6927 32724
rect 6983 32668 7009 32724
rect 7065 32668 7091 32724
rect 7147 32668 7173 32724
rect 7229 32668 7255 32724
rect 7311 32720 7337 32724
rect 7311 32668 7322 32720
rect 7393 32668 7419 32724
rect 7475 32668 7501 32724
rect 7557 32668 7583 32724
rect 7639 32668 7665 32724
rect 7721 32668 7747 32724
rect 7803 32720 7829 32724
rect 7885 32720 7911 32724
rect 7803 32668 7810 32720
rect 7967 32668 7993 32724
rect 8049 32668 8075 32672
rect 8131 32668 8157 32724
rect 8221 32672 8222 32724
rect 8213 32668 8222 32672
rect 2270 32655 8222 32668
rect 2322 32603 2392 32655
rect 2444 32651 8047 32655
rect 2444 32603 2824 32651
rect 2270 32599 2824 32603
rect 2876 32599 2890 32651
rect 2942 32599 3378 32651
rect 3430 32599 3444 32651
rect 3496 32599 3932 32651
rect 3984 32599 3998 32651
rect 4050 32599 4486 32651
rect 4538 32599 4552 32651
rect 4604 32599 5040 32651
rect 5092 32599 5106 32651
rect 5158 32599 5594 32651
rect 5646 32644 5660 32651
rect 5712 32644 6148 32651
rect 6200 32644 6214 32651
rect 6266 32644 6702 32651
rect 6754 32644 6768 32651
rect 6820 32644 7256 32651
rect 7308 32644 7322 32651
rect 7374 32644 7810 32651
rect 7862 32644 7876 32651
rect 7928 32644 8047 32651
rect 8099 32644 8169 32655
rect 2270 32588 5613 32599
rect 5669 32588 5696 32599
rect 5752 32588 5779 32644
rect 5835 32588 5861 32644
rect 5917 32588 5943 32644
rect 5999 32588 6025 32644
rect 6081 32588 6107 32644
rect 6266 32599 6271 32644
rect 6163 32588 6189 32599
rect 6245 32588 6271 32599
rect 6327 32588 6353 32644
rect 6409 32588 6435 32644
rect 6491 32588 6517 32644
rect 6573 32588 6599 32644
rect 6655 32588 6681 32644
rect 6754 32599 6763 32644
rect 6820 32599 6845 32644
rect 6737 32588 6763 32599
rect 6819 32588 6845 32599
rect 6901 32588 6927 32644
rect 6983 32588 7009 32644
rect 7065 32588 7091 32644
rect 7147 32588 7173 32644
rect 7229 32588 7255 32644
rect 7311 32599 7322 32644
rect 7311 32588 7337 32599
rect 7393 32588 7419 32644
rect 7475 32588 7501 32644
rect 7557 32588 7583 32644
rect 7639 32588 7665 32644
rect 7721 32588 7747 32644
rect 7803 32599 7810 32644
rect 7803 32588 7829 32599
rect 7885 32588 7911 32599
rect 7967 32588 7993 32644
rect 8049 32588 8075 32603
rect 8131 32588 8157 32644
rect 8221 32603 8222 32655
rect 8213 32588 8222 32603
rect 2270 32586 8222 32588
rect 2322 32534 2392 32586
rect 2444 32582 8047 32586
rect 2444 32534 2824 32582
rect 2270 32530 2824 32534
rect 2876 32530 2890 32582
rect 2942 32530 3378 32582
rect 3430 32530 3444 32582
rect 3496 32530 3932 32582
rect 3984 32530 3998 32582
rect 4050 32530 4486 32582
rect 4538 32530 4552 32582
rect 4604 32530 5040 32582
rect 5092 32530 5106 32582
rect 5158 32530 5594 32582
rect 5646 32564 5660 32582
rect 5712 32564 6148 32582
rect 6200 32564 6214 32582
rect 6266 32564 6702 32582
rect 6754 32564 6768 32582
rect 6820 32564 7256 32582
rect 7308 32564 7322 32582
rect 7374 32564 7810 32582
rect 7862 32564 7876 32582
rect 7928 32564 8047 32582
rect 8099 32564 8169 32586
rect 2270 32517 5613 32530
rect 2322 32465 2392 32517
rect 2444 32513 5613 32517
rect 5669 32513 5696 32530
rect 2444 32465 2824 32513
rect 2270 32461 2824 32465
rect 2876 32461 2890 32513
rect 2942 32461 3378 32513
rect 3430 32461 3444 32513
rect 3496 32461 3932 32513
rect 3984 32461 3998 32513
rect 4050 32461 4486 32513
rect 4538 32461 4552 32513
rect 4604 32461 5040 32513
rect 5092 32461 5106 32513
rect 5158 32461 5594 32513
rect 5752 32508 5779 32564
rect 5835 32508 5861 32564
rect 5917 32508 5943 32564
rect 5999 32508 6025 32564
rect 6081 32508 6107 32564
rect 6266 32530 6271 32564
rect 6163 32513 6189 32530
rect 6245 32513 6271 32530
rect 6266 32508 6271 32513
rect 6327 32508 6353 32564
rect 6409 32508 6435 32564
rect 6491 32508 6517 32564
rect 6573 32508 6599 32564
rect 6655 32508 6681 32564
rect 6754 32530 6763 32564
rect 6820 32530 6845 32564
rect 6737 32513 6763 32530
rect 6819 32513 6845 32530
rect 6754 32508 6763 32513
rect 6820 32508 6845 32513
rect 6901 32508 6927 32564
rect 6983 32508 7009 32564
rect 7065 32508 7091 32564
rect 7147 32508 7173 32564
rect 7229 32508 7255 32564
rect 7311 32530 7322 32564
rect 7311 32513 7337 32530
rect 7311 32508 7322 32513
rect 7393 32508 7419 32564
rect 7475 32508 7501 32564
rect 7557 32508 7583 32564
rect 7639 32508 7665 32564
rect 7721 32508 7747 32564
rect 7803 32530 7810 32564
rect 7803 32513 7829 32530
rect 7885 32513 7911 32530
rect 7803 32508 7810 32513
rect 7967 32508 7993 32564
rect 8049 32517 8075 32534
rect 8131 32508 8157 32564
rect 8221 32534 8222 32586
rect 8213 32517 8222 32534
rect 5646 32484 5660 32508
rect 5712 32484 6148 32508
rect 6200 32484 6214 32508
rect 6266 32484 6702 32508
rect 6754 32484 6768 32508
rect 6820 32484 7256 32508
rect 7308 32484 7322 32508
rect 7374 32484 7810 32508
rect 7862 32484 7876 32508
rect 7928 32484 8047 32508
rect 8099 32484 8169 32508
rect 2270 32448 5613 32461
rect 2322 32396 2392 32448
rect 2444 32444 5613 32448
rect 5669 32444 5696 32461
rect 2444 32396 2824 32444
rect 2270 32392 2824 32396
rect 2876 32392 2890 32444
rect 2942 32392 3378 32444
rect 3430 32392 3444 32444
rect 3496 32392 3932 32444
rect 3984 32392 3998 32444
rect 4050 32392 4486 32444
rect 4538 32392 4552 32444
rect 4604 32392 5040 32444
rect 5092 32392 5106 32444
rect 5158 32392 5594 32444
rect 5752 32428 5779 32484
rect 5835 32428 5861 32484
rect 5917 32428 5943 32484
rect 5999 32428 6025 32484
rect 6081 32428 6107 32484
rect 6266 32461 6271 32484
rect 6163 32444 6189 32461
rect 6245 32444 6271 32461
rect 6266 32428 6271 32444
rect 6327 32428 6353 32484
rect 6409 32428 6435 32484
rect 6491 32428 6517 32484
rect 6573 32428 6599 32484
rect 6655 32428 6681 32484
rect 6754 32461 6763 32484
rect 6820 32461 6845 32484
rect 6737 32444 6763 32461
rect 6819 32444 6845 32461
rect 6754 32428 6763 32444
rect 6820 32428 6845 32444
rect 6901 32428 6927 32484
rect 6983 32428 7009 32484
rect 7065 32428 7091 32484
rect 7147 32428 7173 32484
rect 7229 32428 7255 32484
rect 7311 32461 7322 32484
rect 7311 32444 7337 32461
rect 7311 32428 7322 32444
rect 7393 32428 7419 32484
rect 7475 32428 7501 32484
rect 7557 32428 7583 32484
rect 7639 32428 7665 32484
rect 7721 32428 7747 32484
rect 7803 32461 7810 32484
rect 7803 32444 7829 32461
rect 7885 32444 7911 32461
rect 7803 32428 7810 32444
rect 7967 32428 7993 32484
rect 8049 32448 8075 32465
rect 8131 32428 8157 32484
rect 8221 32465 8222 32517
rect 8213 32448 8222 32465
rect 5646 32404 5660 32428
rect 5712 32404 6148 32428
rect 6200 32404 6214 32428
rect 6266 32404 6702 32428
rect 6754 32404 6768 32428
rect 6820 32404 7256 32428
rect 7308 32404 7322 32428
rect 7374 32404 7810 32428
rect 7862 32404 7876 32428
rect 7928 32404 8047 32428
rect 8099 32404 8169 32428
rect 2270 32378 5613 32392
rect 2322 32326 2392 32378
rect 2444 32375 5613 32378
rect 5669 32375 5696 32392
rect 2444 32326 2824 32375
rect 2270 32323 2824 32326
rect 2876 32323 2890 32375
rect 2942 32323 3378 32375
rect 3430 32323 3444 32375
rect 3496 32323 3932 32375
rect 3984 32323 3998 32375
rect 4050 32323 4486 32375
rect 4538 32323 4552 32375
rect 4604 32323 5040 32375
rect 5092 32323 5106 32375
rect 5158 32323 5594 32375
rect 5752 32348 5779 32404
rect 5835 32348 5861 32404
rect 5917 32348 5943 32404
rect 5999 32348 6025 32404
rect 6081 32348 6107 32404
rect 6266 32392 6271 32404
rect 6163 32375 6189 32392
rect 6245 32375 6271 32392
rect 6266 32348 6271 32375
rect 6327 32348 6353 32404
rect 6409 32348 6435 32404
rect 6491 32348 6517 32404
rect 6573 32348 6599 32404
rect 6655 32348 6681 32404
rect 6754 32392 6763 32404
rect 6820 32392 6845 32404
rect 6737 32375 6763 32392
rect 6819 32375 6845 32392
rect 6754 32348 6763 32375
rect 6820 32348 6845 32375
rect 6901 32348 6927 32404
rect 6983 32348 7009 32404
rect 7065 32348 7091 32404
rect 7147 32348 7173 32404
rect 7229 32348 7255 32404
rect 7311 32392 7322 32404
rect 7311 32375 7337 32392
rect 7311 32348 7322 32375
rect 7393 32348 7419 32404
rect 7475 32348 7501 32404
rect 7557 32348 7583 32404
rect 7639 32348 7665 32404
rect 7721 32348 7747 32404
rect 7803 32392 7810 32404
rect 7803 32375 7829 32392
rect 7885 32375 7911 32392
rect 7803 32348 7810 32375
rect 7967 32348 7993 32404
rect 8049 32378 8075 32396
rect 8131 32348 8157 32404
rect 8221 32396 8222 32448
rect 8213 32378 8222 32396
rect 5646 32324 5660 32348
rect 5712 32324 6148 32348
rect 6200 32324 6214 32348
rect 6266 32324 6702 32348
rect 6754 32324 6768 32348
rect 6820 32324 7256 32348
rect 7308 32324 7322 32348
rect 7374 32324 7810 32348
rect 7862 32324 7876 32348
rect 7928 32326 8047 32348
rect 8099 32326 8169 32348
rect 8221 32326 8222 32378
rect 7928 32324 8222 32326
rect 2270 32308 5613 32323
rect 2322 32256 2392 32308
rect 2444 32306 5613 32308
rect 5669 32306 5696 32323
rect 2444 32256 2824 32306
rect 2270 32254 2824 32256
rect 2876 32254 2890 32306
rect 2942 32254 3378 32306
rect 3430 32254 3444 32306
rect 3496 32254 3932 32306
rect 3984 32254 3998 32306
rect 4050 32254 4486 32306
rect 4538 32254 4552 32306
rect 4604 32254 5040 32306
rect 5092 32254 5106 32306
rect 5158 32254 5594 32306
rect 5752 32268 5779 32324
rect 5835 32268 5861 32324
rect 5917 32268 5943 32324
rect 5999 32268 6025 32324
rect 6081 32268 6107 32324
rect 6266 32323 6271 32324
rect 6163 32306 6189 32323
rect 6245 32306 6271 32323
rect 6266 32268 6271 32306
rect 6327 32268 6353 32324
rect 6409 32268 6435 32324
rect 6491 32268 6517 32324
rect 6573 32268 6599 32324
rect 6655 32268 6681 32324
rect 6754 32323 6763 32324
rect 6820 32323 6845 32324
rect 6737 32306 6763 32323
rect 6819 32306 6845 32323
rect 6754 32268 6763 32306
rect 6820 32268 6845 32306
rect 6901 32268 6927 32324
rect 6983 32268 7009 32324
rect 7065 32268 7091 32324
rect 7147 32268 7173 32324
rect 7229 32268 7255 32324
rect 7311 32323 7322 32324
rect 7311 32306 7337 32323
rect 7311 32268 7322 32306
rect 7393 32268 7419 32324
rect 7475 32268 7501 32324
rect 7557 32268 7583 32324
rect 7639 32268 7665 32324
rect 7721 32268 7747 32324
rect 7803 32323 7810 32324
rect 7803 32306 7829 32323
rect 7885 32306 7911 32323
rect 7803 32268 7810 32306
rect 7967 32268 7993 32324
rect 8049 32308 8075 32324
rect 8131 32268 8157 32324
rect 8213 32308 8222 32324
rect 5646 32254 5660 32268
rect 5712 32254 6148 32268
rect 6200 32254 6214 32268
rect 6266 32254 6702 32268
rect 6754 32254 6768 32268
rect 6820 32254 7256 32268
rect 7308 32254 7322 32268
rect 7374 32254 7810 32268
rect 7862 32254 7876 32268
rect 7928 32256 8047 32268
rect 8099 32256 8169 32268
rect 8221 32256 8222 32308
rect 7928 32254 8222 32256
rect 2270 32244 8222 32254
rect 2270 32238 5613 32244
rect 2322 32186 2392 32238
rect 2444 32236 5613 32238
rect 5669 32236 5696 32244
rect 2444 32186 2824 32236
rect 2270 32184 2824 32186
rect 2876 32184 2890 32236
rect 2942 32184 3378 32236
rect 3430 32184 3444 32236
rect 3496 32184 3932 32236
rect 3984 32184 3998 32236
rect 4050 32184 4486 32236
rect 4538 32184 4552 32236
rect 4604 32184 5040 32236
rect 5092 32184 5106 32236
rect 5158 32184 5594 32236
rect 5752 32188 5779 32244
rect 5835 32188 5861 32244
rect 5917 32188 5943 32244
rect 5999 32188 6025 32244
rect 6081 32188 6107 32244
rect 6163 32236 6189 32244
rect 6245 32236 6271 32244
rect 6266 32188 6271 32236
rect 6327 32188 6353 32244
rect 6409 32188 6435 32244
rect 6491 32188 6517 32244
rect 6573 32188 6599 32244
rect 6655 32188 6681 32244
rect 6737 32236 6763 32244
rect 6819 32236 6845 32244
rect 6754 32188 6763 32236
rect 6820 32188 6845 32236
rect 6901 32188 6927 32244
rect 6983 32188 7009 32244
rect 7065 32188 7091 32244
rect 7147 32188 7173 32244
rect 7229 32188 7255 32244
rect 7311 32236 7337 32244
rect 7311 32188 7322 32236
rect 7393 32188 7419 32244
rect 7475 32188 7501 32244
rect 7557 32188 7583 32244
rect 7639 32188 7665 32244
rect 7721 32188 7747 32244
rect 7803 32236 7829 32244
rect 7885 32236 7911 32244
rect 7803 32188 7810 32236
rect 7967 32188 7993 32244
rect 8049 32238 8075 32244
rect 8131 32188 8157 32244
rect 8213 32238 8222 32244
rect 5646 32184 5660 32188
rect 5712 32184 6148 32188
rect 6200 32184 6214 32188
rect 6266 32184 6702 32188
rect 6754 32184 6768 32188
rect 6820 32184 7256 32188
rect 7308 32184 7322 32188
rect 7374 32184 7810 32188
rect 7862 32184 7876 32188
rect 7928 32186 8047 32188
rect 8099 32186 8169 32188
rect 8221 32186 8222 32238
rect 7928 32184 8222 32186
rect 2270 32168 8222 32184
rect 2322 32116 2392 32168
rect 2444 32166 8047 32168
rect 2444 32116 2824 32166
rect 2270 32114 2824 32116
rect 2876 32114 2890 32166
rect 2942 32114 3378 32166
rect 3430 32114 3444 32166
rect 3496 32114 3932 32166
rect 3984 32114 3998 32166
rect 4050 32114 4486 32166
rect 4538 32114 4552 32166
rect 4604 32114 5040 32166
rect 5092 32114 5106 32166
rect 5158 32114 5594 32166
rect 5646 32164 5660 32166
rect 5712 32164 6148 32166
rect 6200 32164 6214 32166
rect 6266 32164 6702 32166
rect 6754 32164 6768 32166
rect 6820 32164 7256 32166
rect 7308 32164 7322 32166
rect 7374 32164 7810 32166
rect 7862 32164 7876 32166
rect 7928 32164 8047 32166
rect 8099 32164 8169 32168
rect 2270 32108 5613 32114
rect 5669 32108 5696 32114
rect 5752 32108 5779 32164
rect 5835 32108 5861 32164
rect 5917 32108 5943 32164
rect 5999 32108 6025 32164
rect 6081 32108 6107 32164
rect 6266 32114 6271 32164
rect 6163 32108 6189 32114
rect 6245 32108 6271 32114
rect 6327 32108 6353 32164
rect 6409 32108 6435 32164
rect 6491 32108 6517 32164
rect 6573 32108 6599 32164
rect 6655 32108 6681 32164
rect 6754 32114 6763 32164
rect 6820 32114 6845 32164
rect 6737 32108 6763 32114
rect 6819 32108 6845 32114
rect 6901 32108 6927 32164
rect 6983 32108 7009 32164
rect 7065 32108 7091 32164
rect 7147 32108 7173 32164
rect 7229 32108 7255 32164
rect 7311 32114 7322 32164
rect 7311 32108 7337 32114
rect 7393 32108 7419 32164
rect 7475 32108 7501 32164
rect 7557 32108 7583 32164
rect 7639 32108 7665 32164
rect 7721 32108 7747 32164
rect 7803 32114 7810 32164
rect 7803 32108 7829 32114
rect 7885 32108 7911 32114
rect 7967 32108 7993 32164
rect 8049 32108 8075 32116
rect 8131 32108 8157 32164
rect 8221 32116 8222 32168
rect 8213 32108 8222 32116
rect 2724 31987 7651 31988
rect 2724 31931 2733 31987
rect 2789 31931 2814 31987
rect 2870 31931 2895 31987
rect 2951 31931 2976 31987
rect 3032 31931 3057 31987
rect 3113 31982 3138 31987
rect 3194 31982 3219 31987
rect 3275 31931 3300 31987
rect 3356 31931 3381 31987
rect 3437 31931 3462 31987
rect 3518 31931 3543 31987
rect 3599 31931 3624 31987
rect 3680 31982 3705 31987
rect 3761 31982 3786 31987
rect 3773 31931 3786 31982
rect 3842 31931 3867 31987
rect 3923 31931 3948 31987
rect 4004 31931 4029 31987
rect 4085 31931 4110 31987
rect 4166 31931 4191 31987
rect 4247 31982 4272 31987
rect 4261 31931 4272 31982
rect 4328 31931 4353 31987
rect 4409 31931 4434 31987
rect 4490 31931 4515 31987
rect 4571 31931 4596 31987
rect 4652 31931 4677 31987
rect 4733 31931 4758 31987
rect 4814 31982 4839 31987
rect 2724 31930 3101 31931
rect 3153 31930 3167 31931
rect 3219 31930 3655 31931
rect 3707 31930 3721 31931
rect 3773 31930 4209 31931
rect 4261 31930 4275 31931
rect 4327 31930 4763 31931
rect 4815 31930 4829 31982
rect 4895 31931 4920 31987
rect 4976 31931 5001 31987
rect 5057 31931 5082 31987
rect 5138 31931 5163 31987
rect 4881 31930 5163 31931
rect 2724 31913 5163 31930
rect 2724 31907 3101 31913
rect 3153 31907 3167 31913
rect 3219 31907 3655 31913
rect 3707 31907 3721 31913
rect 3773 31907 4209 31913
rect 4261 31907 4275 31913
rect 4327 31907 4763 31913
rect 2724 31851 2733 31907
rect 2789 31851 2814 31907
rect 2870 31851 2895 31907
rect 2951 31851 2976 31907
rect 3032 31851 3057 31907
rect 3113 31851 3138 31861
rect 3194 31851 3219 31861
rect 3275 31851 3300 31907
rect 3356 31851 3381 31907
rect 3437 31851 3462 31907
rect 3518 31851 3543 31907
rect 3599 31851 3624 31907
rect 3773 31861 3786 31907
rect 3680 31851 3705 31861
rect 3761 31851 3786 31861
rect 3842 31851 3867 31907
rect 3923 31851 3948 31907
rect 4004 31851 4029 31907
rect 4085 31851 4110 31907
rect 4166 31851 4191 31907
rect 4261 31861 4272 31907
rect 4247 31851 4272 31861
rect 4328 31851 4353 31907
rect 4409 31851 4434 31907
rect 4490 31851 4515 31907
rect 4571 31851 4596 31907
rect 4652 31851 4677 31907
rect 4733 31851 4758 31907
rect 4815 31861 4829 31913
rect 4881 31907 5163 31913
rect 4814 31851 4839 31861
rect 4895 31851 4920 31907
rect 4976 31851 5001 31907
rect 5057 31851 5082 31907
rect 5138 31851 5163 31907
rect 2724 31844 5163 31851
rect 2724 31827 3101 31844
rect 3153 31827 3167 31844
rect 3219 31827 3655 31844
rect 3707 31827 3721 31844
rect 3773 31827 4209 31844
rect 4261 31827 4275 31844
rect 4327 31827 4763 31844
rect 2724 31771 2733 31827
rect 2789 31771 2814 31827
rect 2870 31771 2895 31827
rect 2951 31771 2976 31827
rect 3032 31771 3057 31827
rect 3113 31775 3138 31792
rect 3194 31775 3219 31792
rect 3275 31771 3300 31827
rect 3356 31771 3381 31827
rect 3437 31771 3462 31827
rect 3518 31771 3543 31827
rect 3599 31771 3624 31827
rect 3773 31792 3786 31827
rect 3680 31775 3705 31792
rect 3761 31775 3786 31792
rect 3773 31771 3786 31775
rect 3842 31771 3867 31827
rect 3923 31771 3948 31827
rect 4004 31771 4029 31827
rect 4085 31771 4110 31827
rect 4166 31771 4191 31827
rect 4261 31792 4272 31827
rect 4247 31775 4272 31792
rect 4261 31771 4272 31775
rect 4328 31771 4353 31827
rect 4409 31771 4434 31827
rect 4490 31771 4515 31827
rect 4571 31771 4596 31827
rect 4652 31771 4677 31827
rect 4733 31771 4758 31827
rect 4815 31792 4829 31844
rect 4881 31827 5163 31844
rect 4814 31775 4839 31792
rect 2724 31747 3101 31771
rect 3153 31747 3167 31771
rect 3219 31747 3655 31771
rect 3707 31747 3721 31771
rect 3773 31747 4209 31771
rect 4261 31747 4275 31771
rect 4327 31747 4763 31771
rect 2724 31691 2733 31747
rect 2789 31691 2814 31747
rect 2870 31691 2895 31747
rect 2951 31691 2976 31747
rect 3032 31691 3057 31747
rect 3113 31706 3138 31723
rect 3194 31706 3219 31723
rect 3275 31691 3300 31747
rect 3356 31691 3381 31747
rect 3437 31691 3462 31747
rect 3518 31691 3543 31747
rect 3599 31691 3624 31747
rect 3773 31723 3786 31747
rect 3680 31706 3705 31723
rect 3761 31706 3786 31723
rect 3773 31691 3786 31706
rect 3842 31691 3867 31747
rect 3923 31691 3948 31747
rect 4004 31691 4029 31747
rect 4085 31691 4110 31747
rect 4166 31691 4191 31747
rect 4261 31723 4272 31747
rect 4247 31706 4272 31723
rect 4261 31691 4272 31706
rect 4328 31691 4353 31747
rect 4409 31691 4434 31747
rect 4490 31691 4515 31747
rect 4571 31691 4596 31747
rect 4652 31691 4677 31747
rect 4733 31691 4758 31747
rect 4815 31723 4829 31775
rect 4895 31771 4920 31827
rect 4976 31771 5001 31827
rect 5057 31771 5082 31827
rect 5138 31771 5163 31827
rect 4881 31747 5163 31771
rect 4814 31706 4839 31723
rect 2724 31667 3101 31691
rect 3153 31667 3167 31691
rect 3219 31667 3655 31691
rect 3707 31667 3721 31691
rect 3773 31667 4209 31691
rect 4261 31667 4275 31691
rect 4327 31667 4763 31691
rect 2724 31611 2733 31667
rect 2789 31611 2814 31667
rect 2870 31611 2895 31667
rect 2951 31611 2976 31667
rect 3032 31611 3057 31667
rect 3113 31636 3138 31654
rect 3194 31636 3219 31654
rect 3275 31611 3300 31667
rect 3356 31611 3381 31667
rect 3437 31611 3462 31667
rect 3518 31611 3543 31667
rect 3599 31611 3624 31667
rect 3773 31654 3786 31667
rect 3680 31636 3705 31654
rect 3761 31636 3786 31654
rect 3773 31611 3786 31636
rect 3842 31611 3867 31667
rect 3923 31611 3948 31667
rect 4004 31611 4029 31667
rect 4085 31611 4110 31667
rect 4166 31611 4191 31667
rect 4261 31654 4272 31667
rect 4247 31636 4272 31654
rect 4261 31611 4272 31636
rect 4328 31611 4353 31667
rect 4409 31611 4434 31667
rect 4490 31611 4515 31667
rect 4571 31611 4596 31667
rect 4652 31611 4677 31667
rect 4733 31611 4758 31667
rect 4815 31654 4829 31706
rect 4895 31691 4920 31747
rect 4976 31691 5001 31747
rect 5057 31691 5082 31747
rect 5138 31691 5163 31747
rect 4881 31667 5163 31691
rect 4814 31636 4839 31654
rect 2724 31587 3101 31611
rect 3153 31587 3167 31611
rect 3219 31587 3655 31611
rect 3707 31587 3721 31611
rect 3773 31587 4209 31611
rect 4261 31587 4275 31611
rect 4327 31587 4763 31611
rect 2724 31531 2733 31587
rect 2789 31531 2814 31587
rect 2870 31531 2895 31587
rect 2951 31531 2976 31587
rect 3032 31531 3057 31587
rect 3113 31566 3138 31584
rect 3194 31566 3219 31584
rect 3275 31531 3300 31587
rect 3356 31531 3381 31587
rect 3437 31531 3462 31587
rect 3518 31531 3543 31587
rect 3599 31531 3624 31587
rect 3773 31584 3786 31587
rect 3680 31566 3705 31584
rect 3761 31566 3786 31584
rect 3773 31531 3786 31566
rect 3842 31531 3867 31587
rect 3923 31531 3948 31587
rect 4004 31531 4029 31587
rect 4085 31531 4110 31587
rect 4166 31531 4191 31587
rect 4261 31584 4272 31587
rect 4247 31566 4272 31584
rect 4261 31531 4272 31566
rect 4328 31531 4353 31587
rect 4409 31531 4434 31587
rect 4490 31531 4515 31587
rect 4571 31531 4596 31587
rect 4652 31531 4677 31587
rect 4733 31531 4758 31587
rect 4815 31584 4829 31636
rect 4895 31611 4920 31667
rect 4976 31611 5001 31667
rect 5057 31611 5082 31667
rect 5138 31611 5163 31667
rect 4881 31587 5163 31611
rect 4814 31566 4839 31584
rect 2724 31514 3101 31531
rect 3153 31514 3167 31531
rect 3219 31514 3655 31531
rect 3707 31514 3721 31531
rect 3773 31514 4209 31531
rect 4261 31514 4275 31531
rect 4327 31514 4763 31531
rect 4815 31514 4829 31566
rect 4895 31531 4920 31587
rect 4976 31531 5001 31587
rect 5057 31531 5082 31587
rect 5138 31531 5163 31587
rect 4881 31514 5163 31531
rect 2724 31507 5163 31514
rect 2724 31451 2733 31507
rect 2789 31451 2814 31507
rect 2870 31451 2895 31507
rect 2951 31451 2976 31507
rect 3032 31451 3057 31507
rect 3113 31496 3138 31507
rect 3194 31496 3219 31507
rect 3275 31451 3300 31507
rect 3356 31451 3381 31507
rect 3437 31451 3462 31507
rect 3518 31451 3543 31507
rect 3599 31451 3624 31507
rect 3680 31496 3705 31507
rect 3761 31496 3786 31507
rect 3773 31451 3786 31496
rect 3842 31451 3867 31507
rect 3923 31451 3948 31507
rect 4004 31451 4029 31507
rect 4085 31451 4110 31507
rect 4166 31451 4191 31507
rect 4247 31496 4272 31507
rect 4261 31451 4272 31496
rect 4328 31451 4353 31507
rect 4409 31451 4434 31507
rect 4490 31451 4515 31507
rect 4571 31451 4596 31507
rect 4652 31451 4677 31507
rect 4733 31451 4758 31507
rect 4814 31496 4839 31507
rect 2724 31444 3101 31451
rect 3153 31444 3167 31451
rect 3219 31444 3655 31451
rect 3707 31444 3721 31451
rect 3773 31444 4209 31451
rect 4261 31444 4275 31451
rect 4327 31444 4763 31451
rect 4815 31444 4829 31496
rect 4895 31451 4920 31507
rect 4976 31451 5001 31507
rect 5057 31451 5082 31507
rect 5138 31451 5163 31507
rect 4881 31444 5163 31451
rect 2724 31427 5163 31444
rect 2724 31371 2733 31427
rect 2789 31371 2814 31427
rect 2870 31371 2895 31427
rect 2951 31371 2976 31427
rect 3032 31371 3057 31427
rect 3113 31426 3138 31427
rect 3194 31426 3219 31427
rect 3113 31371 3138 31374
rect 3194 31371 3219 31374
rect 3275 31371 3300 31427
rect 3356 31371 3381 31427
rect 3437 31371 3462 31427
rect 3518 31371 3543 31427
rect 3599 31371 3624 31427
rect 3680 31426 3705 31427
rect 3761 31426 3786 31427
rect 3773 31374 3786 31426
rect 3680 31371 3705 31374
rect 3761 31371 3786 31374
rect 3842 31371 3867 31427
rect 3923 31371 3948 31427
rect 4004 31371 4029 31427
rect 4085 31371 4110 31427
rect 4166 31371 4191 31427
rect 4247 31426 4272 31427
rect 4261 31374 4272 31426
rect 4247 31371 4272 31374
rect 4328 31371 4353 31427
rect 4409 31371 4434 31427
rect 4490 31371 4515 31427
rect 4571 31371 4596 31427
rect 4652 31371 4677 31427
rect 4733 31371 4758 31427
rect 4814 31426 4839 31427
rect 4815 31374 4829 31426
rect 4814 31371 4839 31374
rect 4895 31371 4920 31427
rect 4976 31371 5001 31427
rect 5057 31371 5082 31427
rect 5138 31371 5163 31427
rect 5299 31982 7651 31987
rect 5299 31930 5317 31982
rect 5369 31930 5383 31982
rect 5435 31930 5871 31982
rect 5923 31930 5937 31982
rect 5989 31930 6425 31982
rect 6477 31930 6491 31982
rect 6543 31930 6979 31982
rect 7031 31930 7045 31982
rect 7097 31930 7533 31982
rect 7585 31930 7599 31982
rect 5299 31913 7651 31930
rect 5299 31861 5317 31913
rect 5369 31861 5383 31913
rect 5435 31861 5871 31913
rect 5923 31861 5937 31913
rect 5989 31861 6425 31913
rect 6477 31861 6491 31913
rect 6543 31861 6979 31913
rect 7031 31861 7045 31913
rect 7097 31861 7533 31913
rect 7585 31861 7599 31913
rect 5299 31844 7651 31861
rect 5299 31792 5317 31844
rect 5369 31792 5383 31844
rect 5435 31792 5871 31844
rect 5923 31792 5937 31844
rect 5989 31792 6425 31844
rect 6477 31792 6491 31844
rect 6543 31792 6979 31844
rect 7031 31792 7045 31844
rect 7097 31792 7533 31844
rect 7585 31792 7599 31844
rect 5299 31775 7651 31792
rect 5299 31723 5317 31775
rect 5369 31723 5383 31775
rect 5435 31723 5871 31775
rect 5923 31723 5937 31775
rect 5989 31723 6425 31775
rect 6477 31723 6491 31775
rect 6543 31723 6979 31775
rect 7031 31723 7045 31775
rect 7097 31723 7533 31775
rect 7585 31723 7599 31775
rect 5299 31706 7651 31723
rect 5299 31654 5317 31706
rect 5369 31654 5383 31706
rect 5435 31654 5871 31706
rect 5923 31654 5937 31706
rect 5989 31654 6425 31706
rect 6477 31654 6491 31706
rect 6543 31654 6979 31706
rect 7031 31654 7045 31706
rect 7097 31654 7533 31706
rect 7585 31654 7599 31706
rect 5299 31636 7651 31654
rect 5299 31584 5317 31636
rect 5369 31584 5383 31636
rect 5435 31584 5871 31636
rect 5923 31584 5937 31636
rect 5989 31584 6425 31636
rect 6477 31584 6491 31636
rect 6543 31584 6979 31636
rect 7031 31584 7045 31636
rect 7097 31584 7533 31636
rect 7585 31584 7599 31636
rect 5299 31566 7651 31584
rect 5299 31514 5317 31566
rect 5369 31514 5383 31566
rect 5435 31514 5871 31566
rect 5923 31514 5937 31566
rect 5989 31514 6425 31566
rect 6477 31514 6491 31566
rect 6543 31514 6979 31566
rect 7031 31514 7045 31566
rect 7097 31514 7533 31566
rect 7585 31514 7599 31566
rect 5299 31496 7651 31514
rect 5299 31444 5317 31496
rect 5369 31444 5383 31496
rect 5435 31444 5871 31496
rect 5923 31444 5937 31496
rect 5989 31444 6425 31496
rect 6477 31444 6491 31496
rect 6543 31444 6979 31496
rect 7031 31444 7045 31496
rect 7097 31444 7533 31496
rect 7585 31444 7599 31496
rect 5299 31426 7651 31444
rect 5299 31374 5317 31426
rect 5369 31374 5383 31426
rect 5435 31374 5871 31426
rect 5923 31374 5937 31426
rect 5989 31374 6425 31426
rect 6477 31374 6491 31426
rect 6543 31374 6979 31426
rect 7031 31374 7045 31426
rect 7097 31374 7533 31426
rect 7585 31374 7599 31426
rect 5299 31371 7651 31374
rect 2724 31368 7651 31371
rect 2270 30724 8222 30730
rect 2322 30672 2392 30724
rect 2444 30720 5613 30724
rect 5669 30720 5696 30724
rect 2444 30672 2824 30720
rect 2270 30668 2824 30672
rect 2876 30668 2890 30720
rect 2942 30668 3378 30720
rect 3430 30668 3444 30720
rect 3496 30668 3932 30720
rect 3984 30668 3998 30720
rect 4050 30668 4486 30720
rect 4538 30668 4552 30720
rect 4604 30668 5040 30720
rect 5092 30668 5106 30720
rect 5158 30668 5594 30720
rect 5752 30668 5779 30724
rect 5835 30668 5861 30724
rect 5917 30668 5943 30724
rect 5999 30668 6025 30724
rect 6081 30668 6107 30724
rect 6163 30720 6189 30724
rect 6245 30720 6271 30724
rect 6266 30668 6271 30720
rect 6327 30668 6353 30724
rect 6409 30668 6435 30724
rect 6491 30668 6517 30724
rect 6573 30668 6599 30724
rect 6655 30668 6681 30724
rect 6737 30720 6763 30724
rect 6819 30720 6845 30724
rect 6754 30668 6763 30720
rect 6820 30668 6845 30720
rect 6901 30668 6927 30724
rect 6983 30668 7009 30724
rect 7065 30668 7091 30724
rect 7147 30668 7173 30724
rect 7229 30668 7255 30724
rect 7311 30720 7337 30724
rect 7311 30668 7322 30720
rect 7393 30668 7419 30724
rect 7475 30668 7501 30724
rect 7557 30668 7583 30724
rect 7639 30668 7665 30724
rect 7721 30668 7747 30724
rect 7803 30720 7829 30724
rect 7885 30720 7911 30724
rect 7803 30668 7810 30720
rect 7967 30668 7993 30724
rect 8049 30668 8075 30672
rect 8131 30668 8157 30724
rect 8221 30672 8222 30724
rect 8213 30668 8222 30672
rect 2270 30655 8222 30668
rect 2322 30603 2392 30655
rect 2444 30651 8047 30655
rect 2444 30603 2824 30651
rect 2270 30599 2824 30603
rect 2876 30599 2890 30651
rect 2942 30599 3378 30651
rect 3430 30599 3444 30651
rect 3496 30599 3932 30651
rect 3984 30599 3998 30651
rect 4050 30599 4486 30651
rect 4538 30599 4552 30651
rect 4604 30599 5040 30651
rect 5092 30599 5106 30651
rect 5158 30599 5594 30651
rect 5646 30644 5660 30651
rect 5712 30644 6148 30651
rect 6200 30644 6214 30651
rect 6266 30644 6702 30651
rect 6754 30644 6768 30651
rect 6820 30644 7256 30651
rect 7308 30644 7322 30651
rect 7374 30644 7810 30651
rect 7862 30644 7876 30651
rect 7928 30644 8047 30651
rect 8099 30644 8169 30655
rect 2270 30588 5613 30599
rect 5669 30588 5696 30599
rect 5752 30588 5779 30644
rect 5835 30588 5861 30644
rect 5917 30588 5943 30644
rect 5999 30588 6025 30644
rect 6081 30588 6107 30644
rect 6266 30599 6271 30644
rect 6163 30588 6189 30599
rect 6245 30588 6271 30599
rect 6327 30588 6353 30644
rect 6409 30588 6435 30644
rect 6491 30588 6517 30644
rect 6573 30588 6599 30644
rect 6655 30588 6681 30644
rect 6754 30599 6763 30644
rect 6820 30599 6845 30644
rect 6737 30588 6763 30599
rect 6819 30588 6845 30599
rect 6901 30588 6927 30644
rect 6983 30588 7009 30644
rect 7065 30588 7091 30644
rect 7147 30588 7173 30644
rect 7229 30588 7255 30644
rect 7311 30599 7322 30644
rect 7311 30588 7337 30599
rect 7393 30588 7419 30644
rect 7475 30588 7501 30644
rect 7557 30588 7583 30644
rect 7639 30588 7665 30644
rect 7721 30588 7747 30644
rect 7803 30599 7810 30644
rect 7803 30588 7829 30599
rect 7885 30588 7911 30599
rect 7967 30588 7993 30644
rect 8049 30588 8075 30603
rect 8131 30588 8157 30644
rect 8221 30603 8222 30655
rect 8213 30588 8222 30603
rect 2270 30586 8222 30588
rect 2322 30534 2392 30586
rect 2444 30582 8047 30586
rect 2444 30534 2824 30582
rect 2270 30530 2824 30534
rect 2876 30530 2890 30582
rect 2942 30530 3378 30582
rect 3430 30530 3444 30582
rect 3496 30530 3932 30582
rect 3984 30530 3998 30582
rect 4050 30530 4486 30582
rect 4538 30530 4552 30582
rect 4604 30530 5040 30582
rect 5092 30530 5106 30582
rect 5158 30530 5594 30582
rect 5646 30564 5660 30582
rect 5712 30564 6148 30582
rect 6200 30564 6214 30582
rect 6266 30564 6702 30582
rect 6754 30564 6768 30582
rect 6820 30564 7256 30582
rect 7308 30564 7322 30582
rect 7374 30564 7810 30582
rect 7862 30564 7876 30582
rect 7928 30564 8047 30582
rect 8099 30564 8169 30586
rect 2270 30517 5613 30530
rect 2322 30465 2392 30517
rect 2444 30513 5613 30517
rect 5669 30513 5696 30530
rect 2444 30465 2824 30513
rect 2270 30461 2824 30465
rect 2876 30461 2890 30513
rect 2942 30461 3378 30513
rect 3430 30461 3444 30513
rect 3496 30461 3932 30513
rect 3984 30461 3998 30513
rect 4050 30461 4486 30513
rect 4538 30461 4552 30513
rect 4604 30461 5040 30513
rect 5092 30461 5106 30513
rect 5158 30461 5594 30513
rect 5752 30508 5779 30564
rect 5835 30508 5861 30564
rect 5917 30508 5943 30564
rect 5999 30508 6025 30564
rect 6081 30508 6107 30564
rect 6266 30530 6271 30564
rect 6163 30513 6189 30530
rect 6245 30513 6271 30530
rect 6266 30508 6271 30513
rect 6327 30508 6353 30564
rect 6409 30508 6435 30564
rect 6491 30508 6517 30564
rect 6573 30508 6599 30564
rect 6655 30508 6681 30564
rect 6754 30530 6763 30564
rect 6820 30530 6845 30564
rect 6737 30513 6763 30530
rect 6819 30513 6845 30530
rect 6754 30508 6763 30513
rect 6820 30508 6845 30513
rect 6901 30508 6927 30564
rect 6983 30508 7009 30564
rect 7065 30508 7091 30564
rect 7147 30508 7173 30564
rect 7229 30508 7255 30564
rect 7311 30530 7322 30564
rect 7311 30513 7337 30530
rect 7311 30508 7322 30513
rect 7393 30508 7419 30564
rect 7475 30508 7501 30564
rect 7557 30508 7583 30564
rect 7639 30508 7665 30564
rect 7721 30508 7747 30564
rect 7803 30530 7810 30564
rect 7803 30513 7829 30530
rect 7885 30513 7911 30530
rect 7803 30508 7810 30513
rect 7967 30508 7993 30564
rect 8049 30517 8075 30534
rect 8131 30508 8157 30564
rect 8221 30534 8222 30586
rect 8213 30517 8222 30534
rect 5646 30484 5660 30508
rect 5712 30484 6148 30508
rect 6200 30484 6214 30508
rect 6266 30484 6702 30508
rect 6754 30484 6768 30508
rect 6820 30484 7256 30508
rect 7308 30484 7322 30508
rect 7374 30484 7810 30508
rect 7862 30484 7876 30508
rect 7928 30484 8047 30508
rect 8099 30484 8169 30508
rect 2270 30448 5613 30461
rect 2322 30396 2392 30448
rect 2444 30444 5613 30448
rect 5669 30444 5696 30461
rect 2444 30396 2824 30444
rect 2270 30392 2824 30396
rect 2876 30392 2890 30444
rect 2942 30392 3378 30444
rect 3430 30392 3444 30444
rect 3496 30392 3932 30444
rect 3984 30392 3998 30444
rect 4050 30392 4486 30444
rect 4538 30392 4552 30444
rect 4604 30392 5040 30444
rect 5092 30392 5106 30444
rect 5158 30392 5594 30444
rect 5752 30428 5779 30484
rect 5835 30428 5861 30484
rect 5917 30428 5943 30484
rect 5999 30428 6025 30484
rect 6081 30428 6107 30484
rect 6266 30461 6271 30484
rect 6163 30444 6189 30461
rect 6245 30444 6271 30461
rect 6266 30428 6271 30444
rect 6327 30428 6353 30484
rect 6409 30428 6435 30484
rect 6491 30428 6517 30484
rect 6573 30428 6599 30484
rect 6655 30428 6681 30484
rect 6754 30461 6763 30484
rect 6820 30461 6845 30484
rect 6737 30444 6763 30461
rect 6819 30444 6845 30461
rect 6754 30428 6763 30444
rect 6820 30428 6845 30444
rect 6901 30428 6927 30484
rect 6983 30428 7009 30484
rect 7065 30428 7091 30484
rect 7147 30428 7173 30484
rect 7229 30428 7255 30484
rect 7311 30461 7322 30484
rect 7311 30444 7337 30461
rect 7311 30428 7322 30444
rect 7393 30428 7419 30484
rect 7475 30428 7501 30484
rect 7557 30428 7583 30484
rect 7639 30428 7665 30484
rect 7721 30428 7747 30484
rect 7803 30461 7810 30484
rect 7803 30444 7829 30461
rect 7885 30444 7911 30461
rect 7803 30428 7810 30444
rect 7967 30428 7993 30484
rect 8049 30448 8075 30465
rect 8131 30428 8157 30484
rect 8221 30465 8222 30517
rect 8213 30448 8222 30465
rect 5646 30404 5660 30428
rect 5712 30404 6148 30428
rect 6200 30404 6214 30428
rect 6266 30404 6702 30428
rect 6754 30404 6768 30428
rect 6820 30404 7256 30428
rect 7308 30404 7322 30428
rect 7374 30404 7810 30428
rect 7862 30404 7876 30428
rect 7928 30404 8047 30428
rect 8099 30404 8169 30428
rect 2270 30378 5613 30392
rect 2322 30326 2392 30378
rect 2444 30375 5613 30378
rect 5669 30375 5696 30392
rect 2444 30326 2824 30375
rect 2270 30323 2824 30326
rect 2876 30323 2890 30375
rect 2942 30323 3378 30375
rect 3430 30323 3444 30375
rect 3496 30323 3932 30375
rect 3984 30323 3998 30375
rect 4050 30323 4486 30375
rect 4538 30323 4552 30375
rect 4604 30323 5040 30375
rect 5092 30323 5106 30375
rect 5158 30323 5594 30375
rect 5752 30348 5779 30404
rect 5835 30348 5861 30404
rect 5917 30348 5943 30404
rect 5999 30348 6025 30404
rect 6081 30348 6107 30404
rect 6266 30392 6271 30404
rect 6163 30375 6189 30392
rect 6245 30375 6271 30392
rect 6266 30348 6271 30375
rect 6327 30348 6353 30404
rect 6409 30348 6435 30404
rect 6491 30348 6517 30404
rect 6573 30348 6599 30404
rect 6655 30348 6681 30404
rect 6754 30392 6763 30404
rect 6820 30392 6845 30404
rect 6737 30375 6763 30392
rect 6819 30375 6845 30392
rect 6754 30348 6763 30375
rect 6820 30348 6845 30375
rect 6901 30348 6927 30404
rect 6983 30348 7009 30404
rect 7065 30348 7091 30404
rect 7147 30348 7173 30404
rect 7229 30348 7255 30404
rect 7311 30392 7322 30404
rect 7311 30375 7337 30392
rect 7311 30348 7322 30375
rect 7393 30348 7419 30404
rect 7475 30348 7501 30404
rect 7557 30348 7583 30404
rect 7639 30348 7665 30404
rect 7721 30348 7747 30404
rect 7803 30392 7810 30404
rect 7803 30375 7829 30392
rect 7885 30375 7911 30392
rect 7803 30348 7810 30375
rect 7967 30348 7993 30404
rect 8049 30378 8075 30396
rect 8131 30348 8157 30404
rect 8221 30396 8222 30448
rect 8213 30378 8222 30396
rect 5646 30324 5660 30348
rect 5712 30324 6148 30348
rect 6200 30324 6214 30348
rect 6266 30324 6702 30348
rect 6754 30324 6768 30348
rect 6820 30324 7256 30348
rect 7308 30324 7322 30348
rect 7374 30324 7810 30348
rect 7862 30324 7876 30348
rect 7928 30326 8047 30348
rect 8099 30326 8169 30348
rect 8221 30326 8222 30378
rect 7928 30324 8222 30326
rect 2270 30308 5613 30323
rect 2322 30256 2392 30308
rect 2444 30306 5613 30308
rect 5669 30306 5696 30323
rect 2444 30256 2824 30306
rect 2270 30254 2824 30256
rect 2876 30254 2890 30306
rect 2942 30254 3378 30306
rect 3430 30254 3444 30306
rect 3496 30254 3932 30306
rect 3984 30254 3998 30306
rect 4050 30254 4486 30306
rect 4538 30254 4552 30306
rect 4604 30254 5040 30306
rect 5092 30254 5106 30306
rect 5158 30254 5594 30306
rect 5752 30268 5779 30324
rect 5835 30268 5861 30324
rect 5917 30268 5943 30324
rect 5999 30268 6025 30324
rect 6081 30268 6107 30324
rect 6266 30323 6271 30324
rect 6163 30306 6189 30323
rect 6245 30306 6271 30323
rect 6266 30268 6271 30306
rect 6327 30268 6353 30324
rect 6409 30268 6435 30324
rect 6491 30268 6517 30324
rect 6573 30268 6599 30324
rect 6655 30268 6681 30324
rect 6754 30323 6763 30324
rect 6820 30323 6845 30324
rect 6737 30306 6763 30323
rect 6819 30306 6845 30323
rect 6754 30268 6763 30306
rect 6820 30268 6845 30306
rect 6901 30268 6927 30324
rect 6983 30268 7009 30324
rect 7065 30268 7091 30324
rect 7147 30268 7173 30324
rect 7229 30268 7255 30324
rect 7311 30323 7322 30324
rect 7311 30306 7337 30323
rect 7311 30268 7322 30306
rect 7393 30268 7419 30324
rect 7475 30268 7501 30324
rect 7557 30268 7583 30324
rect 7639 30268 7665 30324
rect 7721 30268 7747 30324
rect 7803 30323 7810 30324
rect 7803 30306 7829 30323
rect 7885 30306 7911 30323
rect 7803 30268 7810 30306
rect 7967 30268 7993 30324
rect 8049 30308 8075 30324
rect 8131 30268 8157 30324
rect 8213 30308 8222 30324
rect 5646 30254 5660 30268
rect 5712 30254 6148 30268
rect 6200 30254 6214 30268
rect 6266 30254 6702 30268
rect 6754 30254 6768 30268
rect 6820 30254 7256 30268
rect 7308 30254 7322 30268
rect 7374 30254 7810 30268
rect 7862 30254 7876 30268
rect 7928 30256 8047 30268
rect 8099 30256 8169 30268
rect 8221 30256 8222 30308
rect 7928 30254 8222 30256
rect 2270 30244 8222 30254
rect 2270 30238 5613 30244
rect 2322 30186 2392 30238
rect 2444 30236 5613 30238
rect 5669 30236 5696 30244
rect 2444 30186 2824 30236
rect 2270 30184 2824 30186
rect 2876 30184 2890 30236
rect 2942 30184 3378 30236
rect 3430 30184 3444 30236
rect 3496 30184 3932 30236
rect 3984 30184 3998 30236
rect 4050 30184 4486 30236
rect 4538 30184 4552 30236
rect 4604 30184 5040 30236
rect 5092 30184 5106 30236
rect 5158 30184 5594 30236
rect 5752 30188 5779 30244
rect 5835 30188 5861 30244
rect 5917 30188 5943 30244
rect 5999 30188 6025 30244
rect 6081 30188 6107 30244
rect 6163 30236 6189 30244
rect 6245 30236 6271 30244
rect 6266 30188 6271 30236
rect 6327 30188 6353 30244
rect 6409 30188 6435 30244
rect 6491 30188 6517 30244
rect 6573 30188 6599 30244
rect 6655 30188 6681 30244
rect 6737 30236 6763 30244
rect 6819 30236 6845 30244
rect 6754 30188 6763 30236
rect 6820 30188 6845 30236
rect 6901 30188 6927 30244
rect 6983 30188 7009 30244
rect 7065 30188 7091 30244
rect 7147 30188 7173 30244
rect 7229 30188 7255 30244
rect 7311 30236 7337 30244
rect 7311 30188 7322 30236
rect 7393 30188 7419 30244
rect 7475 30188 7501 30244
rect 7557 30188 7583 30244
rect 7639 30188 7665 30244
rect 7721 30188 7747 30244
rect 7803 30236 7829 30244
rect 7885 30236 7911 30244
rect 7803 30188 7810 30236
rect 7967 30188 7993 30244
rect 8049 30238 8075 30244
rect 8131 30188 8157 30244
rect 8213 30238 8222 30244
rect 5646 30184 5660 30188
rect 5712 30184 6148 30188
rect 6200 30184 6214 30188
rect 6266 30184 6702 30188
rect 6754 30184 6768 30188
rect 6820 30184 7256 30188
rect 7308 30184 7322 30188
rect 7374 30184 7810 30188
rect 7862 30184 7876 30188
rect 7928 30186 8047 30188
rect 8099 30186 8169 30188
rect 8221 30186 8222 30238
rect 7928 30184 8222 30186
rect 2270 30168 8222 30184
rect 2322 30116 2392 30168
rect 2444 30166 8047 30168
rect 2444 30116 2824 30166
rect 2270 30114 2824 30116
rect 2876 30114 2890 30166
rect 2942 30114 3378 30166
rect 3430 30114 3444 30166
rect 3496 30114 3932 30166
rect 3984 30114 3998 30166
rect 4050 30114 4486 30166
rect 4538 30114 4552 30166
rect 4604 30114 5040 30166
rect 5092 30114 5106 30166
rect 5158 30114 5594 30166
rect 5646 30164 5660 30166
rect 5712 30164 6148 30166
rect 6200 30164 6214 30166
rect 6266 30164 6702 30166
rect 6754 30164 6768 30166
rect 6820 30164 7256 30166
rect 7308 30164 7322 30166
rect 7374 30164 7810 30166
rect 7862 30164 7876 30166
rect 7928 30164 8047 30166
rect 8099 30164 8169 30168
rect 2270 30108 5613 30114
rect 5669 30108 5696 30114
rect 5752 30108 5779 30164
rect 5835 30108 5861 30164
rect 5917 30108 5943 30164
rect 5999 30108 6025 30164
rect 6081 30108 6107 30164
rect 6266 30114 6271 30164
rect 6163 30108 6189 30114
rect 6245 30108 6271 30114
rect 6327 30108 6353 30164
rect 6409 30108 6435 30164
rect 6491 30108 6517 30164
rect 6573 30108 6599 30164
rect 6655 30108 6681 30164
rect 6754 30114 6763 30164
rect 6820 30114 6845 30164
rect 6737 30108 6763 30114
rect 6819 30108 6845 30114
rect 6901 30108 6927 30164
rect 6983 30108 7009 30164
rect 7065 30108 7091 30164
rect 7147 30108 7173 30164
rect 7229 30108 7255 30164
rect 7311 30114 7322 30164
rect 7311 30108 7337 30114
rect 7393 30108 7419 30164
rect 7475 30108 7501 30164
rect 7557 30108 7583 30164
rect 7639 30108 7665 30164
rect 7721 30108 7747 30164
rect 7803 30114 7810 30164
rect 7803 30108 7829 30114
rect 7885 30108 7911 30114
rect 7967 30108 7993 30164
rect 8049 30108 8075 30116
rect 8131 30108 8157 30164
rect 8221 30116 8222 30168
rect 8213 30108 8222 30116
rect 2724 29987 7651 29988
rect 2724 29931 2733 29987
rect 2789 29931 2814 29987
rect 2870 29931 2895 29987
rect 2951 29931 2976 29987
rect 3032 29931 3057 29987
rect 3113 29982 3138 29987
rect 3194 29982 3219 29987
rect 3275 29931 3300 29987
rect 3356 29931 3381 29987
rect 3437 29931 3462 29987
rect 3518 29931 3543 29987
rect 3599 29931 3624 29987
rect 3680 29982 3705 29987
rect 3761 29982 3786 29987
rect 3773 29931 3786 29982
rect 3842 29931 3867 29987
rect 3923 29931 3948 29987
rect 4004 29931 4029 29987
rect 4085 29931 4110 29987
rect 4166 29931 4191 29987
rect 4247 29982 4272 29987
rect 4261 29931 4272 29982
rect 4328 29931 4353 29987
rect 4409 29931 4434 29987
rect 4490 29931 4515 29987
rect 4571 29931 4596 29987
rect 4652 29931 4677 29987
rect 4733 29931 4758 29987
rect 4814 29982 4839 29987
rect 2724 29930 3101 29931
rect 3153 29930 3167 29931
rect 3219 29930 3655 29931
rect 3707 29930 3721 29931
rect 3773 29930 4209 29931
rect 4261 29930 4275 29931
rect 4327 29930 4763 29931
rect 4815 29930 4829 29982
rect 4895 29931 4920 29987
rect 4976 29931 5001 29987
rect 5057 29931 5082 29987
rect 5138 29931 5163 29987
rect 4881 29930 5163 29931
rect 2724 29913 5163 29930
rect 2724 29907 3101 29913
rect 3153 29907 3167 29913
rect 3219 29907 3655 29913
rect 3707 29907 3721 29913
rect 3773 29907 4209 29913
rect 4261 29907 4275 29913
rect 4327 29907 4763 29913
rect 2724 29851 2733 29907
rect 2789 29851 2814 29907
rect 2870 29851 2895 29907
rect 2951 29851 2976 29907
rect 3032 29851 3057 29907
rect 3113 29851 3138 29861
rect 3194 29851 3219 29861
rect 3275 29851 3300 29907
rect 3356 29851 3381 29907
rect 3437 29851 3462 29907
rect 3518 29851 3543 29907
rect 3599 29851 3624 29907
rect 3773 29861 3786 29907
rect 3680 29851 3705 29861
rect 3761 29851 3786 29861
rect 3842 29851 3867 29907
rect 3923 29851 3948 29907
rect 4004 29851 4029 29907
rect 4085 29851 4110 29907
rect 4166 29851 4191 29907
rect 4261 29861 4272 29907
rect 4247 29851 4272 29861
rect 4328 29851 4353 29907
rect 4409 29851 4434 29907
rect 4490 29851 4515 29907
rect 4571 29851 4596 29907
rect 4652 29851 4677 29907
rect 4733 29851 4758 29907
rect 4815 29861 4829 29913
rect 4881 29907 5163 29913
rect 4814 29851 4839 29861
rect 4895 29851 4920 29907
rect 4976 29851 5001 29907
rect 5057 29851 5082 29907
rect 5138 29851 5163 29907
rect 2724 29844 5163 29851
rect 2724 29827 3101 29844
rect 3153 29827 3167 29844
rect 3219 29827 3655 29844
rect 3707 29827 3721 29844
rect 3773 29827 4209 29844
rect 4261 29827 4275 29844
rect 4327 29827 4763 29844
rect 2724 29771 2733 29827
rect 2789 29771 2814 29827
rect 2870 29771 2895 29827
rect 2951 29771 2976 29827
rect 3032 29771 3057 29827
rect 3113 29775 3138 29792
rect 3194 29775 3219 29792
rect 3275 29771 3300 29827
rect 3356 29771 3381 29827
rect 3437 29771 3462 29827
rect 3518 29771 3543 29827
rect 3599 29771 3624 29827
rect 3773 29792 3786 29827
rect 3680 29775 3705 29792
rect 3761 29775 3786 29792
rect 3773 29771 3786 29775
rect 3842 29771 3867 29827
rect 3923 29771 3948 29827
rect 4004 29771 4029 29827
rect 4085 29771 4110 29827
rect 4166 29771 4191 29827
rect 4261 29792 4272 29827
rect 4247 29775 4272 29792
rect 4261 29771 4272 29775
rect 4328 29771 4353 29827
rect 4409 29771 4434 29827
rect 4490 29771 4515 29827
rect 4571 29771 4596 29827
rect 4652 29771 4677 29827
rect 4733 29771 4758 29827
rect 4815 29792 4829 29844
rect 4881 29827 5163 29844
rect 4814 29775 4839 29792
rect 2724 29747 3101 29771
rect 3153 29747 3167 29771
rect 3219 29747 3655 29771
rect 3707 29747 3721 29771
rect 3773 29747 4209 29771
rect 4261 29747 4275 29771
rect 4327 29747 4763 29771
rect 2724 29691 2733 29747
rect 2789 29691 2814 29747
rect 2870 29691 2895 29747
rect 2951 29691 2976 29747
rect 3032 29691 3057 29747
rect 3113 29706 3138 29723
rect 3194 29706 3219 29723
rect 3275 29691 3300 29747
rect 3356 29691 3381 29747
rect 3437 29691 3462 29747
rect 3518 29691 3543 29747
rect 3599 29691 3624 29747
rect 3773 29723 3786 29747
rect 3680 29706 3705 29723
rect 3761 29706 3786 29723
rect 3773 29691 3786 29706
rect 3842 29691 3867 29747
rect 3923 29691 3948 29747
rect 4004 29691 4029 29747
rect 4085 29691 4110 29747
rect 4166 29691 4191 29747
rect 4261 29723 4272 29747
rect 4247 29706 4272 29723
rect 4261 29691 4272 29706
rect 4328 29691 4353 29747
rect 4409 29691 4434 29747
rect 4490 29691 4515 29747
rect 4571 29691 4596 29747
rect 4652 29691 4677 29747
rect 4733 29691 4758 29747
rect 4815 29723 4829 29775
rect 4895 29771 4920 29827
rect 4976 29771 5001 29827
rect 5057 29771 5082 29827
rect 5138 29771 5163 29827
rect 4881 29747 5163 29771
rect 4814 29706 4839 29723
rect 2724 29667 3101 29691
rect 3153 29667 3167 29691
rect 3219 29667 3655 29691
rect 3707 29667 3721 29691
rect 3773 29667 4209 29691
rect 4261 29667 4275 29691
rect 4327 29667 4763 29691
rect 2724 29611 2733 29667
rect 2789 29611 2814 29667
rect 2870 29611 2895 29667
rect 2951 29611 2976 29667
rect 3032 29611 3057 29667
rect 3113 29636 3138 29654
rect 3194 29636 3219 29654
rect 3275 29611 3300 29667
rect 3356 29611 3381 29667
rect 3437 29611 3462 29667
rect 3518 29611 3543 29667
rect 3599 29611 3624 29667
rect 3773 29654 3786 29667
rect 3680 29636 3705 29654
rect 3761 29636 3786 29654
rect 3773 29611 3786 29636
rect 3842 29611 3867 29667
rect 3923 29611 3948 29667
rect 4004 29611 4029 29667
rect 4085 29611 4110 29667
rect 4166 29611 4191 29667
rect 4261 29654 4272 29667
rect 4247 29636 4272 29654
rect 4261 29611 4272 29636
rect 4328 29611 4353 29667
rect 4409 29611 4434 29667
rect 4490 29611 4515 29667
rect 4571 29611 4596 29667
rect 4652 29611 4677 29667
rect 4733 29611 4758 29667
rect 4815 29654 4829 29706
rect 4895 29691 4920 29747
rect 4976 29691 5001 29747
rect 5057 29691 5082 29747
rect 5138 29691 5163 29747
rect 4881 29667 5163 29691
rect 4814 29636 4839 29654
rect 2724 29587 3101 29611
rect 3153 29587 3167 29611
rect 3219 29587 3655 29611
rect 3707 29587 3721 29611
rect 3773 29587 4209 29611
rect 4261 29587 4275 29611
rect 4327 29587 4763 29611
rect 2724 29531 2733 29587
rect 2789 29531 2814 29587
rect 2870 29531 2895 29587
rect 2951 29531 2976 29587
rect 3032 29531 3057 29587
rect 3113 29566 3138 29584
rect 3194 29566 3219 29584
rect 3275 29531 3300 29587
rect 3356 29531 3381 29587
rect 3437 29531 3462 29587
rect 3518 29531 3543 29587
rect 3599 29531 3624 29587
rect 3773 29584 3786 29587
rect 3680 29566 3705 29584
rect 3761 29566 3786 29584
rect 3773 29531 3786 29566
rect 3842 29531 3867 29587
rect 3923 29531 3948 29587
rect 4004 29531 4029 29587
rect 4085 29531 4110 29587
rect 4166 29531 4191 29587
rect 4261 29584 4272 29587
rect 4247 29566 4272 29584
rect 4261 29531 4272 29566
rect 4328 29531 4353 29587
rect 4409 29531 4434 29587
rect 4490 29531 4515 29587
rect 4571 29531 4596 29587
rect 4652 29531 4677 29587
rect 4733 29531 4758 29587
rect 4815 29584 4829 29636
rect 4895 29611 4920 29667
rect 4976 29611 5001 29667
rect 5057 29611 5082 29667
rect 5138 29611 5163 29667
rect 4881 29587 5163 29611
rect 4814 29566 4839 29584
rect 2724 29514 3101 29531
rect 3153 29514 3167 29531
rect 3219 29514 3655 29531
rect 3707 29514 3721 29531
rect 3773 29514 4209 29531
rect 4261 29514 4275 29531
rect 4327 29514 4763 29531
rect 4815 29514 4829 29566
rect 4895 29531 4920 29587
rect 4976 29531 5001 29587
rect 5057 29531 5082 29587
rect 5138 29531 5163 29587
rect 4881 29514 5163 29531
rect 2724 29507 5163 29514
rect 2724 29451 2733 29507
rect 2789 29451 2814 29507
rect 2870 29451 2895 29507
rect 2951 29451 2976 29507
rect 3032 29451 3057 29507
rect 3113 29496 3138 29507
rect 3194 29496 3219 29507
rect 3275 29451 3300 29507
rect 3356 29451 3381 29507
rect 3437 29451 3462 29507
rect 3518 29451 3543 29507
rect 3599 29451 3624 29507
rect 3680 29496 3705 29507
rect 3761 29496 3786 29507
rect 3773 29451 3786 29496
rect 3842 29451 3867 29507
rect 3923 29451 3948 29507
rect 4004 29451 4029 29507
rect 4085 29451 4110 29507
rect 4166 29451 4191 29507
rect 4247 29496 4272 29507
rect 4261 29451 4272 29496
rect 4328 29451 4353 29507
rect 4409 29451 4434 29507
rect 4490 29451 4515 29507
rect 4571 29451 4596 29507
rect 4652 29451 4677 29507
rect 4733 29451 4758 29507
rect 4814 29496 4839 29507
rect 2724 29444 3101 29451
rect 3153 29444 3167 29451
rect 3219 29444 3655 29451
rect 3707 29444 3721 29451
rect 3773 29444 4209 29451
rect 4261 29444 4275 29451
rect 4327 29444 4763 29451
rect 4815 29444 4829 29496
rect 4895 29451 4920 29507
rect 4976 29451 5001 29507
rect 5057 29451 5082 29507
rect 5138 29451 5163 29507
rect 4881 29444 5163 29451
rect 2724 29427 5163 29444
rect 2724 29371 2733 29427
rect 2789 29371 2814 29427
rect 2870 29371 2895 29427
rect 2951 29371 2976 29427
rect 3032 29371 3057 29427
rect 3113 29426 3138 29427
rect 3194 29426 3219 29427
rect 3113 29371 3138 29374
rect 3194 29371 3219 29374
rect 3275 29371 3300 29427
rect 3356 29371 3381 29427
rect 3437 29371 3462 29427
rect 3518 29371 3543 29427
rect 3599 29371 3624 29427
rect 3680 29426 3705 29427
rect 3761 29426 3786 29427
rect 3773 29374 3786 29426
rect 3680 29371 3705 29374
rect 3761 29371 3786 29374
rect 3842 29371 3867 29427
rect 3923 29371 3948 29427
rect 4004 29371 4029 29427
rect 4085 29371 4110 29427
rect 4166 29371 4191 29427
rect 4247 29426 4272 29427
rect 4261 29374 4272 29426
rect 4247 29371 4272 29374
rect 4328 29371 4353 29427
rect 4409 29371 4434 29427
rect 4490 29371 4515 29427
rect 4571 29371 4596 29427
rect 4652 29371 4677 29427
rect 4733 29371 4758 29427
rect 4814 29426 4839 29427
rect 4815 29374 4829 29426
rect 4814 29371 4839 29374
rect 4895 29371 4920 29427
rect 4976 29371 5001 29427
rect 5057 29371 5082 29427
rect 5138 29371 5163 29427
rect 5299 29982 7651 29987
rect 5299 29930 5317 29982
rect 5369 29930 5383 29982
rect 5435 29930 5871 29982
rect 5923 29930 5937 29982
rect 5989 29930 6425 29982
rect 6477 29930 6491 29982
rect 6543 29930 6979 29982
rect 7031 29930 7045 29982
rect 7097 29930 7533 29982
rect 7585 29930 7599 29982
rect 5299 29913 7651 29930
rect 5299 29861 5317 29913
rect 5369 29861 5383 29913
rect 5435 29861 5871 29913
rect 5923 29861 5937 29913
rect 5989 29861 6425 29913
rect 6477 29861 6491 29913
rect 6543 29861 6979 29913
rect 7031 29861 7045 29913
rect 7097 29861 7533 29913
rect 7585 29861 7599 29913
rect 5299 29844 7651 29861
rect 5299 29792 5317 29844
rect 5369 29792 5383 29844
rect 5435 29792 5871 29844
rect 5923 29792 5937 29844
rect 5989 29792 6425 29844
rect 6477 29792 6491 29844
rect 6543 29792 6979 29844
rect 7031 29792 7045 29844
rect 7097 29792 7533 29844
rect 7585 29792 7599 29844
rect 5299 29775 7651 29792
rect 5299 29723 5317 29775
rect 5369 29723 5383 29775
rect 5435 29723 5871 29775
rect 5923 29723 5937 29775
rect 5989 29723 6425 29775
rect 6477 29723 6491 29775
rect 6543 29723 6979 29775
rect 7031 29723 7045 29775
rect 7097 29723 7533 29775
rect 7585 29723 7599 29775
rect 5299 29706 7651 29723
rect 5299 29654 5317 29706
rect 5369 29654 5383 29706
rect 5435 29654 5871 29706
rect 5923 29654 5937 29706
rect 5989 29654 6425 29706
rect 6477 29654 6491 29706
rect 6543 29654 6979 29706
rect 7031 29654 7045 29706
rect 7097 29654 7533 29706
rect 7585 29654 7599 29706
rect 5299 29636 7651 29654
rect 5299 29584 5317 29636
rect 5369 29584 5383 29636
rect 5435 29584 5871 29636
rect 5923 29584 5937 29636
rect 5989 29584 6425 29636
rect 6477 29584 6491 29636
rect 6543 29584 6979 29636
rect 7031 29584 7045 29636
rect 7097 29584 7533 29636
rect 7585 29584 7599 29636
rect 5299 29566 7651 29584
rect 5299 29514 5317 29566
rect 5369 29514 5383 29566
rect 5435 29514 5871 29566
rect 5923 29514 5937 29566
rect 5989 29514 6425 29566
rect 6477 29514 6491 29566
rect 6543 29514 6979 29566
rect 7031 29514 7045 29566
rect 7097 29514 7533 29566
rect 7585 29514 7599 29566
rect 5299 29496 7651 29514
rect 5299 29444 5317 29496
rect 5369 29444 5383 29496
rect 5435 29444 5871 29496
rect 5923 29444 5937 29496
rect 5989 29444 6425 29496
rect 6477 29444 6491 29496
rect 6543 29444 6979 29496
rect 7031 29444 7045 29496
rect 7097 29444 7533 29496
rect 7585 29444 7599 29496
rect 5299 29426 7651 29444
rect 5299 29374 5317 29426
rect 5369 29374 5383 29426
rect 5435 29374 5871 29426
rect 5923 29374 5937 29426
rect 5989 29374 6425 29426
rect 6477 29374 6491 29426
rect 6543 29374 6979 29426
rect 7031 29374 7045 29426
rect 7097 29374 7533 29426
rect 7585 29374 7599 29426
rect 5299 29371 7651 29374
rect 2724 29368 7651 29371
rect 2270 28724 8222 28730
rect 2322 28672 2392 28724
rect 2444 28720 5613 28724
rect 5669 28720 5696 28724
rect 2444 28672 5040 28720
rect 2270 28668 5040 28672
rect 5092 28668 5106 28720
rect 5158 28668 5594 28720
rect 5752 28668 5779 28724
rect 5835 28668 5861 28724
rect 5917 28668 5943 28724
rect 5999 28668 6025 28724
rect 6081 28668 6107 28724
rect 6163 28720 6189 28724
rect 6245 28720 6271 28724
rect 6266 28668 6271 28720
rect 6327 28668 6353 28724
rect 6409 28668 6435 28724
rect 6491 28668 6517 28724
rect 6573 28668 6599 28724
rect 6655 28668 6681 28724
rect 6737 28720 6763 28724
rect 6819 28720 6845 28724
rect 6754 28668 6763 28720
rect 6820 28668 6845 28720
rect 6901 28668 6927 28724
rect 6983 28668 7009 28724
rect 7065 28668 7091 28724
rect 7147 28668 7173 28724
rect 7229 28668 7255 28724
rect 7311 28720 7337 28724
rect 7311 28668 7322 28720
rect 7393 28668 7419 28724
rect 7475 28668 7501 28724
rect 7557 28668 7583 28724
rect 7639 28668 7665 28724
rect 7721 28668 7747 28724
rect 7803 28720 7829 28724
rect 7885 28720 7911 28724
rect 7803 28668 7810 28720
rect 7967 28668 7993 28724
rect 8049 28668 8075 28672
rect 8131 28668 8157 28724
rect 8221 28672 8222 28724
rect 8213 28668 8222 28672
rect 2270 28655 8222 28668
rect 2322 28603 2392 28655
rect 2444 28651 8047 28655
rect 2444 28603 5040 28651
rect 2270 28599 5040 28603
rect 5092 28599 5106 28651
rect 5158 28599 5594 28651
rect 5646 28644 5660 28651
rect 5712 28644 6148 28651
rect 6200 28644 6214 28651
rect 6266 28644 6702 28651
rect 6754 28644 6768 28651
rect 6820 28644 7256 28651
rect 7308 28644 7322 28651
rect 7374 28644 7810 28651
rect 7862 28644 7876 28651
rect 7928 28644 8047 28651
rect 8099 28644 8169 28655
rect 2270 28588 5613 28599
rect 5669 28588 5696 28599
rect 5752 28588 5779 28644
rect 5835 28588 5861 28644
rect 5917 28588 5943 28644
rect 5999 28588 6025 28644
rect 6081 28588 6107 28644
rect 6266 28599 6271 28644
rect 6163 28588 6189 28599
rect 6245 28588 6271 28599
rect 6327 28588 6353 28644
rect 6409 28588 6435 28644
rect 6491 28588 6517 28644
rect 6573 28588 6599 28644
rect 6655 28588 6681 28644
rect 6754 28599 6763 28644
rect 6820 28599 6845 28644
rect 6737 28588 6763 28599
rect 6819 28588 6845 28599
rect 6901 28588 6927 28644
rect 6983 28588 7009 28644
rect 7065 28588 7091 28644
rect 7147 28588 7173 28644
rect 7229 28588 7255 28644
rect 7311 28599 7322 28644
rect 7311 28588 7337 28599
rect 7393 28588 7419 28644
rect 7475 28588 7501 28644
rect 7557 28588 7583 28644
rect 7639 28588 7665 28644
rect 7721 28588 7747 28644
rect 7803 28599 7810 28644
rect 7803 28588 7829 28599
rect 7885 28588 7911 28599
rect 7967 28588 7993 28644
rect 8049 28588 8075 28603
rect 8131 28588 8157 28644
rect 8221 28603 8222 28655
rect 8213 28588 8222 28603
rect 2270 28586 8222 28588
rect 2322 28534 2392 28586
rect 2444 28582 8047 28586
rect 2444 28534 5040 28582
rect 2270 28530 5040 28534
rect 5092 28530 5106 28582
rect 5158 28530 5594 28582
rect 5646 28564 5660 28582
rect 5712 28564 6148 28582
rect 6200 28564 6214 28582
rect 6266 28564 6702 28582
rect 6754 28564 6768 28582
rect 6820 28564 7256 28582
rect 7308 28564 7322 28582
rect 7374 28564 7810 28582
rect 7862 28564 7876 28582
rect 7928 28564 8047 28582
rect 8099 28564 8169 28586
rect 2270 28517 5613 28530
rect 2322 28465 2392 28517
rect 2444 28513 5613 28517
rect 5669 28513 5696 28530
rect 2444 28465 5040 28513
rect 2270 28461 5040 28465
rect 5092 28461 5106 28513
rect 5158 28461 5594 28513
rect 5752 28508 5779 28564
rect 5835 28508 5861 28564
rect 5917 28508 5943 28564
rect 5999 28508 6025 28564
rect 6081 28508 6107 28564
rect 6266 28530 6271 28564
rect 6163 28513 6189 28530
rect 6245 28513 6271 28530
rect 6266 28508 6271 28513
rect 6327 28508 6353 28564
rect 6409 28508 6435 28564
rect 6491 28508 6517 28564
rect 6573 28508 6599 28564
rect 6655 28508 6681 28564
rect 6754 28530 6763 28564
rect 6820 28530 6845 28564
rect 6737 28513 6763 28530
rect 6819 28513 6845 28530
rect 6754 28508 6763 28513
rect 6820 28508 6845 28513
rect 6901 28508 6927 28564
rect 6983 28508 7009 28564
rect 7065 28508 7091 28564
rect 7147 28508 7173 28564
rect 7229 28508 7255 28564
rect 7311 28530 7322 28564
rect 7311 28513 7337 28530
rect 7311 28508 7322 28513
rect 7393 28508 7419 28564
rect 7475 28508 7501 28564
rect 7557 28508 7583 28564
rect 7639 28508 7665 28564
rect 7721 28508 7747 28564
rect 7803 28530 7810 28564
rect 7803 28513 7829 28530
rect 7885 28513 7911 28530
rect 7803 28508 7810 28513
rect 7967 28508 7993 28564
rect 8049 28517 8075 28534
rect 8131 28508 8157 28564
rect 8221 28534 8222 28586
rect 8213 28517 8222 28534
rect 5646 28484 5660 28508
rect 5712 28484 6148 28508
rect 6200 28484 6214 28508
rect 6266 28484 6702 28508
rect 6754 28484 6768 28508
rect 6820 28484 7256 28508
rect 7308 28484 7322 28508
rect 7374 28484 7810 28508
rect 7862 28484 7876 28508
rect 7928 28484 8047 28508
rect 8099 28484 8169 28508
rect 2270 28448 5613 28461
rect 2322 28396 2392 28448
rect 2444 28444 5613 28448
rect 5669 28444 5696 28461
rect 2444 28396 5040 28444
rect 2270 28392 5040 28396
rect 5092 28392 5106 28444
rect 5158 28392 5594 28444
rect 5752 28428 5779 28484
rect 5835 28428 5861 28484
rect 5917 28428 5943 28484
rect 5999 28428 6025 28484
rect 6081 28428 6107 28484
rect 6266 28461 6271 28484
rect 6163 28444 6189 28461
rect 6245 28444 6271 28461
rect 6266 28428 6271 28444
rect 6327 28428 6353 28484
rect 6409 28428 6435 28484
rect 6491 28428 6517 28484
rect 6573 28428 6599 28484
rect 6655 28428 6681 28484
rect 6754 28461 6763 28484
rect 6820 28461 6845 28484
rect 6737 28444 6763 28461
rect 6819 28444 6845 28461
rect 6754 28428 6763 28444
rect 6820 28428 6845 28444
rect 6901 28428 6927 28484
rect 6983 28428 7009 28484
rect 7065 28428 7091 28484
rect 7147 28428 7173 28484
rect 7229 28428 7255 28484
rect 7311 28461 7322 28484
rect 7311 28444 7337 28461
rect 7311 28428 7322 28444
rect 7393 28428 7419 28484
rect 7475 28428 7501 28484
rect 7557 28428 7583 28484
rect 7639 28428 7665 28484
rect 7721 28428 7747 28484
rect 7803 28461 7810 28484
rect 7803 28444 7829 28461
rect 7885 28444 7911 28461
rect 7803 28428 7810 28444
rect 7967 28428 7993 28484
rect 8049 28448 8075 28465
rect 8131 28428 8157 28484
rect 8221 28465 8222 28517
rect 8213 28448 8222 28465
rect 5646 28404 5660 28428
rect 5712 28404 6148 28428
rect 6200 28404 6214 28428
rect 6266 28404 6702 28428
rect 6754 28404 6768 28428
rect 6820 28404 7256 28428
rect 7308 28404 7322 28428
rect 7374 28404 7810 28428
rect 7862 28404 7876 28428
rect 7928 28404 8047 28428
rect 8099 28404 8169 28428
rect 2270 28378 5613 28392
rect 2322 28326 2392 28378
rect 2444 28375 5613 28378
rect 5669 28375 5696 28392
rect 2444 28326 5040 28375
rect 2270 28323 5040 28326
rect 5092 28323 5106 28375
rect 5158 28323 5594 28375
rect 5752 28348 5779 28404
rect 5835 28348 5861 28404
rect 5917 28348 5943 28404
rect 5999 28348 6025 28404
rect 6081 28348 6107 28404
rect 6266 28392 6271 28404
rect 6163 28375 6189 28392
rect 6245 28375 6271 28392
rect 6266 28348 6271 28375
rect 6327 28348 6353 28404
rect 6409 28348 6435 28404
rect 6491 28348 6517 28404
rect 6573 28348 6599 28404
rect 6655 28348 6681 28404
rect 6754 28392 6763 28404
rect 6820 28392 6845 28404
rect 6737 28375 6763 28392
rect 6819 28375 6845 28392
rect 6754 28348 6763 28375
rect 6820 28348 6845 28375
rect 6901 28348 6927 28404
rect 6983 28348 7009 28404
rect 7065 28348 7091 28404
rect 7147 28348 7173 28404
rect 7229 28348 7255 28404
rect 7311 28392 7322 28404
rect 7311 28375 7337 28392
rect 7311 28348 7322 28375
rect 7393 28348 7419 28404
rect 7475 28348 7501 28404
rect 7557 28348 7583 28404
rect 7639 28348 7665 28404
rect 7721 28348 7747 28404
rect 7803 28392 7810 28404
rect 7803 28375 7829 28392
rect 7885 28375 7911 28392
rect 7803 28348 7810 28375
rect 7967 28348 7993 28404
rect 8049 28378 8075 28396
rect 8131 28348 8157 28404
rect 8221 28396 8222 28448
rect 8213 28378 8222 28396
rect 5646 28324 5660 28348
rect 5712 28324 6148 28348
rect 6200 28324 6214 28348
rect 6266 28324 6702 28348
rect 6754 28324 6768 28348
rect 6820 28324 7256 28348
rect 7308 28324 7322 28348
rect 7374 28324 7810 28348
rect 7862 28324 7876 28348
rect 7928 28326 8047 28348
rect 8099 28326 8169 28348
rect 8221 28326 8222 28378
rect 7928 28324 8222 28326
rect 2270 28308 5613 28323
rect 2322 28256 2392 28308
rect 2444 28306 5613 28308
rect 5669 28306 5696 28323
rect 2444 28256 5040 28306
rect 2270 28254 5040 28256
rect 5092 28254 5106 28306
rect 5158 28254 5594 28306
rect 5752 28268 5779 28324
rect 5835 28268 5861 28324
rect 5917 28268 5943 28324
rect 5999 28268 6025 28324
rect 6081 28268 6107 28324
rect 6266 28323 6271 28324
rect 6163 28306 6189 28323
rect 6245 28306 6271 28323
rect 6266 28268 6271 28306
rect 6327 28268 6353 28324
rect 6409 28268 6435 28324
rect 6491 28268 6517 28324
rect 6573 28268 6599 28324
rect 6655 28268 6681 28324
rect 6754 28323 6763 28324
rect 6820 28323 6845 28324
rect 6737 28306 6763 28323
rect 6819 28306 6845 28323
rect 6754 28268 6763 28306
rect 6820 28268 6845 28306
rect 6901 28268 6927 28324
rect 6983 28268 7009 28324
rect 7065 28268 7091 28324
rect 7147 28268 7173 28324
rect 7229 28268 7255 28324
rect 7311 28323 7322 28324
rect 7311 28306 7337 28323
rect 7311 28268 7322 28306
rect 7393 28268 7419 28324
rect 7475 28268 7501 28324
rect 7557 28268 7583 28324
rect 7639 28268 7665 28324
rect 7721 28268 7747 28324
rect 7803 28323 7810 28324
rect 7803 28306 7829 28323
rect 7885 28306 7911 28323
rect 7803 28268 7810 28306
rect 7967 28268 7993 28324
rect 8049 28308 8075 28324
rect 8131 28268 8157 28324
rect 8213 28308 8222 28324
rect 5646 28254 5660 28268
rect 5712 28254 6148 28268
rect 6200 28254 6214 28268
rect 6266 28254 6702 28268
rect 6754 28254 6768 28268
rect 6820 28254 7256 28268
rect 7308 28254 7322 28268
rect 7374 28254 7810 28268
rect 7862 28254 7876 28268
rect 7928 28256 8047 28268
rect 8099 28256 8169 28268
rect 8221 28256 8222 28308
rect 7928 28254 8222 28256
rect 2270 28244 8222 28254
rect 2270 28238 5613 28244
rect 2322 28186 2392 28238
rect 2444 28236 5613 28238
rect 5669 28236 5696 28244
rect 2444 28186 5040 28236
rect 2270 28184 5040 28186
rect 5092 28184 5106 28236
rect 5158 28184 5594 28236
rect 5752 28188 5779 28244
rect 5835 28188 5861 28244
rect 5917 28188 5943 28244
rect 5999 28188 6025 28244
rect 6081 28188 6107 28244
rect 6163 28236 6189 28244
rect 6245 28236 6271 28244
rect 6266 28188 6271 28236
rect 6327 28188 6353 28244
rect 6409 28188 6435 28244
rect 6491 28188 6517 28244
rect 6573 28188 6599 28244
rect 6655 28188 6681 28244
rect 6737 28236 6763 28244
rect 6819 28236 6845 28244
rect 6754 28188 6763 28236
rect 6820 28188 6845 28236
rect 6901 28188 6927 28244
rect 6983 28188 7009 28244
rect 7065 28188 7091 28244
rect 7147 28188 7173 28244
rect 7229 28188 7255 28244
rect 7311 28236 7337 28244
rect 7311 28188 7322 28236
rect 7393 28188 7419 28244
rect 7475 28188 7501 28244
rect 7557 28188 7583 28244
rect 7639 28188 7665 28244
rect 7721 28188 7747 28244
rect 7803 28236 7829 28244
rect 7885 28236 7911 28244
rect 7803 28188 7810 28236
rect 7967 28188 7993 28244
rect 8049 28238 8075 28244
rect 8131 28188 8157 28244
rect 8213 28238 8222 28244
rect 5646 28184 5660 28188
rect 5712 28184 6148 28188
rect 6200 28184 6214 28188
rect 6266 28184 6702 28188
rect 6754 28184 6768 28188
rect 6820 28184 7256 28188
rect 7308 28184 7322 28188
rect 7374 28184 7810 28188
rect 7862 28184 7876 28188
rect 7928 28186 8047 28188
rect 8099 28186 8169 28188
rect 8221 28186 8222 28238
rect 7928 28184 8222 28186
rect 2270 28168 8222 28184
rect 2322 28116 2392 28168
rect 2444 28166 8047 28168
rect 2444 28116 5040 28166
rect 2270 28114 5040 28116
rect 5092 28114 5106 28166
rect 5158 28114 5594 28166
rect 5646 28164 5660 28166
rect 5712 28164 6148 28166
rect 6200 28164 6214 28166
rect 6266 28164 6702 28166
rect 6754 28164 6768 28166
rect 6820 28164 7256 28166
rect 7308 28164 7322 28166
rect 7374 28164 7810 28166
rect 7862 28164 7876 28166
rect 7928 28164 8047 28166
rect 8099 28164 8169 28168
rect 2270 28108 5613 28114
rect 5669 28108 5696 28114
rect 5752 28108 5779 28164
rect 5835 28108 5861 28164
rect 5917 28108 5943 28164
rect 5999 28108 6025 28164
rect 6081 28108 6107 28164
rect 6266 28114 6271 28164
rect 6163 28108 6189 28114
rect 6245 28108 6271 28114
rect 6327 28108 6353 28164
rect 6409 28108 6435 28164
rect 6491 28108 6517 28164
rect 6573 28108 6599 28164
rect 6655 28108 6681 28164
rect 6754 28114 6763 28164
rect 6820 28114 6845 28164
rect 6737 28108 6763 28114
rect 6819 28108 6845 28114
rect 6901 28108 6927 28164
rect 6983 28108 7009 28164
rect 7065 28108 7091 28164
rect 7147 28108 7173 28164
rect 7229 28108 7255 28164
rect 7311 28114 7322 28164
rect 7311 28108 7337 28114
rect 7393 28108 7419 28164
rect 7475 28108 7501 28164
rect 7557 28108 7583 28164
rect 7639 28108 7665 28164
rect 7721 28108 7747 28164
rect 7803 28114 7810 28164
rect 7803 28108 7829 28114
rect 7885 28108 7911 28114
rect 7967 28108 7993 28164
rect 8049 28108 8075 28116
rect 8131 28108 8157 28164
rect 8221 28116 8222 28168
rect 8213 28108 8222 28116
rect 2724 27987 7651 27988
rect 2724 27931 2733 27987
rect 2789 27931 2814 27987
rect 2870 27931 2895 27987
rect 2951 27931 2976 27987
rect 3032 27931 3057 27987
rect 3113 27931 3138 27987
rect 3194 27931 3219 27987
rect 3275 27931 3300 27987
rect 3356 27931 3381 27987
rect 3437 27931 3462 27987
rect 3518 27931 3543 27987
rect 3599 27931 3624 27987
rect 3680 27931 3705 27987
rect 3761 27931 3786 27987
rect 3842 27931 3867 27987
rect 3923 27931 3948 27987
rect 4004 27931 4029 27987
rect 4085 27931 4110 27987
rect 4166 27931 4191 27987
rect 4247 27931 4272 27987
rect 4328 27931 4353 27987
rect 4409 27931 4434 27987
rect 4490 27931 4515 27987
rect 4571 27931 4596 27987
rect 4652 27931 4677 27987
rect 4733 27931 4758 27987
rect 4814 27931 4839 27987
rect 4895 27931 4920 27987
rect 4976 27931 5001 27987
rect 5057 27931 5082 27987
rect 5138 27931 5163 27987
rect 2724 27907 5163 27931
rect 2724 27851 2733 27907
rect 2789 27851 2814 27907
rect 2870 27851 2895 27907
rect 2951 27851 2976 27907
rect 3032 27851 3057 27907
rect 3113 27851 3138 27907
rect 3194 27851 3219 27907
rect 3275 27851 3300 27907
rect 3356 27851 3381 27907
rect 3437 27851 3462 27907
rect 3518 27851 3543 27907
rect 3599 27851 3624 27907
rect 3680 27851 3705 27907
rect 3761 27851 3786 27907
rect 3842 27851 3867 27907
rect 3923 27851 3948 27907
rect 4004 27851 4029 27907
rect 4085 27851 4110 27907
rect 4166 27851 4191 27907
rect 4247 27851 4272 27907
rect 4328 27851 4353 27907
rect 4409 27851 4434 27907
rect 4490 27851 4515 27907
rect 4571 27851 4596 27907
rect 4652 27851 4677 27907
rect 4733 27851 4758 27907
rect 4814 27851 4839 27907
rect 4895 27851 4920 27907
rect 4976 27851 5001 27907
rect 5057 27851 5082 27907
rect 5138 27851 5163 27907
rect 2724 27827 5163 27851
rect 2724 27771 2733 27827
rect 2789 27771 2814 27827
rect 2870 27771 2895 27827
rect 2951 27771 2976 27827
rect 3032 27771 3057 27827
rect 3113 27771 3138 27827
rect 3194 27771 3219 27827
rect 3275 27771 3300 27827
rect 3356 27771 3381 27827
rect 3437 27771 3462 27827
rect 3518 27771 3543 27827
rect 3599 27771 3624 27827
rect 3680 27771 3705 27827
rect 3761 27771 3786 27827
rect 3842 27771 3867 27827
rect 3923 27771 3948 27827
rect 4004 27771 4029 27827
rect 4085 27771 4110 27827
rect 4166 27771 4191 27827
rect 4247 27771 4272 27827
rect 4328 27771 4353 27827
rect 4409 27771 4434 27827
rect 4490 27771 4515 27827
rect 4571 27771 4596 27827
rect 4652 27771 4677 27827
rect 4733 27771 4758 27827
rect 4814 27771 4839 27827
rect 4895 27771 4920 27827
rect 4976 27771 5001 27827
rect 5057 27771 5082 27827
rect 5138 27771 5163 27827
rect 2724 27747 5163 27771
rect 2724 27691 2733 27747
rect 2789 27691 2814 27747
rect 2870 27691 2895 27747
rect 2951 27691 2976 27747
rect 3032 27691 3057 27747
rect 3113 27691 3138 27747
rect 3194 27691 3219 27747
rect 3275 27691 3300 27747
rect 3356 27691 3381 27747
rect 3437 27691 3462 27747
rect 3518 27691 3543 27747
rect 3599 27691 3624 27747
rect 3680 27691 3705 27747
rect 3761 27691 3786 27747
rect 3842 27691 3867 27747
rect 3923 27691 3948 27747
rect 4004 27691 4029 27747
rect 4085 27691 4110 27747
rect 4166 27691 4191 27747
rect 4247 27691 4272 27747
rect 4328 27691 4353 27747
rect 4409 27691 4434 27747
rect 4490 27691 4515 27747
rect 4571 27691 4596 27747
rect 4652 27691 4677 27747
rect 4733 27691 4758 27747
rect 4814 27691 4839 27747
rect 4895 27691 4920 27747
rect 4976 27691 5001 27747
rect 5057 27691 5082 27747
rect 5138 27691 5163 27747
rect 2724 27667 5163 27691
rect 2724 27611 2733 27667
rect 2789 27611 2814 27667
rect 2870 27611 2895 27667
rect 2951 27611 2976 27667
rect 3032 27611 3057 27667
rect 3113 27611 3138 27667
rect 3194 27611 3219 27667
rect 3275 27611 3300 27667
rect 3356 27611 3381 27667
rect 3437 27611 3462 27667
rect 3518 27611 3543 27667
rect 3599 27611 3624 27667
rect 3680 27611 3705 27667
rect 3761 27611 3786 27667
rect 3842 27611 3867 27667
rect 3923 27611 3948 27667
rect 4004 27611 4029 27667
rect 4085 27611 4110 27667
rect 4166 27611 4191 27667
rect 4247 27611 4272 27667
rect 4328 27611 4353 27667
rect 4409 27611 4434 27667
rect 4490 27611 4515 27667
rect 4571 27611 4596 27667
rect 4652 27611 4677 27667
rect 4733 27611 4758 27667
rect 4814 27611 4839 27667
rect 4895 27611 4920 27667
rect 4976 27611 5001 27667
rect 5057 27611 5082 27667
rect 5138 27611 5163 27667
rect 2724 27587 5163 27611
rect 2724 27531 2733 27587
rect 2789 27531 2814 27587
rect 2870 27531 2895 27587
rect 2951 27531 2976 27587
rect 3032 27531 3057 27587
rect 3113 27531 3138 27587
rect 3194 27531 3219 27587
rect 3275 27531 3300 27587
rect 3356 27531 3381 27587
rect 3437 27531 3462 27587
rect 3518 27531 3543 27587
rect 3599 27531 3624 27587
rect 3680 27531 3705 27587
rect 3761 27531 3786 27587
rect 3842 27531 3867 27587
rect 3923 27531 3948 27587
rect 4004 27531 4029 27587
rect 4085 27531 4110 27587
rect 4166 27531 4191 27587
rect 4247 27531 4272 27587
rect 4328 27531 4353 27587
rect 4409 27531 4434 27587
rect 4490 27531 4515 27587
rect 4571 27531 4596 27587
rect 4652 27531 4677 27587
rect 4733 27531 4758 27587
rect 4814 27531 4839 27587
rect 4895 27531 4920 27587
rect 4976 27531 5001 27587
rect 5057 27531 5082 27587
rect 5138 27531 5163 27587
rect 2724 27507 5163 27531
rect 2724 27451 2733 27507
rect 2789 27451 2814 27507
rect 2870 27451 2895 27507
rect 2951 27451 2976 27507
rect 3032 27451 3057 27507
rect 3113 27451 3138 27507
rect 3194 27451 3219 27507
rect 3275 27451 3300 27507
rect 3356 27451 3381 27507
rect 3437 27451 3462 27507
rect 3518 27451 3543 27507
rect 3599 27451 3624 27507
rect 3680 27451 3705 27507
rect 3761 27451 3786 27507
rect 3842 27451 3867 27507
rect 3923 27451 3948 27507
rect 4004 27451 4029 27507
rect 4085 27451 4110 27507
rect 4166 27451 4191 27507
rect 4247 27451 4272 27507
rect 4328 27451 4353 27507
rect 4409 27451 4434 27507
rect 4490 27451 4515 27507
rect 4571 27451 4596 27507
rect 4652 27451 4677 27507
rect 4733 27451 4758 27507
rect 4814 27451 4839 27507
rect 4895 27451 4920 27507
rect 4976 27451 5001 27507
rect 5057 27451 5082 27507
rect 5138 27451 5163 27507
rect 2724 27427 5163 27451
rect 2724 27371 2733 27427
rect 2789 27371 2814 27427
rect 2870 27371 2895 27427
rect 2951 27371 2976 27427
rect 3032 27371 3057 27427
rect 3113 27371 3138 27427
rect 3194 27371 3219 27427
rect 3275 27371 3300 27427
rect 3356 27371 3381 27427
rect 3437 27371 3462 27427
rect 3518 27371 3543 27427
rect 3599 27371 3624 27427
rect 3680 27371 3705 27427
rect 3761 27371 3786 27427
rect 3842 27371 3867 27427
rect 3923 27371 3948 27427
rect 4004 27371 4029 27427
rect 4085 27371 4110 27427
rect 4166 27371 4191 27427
rect 4247 27371 4272 27427
rect 4328 27371 4353 27427
rect 4409 27371 4434 27427
rect 4490 27371 4515 27427
rect 4571 27371 4596 27427
rect 4652 27371 4677 27427
rect 4733 27371 4758 27427
rect 4814 27371 4839 27427
rect 4895 27371 4920 27427
rect 4976 27371 5001 27427
rect 5057 27371 5082 27427
rect 5138 27371 5163 27427
rect 5299 27982 7651 27987
rect 5299 27930 5317 27982
rect 5369 27930 5383 27982
rect 5435 27930 5871 27982
rect 5923 27930 5937 27982
rect 5989 27930 6425 27982
rect 6477 27930 6491 27982
rect 6543 27930 6979 27982
rect 7031 27930 7045 27982
rect 7097 27930 7533 27982
rect 7585 27930 7599 27982
rect 5299 27913 7651 27930
rect 5299 27861 5317 27913
rect 5369 27861 5383 27913
rect 5435 27861 5871 27913
rect 5923 27861 5937 27913
rect 5989 27861 6425 27913
rect 6477 27861 6491 27913
rect 6543 27861 6979 27913
rect 7031 27861 7045 27913
rect 7097 27861 7533 27913
rect 7585 27861 7599 27913
rect 5299 27844 7651 27861
rect 5299 27792 5317 27844
rect 5369 27792 5383 27844
rect 5435 27792 5871 27844
rect 5923 27792 5937 27844
rect 5989 27792 6425 27844
rect 6477 27792 6491 27844
rect 6543 27792 6979 27844
rect 7031 27792 7045 27844
rect 7097 27792 7533 27844
rect 7585 27792 7599 27844
rect 5299 27775 7651 27792
rect 5299 27723 5317 27775
rect 5369 27723 5383 27775
rect 5435 27723 5871 27775
rect 5923 27723 5937 27775
rect 5989 27723 6425 27775
rect 6477 27723 6491 27775
rect 6543 27723 6979 27775
rect 7031 27723 7045 27775
rect 7097 27723 7533 27775
rect 7585 27723 7599 27775
rect 5299 27706 7651 27723
rect 5299 27654 5317 27706
rect 5369 27654 5383 27706
rect 5435 27654 5871 27706
rect 5923 27654 5937 27706
rect 5989 27654 6425 27706
rect 6477 27654 6491 27706
rect 6543 27654 6979 27706
rect 7031 27654 7045 27706
rect 7097 27654 7533 27706
rect 7585 27654 7599 27706
rect 5299 27636 7651 27654
rect 5299 27584 5317 27636
rect 5369 27584 5383 27636
rect 5435 27584 5871 27636
rect 5923 27584 5937 27636
rect 5989 27584 6425 27636
rect 6477 27584 6491 27636
rect 6543 27584 6979 27636
rect 7031 27584 7045 27636
rect 7097 27584 7533 27636
rect 7585 27584 7599 27636
rect 5299 27566 7651 27584
rect 5299 27514 5317 27566
rect 5369 27514 5383 27566
rect 5435 27514 5871 27566
rect 5923 27514 5937 27566
rect 5989 27514 6425 27566
rect 6477 27514 6491 27566
rect 6543 27514 6979 27566
rect 7031 27514 7045 27566
rect 7097 27514 7533 27566
rect 7585 27514 7599 27566
rect 5299 27496 7651 27514
rect 5299 27444 5317 27496
rect 5369 27444 5383 27496
rect 5435 27444 5871 27496
rect 5923 27444 5937 27496
rect 5989 27444 6425 27496
rect 6477 27444 6491 27496
rect 6543 27444 6979 27496
rect 7031 27444 7045 27496
rect 7097 27444 7533 27496
rect 7585 27444 7599 27496
rect 5299 27426 7651 27444
rect 5299 27374 5317 27426
rect 5369 27374 5383 27426
rect 5435 27374 5871 27426
rect 5923 27374 5937 27426
rect 5989 27374 6425 27426
rect 6477 27374 6491 27426
rect 6543 27374 6979 27426
rect 7031 27374 7045 27426
rect 7097 27374 7533 27426
rect 7585 27374 7599 27426
rect 5299 27371 7651 27374
rect 2724 27368 7651 27371
rect 1938 27020 2056 27026
rect 1990 26968 2004 27020
tri 2056 27019 2063 27026 sw
rect 2056 26968 8429 27019
rect 1938 26967 8429 26968
rect 8481 26967 8515 27019
rect 8567 26967 8573 27019
rect 1938 26956 8573 26967
rect 1990 26904 2004 26956
rect 2056 26951 8573 26956
rect 2056 26904 8429 26951
rect 1938 26899 8429 26904
rect 8481 26899 8515 26951
rect 8567 26899 8573 26951
rect 1938 26898 8573 26899
rect 2270 26728 8222 26730
rect 2270 26724 2648 26728
rect 2322 26672 2392 26724
rect 2444 26676 2648 26724
rect 2700 26676 2713 26728
rect 2765 26676 2778 26728
rect 2830 26676 2843 26728
rect 2895 26676 2908 26728
rect 2960 26676 2973 26728
rect 3025 26676 3038 26728
rect 3090 26676 3103 26728
rect 3155 26676 3168 26728
rect 3220 26676 3233 26728
rect 3285 26676 3298 26728
rect 3350 26676 3363 26728
rect 3415 26676 3428 26728
rect 3480 26676 3493 26728
rect 3545 26676 3558 26728
rect 3610 26676 3623 26728
rect 3675 26676 3688 26728
rect 3740 26676 3753 26728
rect 3805 26676 3818 26728
rect 3870 26676 3883 26728
rect 3935 26676 3948 26728
rect 4000 26676 4013 26728
rect 4065 26676 4078 26728
rect 4130 26676 4143 26728
rect 4195 26676 4208 26728
rect 4260 26676 4273 26728
rect 4325 26676 4338 26728
rect 4390 26676 4403 26728
rect 4455 26676 4468 26728
rect 4520 26676 4532 26728
rect 4584 26724 8222 26728
rect 4584 26720 5613 26724
rect 5669 26720 5696 26724
rect 4584 26676 5040 26720
rect 2444 26672 5040 26676
rect 2270 26668 5040 26672
rect 5092 26668 5106 26720
rect 5158 26668 5594 26720
rect 5752 26668 5779 26724
rect 5835 26668 5861 26724
rect 5917 26668 5943 26724
rect 5999 26668 6025 26724
rect 6081 26668 6107 26724
rect 6163 26720 6189 26724
rect 6245 26720 6271 26724
rect 6266 26668 6271 26720
rect 6327 26668 6353 26724
rect 6409 26668 6435 26724
rect 6491 26668 6517 26724
rect 6573 26668 6599 26724
rect 6655 26668 6681 26724
rect 6737 26720 6763 26724
rect 6819 26720 6845 26724
rect 6754 26668 6763 26720
rect 6820 26668 6845 26720
rect 6901 26668 6927 26724
rect 6983 26668 7009 26724
rect 7065 26668 7091 26724
rect 7147 26668 7173 26724
rect 7229 26668 7255 26724
rect 7311 26720 7337 26724
rect 7311 26668 7322 26720
rect 7393 26668 7419 26724
rect 7475 26668 7501 26724
rect 7557 26668 7583 26724
rect 7639 26668 7665 26724
rect 7721 26668 7747 26724
rect 7803 26720 7829 26724
rect 7885 26720 7911 26724
rect 7803 26668 7810 26720
rect 7967 26668 7993 26724
rect 8049 26668 8075 26672
rect 8131 26668 8157 26724
rect 8221 26672 8222 26724
rect 8213 26668 8222 26672
rect 2270 26660 8222 26668
rect 2270 26655 2648 26660
rect 2322 26603 2392 26655
rect 2444 26608 2648 26655
rect 2700 26608 2713 26660
rect 2765 26608 2778 26660
rect 2830 26608 2843 26660
rect 2895 26608 2908 26660
rect 2960 26608 2973 26660
rect 3025 26608 3038 26660
rect 3090 26608 3103 26660
rect 3155 26608 3168 26660
rect 3220 26608 3233 26660
rect 3285 26608 3298 26660
rect 3350 26608 3363 26660
rect 3415 26608 3428 26660
rect 3480 26608 3493 26660
rect 3545 26608 3558 26660
rect 3610 26608 3623 26660
rect 3675 26608 3688 26660
rect 3740 26608 3753 26660
rect 3805 26608 3818 26660
rect 3870 26608 3883 26660
rect 3935 26608 3948 26660
rect 4000 26608 4013 26660
rect 4065 26608 4078 26660
rect 4130 26608 4143 26660
rect 4195 26608 4208 26660
rect 4260 26608 4273 26660
rect 4325 26608 4338 26660
rect 4390 26608 4403 26660
rect 4455 26608 4468 26660
rect 4520 26608 4532 26660
rect 4584 26655 8222 26660
rect 4584 26651 8047 26655
rect 4584 26608 5040 26651
rect 2444 26603 5040 26608
rect 2270 26599 5040 26603
rect 5092 26599 5106 26651
rect 5158 26599 5594 26651
rect 5646 26644 5660 26651
rect 5712 26644 6148 26651
rect 6200 26644 6214 26651
rect 6266 26644 6702 26651
rect 6754 26644 6768 26651
rect 6820 26644 7256 26651
rect 7308 26644 7322 26651
rect 7374 26644 7810 26651
rect 7862 26644 7876 26651
rect 7928 26644 8047 26651
rect 8099 26644 8169 26655
rect 2270 26592 5613 26599
rect 2270 26586 2648 26592
rect 2322 26534 2392 26586
rect 2444 26540 2648 26586
rect 2700 26540 2713 26592
rect 2765 26540 2778 26592
rect 2830 26540 2843 26592
rect 2895 26540 2908 26592
rect 2960 26540 2973 26592
rect 3025 26540 3038 26592
rect 3090 26540 3103 26592
rect 3155 26540 3168 26592
rect 3220 26540 3233 26592
rect 3285 26540 3298 26592
rect 3350 26540 3363 26592
rect 3415 26540 3428 26592
rect 3480 26540 3493 26592
rect 3545 26540 3558 26592
rect 3610 26540 3623 26592
rect 3675 26540 3688 26592
rect 3740 26540 3753 26592
rect 3805 26540 3818 26592
rect 3870 26540 3883 26592
rect 3935 26540 3948 26592
rect 4000 26540 4013 26592
rect 4065 26540 4078 26592
rect 4130 26540 4143 26592
rect 4195 26540 4208 26592
rect 4260 26540 4273 26592
rect 4325 26540 4338 26592
rect 4390 26540 4403 26592
rect 4455 26540 4468 26592
rect 4520 26540 4532 26592
rect 4584 26588 5613 26592
rect 5669 26588 5696 26599
rect 5752 26588 5779 26644
rect 5835 26588 5861 26644
rect 5917 26588 5943 26644
rect 5999 26588 6025 26644
rect 6081 26588 6107 26644
rect 6266 26599 6271 26644
rect 6163 26588 6189 26599
rect 6245 26588 6271 26599
rect 6327 26588 6353 26644
rect 6409 26588 6435 26644
rect 6491 26588 6517 26644
rect 6573 26588 6599 26644
rect 6655 26588 6681 26644
rect 6754 26599 6763 26644
rect 6820 26599 6845 26644
rect 6737 26588 6763 26599
rect 6819 26588 6845 26599
rect 6901 26588 6927 26644
rect 6983 26588 7009 26644
rect 7065 26588 7091 26644
rect 7147 26588 7173 26644
rect 7229 26588 7255 26644
rect 7311 26599 7322 26644
rect 7311 26588 7337 26599
rect 7393 26588 7419 26644
rect 7475 26588 7501 26644
rect 7557 26588 7583 26644
rect 7639 26588 7665 26644
rect 7721 26588 7747 26644
rect 7803 26599 7810 26644
rect 7803 26588 7829 26599
rect 7885 26588 7911 26599
rect 7967 26588 7993 26644
rect 8049 26588 8075 26603
rect 8131 26588 8157 26644
rect 8221 26603 8222 26655
rect 8213 26588 8222 26603
rect 4584 26586 8222 26588
rect 4584 26582 8047 26586
rect 4584 26540 5040 26582
rect 2444 26534 5040 26540
rect 2270 26530 5040 26534
rect 5092 26530 5106 26582
rect 5158 26530 5594 26582
rect 5646 26564 5660 26582
rect 5712 26564 6148 26582
rect 6200 26564 6214 26582
rect 6266 26564 6702 26582
rect 6754 26564 6768 26582
rect 6820 26564 7256 26582
rect 7308 26564 7322 26582
rect 7374 26564 7810 26582
rect 7862 26564 7876 26582
rect 7928 26564 8047 26582
rect 8099 26564 8169 26586
rect 2270 26524 5613 26530
rect 2270 26517 2648 26524
rect 2322 26465 2392 26517
rect 2444 26472 2648 26517
rect 2700 26472 2713 26524
rect 2765 26472 2778 26524
rect 2830 26472 2843 26524
rect 2895 26472 2908 26524
rect 2960 26472 2973 26524
rect 3025 26472 3038 26524
rect 3090 26472 3103 26524
rect 3155 26472 3168 26524
rect 3220 26472 3233 26524
rect 3285 26472 3298 26524
rect 3350 26472 3363 26524
rect 3415 26472 3428 26524
rect 3480 26472 3493 26524
rect 3545 26472 3558 26524
rect 3610 26472 3623 26524
rect 3675 26472 3688 26524
rect 3740 26472 3753 26524
rect 3805 26472 3818 26524
rect 3870 26472 3883 26524
rect 3935 26472 3948 26524
rect 4000 26472 4013 26524
rect 4065 26472 4078 26524
rect 4130 26472 4143 26524
rect 4195 26472 4208 26524
rect 4260 26472 4273 26524
rect 4325 26472 4338 26524
rect 4390 26472 4403 26524
rect 4455 26472 4468 26524
rect 4520 26472 4532 26524
rect 4584 26513 5613 26524
rect 5669 26513 5696 26530
rect 4584 26472 5040 26513
rect 2444 26465 5040 26472
rect 2270 26461 5040 26465
rect 5092 26461 5106 26513
rect 5158 26461 5594 26513
rect 5752 26508 5779 26564
rect 5835 26508 5861 26564
rect 5917 26508 5943 26564
rect 5999 26508 6025 26564
rect 6081 26508 6107 26564
rect 6266 26530 6271 26564
rect 6163 26513 6189 26530
rect 6245 26513 6271 26530
rect 6266 26508 6271 26513
rect 6327 26508 6353 26564
rect 6409 26508 6435 26564
rect 6491 26508 6517 26564
rect 6573 26508 6599 26564
rect 6655 26508 6681 26564
rect 6754 26530 6763 26564
rect 6820 26530 6845 26564
rect 6737 26513 6763 26530
rect 6819 26513 6845 26530
rect 6754 26508 6763 26513
rect 6820 26508 6845 26513
rect 6901 26508 6927 26564
rect 6983 26508 7009 26564
rect 7065 26508 7091 26564
rect 7147 26508 7173 26564
rect 7229 26508 7255 26564
rect 7311 26530 7322 26564
rect 7311 26513 7337 26530
rect 7311 26508 7322 26513
rect 7393 26508 7419 26564
rect 7475 26508 7501 26564
rect 7557 26508 7583 26564
rect 7639 26508 7665 26564
rect 7721 26508 7747 26564
rect 7803 26530 7810 26564
rect 7803 26513 7829 26530
rect 7885 26513 7911 26530
rect 7803 26508 7810 26513
rect 7967 26508 7993 26564
rect 8049 26517 8075 26534
rect 8131 26508 8157 26564
rect 8221 26534 8222 26586
rect 8213 26517 8222 26534
rect 5646 26484 5660 26508
rect 5712 26484 6148 26508
rect 6200 26484 6214 26508
rect 6266 26484 6702 26508
rect 6754 26484 6768 26508
rect 6820 26484 7256 26508
rect 7308 26484 7322 26508
rect 7374 26484 7810 26508
rect 7862 26484 7876 26508
rect 7928 26484 8047 26508
rect 8099 26484 8169 26508
rect 2270 26456 5613 26461
rect 2270 26448 2648 26456
rect 2322 26396 2392 26448
rect 2444 26404 2648 26448
rect 2700 26404 2713 26456
rect 2765 26404 2778 26456
rect 2830 26404 2843 26456
rect 2895 26404 2908 26456
rect 2960 26404 2973 26456
rect 3025 26404 3038 26456
rect 3090 26404 3103 26456
rect 3155 26404 3168 26456
rect 3220 26404 3233 26456
rect 3285 26404 3298 26456
rect 3350 26404 3363 26456
rect 3415 26404 3428 26456
rect 3480 26404 3493 26456
rect 3545 26404 3558 26456
rect 3610 26404 3623 26456
rect 3675 26404 3688 26456
rect 3740 26404 3753 26456
rect 3805 26404 3818 26456
rect 3870 26404 3883 26456
rect 3935 26404 3948 26456
rect 4000 26404 4013 26456
rect 4065 26404 4078 26456
rect 4130 26404 4143 26456
rect 4195 26404 4208 26456
rect 4260 26404 4273 26456
rect 4325 26404 4338 26456
rect 4390 26404 4403 26456
rect 4455 26404 4468 26456
rect 4520 26404 4532 26456
rect 4584 26444 5613 26456
rect 5669 26444 5696 26461
rect 4584 26404 5040 26444
rect 2444 26396 5040 26404
rect 2270 26392 5040 26396
rect 5092 26392 5106 26444
rect 5158 26392 5594 26444
rect 5752 26428 5779 26484
rect 5835 26428 5861 26484
rect 5917 26428 5943 26484
rect 5999 26428 6025 26484
rect 6081 26428 6107 26484
rect 6266 26461 6271 26484
rect 6163 26444 6189 26461
rect 6245 26444 6271 26461
rect 6266 26428 6271 26444
rect 6327 26428 6353 26484
rect 6409 26428 6435 26484
rect 6491 26428 6517 26484
rect 6573 26428 6599 26484
rect 6655 26428 6681 26484
rect 6754 26461 6763 26484
rect 6820 26461 6845 26484
rect 6737 26444 6763 26461
rect 6819 26444 6845 26461
rect 6754 26428 6763 26444
rect 6820 26428 6845 26444
rect 6901 26428 6927 26484
rect 6983 26428 7009 26484
rect 7065 26428 7091 26484
rect 7147 26428 7173 26484
rect 7229 26428 7255 26484
rect 7311 26461 7322 26484
rect 7311 26444 7337 26461
rect 7311 26428 7322 26444
rect 7393 26428 7419 26484
rect 7475 26428 7501 26484
rect 7557 26428 7583 26484
rect 7639 26428 7665 26484
rect 7721 26428 7747 26484
rect 7803 26461 7810 26484
rect 7803 26444 7829 26461
rect 7885 26444 7911 26461
rect 7803 26428 7810 26444
rect 7967 26428 7993 26484
rect 8049 26448 8075 26465
rect 8131 26428 8157 26484
rect 8221 26465 8222 26517
rect 8213 26448 8222 26465
rect 5646 26404 5660 26428
rect 5712 26404 6148 26428
rect 6200 26404 6214 26428
rect 6266 26404 6702 26428
rect 6754 26404 6768 26428
rect 6820 26404 7256 26428
rect 7308 26404 7322 26428
rect 7374 26404 7810 26428
rect 7862 26404 7876 26428
rect 7928 26404 8047 26428
rect 8099 26404 8169 26428
rect 2270 26388 5613 26392
rect 2270 26378 2648 26388
rect 2322 26326 2392 26378
rect 2444 26336 2648 26378
rect 2700 26336 2713 26388
rect 2765 26336 2778 26388
rect 2830 26336 2843 26388
rect 2895 26336 2908 26388
rect 2960 26336 2973 26388
rect 3025 26336 3038 26388
rect 3090 26336 3103 26388
rect 3155 26336 3168 26388
rect 3220 26336 3233 26388
rect 3285 26336 3298 26388
rect 3350 26336 3363 26388
rect 3415 26336 3428 26388
rect 3480 26336 3493 26388
rect 3545 26336 3558 26388
rect 3610 26336 3623 26388
rect 3675 26336 3688 26388
rect 3740 26336 3753 26388
rect 3805 26336 3818 26388
rect 3870 26336 3883 26388
rect 3935 26336 3948 26388
rect 4000 26336 4013 26388
rect 4065 26336 4078 26388
rect 4130 26336 4143 26388
rect 4195 26336 4208 26388
rect 4260 26336 4273 26388
rect 4325 26336 4338 26388
rect 4390 26336 4403 26388
rect 4455 26336 4468 26388
rect 4520 26336 4532 26388
rect 4584 26375 5613 26388
rect 5669 26375 5696 26392
rect 4584 26336 5040 26375
rect 2444 26326 5040 26336
rect 2270 26323 5040 26326
rect 5092 26323 5106 26375
rect 5158 26323 5594 26375
rect 5752 26348 5779 26404
rect 5835 26348 5861 26404
rect 5917 26348 5943 26404
rect 5999 26348 6025 26404
rect 6081 26348 6107 26404
rect 6266 26392 6271 26404
rect 6163 26375 6189 26392
rect 6245 26375 6271 26392
rect 6266 26348 6271 26375
rect 6327 26348 6353 26404
rect 6409 26348 6435 26404
rect 6491 26348 6517 26404
rect 6573 26348 6599 26404
rect 6655 26348 6681 26404
rect 6754 26392 6763 26404
rect 6820 26392 6845 26404
rect 6737 26375 6763 26392
rect 6819 26375 6845 26392
rect 6754 26348 6763 26375
rect 6820 26348 6845 26375
rect 6901 26348 6927 26404
rect 6983 26348 7009 26404
rect 7065 26348 7091 26404
rect 7147 26348 7173 26404
rect 7229 26348 7255 26404
rect 7311 26392 7322 26404
rect 7311 26375 7337 26392
rect 7311 26348 7322 26375
rect 7393 26348 7419 26404
rect 7475 26348 7501 26404
rect 7557 26348 7583 26404
rect 7639 26348 7665 26404
rect 7721 26348 7747 26404
rect 7803 26392 7810 26404
rect 7803 26375 7829 26392
rect 7885 26375 7911 26392
rect 7803 26348 7810 26375
rect 7967 26348 7993 26404
rect 8049 26378 8075 26396
rect 8131 26348 8157 26404
rect 8221 26396 8222 26448
rect 8213 26378 8222 26396
rect 5646 26324 5660 26348
rect 5712 26324 6148 26348
rect 6200 26324 6214 26348
rect 6266 26324 6702 26348
rect 6754 26324 6768 26348
rect 6820 26324 7256 26348
rect 7308 26324 7322 26348
rect 7374 26324 7810 26348
rect 7862 26324 7876 26348
rect 7928 26326 8047 26348
rect 8099 26326 8169 26348
rect 8221 26326 8222 26378
rect 7928 26324 8222 26326
rect 2270 26320 5613 26323
rect 2270 26308 2648 26320
rect 2322 26256 2392 26308
rect 2444 26268 2648 26308
rect 2700 26268 2713 26320
rect 2765 26268 2778 26320
rect 2830 26268 2843 26320
rect 2895 26268 2908 26320
rect 2960 26268 2973 26320
rect 3025 26268 3038 26320
rect 3090 26268 3103 26320
rect 3155 26268 3168 26320
rect 3220 26268 3233 26320
rect 3285 26268 3298 26320
rect 3350 26268 3363 26320
rect 3415 26268 3428 26320
rect 3480 26268 3493 26320
rect 3545 26268 3558 26320
rect 3610 26268 3623 26320
rect 3675 26268 3688 26320
rect 3740 26268 3753 26320
rect 3805 26268 3818 26320
rect 3870 26268 3883 26320
rect 3935 26268 3948 26320
rect 4000 26268 4013 26320
rect 4065 26268 4078 26320
rect 4130 26268 4143 26320
rect 4195 26268 4208 26320
rect 4260 26268 4273 26320
rect 4325 26268 4338 26320
rect 4390 26268 4403 26320
rect 4455 26268 4468 26320
rect 4520 26268 4532 26320
rect 4584 26306 5613 26320
rect 5669 26306 5696 26323
rect 4584 26268 5040 26306
rect 2444 26256 5040 26268
rect 2270 26254 5040 26256
rect 5092 26254 5106 26306
rect 5158 26254 5594 26306
rect 5752 26268 5779 26324
rect 5835 26268 5861 26324
rect 5917 26268 5943 26324
rect 5999 26268 6025 26324
rect 6081 26268 6107 26324
rect 6266 26323 6271 26324
rect 6163 26306 6189 26323
rect 6245 26306 6271 26323
rect 6266 26268 6271 26306
rect 6327 26268 6353 26324
rect 6409 26268 6435 26324
rect 6491 26268 6517 26324
rect 6573 26268 6599 26324
rect 6655 26268 6681 26324
rect 6754 26323 6763 26324
rect 6820 26323 6845 26324
rect 6737 26306 6763 26323
rect 6819 26306 6845 26323
rect 6754 26268 6763 26306
rect 6820 26268 6845 26306
rect 6901 26268 6927 26324
rect 6983 26268 7009 26324
rect 7065 26268 7091 26324
rect 7147 26268 7173 26324
rect 7229 26268 7255 26324
rect 7311 26323 7322 26324
rect 7311 26306 7337 26323
rect 7311 26268 7322 26306
rect 7393 26268 7419 26324
rect 7475 26268 7501 26324
rect 7557 26268 7583 26324
rect 7639 26268 7665 26324
rect 7721 26268 7747 26324
rect 7803 26323 7810 26324
rect 7803 26306 7829 26323
rect 7885 26306 7911 26323
rect 7803 26268 7810 26306
rect 7967 26268 7993 26324
rect 8049 26308 8075 26324
rect 8131 26268 8157 26324
rect 8213 26308 8222 26324
rect 5646 26254 5660 26268
rect 5712 26254 6148 26268
rect 6200 26254 6214 26268
rect 6266 26254 6702 26268
rect 6754 26254 6768 26268
rect 6820 26254 7256 26268
rect 7308 26254 7322 26268
rect 7374 26254 7810 26268
rect 7862 26254 7876 26268
rect 7928 26256 8047 26268
rect 8099 26256 8169 26268
rect 8221 26256 8222 26308
rect 7928 26254 8222 26256
rect 2270 26252 8222 26254
rect 2270 26238 2648 26252
rect 2322 26186 2392 26238
rect 2444 26200 2648 26238
rect 2700 26200 2713 26252
rect 2765 26200 2778 26252
rect 2830 26200 2843 26252
rect 2895 26200 2908 26252
rect 2960 26200 2973 26252
rect 3025 26200 3038 26252
rect 3090 26200 3103 26252
rect 3155 26200 3168 26252
rect 3220 26200 3233 26252
rect 3285 26200 3298 26252
rect 3350 26200 3363 26252
rect 3415 26200 3428 26252
rect 3480 26200 3493 26252
rect 3545 26200 3558 26252
rect 3610 26200 3623 26252
rect 3675 26200 3688 26252
rect 3740 26200 3753 26252
rect 3805 26200 3818 26252
rect 3870 26200 3883 26252
rect 3935 26200 3948 26252
rect 4000 26200 4013 26252
rect 4065 26200 4078 26252
rect 4130 26200 4143 26252
rect 4195 26200 4208 26252
rect 4260 26200 4273 26252
rect 4325 26200 4338 26252
rect 4390 26200 4403 26252
rect 4455 26200 4468 26252
rect 4520 26200 4532 26252
rect 4584 26244 8222 26252
rect 4584 26236 5613 26244
rect 5669 26236 5696 26244
rect 4584 26200 5040 26236
rect 2444 26186 5040 26200
rect 2270 26184 5040 26186
rect 5092 26184 5106 26236
rect 5158 26184 5594 26236
rect 5752 26188 5779 26244
rect 5835 26188 5861 26244
rect 5917 26188 5943 26244
rect 5999 26188 6025 26244
rect 6081 26188 6107 26244
rect 6163 26236 6189 26244
rect 6245 26236 6271 26244
rect 6266 26188 6271 26236
rect 6327 26188 6353 26244
rect 6409 26188 6435 26244
rect 6491 26188 6517 26244
rect 6573 26188 6599 26244
rect 6655 26188 6681 26244
rect 6737 26236 6763 26244
rect 6819 26236 6845 26244
rect 6754 26188 6763 26236
rect 6820 26188 6845 26236
rect 6901 26188 6927 26244
rect 6983 26188 7009 26244
rect 7065 26188 7091 26244
rect 7147 26188 7173 26244
rect 7229 26188 7255 26244
rect 7311 26236 7337 26244
rect 7311 26188 7322 26236
rect 7393 26188 7419 26244
rect 7475 26188 7501 26244
rect 7557 26188 7583 26244
rect 7639 26188 7665 26244
rect 7721 26188 7747 26244
rect 7803 26236 7829 26244
rect 7885 26236 7911 26244
rect 7803 26188 7810 26236
rect 7967 26188 7993 26244
rect 8049 26238 8075 26244
rect 8131 26188 8157 26244
rect 8213 26238 8222 26244
rect 5646 26184 5660 26188
rect 5712 26184 6148 26188
rect 6200 26184 6214 26188
rect 6266 26184 6702 26188
rect 6754 26184 6768 26188
rect 6820 26184 7256 26188
rect 7308 26184 7322 26188
rect 7374 26184 7810 26188
rect 7862 26184 7876 26188
rect 7928 26186 8047 26188
rect 8099 26186 8169 26188
rect 8221 26186 8222 26238
rect 7928 26184 8222 26186
rect 2270 26168 8222 26184
rect 2322 26116 2392 26168
rect 2444 26166 8047 26168
rect 2444 26116 5040 26166
rect 2270 26114 5040 26116
rect 5092 26114 5106 26166
rect 5158 26114 5594 26166
rect 5646 26164 5660 26166
rect 5712 26164 6148 26166
rect 6200 26164 6214 26166
rect 6266 26164 6702 26166
rect 6754 26164 6768 26166
rect 6820 26164 7256 26166
rect 7308 26164 7322 26166
rect 7374 26164 7810 26166
rect 7862 26164 7876 26166
rect 7928 26164 8047 26166
rect 8099 26164 8169 26168
rect 2270 26108 5613 26114
rect 5669 26108 5696 26114
rect 5752 26108 5779 26164
rect 5835 26108 5861 26164
rect 5917 26108 5943 26164
rect 5999 26108 6025 26164
rect 6081 26108 6107 26164
rect 6266 26114 6271 26164
rect 6163 26108 6189 26114
rect 6245 26108 6271 26114
rect 6327 26108 6353 26164
rect 6409 26108 6435 26164
rect 6491 26108 6517 26164
rect 6573 26108 6599 26164
rect 6655 26108 6681 26164
rect 6754 26114 6763 26164
rect 6820 26114 6845 26164
rect 6737 26108 6763 26114
rect 6819 26108 6845 26114
rect 6901 26108 6927 26164
rect 6983 26108 7009 26164
rect 7065 26108 7091 26164
rect 7147 26108 7173 26164
rect 7229 26108 7255 26164
rect 7311 26114 7322 26164
rect 7311 26108 7337 26114
rect 7393 26108 7419 26164
rect 7475 26108 7501 26164
rect 7557 26108 7583 26164
rect 7639 26108 7665 26164
rect 7721 26108 7747 26164
rect 7803 26114 7810 26164
rect 7803 26108 7829 26114
rect 7885 26108 7911 26114
rect 7967 26108 7993 26164
rect 8049 26108 8075 26116
rect 8131 26108 8157 26164
rect 8221 26116 8222 26168
rect 8213 26108 8222 26116
rect 2724 25987 7651 25988
rect 2724 25931 2733 25987
rect 2789 25931 2814 25987
rect 2870 25931 2895 25987
rect 2951 25931 2976 25987
rect 3032 25931 3057 25987
rect 3113 25931 3138 25987
rect 3194 25931 3219 25987
rect 3275 25931 3300 25987
rect 3356 25931 3381 25987
rect 3437 25931 3462 25987
rect 3518 25931 3543 25987
rect 3599 25931 3624 25987
rect 3680 25931 3705 25987
rect 3761 25931 3786 25987
rect 3842 25931 3867 25987
rect 3923 25931 3948 25987
rect 4004 25931 4029 25987
rect 4085 25931 4110 25987
rect 4166 25931 4191 25987
rect 4247 25931 4272 25987
rect 4328 25931 4353 25987
rect 4409 25931 4434 25987
rect 4490 25931 4515 25987
rect 4571 25931 4596 25987
rect 4652 25931 4677 25987
rect 4733 25931 4758 25987
rect 4814 25931 4839 25987
rect 4895 25931 4920 25987
rect 4976 25931 5001 25987
rect 5057 25931 5082 25987
rect 5138 25931 5163 25987
rect 2724 25907 5163 25931
rect 2724 25851 2733 25907
rect 2789 25851 2814 25907
rect 2870 25851 2895 25907
rect 2951 25851 2976 25907
rect 3032 25851 3057 25907
rect 3113 25851 3138 25907
rect 3194 25851 3219 25907
rect 3275 25851 3300 25907
rect 3356 25851 3381 25907
rect 3437 25851 3462 25907
rect 3518 25851 3543 25907
rect 3599 25851 3624 25907
rect 3680 25851 3705 25907
rect 3761 25851 3786 25907
rect 3842 25851 3867 25907
rect 3923 25851 3948 25907
rect 4004 25851 4029 25907
rect 4085 25851 4110 25907
rect 4166 25851 4191 25907
rect 4247 25851 4272 25907
rect 4328 25851 4353 25907
rect 4409 25851 4434 25907
rect 4490 25851 4515 25907
rect 4571 25851 4596 25907
rect 4652 25851 4677 25907
rect 4733 25851 4758 25907
rect 4814 25851 4839 25907
rect 4895 25851 4920 25907
rect 4976 25851 5001 25907
rect 5057 25851 5082 25907
rect 5138 25851 5163 25907
rect 2724 25827 5163 25851
rect 2724 25771 2733 25827
rect 2789 25771 2814 25827
rect 2870 25771 2895 25827
rect 2951 25771 2976 25827
rect 3032 25771 3057 25827
rect 3113 25771 3138 25827
rect 3194 25771 3219 25827
rect 3275 25771 3300 25827
rect 3356 25771 3381 25827
rect 3437 25771 3462 25827
rect 3518 25771 3543 25827
rect 3599 25771 3624 25827
rect 3680 25771 3705 25827
rect 3761 25771 3786 25827
rect 3842 25771 3867 25827
rect 3923 25771 3948 25827
rect 4004 25771 4029 25827
rect 4085 25771 4110 25827
rect 4166 25771 4191 25827
rect 4247 25771 4272 25827
rect 4328 25771 4353 25827
rect 4409 25771 4434 25827
rect 4490 25771 4515 25827
rect 4571 25771 4596 25827
rect 4652 25771 4677 25827
rect 4733 25771 4758 25827
rect 4814 25771 4839 25827
rect 4895 25771 4920 25827
rect 4976 25771 5001 25827
rect 5057 25771 5082 25827
rect 5138 25771 5163 25827
rect 2724 25747 5163 25771
rect 2724 25691 2733 25747
rect 2789 25691 2814 25747
rect 2870 25691 2895 25747
rect 2951 25691 2976 25747
rect 3032 25691 3057 25747
rect 3113 25691 3138 25747
rect 3194 25691 3219 25747
rect 3275 25691 3300 25747
rect 3356 25691 3381 25747
rect 3437 25691 3462 25747
rect 3518 25691 3543 25747
rect 3599 25691 3624 25747
rect 3680 25691 3705 25747
rect 3761 25691 3786 25747
rect 3842 25691 3867 25747
rect 3923 25691 3948 25747
rect 4004 25691 4029 25747
rect 4085 25691 4110 25747
rect 4166 25691 4191 25747
rect 4247 25691 4272 25747
rect 4328 25691 4353 25747
rect 4409 25691 4434 25747
rect 4490 25691 4515 25747
rect 4571 25691 4596 25747
rect 4652 25691 4677 25747
rect 4733 25691 4758 25747
rect 4814 25691 4839 25747
rect 4895 25691 4920 25747
rect 4976 25691 5001 25747
rect 5057 25691 5082 25747
rect 5138 25691 5163 25747
rect 2724 25667 5163 25691
rect 2724 25611 2733 25667
rect 2789 25611 2814 25667
rect 2870 25611 2895 25667
rect 2951 25611 2976 25667
rect 3032 25611 3057 25667
rect 3113 25611 3138 25667
rect 3194 25611 3219 25667
rect 3275 25611 3300 25667
rect 3356 25611 3381 25667
rect 3437 25611 3462 25667
rect 3518 25611 3543 25667
rect 3599 25611 3624 25667
rect 3680 25611 3705 25667
rect 3761 25611 3786 25667
rect 3842 25611 3867 25667
rect 3923 25611 3948 25667
rect 4004 25611 4029 25667
rect 4085 25611 4110 25667
rect 4166 25611 4191 25667
rect 4247 25611 4272 25667
rect 4328 25611 4353 25667
rect 4409 25611 4434 25667
rect 4490 25611 4515 25667
rect 4571 25611 4596 25667
rect 4652 25611 4677 25667
rect 4733 25611 4758 25667
rect 4814 25611 4839 25667
rect 4895 25611 4920 25667
rect 4976 25611 5001 25667
rect 5057 25611 5082 25667
rect 5138 25611 5163 25667
rect 2724 25587 5163 25611
rect 2724 25531 2733 25587
rect 2789 25531 2814 25587
rect 2870 25531 2895 25587
rect 2951 25531 2976 25587
rect 3032 25531 3057 25587
rect 3113 25531 3138 25587
rect 3194 25531 3219 25587
rect 3275 25531 3300 25587
rect 3356 25531 3381 25587
rect 3437 25531 3462 25587
rect 3518 25531 3543 25587
rect 3599 25531 3624 25587
rect 3680 25531 3705 25587
rect 3761 25531 3786 25587
rect 3842 25531 3867 25587
rect 3923 25531 3948 25587
rect 4004 25531 4029 25587
rect 4085 25531 4110 25587
rect 4166 25531 4191 25587
rect 4247 25531 4272 25587
rect 4328 25531 4353 25587
rect 4409 25531 4434 25587
rect 4490 25531 4515 25587
rect 4571 25531 4596 25587
rect 4652 25531 4677 25587
rect 4733 25531 4758 25587
rect 4814 25531 4839 25587
rect 4895 25531 4920 25587
rect 4976 25531 5001 25587
rect 5057 25531 5082 25587
rect 5138 25531 5163 25587
rect 2724 25507 5163 25531
rect 2724 25451 2733 25507
rect 2789 25451 2814 25507
rect 2870 25451 2895 25507
rect 2951 25451 2976 25507
rect 3032 25451 3057 25507
rect 3113 25451 3138 25507
rect 3194 25451 3219 25507
rect 3275 25451 3300 25507
rect 3356 25451 3381 25507
rect 3437 25451 3462 25507
rect 3518 25451 3543 25507
rect 3599 25451 3624 25507
rect 3680 25451 3705 25507
rect 3761 25451 3786 25507
rect 3842 25451 3867 25507
rect 3923 25451 3948 25507
rect 4004 25451 4029 25507
rect 4085 25451 4110 25507
rect 4166 25451 4191 25507
rect 4247 25451 4272 25507
rect 4328 25451 4353 25507
rect 4409 25451 4434 25507
rect 4490 25451 4515 25507
rect 4571 25451 4596 25507
rect 4652 25451 4677 25507
rect 4733 25451 4758 25507
rect 4814 25451 4839 25507
rect 4895 25451 4920 25507
rect 4976 25451 5001 25507
rect 5057 25451 5082 25507
rect 5138 25451 5163 25507
rect 2724 25427 5163 25451
rect 2724 25371 2733 25427
rect 2789 25371 2814 25427
rect 2870 25371 2895 25427
rect 2951 25371 2976 25427
rect 3032 25371 3057 25427
rect 3113 25371 3138 25427
rect 3194 25371 3219 25427
rect 3275 25371 3300 25427
rect 3356 25371 3381 25427
rect 3437 25371 3462 25427
rect 3518 25371 3543 25427
rect 3599 25371 3624 25427
rect 3680 25371 3705 25427
rect 3761 25371 3786 25427
rect 3842 25371 3867 25427
rect 3923 25371 3948 25427
rect 4004 25371 4029 25427
rect 4085 25371 4110 25427
rect 4166 25371 4191 25427
rect 4247 25371 4272 25427
rect 4328 25371 4353 25427
rect 4409 25371 4434 25427
rect 4490 25371 4515 25427
rect 4571 25371 4596 25427
rect 4652 25371 4677 25427
rect 4733 25371 4758 25427
rect 4814 25371 4839 25427
rect 4895 25371 4920 25427
rect 4976 25371 5001 25427
rect 5057 25371 5082 25427
rect 5138 25371 5163 25427
rect 5299 25982 7651 25987
rect 5299 25930 5317 25982
rect 5369 25930 5383 25982
rect 5435 25930 5871 25982
rect 5923 25930 5937 25982
rect 5989 25930 6425 25982
rect 6477 25930 6491 25982
rect 6543 25930 6979 25982
rect 7031 25930 7045 25982
rect 7097 25930 7533 25982
rect 7585 25930 7599 25982
rect 5299 25913 7651 25930
rect 5299 25861 5317 25913
rect 5369 25861 5383 25913
rect 5435 25861 5871 25913
rect 5923 25861 5937 25913
rect 5989 25861 6425 25913
rect 6477 25861 6491 25913
rect 6543 25861 6979 25913
rect 7031 25861 7045 25913
rect 7097 25861 7533 25913
rect 7585 25861 7599 25913
rect 5299 25844 7651 25861
rect 5299 25792 5317 25844
rect 5369 25792 5383 25844
rect 5435 25792 5871 25844
rect 5923 25792 5937 25844
rect 5989 25792 6425 25844
rect 6477 25792 6491 25844
rect 6543 25792 6979 25844
rect 7031 25792 7045 25844
rect 7097 25792 7533 25844
rect 7585 25792 7599 25844
rect 5299 25775 7651 25792
rect 5299 25723 5317 25775
rect 5369 25723 5383 25775
rect 5435 25723 5871 25775
rect 5923 25723 5937 25775
rect 5989 25723 6425 25775
rect 6477 25723 6491 25775
rect 6543 25723 6979 25775
rect 7031 25723 7045 25775
rect 7097 25723 7533 25775
rect 7585 25723 7599 25775
rect 5299 25706 7651 25723
rect 5299 25654 5317 25706
rect 5369 25654 5383 25706
rect 5435 25654 5871 25706
rect 5923 25654 5937 25706
rect 5989 25654 6425 25706
rect 6477 25654 6491 25706
rect 6543 25654 6979 25706
rect 7031 25654 7045 25706
rect 7097 25654 7533 25706
rect 7585 25654 7599 25706
rect 5299 25636 7651 25654
rect 5299 25584 5317 25636
rect 5369 25584 5383 25636
rect 5435 25584 5871 25636
rect 5923 25584 5937 25636
rect 5989 25584 6425 25636
rect 6477 25584 6491 25636
rect 6543 25584 6979 25636
rect 7031 25584 7045 25636
rect 7097 25584 7533 25636
rect 7585 25584 7599 25636
rect 5299 25566 7651 25584
rect 5299 25514 5317 25566
rect 5369 25514 5383 25566
rect 5435 25514 5871 25566
rect 5923 25514 5937 25566
rect 5989 25514 6425 25566
rect 6477 25514 6491 25566
rect 6543 25514 6979 25566
rect 7031 25514 7045 25566
rect 7097 25514 7533 25566
rect 7585 25514 7599 25566
rect 5299 25496 7651 25514
rect 5299 25444 5317 25496
rect 5369 25444 5383 25496
rect 5435 25444 5871 25496
rect 5923 25444 5937 25496
rect 5989 25444 6425 25496
rect 6477 25444 6491 25496
rect 6543 25444 6979 25496
rect 7031 25444 7045 25496
rect 7097 25444 7533 25496
rect 7585 25444 7599 25496
rect 5299 25426 7651 25444
rect 5299 25374 5317 25426
rect 5369 25374 5383 25426
rect 5435 25374 5871 25426
rect 5923 25374 5937 25426
rect 5989 25374 6425 25426
rect 6477 25374 6491 25426
rect 6543 25374 6979 25426
rect 7031 25374 7045 25426
rect 7097 25374 7533 25426
rect 7585 25374 7599 25426
rect 5299 25371 7651 25374
rect 2724 25368 7651 25371
rect 2270 24728 8222 24730
rect 2270 24724 2648 24728
rect 2322 24672 2392 24724
rect 2444 24676 2648 24724
rect 2700 24676 2713 24728
rect 2765 24676 2778 24728
rect 2830 24676 2843 24728
rect 2895 24676 2908 24728
rect 2960 24676 2973 24728
rect 3025 24676 3038 24728
rect 3090 24676 3103 24728
rect 3155 24676 3168 24728
rect 3220 24676 3233 24728
rect 3285 24676 3298 24728
rect 3350 24676 3363 24728
rect 3415 24676 3428 24728
rect 3480 24676 3493 24728
rect 3545 24676 3558 24728
rect 3610 24676 3623 24728
rect 3675 24676 3688 24728
rect 3740 24676 3753 24728
rect 3805 24676 3818 24728
rect 3870 24676 3883 24728
rect 3935 24676 3948 24728
rect 4000 24676 4013 24728
rect 4065 24676 4078 24728
rect 4130 24676 4143 24728
rect 4195 24676 4208 24728
rect 4260 24676 4273 24728
rect 4325 24676 4338 24728
rect 4390 24676 4403 24728
rect 4455 24676 4468 24728
rect 4520 24676 4532 24728
rect 4584 24724 8222 24728
rect 4584 24720 5613 24724
rect 5669 24720 5696 24724
rect 4584 24676 5040 24720
rect 2444 24672 5040 24676
rect 2270 24668 5040 24672
rect 5092 24668 5106 24720
rect 5158 24668 5594 24720
rect 5752 24668 5779 24724
rect 5835 24668 5861 24724
rect 5917 24668 5943 24724
rect 5999 24668 6025 24724
rect 6081 24668 6107 24724
rect 6163 24720 6189 24724
rect 6245 24720 6271 24724
rect 6266 24668 6271 24720
rect 6327 24668 6353 24724
rect 6409 24668 6435 24724
rect 6491 24668 6517 24724
rect 6573 24668 6599 24724
rect 6655 24668 6681 24724
rect 6737 24720 6763 24724
rect 6819 24720 6845 24724
rect 6754 24668 6763 24720
rect 6820 24668 6845 24720
rect 6901 24668 6927 24724
rect 6983 24668 7009 24724
rect 7065 24668 7091 24724
rect 7147 24668 7173 24724
rect 7229 24668 7255 24724
rect 7311 24720 7337 24724
rect 7311 24668 7322 24720
rect 7393 24668 7419 24724
rect 7475 24668 7501 24724
rect 7557 24668 7583 24724
rect 7639 24668 7665 24724
rect 7721 24668 7747 24724
rect 7803 24720 7829 24724
rect 7885 24720 7911 24724
rect 7803 24668 7810 24720
rect 7967 24668 7993 24724
rect 8049 24668 8075 24672
rect 8131 24668 8157 24724
rect 8221 24672 8222 24724
rect 8213 24668 8222 24672
rect 2270 24660 8222 24668
rect 2270 24655 2648 24660
rect 2322 24603 2392 24655
rect 2444 24608 2648 24655
rect 2700 24608 2713 24660
rect 2765 24608 2778 24660
rect 2830 24608 2843 24660
rect 2895 24608 2908 24660
rect 2960 24608 2973 24660
rect 3025 24608 3038 24660
rect 3090 24608 3103 24660
rect 3155 24608 3168 24660
rect 3220 24608 3233 24660
rect 3285 24608 3298 24660
rect 3350 24608 3363 24660
rect 3415 24608 3428 24660
rect 3480 24608 3493 24660
rect 3545 24608 3558 24660
rect 3610 24608 3623 24660
rect 3675 24608 3688 24660
rect 3740 24608 3753 24660
rect 3805 24608 3818 24660
rect 3870 24608 3883 24660
rect 3935 24608 3948 24660
rect 4000 24608 4013 24660
rect 4065 24608 4078 24660
rect 4130 24608 4143 24660
rect 4195 24608 4208 24660
rect 4260 24608 4273 24660
rect 4325 24608 4338 24660
rect 4390 24608 4403 24660
rect 4455 24608 4468 24660
rect 4520 24608 4532 24660
rect 4584 24655 8222 24660
rect 4584 24651 8047 24655
rect 4584 24608 5040 24651
rect 2444 24603 5040 24608
rect 2270 24599 5040 24603
rect 5092 24599 5106 24651
rect 5158 24599 5594 24651
rect 5646 24644 5660 24651
rect 5712 24644 6148 24651
rect 6200 24644 6214 24651
rect 6266 24644 6702 24651
rect 6754 24644 6768 24651
rect 6820 24644 7256 24651
rect 7308 24644 7322 24651
rect 7374 24644 7810 24651
rect 7862 24644 7876 24651
rect 7928 24644 8047 24651
rect 8099 24644 8169 24655
rect 2270 24592 5613 24599
rect 2270 24586 2648 24592
rect 2322 24534 2392 24586
rect 2444 24540 2648 24586
rect 2700 24540 2713 24592
rect 2765 24540 2778 24592
rect 2830 24540 2843 24592
rect 2895 24540 2908 24592
rect 2960 24540 2973 24592
rect 3025 24540 3038 24592
rect 3090 24540 3103 24592
rect 3155 24540 3168 24592
rect 3220 24540 3233 24592
rect 3285 24540 3298 24592
rect 3350 24540 3363 24592
rect 3415 24540 3428 24592
rect 3480 24540 3493 24592
rect 3545 24540 3558 24592
rect 3610 24540 3623 24592
rect 3675 24540 3688 24592
rect 3740 24540 3753 24592
rect 3805 24540 3818 24592
rect 3870 24540 3883 24592
rect 3935 24540 3948 24592
rect 4000 24540 4013 24592
rect 4065 24540 4078 24592
rect 4130 24540 4143 24592
rect 4195 24540 4208 24592
rect 4260 24540 4273 24592
rect 4325 24540 4338 24592
rect 4390 24540 4403 24592
rect 4455 24540 4468 24592
rect 4520 24540 4532 24592
rect 4584 24588 5613 24592
rect 5669 24588 5696 24599
rect 5752 24588 5779 24644
rect 5835 24588 5861 24644
rect 5917 24588 5943 24644
rect 5999 24588 6025 24644
rect 6081 24588 6107 24644
rect 6266 24599 6271 24644
rect 6163 24588 6189 24599
rect 6245 24588 6271 24599
rect 6327 24588 6353 24644
rect 6409 24588 6435 24644
rect 6491 24588 6517 24644
rect 6573 24588 6599 24644
rect 6655 24588 6681 24644
rect 6754 24599 6763 24644
rect 6820 24599 6845 24644
rect 6737 24588 6763 24599
rect 6819 24588 6845 24599
rect 6901 24588 6927 24644
rect 6983 24588 7009 24644
rect 7065 24588 7091 24644
rect 7147 24588 7173 24644
rect 7229 24588 7255 24644
rect 7311 24599 7322 24644
rect 7311 24588 7337 24599
rect 7393 24588 7419 24644
rect 7475 24588 7501 24644
rect 7557 24588 7583 24644
rect 7639 24588 7665 24644
rect 7721 24588 7747 24644
rect 7803 24599 7810 24644
rect 7803 24588 7829 24599
rect 7885 24588 7911 24599
rect 7967 24588 7993 24644
rect 8049 24588 8075 24603
rect 8131 24588 8157 24644
rect 8221 24603 8222 24655
rect 8213 24588 8222 24603
rect 4584 24586 8222 24588
rect 4584 24582 8047 24586
rect 4584 24540 5040 24582
rect 2444 24534 5040 24540
rect 2270 24530 5040 24534
rect 5092 24530 5106 24582
rect 5158 24530 5594 24582
rect 5646 24564 5660 24582
rect 5712 24564 6148 24582
rect 6200 24564 6214 24582
rect 6266 24564 6702 24582
rect 6754 24564 6768 24582
rect 6820 24564 7256 24582
rect 7308 24564 7322 24582
rect 7374 24564 7810 24582
rect 7862 24564 7876 24582
rect 7928 24564 8047 24582
rect 8099 24564 8169 24586
rect 2270 24524 5613 24530
rect 2270 24517 2648 24524
rect 2322 24465 2392 24517
rect 2444 24472 2648 24517
rect 2700 24472 2713 24524
rect 2765 24472 2778 24524
rect 2830 24472 2843 24524
rect 2895 24472 2908 24524
rect 2960 24472 2973 24524
rect 3025 24472 3038 24524
rect 3090 24472 3103 24524
rect 3155 24472 3168 24524
rect 3220 24472 3233 24524
rect 3285 24472 3298 24524
rect 3350 24472 3363 24524
rect 3415 24472 3428 24524
rect 3480 24472 3493 24524
rect 3545 24472 3558 24524
rect 3610 24472 3623 24524
rect 3675 24472 3688 24524
rect 3740 24472 3753 24524
rect 3805 24472 3818 24524
rect 3870 24472 3883 24524
rect 3935 24472 3948 24524
rect 4000 24472 4013 24524
rect 4065 24472 4078 24524
rect 4130 24472 4143 24524
rect 4195 24472 4208 24524
rect 4260 24472 4273 24524
rect 4325 24472 4338 24524
rect 4390 24472 4403 24524
rect 4455 24472 4468 24524
rect 4520 24472 4532 24524
rect 4584 24513 5613 24524
rect 5669 24513 5696 24530
rect 4584 24472 5040 24513
rect 2444 24465 5040 24472
rect 2270 24461 5040 24465
rect 5092 24461 5106 24513
rect 5158 24461 5594 24513
rect 5752 24508 5779 24564
rect 5835 24508 5861 24564
rect 5917 24508 5943 24564
rect 5999 24508 6025 24564
rect 6081 24508 6107 24564
rect 6266 24530 6271 24564
rect 6163 24513 6189 24530
rect 6245 24513 6271 24530
rect 6266 24508 6271 24513
rect 6327 24508 6353 24564
rect 6409 24508 6435 24564
rect 6491 24508 6517 24564
rect 6573 24508 6599 24564
rect 6655 24508 6681 24564
rect 6754 24530 6763 24564
rect 6820 24530 6845 24564
rect 6737 24513 6763 24530
rect 6819 24513 6845 24530
rect 6754 24508 6763 24513
rect 6820 24508 6845 24513
rect 6901 24508 6927 24564
rect 6983 24508 7009 24564
rect 7065 24508 7091 24564
rect 7147 24508 7173 24564
rect 7229 24508 7255 24564
rect 7311 24530 7322 24564
rect 7311 24513 7337 24530
rect 7311 24508 7322 24513
rect 7393 24508 7419 24564
rect 7475 24508 7501 24564
rect 7557 24508 7583 24564
rect 7639 24508 7665 24564
rect 7721 24508 7747 24564
rect 7803 24530 7810 24564
rect 7803 24513 7829 24530
rect 7885 24513 7911 24530
rect 7803 24508 7810 24513
rect 7967 24508 7993 24564
rect 8049 24517 8075 24534
rect 8131 24508 8157 24564
rect 8221 24534 8222 24586
rect 8213 24517 8222 24534
rect 5646 24484 5660 24508
rect 5712 24484 6148 24508
rect 6200 24484 6214 24508
rect 6266 24484 6702 24508
rect 6754 24484 6768 24508
rect 6820 24484 7256 24508
rect 7308 24484 7322 24508
rect 7374 24484 7810 24508
rect 7862 24484 7876 24508
rect 7928 24484 8047 24508
rect 8099 24484 8169 24508
rect 2270 24456 5613 24461
rect 2270 24448 2648 24456
rect 2322 24396 2392 24448
rect 2444 24404 2648 24448
rect 2700 24404 2713 24456
rect 2765 24404 2778 24456
rect 2830 24404 2843 24456
rect 2895 24404 2908 24456
rect 2960 24404 2973 24456
rect 3025 24404 3038 24456
rect 3090 24404 3103 24456
rect 3155 24404 3168 24456
rect 3220 24404 3233 24456
rect 3285 24404 3298 24456
rect 3350 24404 3363 24456
rect 3415 24404 3428 24456
rect 3480 24404 3493 24456
rect 3545 24404 3558 24456
rect 3610 24404 3623 24456
rect 3675 24404 3688 24456
rect 3740 24404 3753 24456
rect 3805 24404 3818 24456
rect 3870 24404 3883 24456
rect 3935 24404 3948 24456
rect 4000 24404 4013 24456
rect 4065 24404 4078 24456
rect 4130 24404 4143 24456
rect 4195 24404 4208 24456
rect 4260 24404 4273 24456
rect 4325 24404 4338 24456
rect 4390 24404 4403 24456
rect 4455 24404 4468 24456
rect 4520 24404 4532 24456
rect 4584 24444 5613 24456
rect 5669 24444 5696 24461
rect 4584 24404 5040 24444
rect 2444 24396 5040 24404
rect 2270 24392 5040 24396
rect 5092 24392 5106 24444
rect 5158 24392 5594 24444
rect 5752 24428 5779 24484
rect 5835 24428 5861 24484
rect 5917 24428 5943 24484
rect 5999 24428 6025 24484
rect 6081 24428 6107 24484
rect 6266 24461 6271 24484
rect 6163 24444 6189 24461
rect 6245 24444 6271 24461
rect 6266 24428 6271 24444
rect 6327 24428 6353 24484
rect 6409 24428 6435 24484
rect 6491 24428 6517 24484
rect 6573 24428 6599 24484
rect 6655 24428 6681 24484
rect 6754 24461 6763 24484
rect 6820 24461 6845 24484
rect 6737 24444 6763 24461
rect 6819 24444 6845 24461
rect 6754 24428 6763 24444
rect 6820 24428 6845 24444
rect 6901 24428 6927 24484
rect 6983 24428 7009 24484
rect 7065 24428 7091 24484
rect 7147 24428 7173 24484
rect 7229 24428 7255 24484
rect 7311 24461 7322 24484
rect 7311 24444 7337 24461
rect 7311 24428 7322 24444
rect 7393 24428 7419 24484
rect 7475 24428 7501 24484
rect 7557 24428 7583 24484
rect 7639 24428 7665 24484
rect 7721 24428 7747 24484
rect 7803 24461 7810 24484
rect 7803 24444 7829 24461
rect 7885 24444 7911 24461
rect 7803 24428 7810 24444
rect 7967 24428 7993 24484
rect 8049 24448 8075 24465
rect 8131 24428 8157 24484
rect 8221 24465 8222 24517
rect 8213 24448 8222 24465
rect 5646 24404 5660 24428
rect 5712 24404 6148 24428
rect 6200 24404 6214 24428
rect 6266 24404 6702 24428
rect 6754 24404 6768 24428
rect 6820 24404 7256 24428
rect 7308 24404 7322 24428
rect 7374 24404 7810 24428
rect 7862 24404 7876 24428
rect 7928 24404 8047 24428
rect 8099 24404 8169 24428
rect 2270 24388 5613 24392
rect 2270 24378 2648 24388
rect 2322 24326 2392 24378
rect 2444 24336 2648 24378
rect 2700 24336 2713 24388
rect 2765 24336 2778 24388
rect 2830 24336 2843 24388
rect 2895 24336 2908 24388
rect 2960 24336 2973 24388
rect 3025 24336 3038 24388
rect 3090 24336 3103 24388
rect 3155 24336 3168 24388
rect 3220 24336 3233 24388
rect 3285 24336 3298 24388
rect 3350 24336 3363 24388
rect 3415 24336 3428 24388
rect 3480 24336 3493 24388
rect 3545 24336 3558 24388
rect 3610 24336 3623 24388
rect 3675 24336 3688 24388
rect 3740 24336 3753 24388
rect 3805 24336 3818 24388
rect 3870 24336 3883 24388
rect 3935 24336 3948 24388
rect 4000 24336 4013 24388
rect 4065 24336 4078 24388
rect 4130 24336 4143 24388
rect 4195 24336 4208 24388
rect 4260 24336 4273 24388
rect 4325 24336 4338 24388
rect 4390 24336 4403 24388
rect 4455 24336 4468 24388
rect 4520 24336 4532 24388
rect 4584 24375 5613 24388
rect 5669 24375 5696 24392
rect 4584 24336 5040 24375
rect 2444 24326 5040 24336
rect 2270 24323 5040 24326
rect 5092 24323 5106 24375
rect 5158 24323 5594 24375
rect 5752 24348 5779 24404
rect 5835 24348 5861 24404
rect 5917 24348 5943 24404
rect 5999 24348 6025 24404
rect 6081 24348 6107 24404
rect 6266 24392 6271 24404
rect 6163 24375 6189 24392
rect 6245 24375 6271 24392
rect 6266 24348 6271 24375
rect 6327 24348 6353 24404
rect 6409 24348 6435 24404
rect 6491 24348 6517 24404
rect 6573 24348 6599 24404
rect 6655 24348 6681 24404
rect 6754 24392 6763 24404
rect 6820 24392 6845 24404
rect 6737 24375 6763 24392
rect 6819 24375 6845 24392
rect 6754 24348 6763 24375
rect 6820 24348 6845 24375
rect 6901 24348 6927 24404
rect 6983 24348 7009 24404
rect 7065 24348 7091 24404
rect 7147 24348 7173 24404
rect 7229 24348 7255 24404
rect 7311 24392 7322 24404
rect 7311 24375 7337 24392
rect 7311 24348 7322 24375
rect 7393 24348 7419 24404
rect 7475 24348 7501 24404
rect 7557 24348 7583 24404
rect 7639 24348 7665 24404
rect 7721 24348 7747 24404
rect 7803 24392 7810 24404
rect 7803 24375 7829 24392
rect 7885 24375 7911 24392
rect 7803 24348 7810 24375
rect 7967 24348 7993 24404
rect 8049 24378 8075 24396
rect 8131 24348 8157 24404
rect 8221 24396 8222 24448
rect 8213 24378 8222 24396
rect 5646 24324 5660 24348
rect 5712 24324 6148 24348
rect 6200 24324 6214 24348
rect 6266 24324 6702 24348
rect 6754 24324 6768 24348
rect 6820 24324 7256 24348
rect 7308 24324 7322 24348
rect 7374 24324 7810 24348
rect 7862 24324 7876 24348
rect 7928 24326 8047 24348
rect 8099 24326 8169 24348
rect 8221 24326 8222 24378
rect 7928 24324 8222 24326
rect 2270 24320 5613 24323
rect 2270 24308 2648 24320
rect 2322 24256 2392 24308
rect 2444 24268 2648 24308
rect 2700 24268 2713 24320
rect 2765 24268 2778 24320
rect 2830 24268 2843 24320
rect 2895 24268 2908 24320
rect 2960 24268 2973 24320
rect 3025 24268 3038 24320
rect 3090 24268 3103 24320
rect 3155 24268 3168 24320
rect 3220 24268 3233 24320
rect 3285 24268 3298 24320
rect 3350 24268 3363 24320
rect 3415 24268 3428 24320
rect 3480 24268 3493 24320
rect 3545 24268 3558 24320
rect 3610 24268 3623 24320
rect 3675 24268 3688 24320
rect 3740 24268 3753 24320
rect 3805 24268 3818 24320
rect 3870 24268 3883 24320
rect 3935 24268 3948 24320
rect 4000 24268 4013 24320
rect 4065 24268 4078 24320
rect 4130 24268 4143 24320
rect 4195 24268 4208 24320
rect 4260 24268 4273 24320
rect 4325 24268 4338 24320
rect 4390 24268 4403 24320
rect 4455 24268 4468 24320
rect 4520 24268 4532 24320
rect 4584 24306 5613 24320
rect 5669 24306 5696 24323
rect 4584 24268 5040 24306
rect 2444 24256 5040 24268
rect 2270 24254 5040 24256
rect 5092 24254 5106 24306
rect 5158 24254 5594 24306
rect 5752 24268 5779 24324
rect 5835 24268 5861 24324
rect 5917 24268 5943 24324
rect 5999 24268 6025 24324
rect 6081 24268 6107 24324
rect 6266 24323 6271 24324
rect 6163 24306 6189 24323
rect 6245 24306 6271 24323
rect 6266 24268 6271 24306
rect 6327 24268 6353 24324
rect 6409 24268 6435 24324
rect 6491 24268 6517 24324
rect 6573 24268 6599 24324
rect 6655 24268 6681 24324
rect 6754 24323 6763 24324
rect 6820 24323 6845 24324
rect 6737 24306 6763 24323
rect 6819 24306 6845 24323
rect 6754 24268 6763 24306
rect 6820 24268 6845 24306
rect 6901 24268 6927 24324
rect 6983 24268 7009 24324
rect 7065 24268 7091 24324
rect 7147 24268 7173 24324
rect 7229 24268 7255 24324
rect 7311 24323 7322 24324
rect 7311 24306 7337 24323
rect 7311 24268 7322 24306
rect 7393 24268 7419 24324
rect 7475 24268 7501 24324
rect 7557 24268 7583 24324
rect 7639 24268 7665 24324
rect 7721 24268 7747 24324
rect 7803 24323 7810 24324
rect 7803 24306 7829 24323
rect 7885 24306 7911 24323
rect 7803 24268 7810 24306
rect 7967 24268 7993 24324
rect 8049 24308 8075 24324
rect 8131 24268 8157 24324
rect 8213 24308 8222 24324
rect 5646 24254 5660 24268
rect 5712 24254 6148 24268
rect 6200 24254 6214 24268
rect 6266 24254 6702 24268
rect 6754 24254 6768 24268
rect 6820 24254 7256 24268
rect 7308 24254 7322 24268
rect 7374 24254 7810 24268
rect 7862 24254 7876 24268
rect 7928 24256 8047 24268
rect 8099 24256 8169 24268
rect 8221 24256 8222 24308
rect 7928 24254 8222 24256
rect 2270 24252 8222 24254
rect 2270 24238 2648 24252
rect 2322 24186 2392 24238
rect 2444 24200 2648 24238
rect 2700 24200 2713 24252
rect 2765 24200 2778 24252
rect 2830 24200 2843 24252
rect 2895 24200 2908 24252
rect 2960 24200 2973 24252
rect 3025 24200 3038 24252
rect 3090 24200 3103 24252
rect 3155 24200 3168 24252
rect 3220 24200 3233 24252
rect 3285 24200 3298 24252
rect 3350 24200 3363 24252
rect 3415 24200 3428 24252
rect 3480 24200 3493 24252
rect 3545 24200 3558 24252
rect 3610 24200 3623 24252
rect 3675 24200 3688 24252
rect 3740 24200 3753 24252
rect 3805 24200 3818 24252
rect 3870 24200 3883 24252
rect 3935 24200 3948 24252
rect 4000 24200 4013 24252
rect 4065 24200 4078 24252
rect 4130 24200 4143 24252
rect 4195 24200 4208 24252
rect 4260 24200 4273 24252
rect 4325 24200 4338 24252
rect 4390 24200 4403 24252
rect 4455 24200 4468 24252
rect 4520 24200 4532 24252
rect 4584 24244 8222 24252
rect 4584 24236 5613 24244
rect 5669 24236 5696 24244
rect 4584 24200 5040 24236
rect 2444 24186 5040 24200
rect 2270 24184 5040 24186
rect 5092 24184 5106 24236
rect 5158 24184 5594 24236
rect 5752 24188 5779 24244
rect 5835 24188 5861 24244
rect 5917 24188 5943 24244
rect 5999 24188 6025 24244
rect 6081 24188 6107 24244
rect 6163 24236 6189 24244
rect 6245 24236 6271 24244
rect 6266 24188 6271 24236
rect 6327 24188 6353 24244
rect 6409 24188 6435 24244
rect 6491 24188 6517 24244
rect 6573 24188 6599 24244
rect 6655 24188 6681 24244
rect 6737 24236 6763 24244
rect 6819 24236 6845 24244
rect 6754 24188 6763 24236
rect 6820 24188 6845 24236
rect 6901 24188 6927 24244
rect 6983 24188 7009 24244
rect 7065 24188 7091 24244
rect 7147 24188 7173 24244
rect 7229 24188 7255 24244
rect 7311 24236 7337 24244
rect 7311 24188 7322 24236
rect 7393 24188 7419 24244
rect 7475 24188 7501 24244
rect 7557 24188 7583 24244
rect 7639 24188 7665 24244
rect 7721 24188 7747 24244
rect 7803 24236 7829 24244
rect 7885 24236 7911 24244
rect 7803 24188 7810 24236
rect 7967 24188 7993 24244
rect 8049 24238 8075 24244
rect 8131 24188 8157 24244
rect 8213 24238 8222 24244
rect 5646 24184 5660 24188
rect 5712 24184 6148 24188
rect 6200 24184 6214 24188
rect 6266 24184 6702 24188
rect 6754 24184 6768 24188
rect 6820 24184 7256 24188
rect 7308 24184 7322 24188
rect 7374 24184 7810 24188
rect 7862 24184 7876 24188
rect 7928 24186 8047 24188
rect 8099 24186 8169 24188
rect 8221 24186 8222 24238
rect 7928 24184 8222 24186
rect 2270 24168 8222 24184
rect 2322 24116 2392 24168
rect 2444 24166 8047 24168
rect 2444 24116 5040 24166
rect 2270 24114 5040 24116
rect 5092 24114 5106 24166
rect 5158 24114 5594 24166
rect 5646 24164 5660 24166
rect 5712 24164 6148 24166
rect 6200 24164 6214 24166
rect 6266 24164 6702 24166
rect 6754 24164 6768 24166
rect 6820 24164 7256 24166
rect 7308 24164 7322 24166
rect 7374 24164 7810 24166
rect 7862 24164 7876 24166
rect 7928 24164 8047 24166
rect 8099 24164 8169 24168
rect 2270 24108 5613 24114
rect 5669 24108 5696 24114
rect 5752 24108 5779 24164
rect 5835 24108 5861 24164
rect 5917 24108 5943 24164
rect 5999 24108 6025 24164
rect 6081 24108 6107 24164
rect 6266 24114 6271 24164
rect 6163 24108 6189 24114
rect 6245 24108 6271 24114
rect 6327 24108 6353 24164
rect 6409 24108 6435 24164
rect 6491 24108 6517 24164
rect 6573 24108 6599 24164
rect 6655 24108 6681 24164
rect 6754 24114 6763 24164
rect 6820 24114 6845 24164
rect 6737 24108 6763 24114
rect 6819 24108 6845 24114
rect 6901 24108 6927 24164
rect 6983 24108 7009 24164
rect 7065 24108 7091 24164
rect 7147 24108 7173 24164
rect 7229 24108 7255 24164
rect 7311 24114 7322 24164
rect 7311 24108 7337 24114
rect 7393 24108 7419 24164
rect 7475 24108 7501 24164
rect 7557 24108 7583 24164
rect 7639 24108 7665 24164
rect 7721 24108 7747 24164
rect 7803 24114 7810 24164
rect 7803 24108 7829 24114
rect 7885 24108 7911 24114
rect 7967 24108 7993 24164
rect 8049 24108 8075 24116
rect 8131 24108 8157 24164
rect 8221 24116 8222 24168
rect 8213 24108 8222 24116
rect 2724 23987 7651 23988
rect 2724 23931 2733 23987
rect 2789 23931 2814 23987
rect 2870 23931 2895 23987
rect 2951 23931 2976 23987
rect 3032 23931 3057 23987
rect 3113 23931 3138 23987
rect 3194 23931 3219 23987
rect 3275 23931 3300 23987
rect 3356 23931 3381 23987
rect 3437 23931 3462 23987
rect 3518 23931 3543 23987
rect 3599 23931 3624 23987
rect 3680 23931 3705 23987
rect 3761 23931 3786 23987
rect 3842 23931 3867 23987
rect 3923 23931 3948 23987
rect 4004 23931 4029 23987
rect 4085 23931 4110 23987
rect 4166 23931 4191 23987
rect 4247 23931 4272 23987
rect 4328 23931 4353 23987
rect 4409 23931 4434 23987
rect 4490 23931 4515 23987
rect 4571 23931 4596 23987
rect 4652 23931 4677 23987
rect 4733 23931 4758 23987
rect 4814 23931 4839 23987
rect 4895 23931 4920 23987
rect 4976 23931 5001 23987
rect 5057 23931 5082 23987
rect 5138 23931 5163 23987
rect 2724 23907 5163 23931
rect 2724 23851 2733 23907
rect 2789 23851 2814 23907
rect 2870 23851 2895 23907
rect 2951 23851 2976 23907
rect 3032 23851 3057 23907
rect 3113 23851 3138 23907
rect 3194 23851 3219 23907
rect 3275 23851 3300 23907
rect 3356 23851 3381 23907
rect 3437 23851 3462 23907
rect 3518 23851 3543 23907
rect 3599 23851 3624 23907
rect 3680 23851 3705 23907
rect 3761 23851 3786 23907
rect 3842 23851 3867 23907
rect 3923 23851 3948 23907
rect 4004 23851 4029 23907
rect 4085 23851 4110 23907
rect 4166 23851 4191 23907
rect 4247 23851 4272 23907
rect 4328 23851 4353 23907
rect 4409 23851 4434 23907
rect 4490 23851 4515 23907
rect 4571 23851 4596 23907
rect 4652 23851 4677 23907
rect 4733 23851 4758 23907
rect 4814 23851 4839 23907
rect 4895 23851 4920 23907
rect 4976 23851 5001 23907
rect 5057 23851 5082 23907
rect 5138 23851 5163 23907
rect 2724 23827 5163 23851
rect 2724 23771 2733 23827
rect 2789 23771 2814 23827
rect 2870 23771 2895 23827
rect 2951 23771 2976 23827
rect 3032 23771 3057 23827
rect 3113 23771 3138 23827
rect 3194 23771 3219 23827
rect 3275 23771 3300 23827
rect 3356 23771 3381 23827
rect 3437 23771 3462 23827
rect 3518 23771 3543 23827
rect 3599 23771 3624 23827
rect 3680 23771 3705 23827
rect 3761 23771 3786 23827
rect 3842 23771 3867 23827
rect 3923 23771 3948 23827
rect 4004 23771 4029 23827
rect 4085 23771 4110 23827
rect 4166 23771 4191 23827
rect 4247 23771 4272 23827
rect 4328 23771 4353 23827
rect 4409 23771 4434 23827
rect 4490 23771 4515 23827
rect 4571 23771 4596 23827
rect 4652 23771 4677 23827
rect 4733 23771 4758 23827
rect 4814 23771 4839 23827
rect 4895 23771 4920 23827
rect 4976 23771 5001 23827
rect 5057 23771 5082 23827
rect 5138 23771 5163 23827
rect 2724 23747 5163 23771
rect 2724 23691 2733 23747
rect 2789 23691 2814 23747
rect 2870 23691 2895 23747
rect 2951 23691 2976 23747
rect 3032 23691 3057 23747
rect 3113 23691 3138 23747
rect 3194 23691 3219 23747
rect 3275 23691 3300 23747
rect 3356 23691 3381 23747
rect 3437 23691 3462 23747
rect 3518 23691 3543 23747
rect 3599 23691 3624 23747
rect 3680 23691 3705 23747
rect 3761 23691 3786 23747
rect 3842 23691 3867 23747
rect 3923 23691 3948 23747
rect 4004 23691 4029 23747
rect 4085 23691 4110 23747
rect 4166 23691 4191 23747
rect 4247 23691 4272 23747
rect 4328 23691 4353 23747
rect 4409 23691 4434 23747
rect 4490 23691 4515 23747
rect 4571 23691 4596 23747
rect 4652 23691 4677 23747
rect 4733 23691 4758 23747
rect 4814 23691 4839 23747
rect 4895 23691 4920 23747
rect 4976 23691 5001 23747
rect 5057 23691 5082 23747
rect 5138 23691 5163 23747
rect 2724 23667 5163 23691
rect 2724 23611 2733 23667
rect 2789 23611 2814 23667
rect 2870 23611 2895 23667
rect 2951 23611 2976 23667
rect 3032 23611 3057 23667
rect 3113 23611 3138 23667
rect 3194 23611 3219 23667
rect 3275 23611 3300 23667
rect 3356 23611 3381 23667
rect 3437 23611 3462 23667
rect 3518 23611 3543 23667
rect 3599 23611 3624 23667
rect 3680 23611 3705 23667
rect 3761 23611 3786 23667
rect 3842 23611 3867 23667
rect 3923 23611 3948 23667
rect 4004 23611 4029 23667
rect 4085 23611 4110 23667
rect 4166 23611 4191 23667
rect 4247 23611 4272 23667
rect 4328 23611 4353 23667
rect 4409 23611 4434 23667
rect 4490 23611 4515 23667
rect 4571 23611 4596 23667
rect 4652 23611 4677 23667
rect 4733 23611 4758 23667
rect 4814 23611 4839 23667
rect 4895 23611 4920 23667
rect 4976 23611 5001 23667
rect 5057 23611 5082 23667
rect 5138 23611 5163 23667
rect 2724 23587 5163 23611
rect 2724 23531 2733 23587
rect 2789 23531 2814 23587
rect 2870 23531 2895 23587
rect 2951 23531 2976 23587
rect 3032 23531 3057 23587
rect 3113 23531 3138 23587
rect 3194 23531 3219 23587
rect 3275 23531 3300 23587
rect 3356 23531 3381 23587
rect 3437 23531 3462 23587
rect 3518 23531 3543 23587
rect 3599 23531 3624 23587
rect 3680 23531 3705 23587
rect 3761 23531 3786 23587
rect 3842 23531 3867 23587
rect 3923 23531 3948 23587
rect 4004 23531 4029 23587
rect 4085 23531 4110 23587
rect 4166 23531 4191 23587
rect 4247 23531 4272 23587
rect 4328 23531 4353 23587
rect 4409 23531 4434 23587
rect 4490 23531 4515 23587
rect 4571 23531 4596 23587
rect 4652 23531 4677 23587
rect 4733 23531 4758 23587
rect 4814 23531 4839 23587
rect 4895 23531 4920 23587
rect 4976 23531 5001 23587
rect 5057 23531 5082 23587
rect 5138 23531 5163 23587
rect 2724 23507 5163 23531
rect 2724 23451 2733 23507
rect 2789 23451 2814 23507
rect 2870 23451 2895 23507
rect 2951 23451 2976 23507
rect 3032 23451 3057 23507
rect 3113 23451 3138 23507
rect 3194 23451 3219 23507
rect 3275 23451 3300 23507
rect 3356 23451 3381 23507
rect 3437 23451 3462 23507
rect 3518 23451 3543 23507
rect 3599 23451 3624 23507
rect 3680 23451 3705 23507
rect 3761 23451 3786 23507
rect 3842 23451 3867 23507
rect 3923 23451 3948 23507
rect 4004 23451 4029 23507
rect 4085 23451 4110 23507
rect 4166 23451 4191 23507
rect 4247 23451 4272 23507
rect 4328 23451 4353 23507
rect 4409 23451 4434 23507
rect 4490 23451 4515 23507
rect 4571 23451 4596 23507
rect 4652 23451 4677 23507
rect 4733 23451 4758 23507
rect 4814 23451 4839 23507
rect 4895 23451 4920 23507
rect 4976 23451 5001 23507
rect 5057 23451 5082 23507
rect 5138 23451 5163 23507
rect 2724 23427 5163 23451
rect 2724 23371 2733 23427
rect 2789 23371 2814 23427
rect 2870 23371 2895 23427
rect 2951 23371 2976 23427
rect 3032 23371 3057 23427
rect 3113 23371 3138 23427
rect 3194 23371 3219 23427
rect 3275 23371 3300 23427
rect 3356 23371 3381 23427
rect 3437 23371 3462 23427
rect 3518 23371 3543 23427
rect 3599 23371 3624 23427
rect 3680 23371 3705 23427
rect 3761 23371 3786 23427
rect 3842 23371 3867 23427
rect 3923 23371 3948 23427
rect 4004 23371 4029 23427
rect 4085 23371 4110 23427
rect 4166 23371 4191 23427
rect 4247 23371 4272 23427
rect 4328 23371 4353 23427
rect 4409 23371 4434 23427
rect 4490 23371 4515 23427
rect 4571 23371 4596 23427
rect 4652 23371 4677 23427
rect 4733 23371 4758 23427
rect 4814 23371 4839 23427
rect 4895 23371 4920 23427
rect 4976 23371 5001 23427
rect 5057 23371 5082 23427
rect 5138 23371 5163 23427
rect 5299 23982 7651 23987
rect 5299 23930 5317 23982
rect 5369 23930 5383 23982
rect 5435 23930 5871 23982
rect 5923 23930 5937 23982
rect 5989 23930 6425 23982
rect 6477 23930 6491 23982
rect 6543 23930 6979 23982
rect 7031 23930 7045 23982
rect 7097 23930 7533 23982
rect 7585 23930 7599 23982
rect 5299 23913 7651 23930
rect 5299 23861 5317 23913
rect 5369 23861 5383 23913
rect 5435 23861 5871 23913
rect 5923 23861 5937 23913
rect 5989 23861 6425 23913
rect 6477 23861 6491 23913
rect 6543 23861 6979 23913
rect 7031 23861 7045 23913
rect 7097 23861 7533 23913
rect 7585 23861 7599 23913
rect 5299 23844 7651 23861
rect 5299 23792 5317 23844
rect 5369 23792 5383 23844
rect 5435 23792 5871 23844
rect 5923 23792 5937 23844
rect 5989 23792 6425 23844
rect 6477 23792 6491 23844
rect 6543 23792 6979 23844
rect 7031 23792 7045 23844
rect 7097 23792 7533 23844
rect 7585 23792 7599 23844
rect 5299 23775 7651 23792
rect 5299 23723 5317 23775
rect 5369 23723 5383 23775
rect 5435 23723 5871 23775
rect 5923 23723 5937 23775
rect 5989 23723 6425 23775
rect 6477 23723 6491 23775
rect 6543 23723 6979 23775
rect 7031 23723 7045 23775
rect 7097 23723 7533 23775
rect 7585 23723 7599 23775
rect 5299 23706 7651 23723
rect 5299 23654 5317 23706
rect 5369 23654 5383 23706
rect 5435 23654 5871 23706
rect 5923 23654 5937 23706
rect 5989 23654 6425 23706
rect 6477 23654 6491 23706
rect 6543 23654 6979 23706
rect 7031 23654 7045 23706
rect 7097 23654 7533 23706
rect 7585 23654 7599 23706
rect 5299 23636 7651 23654
rect 5299 23584 5317 23636
rect 5369 23584 5383 23636
rect 5435 23584 5871 23636
rect 5923 23584 5937 23636
rect 5989 23584 6425 23636
rect 6477 23584 6491 23636
rect 6543 23584 6979 23636
rect 7031 23584 7045 23636
rect 7097 23584 7533 23636
rect 7585 23584 7599 23636
rect 5299 23566 7651 23584
rect 5299 23514 5317 23566
rect 5369 23514 5383 23566
rect 5435 23514 5871 23566
rect 5923 23514 5937 23566
rect 5989 23514 6425 23566
rect 6477 23514 6491 23566
rect 6543 23514 6979 23566
rect 7031 23514 7045 23566
rect 7097 23514 7533 23566
rect 7585 23514 7599 23566
rect 5299 23496 7651 23514
rect 5299 23444 5317 23496
rect 5369 23444 5383 23496
rect 5435 23444 5871 23496
rect 5923 23444 5937 23496
rect 5989 23444 6425 23496
rect 6477 23444 6491 23496
rect 6543 23444 6979 23496
rect 7031 23444 7045 23496
rect 7097 23444 7533 23496
rect 7585 23444 7599 23496
rect 5299 23426 7651 23444
rect 5299 23374 5317 23426
rect 5369 23374 5383 23426
rect 5435 23374 5871 23426
rect 5923 23374 5937 23426
rect 5989 23374 6425 23426
rect 6477 23374 6491 23426
rect 6543 23374 6979 23426
rect 7031 23374 7045 23426
rect 7097 23374 7533 23426
rect 7585 23374 7599 23426
rect 5299 23371 7651 23374
rect 2724 23368 7651 23371
rect 2270 22728 8222 22730
rect 2270 22724 2648 22728
rect 2322 22672 2392 22724
rect 2444 22676 2648 22724
rect 2700 22676 2713 22728
rect 2765 22676 2778 22728
rect 2830 22676 2843 22728
rect 2895 22676 2908 22728
rect 2960 22676 2973 22728
rect 3025 22676 3038 22728
rect 3090 22676 3103 22728
rect 3155 22676 3168 22728
rect 3220 22676 3233 22728
rect 3285 22676 3298 22728
rect 3350 22676 3363 22728
rect 3415 22676 3428 22728
rect 3480 22676 3493 22728
rect 3545 22676 3558 22728
rect 3610 22676 3623 22728
rect 3675 22676 3688 22728
rect 3740 22676 3753 22728
rect 3805 22676 3818 22728
rect 3870 22676 3883 22728
rect 3935 22676 3948 22728
rect 4000 22676 4013 22728
rect 4065 22676 4078 22728
rect 4130 22676 4143 22728
rect 4195 22676 4208 22728
rect 4260 22676 4273 22728
rect 4325 22676 4338 22728
rect 4390 22676 4403 22728
rect 4455 22676 4468 22728
rect 4520 22676 4532 22728
rect 4584 22724 8222 22728
rect 4584 22720 5613 22724
rect 5669 22720 5696 22724
rect 4584 22676 5040 22720
rect 2444 22672 5040 22676
rect 2270 22668 5040 22672
rect 5092 22668 5106 22720
rect 5158 22668 5594 22720
rect 5752 22668 5779 22724
rect 5835 22668 5861 22724
rect 5917 22668 5943 22724
rect 5999 22668 6025 22724
rect 6081 22668 6107 22724
rect 6163 22720 6189 22724
rect 6245 22720 6271 22724
rect 6266 22668 6271 22720
rect 6327 22668 6353 22724
rect 6409 22668 6435 22724
rect 6491 22668 6517 22724
rect 6573 22668 6599 22724
rect 6655 22668 6681 22724
rect 6737 22720 6763 22724
rect 6819 22720 6845 22724
rect 6754 22668 6763 22720
rect 6820 22668 6845 22720
rect 6901 22668 6927 22724
rect 6983 22668 7009 22724
rect 7065 22668 7091 22724
rect 7147 22668 7173 22724
rect 7229 22668 7255 22724
rect 7311 22720 7337 22724
rect 7311 22668 7322 22720
rect 7393 22668 7419 22724
rect 7475 22668 7501 22724
rect 7557 22668 7583 22724
rect 7639 22668 7665 22724
rect 7721 22668 7747 22724
rect 7803 22720 7829 22724
rect 7885 22720 7911 22724
rect 7803 22668 7810 22720
rect 7967 22668 7993 22724
rect 8049 22668 8075 22672
rect 8131 22668 8157 22724
rect 8221 22672 8222 22724
rect 8213 22668 8222 22672
rect 2270 22660 8222 22668
rect 2270 22655 2648 22660
rect 2322 22603 2392 22655
rect 2444 22608 2648 22655
rect 2700 22608 2713 22660
rect 2765 22608 2778 22660
rect 2830 22608 2843 22660
rect 2895 22608 2908 22660
rect 2960 22608 2973 22660
rect 3025 22608 3038 22660
rect 3090 22608 3103 22660
rect 3155 22608 3168 22660
rect 3220 22608 3233 22660
rect 3285 22608 3298 22660
rect 3350 22608 3363 22660
rect 3415 22608 3428 22660
rect 3480 22608 3493 22660
rect 3545 22608 3558 22660
rect 3610 22608 3623 22660
rect 3675 22608 3688 22660
rect 3740 22608 3753 22660
rect 3805 22608 3818 22660
rect 3870 22608 3883 22660
rect 3935 22608 3948 22660
rect 4000 22608 4013 22660
rect 4065 22608 4078 22660
rect 4130 22608 4143 22660
rect 4195 22608 4208 22660
rect 4260 22608 4273 22660
rect 4325 22608 4338 22660
rect 4390 22608 4403 22660
rect 4455 22608 4468 22660
rect 4520 22608 4532 22660
rect 4584 22655 8222 22660
rect 4584 22651 8047 22655
rect 4584 22608 5040 22651
rect 2444 22603 5040 22608
rect 2270 22599 5040 22603
rect 5092 22599 5106 22651
rect 5158 22599 5594 22651
rect 5646 22644 5660 22651
rect 5712 22644 6148 22651
rect 6200 22644 6214 22651
rect 6266 22644 6702 22651
rect 6754 22644 6768 22651
rect 6820 22644 7256 22651
rect 7308 22644 7322 22651
rect 7374 22644 7810 22651
rect 7862 22644 7876 22651
rect 7928 22644 8047 22651
rect 8099 22644 8169 22655
rect 2270 22592 5613 22599
rect 2270 22586 2648 22592
rect 2322 22534 2392 22586
rect 2444 22540 2648 22586
rect 2700 22540 2713 22592
rect 2765 22540 2778 22592
rect 2830 22540 2843 22592
rect 2895 22540 2908 22592
rect 2960 22540 2973 22592
rect 3025 22540 3038 22592
rect 3090 22540 3103 22592
rect 3155 22540 3168 22592
rect 3220 22540 3233 22592
rect 3285 22540 3298 22592
rect 3350 22540 3363 22592
rect 3415 22540 3428 22592
rect 3480 22540 3493 22592
rect 3545 22540 3558 22592
rect 3610 22540 3623 22592
rect 3675 22540 3688 22592
rect 3740 22540 3753 22592
rect 3805 22540 3818 22592
rect 3870 22540 3883 22592
rect 3935 22540 3948 22592
rect 4000 22540 4013 22592
rect 4065 22540 4078 22592
rect 4130 22540 4143 22592
rect 4195 22540 4208 22592
rect 4260 22540 4273 22592
rect 4325 22540 4338 22592
rect 4390 22540 4403 22592
rect 4455 22540 4468 22592
rect 4520 22540 4532 22592
rect 4584 22588 5613 22592
rect 5669 22588 5696 22599
rect 5752 22588 5779 22644
rect 5835 22588 5861 22644
rect 5917 22588 5943 22644
rect 5999 22588 6025 22644
rect 6081 22588 6107 22644
rect 6266 22599 6271 22644
rect 6163 22588 6189 22599
rect 6245 22588 6271 22599
rect 6327 22588 6353 22644
rect 6409 22588 6435 22644
rect 6491 22588 6517 22644
rect 6573 22588 6599 22644
rect 6655 22588 6681 22644
rect 6754 22599 6763 22644
rect 6820 22599 6845 22644
rect 6737 22588 6763 22599
rect 6819 22588 6845 22599
rect 6901 22588 6927 22644
rect 6983 22588 7009 22644
rect 7065 22588 7091 22644
rect 7147 22588 7173 22644
rect 7229 22588 7255 22644
rect 7311 22599 7322 22644
rect 7311 22588 7337 22599
rect 7393 22588 7419 22644
rect 7475 22588 7501 22644
rect 7557 22588 7583 22644
rect 7639 22588 7665 22644
rect 7721 22588 7747 22644
rect 7803 22599 7810 22644
rect 7803 22588 7829 22599
rect 7885 22588 7911 22599
rect 7967 22588 7993 22644
rect 8049 22588 8075 22603
rect 8131 22588 8157 22644
rect 8221 22603 8222 22655
rect 8213 22588 8222 22603
rect 4584 22586 8222 22588
rect 4584 22582 8047 22586
rect 4584 22540 5040 22582
rect 2444 22534 5040 22540
rect 2270 22530 5040 22534
rect 5092 22530 5106 22582
rect 5158 22530 5594 22582
rect 5646 22564 5660 22582
rect 5712 22564 6148 22582
rect 6200 22564 6214 22582
rect 6266 22564 6702 22582
rect 6754 22564 6768 22582
rect 6820 22564 7256 22582
rect 7308 22564 7322 22582
rect 7374 22564 7810 22582
rect 7862 22564 7876 22582
rect 7928 22564 8047 22582
rect 8099 22564 8169 22586
rect 2270 22524 5613 22530
rect 2270 22517 2648 22524
rect 2322 22465 2392 22517
rect 2444 22472 2648 22517
rect 2700 22472 2713 22524
rect 2765 22472 2778 22524
rect 2830 22472 2843 22524
rect 2895 22472 2908 22524
rect 2960 22472 2973 22524
rect 3025 22472 3038 22524
rect 3090 22472 3103 22524
rect 3155 22472 3168 22524
rect 3220 22472 3233 22524
rect 3285 22472 3298 22524
rect 3350 22472 3363 22524
rect 3415 22472 3428 22524
rect 3480 22472 3493 22524
rect 3545 22472 3558 22524
rect 3610 22472 3623 22524
rect 3675 22472 3688 22524
rect 3740 22472 3753 22524
rect 3805 22472 3818 22524
rect 3870 22472 3883 22524
rect 3935 22472 3948 22524
rect 4000 22472 4013 22524
rect 4065 22472 4078 22524
rect 4130 22472 4143 22524
rect 4195 22472 4208 22524
rect 4260 22472 4273 22524
rect 4325 22472 4338 22524
rect 4390 22472 4403 22524
rect 4455 22472 4468 22524
rect 4520 22472 4532 22524
rect 4584 22513 5613 22524
rect 5669 22513 5696 22530
rect 4584 22472 5040 22513
rect 2444 22465 5040 22472
rect 2270 22461 5040 22465
rect 5092 22461 5106 22513
rect 5158 22461 5594 22513
rect 5752 22508 5779 22564
rect 5835 22508 5861 22564
rect 5917 22508 5943 22564
rect 5999 22508 6025 22564
rect 6081 22508 6107 22564
rect 6266 22530 6271 22564
rect 6163 22513 6189 22530
rect 6245 22513 6271 22530
rect 6266 22508 6271 22513
rect 6327 22508 6353 22564
rect 6409 22508 6435 22564
rect 6491 22508 6517 22564
rect 6573 22508 6599 22564
rect 6655 22508 6681 22564
rect 6754 22530 6763 22564
rect 6820 22530 6845 22564
rect 6737 22513 6763 22530
rect 6819 22513 6845 22530
rect 6754 22508 6763 22513
rect 6820 22508 6845 22513
rect 6901 22508 6927 22564
rect 6983 22508 7009 22564
rect 7065 22508 7091 22564
rect 7147 22508 7173 22564
rect 7229 22508 7255 22564
rect 7311 22530 7322 22564
rect 7311 22513 7337 22530
rect 7311 22508 7322 22513
rect 7393 22508 7419 22564
rect 7475 22508 7501 22564
rect 7557 22508 7583 22564
rect 7639 22508 7665 22564
rect 7721 22508 7747 22564
rect 7803 22530 7810 22564
rect 7803 22513 7829 22530
rect 7885 22513 7911 22530
rect 7803 22508 7810 22513
rect 7967 22508 7993 22564
rect 8049 22517 8075 22534
rect 8131 22508 8157 22564
rect 8221 22534 8222 22586
rect 8213 22517 8222 22534
rect 5646 22484 5660 22508
rect 5712 22484 6148 22508
rect 6200 22484 6214 22508
rect 6266 22484 6702 22508
rect 6754 22484 6768 22508
rect 6820 22484 7256 22508
rect 7308 22484 7322 22508
rect 7374 22484 7810 22508
rect 7862 22484 7876 22508
rect 7928 22484 8047 22508
rect 8099 22484 8169 22508
rect 2270 22456 5613 22461
rect 2270 22448 2648 22456
rect 2322 22396 2392 22448
rect 2444 22404 2648 22448
rect 2700 22404 2713 22456
rect 2765 22404 2778 22456
rect 2830 22404 2843 22456
rect 2895 22404 2908 22456
rect 2960 22404 2973 22456
rect 3025 22404 3038 22456
rect 3090 22404 3103 22456
rect 3155 22404 3168 22456
rect 3220 22404 3233 22456
rect 3285 22404 3298 22456
rect 3350 22404 3363 22456
rect 3415 22404 3428 22456
rect 3480 22404 3493 22456
rect 3545 22404 3558 22456
rect 3610 22404 3623 22456
rect 3675 22404 3688 22456
rect 3740 22404 3753 22456
rect 3805 22404 3818 22456
rect 3870 22404 3883 22456
rect 3935 22404 3948 22456
rect 4000 22404 4013 22456
rect 4065 22404 4078 22456
rect 4130 22404 4143 22456
rect 4195 22404 4208 22456
rect 4260 22404 4273 22456
rect 4325 22404 4338 22456
rect 4390 22404 4403 22456
rect 4455 22404 4468 22456
rect 4520 22404 4532 22456
rect 4584 22444 5613 22456
rect 5669 22444 5696 22461
rect 4584 22404 5040 22444
rect 2444 22396 5040 22404
rect 2270 22392 5040 22396
rect 5092 22392 5106 22444
rect 5158 22392 5594 22444
rect 5752 22428 5779 22484
rect 5835 22428 5861 22484
rect 5917 22428 5943 22484
rect 5999 22428 6025 22484
rect 6081 22428 6107 22484
rect 6266 22461 6271 22484
rect 6163 22444 6189 22461
rect 6245 22444 6271 22461
rect 6266 22428 6271 22444
rect 6327 22428 6353 22484
rect 6409 22428 6435 22484
rect 6491 22428 6517 22484
rect 6573 22428 6599 22484
rect 6655 22428 6681 22484
rect 6754 22461 6763 22484
rect 6820 22461 6845 22484
rect 6737 22444 6763 22461
rect 6819 22444 6845 22461
rect 6754 22428 6763 22444
rect 6820 22428 6845 22444
rect 6901 22428 6927 22484
rect 6983 22428 7009 22484
rect 7065 22428 7091 22484
rect 7147 22428 7173 22484
rect 7229 22428 7255 22484
rect 7311 22461 7322 22484
rect 7311 22444 7337 22461
rect 7311 22428 7322 22444
rect 7393 22428 7419 22484
rect 7475 22428 7501 22484
rect 7557 22428 7583 22484
rect 7639 22428 7665 22484
rect 7721 22428 7747 22484
rect 7803 22461 7810 22484
rect 7803 22444 7829 22461
rect 7885 22444 7911 22461
rect 7803 22428 7810 22444
rect 7967 22428 7993 22484
rect 8049 22448 8075 22465
rect 8131 22428 8157 22484
rect 8221 22465 8222 22517
rect 8213 22448 8222 22465
rect 5646 22404 5660 22428
rect 5712 22404 6148 22428
rect 6200 22404 6214 22428
rect 6266 22404 6702 22428
rect 6754 22404 6768 22428
rect 6820 22404 7256 22428
rect 7308 22404 7322 22428
rect 7374 22404 7810 22428
rect 7862 22404 7876 22428
rect 7928 22404 8047 22428
rect 8099 22404 8169 22428
rect 2270 22388 5613 22392
rect 2270 22378 2648 22388
rect 2322 22326 2392 22378
rect 2444 22336 2648 22378
rect 2700 22336 2713 22388
rect 2765 22336 2778 22388
rect 2830 22336 2843 22388
rect 2895 22336 2908 22388
rect 2960 22336 2973 22388
rect 3025 22336 3038 22388
rect 3090 22336 3103 22388
rect 3155 22336 3168 22388
rect 3220 22336 3233 22388
rect 3285 22336 3298 22388
rect 3350 22336 3363 22388
rect 3415 22336 3428 22388
rect 3480 22336 3493 22388
rect 3545 22336 3558 22388
rect 3610 22336 3623 22388
rect 3675 22336 3688 22388
rect 3740 22336 3753 22388
rect 3805 22336 3818 22388
rect 3870 22336 3883 22388
rect 3935 22336 3948 22388
rect 4000 22336 4013 22388
rect 4065 22336 4078 22388
rect 4130 22336 4143 22388
rect 4195 22336 4208 22388
rect 4260 22336 4273 22388
rect 4325 22336 4338 22388
rect 4390 22336 4403 22388
rect 4455 22336 4468 22388
rect 4520 22336 4532 22388
rect 4584 22375 5613 22388
rect 5669 22375 5696 22392
rect 4584 22336 5040 22375
rect 2444 22326 5040 22336
rect 2270 22323 5040 22326
rect 5092 22323 5106 22375
rect 5158 22323 5594 22375
rect 5752 22348 5779 22404
rect 5835 22348 5861 22404
rect 5917 22348 5943 22404
rect 5999 22348 6025 22404
rect 6081 22348 6107 22404
rect 6266 22392 6271 22404
rect 6163 22375 6189 22392
rect 6245 22375 6271 22392
rect 6266 22348 6271 22375
rect 6327 22348 6353 22404
rect 6409 22348 6435 22404
rect 6491 22348 6517 22404
rect 6573 22348 6599 22404
rect 6655 22348 6681 22404
rect 6754 22392 6763 22404
rect 6820 22392 6845 22404
rect 6737 22375 6763 22392
rect 6819 22375 6845 22392
rect 6754 22348 6763 22375
rect 6820 22348 6845 22375
rect 6901 22348 6927 22404
rect 6983 22348 7009 22404
rect 7065 22348 7091 22404
rect 7147 22348 7173 22404
rect 7229 22348 7255 22404
rect 7311 22392 7322 22404
rect 7311 22375 7337 22392
rect 7311 22348 7322 22375
rect 7393 22348 7419 22404
rect 7475 22348 7501 22404
rect 7557 22348 7583 22404
rect 7639 22348 7665 22404
rect 7721 22348 7747 22404
rect 7803 22392 7810 22404
rect 7803 22375 7829 22392
rect 7885 22375 7911 22392
rect 7803 22348 7810 22375
rect 7967 22348 7993 22404
rect 8049 22378 8075 22396
rect 8131 22348 8157 22404
rect 8221 22396 8222 22448
rect 8213 22378 8222 22396
rect 5646 22324 5660 22348
rect 5712 22324 6148 22348
rect 6200 22324 6214 22348
rect 6266 22324 6702 22348
rect 6754 22324 6768 22348
rect 6820 22324 7256 22348
rect 7308 22324 7322 22348
rect 7374 22324 7810 22348
rect 7862 22324 7876 22348
rect 7928 22326 8047 22348
rect 8099 22326 8169 22348
rect 8221 22326 8222 22378
rect 7928 22324 8222 22326
rect 2270 22320 5613 22323
rect 2270 22308 2648 22320
rect 2322 22256 2392 22308
rect 2444 22268 2648 22308
rect 2700 22268 2713 22320
rect 2765 22268 2778 22320
rect 2830 22268 2843 22320
rect 2895 22268 2908 22320
rect 2960 22268 2973 22320
rect 3025 22268 3038 22320
rect 3090 22268 3103 22320
rect 3155 22268 3168 22320
rect 3220 22268 3233 22320
rect 3285 22268 3298 22320
rect 3350 22268 3363 22320
rect 3415 22268 3428 22320
rect 3480 22268 3493 22320
rect 3545 22268 3558 22320
rect 3610 22268 3623 22320
rect 3675 22268 3688 22320
rect 3740 22268 3753 22320
rect 3805 22268 3818 22320
rect 3870 22268 3883 22320
rect 3935 22268 3948 22320
rect 4000 22268 4013 22320
rect 4065 22268 4078 22320
rect 4130 22268 4143 22320
rect 4195 22268 4208 22320
rect 4260 22268 4273 22320
rect 4325 22268 4338 22320
rect 4390 22268 4403 22320
rect 4455 22268 4468 22320
rect 4520 22268 4532 22320
rect 4584 22306 5613 22320
rect 5669 22306 5696 22323
rect 4584 22268 5040 22306
rect 2444 22256 5040 22268
rect 2270 22254 5040 22256
rect 5092 22254 5106 22306
rect 5158 22254 5594 22306
rect 5752 22268 5779 22324
rect 5835 22268 5861 22324
rect 5917 22268 5943 22324
rect 5999 22268 6025 22324
rect 6081 22268 6107 22324
rect 6266 22323 6271 22324
rect 6163 22306 6189 22323
rect 6245 22306 6271 22323
rect 6266 22268 6271 22306
rect 6327 22268 6353 22324
rect 6409 22268 6435 22324
rect 6491 22268 6517 22324
rect 6573 22268 6599 22324
rect 6655 22268 6681 22324
rect 6754 22323 6763 22324
rect 6820 22323 6845 22324
rect 6737 22306 6763 22323
rect 6819 22306 6845 22323
rect 6754 22268 6763 22306
rect 6820 22268 6845 22306
rect 6901 22268 6927 22324
rect 6983 22268 7009 22324
rect 7065 22268 7091 22324
rect 7147 22268 7173 22324
rect 7229 22268 7255 22324
rect 7311 22323 7322 22324
rect 7311 22306 7337 22323
rect 7311 22268 7322 22306
rect 7393 22268 7419 22324
rect 7475 22268 7501 22324
rect 7557 22268 7583 22324
rect 7639 22268 7665 22324
rect 7721 22268 7747 22324
rect 7803 22323 7810 22324
rect 7803 22306 7829 22323
rect 7885 22306 7911 22323
rect 7803 22268 7810 22306
rect 7967 22268 7993 22324
rect 8049 22308 8075 22324
rect 8131 22268 8157 22324
rect 8213 22308 8222 22324
rect 5646 22254 5660 22268
rect 5712 22254 6148 22268
rect 6200 22254 6214 22268
rect 6266 22254 6702 22268
rect 6754 22254 6768 22268
rect 6820 22254 7256 22268
rect 7308 22254 7322 22268
rect 7374 22254 7810 22268
rect 7862 22254 7876 22268
rect 7928 22256 8047 22268
rect 8099 22256 8169 22268
rect 8221 22256 8222 22308
rect 7928 22254 8222 22256
rect 2270 22252 8222 22254
rect 2270 22238 2648 22252
rect 2322 22186 2392 22238
rect 2444 22200 2648 22238
rect 2700 22200 2713 22252
rect 2765 22200 2778 22252
rect 2830 22200 2843 22252
rect 2895 22200 2908 22252
rect 2960 22200 2973 22252
rect 3025 22200 3038 22252
rect 3090 22200 3103 22252
rect 3155 22200 3168 22252
rect 3220 22200 3233 22252
rect 3285 22200 3298 22252
rect 3350 22200 3363 22252
rect 3415 22200 3428 22252
rect 3480 22200 3493 22252
rect 3545 22200 3558 22252
rect 3610 22200 3623 22252
rect 3675 22200 3688 22252
rect 3740 22200 3753 22252
rect 3805 22200 3818 22252
rect 3870 22200 3883 22252
rect 3935 22200 3948 22252
rect 4000 22200 4013 22252
rect 4065 22200 4078 22252
rect 4130 22200 4143 22252
rect 4195 22200 4208 22252
rect 4260 22200 4273 22252
rect 4325 22200 4338 22252
rect 4390 22200 4403 22252
rect 4455 22200 4468 22252
rect 4520 22200 4532 22252
rect 4584 22244 8222 22252
rect 4584 22236 5613 22244
rect 5669 22236 5696 22244
rect 4584 22200 5040 22236
rect 2444 22186 5040 22200
rect 2270 22184 5040 22186
rect 5092 22184 5106 22236
rect 5158 22184 5594 22236
rect 5752 22188 5779 22244
rect 5835 22188 5861 22244
rect 5917 22188 5943 22244
rect 5999 22188 6025 22244
rect 6081 22188 6107 22244
rect 6163 22236 6189 22244
rect 6245 22236 6271 22244
rect 6266 22188 6271 22236
rect 6327 22188 6353 22244
rect 6409 22188 6435 22244
rect 6491 22188 6517 22244
rect 6573 22188 6599 22244
rect 6655 22188 6681 22244
rect 6737 22236 6763 22244
rect 6819 22236 6845 22244
rect 6754 22188 6763 22236
rect 6820 22188 6845 22236
rect 6901 22188 6927 22244
rect 6983 22188 7009 22244
rect 7065 22188 7091 22244
rect 7147 22188 7173 22244
rect 7229 22188 7255 22244
rect 7311 22236 7337 22244
rect 7311 22188 7322 22236
rect 7393 22188 7419 22244
rect 7475 22188 7501 22244
rect 7557 22188 7583 22244
rect 7639 22188 7665 22244
rect 7721 22188 7747 22244
rect 7803 22236 7829 22244
rect 7885 22236 7911 22244
rect 7803 22188 7810 22236
rect 7967 22188 7993 22244
rect 8049 22238 8075 22244
rect 8131 22188 8157 22244
rect 8213 22238 8222 22244
rect 5646 22184 5660 22188
rect 5712 22184 6148 22188
rect 6200 22184 6214 22188
rect 6266 22184 6702 22188
rect 6754 22184 6768 22188
rect 6820 22184 7256 22188
rect 7308 22184 7322 22188
rect 7374 22184 7810 22188
rect 7862 22184 7876 22188
rect 7928 22186 8047 22188
rect 8099 22186 8169 22188
rect 8221 22186 8222 22238
rect 7928 22184 8222 22186
rect 2270 22168 8222 22184
rect 2322 22116 2392 22168
rect 2444 22166 8047 22168
rect 2444 22116 5040 22166
rect 2270 22114 5040 22116
rect 5092 22114 5106 22166
rect 5158 22114 5594 22166
rect 5646 22164 5660 22166
rect 5712 22164 6148 22166
rect 6200 22164 6214 22166
rect 6266 22164 6702 22166
rect 6754 22164 6768 22166
rect 6820 22164 7256 22166
rect 7308 22164 7322 22166
rect 7374 22164 7810 22166
rect 7862 22164 7876 22166
rect 7928 22164 8047 22166
rect 8099 22164 8169 22168
rect 2270 22108 5613 22114
rect 5669 22108 5696 22114
rect 5752 22108 5779 22164
rect 5835 22108 5861 22164
rect 5917 22108 5943 22164
rect 5999 22108 6025 22164
rect 6081 22108 6107 22164
rect 6266 22114 6271 22164
rect 6163 22108 6189 22114
rect 6245 22108 6271 22114
rect 6327 22108 6353 22164
rect 6409 22108 6435 22164
rect 6491 22108 6517 22164
rect 6573 22108 6599 22164
rect 6655 22108 6681 22164
rect 6754 22114 6763 22164
rect 6820 22114 6845 22164
rect 6737 22108 6763 22114
rect 6819 22108 6845 22114
rect 6901 22108 6927 22164
rect 6983 22108 7009 22164
rect 7065 22108 7091 22164
rect 7147 22108 7173 22164
rect 7229 22108 7255 22164
rect 7311 22114 7322 22164
rect 7311 22108 7337 22114
rect 7393 22108 7419 22164
rect 7475 22108 7501 22164
rect 7557 22108 7583 22164
rect 7639 22108 7665 22164
rect 7721 22108 7747 22164
rect 7803 22114 7810 22164
rect 7803 22108 7829 22114
rect 7885 22108 7911 22114
rect 7967 22108 7993 22164
rect 8049 22108 8075 22116
rect 8131 22108 8157 22164
rect 8221 22116 8222 22168
rect 8213 22108 8222 22116
rect 2724 21987 7651 21988
rect 2724 21931 2733 21987
rect 2789 21931 2814 21987
rect 2870 21931 2895 21987
rect 2951 21931 2976 21987
rect 3032 21931 3057 21987
rect 3113 21931 3138 21987
rect 3194 21931 3219 21987
rect 3275 21931 3300 21987
rect 3356 21931 3381 21987
rect 3437 21931 3462 21987
rect 3518 21931 3543 21987
rect 3599 21931 3624 21987
rect 3680 21931 3705 21987
rect 3761 21931 3786 21987
rect 3842 21931 3867 21987
rect 3923 21931 3948 21987
rect 4004 21931 4029 21987
rect 4085 21931 4110 21987
rect 4166 21931 4191 21987
rect 4247 21931 4272 21987
rect 4328 21931 4353 21987
rect 4409 21931 4434 21987
rect 4490 21931 4515 21987
rect 4571 21931 4596 21987
rect 4652 21931 4677 21987
rect 4733 21931 4758 21987
rect 4814 21931 4839 21987
rect 4895 21931 4920 21987
rect 4976 21931 5001 21987
rect 5057 21931 5082 21987
rect 5138 21931 5163 21987
rect 2724 21907 5163 21931
rect 2724 21851 2733 21907
rect 2789 21851 2814 21907
rect 2870 21851 2895 21907
rect 2951 21851 2976 21907
rect 3032 21851 3057 21907
rect 3113 21851 3138 21907
rect 3194 21851 3219 21907
rect 3275 21851 3300 21907
rect 3356 21851 3381 21907
rect 3437 21851 3462 21907
rect 3518 21851 3543 21907
rect 3599 21851 3624 21907
rect 3680 21851 3705 21907
rect 3761 21851 3786 21907
rect 3842 21851 3867 21907
rect 3923 21851 3948 21907
rect 4004 21851 4029 21907
rect 4085 21851 4110 21907
rect 4166 21851 4191 21907
rect 4247 21851 4272 21907
rect 4328 21851 4353 21907
rect 4409 21851 4434 21907
rect 4490 21851 4515 21907
rect 4571 21851 4596 21907
rect 4652 21851 4677 21907
rect 4733 21851 4758 21907
rect 4814 21851 4839 21907
rect 4895 21851 4920 21907
rect 4976 21851 5001 21907
rect 5057 21851 5082 21907
rect 5138 21851 5163 21907
rect 2724 21827 5163 21851
rect 2724 21771 2733 21827
rect 2789 21771 2814 21827
rect 2870 21771 2895 21827
rect 2951 21771 2976 21827
rect 3032 21771 3057 21827
rect 3113 21771 3138 21827
rect 3194 21771 3219 21827
rect 3275 21771 3300 21827
rect 3356 21771 3381 21827
rect 3437 21771 3462 21827
rect 3518 21771 3543 21827
rect 3599 21771 3624 21827
rect 3680 21771 3705 21827
rect 3761 21771 3786 21827
rect 3842 21771 3867 21827
rect 3923 21771 3948 21827
rect 4004 21771 4029 21827
rect 4085 21771 4110 21827
rect 4166 21771 4191 21827
rect 4247 21771 4272 21827
rect 4328 21771 4353 21827
rect 4409 21771 4434 21827
rect 4490 21771 4515 21827
rect 4571 21771 4596 21827
rect 4652 21771 4677 21827
rect 4733 21771 4758 21827
rect 4814 21771 4839 21827
rect 4895 21771 4920 21827
rect 4976 21771 5001 21827
rect 5057 21771 5082 21827
rect 5138 21771 5163 21827
rect 2724 21747 5163 21771
rect 2724 21691 2733 21747
rect 2789 21691 2814 21747
rect 2870 21691 2895 21747
rect 2951 21691 2976 21747
rect 3032 21691 3057 21747
rect 3113 21691 3138 21747
rect 3194 21691 3219 21747
rect 3275 21691 3300 21747
rect 3356 21691 3381 21747
rect 3437 21691 3462 21747
rect 3518 21691 3543 21747
rect 3599 21691 3624 21747
rect 3680 21691 3705 21747
rect 3761 21691 3786 21747
rect 3842 21691 3867 21747
rect 3923 21691 3948 21747
rect 4004 21691 4029 21747
rect 4085 21691 4110 21747
rect 4166 21691 4191 21747
rect 4247 21691 4272 21747
rect 4328 21691 4353 21747
rect 4409 21691 4434 21747
rect 4490 21691 4515 21747
rect 4571 21691 4596 21747
rect 4652 21691 4677 21747
rect 4733 21691 4758 21747
rect 4814 21691 4839 21747
rect 4895 21691 4920 21747
rect 4976 21691 5001 21747
rect 5057 21691 5082 21747
rect 5138 21691 5163 21747
rect 2724 21667 5163 21691
rect 2724 21611 2733 21667
rect 2789 21611 2814 21667
rect 2870 21611 2895 21667
rect 2951 21611 2976 21667
rect 3032 21611 3057 21667
rect 3113 21611 3138 21667
rect 3194 21611 3219 21667
rect 3275 21611 3300 21667
rect 3356 21611 3381 21667
rect 3437 21611 3462 21667
rect 3518 21611 3543 21667
rect 3599 21611 3624 21667
rect 3680 21611 3705 21667
rect 3761 21611 3786 21667
rect 3842 21611 3867 21667
rect 3923 21611 3948 21667
rect 4004 21611 4029 21667
rect 4085 21611 4110 21667
rect 4166 21611 4191 21667
rect 4247 21611 4272 21667
rect 4328 21611 4353 21667
rect 4409 21611 4434 21667
rect 4490 21611 4515 21667
rect 4571 21611 4596 21667
rect 4652 21611 4677 21667
rect 4733 21611 4758 21667
rect 4814 21611 4839 21667
rect 4895 21611 4920 21667
rect 4976 21611 5001 21667
rect 5057 21611 5082 21667
rect 5138 21611 5163 21667
rect 2724 21587 5163 21611
rect 2724 21531 2733 21587
rect 2789 21531 2814 21587
rect 2870 21531 2895 21587
rect 2951 21531 2976 21587
rect 3032 21531 3057 21587
rect 3113 21531 3138 21587
rect 3194 21531 3219 21587
rect 3275 21531 3300 21587
rect 3356 21531 3381 21587
rect 3437 21531 3462 21587
rect 3518 21531 3543 21587
rect 3599 21531 3624 21587
rect 3680 21531 3705 21587
rect 3761 21531 3786 21587
rect 3842 21531 3867 21587
rect 3923 21531 3948 21587
rect 4004 21531 4029 21587
rect 4085 21531 4110 21587
rect 4166 21531 4191 21587
rect 4247 21531 4272 21587
rect 4328 21531 4353 21587
rect 4409 21531 4434 21587
rect 4490 21531 4515 21587
rect 4571 21531 4596 21587
rect 4652 21531 4677 21587
rect 4733 21531 4758 21587
rect 4814 21531 4839 21587
rect 4895 21531 4920 21587
rect 4976 21531 5001 21587
rect 5057 21531 5082 21587
rect 5138 21531 5163 21587
rect 2724 21507 5163 21531
rect 2724 21451 2733 21507
rect 2789 21451 2814 21507
rect 2870 21451 2895 21507
rect 2951 21451 2976 21507
rect 3032 21451 3057 21507
rect 3113 21451 3138 21507
rect 3194 21451 3219 21507
rect 3275 21451 3300 21507
rect 3356 21451 3381 21507
rect 3437 21451 3462 21507
rect 3518 21451 3543 21507
rect 3599 21451 3624 21507
rect 3680 21451 3705 21507
rect 3761 21451 3786 21507
rect 3842 21451 3867 21507
rect 3923 21451 3948 21507
rect 4004 21451 4029 21507
rect 4085 21451 4110 21507
rect 4166 21451 4191 21507
rect 4247 21451 4272 21507
rect 4328 21451 4353 21507
rect 4409 21451 4434 21507
rect 4490 21451 4515 21507
rect 4571 21451 4596 21507
rect 4652 21451 4677 21507
rect 4733 21451 4758 21507
rect 4814 21451 4839 21507
rect 4895 21451 4920 21507
rect 4976 21451 5001 21507
rect 5057 21451 5082 21507
rect 5138 21451 5163 21507
rect 2724 21427 5163 21451
rect 2724 21371 2733 21427
rect 2789 21371 2814 21427
rect 2870 21371 2895 21427
rect 2951 21371 2976 21427
rect 3032 21371 3057 21427
rect 3113 21371 3138 21427
rect 3194 21371 3219 21427
rect 3275 21371 3300 21427
rect 3356 21371 3381 21427
rect 3437 21371 3462 21427
rect 3518 21371 3543 21427
rect 3599 21371 3624 21427
rect 3680 21371 3705 21427
rect 3761 21371 3786 21427
rect 3842 21371 3867 21427
rect 3923 21371 3948 21427
rect 4004 21371 4029 21427
rect 4085 21371 4110 21427
rect 4166 21371 4191 21427
rect 4247 21371 4272 21427
rect 4328 21371 4353 21427
rect 4409 21371 4434 21427
rect 4490 21371 4515 21427
rect 4571 21371 4596 21427
rect 4652 21371 4677 21427
rect 4733 21371 4758 21427
rect 4814 21371 4839 21427
rect 4895 21371 4920 21427
rect 4976 21371 5001 21427
rect 5057 21371 5082 21427
rect 5138 21371 5163 21427
rect 5299 21982 7651 21987
rect 5299 21930 5317 21982
rect 5369 21930 5383 21982
rect 5435 21930 5871 21982
rect 5923 21930 5937 21982
rect 5989 21930 6425 21982
rect 6477 21930 6491 21982
rect 6543 21930 6979 21982
rect 7031 21930 7045 21982
rect 7097 21930 7533 21982
rect 7585 21930 7599 21982
rect 5299 21913 7651 21930
rect 5299 21861 5317 21913
rect 5369 21861 5383 21913
rect 5435 21861 5871 21913
rect 5923 21861 5937 21913
rect 5989 21861 6425 21913
rect 6477 21861 6491 21913
rect 6543 21861 6979 21913
rect 7031 21861 7045 21913
rect 7097 21861 7533 21913
rect 7585 21861 7599 21913
rect 5299 21844 7651 21861
rect 5299 21792 5317 21844
rect 5369 21792 5383 21844
rect 5435 21792 5871 21844
rect 5923 21792 5937 21844
rect 5989 21792 6425 21844
rect 6477 21792 6491 21844
rect 6543 21792 6979 21844
rect 7031 21792 7045 21844
rect 7097 21792 7533 21844
rect 7585 21792 7599 21844
rect 5299 21775 7651 21792
rect 5299 21723 5317 21775
rect 5369 21723 5383 21775
rect 5435 21723 5871 21775
rect 5923 21723 5937 21775
rect 5989 21723 6425 21775
rect 6477 21723 6491 21775
rect 6543 21723 6979 21775
rect 7031 21723 7045 21775
rect 7097 21723 7533 21775
rect 7585 21723 7599 21775
rect 5299 21706 7651 21723
rect 5299 21654 5317 21706
rect 5369 21654 5383 21706
rect 5435 21654 5871 21706
rect 5923 21654 5937 21706
rect 5989 21654 6425 21706
rect 6477 21654 6491 21706
rect 6543 21654 6979 21706
rect 7031 21654 7045 21706
rect 7097 21654 7533 21706
rect 7585 21654 7599 21706
rect 5299 21636 7651 21654
rect 5299 21584 5317 21636
rect 5369 21584 5383 21636
rect 5435 21584 5871 21636
rect 5923 21584 5937 21636
rect 5989 21584 6425 21636
rect 6477 21584 6491 21636
rect 6543 21584 6979 21636
rect 7031 21584 7045 21636
rect 7097 21584 7533 21636
rect 7585 21584 7599 21636
rect 5299 21566 7651 21584
rect 5299 21514 5317 21566
rect 5369 21514 5383 21566
rect 5435 21514 5871 21566
rect 5923 21514 5937 21566
rect 5989 21514 6425 21566
rect 6477 21514 6491 21566
rect 6543 21514 6979 21566
rect 7031 21514 7045 21566
rect 7097 21514 7533 21566
rect 7585 21514 7599 21566
rect 5299 21496 7651 21514
rect 5299 21444 5317 21496
rect 5369 21444 5383 21496
rect 5435 21444 5871 21496
rect 5923 21444 5937 21496
rect 5989 21444 6425 21496
rect 6477 21444 6491 21496
rect 6543 21444 6979 21496
rect 7031 21444 7045 21496
rect 7097 21444 7533 21496
rect 7585 21444 7599 21496
rect 5299 21426 7651 21444
rect 5299 21374 5317 21426
rect 5369 21374 5383 21426
rect 5435 21374 5871 21426
rect 5923 21374 5937 21426
rect 5989 21374 6425 21426
rect 6477 21374 6491 21426
rect 6543 21374 6979 21426
rect 7031 21374 7045 21426
rect 7097 21374 7533 21426
rect 7585 21374 7599 21426
rect 5299 21371 7651 21374
rect 2724 21368 7651 21371
rect 2270 20728 8222 20730
rect 2270 20724 2648 20728
rect 2322 20672 2392 20724
rect 2444 20676 2648 20724
rect 2700 20676 2713 20728
rect 2765 20676 2778 20728
rect 2830 20676 2843 20728
rect 2895 20676 2908 20728
rect 2960 20676 2973 20728
rect 3025 20676 3038 20728
rect 3090 20676 3103 20728
rect 3155 20676 3168 20728
rect 3220 20676 3233 20728
rect 3285 20676 3298 20728
rect 3350 20676 3363 20728
rect 3415 20676 3428 20728
rect 3480 20676 3493 20728
rect 3545 20676 3558 20728
rect 3610 20676 3623 20728
rect 3675 20676 3688 20728
rect 3740 20676 3753 20728
rect 3805 20676 3818 20728
rect 3870 20676 3883 20728
rect 3935 20676 3948 20728
rect 4000 20676 4013 20728
rect 4065 20676 4078 20728
rect 4130 20676 4143 20728
rect 4195 20676 4208 20728
rect 4260 20676 4273 20728
rect 4325 20676 4338 20728
rect 4390 20676 4403 20728
rect 4455 20676 4468 20728
rect 4520 20676 4532 20728
rect 4584 20724 8222 20728
rect 4584 20720 5613 20724
rect 5669 20720 5696 20724
rect 4584 20676 5040 20720
rect 2444 20672 5040 20676
rect 2270 20668 5040 20672
rect 5092 20668 5106 20720
rect 5158 20668 5594 20720
rect 5752 20668 5779 20724
rect 5835 20668 5861 20724
rect 5917 20668 5943 20724
rect 5999 20668 6025 20724
rect 6081 20668 6107 20724
rect 6163 20720 6189 20724
rect 6245 20720 6271 20724
rect 6266 20668 6271 20720
rect 6327 20668 6353 20724
rect 6409 20668 6435 20724
rect 6491 20668 6517 20724
rect 6573 20668 6599 20724
rect 6655 20668 6681 20724
rect 6737 20720 6763 20724
rect 6819 20720 6845 20724
rect 6754 20668 6763 20720
rect 6820 20668 6845 20720
rect 6901 20668 6927 20724
rect 6983 20668 7009 20724
rect 7065 20668 7091 20724
rect 7147 20668 7173 20724
rect 7229 20668 7255 20724
rect 7311 20720 7337 20724
rect 7311 20668 7322 20720
rect 7393 20668 7419 20724
rect 7475 20668 7501 20724
rect 7557 20668 7583 20724
rect 7639 20668 7665 20724
rect 7721 20668 7747 20724
rect 7803 20720 7829 20724
rect 7885 20720 7911 20724
rect 7803 20668 7810 20720
rect 7967 20668 7993 20724
rect 8049 20668 8075 20672
rect 8131 20668 8157 20724
rect 8221 20672 8222 20724
rect 8213 20668 8222 20672
rect 2270 20660 8222 20668
rect 2270 20655 2648 20660
rect 2322 20603 2392 20655
rect 2444 20608 2648 20655
rect 2700 20608 2713 20660
rect 2765 20608 2778 20660
rect 2830 20608 2843 20660
rect 2895 20608 2908 20660
rect 2960 20608 2973 20660
rect 3025 20608 3038 20660
rect 3090 20608 3103 20660
rect 3155 20608 3168 20660
rect 3220 20608 3233 20660
rect 3285 20608 3298 20660
rect 3350 20608 3363 20660
rect 3415 20608 3428 20660
rect 3480 20608 3493 20660
rect 3545 20608 3558 20660
rect 3610 20608 3623 20660
rect 3675 20608 3688 20660
rect 3740 20608 3753 20660
rect 3805 20608 3818 20660
rect 3870 20608 3883 20660
rect 3935 20608 3948 20660
rect 4000 20608 4013 20660
rect 4065 20608 4078 20660
rect 4130 20608 4143 20660
rect 4195 20608 4208 20660
rect 4260 20608 4273 20660
rect 4325 20608 4338 20660
rect 4390 20608 4403 20660
rect 4455 20608 4468 20660
rect 4520 20608 4532 20660
rect 4584 20655 8222 20660
rect 4584 20651 8047 20655
rect 4584 20608 5040 20651
rect 2444 20603 5040 20608
rect 2270 20599 5040 20603
rect 5092 20599 5106 20651
rect 5158 20599 5594 20651
rect 5646 20644 5660 20651
rect 5712 20644 6148 20651
rect 6200 20644 6214 20651
rect 6266 20644 6702 20651
rect 6754 20644 6768 20651
rect 6820 20644 7256 20651
rect 7308 20644 7322 20651
rect 7374 20644 7810 20651
rect 7862 20644 7876 20651
rect 7928 20644 8047 20651
rect 8099 20644 8169 20655
rect 2270 20592 5613 20599
rect 2270 20586 2648 20592
rect 2322 20534 2392 20586
rect 2444 20540 2648 20586
rect 2700 20540 2713 20592
rect 2765 20540 2778 20592
rect 2830 20540 2843 20592
rect 2895 20540 2908 20592
rect 2960 20540 2973 20592
rect 3025 20540 3038 20592
rect 3090 20540 3103 20592
rect 3155 20540 3168 20592
rect 3220 20540 3233 20592
rect 3285 20540 3298 20592
rect 3350 20540 3363 20592
rect 3415 20540 3428 20592
rect 3480 20540 3493 20592
rect 3545 20540 3558 20592
rect 3610 20540 3623 20592
rect 3675 20540 3688 20592
rect 3740 20540 3753 20592
rect 3805 20540 3818 20592
rect 3870 20540 3883 20592
rect 3935 20540 3948 20592
rect 4000 20540 4013 20592
rect 4065 20540 4078 20592
rect 4130 20540 4143 20592
rect 4195 20540 4208 20592
rect 4260 20540 4273 20592
rect 4325 20540 4338 20592
rect 4390 20540 4403 20592
rect 4455 20540 4468 20592
rect 4520 20540 4532 20592
rect 4584 20588 5613 20592
rect 5669 20588 5696 20599
rect 5752 20588 5779 20644
rect 5835 20588 5861 20644
rect 5917 20588 5943 20644
rect 5999 20588 6025 20644
rect 6081 20588 6107 20644
rect 6266 20599 6271 20644
rect 6163 20588 6189 20599
rect 6245 20588 6271 20599
rect 6327 20588 6353 20644
rect 6409 20588 6435 20644
rect 6491 20588 6517 20644
rect 6573 20588 6599 20644
rect 6655 20588 6681 20644
rect 6754 20599 6763 20644
rect 6820 20599 6845 20644
rect 6737 20588 6763 20599
rect 6819 20588 6845 20599
rect 6901 20588 6927 20644
rect 6983 20588 7009 20644
rect 7065 20588 7091 20644
rect 7147 20588 7173 20644
rect 7229 20588 7255 20644
rect 7311 20599 7322 20644
rect 7311 20588 7337 20599
rect 7393 20588 7419 20644
rect 7475 20588 7501 20644
rect 7557 20588 7583 20644
rect 7639 20588 7665 20644
rect 7721 20588 7747 20644
rect 7803 20599 7810 20644
rect 7803 20588 7829 20599
rect 7885 20588 7911 20599
rect 7967 20588 7993 20644
rect 8049 20588 8075 20603
rect 8131 20588 8157 20644
rect 8221 20603 8222 20655
rect 8213 20588 8222 20603
rect 4584 20586 8222 20588
rect 4584 20582 8047 20586
rect 4584 20540 5040 20582
rect 2444 20534 5040 20540
rect 2270 20530 5040 20534
rect 5092 20530 5106 20582
rect 5158 20530 5594 20582
rect 5646 20564 5660 20582
rect 5712 20564 6148 20582
rect 6200 20564 6214 20582
rect 6266 20564 6702 20582
rect 6754 20564 6768 20582
rect 6820 20564 7256 20582
rect 7308 20564 7322 20582
rect 7374 20564 7810 20582
rect 7862 20564 7876 20582
rect 7928 20564 8047 20582
rect 8099 20564 8169 20586
rect 2270 20524 5613 20530
rect 2270 20517 2648 20524
rect 2322 20465 2392 20517
rect 2444 20472 2648 20517
rect 2700 20472 2713 20524
rect 2765 20472 2778 20524
rect 2830 20472 2843 20524
rect 2895 20472 2908 20524
rect 2960 20472 2973 20524
rect 3025 20472 3038 20524
rect 3090 20472 3103 20524
rect 3155 20472 3168 20524
rect 3220 20472 3233 20524
rect 3285 20472 3298 20524
rect 3350 20472 3363 20524
rect 3415 20472 3428 20524
rect 3480 20472 3493 20524
rect 3545 20472 3558 20524
rect 3610 20472 3623 20524
rect 3675 20472 3688 20524
rect 3740 20472 3753 20524
rect 3805 20472 3818 20524
rect 3870 20472 3883 20524
rect 3935 20472 3948 20524
rect 4000 20472 4013 20524
rect 4065 20472 4078 20524
rect 4130 20472 4143 20524
rect 4195 20472 4208 20524
rect 4260 20472 4273 20524
rect 4325 20472 4338 20524
rect 4390 20472 4403 20524
rect 4455 20472 4468 20524
rect 4520 20472 4532 20524
rect 4584 20513 5613 20524
rect 5669 20513 5696 20530
rect 4584 20472 5040 20513
rect 2444 20465 5040 20472
rect 2270 20461 5040 20465
rect 5092 20461 5106 20513
rect 5158 20461 5594 20513
rect 5752 20508 5779 20564
rect 5835 20508 5861 20564
rect 5917 20508 5943 20564
rect 5999 20508 6025 20564
rect 6081 20508 6107 20564
rect 6266 20530 6271 20564
rect 6163 20513 6189 20530
rect 6245 20513 6271 20530
rect 6266 20508 6271 20513
rect 6327 20508 6353 20564
rect 6409 20508 6435 20564
rect 6491 20508 6517 20564
rect 6573 20508 6599 20564
rect 6655 20508 6681 20564
rect 6754 20530 6763 20564
rect 6820 20530 6845 20564
rect 6737 20513 6763 20530
rect 6819 20513 6845 20530
rect 6754 20508 6763 20513
rect 6820 20508 6845 20513
rect 6901 20508 6927 20564
rect 6983 20508 7009 20564
rect 7065 20508 7091 20564
rect 7147 20508 7173 20564
rect 7229 20508 7255 20564
rect 7311 20530 7322 20564
rect 7311 20513 7337 20530
rect 7311 20508 7322 20513
rect 7393 20508 7419 20564
rect 7475 20508 7501 20564
rect 7557 20508 7583 20564
rect 7639 20508 7665 20564
rect 7721 20508 7747 20564
rect 7803 20530 7810 20564
rect 7803 20513 7829 20530
rect 7885 20513 7911 20530
rect 7803 20508 7810 20513
rect 7967 20508 7993 20564
rect 8049 20517 8075 20534
rect 8131 20508 8157 20564
rect 8221 20534 8222 20586
rect 8213 20517 8222 20534
rect 5646 20484 5660 20508
rect 5712 20484 6148 20508
rect 6200 20484 6214 20508
rect 6266 20484 6702 20508
rect 6754 20484 6768 20508
rect 6820 20484 7256 20508
rect 7308 20484 7322 20508
rect 7374 20484 7810 20508
rect 7862 20484 7876 20508
rect 7928 20484 8047 20508
rect 8099 20484 8169 20508
rect 2270 20456 5613 20461
rect 2270 20448 2648 20456
rect 2322 20396 2392 20448
rect 2444 20404 2648 20448
rect 2700 20404 2713 20456
rect 2765 20404 2778 20456
rect 2830 20404 2843 20456
rect 2895 20404 2908 20456
rect 2960 20404 2973 20456
rect 3025 20404 3038 20456
rect 3090 20404 3103 20456
rect 3155 20404 3168 20456
rect 3220 20404 3233 20456
rect 3285 20404 3298 20456
rect 3350 20404 3363 20456
rect 3415 20404 3428 20456
rect 3480 20404 3493 20456
rect 3545 20404 3558 20456
rect 3610 20404 3623 20456
rect 3675 20404 3688 20456
rect 3740 20404 3753 20456
rect 3805 20404 3818 20456
rect 3870 20404 3883 20456
rect 3935 20404 3948 20456
rect 4000 20404 4013 20456
rect 4065 20404 4078 20456
rect 4130 20404 4143 20456
rect 4195 20404 4208 20456
rect 4260 20404 4273 20456
rect 4325 20404 4338 20456
rect 4390 20404 4403 20456
rect 4455 20404 4468 20456
rect 4520 20404 4532 20456
rect 4584 20444 5613 20456
rect 5669 20444 5696 20461
rect 4584 20404 5040 20444
rect 2444 20396 5040 20404
rect 2270 20392 5040 20396
rect 5092 20392 5106 20444
rect 5158 20392 5594 20444
rect 5752 20428 5779 20484
rect 5835 20428 5861 20484
rect 5917 20428 5943 20484
rect 5999 20428 6025 20484
rect 6081 20428 6107 20484
rect 6266 20461 6271 20484
rect 6163 20444 6189 20461
rect 6245 20444 6271 20461
rect 6266 20428 6271 20444
rect 6327 20428 6353 20484
rect 6409 20428 6435 20484
rect 6491 20428 6517 20484
rect 6573 20428 6599 20484
rect 6655 20428 6681 20484
rect 6754 20461 6763 20484
rect 6820 20461 6845 20484
rect 6737 20444 6763 20461
rect 6819 20444 6845 20461
rect 6754 20428 6763 20444
rect 6820 20428 6845 20444
rect 6901 20428 6927 20484
rect 6983 20428 7009 20484
rect 7065 20428 7091 20484
rect 7147 20428 7173 20484
rect 7229 20428 7255 20484
rect 7311 20461 7322 20484
rect 7311 20444 7337 20461
rect 7311 20428 7322 20444
rect 7393 20428 7419 20484
rect 7475 20428 7501 20484
rect 7557 20428 7583 20484
rect 7639 20428 7665 20484
rect 7721 20428 7747 20484
rect 7803 20461 7810 20484
rect 7803 20444 7829 20461
rect 7885 20444 7911 20461
rect 7803 20428 7810 20444
rect 7967 20428 7993 20484
rect 8049 20448 8075 20465
rect 8131 20428 8157 20484
rect 8221 20465 8222 20517
rect 8213 20448 8222 20465
rect 5646 20404 5660 20428
rect 5712 20404 6148 20428
rect 6200 20404 6214 20428
rect 6266 20404 6702 20428
rect 6754 20404 6768 20428
rect 6820 20404 7256 20428
rect 7308 20404 7322 20428
rect 7374 20404 7810 20428
rect 7862 20404 7876 20428
rect 7928 20404 8047 20428
rect 8099 20404 8169 20428
rect 2270 20388 5613 20392
rect 2270 20378 2648 20388
rect 2322 20326 2392 20378
rect 2444 20336 2648 20378
rect 2700 20336 2713 20388
rect 2765 20336 2778 20388
rect 2830 20336 2843 20388
rect 2895 20336 2908 20388
rect 2960 20336 2973 20388
rect 3025 20336 3038 20388
rect 3090 20336 3103 20388
rect 3155 20336 3168 20388
rect 3220 20336 3233 20388
rect 3285 20336 3298 20388
rect 3350 20336 3363 20388
rect 3415 20336 3428 20388
rect 3480 20336 3493 20388
rect 3545 20336 3558 20388
rect 3610 20336 3623 20388
rect 3675 20336 3688 20388
rect 3740 20336 3753 20388
rect 3805 20336 3818 20388
rect 3870 20336 3883 20388
rect 3935 20336 3948 20388
rect 4000 20336 4013 20388
rect 4065 20336 4078 20388
rect 4130 20336 4143 20388
rect 4195 20336 4208 20388
rect 4260 20336 4273 20388
rect 4325 20336 4338 20388
rect 4390 20336 4403 20388
rect 4455 20336 4468 20388
rect 4520 20336 4532 20388
rect 4584 20375 5613 20388
rect 5669 20375 5696 20392
rect 4584 20336 5040 20375
rect 2444 20326 5040 20336
rect 2270 20323 5040 20326
rect 5092 20323 5106 20375
rect 5158 20323 5594 20375
rect 5752 20348 5779 20404
rect 5835 20348 5861 20404
rect 5917 20348 5943 20404
rect 5999 20348 6025 20404
rect 6081 20348 6107 20404
rect 6266 20392 6271 20404
rect 6163 20375 6189 20392
rect 6245 20375 6271 20392
rect 6266 20348 6271 20375
rect 6327 20348 6353 20404
rect 6409 20348 6435 20404
rect 6491 20348 6517 20404
rect 6573 20348 6599 20404
rect 6655 20348 6681 20404
rect 6754 20392 6763 20404
rect 6820 20392 6845 20404
rect 6737 20375 6763 20392
rect 6819 20375 6845 20392
rect 6754 20348 6763 20375
rect 6820 20348 6845 20375
rect 6901 20348 6927 20404
rect 6983 20348 7009 20404
rect 7065 20348 7091 20404
rect 7147 20348 7173 20404
rect 7229 20348 7255 20404
rect 7311 20392 7322 20404
rect 7311 20375 7337 20392
rect 7311 20348 7322 20375
rect 7393 20348 7419 20404
rect 7475 20348 7501 20404
rect 7557 20348 7583 20404
rect 7639 20348 7665 20404
rect 7721 20348 7747 20404
rect 7803 20392 7810 20404
rect 7803 20375 7829 20392
rect 7885 20375 7911 20392
rect 7803 20348 7810 20375
rect 7967 20348 7993 20404
rect 8049 20378 8075 20396
rect 8131 20348 8157 20404
rect 8221 20396 8222 20448
rect 8213 20378 8222 20396
rect 5646 20324 5660 20348
rect 5712 20324 6148 20348
rect 6200 20324 6214 20348
rect 6266 20324 6702 20348
rect 6754 20324 6768 20348
rect 6820 20324 7256 20348
rect 7308 20324 7322 20348
rect 7374 20324 7810 20348
rect 7862 20324 7876 20348
rect 7928 20326 8047 20348
rect 8099 20326 8169 20348
rect 8221 20326 8222 20378
rect 7928 20324 8222 20326
rect 2270 20320 5613 20323
rect 2270 20308 2648 20320
rect 2322 20256 2392 20308
rect 2444 20268 2648 20308
rect 2700 20268 2713 20320
rect 2765 20268 2778 20320
rect 2830 20268 2843 20320
rect 2895 20268 2908 20320
rect 2960 20268 2973 20320
rect 3025 20268 3038 20320
rect 3090 20268 3103 20320
rect 3155 20268 3168 20320
rect 3220 20268 3233 20320
rect 3285 20268 3298 20320
rect 3350 20268 3363 20320
rect 3415 20268 3428 20320
rect 3480 20268 3493 20320
rect 3545 20268 3558 20320
rect 3610 20268 3623 20320
rect 3675 20268 3688 20320
rect 3740 20268 3753 20320
rect 3805 20268 3818 20320
rect 3870 20268 3883 20320
rect 3935 20268 3948 20320
rect 4000 20268 4013 20320
rect 4065 20268 4078 20320
rect 4130 20268 4143 20320
rect 4195 20268 4208 20320
rect 4260 20268 4273 20320
rect 4325 20268 4338 20320
rect 4390 20268 4403 20320
rect 4455 20268 4468 20320
rect 4520 20268 4532 20320
rect 4584 20306 5613 20320
rect 5669 20306 5696 20323
rect 4584 20268 5040 20306
rect 2444 20256 5040 20268
rect 2270 20254 5040 20256
rect 5092 20254 5106 20306
rect 5158 20254 5594 20306
rect 5752 20268 5779 20324
rect 5835 20268 5861 20324
rect 5917 20268 5943 20324
rect 5999 20268 6025 20324
rect 6081 20268 6107 20324
rect 6266 20323 6271 20324
rect 6163 20306 6189 20323
rect 6245 20306 6271 20323
rect 6266 20268 6271 20306
rect 6327 20268 6353 20324
rect 6409 20268 6435 20324
rect 6491 20268 6517 20324
rect 6573 20268 6599 20324
rect 6655 20268 6681 20324
rect 6754 20323 6763 20324
rect 6820 20323 6845 20324
rect 6737 20306 6763 20323
rect 6819 20306 6845 20323
rect 6754 20268 6763 20306
rect 6820 20268 6845 20306
rect 6901 20268 6927 20324
rect 6983 20268 7009 20324
rect 7065 20268 7091 20324
rect 7147 20268 7173 20324
rect 7229 20268 7255 20324
rect 7311 20323 7322 20324
rect 7311 20306 7337 20323
rect 7311 20268 7322 20306
rect 7393 20268 7419 20324
rect 7475 20268 7501 20324
rect 7557 20268 7583 20324
rect 7639 20268 7665 20324
rect 7721 20268 7747 20324
rect 7803 20323 7810 20324
rect 7803 20306 7829 20323
rect 7885 20306 7911 20323
rect 7803 20268 7810 20306
rect 7967 20268 7993 20324
rect 8049 20308 8075 20324
rect 8131 20268 8157 20324
rect 8213 20308 8222 20324
rect 5646 20254 5660 20268
rect 5712 20254 6148 20268
rect 6200 20254 6214 20268
rect 6266 20254 6702 20268
rect 6754 20254 6768 20268
rect 6820 20254 7256 20268
rect 7308 20254 7322 20268
rect 7374 20254 7810 20268
rect 7862 20254 7876 20268
rect 7928 20256 8047 20268
rect 8099 20256 8169 20268
rect 8221 20256 8222 20308
rect 7928 20254 8222 20256
rect 2270 20252 8222 20254
rect 2270 20238 2648 20252
rect 2322 20186 2392 20238
rect 2444 20200 2648 20238
rect 2700 20200 2713 20252
rect 2765 20200 2778 20252
rect 2830 20200 2843 20252
rect 2895 20200 2908 20252
rect 2960 20200 2973 20252
rect 3025 20200 3038 20252
rect 3090 20200 3103 20252
rect 3155 20200 3168 20252
rect 3220 20200 3233 20252
rect 3285 20200 3298 20252
rect 3350 20200 3363 20252
rect 3415 20200 3428 20252
rect 3480 20200 3493 20252
rect 3545 20200 3558 20252
rect 3610 20200 3623 20252
rect 3675 20200 3688 20252
rect 3740 20200 3753 20252
rect 3805 20200 3818 20252
rect 3870 20200 3883 20252
rect 3935 20200 3948 20252
rect 4000 20200 4013 20252
rect 4065 20200 4078 20252
rect 4130 20200 4143 20252
rect 4195 20200 4208 20252
rect 4260 20200 4273 20252
rect 4325 20200 4338 20252
rect 4390 20200 4403 20252
rect 4455 20200 4468 20252
rect 4520 20200 4532 20252
rect 4584 20244 8222 20252
rect 4584 20236 5613 20244
rect 5669 20236 5696 20244
rect 4584 20200 5040 20236
rect 2444 20186 5040 20200
rect 2270 20184 5040 20186
rect 5092 20184 5106 20236
rect 5158 20184 5594 20236
rect 5752 20188 5779 20244
rect 5835 20188 5861 20244
rect 5917 20188 5943 20244
rect 5999 20188 6025 20244
rect 6081 20188 6107 20244
rect 6163 20236 6189 20244
rect 6245 20236 6271 20244
rect 6266 20188 6271 20236
rect 6327 20188 6353 20244
rect 6409 20188 6435 20244
rect 6491 20188 6517 20244
rect 6573 20188 6599 20244
rect 6655 20188 6681 20244
rect 6737 20236 6763 20244
rect 6819 20236 6845 20244
rect 6754 20188 6763 20236
rect 6820 20188 6845 20236
rect 6901 20188 6927 20244
rect 6983 20188 7009 20244
rect 7065 20188 7091 20244
rect 7147 20188 7173 20244
rect 7229 20188 7255 20244
rect 7311 20236 7337 20244
rect 7311 20188 7322 20236
rect 7393 20188 7419 20244
rect 7475 20188 7501 20244
rect 7557 20188 7583 20244
rect 7639 20188 7665 20244
rect 7721 20188 7747 20244
rect 7803 20236 7829 20244
rect 7885 20236 7911 20244
rect 7803 20188 7810 20236
rect 7967 20188 7993 20244
rect 8049 20238 8075 20244
rect 8131 20188 8157 20244
rect 8213 20238 8222 20244
rect 5646 20184 5660 20188
rect 5712 20184 6148 20188
rect 6200 20184 6214 20188
rect 6266 20184 6702 20188
rect 6754 20184 6768 20188
rect 6820 20184 7256 20188
rect 7308 20184 7322 20188
rect 7374 20184 7810 20188
rect 7862 20184 7876 20188
rect 7928 20186 8047 20188
rect 8099 20186 8169 20188
rect 8221 20186 8222 20238
rect 7928 20184 8222 20186
rect 2270 20168 8222 20184
rect 2322 20116 2392 20168
rect 2444 20166 8047 20168
rect 2444 20116 5040 20166
rect 2270 20114 5040 20116
rect 5092 20114 5106 20166
rect 5158 20114 5594 20166
rect 5646 20164 5660 20166
rect 5712 20164 6148 20166
rect 6200 20164 6214 20166
rect 6266 20164 6702 20166
rect 6754 20164 6768 20166
rect 6820 20164 7256 20166
rect 7308 20164 7322 20166
rect 7374 20164 7810 20166
rect 7862 20164 7876 20166
rect 7928 20164 8047 20166
rect 8099 20164 8169 20168
rect 2270 20108 5613 20114
rect 5669 20108 5696 20114
rect 5752 20108 5779 20164
rect 5835 20108 5861 20164
rect 5917 20108 5943 20164
rect 5999 20108 6025 20164
rect 6081 20108 6107 20164
rect 6266 20114 6271 20164
rect 6163 20108 6189 20114
rect 6245 20108 6271 20114
rect 6327 20108 6353 20164
rect 6409 20108 6435 20164
rect 6491 20108 6517 20164
rect 6573 20108 6599 20164
rect 6655 20108 6681 20164
rect 6754 20114 6763 20164
rect 6820 20114 6845 20164
rect 6737 20108 6763 20114
rect 6819 20108 6845 20114
rect 6901 20108 6927 20164
rect 6983 20108 7009 20164
rect 7065 20108 7091 20164
rect 7147 20108 7173 20164
rect 7229 20108 7255 20164
rect 7311 20114 7322 20164
rect 7311 20108 7337 20114
rect 7393 20108 7419 20164
rect 7475 20108 7501 20164
rect 7557 20108 7583 20164
rect 7639 20108 7665 20164
rect 7721 20108 7747 20164
rect 7803 20114 7810 20164
rect 7803 20108 7829 20114
rect 7885 20108 7911 20114
rect 7967 20108 7993 20164
rect 8049 20108 8075 20116
rect 8131 20108 8157 20164
rect 8221 20116 8222 20168
rect 8213 20108 8222 20116
rect 2724 19987 7651 19988
rect 2724 19931 2733 19987
rect 2789 19931 2814 19987
rect 2870 19931 2895 19987
rect 2951 19931 2976 19987
rect 3032 19931 3057 19987
rect 3113 19931 3138 19987
rect 3194 19931 3219 19987
rect 3275 19931 3300 19987
rect 3356 19931 3381 19987
rect 3437 19931 3462 19987
rect 3518 19931 3543 19987
rect 3599 19931 3624 19987
rect 3680 19931 3705 19987
rect 3761 19931 3786 19987
rect 3842 19931 3867 19987
rect 3923 19931 3948 19987
rect 4004 19931 4029 19987
rect 4085 19931 4110 19987
rect 4166 19931 4191 19987
rect 4247 19931 4272 19987
rect 4328 19931 4353 19987
rect 4409 19931 4434 19987
rect 4490 19931 4515 19987
rect 4571 19931 4596 19987
rect 4652 19931 4677 19987
rect 4733 19931 4758 19987
rect 4814 19931 4839 19987
rect 4895 19931 4920 19987
rect 4976 19931 5001 19987
rect 5057 19931 5082 19987
rect 5138 19931 5163 19987
rect 2724 19907 5163 19931
rect 2724 19851 2733 19907
rect 2789 19851 2814 19907
rect 2870 19851 2895 19907
rect 2951 19851 2976 19907
rect 3032 19851 3057 19907
rect 3113 19851 3138 19907
rect 3194 19851 3219 19907
rect 3275 19851 3300 19907
rect 3356 19851 3381 19907
rect 3437 19851 3462 19907
rect 3518 19851 3543 19907
rect 3599 19851 3624 19907
rect 3680 19851 3705 19907
rect 3761 19851 3786 19907
rect 3842 19851 3867 19907
rect 3923 19851 3948 19907
rect 4004 19851 4029 19907
rect 4085 19851 4110 19907
rect 4166 19851 4191 19907
rect 4247 19851 4272 19907
rect 4328 19851 4353 19907
rect 4409 19851 4434 19907
rect 4490 19851 4515 19907
rect 4571 19851 4596 19907
rect 4652 19851 4677 19907
rect 4733 19851 4758 19907
rect 4814 19851 4839 19907
rect 4895 19851 4920 19907
rect 4976 19851 5001 19907
rect 5057 19851 5082 19907
rect 5138 19851 5163 19907
rect 2724 19827 5163 19851
rect 2724 19771 2733 19827
rect 2789 19771 2814 19827
rect 2870 19771 2895 19827
rect 2951 19771 2976 19827
rect 3032 19771 3057 19827
rect 3113 19771 3138 19827
rect 3194 19771 3219 19827
rect 3275 19771 3300 19827
rect 3356 19771 3381 19827
rect 3437 19771 3462 19827
rect 3518 19771 3543 19827
rect 3599 19771 3624 19827
rect 3680 19771 3705 19827
rect 3761 19771 3786 19827
rect 3842 19771 3867 19827
rect 3923 19771 3948 19827
rect 4004 19771 4029 19827
rect 4085 19771 4110 19827
rect 4166 19771 4191 19827
rect 4247 19771 4272 19827
rect 4328 19771 4353 19827
rect 4409 19771 4434 19827
rect 4490 19771 4515 19827
rect 4571 19771 4596 19827
rect 4652 19771 4677 19827
rect 4733 19771 4758 19827
rect 4814 19771 4839 19827
rect 4895 19771 4920 19827
rect 4976 19771 5001 19827
rect 5057 19771 5082 19827
rect 5138 19771 5163 19827
rect 2724 19747 5163 19771
rect 2724 19691 2733 19747
rect 2789 19691 2814 19747
rect 2870 19691 2895 19747
rect 2951 19691 2976 19747
rect 3032 19691 3057 19747
rect 3113 19691 3138 19747
rect 3194 19691 3219 19747
rect 3275 19691 3300 19747
rect 3356 19691 3381 19747
rect 3437 19691 3462 19747
rect 3518 19691 3543 19747
rect 3599 19691 3624 19747
rect 3680 19691 3705 19747
rect 3761 19691 3786 19747
rect 3842 19691 3867 19747
rect 3923 19691 3948 19747
rect 4004 19691 4029 19747
rect 4085 19691 4110 19747
rect 4166 19691 4191 19747
rect 4247 19691 4272 19747
rect 4328 19691 4353 19747
rect 4409 19691 4434 19747
rect 4490 19691 4515 19747
rect 4571 19691 4596 19747
rect 4652 19691 4677 19747
rect 4733 19691 4758 19747
rect 4814 19691 4839 19747
rect 4895 19691 4920 19747
rect 4976 19691 5001 19747
rect 5057 19691 5082 19747
rect 5138 19691 5163 19747
rect 2724 19667 5163 19691
rect 2724 19611 2733 19667
rect 2789 19611 2814 19667
rect 2870 19611 2895 19667
rect 2951 19611 2976 19667
rect 3032 19611 3057 19667
rect 3113 19611 3138 19667
rect 3194 19611 3219 19667
rect 3275 19611 3300 19667
rect 3356 19611 3381 19667
rect 3437 19611 3462 19667
rect 3518 19611 3543 19667
rect 3599 19611 3624 19667
rect 3680 19611 3705 19667
rect 3761 19611 3786 19667
rect 3842 19611 3867 19667
rect 3923 19611 3948 19667
rect 4004 19611 4029 19667
rect 4085 19611 4110 19667
rect 4166 19611 4191 19667
rect 4247 19611 4272 19667
rect 4328 19611 4353 19667
rect 4409 19611 4434 19667
rect 4490 19611 4515 19667
rect 4571 19611 4596 19667
rect 4652 19611 4677 19667
rect 4733 19611 4758 19667
rect 4814 19611 4839 19667
rect 4895 19611 4920 19667
rect 4976 19611 5001 19667
rect 5057 19611 5082 19667
rect 5138 19611 5163 19667
rect 2724 19587 5163 19611
rect 2724 19531 2733 19587
rect 2789 19531 2814 19587
rect 2870 19531 2895 19587
rect 2951 19531 2976 19587
rect 3032 19531 3057 19587
rect 3113 19531 3138 19587
rect 3194 19531 3219 19587
rect 3275 19531 3300 19587
rect 3356 19531 3381 19587
rect 3437 19531 3462 19587
rect 3518 19531 3543 19587
rect 3599 19531 3624 19587
rect 3680 19531 3705 19587
rect 3761 19531 3786 19587
rect 3842 19531 3867 19587
rect 3923 19531 3948 19587
rect 4004 19531 4029 19587
rect 4085 19531 4110 19587
rect 4166 19531 4191 19587
rect 4247 19531 4272 19587
rect 4328 19531 4353 19587
rect 4409 19531 4434 19587
rect 4490 19531 4515 19587
rect 4571 19531 4596 19587
rect 4652 19531 4677 19587
rect 4733 19531 4758 19587
rect 4814 19531 4839 19587
rect 4895 19531 4920 19587
rect 4976 19531 5001 19587
rect 5057 19531 5082 19587
rect 5138 19531 5163 19587
rect 2724 19507 5163 19531
rect 2724 19451 2733 19507
rect 2789 19451 2814 19507
rect 2870 19451 2895 19507
rect 2951 19451 2976 19507
rect 3032 19451 3057 19507
rect 3113 19451 3138 19507
rect 3194 19451 3219 19507
rect 3275 19451 3300 19507
rect 3356 19451 3381 19507
rect 3437 19451 3462 19507
rect 3518 19451 3543 19507
rect 3599 19451 3624 19507
rect 3680 19451 3705 19507
rect 3761 19451 3786 19507
rect 3842 19451 3867 19507
rect 3923 19451 3948 19507
rect 4004 19451 4029 19507
rect 4085 19451 4110 19507
rect 4166 19451 4191 19507
rect 4247 19451 4272 19507
rect 4328 19451 4353 19507
rect 4409 19451 4434 19507
rect 4490 19451 4515 19507
rect 4571 19451 4596 19507
rect 4652 19451 4677 19507
rect 4733 19451 4758 19507
rect 4814 19451 4839 19507
rect 4895 19451 4920 19507
rect 4976 19451 5001 19507
rect 5057 19451 5082 19507
rect 5138 19451 5163 19507
rect 2724 19427 5163 19451
rect 2724 19371 2733 19427
rect 2789 19371 2814 19427
rect 2870 19371 2895 19427
rect 2951 19371 2976 19427
rect 3032 19371 3057 19427
rect 3113 19371 3138 19427
rect 3194 19371 3219 19427
rect 3275 19371 3300 19427
rect 3356 19371 3381 19427
rect 3437 19371 3462 19427
rect 3518 19371 3543 19427
rect 3599 19371 3624 19427
rect 3680 19371 3705 19427
rect 3761 19371 3786 19427
rect 3842 19371 3867 19427
rect 3923 19371 3948 19427
rect 4004 19371 4029 19427
rect 4085 19371 4110 19427
rect 4166 19371 4191 19427
rect 4247 19371 4272 19427
rect 4328 19371 4353 19427
rect 4409 19371 4434 19427
rect 4490 19371 4515 19427
rect 4571 19371 4596 19427
rect 4652 19371 4677 19427
rect 4733 19371 4758 19427
rect 4814 19371 4839 19427
rect 4895 19371 4920 19427
rect 4976 19371 5001 19427
rect 5057 19371 5082 19427
rect 5138 19371 5163 19427
rect 5299 19982 7651 19987
rect 5299 19930 5317 19982
rect 5369 19930 5383 19982
rect 5435 19930 5871 19982
rect 5923 19930 5937 19982
rect 5989 19930 6425 19982
rect 6477 19930 6491 19982
rect 6543 19930 6979 19982
rect 7031 19930 7045 19982
rect 7097 19930 7533 19982
rect 7585 19930 7599 19982
rect 5299 19913 7651 19930
rect 5299 19861 5317 19913
rect 5369 19861 5383 19913
rect 5435 19861 5871 19913
rect 5923 19861 5937 19913
rect 5989 19861 6425 19913
rect 6477 19861 6491 19913
rect 6543 19861 6979 19913
rect 7031 19861 7045 19913
rect 7097 19861 7533 19913
rect 7585 19861 7599 19913
rect 5299 19844 7651 19861
rect 5299 19792 5317 19844
rect 5369 19792 5383 19844
rect 5435 19792 5871 19844
rect 5923 19792 5937 19844
rect 5989 19792 6425 19844
rect 6477 19792 6491 19844
rect 6543 19792 6979 19844
rect 7031 19792 7045 19844
rect 7097 19792 7533 19844
rect 7585 19792 7599 19844
rect 5299 19775 7651 19792
rect 5299 19723 5317 19775
rect 5369 19723 5383 19775
rect 5435 19723 5871 19775
rect 5923 19723 5937 19775
rect 5989 19723 6425 19775
rect 6477 19723 6491 19775
rect 6543 19723 6979 19775
rect 7031 19723 7045 19775
rect 7097 19723 7533 19775
rect 7585 19723 7599 19775
rect 5299 19706 7651 19723
rect 5299 19654 5317 19706
rect 5369 19654 5383 19706
rect 5435 19654 5871 19706
rect 5923 19654 5937 19706
rect 5989 19654 6425 19706
rect 6477 19654 6491 19706
rect 6543 19654 6979 19706
rect 7031 19654 7045 19706
rect 7097 19654 7533 19706
rect 7585 19654 7599 19706
rect 5299 19636 7651 19654
rect 5299 19584 5317 19636
rect 5369 19584 5383 19636
rect 5435 19584 5871 19636
rect 5923 19584 5937 19636
rect 5989 19584 6425 19636
rect 6477 19584 6491 19636
rect 6543 19584 6979 19636
rect 7031 19584 7045 19636
rect 7097 19584 7533 19636
rect 7585 19584 7599 19636
rect 5299 19566 7651 19584
rect 5299 19514 5317 19566
rect 5369 19514 5383 19566
rect 5435 19514 5871 19566
rect 5923 19514 5937 19566
rect 5989 19514 6425 19566
rect 6477 19514 6491 19566
rect 6543 19514 6979 19566
rect 7031 19514 7045 19566
rect 7097 19514 7533 19566
rect 7585 19514 7599 19566
rect 5299 19496 7651 19514
rect 5299 19444 5317 19496
rect 5369 19444 5383 19496
rect 5435 19444 5871 19496
rect 5923 19444 5937 19496
rect 5989 19444 6425 19496
rect 6477 19444 6491 19496
rect 6543 19444 6979 19496
rect 7031 19444 7045 19496
rect 7097 19444 7533 19496
rect 7585 19444 7599 19496
rect 5299 19426 7651 19444
rect 5299 19374 5317 19426
rect 5369 19374 5383 19426
rect 5435 19374 5871 19426
rect 5923 19374 5937 19426
rect 5989 19374 6425 19426
rect 6477 19374 6491 19426
rect 6543 19374 6979 19426
rect 7031 19374 7045 19426
rect 7097 19374 7533 19426
rect 7585 19374 7599 19426
rect 5299 19371 7651 19374
rect 2724 19368 7651 19371
rect 2270 18728 8222 18730
rect 2270 18724 2648 18728
rect 2322 18672 2392 18724
rect 2444 18676 2648 18724
rect 2700 18676 2713 18728
rect 2765 18676 2778 18728
rect 2830 18676 2843 18728
rect 2895 18676 2908 18728
rect 2960 18676 2973 18728
rect 3025 18676 3038 18728
rect 3090 18676 3103 18728
rect 3155 18676 3168 18728
rect 3220 18676 3233 18728
rect 3285 18676 3298 18728
rect 3350 18676 3363 18728
rect 3415 18676 3428 18728
rect 3480 18676 3493 18728
rect 3545 18676 3558 18728
rect 3610 18676 3623 18728
rect 3675 18676 3688 18728
rect 3740 18676 3753 18728
rect 3805 18676 3818 18728
rect 3870 18676 3883 18728
rect 3935 18676 3948 18728
rect 4000 18676 4013 18728
rect 4065 18676 4078 18728
rect 4130 18676 4143 18728
rect 4195 18676 4208 18728
rect 4260 18676 4273 18728
rect 4325 18676 4338 18728
rect 4390 18676 4403 18728
rect 4455 18676 4468 18728
rect 4520 18676 4532 18728
rect 4584 18724 8222 18728
rect 4584 18720 5613 18724
rect 5669 18720 5696 18724
rect 4584 18676 5040 18720
rect 2444 18672 5040 18676
rect 2270 18668 5040 18672
rect 5092 18668 5106 18720
rect 5158 18668 5594 18720
rect 5752 18668 5779 18724
rect 5835 18668 5861 18724
rect 5917 18668 5943 18724
rect 5999 18668 6025 18724
rect 6081 18668 6107 18724
rect 6163 18720 6189 18724
rect 6245 18720 6271 18724
rect 6266 18668 6271 18720
rect 6327 18668 6353 18724
rect 6409 18668 6435 18724
rect 6491 18668 6517 18724
rect 6573 18668 6599 18724
rect 6655 18668 6681 18724
rect 6737 18720 6763 18724
rect 6819 18720 6845 18724
rect 6754 18668 6763 18720
rect 6820 18668 6845 18720
rect 6901 18668 6927 18724
rect 6983 18668 7009 18724
rect 7065 18668 7091 18724
rect 7147 18668 7173 18724
rect 7229 18668 7255 18724
rect 7311 18720 7337 18724
rect 7311 18668 7322 18720
rect 7393 18668 7419 18724
rect 7475 18668 7501 18724
rect 7557 18668 7583 18724
rect 7639 18668 7665 18724
rect 7721 18668 7747 18724
rect 7803 18720 7829 18724
rect 7885 18720 7911 18724
rect 7803 18668 7810 18720
rect 7967 18668 7993 18724
rect 8049 18668 8075 18672
rect 8131 18668 8157 18724
rect 8221 18672 8222 18724
rect 8213 18668 8222 18672
rect 2270 18660 8222 18668
rect 2270 18655 2648 18660
rect 2322 18603 2392 18655
rect 2444 18608 2648 18655
rect 2700 18608 2713 18660
rect 2765 18608 2778 18660
rect 2830 18608 2843 18660
rect 2895 18608 2908 18660
rect 2960 18608 2973 18660
rect 3025 18608 3038 18660
rect 3090 18608 3103 18660
rect 3155 18608 3168 18660
rect 3220 18608 3233 18660
rect 3285 18608 3298 18660
rect 3350 18608 3363 18660
rect 3415 18608 3428 18660
rect 3480 18608 3493 18660
rect 3545 18608 3558 18660
rect 3610 18608 3623 18660
rect 3675 18608 3688 18660
rect 3740 18608 3753 18660
rect 3805 18608 3818 18660
rect 3870 18608 3883 18660
rect 3935 18608 3948 18660
rect 4000 18608 4013 18660
rect 4065 18608 4078 18660
rect 4130 18608 4143 18660
rect 4195 18608 4208 18660
rect 4260 18608 4273 18660
rect 4325 18608 4338 18660
rect 4390 18608 4403 18660
rect 4455 18608 4468 18660
rect 4520 18608 4532 18660
rect 4584 18655 8222 18660
rect 4584 18651 8047 18655
rect 4584 18608 5040 18651
rect 2444 18603 5040 18608
rect 2270 18599 5040 18603
rect 5092 18599 5106 18651
rect 5158 18599 5594 18651
rect 5646 18644 5660 18651
rect 5712 18644 6148 18651
rect 6200 18644 6214 18651
rect 6266 18644 6702 18651
rect 6754 18644 6768 18651
rect 6820 18644 7256 18651
rect 7308 18644 7322 18651
rect 7374 18644 7810 18651
rect 7862 18644 7876 18651
rect 7928 18644 8047 18651
rect 8099 18644 8169 18655
rect 2270 18592 5613 18599
rect 2270 18586 2648 18592
rect 2322 18534 2392 18586
rect 2444 18540 2648 18586
rect 2700 18540 2713 18592
rect 2765 18540 2778 18592
rect 2830 18540 2843 18592
rect 2895 18540 2908 18592
rect 2960 18540 2973 18592
rect 3025 18540 3038 18592
rect 3090 18540 3103 18592
rect 3155 18540 3168 18592
rect 3220 18540 3233 18592
rect 3285 18540 3298 18592
rect 3350 18540 3363 18592
rect 3415 18540 3428 18592
rect 3480 18540 3493 18592
rect 3545 18540 3558 18592
rect 3610 18540 3623 18592
rect 3675 18540 3688 18592
rect 3740 18540 3753 18592
rect 3805 18540 3818 18592
rect 3870 18540 3883 18592
rect 3935 18540 3948 18592
rect 4000 18540 4013 18592
rect 4065 18540 4078 18592
rect 4130 18540 4143 18592
rect 4195 18540 4208 18592
rect 4260 18540 4273 18592
rect 4325 18540 4338 18592
rect 4390 18540 4403 18592
rect 4455 18540 4468 18592
rect 4520 18540 4532 18592
rect 4584 18588 5613 18592
rect 5669 18588 5696 18599
rect 5752 18588 5779 18644
rect 5835 18588 5861 18644
rect 5917 18588 5943 18644
rect 5999 18588 6025 18644
rect 6081 18588 6107 18644
rect 6266 18599 6271 18644
rect 6163 18588 6189 18599
rect 6245 18588 6271 18599
rect 6327 18588 6353 18644
rect 6409 18588 6435 18644
rect 6491 18588 6517 18644
rect 6573 18588 6599 18644
rect 6655 18588 6681 18644
rect 6754 18599 6763 18644
rect 6820 18599 6845 18644
rect 6737 18588 6763 18599
rect 6819 18588 6845 18599
rect 6901 18588 6927 18644
rect 6983 18588 7009 18644
rect 7065 18588 7091 18644
rect 7147 18588 7173 18644
rect 7229 18588 7255 18644
rect 7311 18599 7322 18644
rect 7311 18588 7337 18599
rect 7393 18588 7419 18644
rect 7475 18588 7501 18644
rect 7557 18588 7583 18644
rect 7639 18588 7665 18644
rect 7721 18588 7747 18644
rect 7803 18599 7810 18644
rect 7803 18588 7829 18599
rect 7885 18588 7911 18599
rect 7967 18588 7993 18644
rect 8049 18588 8075 18603
rect 8131 18588 8157 18644
rect 8221 18603 8222 18655
rect 8213 18588 8222 18603
rect 4584 18586 8222 18588
rect 4584 18582 8047 18586
rect 4584 18540 5040 18582
rect 2444 18534 5040 18540
rect 2270 18530 5040 18534
rect 5092 18530 5106 18582
rect 5158 18530 5594 18582
rect 5646 18564 5660 18582
rect 5712 18564 6148 18582
rect 6200 18564 6214 18582
rect 6266 18564 6702 18582
rect 6754 18564 6768 18582
rect 6820 18564 7256 18582
rect 7308 18564 7322 18582
rect 7374 18564 7810 18582
rect 7862 18564 7876 18582
rect 7928 18564 8047 18582
rect 8099 18564 8169 18586
rect 2270 18524 5613 18530
rect 2270 18517 2648 18524
rect 2322 18465 2392 18517
rect 2444 18472 2648 18517
rect 2700 18472 2713 18524
rect 2765 18472 2778 18524
rect 2830 18472 2843 18524
rect 2895 18472 2908 18524
rect 2960 18472 2973 18524
rect 3025 18472 3038 18524
rect 3090 18472 3103 18524
rect 3155 18472 3168 18524
rect 3220 18472 3233 18524
rect 3285 18472 3298 18524
rect 3350 18472 3363 18524
rect 3415 18472 3428 18524
rect 3480 18472 3493 18524
rect 3545 18472 3558 18524
rect 3610 18472 3623 18524
rect 3675 18472 3688 18524
rect 3740 18472 3753 18524
rect 3805 18472 3818 18524
rect 3870 18472 3883 18524
rect 3935 18472 3948 18524
rect 4000 18472 4013 18524
rect 4065 18472 4078 18524
rect 4130 18472 4143 18524
rect 4195 18472 4208 18524
rect 4260 18472 4273 18524
rect 4325 18472 4338 18524
rect 4390 18472 4403 18524
rect 4455 18472 4468 18524
rect 4520 18472 4532 18524
rect 4584 18513 5613 18524
rect 5669 18513 5696 18530
rect 4584 18472 5040 18513
rect 2444 18465 5040 18472
rect 2270 18461 5040 18465
rect 5092 18461 5106 18513
rect 5158 18461 5594 18513
rect 5752 18508 5779 18564
rect 5835 18508 5861 18564
rect 5917 18508 5943 18564
rect 5999 18508 6025 18564
rect 6081 18508 6107 18564
rect 6266 18530 6271 18564
rect 6163 18513 6189 18530
rect 6245 18513 6271 18530
rect 6266 18508 6271 18513
rect 6327 18508 6353 18564
rect 6409 18508 6435 18564
rect 6491 18508 6517 18564
rect 6573 18508 6599 18564
rect 6655 18508 6681 18564
rect 6754 18530 6763 18564
rect 6820 18530 6845 18564
rect 6737 18513 6763 18530
rect 6819 18513 6845 18530
rect 6754 18508 6763 18513
rect 6820 18508 6845 18513
rect 6901 18508 6927 18564
rect 6983 18508 7009 18564
rect 7065 18508 7091 18564
rect 7147 18508 7173 18564
rect 7229 18508 7255 18564
rect 7311 18530 7322 18564
rect 7311 18513 7337 18530
rect 7311 18508 7322 18513
rect 7393 18508 7419 18564
rect 7475 18508 7501 18564
rect 7557 18508 7583 18564
rect 7639 18508 7665 18564
rect 7721 18508 7747 18564
rect 7803 18530 7810 18564
rect 7803 18513 7829 18530
rect 7885 18513 7911 18530
rect 7803 18508 7810 18513
rect 7967 18508 7993 18564
rect 8049 18517 8075 18534
rect 8131 18508 8157 18564
rect 8221 18534 8222 18586
rect 8213 18517 8222 18534
rect 5646 18484 5660 18508
rect 5712 18484 6148 18508
rect 6200 18484 6214 18508
rect 6266 18484 6702 18508
rect 6754 18484 6768 18508
rect 6820 18484 7256 18508
rect 7308 18484 7322 18508
rect 7374 18484 7810 18508
rect 7862 18484 7876 18508
rect 7928 18484 8047 18508
rect 8099 18484 8169 18508
rect 2270 18456 5613 18461
rect 2270 18448 2648 18456
rect 2322 18396 2392 18448
rect 2444 18404 2648 18448
rect 2700 18404 2713 18456
rect 2765 18404 2778 18456
rect 2830 18404 2843 18456
rect 2895 18404 2908 18456
rect 2960 18404 2973 18456
rect 3025 18404 3038 18456
rect 3090 18404 3103 18456
rect 3155 18404 3168 18456
rect 3220 18404 3233 18456
rect 3285 18404 3298 18456
rect 3350 18404 3363 18456
rect 3415 18404 3428 18456
rect 3480 18404 3493 18456
rect 3545 18404 3558 18456
rect 3610 18404 3623 18456
rect 3675 18404 3688 18456
rect 3740 18404 3753 18456
rect 3805 18404 3818 18456
rect 3870 18404 3883 18456
rect 3935 18404 3948 18456
rect 4000 18404 4013 18456
rect 4065 18404 4078 18456
rect 4130 18404 4143 18456
rect 4195 18404 4208 18456
rect 4260 18404 4273 18456
rect 4325 18404 4338 18456
rect 4390 18404 4403 18456
rect 4455 18404 4468 18456
rect 4520 18404 4532 18456
rect 4584 18444 5613 18456
rect 5669 18444 5696 18461
rect 4584 18404 5040 18444
rect 2444 18396 5040 18404
rect 2270 18392 5040 18396
rect 5092 18392 5106 18444
rect 5158 18392 5594 18444
rect 5752 18428 5779 18484
rect 5835 18428 5861 18484
rect 5917 18428 5943 18484
rect 5999 18428 6025 18484
rect 6081 18428 6107 18484
rect 6266 18461 6271 18484
rect 6163 18444 6189 18461
rect 6245 18444 6271 18461
rect 6266 18428 6271 18444
rect 6327 18428 6353 18484
rect 6409 18428 6435 18484
rect 6491 18428 6517 18484
rect 6573 18428 6599 18484
rect 6655 18428 6681 18484
rect 6754 18461 6763 18484
rect 6820 18461 6845 18484
rect 6737 18444 6763 18461
rect 6819 18444 6845 18461
rect 6754 18428 6763 18444
rect 6820 18428 6845 18444
rect 6901 18428 6927 18484
rect 6983 18428 7009 18484
rect 7065 18428 7091 18484
rect 7147 18428 7173 18484
rect 7229 18428 7255 18484
rect 7311 18461 7322 18484
rect 7311 18444 7337 18461
rect 7311 18428 7322 18444
rect 7393 18428 7419 18484
rect 7475 18428 7501 18484
rect 7557 18428 7583 18484
rect 7639 18428 7665 18484
rect 7721 18428 7747 18484
rect 7803 18461 7810 18484
rect 7803 18444 7829 18461
rect 7885 18444 7911 18461
rect 7803 18428 7810 18444
rect 7967 18428 7993 18484
rect 8049 18448 8075 18465
rect 8131 18428 8157 18484
rect 8221 18465 8222 18517
rect 8213 18448 8222 18465
rect 5646 18404 5660 18428
rect 5712 18404 6148 18428
rect 6200 18404 6214 18428
rect 6266 18404 6702 18428
rect 6754 18404 6768 18428
rect 6820 18404 7256 18428
rect 7308 18404 7322 18428
rect 7374 18404 7810 18428
rect 7862 18404 7876 18428
rect 7928 18404 8047 18428
rect 8099 18404 8169 18428
rect 2270 18388 5613 18392
rect 2270 18378 2648 18388
rect 2322 18326 2392 18378
rect 2444 18336 2648 18378
rect 2700 18336 2713 18388
rect 2765 18336 2778 18388
rect 2830 18336 2843 18388
rect 2895 18336 2908 18388
rect 2960 18336 2973 18388
rect 3025 18336 3038 18388
rect 3090 18336 3103 18388
rect 3155 18336 3168 18388
rect 3220 18336 3233 18388
rect 3285 18336 3298 18388
rect 3350 18336 3363 18388
rect 3415 18336 3428 18388
rect 3480 18336 3493 18388
rect 3545 18336 3558 18388
rect 3610 18336 3623 18388
rect 3675 18336 3688 18388
rect 3740 18336 3753 18388
rect 3805 18336 3818 18388
rect 3870 18336 3883 18388
rect 3935 18336 3948 18388
rect 4000 18336 4013 18388
rect 4065 18336 4078 18388
rect 4130 18336 4143 18388
rect 4195 18336 4208 18388
rect 4260 18336 4273 18388
rect 4325 18336 4338 18388
rect 4390 18336 4403 18388
rect 4455 18336 4468 18388
rect 4520 18336 4532 18388
rect 4584 18375 5613 18388
rect 5669 18375 5696 18392
rect 4584 18336 5040 18375
rect 2444 18326 5040 18336
rect 2270 18323 5040 18326
rect 5092 18323 5106 18375
rect 5158 18323 5594 18375
rect 5752 18348 5779 18404
rect 5835 18348 5861 18404
rect 5917 18348 5943 18404
rect 5999 18348 6025 18404
rect 6081 18348 6107 18404
rect 6266 18392 6271 18404
rect 6163 18375 6189 18392
rect 6245 18375 6271 18392
rect 6266 18348 6271 18375
rect 6327 18348 6353 18404
rect 6409 18348 6435 18404
rect 6491 18348 6517 18404
rect 6573 18348 6599 18404
rect 6655 18348 6681 18404
rect 6754 18392 6763 18404
rect 6820 18392 6845 18404
rect 6737 18375 6763 18392
rect 6819 18375 6845 18392
rect 6754 18348 6763 18375
rect 6820 18348 6845 18375
rect 6901 18348 6927 18404
rect 6983 18348 7009 18404
rect 7065 18348 7091 18404
rect 7147 18348 7173 18404
rect 7229 18348 7255 18404
rect 7311 18392 7322 18404
rect 7311 18375 7337 18392
rect 7311 18348 7322 18375
rect 7393 18348 7419 18404
rect 7475 18348 7501 18404
rect 7557 18348 7583 18404
rect 7639 18348 7665 18404
rect 7721 18348 7747 18404
rect 7803 18392 7810 18404
rect 7803 18375 7829 18392
rect 7885 18375 7911 18392
rect 7803 18348 7810 18375
rect 7967 18348 7993 18404
rect 8049 18378 8075 18396
rect 8131 18348 8157 18404
rect 8221 18396 8222 18448
rect 8213 18378 8222 18396
rect 5646 18324 5660 18348
rect 5712 18324 6148 18348
rect 6200 18324 6214 18348
rect 6266 18324 6702 18348
rect 6754 18324 6768 18348
rect 6820 18324 7256 18348
rect 7308 18324 7322 18348
rect 7374 18324 7810 18348
rect 7862 18324 7876 18348
rect 7928 18326 8047 18348
rect 8099 18326 8169 18348
rect 8221 18326 8222 18378
rect 7928 18324 8222 18326
rect 2270 18320 5613 18323
rect 2270 18308 2648 18320
rect 2322 18256 2392 18308
rect 2444 18268 2648 18308
rect 2700 18268 2713 18320
rect 2765 18268 2778 18320
rect 2830 18268 2843 18320
rect 2895 18268 2908 18320
rect 2960 18268 2973 18320
rect 3025 18268 3038 18320
rect 3090 18268 3103 18320
rect 3155 18268 3168 18320
rect 3220 18268 3233 18320
rect 3285 18268 3298 18320
rect 3350 18268 3363 18320
rect 3415 18268 3428 18320
rect 3480 18268 3493 18320
rect 3545 18268 3558 18320
rect 3610 18268 3623 18320
rect 3675 18268 3688 18320
rect 3740 18268 3753 18320
rect 3805 18268 3818 18320
rect 3870 18268 3883 18320
rect 3935 18268 3948 18320
rect 4000 18268 4013 18320
rect 4065 18268 4078 18320
rect 4130 18268 4143 18320
rect 4195 18268 4208 18320
rect 4260 18268 4273 18320
rect 4325 18268 4338 18320
rect 4390 18268 4403 18320
rect 4455 18268 4468 18320
rect 4520 18268 4532 18320
rect 4584 18306 5613 18320
rect 5669 18306 5696 18323
rect 4584 18268 5040 18306
rect 2444 18256 5040 18268
rect 2270 18254 5040 18256
rect 5092 18254 5106 18306
rect 5158 18254 5594 18306
rect 5752 18268 5779 18324
rect 5835 18268 5861 18324
rect 5917 18268 5943 18324
rect 5999 18268 6025 18324
rect 6081 18268 6107 18324
rect 6266 18323 6271 18324
rect 6163 18306 6189 18323
rect 6245 18306 6271 18323
rect 6266 18268 6271 18306
rect 6327 18268 6353 18324
rect 6409 18268 6435 18324
rect 6491 18268 6517 18324
rect 6573 18268 6599 18324
rect 6655 18268 6681 18324
rect 6754 18323 6763 18324
rect 6820 18323 6845 18324
rect 6737 18306 6763 18323
rect 6819 18306 6845 18323
rect 6754 18268 6763 18306
rect 6820 18268 6845 18306
rect 6901 18268 6927 18324
rect 6983 18268 7009 18324
rect 7065 18268 7091 18324
rect 7147 18268 7173 18324
rect 7229 18268 7255 18324
rect 7311 18323 7322 18324
rect 7311 18306 7337 18323
rect 7311 18268 7322 18306
rect 7393 18268 7419 18324
rect 7475 18268 7501 18324
rect 7557 18268 7583 18324
rect 7639 18268 7665 18324
rect 7721 18268 7747 18324
rect 7803 18323 7810 18324
rect 7803 18306 7829 18323
rect 7885 18306 7911 18323
rect 7803 18268 7810 18306
rect 7967 18268 7993 18324
rect 8049 18308 8075 18324
rect 8131 18268 8157 18324
rect 8213 18308 8222 18324
rect 5646 18254 5660 18268
rect 5712 18254 6148 18268
rect 6200 18254 6214 18268
rect 6266 18254 6702 18268
rect 6754 18254 6768 18268
rect 6820 18254 7256 18268
rect 7308 18254 7322 18268
rect 7374 18254 7810 18268
rect 7862 18254 7876 18268
rect 7928 18256 8047 18268
rect 8099 18256 8169 18268
rect 8221 18256 8222 18308
rect 7928 18254 8222 18256
rect 2270 18252 8222 18254
rect 2270 18238 2648 18252
rect 2322 18186 2392 18238
rect 2444 18200 2648 18238
rect 2700 18200 2713 18252
rect 2765 18200 2778 18252
rect 2830 18200 2843 18252
rect 2895 18200 2908 18252
rect 2960 18200 2973 18252
rect 3025 18200 3038 18252
rect 3090 18200 3103 18252
rect 3155 18200 3168 18252
rect 3220 18200 3233 18252
rect 3285 18200 3298 18252
rect 3350 18200 3363 18252
rect 3415 18200 3428 18252
rect 3480 18200 3493 18252
rect 3545 18200 3558 18252
rect 3610 18200 3623 18252
rect 3675 18200 3688 18252
rect 3740 18200 3753 18252
rect 3805 18200 3818 18252
rect 3870 18200 3883 18252
rect 3935 18200 3948 18252
rect 4000 18200 4013 18252
rect 4065 18200 4078 18252
rect 4130 18200 4143 18252
rect 4195 18200 4208 18252
rect 4260 18200 4273 18252
rect 4325 18200 4338 18252
rect 4390 18200 4403 18252
rect 4455 18200 4468 18252
rect 4520 18200 4532 18252
rect 4584 18244 8222 18252
rect 4584 18236 5613 18244
rect 5669 18236 5696 18244
rect 4584 18200 5040 18236
rect 2444 18186 5040 18200
rect 2270 18184 5040 18186
rect 5092 18184 5106 18236
rect 5158 18184 5594 18236
rect 5752 18188 5779 18244
rect 5835 18188 5861 18244
rect 5917 18188 5943 18244
rect 5999 18188 6025 18244
rect 6081 18188 6107 18244
rect 6163 18236 6189 18244
rect 6245 18236 6271 18244
rect 6266 18188 6271 18236
rect 6327 18188 6353 18244
rect 6409 18188 6435 18244
rect 6491 18188 6517 18244
rect 6573 18188 6599 18244
rect 6655 18188 6681 18244
rect 6737 18236 6763 18244
rect 6819 18236 6845 18244
rect 6754 18188 6763 18236
rect 6820 18188 6845 18236
rect 6901 18188 6927 18244
rect 6983 18188 7009 18244
rect 7065 18188 7091 18244
rect 7147 18188 7173 18244
rect 7229 18188 7255 18244
rect 7311 18236 7337 18244
rect 7311 18188 7322 18236
rect 7393 18188 7419 18244
rect 7475 18188 7501 18244
rect 7557 18188 7583 18244
rect 7639 18188 7665 18244
rect 7721 18188 7747 18244
rect 7803 18236 7829 18244
rect 7885 18236 7911 18244
rect 7803 18188 7810 18236
rect 7967 18188 7993 18244
rect 8049 18238 8075 18244
rect 8131 18188 8157 18244
rect 8213 18238 8222 18244
rect 5646 18184 5660 18188
rect 5712 18184 6148 18188
rect 6200 18184 6214 18188
rect 6266 18184 6702 18188
rect 6754 18184 6768 18188
rect 6820 18184 7256 18188
rect 7308 18184 7322 18188
rect 7374 18184 7810 18188
rect 7862 18184 7876 18188
rect 7928 18186 8047 18188
rect 8099 18186 8169 18188
rect 8221 18186 8222 18238
rect 7928 18184 8222 18186
rect 2270 18168 8222 18184
rect 2322 18116 2392 18168
rect 2444 18166 8047 18168
rect 2444 18116 5040 18166
rect 2270 18114 5040 18116
rect 5092 18114 5106 18166
rect 5158 18114 5594 18166
rect 5646 18164 5660 18166
rect 5712 18164 6148 18166
rect 6200 18164 6214 18166
rect 6266 18164 6702 18166
rect 6754 18164 6768 18166
rect 6820 18164 7256 18166
rect 7308 18164 7322 18166
rect 7374 18164 7810 18166
rect 7862 18164 7876 18166
rect 7928 18164 8047 18166
rect 8099 18164 8169 18168
rect 2270 18108 5613 18114
rect 5669 18108 5696 18114
rect 5752 18108 5779 18164
rect 5835 18108 5861 18164
rect 5917 18108 5943 18164
rect 5999 18108 6025 18164
rect 6081 18108 6107 18164
rect 6266 18114 6271 18164
rect 6163 18108 6189 18114
rect 6245 18108 6271 18114
rect 6327 18108 6353 18164
rect 6409 18108 6435 18164
rect 6491 18108 6517 18164
rect 6573 18108 6599 18164
rect 6655 18108 6681 18164
rect 6754 18114 6763 18164
rect 6820 18114 6845 18164
rect 6737 18108 6763 18114
rect 6819 18108 6845 18114
rect 6901 18108 6927 18164
rect 6983 18108 7009 18164
rect 7065 18108 7091 18164
rect 7147 18108 7173 18164
rect 7229 18108 7255 18164
rect 7311 18114 7322 18164
rect 7311 18108 7337 18114
rect 7393 18108 7419 18164
rect 7475 18108 7501 18164
rect 7557 18108 7583 18164
rect 7639 18108 7665 18164
rect 7721 18108 7747 18164
rect 7803 18114 7810 18164
rect 7803 18108 7829 18114
rect 7885 18108 7911 18114
rect 7967 18108 7993 18164
rect 8049 18108 8075 18116
rect 8131 18108 8157 18164
rect 8221 18116 8222 18168
rect 8213 18108 8222 18116
rect 2724 17987 7651 17988
rect 2724 17931 2733 17987
rect 2789 17931 2814 17987
rect 2870 17931 2895 17987
rect 2951 17931 2976 17987
rect 3032 17931 3057 17987
rect 3113 17931 3138 17987
rect 3194 17931 3219 17987
rect 3275 17931 3300 17987
rect 3356 17931 3381 17987
rect 3437 17931 3462 17987
rect 3518 17931 3543 17987
rect 3599 17931 3624 17987
rect 3680 17931 3705 17987
rect 3761 17931 3786 17987
rect 3842 17931 3867 17987
rect 3923 17931 3948 17987
rect 4004 17931 4029 17987
rect 4085 17931 4110 17987
rect 4166 17931 4191 17987
rect 4247 17931 4272 17987
rect 4328 17931 4353 17987
rect 4409 17931 4434 17987
rect 4490 17931 4515 17987
rect 4571 17931 4596 17987
rect 4652 17931 4677 17987
rect 4733 17931 4758 17987
rect 4814 17931 4839 17987
rect 4895 17931 4920 17987
rect 4976 17931 5001 17987
rect 5057 17931 5082 17987
rect 5138 17931 5163 17987
rect 2724 17907 5163 17931
rect 2724 17851 2733 17907
rect 2789 17851 2814 17907
rect 2870 17851 2895 17907
rect 2951 17851 2976 17907
rect 3032 17851 3057 17907
rect 3113 17851 3138 17907
rect 3194 17851 3219 17907
rect 3275 17851 3300 17907
rect 3356 17851 3381 17907
rect 3437 17851 3462 17907
rect 3518 17851 3543 17907
rect 3599 17851 3624 17907
rect 3680 17851 3705 17907
rect 3761 17851 3786 17907
rect 3842 17851 3867 17907
rect 3923 17851 3948 17907
rect 4004 17851 4029 17907
rect 4085 17851 4110 17907
rect 4166 17851 4191 17907
rect 4247 17851 4272 17907
rect 4328 17851 4353 17907
rect 4409 17851 4434 17907
rect 4490 17851 4515 17907
rect 4571 17851 4596 17907
rect 4652 17851 4677 17907
rect 4733 17851 4758 17907
rect 4814 17851 4839 17907
rect 4895 17851 4920 17907
rect 4976 17851 5001 17907
rect 5057 17851 5082 17907
rect 5138 17851 5163 17907
rect 2724 17827 5163 17851
rect 2724 17771 2733 17827
rect 2789 17771 2814 17827
rect 2870 17771 2895 17827
rect 2951 17771 2976 17827
rect 3032 17771 3057 17827
rect 3113 17771 3138 17827
rect 3194 17771 3219 17827
rect 3275 17771 3300 17827
rect 3356 17771 3381 17827
rect 3437 17771 3462 17827
rect 3518 17771 3543 17827
rect 3599 17771 3624 17827
rect 3680 17771 3705 17827
rect 3761 17771 3786 17827
rect 3842 17771 3867 17827
rect 3923 17771 3948 17827
rect 4004 17771 4029 17827
rect 4085 17771 4110 17827
rect 4166 17771 4191 17827
rect 4247 17771 4272 17827
rect 4328 17771 4353 17827
rect 4409 17771 4434 17827
rect 4490 17771 4515 17827
rect 4571 17771 4596 17827
rect 4652 17771 4677 17827
rect 4733 17771 4758 17827
rect 4814 17771 4839 17827
rect 4895 17771 4920 17827
rect 4976 17771 5001 17827
rect 5057 17771 5082 17827
rect 5138 17771 5163 17827
rect 2724 17747 5163 17771
rect 2724 17691 2733 17747
rect 2789 17691 2814 17747
rect 2870 17691 2895 17747
rect 2951 17691 2976 17747
rect 3032 17691 3057 17747
rect 3113 17691 3138 17747
rect 3194 17691 3219 17747
rect 3275 17691 3300 17747
rect 3356 17691 3381 17747
rect 3437 17691 3462 17747
rect 3518 17691 3543 17747
rect 3599 17691 3624 17747
rect 3680 17691 3705 17747
rect 3761 17691 3786 17747
rect 3842 17691 3867 17747
rect 3923 17691 3948 17747
rect 4004 17691 4029 17747
rect 4085 17691 4110 17747
rect 4166 17691 4191 17747
rect 4247 17691 4272 17747
rect 4328 17691 4353 17747
rect 4409 17691 4434 17747
rect 4490 17691 4515 17747
rect 4571 17691 4596 17747
rect 4652 17691 4677 17747
rect 4733 17691 4758 17747
rect 4814 17691 4839 17747
rect 4895 17691 4920 17747
rect 4976 17691 5001 17747
rect 5057 17691 5082 17747
rect 5138 17691 5163 17747
rect 2724 17667 5163 17691
rect 2724 17611 2733 17667
rect 2789 17611 2814 17667
rect 2870 17611 2895 17667
rect 2951 17611 2976 17667
rect 3032 17611 3057 17667
rect 3113 17611 3138 17667
rect 3194 17611 3219 17667
rect 3275 17611 3300 17667
rect 3356 17611 3381 17667
rect 3437 17611 3462 17667
rect 3518 17611 3543 17667
rect 3599 17611 3624 17667
rect 3680 17611 3705 17667
rect 3761 17611 3786 17667
rect 3842 17611 3867 17667
rect 3923 17611 3948 17667
rect 4004 17611 4029 17667
rect 4085 17611 4110 17667
rect 4166 17611 4191 17667
rect 4247 17611 4272 17667
rect 4328 17611 4353 17667
rect 4409 17611 4434 17667
rect 4490 17611 4515 17667
rect 4571 17611 4596 17667
rect 4652 17611 4677 17667
rect 4733 17611 4758 17667
rect 4814 17611 4839 17667
rect 4895 17611 4920 17667
rect 4976 17611 5001 17667
rect 5057 17611 5082 17667
rect 5138 17611 5163 17667
rect 2724 17587 5163 17611
rect 2724 17531 2733 17587
rect 2789 17531 2814 17587
rect 2870 17531 2895 17587
rect 2951 17531 2976 17587
rect 3032 17531 3057 17587
rect 3113 17531 3138 17587
rect 3194 17531 3219 17587
rect 3275 17531 3300 17587
rect 3356 17531 3381 17587
rect 3437 17531 3462 17587
rect 3518 17531 3543 17587
rect 3599 17531 3624 17587
rect 3680 17531 3705 17587
rect 3761 17531 3786 17587
rect 3842 17531 3867 17587
rect 3923 17531 3948 17587
rect 4004 17531 4029 17587
rect 4085 17531 4110 17587
rect 4166 17531 4191 17587
rect 4247 17531 4272 17587
rect 4328 17531 4353 17587
rect 4409 17531 4434 17587
rect 4490 17531 4515 17587
rect 4571 17531 4596 17587
rect 4652 17531 4677 17587
rect 4733 17531 4758 17587
rect 4814 17531 4839 17587
rect 4895 17531 4920 17587
rect 4976 17531 5001 17587
rect 5057 17531 5082 17587
rect 5138 17531 5163 17587
rect 2724 17507 5163 17531
rect 2724 17451 2733 17507
rect 2789 17451 2814 17507
rect 2870 17451 2895 17507
rect 2951 17451 2976 17507
rect 3032 17451 3057 17507
rect 3113 17451 3138 17507
rect 3194 17451 3219 17507
rect 3275 17451 3300 17507
rect 3356 17451 3381 17507
rect 3437 17451 3462 17507
rect 3518 17451 3543 17507
rect 3599 17451 3624 17507
rect 3680 17451 3705 17507
rect 3761 17451 3786 17507
rect 3842 17451 3867 17507
rect 3923 17451 3948 17507
rect 4004 17451 4029 17507
rect 4085 17451 4110 17507
rect 4166 17451 4191 17507
rect 4247 17451 4272 17507
rect 4328 17451 4353 17507
rect 4409 17451 4434 17507
rect 4490 17451 4515 17507
rect 4571 17451 4596 17507
rect 4652 17451 4677 17507
rect 4733 17451 4758 17507
rect 4814 17451 4839 17507
rect 4895 17451 4920 17507
rect 4976 17451 5001 17507
rect 5057 17451 5082 17507
rect 5138 17451 5163 17507
rect 2724 17427 5163 17451
rect 2724 17371 2733 17427
rect 2789 17371 2814 17427
rect 2870 17371 2895 17427
rect 2951 17371 2976 17427
rect 3032 17371 3057 17427
rect 3113 17371 3138 17427
rect 3194 17371 3219 17427
rect 3275 17371 3300 17427
rect 3356 17371 3381 17427
rect 3437 17371 3462 17427
rect 3518 17371 3543 17427
rect 3599 17371 3624 17427
rect 3680 17371 3705 17427
rect 3761 17371 3786 17427
rect 3842 17371 3867 17427
rect 3923 17371 3948 17427
rect 4004 17371 4029 17427
rect 4085 17371 4110 17427
rect 4166 17371 4191 17427
rect 4247 17371 4272 17427
rect 4328 17371 4353 17427
rect 4409 17371 4434 17427
rect 4490 17371 4515 17427
rect 4571 17371 4596 17427
rect 4652 17371 4677 17427
rect 4733 17371 4758 17427
rect 4814 17371 4839 17427
rect 4895 17371 4920 17427
rect 4976 17371 5001 17427
rect 5057 17371 5082 17427
rect 5138 17371 5163 17427
rect 5299 17982 7651 17987
rect 5299 17930 5317 17982
rect 5369 17930 5383 17982
rect 5435 17930 5871 17982
rect 5923 17930 5937 17982
rect 5989 17930 6425 17982
rect 6477 17930 6491 17982
rect 6543 17930 6979 17982
rect 7031 17930 7045 17982
rect 7097 17930 7533 17982
rect 7585 17930 7599 17982
rect 5299 17913 7651 17930
rect 5299 17861 5317 17913
rect 5369 17861 5383 17913
rect 5435 17861 5871 17913
rect 5923 17861 5937 17913
rect 5989 17861 6425 17913
rect 6477 17861 6491 17913
rect 6543 17861 6979 17913
rect 7031 17861 7045 17913
rect 7097 17861 7533 17913
rect 7585 17861 7599 17913
rect 5299 17844 7651 17861
rect 5299 17792 5317 17844
rect 5369 17792 5383 17844
rect 5435 17792 5871 17844
rect 5923 17792 5937 17844
rect 5989 17792 6425 17844
rect 6477 17792 6491 17844
rect 6543 17792 6979 17844
rect 7031 17792 7045 17844
rect 7097 17792 7533 17844
rect 7585 17792 7599 17844
rect 5299 17775 7651 17792
rect 5299 17723 5317 17775
rect 5369 17723 5383 17775
rect 5435 17723 5871 17775
rect 5923 17723 5937 17775
rect 5989 17723 6425 17775
rect 6477 17723 6491 17775
rect 6543 17723 6979 17775
rect 7031 17723 7045 17775
rect 7097 17723 7533 17775
rect 7585 17723 7599 17775
rect 5299 17706 7651 17723
rect 5299 17654 5317 17706
rect 5369 17654 5383 17706
rect 5435 17654 5871 17706
rect 5923 17654 5937 17706
rect 5989 17654 6425 17706
rect 6477 17654 6491 17706
rect 6543 17654 6979 17706
rect 7031 17654 7045 17706
rect 7097 17654 7533 17706
rect 7585 17654 7599 17706
rect 5299 17636 7651 17654
rect 5299 17584 5317 17636
rect 5369 17584 5383 17636
rect 5435 17584 5871 17636
rect 5923 17584 5937 17636
rect 5989 17584 6425 17636
rect 6477 17584 6491 17636
rect 6543 17584 6979 17636
rect 7031 17584 7045 17636
rect 7097 17584 7533 17636
rect 7585 17584 7599 17636
rect 5299 17566 7651 17584
rect 5299 17514 5317 17566
rect 5369 17514 5383 17566
rect 5435 17514 5871 17566
rect 5923 17514 5937 17566
rect 5989 17514 6425 17566
rect 6477 17514 6491 17566
rect 6543 17514 6979 17566
rect 7031 17514 7045 17566
rect 7097 17514 7533 17566
rect 7585 17514 7599 17566
rect 5299 17496 7651 17514
rect 5299 17444 5317 17496
rect 5369 17444 5383 17496
rect 5435 17444 5871 17496
rect 5923 17444 5937 17496
rect 5989 17444 6425 17496
rect 6477 17444 6491 17496
rect 6543 17444 6979 17496
rect 7031 17444 7045 17496
rect 7097 17444 7533 17496
rect 7585 17444 7599 17496
rect 5299 17426 7651 17444
rect 5299 17374 5317 17426
rect 5369 17374 5383 17426
rect 5435 17374 5871 17426
rect 5923 17374 5937 17426
rect 5989 17374 6425 17426
rect 6477 17374 6491 17426
rect 6543 17374 6979 17426
rect 7031 17374 7045 17426
rect 7097 17374 7533 17426
rect 7585 17374 7599 17426
rect 5299 17371 7651 17374
rect 2724 17368 7651 17371
rect 2270 16973 8222 16979
rect 2322 16921 2392 16973
rect 2444 16970 8047 16973
rect 2444 16921 2746 16970
rect 2270 16918 2746 16921
rect 2798 16918 2813 16970
rect 2865 16918 2880 16970
rect 2932 16918 2946 16970
rect 2998 16918 3012 16970
rect 3064 16918 3078 16970
rect 3130 16918 3144 16970
rect 3196 16918 3210 16970
rect 3262 16918 3276 16970
rect 3328 16918 3342 16970
rect 3394 16918 3408 16970
rect 3460 16918 3474 16970
rect 3526 16918 3540 16970
rect 3592 16918 3606 16970
rect 3658 16918 3672 16970
rect 3724 16918 3738 16970
rect 3790 16918 3804 16970
rect 3856 16918 3870 16970
rect 3922 16918 3936 16970
rect 3988 16918 4002 16970
rect 4054 16918 4068 16970
rect 4120 16918 4134 16970
rect 4186 16918 4200 16970
rect 4252 16918 4266 16970
rect 4318 16918 4332 16970
rect 4384 16918 4398 16970
rect 4450 16918 4464 16970
rect 4516 16918 5116 16970
rect 5168 16918 5182 16970
rect 5234 16918 5248 16970
rect 5300 16918 5314 16970
rect 5366 16918 5380 16970
rect 5432 16918 5446 16970
rect 5498 16918 5512 16970
rect 5564 16918 5578 16970
rect 5630 16918 5644 16970
rect 5696 16918 5710 16970
rect 5762 16918 5776 16970
rect 5828 16918 5842 16970
rect 5894 16918 5908 16970
rect 5960 16918 5974 16970
rect 6026 16918 6040 16970
rect 6092 16918 6106 16970
rect 6158 16918 6172 16970
rect 6224 16918 6238 16970
rect 6290 16918 6304 16970
rect 6356 16918 6370 16970
rect 6422 16918 6436 16970
rect 6488 16918 6501 16970
rect 6553 16918 6566 16970
rect 6618 16918 6631 16970
rect 6683 16918 6696 16970
rect 6748 16918 6761 16970
rect 6813 16918 6826 16970
rect 6878 16918 6891 16970
rect 6943 16918 6956 16970
rect 7008 16918 7021 16970
rect 7073 16918 7086 16970
rect 7138 16918 7151 16970
rect 7203 16918 7216 16970
rect 7268 16918 7281 16970
rect 7333 16918 7346 16970
rect 7398 16918 7411 16970
rect 7463 16918 7476 16970
rect 7528 16918 7541 16970
rect 7593 16918 7606 16970
rect 7658 16918 7671 16970
rect 7723 16918 7736 16970
rect 7788 16918 7801 16970
rect 7853 16921 8047 16970
rect 8099 16921 8169 16973
rect 8221 16921 8222 16973
rect 7853 16918 8222 16921
rect 2270 16907 8222 16918
rect 2322 16855 2392 16907
rect 2444 16904 8047 16907
rect 2444 16855 2746 16904
rect 2270 16852 2746 16855
rect 2798 16852 2813 16904
rect 2865 16852 2880 16904
rect 2932 16852 2946 16904
rect 2998 16852 3012 16904
rect 3064 16852 3078 16904
rect 3130 16852 3144 16904
rect 3196 16852 3210 16904
rect 3262 16852 3276 16904
rect 3328 16852 3342 16904
rect 3394 16852 3408 16904
rect 3460 16852 3474 16904
rect 3526 16852 3540 16904
rect 3592 16852 3606 16904
rect 3658 16852 3672 16904
rect 3724 16852 3738 16904
rect 3790 16852 3804 16904
rect 3856 16852 3870 16904
rect 3922 16852 3936 16904
rect 3988 16852 4002 16904
rect 4054 16852 4068 16904
rect 4120 16852 4134 16904
rect 4186 16852 4200 16904
rect 4252 16852 4266 16904
rect 4318 16852 4332 16904
rect 4384 16852 4398 16904
rect 4450 16852 4464 16904
rect 4516 16852 5116 16904
rect 5168 16852 5182 16904
rect 5234 16852 5248 16904
rect 5300 16852 5314 16904
rect 5366 16852 5380 16904
rect 5432 16852 5446 16904
rect 5498 16852 5512 16904
rect 5564 16852 5578 16904
rect 5630 16852 5644 16904
rect 5696 16852 5710 16904
rect 5762 16852 5776 16904
rect 5828 16852 5842 16904
rect 5894 16852 5908 16904
rect 5960 16852 5974 16904
rect 6026 16852 6040 16904
rect 6092 16852 6106 16904
rect 6158 16852 6172 16904
rect 6224 16852 6238 16904
rect 6290 16852 6304 16904
rect 6356 16852 6370 16904
rect 6422 16852 6436 16904
rect 6488 16852 6501 16904
rect 6553 16852 6566 16904
rect 6618 16852 6631 16904
rect 6683 16852 6696 16904
rect 6748 16852 6761 16904
rect 6813 16852 6826 16904
rect 6878 16852 6891 16904
rect 6943 16852 6956 16904
rect 7008 16852 7021 16904
rect 7073 16852 7086 16904
rect 7138 16852 7151 16904
rect 7203 16852 7216 16904
rect 7268 16852 7281 16904
rect 7333 16852 7346 16904
rect 7398 16852 7411 16904
rect 7463 16852 7476 16904
rect 7528 16852 7541 16904
rect 7593 16852 7606 16904
rect 7658 16852 7671 16904
rect 7723 16852 7736 16904
rect 7788 16852 7801 16904
rect 7853 16855 8047 16904
rect 8099 16855 8169 16907
rect 8221 16855 8222 16907
rect 7853 16852 8222 16855
rect 2270 16841 8222 16852
rect 2322 16789 2392 16841
rect 2444 16838 8047 16841
rect 2444 16789 2746 16838
rect 2270 16786 2746 16789
rect 2798 16786 2813 16838
rect 2865 16786 2880 16838
rect 2932 16786 2946 16838
rect 2998 16786 3012 16838
rect 3064 16786 3078 16838
rect 3130 16786 3144 16838
rect 3196 16786 3210 16838
rect 3262 16786 3276 16838
rect 3328 16786 3342 16838
rect 3394 16786 3408 16838
rect 3460 16786 3474 16838
rect 3526 16786 3540 16838
rect 3592 16786 3606 16838
rect 3658 16786 3672 16838
rect 3724 16786 3738 16838
rect 3790 16786 3804 16838
rect 3856 16786 3870 16838
rect 3922 16786 3936 16838
rect 3988 16786 4002 16838
rect 4054 16786 4068 16838
rect 4120 16786 4134 16838
rect 4186 16786 4200 16838
rect 4252 16786 4266 16838
rect 4318 16786 4332 16838
rect 4384 16786 4398 16838
rect 4450 16786 4464 16838
rect 4516 16786 5116 16838
rect 5168 16786 5182 16838
rect 5234 16786 5248 16838
rect 5300 16786 5314 16838
rect 5366 16786 5380 16838
rect 5432 16786 5446 16838
rect 5498 16786 5512 16838
rect 5564 16786 5578 16838
rect 5630 16786 5644 16838
rect 5696 16786 5710 16838
rect 5762 16786 5776 16838
rect 5828 16786 5842 16838
rect 5894 16786 5908 16838
rect 5960 16786 5974 16838
rect 6026 16786 6040 16838
rect 6092 16786 6106 16838
rect 6158 16786 6172 16838
rect 6224 16786 6238 16838
rect 6290 16786 6304 16838
rect 6356 16786 6370 16838
rect 6422 16786 6436 16838
rect 6488 16786 6501 16838
rect 6553 16786 6566 16838
rect 6618 16786 6631 16838
rect 6683 16786 6696 16838
rect 6748 16786 6761 16838
rect 6813 16786 6826 16838
rect 6878 16786 6891 16838
rect 6943 16786 6956 16838
rect 7008 16786 7021 16838
rect 7073 16786 7086 16838
rect 7138 16786 7151 16838
rect 7203 16786 7216 16838
rect 7268 16786 7281 16838
rect 7333 16786 7346 16838
rect 7398 16786 7411 16838
rect 7463 16786 7476 16838
rect 7528 16786 7541 16838
rect 7593 16786 7606 16838
rect 7658 16786 7671 16838
rect 7723 16786 7736 16838
rect 7788 16786 7801 16838
rect 7853 16789 8047 16838
rect 8099 16789 8169 16841
rect 8221 16789 8222 16841
rect 7853 16786 8222 16789
rect 2270 16775 8222 16786
rect 2322 16723 2392 16775
rect 2444 16772 8047 16775
rect 2444 16723 2746 16772
rect 2270 16720 2746 16723
rect 2798 16720 2813 16772
rect 2865 16720 2880 16772
rect 2932 16720 2946 16772
rect 2998 16720 3012 16772
rect 3064 16720 3078 16772
rect 3130 16720 3144 16772
rect 3196 16720 3210 16772
rect 3262 16720 3276 16772
rect 3328 16720 3342 16772
rect 3394 16720 3408 16772
rect 3460 16720 3474 16772
rect 3526 16720 3540 16772
rect 3592 16720 3606 16772
rect 3658 16720 3672 16772
rect 3724 16720 3738 16772
rect 3790 16720 3804 16772
rect 3856 16720 3870 16772
rect 3922 16720 3936 16772
rect 3988 16720 4002 16772
rect 4054 16720 4068 16772
rect 4120 16720 4134 16772
rect 4186 16720 4200 16772
rect 4252 16720 4266 16772
rect 4318 16720 4332 16772
rect 4384 16720 4398 16772
rect 4450 16720 4464 16772
rect 4516 16720 5116 16772
rect 5168 16720 5182 16772
rect 5234 16720 5248 16772
rect 5300 16720 5314 16772
rect 5366 16720 5380 16772
rect 5432 16720 5446 16772
rect 5498 16720 5512 16772
rect 5564 16720 5578 16772
rect 5630 16720 5644 16772
rect 5696 16720 5710 16772
rect 5762 16720 5776 16772
rect 5828 16720 5842 16772
rect 5894 16720 5908 16772
rect 5960 16720 5974 16772
rect 6026 16720 6040 16772
rect 6092 16720 6106 16772
rect 6158 16720 6172 16772
rect 6224 16720 6238 16772
rect 6290 16720 6304 16772
rect 6356 16720 6370 16772
rect 6422 16720 6436 16772
rect 6488 16720 6501 16772
rect 6553 16720 6566 16772
rect 6618 16720 6631 16772
rect 6683 16720 6696 16772
rect 6748 16720 6761 16772
rect 6813 16720 6826 16772
rect 6878 16720 6891 16772
rect 6943 16720 6956 16772
rect 7008 16720 7021 16772
rect 7073 16720 7086 16772
rect 7138 16720 7151 16772
rect 7203 16720 7216 16772
rect 7268 16720 7281 16772
rect 7333 16720 7346 16772
rect 7398 16720 7411 16772
rect 7463 16720 7476 16772
rect 7528 16720 7541 16772
rect 7593 16720 7606 16772
rect 7658 16720 7671 16772
rect 7723 16720 7736 16772
rect 7788 16720 7801 16772
rect 7853 16723 8047 16772
rect 8099 16723 8169 16775
rect 8221 16723 8222 16775
rect 7853 16720 8222 16723
rect 2270 16709 8222 16720
rect 2322 16657 2392 16709
rect 2444 16706 8047 16709
rect 2444 16657 2746 16706
rect 2270 16654 2746 16657
rect 2798 16654 2813 16706
rect 2865 16654 2880 16706
rect 2932 16654 2946 16706
rect 2998 16654 3012 16706
rect 3064 16654 3078 16706
rect 3130 16654 3144 16706
rect 3196 16654 3210 16706
rect 3262 16654 3276 16706
rect 3328 16654 3342 16706
rect 3394 16654 3408 16706
rect 3460 16654 3474 16706
rect 3526 16654 3540 16706
rect 3592 16654 3606 16706
rect 3658 16654 3672 16706
rect 3724 16654 3738 16706
rect 3790 16654 3804 16706
rect 3856 16654 3870 16706
rect 3922 16654 3936 16706
rect 3988 16654 4002 16706
rect 4054 16654 4068 16706
rect 4120 16654 4134 16706
rect 4186 16654 4200 16706
rect 4252 16654 4266 16706
rect 4318 16654 4332 16706
rect 4384 16654 4398 16706
rect 4450 16654 4464 16706
rect 4516 16654 5116 16706
rect 5168 16654 5182 16706
rect 5234 16654 5248 16706
rect 5300 16654 5314 16706
rect 5366 16654 5380 16706
rect 5432 16654 5446 16706
rect 5498 16654 5512 16706
rect 5564 16654 5578 16706
rect 5630 16654 5644 16706
rect 5696 16654 5710 16706
rect 5762 16654 5776 16706
rect 5828 16654 5842 16706
rect 5894 16654 5908 16706
rect 5960 16654 5974 16706
rect 6026 16654 6040 16706
rect 6092 16654 6106 16706
rect 6158 16654 6172 16706
rect 6224 16654 6238 16706
rect 6290 16654 6304 16706
rect 6356 16654 6370 16706
rect 6422 16654 6436 16706
rect 6488 16654 6501 16706
rect 6553 16654 6566 16706
rect 6618 16654 6631 16706
rect 6683 16654 6696 16706
rect 6748 16654 6761 16706
rect 6813 16654 6826 16706
rect 6878 16654 6891 16706
rect 6943 16654 6956 16706
rect 7008 16654 7021 16706
rect 7073 16654 7086 16706
rect 7138 16654 7151 16706
rect 7203 16654 7216 16706
rect 7268 16654 7281 16706
rect 7333 16654 7346 16706
rect 7398 16654 7411 16706
rect 7463 16654 7476 16706
rect 7528 16654 7541 16706
rect 7593 16654 7606 16706
rect 7658 16654 7671 16706
rect 7723 16654 7736 16706
rect 7788 16654 7801 16706
rect 7853 16657 8047 16706
rect 8099 16657 8169 16709
rect 8221 16657 8222 16709
rect 7853 16654 8222 16657
rect 2270 16643 8222 16654
rect 2322 16591 2392 16643
rect 2444 16640 8047 16643
rect 2444 16591 2746 16640
rect 2270 16588 2746 16591
rect 2798 16588 2813 16640
rect 2865 16588 2880 16640
rect 2932 16588 2946 16640
rect 2998 16588 3012 16640
rect 3064 16588 3078 16640
rect 3130 16588 3144 16640
rect 3196 16588 3210 16640
rect 3262 16588 3276 16640
rect 3328 16588 3342 16640
rect 3394 16588 3408 16640
rect 3460 16588 3474 16640
rect 3526 16588 3540 16640
rect 3592 16588 3606 16640
rect 3658 16588 3672 16640
rect 3724 16588 3738 16640
rect 3790 16588 3804 16640
rect 3856 16588 3870 16640
rect 3922 16588 3936 16640
rect 3988 16588 4002 16640
rect 4054 16588 4068 16640
rect 4120 16588 4134 16640
rect 4186 16588 4200 16640
rect 4252 16588 4266 16640
rect 4318 16588 4332 16640
rect 4384 16588 4398 16640
rect 4450 16588 4464 16640
rect 4516 16588 5116 16640
rect 5168 16588 5182 16640
rect 5234 16588 5248 16640
rect 5300 16588 5314 16640
rect 5366 16588 5380 16640
rect 5432 16588 5446 16640
rect 5498 16588 5512 16640
rect 5564 16588 5578 16640
rect 5630 16588 5644 16640
rect 5696 16588 5710 16640
rect 5762 16588 5776 16640
rect 5828 16588 5842 16640
rect 5894 16588 5908 16640
rect 5960 16588 5974 16640
rect 6026 16588 6040 16640
rect 6092 16588 6106 16640
rect 6158 16588 6172 16640
rect 6224 16588 6238 16640
rect 6290 16588 6304 16640
rect 6356 16588 6370 16640
rect 6422 16588 6436 16640
rect 6488 16588 6501 16640
rect 6553 16588 6566 16640
rect 6618 16588 6631 16640
rect 6683 16588 6696 16640
rect 6748 16588 6761 16640
rect 6813 16588 6826 16640
rect 6878 16588 6891 16640
rect 6943 16588 6956 16640
rect 7008 16588 7021 16640
rect 7073 16588 7086 16640
rect 7138 16588 7151 16640
rect 7203 16588 7216 16640
rect 7268 16588 7281 16640
rect 7333 16588 7346 16640
rect 7398 16588 7411 16640
rect 7463 16588 7476 16640
rect 7528 16588 7541 16640
rect 7593 16588 7606 16640
rect 7658 16588 7671 16640
rect 7723 16588 7736 16640
rect 7788 16588 7801 16640
rect 7853 16591 8047 16640
rect 8099 16591 8169 16643
rect 8221 16591 8222 16643
rect 7853 16588 8222 16591
rect 2270 16577 8222 16588
rect 2322 16525 2392 16577
rect 2444 16574 8047 16577
rect 2444 16525 2746 16574
rect 2270 16522 2746 16525
rect 2798 16522 2813 16574
rect 2865 16522 2880 16574
rect 2932 16522 2946 16574
rect 2998 16522 3012 16574
rect 3064 16522 3078 16574
rect 3130 16522 3144 16574
rect 3196 16522 3210 16574
rect 3262 16522 3276 16574
rect 3328 16522 3342 16574
rect 3394 16522 3408 16574
rect 3460 16522 3474 16574
rect 3526 16522 3540 16574
rect 3592 16522 3606 16574
rect 3658 16522 3672 16574
rect 3724 16522 3738 16574
rect 3790 16522 3804 16574
rect 3856 16522 3870 16574
rect 3922 16522 3936 16574
rect 3988 16522 4002 16574
rect 4054 16522 4068 16574
rect 4120 16522 4134 16574
rect 4186 16522 4200 16574
rect 4252 16522 4266 16574
rect 4318 16522 4332 16574
rect 4384 16522 4398 16574
rect 4450 16522 4464 16574
rect 4516 16522 5116 16574
rect 5168 16522 5182 16574
rect 5234 16522 5248 16574
rect 5300 16522 5314 16574
rect 5366 16522 5380 16574
rect 5432 16522 5446 16574
rect 5498 16522 5512 16574
rect 5564 16522 5578 16574
rect 5630 16522 5644 16574
rect 5696 16522 5710 16574
rect 5762 16522 5776 16574
rect 5828 16522 5842 16574
rect 5894 16522 5908 16574
rect 5960 16522 5974 16574
rect 6026 16522 6040 16574
rect 6092 16522 6106 16574
rect 6158 16522 6172 16574
rect 6224 16522 6238 16574
rect 6290 16522 6304 16574
rect 6356 16522 6370 16574
rect 6422 16522 6436 16574
rect 6488 16522 6501 16574
rect 6553 16522 6566 16574
rect 6618 16522 6631 16574
rect 6683 16522 6696 16574
rect 6748 16522 6761 16574
rect 6813 16522 6826 16574
rect 6878 16522 6891 16574
rect 6943 16522 6956 16574
rect 7008 16522 7021 16574
rect 7073 16522 7086 16574
rect 7138 16522 7151 16574
rect 7203 16522 7216 16574
rect 7268 16522 7281 16574
rect 7333 16522 7346 16574
rect 7398 16522 7411 16574
rect 7463 16522 7476 16574
rect 7528 16522 7541 16574
rect 7593 16522 7606 16574
rect 7658 16522 7671 16574
rect 7723 16522 7736 16574
rect 7788 16522 7801 16574
rect 7853 16525 8047 16574
rect 8099 16525 8169 16577
rect 8221 16525 8222 16577
rect 7853 16522 8222 16525
rect 2270 16511 8222 16522
rect 2322 16459 2392 16511
rect 2444 16508 8047 16511
rect 2444 16459 2746 16508
rect 2270 16456 2746 16459
rect 2798 16456 2813 16508
rect 2865 16456 2880 16508
rect 2932 16456 2946 16508
rect 2998 16456 3012 16508
rect 3064 16456 3078 16508
rect 3130 16456 3144 16508
rect 3196 16456 3210 16508
rect 3262 16456 3276 16508
rect 3328 16456 3342 16508
rect 3394 16456 3408 16508
rect 3460 16456 3474 16508
rect 3526 16456 3540 16508
rect 3592 16456 3606 16508
rect 3658 16456 3672 16508
rect 3724 16456 3738 16508
rect 3790 16456 3804 16508
rect 3856 16456 3870 16508
rect 3922 16456 3936 16508
rect 3988 16456 4002 16508
rect 4054 16456 4068 16508
rect 4120 16456 4134 16508
rect 4186 16456 4200 16508
rect 4252 16456 4266 16508
rect 4318 16456 4332 16508
rect 4384 16456 4398 16508
rect 4450 16456 4464 16508
rect 4516 16456 5116 16508
rect 5168 16456 5182 16508
rect 5234 16456 5248 16508
rect 5300 16456 5314 16508
rect 5366 16456 5380 16508
rect 5432 16456 5446 16508
rect 5498 16456 5512 16508
rect 5564 16456 5578 16508
rect 5630 16456 5644 16508
rect 5696 16456 5710 16508
rect 5762 16456 5776 16508
rect 5828 16456 5842 16508
rect 5894 16456 5908 16508
rect 5960 16456 5974 16508
rect 6026 16456 6040 16508
rect 6092 16456 6106 16508
rect 6158 16456 6172 16508
rect 6224 16456 6238 16508
rect 6290 16456 6304 16508
rect 6356 16456 6370 16508
rect 6422 16456 6436 16508
rect 6488 16456 6501 16508
rect 6553 16456 6566 16508
rect 6618 16456 6631 16508
rect 6683 16456 6696 16508
rect 6748 16456 6761 16508
rect 6813 16456 6826 16508
rect 6878 16456 6891 16508
rect 6943 16456 6956 16508
rect 7008 16456 7021 16508
rect 7073 16456 7086 16508
rect 7138 16456 7151 16508
rect 7203 16456 7216 16508
rect 7268 16456 7281 16508
rect 7333 16456 7346 16508
rect 7398 16456 7411 16508
rect 7463 16456 7476 16508
rect 7528 16456 7541 16508
rect 7593 16456 7606 16508
rect 7658 16456 7671 16508
rect 7723 16456 7736 16508
rect 7788 16456 7801 16508
rect 7853 16459 8047 16508
rect 8099 16459 8169 16511
rect 8221 16459 8222 16511
rect 7853 16456 8222 16459
rect 2270 16445 8222 16456
rect 2322 16393 2392 16445
rect 2444 16442 8047 16445
rect 2444 16393 2746 16442
rect 2270 16390 2746 16393
rect 2798 16390 2813 16442
rect 2865 16390 2880 16442
rect 2932 16390 2946 16442
rect 2998 16390 3012 16442
rect 3064 16390 3078 16442
rect 3130 16390 3144 16442
rect 3196 16390 3210 16442
rect 3262 16390 3276 16442
rect 3328 16390 3342 16442
rect 3394 16390 3408 16442
rect 3460 16390 3474 16442
rect 3526 16390 3540 16442
rect 3592 16390 3606 16442
rect 3658 16390 3672 16442
rect 3724 16390 3738 16442
rect 3790 16390 3804 16442
rect 3856 16390 3870 16442
rect 3922 16390 3936 16442
rect 3988 16390 4002 16442
rect 4054 16390 4068 16442
rect 4120 16390 4134 16442
rect 4186 16390 4200 16442
rect 4252 16390 4266 16442
rect 4318 16390 4332 16442
rect 4384 16390 4398 16442
rect 4450 16390 4464 16442
rect 4516 16390 5116 16442
rect 5168 16390 5182 16442
rect 5234 16390 5248 16442
rect 5300 16390 5314 16442
rect 5366 16390 5380 16442
rect 5432 16390 5446 16442
rect 5498 16390 5512 16442
rect 5564 16390 5578 16442
rect 5630 16390 5644 16442
rect 5696 16390 5710 16442
rect 5762 16390 5776 16442
rect 5828 16390 5842 16442
rect 5894 16390 5908 16442
rect 5960 16390 5974 16442
rect 6026 16390 6040 16442
rect 6092 16390 6106 16442
rect 6158 16390 6172 16442
rect 6224 16390 6238 16442
rect 6290 16390 6304 16442
rect 6356 16390 6370 16442
rect 6422 16390 6436 16442
rect 6488 16390 6501 16442
rect 6553 16390 6566 16442
rect 6618 16390 6631 16442
rect 6683 16390 6696 16442
rect 6748 16390 6761 16442
rect 6813 16390 6826 16442
rect 6878 16390 6891 16442
rect 6943 16390 6956 16442
rect 7008 16390 7021 16442
rect 7073 16390 7086 16442
rect 7138 16390 7151 16442
rect 7203 16390 7216 16442
rect 7268 16390 7281 16442
rect 7333 16390 7346 16442
rect 7398 16390 7411 16442
rect 7463 16390 7476 16442
rect 7528 16390 7541 16442
rect 7593 16390 7606 16442
rect 7658 16390 7671 16442
rect 7723 16390 7736 16442
rect 7788 16390 7801 16442
rect 7853 16393 8047 16442
rect 8099 16393 8169 16445
rect 8221 16393 8222 16445
rect 7853 16390 8222 16393
rect 2270 16378 8222 16390
rect 2322 16326 2392 16378
rect 2444 16376 8047 16378
rect 2444 16326 2746 16376
rect 2270 16324 2746 16326
rect 2798 16324 2813 16376
rect 2865 16324 2880 16376
rect 2932 16324 2946 16376
rect 2998 16324 3012 16376
rect 3064 16324 3078 16376
rect 3130 16324 3144 16376
rect 3196 16324 3210 16376
rect 3262 16324 3276 16376
rect 3328 16324 3342 16376
rect 3394 16324 3408 16376
rect 3460 16324 3474 16376
rect 3526 16324 3540 16376
rect 3592 16324 3606 16376
rect 3658 16324 3672 16376
rect 3724 16324 3738 16376
rect 3790 16324 3804 16376
rect 3856 16324 3870 16376
rect 3922 16324 3936 16376
rect 3988 16324 4002 16376
rect 4054 16324 4068 16376
rect 4120 16324 4134 16376
rect 4186 16324 4200 16376
rect 4252 16324 4266 16376
rect 4318 16324 4332 16376
rect 4384 16324 4398 16376
rect 4450 16324 4464 16376
rect 4516 16324 5116 16376
rect 5168 16324 5182 16376
rect 5234 16324 5248 16376
rect 5300 16324 5314 16376
rect 5366 16324 5380 16376
rect 5432 16324 5446 16376
rect 5498 16324 5512 16376
rect 5564 16324 5578 16376
rect 5630 16324 5644 16376
rect 5696 16324 5710 16376
rect 5762 16324 5776 16376
rect 5828 16324 5842 16376
rect 5894 16324 5908 16376
rect 5960 16324 5974 16376
rect 6026 16324 6040 16376
rect 6092 16324 6106 16376
rect 6158 16324 6172 16376
rect 6224 16324 6238 16376
rect 6290 16324 6304 16376
rect 6356 16324 6370 16376
rect 6422 16324 6436 16376
rect 6488 16324 6501 16376
rect 6553 16324 6566 16376
rect 6618 16324 6631 16376
rect 6683 16324 6696 16376
rect 6748 16324 6761 16376
rect 6813 16324 6826 16376
rect 6878 16324 6891 16376
rect 6943 16324 6956 16376
rect 7008 16324 7021 16376
rect 7073 16324 7086 16376
rect 7138 16324 7151 16376
rect 7203 16324 7216 16376
rect 7268 16324 7281 16376
rect 7333 16324 7346 16376
rect 7398 16324 7411 16376
rect 7463 16324 7476 16376
rect 7528 16324 7541 16376
rect 7593 16324 7606 16376
rect 7658 16324 7671 16376
rect 7723 16324 7736 16376
rect 7788 16324 7801 16376
rect 7853 16326 8047 16376
rect 8099 16326 8169 16378
rect 8221 16326 8222 16378
rect 7853 16324 8222 16326
rect 2270 16311 8222 16324
rect 2322 16259 2392 16311
rect 2444 16310 8047 16311
rect 2444 16259 2746 16310
rect 2270 16258 2746 16259
rect 2798 16258 2813 16310
rect 2865 16258 2880 16310
rect 2932 16258 2946 16310
rect 2998 16258 3012 16310
rect 3064 16258 3078 16310
rect 3130 16258 3144 16310
rect 3196 16258 3210 16310
rect 3262 16258 3276 16310
rect 3328 16258 3342 16310
rect 3394 16258 3408 16310
rect 3460 16258 3474 16310
rect 3526 16258 3540 16310
rect 3592 16258 3606 16310
rect 3658 16258 3672 16310
rect 3724 16258 3738 16310
rect 3790 16258 3804 16310
rect 3856 16258 3870 16310
rect 3922 16258 3936 16310
rect 3988 16258 4002 16310
rect 4054 16258 4068 16310
rect 4120 16258 4134 16310
rect 4186 16258 4200 16310
rect 4252 16258 4266 16310
rect 4318 16258 4332 16310
rect 4384 16258 4398 16310
rect 4450 16258 4464 16310
rect 4516 16258 5116 16310
rect 5168 16258 5182 16310
rect 5234 16258 5248 16310
rect 5300 16258 5314 16310
rect 5366 16258 5380 16310
rect 5432 16258 5446 16310
rect 5498 16258 5512 16310
rect 5564 16258 5578 16310
rect 5630 16258 5644 16310
rect 5696 16258 5710 16310
rect 5762 16258 5776 16310
rect 5828 16258 5842 16310
rect 5894 16258 5908 16310
rect 5960 16258 5974 16310
rect 6026 16258 6040 16310
rect 6092 16258 6106 16310
rect 6158 16258 6172 16310
rect 6224 16258 6238 16310
rect 6290 16258 6304 16310
rect 6356 16258 6370 16310
rect 6422 16258 6436 16310
rect 6488 16258 6501 16310
rect 6553 16258 6566 16310
rect 6618 16258 6631 16310
rect 6683 16258 6696 16310
rect 6748 16258 6761 16310
rect 6813 16258 6826 16310
rect 6878 16258 6891 16310
rect 6943 16258 6956 16310
rect 7008 16258 7021 16310
rect 7073 16258 7086 16310
rect 7138 16258 7151 16310
rect 7203 16258 7216 16310
rect 7268 16258 7281 16310
rect 7333 16258 7346 16310
rect 7398 16258 7411 16310
rect 7463 16258 7476 16310
rect 7528 16258 7541 16310
rect 7593 16258 7606 16310
rect 7658 16258 7671 16310
rect 7723 16258 7736 16310
rect 7788 16258 7801 16310
rect 7853 16259 8047 16310
rect 8099 16259 8169 16311
rect 8221 16259 8222 16311
rect 7853 16258 8222 16259
rect 2270 16244 8222 16258
rect 2322 16192 2392 16244
rect 2444 16192 2746 16244
rect 2798 16192 2813 16244
rect 2865 16192 2880 16244
rect 2932 16192 2946 16244
rect 2998 16192 3012 16244
rect 3064 16192 3078 16244
rect 3130 16192 3144 16244
rect 3196 16192 3210 16244
rect 3262 16192 3276 16244
rect 3328 16192 3342 16244
rect 3394 16192 3408 16244
rect 3460 16192 3474 16244
rect 3526 16192 3540 16244
rect 3592 16192 3606 16244
rect 3658 16192 3672 16244
rect 3724 16192 3738 16244
rect 3790 16192 3804 16244
rect 3856 16192 3870 16244
rect 3922 16192 3936 16244
rect 3988 16192 4002 16244
rect 4054 16192 4068 16244
rect 4120 16192 4134 16244
rect 4186 16192 4200 16244
rect 4252 16192 4266 16244
rect 4318 16192 4332 16244
rect 4384 16192 4398 16244
rect 4450 16192 4464 16244
rect 4516 16192 5116 16244
rect 5168 16192 5182 16244
rect 5234 16192 5248 16244
rect 5300 16192 5314 16244
rect 5366 16192 5380 16244
rect 5432 16192 5446 16244
rect 5498 16192 5512 16244
rect 5564 16192 5578 16244
rect 5630 16192 5644 16244
rect 5696 16192 5710 16244
rect 5762 16192 5776 16244
rect 5828 16192 5842 16244
rect 5894 16192 5908 16244
rect 5960 16192 5974 16244
rect 6026 16192 6040 16244
rect 6092 16192 6106 16244
rect 6158 16192 6172 16244
rect 6224 16192 6238 16244
rect 6290 16192 6304 16244
rect 6356 16192 6370 16244
rect 6422 16192 6436 16244
rect 6488 16192 6501 16244
rect 6553 16192 6566 16244
rect 6618 16192 6631 16244
rect 6683 16192 6696 16244
rect 6748 16192 6761 16244
rect 6813 16192 6826 16244
rect 6878 16192 6891 16244
rect 6943 16192 6956 16244
rect 7008 16192 7021 16244
rect 7073 16192 7086 16244
rect 7138 16192 7151 16244
rect 7203 16192 7216 16244
rect 7268 16192 7281 16244
rect 7333 16192 7346 16244
rect 7398 16192 7411 16244
rect 7463 16192 7476 16244
rect 7528 16192 7541 16244
rect 7593 16192 7606 16244
rect 7658 16192 7671 16244
rect 7723 16192 7736 16244
rect 7788 16192 7801 16244
rect 7853 16192 8047 16244
rect 8099 16192 8169 16244
rect 8221 16192 8222 16244
rect 2270 16178 8222 16192
rect 2270 16177 2746 16178
rect 2322 16125 2392 16177
rect 2444 16126 2746 16177
rect 2798 16126 2813 16178
rect 2865 16126 2880 16178
rect 2932 16126 2946 16178
rect 2998 16126 3012 16178
rect 3064 16126 3078 16178
rect 3130 16126 3144 16178
rect 3196 16126 3210 16178
rect 3262 16126 3276 16178
rect 3328 16126 3342 16178
rect 3394 16126 3408 16178
rect 3460 16126 3474 16178
rect 3526 16126 3540 16178
rect 3592 16126 3606 16178
rect 3658 16126 3672 16178
rect 3724 16126 3738 16178
rect 3790 16126 3804 16178
rect 3856 16126 3870 16178
rect 3922 16126 3936 16178
rect 3988 16126 4002 16178
rect 4054 16126 4068 16178
rect 4120 16126 4134 16178
rect 4186 16126 4200 16178
rect 4252 16126 4266 16178
rect 4318 16126 4332 16178
rect 4384 16126 4398 16178
rect 4450 16126 4464 16178
rect 4516 16126 5116 16178
rect 5168 16126 5182 16178
rect 5234 16126 5248 16178
rect 5300 16126 5314 16178
rect 5366 16126 5380 16178
rect 5432 16126 5446 16178
rect 5498 16126 5512 16178
rect 5564 16126 5578 16178
rect 5630 16126 5644 16178
rect 5696 16126 5710 16178
rect 5762 16126 5776 16178
rect 5828 16126 5842 16178
rect 5894 16126 5908 16178
rect 5960 16126 5974 16178
rect 6026 16126 6040 16178
rect 6092 16126 6106 16178
rect 6158 16126 6172 16178
rect 6224 16126 6238 16178
rect 6290 16126 6304 16178
rect 6356 16126 6370 16178
rect 6422 16126 6436 16178
rect 6488 16126 6501 16178
rect 6553 16126 6566 16178
rect 6618 16126 6631 16178
rect 6683 16126 6696 16178
rect 6748 16126 6761 16178
rect 6813 16126 6826 16178
rect 6878 16126 6891 16178
rect 6943 16126 6956 16178
rect 7008 16126 7021 16178
rect 7073 16126 7086 16178
rect 7138 16126 7151 16178
rect 7203 16126 7216 16178
rect 7268 16126 7281 16178
rect 7333 16126 7346 16178
rect 7398 16126 7411 16178
rect 7463 16126 7476 16178
rect 7528 16126 7541 16178
rect 7593 16126 7606 16178
rect 7658 16126 7671 16178
rect 7723 16126 7736 16178
rect 7788 16126 7801 16178
rect 7853 16177 8222 16178
rect 7853 16126 8047 16177
rect 2444 16125 8047 16126
rect 8099 16125 8169 16177
rect 8221 16125 8222 16177
rect 2270 16112 8222 16125
rect 2270 16110 2746 16112
rect 2322 16058 2392 16110
rect 2444 16060 2746 16110
rect 2798 16060 2813 16112
rect 2865 16060 2880 16112
rect 2932 16060 2946 16112
rect 2998 16060 3012 16112
rect 3064 16060 3078 16112
rect 3130 16060 3144 16112
rect 3196 16060 3210 16112
rect 3262 16060 3276 16112
rect 3328 16060 3342 16112
rect 3394 16060 3408 16112
rect 3460 16060 3474 16112
rect 3526 16060 3540 16112
rect 3592 16060 3606 16112
rect 3658 16060 3672 16112
rect 3724 16060 3738 16112
rect 3790 16060 3804 16112
rect 3856 16060 3870 16112
rect 3922 16060 3936 16112
rect 3988 16060 4002 16112
rect 4054 16060 4068 16112
rect 4120 16060 4134 16112
rect 4186 16060 4200 16112
rect 4252 16060 4266 16112
rect 4318 16060 4332 16112
rect 4384 16060 4398 16112
rect 4450 16060 4464 16112
rect 4516 16060 5116 16112
rect 5168 16060 5182 16112
rect 5234 16060 5248 16112
rect 5300 16060 5314 16112
rect 5366 16060 5380 16112
rect 5432 16060 5446 16112
rect 5498 16060 5512 16112
rect 5564 16060 5578 16112
rect 5630 16060 5644 16112
rect 5696 16060 5710 16112
rect 5762 16060 5776 16112
rect 5828 16060 5842 16112
rect 5894 16060 5908 16112
rect 5960 16060 5974 16112
rect 6026 16060 6040 16112
rect 6092 16060 6106 16112
rect 6158 16060 6172 16112
rect 6224 16060 6238 16112
rect 6290 16060 6304 16112
rect 6356 16060 6370 16112
rect 6422 16060 6436 16112
rect 6488 16060 6501 16112
rect 6553 16060 6566 16112
rect 6618 16060 6631 16112
rect 6683 16060 6696 16112
rect 6748 16060 6761 16112
rect 6813 16060 6826 16112
rect 6878 16060 6891 16112
rect 6943 16060 6956 16112
rect 7008 16060 7021 16112
rect 7073 16060 7086 16112
rect 7138 16060 7151 16112
rect 7203 16060 7216 16112
rect 7268 16060 7281 16112
rect 7333 16060 7346 16112
rect 7398 16060 7411 16112
rect 7463 16060 7476 16112
rect 7528 16060 7541 16112
rect 7593 16060 7606 16112
rect 7658 16060 7671 16112
rect 7723 16060 7736 16112
rect 7788 16060 7801 16112
rect 7853 16110 8222 16112
rect 7853 16060 8047 16110
rect 2444 16058 8047 16060
rect 8099 16058 8169 16110
rect 8221 16058 8222 16110
rect 2270 16046 8222 16058
rect 2270 16043 2746 16046
rect 2322 15991 2392 16043
rect 2444 15994 2746 16043
rect 2798 15994 2813 16046
rect 2865 15994 2880 16046
rect 2932 15994 2946 16046
rect 2998 15994 3012 16046
rect 3064 15994 3078 16046
rect 3130 15994 3144 16046
rect 3196 15994 3210 16046
rect 3262 15994 3276 16046
rect 3328 15994 3342 16046
rect 3394 15994 3408 16046
rect 3460 15994 3474 16046
rect 3526 15994 3540 16046
rect 3592 15994 3606 16046
rect 3658 15994 3672 16046
rect 3724 15994 3738 16046
rect 3790 15994 3804 16046
rect 3856 15994 3870 16046
rect 3922 15994 3936 16046
rect 3988 15994 4002 16046
rect 4054 15994 4068 16046
rect 4120 15994 4134 16046
rect 4186 15994 4200 16046
rect 4252 15994 4266 16046
rect 4318 15994 4332 16046
rect 4384 15994 4398 16046
rect 4450 15994 4464 16046
rect 4516 15994 5116 16046
rect 5168 15994 5182 16046
rect 5234 15994 5248 16046
rect 5300 15994 5314 16046
rect 5366 15994 5380 16046
rect 5432 15994 5446 16046
rect 5498 15994 5512 16046
rect 5564 15994 5578 16046
rect 5630 15994 5644 16046
rect 5696 15994 5710 16046
rect 5762 15994 5776 16046
rect 5828 15994 5842 16046
rect 5894 15994 5908 16046
rect 5960 15994 5974 16046
rect 6026 15994 6040 16046
rect 6092 15994 6106 16046
rect 6158 15994 6172 16046
rect 6224 15994 6238 16046
rect 6290 15994 6304 16046
rect 6356 15994 6370 16046
rect 6422 15994 6436 16046
rect 6488 15994 6501 16046
rect 6553 15994 6566 16046
rect 6618 15994 6631 16046
rect 6683 15994 6696 16046
rect 6748 15994 6761 16046
rect 6813 15994 6826 16046
rect 6878 15994 6891 16046
rect 6943 15994 6956 16046
rect 7008 15994 7021 16046
rect 7073 15994 7086 16046
rect 7138 15994 7151 16046
rect 7203 15994 7216 16046
rect 7268 15994 7281 16046
rect 7333 15994 7346 16046
rect 7398 15994 7411 16046
rect 7463 15994 7476 16046
rect 7528 15994 7541 16046
rect 7593 15994 7606 16046
rect 7658 15994 7671 16046
rect 7723 15994 7736 16046
rect 7788 15994 7801 16046
rect 7853 16043 8222 16046
rect 7853 15994 8047 16043
rect 2444 15991 8047 15994
rect 8099 15991 8169 16043
rect 8221 15991 8222 16043
rect 2270 15985 8222 15991
rect 2270 15456 8222 15462
rect 2322 15404 2392 15456
rect 2444 15452 5613 15456
rect 5669 15452 5696 15456
rect 2444 15404 2824 15452
rect 2270 15400 2824 15404
rect 2876 15400 2890 15452
rect 2942 15400 3378 15452
rect 3430 15400 3444 15452
rect 3496 15400 3932 15452
rect 3984 15400 3998 15452
rect 4050 15400 4486 15452
rect 4538 15400 4552 15452
rect 4604 15400 5040 15452
rect 5092 15400 5106 15452
rect 5158 15400 5594 15452
rect 5752 15400 5779 15456
rect 5835 15400 5861 15456
rect 5917 15400 5943 15456
rect 5999 15400 6025 15456
rect 6081 15400 6107 15456
rect 6163 15452 6189 15456
rect 6245 15452 6271 15456
rect 6266 15400 6271 15452
rect 6327 15400 6353 15456
rect 6409 15400 6435 15456
rect 6491 15400 6517 15456
rect 6573 15400 6599 15456
rect 6655 15400 6681 15456
rect 6737 15452 6763 15456
rect 6819 15452 6845 15456
rect 6754 15400 6763 15452
rect 6820 15400 6845 15452
rect 6901 15400 6927 15456
rect 6983 15400 7009 15456
rect 7065 15400 7091 15456
rect 7147 15400 7173 15456
rect 7229 15400 7255 15456
rect 7311 15452 7337 15456
rect 7311 15400 7322 15452
rect 7393 15400 7419 15456
rect 7475 15400 7501 15456
rect 7557 15400 7583 15456
rect 7639 15400 7665 15456
rect 7721 15400 7747 15456
rect 7803 15452 7829 15456
rect 7885 15452 7911 15456
rect 7803 15400 7810 15452
rect 7967 15400 7993 15456
rect 8049 15400 8075 15404
rect 8131 15400 8157 15456
rect 8221 15404 8222 15456
rect 8213 15400 8222 15404
rect 2270 15387 8222 15400
rect 2322 15335 2392 15387
rect 2444 15383 8047 15387
rect 2444 15335 2824 15383
rect 2270 15331 2824 15335
rect 2876 15331 2890 15383
rect 2942 15331 3378 15383
rect 3430 15331 3444 15383
rect 3496 15331 3932 15383
rect 3984 15331 3998 15383
rect 4050 15331 4486 15383
rect 4538 15331 4552 15383
rect 4604 15331 5040 15383
rect 5092 15331 5106 15383
rect 5158 15331 5594 15383
rect 5646 15376 5660 15383
rect 5712 15376 6148 15383
rect 6200 15376 6214 15383
rect 6266 15376 6702 15383
rect 6754 15376 6768 15383
rect 6820 15376 7256 15383
rect 7308 15376 7322 15383
rect 7374 15376 7810 15383
rect 7862 15376 7876 15383
rect 7928 15376 8047 15383
rect 8099 15376 8169 15387
rect 2270 15320 5613 15331
rect 5669 15320 5696 15331
rect 5752 15320 5779 15376
rect 5835 15320 5861 15376
rect 5917 15320 5943 15376
rect 5999 15320 6025 15376
rect 6081 15320 6107 15376
rect 6266 15331 6271 15376
rect 6163 15320 6189 15331
rect 6245 15320 6271 15331
rect 6327 15320 6353 15376
rect 6409 15320 6435 15376
rect 6491 15320 6517 15376
rect 6573 15320 6599 15376
rect 6655 15320 6681 15376
rect 6754 15331 6763 15376
rect 6820 15331 6845 15376
rect 6737 15320 6763 15331
rect 6819 15320 6845 15331
rect 6901 15320 6927 15376
rect 6983 15320 7009 15376
rect 7065 15320 7091 15376
rect 7147 15320 7173 15376
rect 7229 15320 7255 15376
rect 7311 15331 7322 15376
rect 7311 15320 7337 15331
rect 7393 15320 7419 15376
rect 7475 15320 7501 15376
rect 7557 15320 7583 15376
rect 7639 15320 7665 15376
rect 7721 15320 7747 15376
rect 7803 15331 7810 15376
rect 7803 15320 7829 15331
rect 7885 15320 7911 15331
rect 7967 15320 7993 15376
rect 8049 15320 8075 15335
rect 8131 15320 8157 15376
rect 8221 15335 8222 15387
rect 8213 15320 8222 15335
rect 2270 15318 8222 15320
rect 2322 15266 2392 15318
rect 2444 15314 8047 15318
rect 2444 15266 2824 15314
rect 2270 15262 2824 15266
rect 2876 15262 2890 15314
rect 2942 15262 3378 15314
rect 3430 15262 3444 15314
rect 3496 15262 3932 15314
rect 3984 15262 3998 15314
rect 4050 15262 4486 15314
rect 4538 15262 4552 15314
rect 4604 15262 5040 15314
rect 5092 15262 5106 15314
rect 5158 15262 5594 15314
rect 5646 15296 5660 15314
rect 5712 15296 6148 15314
rect 6200 15296 6214 15314
rect 6266 15296 6702 15314
rect 6754 15296 6768 15314
rect 6820 15296 7256 15314
rect 7308 15296 7322 15314
rect 7374 15296 7810 15314
rect 7862 15296 7876 15314
rect 7928 15296 8047 15314
rect 8099 15296 8169 15318
rect 2270 15249 5613 15262
rect 2322 15197 2392 15249
rect 2444 15245 5613 15249
rect 5669 15245 5696 15262
rect 2444 15197 2824 15245
rect 2270 15193 2824 15197
rect 2876 15193 2890 15245
rect 2942 15193 3378 15245
rect 3430 15193 3444 15245
rect 3496 15193 3932 15245
rect 3984 15193 3998 15245
rect 4050 15193 4486 15245
rect 4538 15193 4552 15245
rect 4604 15193 5040 15245
rect 5092 15193 5106 15245
rect 5158 15193 5594 15245
rect 5752 15240 5779 15296
rect 5835 15240 5861 15296
rect 5917 15240 5943 15296
rect 5999 15240 6025 15296
rect 6081 15240 6107 15296
rect 6266 15262 6271 15296
rect 6163 15245 6189 15262
rect 6245 15245 6271 15262
rect 6266 15240 6271 15245
rect 6327 15240 6353 15296
rect 6409 15240 6435 15296
rect 6491 15240 6517 15296
rect 6573 15240 6599 15296
rect 6655 15240 6681 15296
rect 6754 15262 6763 15296
rect 6820 15262 6845 15296
rect 6737 15245 6763 15262
rect 6819 15245 6845 15262
rect 6754 15240 6763 15245
rect 6820 15240 6845 15245
rect 6901 15240 6927 15296
rect 6983 15240 7009 15296
rect 7065 15240 7091 15296
rect 7147 15240 7173 15296
rect 7229 15240 7255 15296
rect 7311 15262 7322 15296
rect 7311 15245 7337 15262
rect 7311 15240 7322 15245
rect 7393 15240 7419 15296
rect 7475 15240 7501 15296
rect 7557 15240 7583 15296
rect 7639 15240 7665 15296
rect 7721 15240 7747 15296
rect 7803 15262 7810 15296
rect 7803 15245 7829 15262
rect 7885 15245 7911 15262
rect 7803 15240 7810 15245
rect 7967 15240 7993 15296
rect 8049 15249 8075 15266
rect 8131 15240 8157 15296
rect 8221 15266 8222 15318
rect 8213 15249 8222 15266
rect 5646 15216 5660 15240
rect 5712 15216 6148 15240
rect 6200 15216 6214 15240
rect 6266 15216 6702 15240
rect 6754 15216 6768 15240
rect 6820 15216 7256 15240
rect 7308 15216 7322 15240
rect 7374 15216 7810 15240
rect 7862 15216 7876 15240
rect 7928 15216 8047 15240
rect 8099 15216 8169 15240
rect 2270 15180 5613 15193
rect 2322 15128 2392 15180
rect 2444 15176 5613 15180
rect 5669 15176 5696 15193
rect 2444 15128 2824 15176
rect 2270 15124 2824 15128
rect 2876 15124 2890 15176
rect 2942 15124 3378 15176
rect 3430 15124 3444 15176
rect 3496 15124 3932 15176
rect 3984 15124 3998 15176
rect 4050 15124 4486 15176
rect 4538 15124 4552 15176
rect 4604 15124 5040 15176
rect 5092 15124 5106 15176
rect 5158 15124 5594 15176
rect 5752 15160 5779 15216
rect 5835 15160 5861 15216
rect 5917 15160 5943 15216
rect 5999 15160 6025 15216
rect 6081 15160 6107 15216
rect 6266 15193 6271 15216
rect 6163 15176 6189 15193
rect 6245 15176 6271 15193
rect 6266 15160 6271 15176
rect 6327 15160 6353 15216
rect 6409 15160 6435 15216
rect 6491 15160 6517 15216
rect 6573 15160 6599 15216
rect 6655 15160 6681 15216
rect 6754 15193 6763 15216
rect 6820 15193 6845 15216
rect 6737 15176 6763 15193
rect 6819 15176 6845 15193
rect 6754 15160 6763 15176
rect 6820 15160 6845 15176
rect 6901 15160 6927 15216
rect 6983 15160 7009 15216
rect 7065 15160 7091 15216
rect 7147 15160 7173 15216
rect 7229 15160 7255 15216
rect 7311 15193 7322 15216
rect 7311 15176 7337 15193
rect 7311 15160 7322 15176
rect 7393 15160 7419 15216
rect 7475 15160 7501 15216
rect 7557 15160 7583 15216
rect 7639 15160 7665 15216
rect 7721 15160 7747 15216
rect 7803 15193 7810 15216
rect 7803 15176 7829 15193
rect 7885 15176 7911 15193
rect 7803 15160 7810 15176
rect 7967 15160 7993 15216
rect 8049 15180 8075 15197
rect 8131 15160 8157 15216
rect 8221 15197 8222 15249
rect 8213 15180 8222 15197
rect 5646 15136 5660 15160
rect 5712 15136 6148 15160
rect 6200 15136 6214 15160
rect 6266 15136 6702 15160
rect 6754 15136 6768 15160
rect 6820 15136 7256 15160
rect 7308 15136 7322 15160
rect 7374 15136 7810 15160
rect 7862 15136 7876 15160
rect 7928 15136 8047 15160
rect 8099 15136 8169 15160
rect 2270 15110 5613 15124
rect 2322 15058 2392 15110
rect 2444 15107 5613 15110
rect 5669 15107 5696 15124
rect 2444 15058 2824 15107
rect 2270 15055 2824 15058
rect 2876 15055 2890 15107
rect 2942 15055 3378 15107
rect 3430 15055 3444 15107
rect 3496 15055 3932 15107
rect 3984 15055 3998 15107
rect 4050 15055 4486 15107
rect 4538 15055 4552 15107
rect 4604 15055 5040 15107
rect 5092 15055 5106 15107
rect 5158 15055 5594 15107
rect 5752 15080 5779 15136
rect 5835 15080 5861 15136
rect 5917 15080 5943 15136
rect 5999 15080 6025 15136
rect 6081 15080 6107 15136
rect 6266 15124 6271 15136
rect 6163 15107 6189 15124
rect 6245 15107 6271 15124
rect 6266 15080 6271 15107
rect 6327 15080 6353 15136
rect 6409 15080 6435 15136
rect 6491 15080 6517 15136
rect 6573 15080 6599 15136
rect 6655 15080 6681 15136
rect 6754 15124 6763 15136
rect 6820 15124 6845 15136
rect 6737 15107 6763 15124
rect 6819 15107 6845 15124
rect 6754 15080 6763 15107
rect 6820 15080 6845 15107
rect 6901 15080 6927 15136
rect 6983 15080 7009 15136
rect 7065 15080 7091 15136
rect 7147 15080 7173 15136
rect 7229 15080 7255 15136
rect 7311 15124 7322 15136
rect 7311 15107 7337 15124
rect 7311 15080 7322 15107
rect 7393 15080 7419 15136
rect 7475 15080 7501 15136
rect 7557 15080 7583 15136
rect 7639 15080 7665 15136
rect 7721 15080 7747 15136
rect 7803 15124 7810 15136
rect 7803 15107 7829 15124
rect 7885 15107 7911 15124
rect 7803 15080 7810 15107
rect 7967 15080 7993 15136
rect 8049 15110 8075 15128
rect 8131 15080 8157 15136
rect 8221 15128 8222 15180
rect 8213 15110 8222 15128
rect 5646 15056 5660 15080
rect 5712 15056 6148 15080
rect 6200 15056 6214 15080
rect 6266 15056 6702 15080
rect 6754 15056 6768 15080
rect 6820 15056 7256 15080
rect 7308 15056 7322 15080
rect 7374 15056 7810 15080
rect 7862 15056 7876 15080
rect 7928 15058 8047 15080
rect 8099 15058 8169 15080
rect 8221 15058 8222 15110
rect 7928 15056 8222 15058
rect 2270 15040 5613 15055
rect 2322 14988 2392 15040
rect 2444 15038 5613 15040
rect 5669 15038 5696 15055
rect 2444 14988 2824 15038
rect 2270 14986 2824 14988
rect 2876 14986 2890 15038
rect 2942 14986 3378 15038
rect 3430 14986 3444 15038
rect 3496 14986 3932 15038
rect 3984 14986 3998 15038
rect 4050 14986 4486 15038
rect 4538 14986 4552 15038
rect 4604 14986 5040 15038
rect 5092 14986 5106 15038
rect 5158 14986 5594 15038
rect 5752 15000 5779 15056
rect 5835 15000 5861 15056
rect 5917 15000 5943 15056
rect 5999 15000 6025 15056
rect 6081 15000 6107 15056
rect 6266 15055 6271 15056
rect 6163 15038 6189 15055
rect 6245 15038 6271 15055
rect 6266 15000 6271 15038
rect 6327 15000 6353 15056
rect 6409 15000 6435 15056
rect 6491 15000 6517 15056
rect 6573 15000 6599 15056
rect 6655 15000 6681 15056
rect 6754 15055 6763 15056
rect 6820 15055 6845 15056
rect 6737 15038 6763 15055
rect 6819 15038 6845 15055
rect 6754 15000 6763 15038
rect 6820 15000 6845 15038
rect 6901 15000 6927 15056
rect 6983 15000 7009 15056
rect 7065 15000 7091 15056
rect 7147 15000 7173 15056
rect 7229 15000 7255 15056
rect 7311 15055 7322 15056
rect 7311 15038 7337 15055
rect 7311 15000 7322 15038
rect 7393 15000 7419 15056
rect 7475 15000 7501 15056
rect 7557 15000 7583 15056
rect 7639 15000 7665 15056
rect 7721 15000 7747 15056
rect 7803 15055 7810 15056
rect 7803 15038 7829 15055
rect 7885 15038 7911 15055
rect 7803 15000 7810 15038
rect 7967 15000 7993 15056
rect 8049 15040 8075 15056
rect 8131 15000 8157 15056
rect 8213 15040 8222 15056
rect 5646 14986 5660 15000
rect 5712 14986 6148 15000
rect 6200 14986 6214 15000
rect 6266 14986 6702 15000
rect 6754 14986 6768 15000
rect 6820 14986 7256 15000
rect 7308 14986 7322 15000
rect 7374 14986 7810 15000
rect 7862 14986 7876 15000
rect 7928 14988 8047 15000
rect 8099 14988 8169 15000
rect 8221 14988 8222 15040
rect 7928 14986 8222 14988
rect 2270 14976 8222 14986
rect 2270 14970 5613 14976
rect 2322 14918 2392 14970
rect 2444 14968 5613 14970
rect 5669 14968 5696 14976
rect 2444 14918 2824 14968
rect 2270 14916 2824 14918
rect 2876 14916 2890 14968
rect 2942 14916 3378 14968
rect 3430 14916 3444 14968
rect 3496 14916 3932 14968
rect 3984 14916 3998 14968
rect 4050 14916 4486 14968
rect 4538 14916 4552 14968
rect 4604 14916 5040 14968
rect 5092 14916 5106 14968
rect 5158 14916 5594 14968
rect 5752 14920 5779 14976
rect 5835 14920 5861 14976
rect 5917 14920 5943 14976
rect 5999 14920 6025 14976
rect 6081 14920 6107 14976
rect 6163 14968 6189 14976
rect 6245 14968 6271 14976
rect 6266 14920 6271 14968
rect 6327 14920 6353 14976
rect 6409 14920 6435 14976
rect 6491 14920 6517 14976
rect 6573 14920 6599 14976
rect 6655 14920 6681 14976
rect 6737 14968 6763 14976
rect 6819 14968 6845 14976
rect 6754 14920 6763 14968
rect 6820 14920 6845 14968
rect 6901 14920 6927 14976
rect 6983 14920 7009 14976
rect 7065 14920 7091 14976
rect 7147 14920 7173 14976
rect 7229 14920 7255 14976
rect 7311 14968 7337 14976
rect 7311 14920 7322 14968
rect 7393 14920 7419 14976
rect 7475 14920 7501 14976
rect 7557 14920 7583 14976
rect 7639 14920 7665 14976
rect 7721 14920 7747 14976
rect 7803 14968 7829 14976
rect 7885 14968 7911 14976
rect 7803 14920 7810 14968
rect 7967 14920 7993 14976
rect 8049 14970 8075 14976
rect 8131 14920 8157 14976
rect 8213 14970 8222 14976
rect 5646 14916 5660 14920
rect 5712 14916 6148 14920
rect 6200 14916 6214 14920
rect 6266 14916 6702 14920
rect 6754 14916 6768 14920
rect 6820 14916 7256 14920
rect 7308 14916 7322 14920
rect 7374 14916 7810 14920
rect 7862 14916 7876 14920
rect 7928 14918 8047 14920
rect 8099 14918 8169 14920
rect 8221 14918 8222 14970
rect 7928 14916 8222 14918
rect 2270 14900 8222 14916
rect 2322 14848 2392 14900
rect 2444 14898 8047 14900
rect 2444 14848 2824 14898
rect 2270 14846 2824 14848
rect 2876 14846 2890 14898
rect 2942 14846 3378 14898
rect 3430 14846 3444 14898
rect 3496 14846 3932 14898
rect 3984 14846 3998 14898
rect 4050 14846 4486 14898
rect 4538 14846 4552 14898
rect 4604 14846 5040 14898
rect 5092 14846 5106 14898
rect 5158 14846 5594 14898
rect 5646 14896 5660 14898
rect 5712 14896 6148 14898
rect 6200 14896 6214 14898
rect 6266 14896 6702 14898
rect 6754 14896 6768 14898
rect 6820 14896 7256 14898
rect 7308 14896 7322 14898
rect 7374 14896 7810 14898
rect 7862 14896 7876 14898
rect 7928 14896 8047 14898
rect 8099 14896 8169 14900
rect 2270 14840 5613 14846
rect 5669 14840 5696 14846
rect 5752 14840 5779 14896
rect 5835 14840 5861 14896
rect 5917 14840 5943 14896
rect 5999 14840 6025 14896
rect 6081 14840 6107 14896
rect 6266 14846 6271 14896
rect 6163 14840 6189 14846
rect 6245 14840 6271 14846
rect 6327 14840 6353 14896
rect 6409 14840 6435 14896
rect 6491 14840 6517 14896
rect 6573 14840 6599 14896
rect 6655 14840 6681 14896
rect 6754 14846 6763 14896
rect 6820 14846 6845 14896
rect 6737 14840 6763 14846
rect 6819 14840 6845 14846
rect 6901 14840 6927 14896
rect 6983 14840 7009 14896
rect 7065 14840 7091 14896
rect 7147 14840 7173 14896
rect 7229 14840 7255 14896
rect 7311 14846 7322 14896
rect 7311 14840 7337 14846
rect 7393 14840 7419 14896
rect 7475 14840 7501 14896
rect 7557 14840 7583 14896
rect 7639 14840 7665 14896
rect 7721 14840 7747 14896
rect 7803 14846 7810 14896
rect 7803 14840 7829 14846
rect 7885 14840 7911 14846
rect 7967 14840 7993 14896
rect 8049 14840 8075 14848
rect 8131 14840 8157 14896
rect 8221 14848 8222 14900
rect 8213 14840 8222 14848
rect 2724 14719 7651 14720
rect 2724 14663 2733 14719
rect 2789 14663 2814 14719
rect 2870 14663 2895 14719
rect 2951 14663 2976 14719
rect 3032 14663 3057 14719
rect 3113 14714 3138 14719
rect 3194 14714 3219 14719
rect 3275 14663 3300 14719
rect 3356 14663 3381 14719
rect 3437 14663 3462 14719
rect 3518 14663 3543 14719
rect 3599 14663 3624 14719
rect 3680 14714 3705 14719
rect 3761 14714 3786 14719
rect 3773 14663 3786 14714
rect 3842 14663 3867 14719
rect 3923 14663 3948 14719
rect 4004 14663 4029 14719
rect 4085 14663 4110 14719
rect 4166 14663 4191 14719
rect 4247 14714 4272 14719
rect 4261 14663 4272 14714
rect 4328 14663 4353 14719
rect 4409 14663 4434 14719
rect 4490 14663 4515 14719
rect 4571 14663 4596 14719
rect 4652 14663 4677 14719
rect 4733 14663 4758 14719
rect 4814 14714 4839 14719
rect 2724 14662 3101 14663
rect 3153 14662 3167 14663
rect 3219 14662 3655 14663
rect 3707 14662 3721 14663
rect 3773 14662 4209 14663
rect 4261 14662 4275 14663
rect 4327 14662 4763 14663
rect 4815 14662 4829 14714
rect 4895 14663 4920 14719
rect 4976 14663 5001 14719
rect 5057 14663 5082 14719
rect 5138 14663 5163 14719
rect 4881 14662 5163 14663
rect 2724 14645 5163 14662
rect 2724 14639 3101 14645
rect 3153 14639 3167 14645
rect 3219 14639 3655 14645
rect 3707 14639 3721 14645
rect 3773 14639 4209 14645
rect 4261 14639 4275 14645
rect 4327 14639 4763 14645
rect 2724 14583 2733 14639
rect 2789 14583 2814 14639
rect 2870 14583 2895 14639
rect 2951 14583 2976 14639
rect 3032 14583 3057 14639
rect 3113 14583 3138 14593
rect 3194 14583 3219 14593
rect 3275 14583 3300 14639
rect 3356 14583 3381 14639
rect 3437 14583 3462 14639
rect 3518 14583 3543 14639
rect 3599 14583 3624 14639
rect 3773 14593 3786 14639
rect 3680 14583 3705 14593
rect 3761 14583 3786 14593
rect 3842 14583 3867 14639
rect 3923 14583 3948 14639
rect 4004 14583 4029 14639
rect 4085 14583 4110 14639
rect 4166 14583 4191 14639
rect 4261 14593 4272 14639
rect 4247 14583 4272 14593
rect 4328 14583 4353 14639
rect 4409 14583 4434 14639
rect 4490 14583 4515 14639
rect 4571 14583 4596 14639
rect 4652 14583 4677 14639
rect 4733 14583 4758 14639
rect 4815 14593 4829 14645
rect 4881 14639 5163 14645
rect 4814 14583 4839 14593
rect 4895 14583 4920 14639
rect 4976 14583 5001 14639
rect 5057 14583 5082 14639
rect 5138 14583 5163 14639
rect 2724 14576 5163 14583
rect 2724 14559 3101 14576
rect 3153 14559 3167 14576
rect 3219 14559 3655 14576
rect 3707 14559 3721 14576
rect 3773 14559 4209 14576
rect 4261 14559 4275 14576
rect 4327 14559 4763 14576
rect 2724 14503 2733 14559
rect 2789 14503 2814 14559
rect 2870 14503 2895 14559
rect 2951 14503 2976 14559
rect 3032 14503 3057 14559
rect 3113 14507 3138 14524
rect 3194 14507 3219 14524
rect 3275 14503 3300 14559
rect 3356 14503 3381 14559
rect 3437 14503 3462 14559
rect 3518 14503 3543 14559
rect 3599 14503 3624 14559
rect 3773 14524 3786 14559
rect 3680 14507 3705 14524
rect 3761 14507 3786 14524
rect 3773 14503 3786 14507
rect 3842 14503 3867 14559
rect 3923 14503 3948 14559
rect 4004 14503 4029 14559
rect 4085 14503 4110 14559
rect 4166 14503 4191 14559
rect 4261 14524 4272 14559
rect 4247 14507 4272 14524
rect 4261 14503 4272 14507
rect 4328 14503 4353 14559
rect 4409 14503 4434 14559
rect 4490 14503 4515 14559
rect 4571 14503 4596 14559
rect 4652 14503 4677 14559
rect 4733 14503 4758 14559
rect 4815 14524 4829 14576
rect 4881 14559 5163 14576
rect 4814 14507 4839 14524
rect 2724 14479 3101 14503
rect 3153 14479 3167 14503
rect 3219 14479 3655 14503
rect 3707 14479 3721 14503
rect 3773 14479 4209 14503
rect 4261 14479 4275 14503
rect 4327 14479 4763 14503
rect 2724 14423 2733 14479
rect 2789 14423 2814 14479
rect 2870 14423 2895 14479
rect 2951 14423 2976 14479
rect 3032 14423 3057 14479
rect 3113 14438 3138 14455
rect 3194 14438 3219 14455
rect 3275 14423 3300 14479
rect 3356 14423 3381 14479
rect 3437 14423 3462 14479
rect 3518 14423 3543 14479
rect 3599 14423 3624 14479
rect 3773 14455 3786 14479
rect 3680 14438 3705 14455
rect 3761 14438 3786 14455
rect 3773 14423 3786 14438
rect 3842 14423 3867 14479
rect 3923 14423 3948 14479
rect 4004 14423 4029 14479
rect 4085 14423 4110 14479
rect 4166 14423 4191 14479
rect 4261 14455 4272 14479
rect 4247 14438 4272 14455
rect 4261 14423 4272 14438
rect 4328 14423 4353 14479
rect 4409 14423 4434 14479
rect 4490 14423 4515 14479
rect 4571 14423 4596 14479
rect 4652 14423 4677 14479
rect 4733 14423 4758 14479
rect 4815 14455 4829 14507
rect 4895 14503 4920 14559
rect 4976 14503 5001 14559
rect 5057 14503 5082 14559
rect 5138 14503 5163 14559
rect 4881 14479 5163 14503
rect 4814 14438 4839 14455
rect 2724 14399 3101 14423
rect 3153 14399 3167 14423
rect 3219 14399 3655 14423
rect 3707 14399 3721 14423
rect 3773 14399 4209 14423
rect 4261 14399 4275 14423
rect 4327 14399 4763 14423
rect 2724 14343 2733 14399
rect 2789 14343 2814 14399
rect 2870 14343 2895 14399
rect 2951 14343 2976 14399
rect 3032 14343 3057 14399
rect 3113 14368 3138 14386
rect 3194 14368 3219 14386
rect 3275 14343 3300 14399
rect 3356 14343 3381 14399
rect 3437 14343 3462 14399
rect 3518 14343 3543 14399
rect 3599 14343 3624 14399
rect 3773 14386 3786 14399
rect 3680 14368 3705 14386
rect 3761 14368 3786 14386
rect 3773 14343 3786 14368
rect 3842 14343 3867 14399
rect 3923 14343 3948 14399
rect 4004 14343 4029 14399
rect 4085 14343 4110 14399
rect 4166 14343 4191 14399
rect 4261 14386 4272 14399
rect 4247 14368 4272 14386
rect 4261 14343 4272 14368
rect 4328 14343 4353 14399
rect 4409 14343 4434 14399
rect 4490 14343 4515 14399
rect 4571 14343 4596 14399
rect 4652 14343 4677 14399
rect 4733 14343 4758 14399
rect 4815 14386 4829 14438
rect 4895 14423 4920 14479
rect 4976 14423 5001 14479
rect 5057 14423 5082 14479
rect 5138 14423 5163 14479
rect 4881 14399 5163 14423
rect 4814 14368 4839 14386
rect 2724 14319 3101 14343
rect 3153 14319 3167 14343
rect 3219 14319 3655 14343
rect 3707 14319 3721 14343
rect 3773 14319 4209 14343
rect 4261 14319 4275 14343
rect 4327 14319 4763 14343
rect 2724 14263 2733 14319
rect 2789 14263 2814 14319
rect 2870 14263 2895 14319
rect 2951 14263 2976 14319
rect 3032 14263 3057 14319
rect 3113 14298 3138 14316
rect 3194 14298 3219 14316
rect 3275 14263 3300 14319
rect 3356 14263 3381 14319
rect 3437 14263 3462 14319
rect 3518 14263 3543 14319
rect 3599 14263 3624 14319
rect 3773 14316 3786 14319
rect 3680 14298 3705 14316
rect 3761 14298 3786 14316
rect 3773 14263 3786 14298
rect 3842 14263 3867 14319
rect 3923 14263 3948 14319
rect 4004 14263 4029 14319
rect 4085 14263 4110 14319
rect 4166 14263 4191 14319
rect 4261 14316 4272 14319
rect 4247 14298 4272 14316
rect 4261 14263 4272 14298
rect 4328 14263 4353 14319
rect 4409 14263 4434 14319
rect 4490 14263 4515 14319
rect 4571 14263 4596 14319
rect 4652 14263 4677 14319
rect 4733 14263 4758 14319
rect 4815 14316 4829 14368
rect 4895 14343 4920 14399
rect 4976 14343 5001 14399
rect 5057 14343 5082 14399
rect 5138 14343 5163 14399
rect 4881 14319 5163 14343
rect 4814 14298 4839 14316
rect 2724 14246 3101 14263
rect 3153 14246 3167 14263
rect 3219 14246 3655 14263
rect 3707 14246 3721 14263
rect 3773 14246 4209 14263
rect 4261 14246 4275 14263
rect 4327 14246 4763 14263
rect 4815 14246 4829 14298
rect 4895 14263 4920 14319
rect 4976 14263 5001 14319
rect 5057 14263 5082 14319
rect 5138 14263 5163 14319
rect 4881 14246 5163 14263
rect 2724 14239 5163 14246
rect 2724 14183 2733 14239
rect 2789 14183 2814 14239
rect 2870 14183 2895 14239
rect 2951 14183 2976 14239
rect 3032 14183 3057 14239
rect 3113 14228 3138 14239
rect 3194 14228 3219 14239
rect 3275 14183 3300 14239
rect 3356 14183 3381 14239
rect 3437 14183 3462 14239
rect 3518 14183 3543 14239
rect 3599 14183 3624 14239
rect 3680 14228 3705 14239
rect 3761 14228 3786 14239
rect 3773 14183 3786 14228
rect 3842 14183 3867 14239
rect 3923 14183 3948 14239
rect 4004 14183 4029 14239
rect 4085 14183 4110 14239
rect 4166 14183 4191 14239
rect 4247 14228 4272 14239
rect 4261 14183 4272 14228
rect 4328 14183 4353 14239
rect 4409 14183 4434 14239
rect 4490 14183 4515 14239
rect 4571 14183 4596 14239
rect 4652 14183 4677 14239
rect 4733 14183 4758 14239
rect 4814 14228 4839 14239
rect 2724 14176 3101 14183
rect 3153 14176 3167 14183
rect 3219 14176 3655 14183
rect 3707 14176 3721 14183
rect 3773 14176 4209 14183
rect 4261 14176 4275 14183
rect 4327 14176 4763 14183
rect 4815 14176 4829 14228
rect 4895 14183 4920 14239
rect 4976 14183 5001 14239
rect 5057 14183 5082 14239
rect 5138 14183 5163 14239
rect 4881 14176 5163 14183
rect 2724 14159 5163 14176
rect 2724 14103 2733 14159
rect 2789 14103 2814 14159
rect 2870 14103 2895 14159
rect 2951 14103 2976 14159
rect 3032 14103 3057 14159
rect 3113 14158 3138 14159
rect 3194 14158 3219 14159
rect 3113 14103 3138 14106
rect 3194 14103 3219 14106
rect 3275 14103 3300 14159
rect 3356 14103 3381 14159
rect 3437 14103 3462 14159
rect 3518 14103 3543 14159
rect 3599 14103 3624 14159
rect 3680 14158 3705 14159
rect 3761 14158 3786 14159
rect 3773 14106 3786 14158
rect 3680 14103 3705 14106
rect 3761 14103 3786 14106
rect 3842 14103 3867 14159
rect 3923 14103 3948 14159
rect 4004 14103 4029 14159
rect 4085 14103 4110 14159
rect 4166 14103 4191 14159
rect 4247 14158 4272 14159
rect 4261 14106 4272 14158
rect 4247 14103 4272 14106
rect 4328 14103 4353 14159
rect 4409 14103 4434 14159
rect 4490 14103 4515 14159
rect 4571 14103 4596 14159
rect 4652 14103 4677 14159
rect 4733 14103 4758 14159
rect 4814 14158 4839 14159
rect 4815 14106 4829 14158
rect 4814 14103 4839 14106
rect 4895 14103 4920 14159
rect 4976 14103 5001 14159
rect 5057 14103 5082 14159
rect 5138 14103 5163 14159
rect 5299 14714 7651 14719
rect 5299 14662 5317 14714
rect 5369 14662 5383 14714
rect 5435 14662 5871 14714
rect 5923 14662 5937 14714
rect 5989 14662 6425 14714
rect 6477 14662 6491 14714
rect 6543 14662 6979 14714
rect 7031 14662 7045 14714
rect 7097 14662 7533 14714
rect 7585 14662 7599 14714
rect 5299 14645 7651 14662
rect 5299 14593 5317 14645
rect 5369 14593 5383 14645
rect 5435 14593 5871 14645
rect 5923 14593 5937 14645
rect 5989 14593 6425 14645
rect 6477 14593 6491 14645
rect 6543 14593 6979 14645
rect 7031 14593 7045 14645
rect 7097 14593 7533 14645
rect 7585 14593 7599 14645
rect 5299 14576 7651 14593
rect 5299 14524 5317 14576
rect 5369 14524 5383 14576
rect 5435 14524 5871 14576
rect 5923 14524 5937 14576
rect 5989 14524 6425 14576
rect 6477 14524 6491 14576
rect 6543 14524 6979 14576
rect 7031 14524 7045 14576
rect 7097 14524 7533 14576
rect 7585 14524 7599 14576
rect 5299 14507 7651 14524
rect 5299 14455 5317 14507
rect 5369 14455 5383 14507
rect 5435 14455 5871 14507
rect 5923 14455 5937 14507
rect 5989 14455 6425 14507
rect 6477 14455 6491 14507
rect 6543 14455 6979 14507
rect 7031 14455 7045 14507
rect 7097 14455 7533 14507
rect 7585 14455 7599 14507
rect 5299 14438 7651 14455
rect 5299 14386 5317 14438
rect 5369 14386 5383 14438
rect 5435 14386 5871 14438
rect 5923 14386 5937 14438
rect 5989 14386 6425 14438
rect 6477 14386 6491 14438
rect 6543 14386 6979 14438
rect 7031 14386 7045 14438
rect 7097 14386 7533 14438
rect 7585 14386 7599 14438
rect 5299 14368 7651 14386
rect 5299 14316 5317 14368
rect 5369 14316 5383 14368
rect 5435 14316 5871 14368
rect 5923 14316 5937 14368
rect 5989 14316 6425 14368
rect 6477 14316 6491 14368
rect 6543 14316 6979 14368
rect 7031 14316 7045 14368
rect 7097 14316 7533 14368
rect 7585 14316 7599 14368
rect 5299 14298 7651 14316
rect 5299 14246 5317 14298
rect 5369 14246 5383 14298
rect 5435 14246 5871 14298
rect 5923 14246 5937 14298
rect 5989 14246 6425 14298
rect 6477 14246 6491 14298
rect 6543 14246 6979 14298
rect 7031 14246 7045 14298
rect 7097 14246 7533 14298
rect 7585 14246 7599 14298
rect 5299 14228 7651 14246
rect 5299 14176 5317 14228
rect 5369 14176 5383 14228
rect 5435 14176 5871 14228
rect 5923 14176 5937 14228
rect 5989 14176 6425 14228
rect 6477 14176 6491 14228
rect 6543 14176 6979 14228
rect 7031 14176 7045 14228
rect 7097 14176 7533 14228
rect 7585 14176 7599 14228
rect 5299 14158 7651 14176
rect 5299 14106 5317 14158
rect 5369 14106 5383 14158
rect 5435 14106 5871 14158
rect 5923 14106 5937 14158
rect 5989 14106 6425 14158
rect 6477 14106 6491 14158
rect 6543 14106 6979 14158
rect 7031 14106 7045 14158
rect 7097 14106 7533 14158
rect 7585 14106 7599 14158
rect 5299 14103 7651 14106
rect 2724 14100 7651 14103
rect 2270 13456 8222 13462
rect 2322 13404 2392 13456
rect 2444 13452 5613 13456
rect 5669 13452 5696 13456
rect 2444 13404 2824 13452
rect 2270 13400 2824 13404
rect 2876 13400 2890 13452
rect 2942 13400 3378 13452
rect 3430 13400 3444 13452
rect 3496 13400 3932 13452
rect 3984 13400 3998 13452
rect 4050 13400 4486 13452
rect 4538 13400 4552 13452
rect 4604 13400 5040 13452
rect 5092 13400 5106 13452
rect 5158 13400 5594 13452
rect 5752 13400 5779 13456
rect 5835 13400 5861 13456
rect 5917 13400 5943 13456
rect 5999 13400 6025 13456
rect 6081 13400 6107 13456
rect 6163 13452 6189 13456
rect 6245 13452 6271 13456
rect 6266 13400 6271 13452
rect 6327 13400 6353 13456
rect 6409 13400 6435 13456
rect 6491 13400 6517 13456
rect 6573 13400 6599 13456
rect 6655 13400 6681 13456
rect 6737 13452 6763 13456
rect 6819 13452 6845 13456
rect 6754 13400 6763 13452
rect 6820 13400 6845 13452
rect 6901 13400 6927 13456
rect 6983 13400 7009 13456
rect 7065 13400 7091 13456
rect 7147 13400 7173 13456
rect 7229 13400 7255 13456
rect 7311 13452 7337 13456
rect 7311 13400 7322 13452
rect 7393 13400 7419 13456
rect 7475 13400 7501 13456
rect 7557 13400 7583 13456
rect 7639 13400 7665 13456
rect 7721 13400 7747 13456
rect 7803 13452 7829 13456
rect 7885 13452 7911 13456
rect 7803 13400 7810 13452
rect 7967 13400 7993 13456
rect 8049 13400 8075 13404
rect 8131 13400 8157 13456
rect 8221 13404 8222 13456
rect 8213 13400 8222 13404
rect 2270 13387 8222 13400
rect 2322 13335 2392 13387
rect 2444 13383 8047 13387
rect 2444 13335 2824 13383
rect 2270 13331 2824 13335
rect 2876 13331 2890 13383
rect 2942 13331 3378 13383
rect 3430 13331 3444 13383
rect 3496 13331 3932 13383
rect 3984 13331 3998 13383
rect 4050 13331 4486 13383
rect 4538 13331 4552 13383
rect 4604 13331 5040 13383
rect 5092 13331 5106 13383
rect 5158 13331 5594 13383
rect 5646 13376 5660 13383
rect 5712 13376 6148 13383
rect 6200 13376 6214 13383
rect 6266 13376 6702 13383
rect 6754 13376 6768 13383
rect 6820 13376 7256 13383
rect 7308 13376 7322 13383
rect 7374 13376 7810 13383
rect 7862 13376 7876 13383
rect 7928 13376 8047 13383
rect 8099 13376 8169 13387
rect 2270 13320 5613 13331
rect 5669 13320 5696 13331
rect 5752 13320 5779 13376
rect 5835 13320 5861 13376
rect 5917 13320 5943 13376
rect 5999 13320 6025 13376
rect 6081 13320 6107 13376
rect 6266 13331 6271 13376
rect 6163 13320 6189 13331
rect 6245 13320 6271 13331
rect 6327 13320 6353 13376
rect 6409 13320 6435 13376
rect 6491 13320 6517 13376
rect 6573 13320 6599 13376
rect 6655 13320 6681 13376
rect 6754 13331 6763 13376
rect 6820 13331 6845 13376
rect 6737 13320 6763 13331
rect 6819 13320 6845 13331
rect 6901 13320 6927 13376
rect 6983 13320 7009 13376
rect 7065 13320 7091 13376
rect 7147 13320 7173 13376
rect 7229 13320 7255 13376
rect 7311 13331 7322 13376
rect 7311 13320 7337 13331
rect 7393 13320 7419 13376
rect 7475 13320 7501 13376
rect 7557 13320 7583 13376
rect 7639 13320 7665 13376
rect 7721 13320 7747 13376
rect 7803 13331 7810 13376
rect 7803 13320 7829 13331
rect 7885 13320 7911 13331
rect 7967 13320 7993 13376
rect 8049 13320 8075 13335
rect 8131 13320 8157 13376
rect 8221 13335 8222 13387
rect 8213 13320 8222 13335
rect 2270 13318 8222 13320
rect 2322 13266 2392 13318
rect 2444 13314 8047 13318
rect 2444 13266 2824 13314
rect 2270 13262 2824 13266
rect 2876 13262 2890 13314
rect 2942 13262 3378 13314
rect 3430 13262 3444 13314
rect 3496 13262 3932 13314
rect 3984 13262 3998 13314
rect 4050 13262 4486 13314
rect 4538 13262 4552 13314
rect 4604 13262 5040 13314
rect 5092 13262 5106 13314
rect 5158 13262 5594 13314
rect 5646 13296 5660 13314
rect 5712 13296 6148 13314
rect 6200 13296 6214 13314
rect 6266 13296 6702 13314
rect 6754 13296 6768 13314
rect 6820 13296 7256 13314
rect 7308 13296 7322 13314
rect 7374 13296 7810 13314
rect 7862 13296 7876 13314
rect 7928 13296 8047 13314
rect 8099 13296 8169 13318
rect 2270 13249 5613 13262
rect 2322 13197 2392 13249
rect 2444 13245 5613 13249
rect 5669 13245 5696 13262
rect 2444 13197 2824 13245
rect 2270 13193 2824 13197
rect 2876 13193 2890 13245
rect 2942 13193 3378 13245
rect 3430 13193 3444 13245
rect 3496 13193 3932 13245
rect 3984 13193 3998 13245
rect 4050 13193 4486 13245
rect 4538 13193 4552 13245
rect 4604 13193 5040 13245
rect 5092 13193 5106 13245
rect 5158 13193 5594 13245
rect 5752 13240 5779 13296
rect 5835 13240 5861 13296
rect 5917 13240 5943 13296
rect 5999 13240 6025 13296
rect 6081 13240 6107 13296
rect 6266 13262 6271 13296
rect 6163 13245 6189 13262
rect 6245 13245 6271 13262
rect 6266 13240 6271 13245
rect 6327 13240 6353 13296
rect 6409 13240 6435 13296
rect 6491 13240 6517 13296
rect 6573 13240 6599 13296
rect 6655 13240 6681 13296
rect 6754 13262 6763 13296
rect 6820 13262 6845 13296
rect 6737 13245 6763 13262
rect 6819 13245 6845 13262
rect 6754 13240 6763 13245
rect 6820 13240 6845 13245
rect 6901 13240 6927 13296
rect 6983 13240 7009 13296
rect 7065 13240 7091 13296
rect 7147 13240 7173 13296
rect 7229 13240 7255 13296
rect 7311 13262 7322 13296
rect 7311 13245 7337 13262
rect 7311 13240 7322 13245
rect 7393 13240 7419 13296
rect 7475 13240 7501 13296
rect 7557 13240 7583 13296
rect 7639 13240 7665 13296
rect 7721 13240 7747 13296
rect 7803 13262 7810 13296
rect 7803 13245 7829 13262
rect 7885 13245 7911 13262
rect 7803 13240 7810 13245
rect 7967 13240 7993 13296
rect 8049 13249 8075 13266
rect 8131 13240 8157 13296
rect 8221 13266 8222 13318
rect 8213 13249 8222 13266
rect 5646 13216 5660 13240
rect 5712 13216 6148 13240
rect 6200 13216 6214 13240
rect 6266 13216 6702 13240
rect 6754 13216 6768 13240
rect 6820 13216 7256 13240
rect 7308 13216 7322 13240
rect 7374 13216 7810 13240
rect 7862 13216 7876 13240
rect 7928 13216 8047 13240
rect 8099 13216 8169 13240
rect 2270 13180 5613 13193
rect 2322 13128 2392 13180
rect 2444 13176 5613 13180
rect 5669 13176 5696 13193
rect 2444 13128 2824 13176
rect 2270 13124 2824 13128
rect 2876 13124 2890 13176
rect 2942 13124 3378 13176
rect 3430 13124 3444 13176
rect 3496 13124 3932 13176
rect 3984 13124 3998 13176
rect 4050 13124 4486 13176
rect 4538 13124 4552 13176
rect 4604 13124 5040 13176
rect 5092 13124 5106 13176
rect 5158 13124 5594 13176
rect 5752 13160 5779 13216
rect 5835 13160 5861 13216
rect 5917 13160 5943 13216
rect 5999 13160 6025 13216
rect 6081 13160 6107 13216
rect 6266 13193 6271 13216
rect 6163 13176 6189 13193
rect 6245 13176 6271 13193
rect 6266 13160 6271 13176
rect 6327 13160 6353 13216
rect 6409 13160 6435 13216
rect 6491 13160 6517 13216
rect 6573 13160 6599 13216
rect 6655 13160 6681 13216
rect 6754 13193 6763 13216
rect 6820 13193 6845 13216
rect 6737 13176 6763 13193
rect 6819 13176 6845 13193
rect 6754 13160 6763 13176
rect 6820 13160 6845 13176
rect 6901 13160 6927 13216
rect 6983 13160 7009 13216
rect 7065 13160 7091 13216
rect 7147 13160 7173 13216
rect 7229 13160 7255 13216
rect 7311 13193 7322 13216
rect 7311 13176 7337 13193
rect 7311 13160 7322 13176
rect 7393 13160 7419 13216
rect 7475 13160 7501 13216
rect 7557 13160 7583 13216
rect 7639 13160 7665 13216
rect 7721 13160 7747 13216
rect 7803 13193 7810 13216
rect 7803 13176 7829 13193
rect 7885 13176 7911 13193
rect 7803 13160 7810 13176
rect 7967 13160 7993 13216
rect 8049 13180 8075 13197
rect 8131 13160 8157 13216
rect 8221 13197 8222 13249
rect 8213 13180 8222 13197
rect 5646 13136 5660 13160
rect 5712 13136 6148 13160
rect 6200 13136 6214 13160
rect 6266 13136 6702 13160
rect 6754 13136 6768 13160
rect 6820 13136 7256 13160
rect 7308 13136 7322 13160
rect 7374 13136 7810 13160
rect 7862 13136 7876 13160
rect 7928 13136 8047 13160
rect 8099 13136 8169 13160
rect 2270 13110 5613 13124
rect 2322 13058 2392 13110
rect 2444 13107 5613 13110
rect 5669 13107 5696 13124
rect 2444 13058 2824 13107
rect 2270 13055 2824 13058
rect 2876 13055 2890 13107
rect 2942 13055 3378 13107
rect 3430 13055 3444 13107
rect 3496 13055 3932 13107
rect 3984 13055 3998 13107
rect 4050 13055 4486 13107
rect 4538 13055 4552 13107
rect 4604 13055 5040 13107
rect 5092 13055 5106 13107
rect 5158 13055 5594 13107
rect 5752 13080 5779 13136
rect 5835 13080 5861 13136
rect 5917 13080 5943 13136
rect 5999 13080 6025 13136
rect 6081 13080 6107 13136
rect 6266 13124 6271 13136
rect 6163 13107 6189 13124
rect 6245 13107 6271 13124
rect 6266 13080 6271 13107
rect 6327 13080 6353 13136
rect 6409 13080 6435 13136
rect 6491 13080 6517 13136
rect 6573 13080 6599 13136
rect 6655 13080 6681 13136
rect 6754 13124 6763 13136
rect 6820 13124 6845 13136
rect 6737 13107 6763 13124
rect 6819 13107 6845 13124
rect 6754 13080 6763 13107
rect 6820 13080 6845 13107
rect 6901 13080 6927 13136
rect 6983 13080 7009 13136
rect 7065 13080 7091 13136
rect 7147 13080 7173 13136
rect 7229 13080 7255 13136
rect 7311 13124 7322 13136
rect 7311 13107 7337 13124
rect 7311 13080 7322 13107
rect 7393 13080 7419 13136
rect 7475 13080 7501 13136
rect 7557 13080 7583 13136
rect 7639 13080 7665 13136
rect 7721 13080 7747 13136
rect 7803 13124 7810 13136
rect 7803 13107 7829 13124
rect 7885 13107 7911 13124
rect 7803 13080 7810 13107
rect 7967 13080 7993 13136
rect 8049 13110 8075 13128
rect 8131 13080 8157 13136
rect 8221 13128 8222 13180
rect 8213 13110 8222 13128
rect 5646 13056 5660 13080
rect 5712 13056 6148 13080
rect 6200 13056 6214 13080
rect 6266 13056 6702 13080
rect 6754 13056 6768 13080
rect 6820 13056 7256 13080
rect 7308 13056 7322 13080
rect 7374 13056 7810 13080
rect 7862 13056 7876 13080
rect 7928 13058 8047 13080
rect 8099 13058 8169 13080
rect 8221 13058 8222 13110
rect 7928 13056 8222 13058
rect 2270 13040 5613 13055
rect 2322 12988 2392 13040
rect 2444 13038 5613 13040
rect 5669 13038 5696 13055
rect 2444 12988 2824 13038
rect 2270 12986 2824 12988
rect 2876 12986 2890 13038
rect 2942 12986 3378 13038
rect 3430 12986 3444 13038
rect 3496 12986 3932 13038
rect 3984 12986 3998 13038
rect 4050 12986 4486 13038
rect 4538 12986 4552 13038
rect 4604 12986 5040 13038
rect 5092 12986 5106 13038
rect 5158 12986 5594 13038
rect 5752 13000 5779 13056
rect 5835 13000 5861 13056
rect 5917 13000 5943 13056
rect 5999 13000 6025 13056
rect 6081 13000 6107 13056
rect 6266 13055 6271 13056
rect 6163 13038 6189 13055
rect 6245 13038 6271 13055
rect 6266 13000 6271 13038
rect 6327 13000 6353 13056
rect 6409 13000 6435 13056
rect 6491 13000 6517 13056
rect 6573 13000 6599 13056
rect 6655 13000 6681 13056
rect 6754 13055 6763 13056
rect 6820 13055 6845 13056
rect 6737 13038 6763 13055
rect 6819 13038 6845 13055
rect 6754 13000 6763 13038
rect 6820 13000 6845 13038
rect 6901 13000 6927 13056
rect 6983 13000 7009 13056
rect 7065 13000 7091 13056
rect 7147 13000 7173 13056
rect 7229 13000 7255 13056
rect 7311 13055 7322 13056
rect 7311 13038 7337 13055
rect 7311 13000 7322 13038
rect 7393 13000 7419 13056
rect 7475 13000 7501 13056
rect 7557 13000 7583 13056
rect 7639 13000 7665 13056
rect 7721 13000 7747 13056
rect 7803 13055 7810 13056
rect 7803 13038 7829 13055
rect 7885 13038 7911 13055
rect 7803 13000 7810 13038
rect 7967 13000 7993 13056
rect 8049 13040 8075 13056
rect 8131 13000 8157 13056
rect 8213 13040 8222 13056
rect 5646 12986 5660 13000
rect 5712 12986 6148 13000
rect 6200 12986 6214 13000
rect 6266 12986 6702 13000
rect 6754 12986 6768 13000
rect 6820 12986 7256 13000
rect 7308 12986 7322 13000
rect 7374 12986 7810 13000
rect 7862 12986 7876 13000
rect 7928 12988 8047 13000
rect 8099 12988 8169 13000
rect 8221 12988 8222 13040
rect 7928 12986 8222 12988
rect 2270 12976 8222 12986
rect 2270 12970 5613 12976
rect 2322 12918 2392 12970
rect 2444 12968 5613 12970
rect 5669 12968 5696 12976
rect 2444 12918 2824 12968
rect 2270 12916 2824 12918
rect 2876 12916 2890 12968
rect 2942 12916 3378 12968
rect 3430 12916 3444 12968
rect 3496 12916 3932 12968
rect 3984 12916 3998 12968
rect 4050 12916 4486 12968
rect 4538 12916 4552 12968
rect 4604 12916 5040 12968
rect 5092 12916 5106 12968
rect 5158 12916 5594 12968
rect 5752 12920 5779 12976
rect 5835 12920 5861 12976
rect 5917 12920 5943 12976
rect 5999 12920 6025 12976
rect 6081 12920 6107 12976
rect 6163 12968 6189 12976
rect 6245 12968 6271 12976
rect 6266 12920 6271 12968
rect 6327 12920 6353 12976
rect 6409 12920 6435 12976
rect 6491 12920 6517 12976
rect 6573 12920 6599 12976
rect 6655 12920 6681 12976
rect 6737 12968 6763 12976
rect 6819 12968 6845 12976
rect 6754 12920 6763 12968
rect 6820 12920 6845 12968
rect 6901 12920 6927 12976
rect 6983 12920 7009 12976
rect 7065 12920 7091 12976
rect 7147 12920 7173 12976
rect 7229 12920 7255 12976
rect 7311 12968 7337 12976
rect 7311 12920 7322 12968
rect 7393 12920 7419 12976
rect 7475 12920 7501 12976
rect 7557 12920 7583 12976
rect 7639 12920 7665 12976
rect 7721 12920 7747 12976
rect 7803 12968 7829 12976
rect 7885 12968 7911 12976
rect 7803 12920 7810 12968
rect 7967 12920 7993 12976
rect 8049 12970 8075 12976
rect 8131 12920 8157 12976
rect 8213 12970 8222 12976
rect 5646 12916 5660 12920
rect 5712 12916 6148 12920
rect 6200 12916 6214 12920
rect 6266 12916 6702 12920
rect 6754 12916 6768 12920
rect 6820 12916 7256 12920
rect 7308 12916 7322 12920
rect 7374 12916 7810 12920
rect 7862 12916 7876 12920
rect 7928 12918 8047 12920
rect 8099 12918 8169 12920
rect 8221 12918 8222 12970
rect 7928 12916 8222 12918
rect 2270 12900 8222 12916
rect 2322 12848 2392 12900
rect 2444 12898 8047 12900
rect 2444 12848 2824 12898
rect 2270 12846 2824 12848
rect 2876 12846 2890 12898
rect 2942 12846 3378 12898
rect 3430 12846 3444 12898
rect 3496 12846 3932 12898
rect 3984 12846 3998 12898
rect 4050 12846 4486 12898
rect 4538 12846 4552 12898
rect 4604 12846 5040 12898
rect 5092 12846 5106 12898
rect 5158 12846 5594 12898
rect 5646 12896 5660 12898
rect 5712 12896 6148 12898
rect 6200 12896 6214 12898
rect 6266 12896 6702 12898
rect 6754 12896 6768 12898
rect 6820 12896 7256 12898
rect 7308 12896 7322 12898
rect 7374 12896 7810 12898
rect 7862 12896 7876 12898
rect 7928 12896 8047 12898
rect 8099 12896 8169 12900
rect 2270 12840 5613 12846
rect 5669 12840 5696 12846
rect 5752 12840 5779 12896
rect 5835 12840 5861 12896
rect 5917 12840 5943 12896
rect 5999 12840 6025 12896
rect 6081 12840 6107 12896
rect 6266 12846 6271 12896
rect 6163 12840 6189 12846
rect 6245 12840 6271 12846
rect 6327 12840 6353 12896
rect 6409 12840 6435 12896
rect 6491 12840 6517 12896
rect 6573 12840 6599 12896
rect 6655 12840 6681 12896
rect 6754 12846 6763 12896
rect 6820 12846 6845 12896
rect 6737 12840 6763 12846
rect 6819 12840 6845 12846
rect 6901 12840 6927 12896
rect 6983 12840 7009 12896
rect 7065 12840 7091 12896
rect 7147 12840 7173 12896
rect 7229 12840 7255 12896
rect 7311 12846 7322 12896
rect 7311 12840 7337 12846
rect 7393 12840 7419 12896
rect 7475 12840 7501 12896
rect 7557 12840 7583 12896
rect 7639 12840 7665 12896
rect 7721 12840 7747 12896
rect 7803 12846 7810 12896
rect 7803 12840 7829 12846
rect 7885 12840 7911 12846
rect 7967 12840 7993 12896
rect 8049 12840 8075 12848
rect 8131 12840 8157 12896
rect 8221 12848 8222 12900
rect 8213 12840 8222 12848
rect 2724 12719 7651 12720
rect 2724 12663 2733 12719
rect 2789 12663 2814 12719
rect 2870 12663 2895 12719
rect 2951 12663 2976 12719
rect 3032 12663 3057 12719
rect 3113 12714 3138 12719
rect 3194 12714 3219 12719
rect 3275 12663 3300 12719
rect 3356 12663 3381 12719
rect 3437 12663 3462 12719
rect 3518 12663 3543 12719
rect 3599 12663 3624 12719
rect 3680 12714 3705 12719
rect 3761 12714 3786 12719
rect 3773 12663 3786 12714
rect 3842 12663 3867 12719
rect 3923 12663 3948 12719
rect 4004 12663 4029 12719
rect 4085 12663 4110 12719
rect 4166 12663 4191 12719
rect 4247 12714 4272 12719
rect 4261 12663 4272 12714
rect 4328 12663 4353 12719
rect 4409 12663 4434 12719
rect 4490 12663 4515 12719
rect 4571 12663 4596 12719
rect 4652 12663 4677 12719
rect 4733 12663 4758 12719
rect 4814 12714 4839 12719
rect 2724 12662 3101 12663
rect 3153 12662 3167 12663
rect 3219 12662 3655 12663
rect 3707 12662 3721 12663
rect 3773 12662 4209 12663
rect 4261 12662 4275 12663
rect 4327 12662 4763 12663
rect 4815 12662 4829 12714
rect 4895 12663 4920 12719
rect 4976 12663 5001 12719
rect 5057 12663 5082 12719
rect 5138 12663 5163 12719
rect 4881 12662 5163 12663
rect 2724 12645 5163 12662
rect 2724 12639 3101 12645
rect 3153 12639 3167 12645
rect 3219 12639 3655 12645
rect 3707 12639 3721 12645
rect 3773 12639 4209 12645
rect 4261 12639 4275 12645
rect 4327 12639 4763 12645
rect 2724 12583 2733 12639
rect 2789 12583 2814 12639
rect 2870 12583 2895 12639
rect 2951 12583 2976 12639
rect 3032 12583 3057 12639
rect 3113 12583 3138 12593
rect 3194 12583 3219 12593
rect 3275 12583 3300 12639
rect 3356 12583 3381 12639
rect 3437 12583 3462 12639
rect 3518 12583 3543 12639
rect 3599 12583 3624 12639
rect 3773 12593 3786 12639
rect 3680 12583 3705 12593
rect 3761 12583 3786 12593
rect 3842 12583 3867 12639
rect 3923 12583 3948 12639
rect 4004 12583 4029 12639
rect 4085 12583 4110 12639
rect 4166 12583 4191 12639
rect 4261 12593 4272 12639
rect 4247 12583 4272 12593
rect 4328 12583 4353 12639
rect 4409 12583 4434 12639
rect 4490 12583 4515 12639
rect 4571 12583 4596 12639
rect 4652 12583 4677 12639
rect 4733 12583 4758 12639
rect 4815 12593 4829 12645
rect 4881 12639 5163 12645
rect 4814 12583 4839 12593
rect 4895 12583 4920 12639
rect 4976 12583 5001 12639
rect 5057 12583 5082 12639
rect 5138 12583 5163 12639
rect 2724 12576 5163 12583
rect 2724 12559 3101 12576
rect 3153 12559 3167 12576
rect 3219 12559 3655 12576
rect 3707 12559 3721 12576
rect 3773 12559 4209 12576
rect 4261 12559 4275 12576
rect 4327 12559 4763 12576
rect 2724 12503 2733 12559
rect 2789 12503 2814 12559
rect 2870 12503 2895 12559
rect 2951 12503 2976 12559
rect 3032 12503 3057 12559
rect 3113 12507 3138 12524
rect 3194 12507 3219 12524
rect 3275 12503 3300 12559
rect 3356 12503 3381 12559
rect 3437 12503 3462 12559
rect 3518 12503 3543 12559
rect 3599 12503 3624 12559
rect 3773 12524 3786 12559
rect 3680 12507 3705 12524
rect 3761 12507 3786 12524
rect 3773 12503 3786 12507
rect 3842 12503 3867 12559
rect 3923 12503 3948 12559
rect 4004 12503 4029 12559
rect 4085 12503 4110 12559
rect 4166 12503 4191 12559
rect 4261 12524 4272 12559
rect 4247 12507 4272 12524
rect 4261 12503 4272 12507
rect 4328 12503 4353 12559
rect 4409 12503 4434 12559
rect 4490 12503 4515 12559
rect 4571 12503 4596 12559
rect 4652 12503 4677 12559
rect 4733 12503 4758 12559
rect 4815 12524 4829 12576
rect 4881 12559 5163 12576
rect 4814 12507 4839 12524
rect 2724 12479 3101 12503
rect 3153 12479 3167 12503
rect 3219 12479 3655 12503
rect 3707 12479 3721 12503
rect 3773 12479 4209 12503
rect 4261 12479 4275 12503
rect 4327 12479 4763 12503
rect 2724 12423 2733 12479
rect 2789 12423 2814 12479
rect 2870 12423 2895 12479
rect 2951 12423 2976 12479
rect 3032 12423 3057 12479
rect 3113 12438 3138 12455
rect 3194 12438 3219 12455
rect 3275 12423 3300 12479
rect 3356 12423 3381 12479
rect 3437 12423 3462 12479
rect 3518 12423 3543 12479
rect 3599 12423 3624 12479
rect 3773 12455 3786 12479
rect 3680 12438 3705 12455
rect 3761 12438 3786 12455
rect 3773 12423 3786 12438
rect 3842 12423 3867 12479
rect 3923 12423 3948 12479
rect 4004 12423 4029 12479
rect 4085 12423 4110 12479
rect 4166 12423 4191 12479
rect 4261 12455 4272 12479
rect 4247 12438 4272 12455
rect 4261 12423 4272 12438
rect 4328 12423 4353 12479
rect 4409 12423 4434 12479
rect 4490 12423 4515 12479
rect 4571 12423 4596 12479
rect 4652 12423 4677 12479
rect 4733 12423 4758 12479
rect 4815 12455 4829 12507
rect 4895 12503 4920 12559
rect 4976 12503 5001 12559
rect 5057 12503 5082 12559
rect 5138 12503 5163 12559
rect 4881 12479 5163 12503
rect 4814 12438 4839 12455
rect 2724 12399 3101 12423
rect 3153 12399 3167 12423
rect 3219 12399 3655 12423
rect 3707 12399 3721 12423
rect 3773 12399 4209 12423
rect 4261 12399 4275 12423
rect 4327 12399 4763 12423
rect 2724 12343 2733 12399
rect 2789 12343 2814 12399
rect 2870 12343 2895 12399
rect 2951 12343 2976 12399
rect 3032 12343 3057 12399
rect 3113 12368 3138 12386
rect 3194 12368 3219 12386
rect 3275 12343 3300 12399
rect 3356 12343 3381 12399
rect 3437 12343 3462 12399
rect 3518 12343 3543 12399
rect 3599 12343 3624 12399
rect 3773 12386 3786 12399
rect 3680 12368 3705 12386
rect 3761 12368 3786 12386
rect 3773 12343 3786 12368
rect 3842 12343 3867 12399
rect 3923 12343 3948 12399
rect 4004 12343 4029 12399
rect 4085 12343 4110 12399
rect 4166 12343 4191 12399
rect 4261 12386 4272 12399
rect 4247 12368 4272 12386
rect 4261 12343 4272 12368
rect 4328 12343 4353 12399
rect 4409 12343 4434 12399
rect 4490 12343 4515 12399
rect 4571 12343 4596 12399
rect 4652 12343 4677 12399
rect 4733 12343 4758 12399
rect 4815 12386 4829 12438
rect 4895 12423 4920 12479
rect 4976 12423 5001 12479
rect 5057 12423 5082 12479
rect 5138 12423 5163 12479
rect 4881 12399 5163 12423
rect 4814 12368 4839 12386
rect 2724 12319 3101 12343
rect 3153 12319 3167 12343
rect 3219 12319 3655 12343
rect 3707 12319 3721 12343
rect 3773 12319 4209 12343
rect 4261 12319 4275 12343
rect 4327 12319 4763 12343
rect 2724 12263 2733 12319
rect 2789 12263 2814 12319
rect 2870 12263 2895 12319
rect 2951 12263 2976 12319
rect 3032 12263 3057 12319
rect 3113 12298 3138 12316
rect 3194 12298 3219 12316
rect 3275 12263 3300 12319
rect 3356 12263 3381 12319
rect 3437 12263 3462 12319
rect 3518 12263 3543 12319
rect 3599 12263 3624 12319
rect 3773 12316 3786 12319
rect 3680 12298 3705 12316
rect 3761 12298 3786 12316
rect 3773 12263 3786 12298
rect 3842 12263 3867 12319
rect 3923 12263 3948 12319
rect 4004 12263 4029 12319
rect 4085 12263 4110 12319
rect 4166 12263 4191 12319
rect 4261 12316 4272 12319
rect 4247 12298 4272 12316
rect 4261 12263 4272 12298
rect 4328 12263 4353 12319
rect 4409 12263 4434 12319
rect 4490 12263 4515 12319
rect 4571 12263 4596 12319
rect 4652 12263 4677 12319
rect 4733 12263 4758 12319
rect 4815 12316 4829 12368
rect 4895 12343 4920 12399
rect 4976 12343 5001 12399
rect 5057 12343 5082 12399
rect 5138 12343 5163 12399
rect 4881 12319 5163 12343
rect 4814 12298 4839 12316
rect 2724 12246 3101 12263
rect 3153 12246 3167 12263
rect 3219 12246 3655 12263
rect 3707 12246 3721 12263
rect 3773 12246 4209 12263
rect 4261 12246 4275 12263
rect 4327 12246 4763 12263
rect 4815 12246 4829 12298
rect 4895 12263 4920 12319
rect 4976 12263 5001 12319
rect 5057 12263 5082 12319
rect 5138 12263 5163 12319
rect 4881 12246 5163 12263
rect 2724 12239 5163 12246
rect 2724 12183 2733 12239
rect 2789 12183 2814 12239
rect 2870 12183 2895 12239
rect 2951 12183 2976 12239
rect 3032 12183 3057 12239
rect 3113 12228 3138 12239
rect 3194 12228 3219 12239
rect 3275 12183 3300 12239
rect 3356 12183 3381 12239
rect 3437 12183 3462 12239
rect 3518 12183 3543 12239
rect 3599 12183 3624 12239
rect 3680 12228 3705 12239
rect 3761 12228 3786 12239
rect 3773 12183 3786 12228
rect 3842 12183 3867 12239
rect 3923 12183 3948 12239
rect 4004 12183 4029 12239
rect 4085 12183 4110 12239
rect 4166 12183 4191 12239
rect 4247 12228 4272 12239
rect 4261 12183 4272 12228
rect 4328 12183 4353 12239
rect 4409 12183 4434 12239
rect 4490 12183 4515 12239
rect 4571 12183 4596 12239
rect 4652 12183 4677 12239
rect 4733 12183 4758 12239
rect 4814 12228 4839 12239
rect 2724 12176 3101 12183
rect 3153 12176 3167 12183
rect 3219 12176 3655 12183
rect 3707 12176 3721 12183
rect 3773 12176 4209 12183
rect 4261 12176 4275 12183
rect 4327 12176 4763 12183
rect 4815 12176 4829 12228
rect 4895 12183 4920 12239
rect 4976 12183 5001 12239
rect 5057 12183 5082 12239
rect 5138 12183 5163 12239
rect 4881 12176 5163 12183
rect 2724 12159 5163 12176
rect 2724 12103 2733 12159
rect 2789 12103 2814 12159
rect 2870 12103 2895 12159
rect 2951 12103 2976 12159
rect 3032 12103 3057 12159
rect 3113 12158 3138 12159
rect 3194 12158 3219 12159
rect 3113 12103 3138 12106
rect 3194 12103 3219 12106
rect 3275 12103 3300 12159
rect 3356 12103 3381 12159
rect 3437 12103 3462 12159
rect 3518 12103 3543 12159
rect 3599 12103 3624 12159
rect 3680 12158 3705 12159
rect 3761 12158 3786 12159
rect 3773 12106 3786 12158
rect 3680 12103 3705 12106
rect 3761 12103 3786 12106
rect 3842 12103 3867 12159
rect 3923 12103 3948 12159
rect 4004 12103 4029 12159
rect 4085 12103 4110 12159
rect 4166 12103 4191 12159
rect 4247 12158 4272 12159
rect 4261 12106 4272 12158
rect 4247 12103 4272 12106
rect 4328 12103 4353 12159
rect 4409 12103 4434 12159
rect 4490 12103 4515 12159
rect 4571 12103 4596 12159
rect 4652 12103 4677 12159
rect 4733 12103 4758 12159
rect 4814 12158 4839 12159
rect 4815 12106 4829 12158
rect 4814 12103 4839 12106
rect 4895 12103 4920 12159
rect 4976 12103 5001 12159
rect 5057 12103 5082 12159
rect 5138 12103 5163 12159
rect 5299 12714 7651 12719
rect 5299 12662 5317 12714
rect 5369 12662 5383 12714
rect 5435 12662 5871 12714
rect 5923 12662 5937 12714
rect 5989 12662 6425 12714
rect 6477 12662 6491 12714
rect 6543 12662 6979 12714
rect 7031 12662 7045 12714
rect 7097 12662 7533 12714
rect 7585 12662 7599 12714
rect 5299 12645 7651 12662
rect 5299 12593 5317 12645
rect 5369 12593 5383 12645
rect 5435 12593 5871 12645
rect 5923 12593 5937 12645
rect 5989 12593 6425 12645
rect 6477 12593 6491 12645
rect 6543 12593 6979 12645
rect 7031 12593 7045 12645
rect 7097 12593 7533 12645
rect 7585 12593 7599 12645
rect 5299 12576 7651 12593
rect 5299 12524 5317 12576
rect 5369 12524 5383 12576
rect 5435 12524 5871 12576
rect 5923 12524 5937 12576
rect 5989 12524 6425 12576
rect 6477 12524 6491 12576
rect 6543 12524 6979 12576
rect 7031 12524 7045 12576
rect 7097 12524 7533 12576
rect 7585 12524 7599 12576
rect 5299 12507 7651 12524
rect 5299 12455 5317 12507
rect 5369 12455 5383 12507
rect 5435 12455 5871 12507
rect 5923 12455 5937 12507
rect 5989 12455 6425 12507
rect 6477 12455 6491 12507
rect 6543 12455 6979 12507
rect 7031 12455 7045 12507
rect 7097 12455 7533 12507
rect 7585 12455 7599 12507
rect 5299 12438 7651 12455
rect 5299 12386 5317 12438
rect 5369 12386 5383 12438
rect 5435 12386 5871 12438
rect 5923 12386 5937 12438
rect 5989 12386 6425 12438
rect 6477 12386 6491 12438
rect 6543 12386 6979 12438
rect 7031 12386 7045 12438
rect 7097 12386 7533 12438
rect 7585 12386 7599 12438
rect 5299 12368 7651 12386
rect 5299 12316 5317 12368
rect 5369 12316 5383 12368
rect 5435 12316 5871 12368
rect 5923 12316 5937 12368
rect 5989 12316 6425 12368
rect 6477 12316 6491 12368
rect 6543 12316 6979 12368
rect 7031 12316 7045 12368
rect 7097 12316 7533 12368
rect 7585 12316 7599 12368
rect 5299 12298 7651 12316
rect 5299 12246 5317 12298
rect 5369 12246 5383 12298
rect 5435 12246 5871 12298
rect 5923 12246 5937 12298
rect 5989 12246 6425 12298
rect 6477 12246 6491 12298
rect 6543 12246 6979 12298
rect 7031 12246 7045 12298
rect 7097 12246 7533 12298
rect 7585 12246 7599 12298
rect 5299 12228 7651 12246
rect 5299 12176 5317 12228
rect 5369 12176 5383 12228
rect 5435 12176 5871 12228
rect 5923 12176 5937 12228
rect 5989 12176 6425 12228
rect 6477 12176 6491 12228
rect 6543 12176 6979 12228
rect 7031 12176 7045 12228
rect 7097 12176 7533 12228
rect 7585 12176 7599 12228
rect 5299 12158 7651 12176
rect 5299 12106 5317 12158
rect 5369 12106 5383 12158
rect 5435 12106 5871 12158
rect 5923 12106 5937 12158
rect 5989 12106 6425 12158
rect 6477 12106 6491 12158
rect 6543 12106 6979 12158
rect 7031 12106 7045 12158
rect 7097 12106 7533 12158
rect 7585 12106 7599 12158
rect 5299 12103 7651 12106
rect 2724 12100 7651 12103
rect 2270 11456 8222 11462
rect 2322 11404 2392 11456
rect 2444 11452 5613 11456
rect 5669 11452 5696 11456
rect 2444 11404 2824 11452
rect 2270 11400 2824 11404
rect 2876 11400 2890 11452
rect 2942 11400 3378 11452
rect 3430 11400 3444 11452
rect 3496 11400 3932 11452
rect 3984 11400 3998 11452
rect 4050 11400 4486 11452
rect 4538 11400 4552 11452
rect 4604 11400 5040 11452
rect 5092 11400 5106 11452
rect 5158 11400 5594 11452
rect 5752 11400 5779 11456
rect 5835 11400 5861 11456
rect 5917 11400 5943 11456
rect 5999 11400 6025 11456
rect 6081 11400 6107 11456
rect 6163 11452 6189 11456
rect 6245 11452 6271 11456
rect 6266 11400 6271 11452
rect 6327 11400 6353 11456
rect 6409 11400 6435 11456
rect 6491 11400 6517 11456
rect 6573 11400 6599 11456
rect 6655 11400 6681 11456
rect 6737 11452 6763 11456
rect 6819 11452 6845 11456
rect 6754 11400 6763 11452
rect 6820 11400 6845 11452
rect 6901 11400 6927 11456
rect 6983 11400 7009 11456
rect 7065 11400 7091 11456
rect 7147 11400 7173 11456
rect 7229 11400 7255 11456
rect 7311 11452 7337 11456
rect 7311 11400 7322 11452
rect 7393 11400 7419 11456
rect 7475 11400 7501 11456
rect 7557 11400 7583 11456
rect 7639 11400 7665 11456
rect 7721 11400 7747 11456
rect 7803 11452 7829 11456
rect 7885 11452 7911 11456
rect 7803 11400 7810 11452
rect 7967 11400 7993 11456
rect 8049 11400 8075 11404
rect 8131 11400 8157 11456
rect 8221 11404 8222 11456
rect 8213 11400 8222 11404
rect 2270 11387 8222 11400
rect 2322 11335 2392 11387
rect 2444 11383 8047 11387
rect 2444 11335 2824 11383
rect 2270 11331 2824 11335
rect 2876 11331 2890 11383
rect 2942 11331 3378 11383
rect 3430 11331 3444 11383
rect 3496 11331 3932 11383
rect 3984 11331 3998 11383
rect 4050 11331 4486 11383
rect 4538 11331 4552 11383
rect 4604 11331 5040 11383
rect 5092 11331 5106 11383
rect 5158 11331 5594 11383
rect 5646 11376 5660 11383
rect 5712 11376 6148 11383
rect 6200 11376 6214 11383
rect 6266 11376 6702 11383
rect 6754 11376 6768 11383
rect 6820 11376 7256 11383
rect 7308 11376 7322 11383
rect 7374 11376 7810 11383
rect 7862 11376 7876 11383
rect 7928 11376 8047 11383
rect 8099 11376 8169 11387
rect 2270 11320 5613 11331
rect 5669 11320 5696 11331
rect 5752 11320 5779 11376
rect 5835 11320 5861 11376
rect 5917 11320 5943 11376
rect 5999 11320 6025 11376
rect 6081 11320 6107 11376
rect 6266 11331 6271 11376
rect 6163 11320 6189 11331
rect 6245 11320 6271 11331
rect 6327 11320 6353 11376
rect 6409 11320 6435 11376
rect 6491 11320 6517 11376
rect 6573 11320 6599 11376
rect 6655 11320 6681 11376
rect 6754 11331 6763 11376
rect 6820 11331 6845 11376
rect 6737 11320 6763 11331
rect 6819 11320 6845 11331
rect 6901 11320 6927 11376
rect 6983 11320 7009 11376
rect 7065 11320 7091 11376
rect 7147 11320 7173 11376
rect 7229 11320 7255 11376
rect 7311 11331 7322 11376
rect 7311 11320 7337 11331
rect 7393 11320 7419 11376
rect 7475 11320 7501 11376
rect 7557 11320 7583 11376
rect 7639 11320 7665 11376
rect 7721 11320 7747 11376
rect 7803 11331 7810 11376
rect 7803 11320 7829 11331
rect 7885 11320 7911 11331
rect 7967 11320 7993 11376
rect 8049 11320 8075 11335
rect 8131 11320 8157 11376
rect 8221 11335 8222 11387
rect 8213 11320 8222 11335
rect 2270 11318 8222 11320
rect 2322 11266 2392 11318
rect 2444 11314 8047 11318
rect 2444 11266 2824 11314
rect 2270 11262 2824 11266
rect 2876 11262 2890 11314
rect 2942 11262 3378 11314
rect 3430 11262 3444 11314
rect 3496 11262 3932 11314
rect 3984 11262 3998 11314
rect 4050 11262 4486 11314
rect 4538 11262 4552 11314
rect 4604 11262 5040 11314
rect 5092 11262 5106 11314
rect 5158 11262 5594 11314
rect 5646 11296 5660 11314
rect 5712 11296 6148 11314
rect 6200 11296 6214 11314
rect 6266 11296 6702 11314
rect 6754 11296 6768 11314
rect 6820 11296 7256 11314
rect 7308 11296 7322 11314
rect 7374 11296 7810 11314
rect 7862 11296 7876 11314
rect 7928 11296 8047 11314
rect 8099 11296 8169 11318
rect 2270 11249 5613 11262
rect 2322 11197 2392 11249
rect 2444 11245 5613 11249
rect 5669 11245 5696 11262
rect 2444 11197 2824 11245
rect 2270 11193 2824 11197
rect 2876 11193 2890 11245
rect 2942 11193 3378 11245
rect 3430 11193 3444 11245
rect 3496 11193 3932 11245
rect 3984 11193 3998 11245
rect 4050 11193 4486 11245
rect 4538 11193 4552 11245
rect 4604 11193 5040 11245
rect 5092 11193 5106 11245
rect 5158 11193 5594 11245
rect 5752 11240 5779 11296
rect 5835 11240 5861 11296
rect 5917 11240 5943 11296
rect 5999 11240 6025 11296
rect 6081 11240 6107 11296
rect 6266 11262 6271 11296
rect 6163 11245 6189 11262
rect 6245 11245 6271 11262
rect 6266 11240 6271 11245
rect 6327 11240 6353 11296
rect 6409 11240 6435 11296
rect 6491 11240 6517 11296
rect 6573 11240 6599 11296
rect 6655 11240 6681 11296
rect 6754 11262 6763 11296
rect 6820 11262 6845 11296
rect 6737 11245 6763 11262
rect 6819 11245 6845 11262
rect 6754 11240 6763 11245
rect 6820 11240 6845 11245
rect 6901 11240 6927 11296
rect 6983 11240 7009 11296
rect 7065 11240 7091 11296
rect 7147 11240 7173 11296
rect 7229 11240 7255 11296
rect 7311 11262 7322 11296
rect 7311 11245 7337 11262
rect 7311 11240 7322 11245
rect 7393 11240 7419 11296
rect 7475 11240 7501 11296
rect 7557 11240 7583 11296
rect 7639 11240 7665 11296
rect 7721 11240 7747 11296
rect 7803 11262 7810 11296
rect 7803 11245 7829 11262
rect 7885 11245 7911 11262
rect 7803 11240 7810 11245
rect 7967 11240 7993 11296
rect 8049 11249 8075 11266
rect 8131 11240 8157 11296
rect 8221 11266 8222 11318
rect 8213 11249 8222 11266
rect 5646 11216 5660 11240
rect 5712 11216 6148 11240
rect 6200 11216 6214 11240
rect 6266 11216 6702 11240
rect 6754 11216 6768 11240
rect 6820 11216 7256 11240
rect 7308 11216 7322 11240
rect 7374 11216 7810 11240
rect 7862 11216 7876 11240
rect 7928 11216 8047 11240
rect 8099 11216 8169 11240
rect 2270 11180 5613 11193
rect 2322 11128 2392 11180
rect 2444 11176 5613 11180
rect 5669 11176 5696 11193
rect 2444 11128 2824 11176
rect 2270 11124 2824 11128
rect 2876 11124 2890 11176
rect 2942 11124 3378 11176
rect 3430 11124 3444 11176
rect 3496 11124 3932 11176
rect 3984 11124 3998 11176
rect 4050 11124 4486 11176
rect 4538 11124 4552 11176
rect 4604 11124 5040 11176
rect 5092 11124 5106 11176
rect 5158 11124 5594 11176
rect 5752 11160 5779 11216
rect 5835 11160 5861 11216
rect 5917 11160 5943 11216
rect 5999 11160 6025 11216
rect 6081 11160 6107 11216
rect 6266 11193 6271 11216
rect 6163 11176 6189 11193
rect 6245 11176 6271 11193
rect 6266 11160 6271 11176
rect 6327 11160 6353 11216
rect 6409 11160 6435 11216
rect 6491 11160 6517 11216
rect 6573 11160 6599 11216
rect 6655 11160 6681 11216
rect 6754 11193 6763 11216
rect 6820 11193 6845 11216
rect 6737 11176 6763 11193
rect 6819 11176 6845 11193
rect 6754 11160 6763 11176
rect 6820 11160 6845 11176
rect 6901 11160 6927 11216
rect 6983 11160 7009 11216
rect 7065 11160 7091 11216
rect 7147 11160 7173 11216
rect 7229 11160 7255 11216
rect 7311 11193 7322 11216
rect 7311 11176 7337 11193
rect 7311 11160 7322 11176
rect 7393 11160 7419 11216
rect 7475 11160 7501 11216
rect 7557 11160 7583 11216
rect 7639 11160 7665 11216
rect 7721 11160 7747 11216
rect 7803 11193 7810 11216
rect 7803 11176 7829 11193
rect 7885 11176 7911 11193
rect 7803 11160 7810 11176
rect 7967 11160 7993 11216
rect 8049 11180 8075 11197
rect 8131 11160 8157 11216
rect 8221 11197 8222 11249
rect 8213 11180 8222 11197
rect 5646 11136 5660 11160
rect 5712 11136 6148 11160
rect 6200 11136 6214 11160
rect 6266 11136 6702 11160
rect 6754 11136 6768 11160
rect 6820 11136 7256 11160
rect 7308 11136 7322 11160
rect 7374 11136 7810 11160
rect 7862 11136 7876 11160
rect 7928 11136 8047 11160
rect 8099 11136 8169 11160
rect 2270 11110 5613 11124
rect 2322 11058 2392 11110
rect 2444 11107 5613 11110
rect 5669 11107 5696 11124
rect 2444 11058 2824 11107
rect 2270 11055 2824 11058
rect 2876 11055 2890 11107
rect 2942 11055 3378 11107
rect 3430 11055 3444 11107
rect 3496 11055 3932 11107
rect 3984 11055 3998 11107
rect 4050 11055 4486 11107
rect 4538 11055 4552 11107
rect 4604 11055 5040 11107
rect 5092 11055 5106 11107
rect 5158 11055 5594 11107
rect 5752 11080 5779 11136
rect 5835 11080 5861 11136
rect 5917 11080 5943 11136
rect 5999 11080 6025 11136
rect 6081 11080 6107 11136
rect 6266 11124 6271 11136
rect 6163 11107 6189 11124
rect 6245 11107 6271 11124
rect 6266 11080 6271 11107
rect 6327 11080 6353 11136
rect 6409 11080 6435 11136
rect 6491 11080 6517 11136
rect 6573 11080 6599 11136
rect 6655 11080 6681 11136
rect 6754 11124 6763 11136
rect 6820 11124 6845 11136
rect 6737 11107 6763 11124
rect 6819 11107 6845 11124
rect 6754 11080 6763 11107
rect 6820 11080 6845 11107
rect 6901 11080 6927 11136
rect 6983 11080 7009 11136
rect 7065 11080 7091 11136
rect 7147 11080 7173 11136
rect 7229 11080 7255 11136
rect 7311 11124 7322 11136
rect 7311 11107 7337 11124
rect 7311 11080 7322 11107
rect 7393 11080 7419 11136
rect 7475 11080 7501 11136
rect 7557 11080 7583 11136
rect 7639 11080 7665 11136
rect 7721 11080 7747 11136
rect 7803 11124 7810 11136
rect 7803 11107 7829 11124
rect 7885 11107 7911 11124
rect 7803 11080 7810 11107
rect 7967 11080 7993 11136
rect 8049 11110 8075 11128
rect 8131 11080 8157 11136
rect 8221 11128 8222 11180
rect 8213 11110 8222 11128
rect 5646 11056 5660 11080
rect 5712 11056 6148 11080
rect 6200 11056 6214 11080
rect 6266 11056 6702 11080
rect 6754 11056 6768 11080
rect 6820 11056 7256 11080
rect 7308 11056 7322 11080
rect 7374 11056 7810 11080
rect 7862 11056 7876 11080
rect 7928 11058 8047 11080
rect 8099 11058 8169 11080
rect 8221 11058 8222 11110
rect 7928 11056 8222 11058
rect 2270 11040 5613 11055
rect 2322 10988 2392 11040
rect 2444 11038 5613 11040
rect 5669 11038 5696 11055
rect 2444 10988 2824 11038
rect 2270 10986 2824 10988
rect 2876 10986 2890 11038
rect 2942 10986 3378 11038
rect 3430 10986 3444 11038
rect 3496 10986 3932 11038
rect 3984 10986 3998 11038
rect 4050 10986 4486 11038
rect 4538 10986 4552 11038
rect 4604 10986 5040 11038
rect 5092 10986 5106 11038
rect 5158 10986 5594 11038
rect 5752 11000 5779 11056
rect 5835 11000 5861 11056
rect 5917 11000 5943 11056
rect 5999 11000 6025 11056
rect 6081 11000 6107 11056
rect 6266 11055 6271 11056
rect 6163 11038 6189 11055
rect 6245 11038 6271 11055
rect 6266 11000 6271 11038
rect 6327 11000 6353 11056
rect 6409 11000 6435 11056
rect 6491 11000 6517 11056
rect 6573 11000 6599 11056
rect 6655 11000 6681 11056
rect 6754 11055 6763 11056
rect 6820 11055 6845 11056
rect 6737 11038 6763 11055
rect 6819 11038 6845 11055
rect 6754 11000 6763 11038
rect 6820 11000 6845 11038
rect 6901 11000 6927 11056
rect 6983 11000 7009 11056
rect 7065 11000 7091 11056
rect 7147 11000 7173 11056
rect 7229 11000 7255 11056
rect 7311 11055 7322 11056
rect 7311 11038 7337 11055
rect 7311 11000 7322 11038
rect 7393 11000 7419 11056
rect 7475 11000 7501 11056
rect 7557 11000 7583 11056
rect 7639 11000 7665 11056
rect 7721 11000 7747 11056
rect 7803 11055 7810 11056
rect 7803 11038 7829 11055
rect 7885 11038 7911 11055
rect 7803 11000 7810 11038
rect 7967 11000 7993 11056
rect 8049 11040 8075 11056
rect 8131 11000 8157 11056
rect 8213 11040 8222 11056
rect 5646 10986 5660 11000
rect 5712 10986 6148 11000
rect 6200 10986 6214 11000
rect 6266 10986 6702 11000
rect 6754 10986 6768 11000
rect 6820 10986 7256 11000
rect 7308 10986 7322 11000
rect 7374 10986 7810 11000
rect 7862 10986 7876 11000
rect 7928 10988 8047 11000
rect 8099 10988 8169 11000
rect 8221 10988 8222 11040
rect 7928 10986 8222 10988
rect 2270 10976 8222 10986
rect 2270 10970 5613 10976
rect 2322 10918 2392 10970
rect 2444 10968 5613 10970
rect 5669 10968 5696 10976
rect 2444 10918 2824 10968
rect 2270 10916 2824 10918
rect 2876 10916 2890 10968
rect 2942 10916 3378 10968
rect 3430 10916 3444 10968
rect 3496 10916 3932 10968
rect 3984 10916 3998 10968
rect 4050 10916 4486 10968
rect 4538 10916 4552 10968
rect 4604 10916 5040 10968
rect 5092 10916 5106 10968
rect 5158 10916 5594 10968
rect 5752 10920 5779 10976
rect 5835 10920 5861 10976
rect 5917 10920 5943 10976
rect 5999 10920 6025 10976
rect 6081 10920 6107 10976
rect 6163 10968 6189 10976
rect 6245 10968 6271 10976
rect 6266 10920 6271 10968
rect 6327 10920 6353 10976
rect 6409 10920 6435 10976
rect 6491 10920 6517 10976
rect 6573 10920 6599 10976
rect 6655 10920 6681 10976
rect 6737 10968 6763 10976
rect 6819 10968 6845 10976
rect 6754 10920 6763 10968
rect 6820 10920 6845 10968
rect 6901 10920 6927 10976
rect 6983 10920 7009 10976
rect 7065 10920 7091 10976
rect 7147 10920 7173 10976
rect 7229 10920 7255 10976
rect 7311 10968 7337 10976
rect 7311 10920 7322 10968
rect 7393 10920 7419 10976
rect 7475 10920 7501 10976
rect 7557 10920 7583 10976
rect 7639 10920 7665 10976
rect 7721 10920 7747 10976
rect 7803 10968 7829 10976
rect 7885 10968 7911 10976
rect 7803 10920 7810 10968
rect 7967 10920 7993 10976
rect 8049 10970 8075 10976
rect 8131 10920 8157 10976
rect 8213 10970 8222 10976
rect 5646 10916 5660 10920
rect 5712 10916 6148 10920
rect 6200 10916 6214 10920
rect 6266 10916 6702 10920
rect 6754 10916 6768 10920
rect 6820 10916 7256 10920
rect 7308 10916 7322 10920
rect 7374 10916 7810 10920
rect 7862 10916 7876 10920
rect 7928 10918 8047 10920
rect 8099 10918 8169 10920
rect 8221 10918 8222 10970
rect 7928 10916 8222 10918
rect 2270 10900 8222 10916
rect 2322 10848 2392 10900
rect 2444 10898 8047 10900
rect 2444 10848 2824 10898
rect 2270 10846 2824 10848
rect 2876 10846 2890 10898
rect 2942 10846 3378 10898
rect 3430 10846 3444 10898
rect 3496 10846 3932 10898
rect 3984 10846 3998 10898
rect 4050 10846 4486 10898
rect 4538 10846 4552 10898
rect 4604 10846 5040 10898
rect 5092 10846 5106 10898
rect 5158 10846 5594 10898
rect 5646 10896 5660 10898
rect 5712 10896 6148 10898
rect 6200 10896 6214 10898
rect 6266 10896 6702 10898
rect 6754 10896 6768 10898
rect 6820 10896 7256 10898
rect 7308 10896 7322 10898
rect 7374 10896 7810 10898
rect 7862 10896 7876 10898
rect 7928 10896 8047 10898
rect 8099 10896 8169 10900
rect 2270 10840 5613 10846
rect 5669 10840 5696 10846
rect 5752 10840 5779 10896
rect 5835 10840 5861 10896
rect 5917 10840 5943 10896
rect 5999 10840 6025 10896
rect 6081 10840 6107 10896
rect 6266 10846 6271 10896
rect 6163 10840 6189 10846
rect 6245 10840 6271 10846
rect 6327 10840 6353 10896
rect 6409 10840 6435 10896
rect 6491 10840 6517 10896
rect 6573 10840 6599 10896
rect 6655 10840 6681 10896
rect 6754 10846 6763 10896
rect 6820 10846 6845 10896
rect 6737 10840 6763 10846
rect 6819 10840 6845 10846
rect 6901 10840 6927 10896
rect 6983 10840 7009 10896
rect 7065 10840 7091 10896
rect 7147 10840 7173 10896
rect 7229 10840 7255 10896
rect 7311 10846 7322 10896
rect 7311 10840 7337 10846
rect 7393 10840 7419 10896
rect 7475 10840 7501 10896
rect 7557 10840 7583 10896
rect 7639 10840 7665 10896
rect 7721 10840 7747 10896
rect 7803 10846 7810 10896
rect 7803 10840 7829 10846
rect 7885 10840 7911 10846
rect 7967 10840 7993 10896
rect 8049 10840 8075 10848
rect 8131 10840 8157 10896
rect 8221 10848 8222 10900
rect 8213 10840 8222 10848
rect 2850 10664 2859 10720
rect 2915 10664 2942 10720
rect 2998 10664 3025 10720
rect 3081 10714 3108 10720
rect 3164 10714 3191 10720
rect 3081 10664 3101 10714
rect 3164 10664 3167 10714
rect 3247 10664 3274 10720
rect 3330 10664 3357 10720
rect 3413 10664 3439 10720
rect 3495 10664 3521 10720
rect 3577 10664 3603 10720
rect 3659 10714 3685 10720
rect 3741 10714 3767 10720
rect 3823 10664 3849 10720
rect 3905 10664 3931 10720
rect 3987 10664 4013 10720
rect 4069 10664 4095 10720
rect 4151 10664 4177 10720
rect 4233 10714 4259 10720
rect 4315 10714 4341 10720
rect 4327 10664 4341 10714
rect 4397 10664 4423 10720
rect 4479 10664 4505 10720
rect 4561 10664 4587 10720
rect 4643 10664 4669 10720
rect 4725 10664 4751 10720
rect 4807 10714 4833 10720
rect 2850 10662 3101 10664
rect 3153 10662 3167 10664
rect 3219 10662 3655 10664
rect 3707 10662 3721 10664
rect 3773 10662 4209 10664
rect 4261 10662 4275 10664
rect 4327 10662 4763 10664
rect 4815 10662 4829 10714
rect 4889 10664 4915 10720
rect 4971 10664 4997 10720
rect 5053 10664 5079 10720
rect 5135 10664 5161 10720
rect 5217 10664 5243 10720
rect 5299 10714 7651 10720
rect 5299 10664 5317 10714
rect 4881 10662 5317 10664
rect 5369 10662 5383 10714
rect 5435 10662 5871 10714
rect 5923 10662 5937 10714
rect 5989 10662 6425 10714
rect 6477 10662 6491 10714
rect 6543 10662 6979 10714
rect 7031 10662 7045 10714
rect 7097 10662 7533 10714
rect 7585 10662 7599 10714
rect 2850 10645 7651 10662
rect 2850 10640 3101 10645
rect 3153 10640 3167 10645
rect 3219 10640 3655 10645
rect 3707 10640 3721 10645
rect 3773 10640 4209 10645
rect 4261 10640 4275 10645
rect 4327 10640 4763 10645
rect 2850 10584 2859 10640
rect 2915 10584 2942 10640
rect 2998 10584 3025 10640
rect 3081 10593 3101 10640
rect 3164 10593 3167 10640
rect 3081 10584 3108 10593
rect 3164 10584 3191 10593
rect 3247 10584 3274 10640
rect 3330 10584 3357 10640
rect 3413 10584 3439 10640
rect 3495 10584 3521 10640
rect 3577 10584 3603 10640
rect 3659 10584 3685 10593
rect 3741 10584 3767 10593
rect 3823 10584 3849 10640
rect 3905 10584 3931 10640
rect 3987 10584 4013 10640
rect 4069 10584 4095 10640
rect 4151 10584 4177 10640
rect 4327 10593 4341 10640
rect 4233 10584 4259 10593
rect 4315 10584 4341 10593
rect 4397 10584 4423 10640
rect 4479 10584 4505 10640
rect 4561 10584 4587 10640
rect 4643 10584 4669 10640
rect 4725 10584 4751 10640
rect 4815 10593 4829 10645
rect 4881 10640 5317 10645
rect 4807 10584 4833 10593
rect 4889 10584 4915 10640
rect 4971 10584 4997 10640
rect 5053 10584 5079 10640
rect 5135 10584 5161 10640
rect 5217 10584 5243 10640
rect 5299 10593 5317 10640
rect 5369 10593 5383 10645
rect 5435 10593 5871 10645
rect 5923 10593 5937 10645
rect 5989 10593 6425 10645
rect 6477 10593 6491 10645
rect 6543 10593 6979 10645
rect 7031 10593 7045 10645
rect 7097 10593 7533 10645
rect 7585 10593 7599 10645
rect 5299 10584 7651 10593
rect 2850 10576 7651 10584
rect 2850 10560 3101 10576
rect 3153 10560 3167 10576
rect 3219 10560 3655 10576
rect 3707 10560 3721 10576
rect 3773 10560 4209 10576
rect 4261 10560 4275 10576
rect 4327 10560 4763 10576
rect 2528 10522 2712 10528
rect 2528 10470 2580 10522
rect 2632 10470 2660 10522
rect 2528 10456 2712 10470
rect 2528 10404 2580 10456
rect 2632 10404 2660 10456
rect 2528 10390 2712 10404
rect 2528 10338 2580 10390
rect 2632 10338 2660 10390
rect 2528 10324 2712 10338
rect 2528 10272 2580 10324
rect 2632 10272 2660 10324
rect 2528 10258 2712 10272
rect 2528 10206 2580 10258
rect 2632 10206 2660 10258
rect 2528 10192 2712 10206
rect 2528 10140 2580 10192
rect 2632 10140 2660 10192
rect 2528 10126 2712 10140
rect 2528 10074 2580 10126
rect 2632 10074 2660 10126
rect 2850 10504 2859 10560
rect 2915 10504 2942 10560
rect 2998 10504 3025 10560
rect 3081 10524 3101 10560
rect 3164 10524 3167 10560
rect 3081 10507 3108 10524
rect 3164 10507 3191 10524
rect 3081 10504 3101 10507
rect 3164 10504 3167 10507
rect 3247 10504 3274 10560
rect 3330 10504 3357 10560
rect 3413 10504 3439 10560
rect 3495 10504 3521 10560
rect 3577 10504 3603 10560
rect 3659 10507 3685 10524
rect 3741 10507 3767 10524
rect 3823 10504 3849 10560
rect 3905 10504 3931 10560
rect 3987 10504 4013 10560
rect 4069 10504 4095 10560
rect 4151 10504 4177 10560
rect 4327 10524 4341 10560
rect 4233 10507 4259 10524
rect 4315 10507 4341 10524
rect 4327 10504 4341 10507
rect 4397 10504 4423 10560
rect 4479 10504 4505 10560
rect 4561 10504 4587 10560
rect 4643 10504 4669 10560
rect 4725 10504 4751 10560
rect 4815 10524 4829 10576
rect 4881 10560 5317 10576
rect 4807 10507 4833 10524
rect 2850 10480 3101 10504
rect 3153 10480 3167 10504
rect 3219 10480 3655 10504
rect 3707 10480 3721 10504
rect 3773 10480 4209 10504
rect 4261 10480 4275 10504
rect 4327 10480 4763 10504
rect 2850 10424 2859 10480
rect 2915 10424 2942 10480
rect 2998 10424 3025 10480
rect 3081 10455 3101 10480
rect 3164 10455 3167 10480
rect 3081 10438 3108 10455
rect 3164 10438 3191 10455
rect 3081 10424 3101 10438
rect 3164 10424 3167 10438
rect 3247 10424 3274 10480
rect 3330 10424 3357 10480
rect 3413 10424 3439 10480
rect 3495 10424 3521 10480
rect 3577 10424 3603 10480
rect 3659 10438 3685 10455
rect 3741 10438 3767 10455
rect 3823 10424 3849 10480
rect 3905 10424 3931 10480
rect 3987 10424 4013 10480
rect 4069 10424 4095 10480
rect 4151 10424 4177 10480
rect 4327 10455 4341 10480
rect 4233 10438 4259 10455
rect 4315 10438 4341 10455
rect 4327 10424 4341 10438
rect 4397 10424 4423 10480
rect 4479 10424 4505 10480
rect 4561 10424 4587 10480
rect 4643 10424 4669 10480
rect 4725 10424 4751 10480
rect 4815 10455 4829 10507
rect 4889 10504 4915 10560
rect 4971 10504 4997 10560
rect 5053 10504 5079 10560
rect 5135 10504 5161 10560
rect 5217 10504 5243 10560
rect 5299 10524 5317 10560
rect 5369 10524 5383 10576
rect 5435 10524 5871 10576
rect 5923 10524 5937 10576
rect 5989 10524 6425 10576
rect 6477 10524 6491 10576
rect 6543 10524 6979 10576
rect 7031 10524 7045 10576
rect 7097 10524 7533 10576
rect 7585 10524 7599 10576
rect 5299 10507 7651 10524
rect 5299 10504 5317 10507
rect 4881 10480 5317 10504
rect 4807 10438 4833 10455
rect 2850 10400 3101 10424
rect 3153 10400 3167 10424
rect 3219 10400 3655 10424
rect 3707 10400 3721 10424
rect 3773 10400 4209 10424
rect 4261 10400 4275 10424
rect 4327 10400 4763 10424
rect 2850 10344 2859 10400
rect 2915 10344 2942 10400
rect 2998 10344 3025 10400
rect 3081 10386 3101 10400
rect 3164 10386 3167 10400
rect 3081 10368 3108 10386
rect 3164 10368 3191 10386
rect 3081 10344 3101 10368
rect 3164 10344 3167 10368
rect 3247 10344 3274 10400
rect 3330 10344 3357 10400
rect 3413 10344 3439 10400
rect 3495 10344 3521 10400
rect 3577 10344 3603 10400
rect 3659 10368 3685 10386
rect 3741 10368 3767 10386
rect 3823 10344 3849 10400
rect 3905 10344 3931 10400
rect 3987 10344 4013 10400
rect 4069 10344 4095 10400
rect 4151 10344 4177 10400
rect 4327 10386 4341 10400
rect 4233 10368 4259 10386
rect 4315 10368 4341 10386
rect 4327 10344 4341 10368
rect 4397 10344 4423 10400
rect 4479 10344 4505 10400
rect 4561 10344 4587 10400
rect 4643 10344 4669 10400
rect 4725 10344 4751 10400
rect 4815 10386 4829 10438
rect 4889 10424 4915 10480
rect 4971 10424 4997 10480
rect 5053 10424 5079 10480
rect 5135 10424 5161 10480
rect 5217 10424 5243 10480
rect 5299 10455 5317 10480
rect 5369 10455 5383 10507
rect 5435 10455 5871 10507
rect 5923 10455 5937 10507
rect 5989 10455 6425 10507
rect 6477 10455 6491 10507
rect 6543 10455 6979 10507
rect 7031 10455 7045 10507
rect 7097 10455 7533 10507
rect 7585 10455 7599 10507
rect 5299 10438 7651 10455
rect 5299 10424 5317 10438
rect 4881 10400 5317 10424
rect 4807 10368 4833 10386
rect 2850 10320 3101 10344
rect 3153 10320 3167 10344
rect 3219 10320 3655 10344
rect 3707 10320 3721 10344
rect 3773 10320 4209 10344
rect 4261 10320 4275 10344
rect 4327 10320 4763 10344
rect 2850 10264 2859 10320
rect 2915 10264 2942 10320
rect 2998 10264 3025 10320
rect 3081 10316 3101 10320
rect 3164 10316 3167 10320
rect 3081 10298 3108 10316
rect 3164 10298 3191 10316
rect 3081 10264 3101 10298
rect 3164 10264 3167 10298
rect 3247 10264 3274 10320
rect 3330 10264 3357 10320
rect 3413 10264 3439 10320
rect 3495 10264 3521 10320
rect 3577 10264 3603 10320
rect 3659 10298 3685 10316
rect 3741 10298 3767 10316
rect 3823 10264 3849 10320
rect 3905 10264 3931 10320
rect 3987 10264 4013 10320
rect 4069 10264 4095 10320
rect 4151 10264 4177 10320
rect 4327 10316 4341 10320
rect 4233 10298 4259 10316
rect 4315 10298 4341 10316
rect 4327 10264 4341 10298
rect 4397 10264 4423 10320
rect 4479 10264 4505 10320
rect 4561 10264 4587 10320
rect 4643 10264 4669 10320
rect 4725 10264 4751 10320
rect 4815 10316 4829 10368
rect 4889 10344 4915 10400
rect 4971 10344 4997 10400
rect 5053 10344 5079 10400
rect 5135 10344 5161 10400
rect 5217 10344 5243 10400
rect 5299 10386 5317 10400
rect 5369 10386 5383 10438
rect 5435 10386 5871 10438
rect 5923 10386 5937 10438
rect 5989 10386 6425 10438
rect 6477 10386 6491 10438
rect 6543 10386 6979 10438
rect 7031 10386 7045 10438
rect 7097 10386 7533 10438
rect 7585 10386 7599 10438
rect 5299 10368 7651 10386
rect 5299 10344 5317 10368
rect 4881 10320 5317 10344
rect 4807 10298 4833 10316
rect 2850 10246 3101 10264
rect 3153 10246 3167 10264
rect 3219 10246 3655 10264
rect 3707 10246 3721 10264
rect 3773 10246 4209 10264
rect 4261 10246 4275 10264
rect 4327 10246 4763 10264
rect 4815 10246 4829 10298
rect 4889 10264 4915 10320
rect 4971 10264 4997 10320
rect 5053 10264 5079 10320
rect 5135 10264 5161 10320
rect 5217 10264 5243 10320
rect 5299 10316 5317 10320
rect 5369 10316 5383 10368
rect 5435 10316 5871 10368
rect 5923 10316 5937 10368
rect 5989 10316 6425 10368
rect 6477 10316 6491 10368
rect 6543 10316 6979 10368
rect 7031 10316 7045 10368
rect 7097 10316 7533 10368
rect 7585 10316 7599 10368
rect 5299 10298 7651 10316
rect 5299 10264 5317 10298
rect 4881 10246 5317 10264
rect 5369 10246 5383 10298
rect 5435 10246 5871 10298
rect 5923 10246 5937 10298
rect 5989 10246 6425 10298
rect 6477 10246 6491 10298
rect 6543 10246 6979 10298
rect 7031 10246 7045 10298
rect 7097 10246 7533 10298
rect 7585 10246 7599 10298
rect 2850 10240 7651 10246
rect 2850 10184 2859 10240
rect 2915 10184 2942 10240
rect 2998 10184 3025 10240
rect 3081 10228 3108 10240
rect 3164 10228 3191 10240
rect 3081 10184 3101 10228
rect 3164 10184 3167 10228
rect 3247 10184 3274 10240
rect 3330 10184 3357 10240
rect 3413 10184 3439 10240
rect 3495 10184 3521 10240
rect 3577 10184 3603 10240
rect 3659 10228 3685 10240
rect 3741 10228 3767 10240
rect 3823 10184 3849 10240
rect 3905 10184 3931 10240
rect 3987 10184 4013 10240
rect 4069 10184 4095 10240
rect 4151 10184 4177 10240
rect 4233 10228 4259 10240
rect 4315 10228 4341 10240
rect 4327 10184 4341 10228
rect 4397 10184 4423 10240
rect 4479 10184 4505 10240
rect 4561 10184 4587 10240
rect 4643 10184 4669 10240
rect 4725 10184 4751 10240
rect 4807 10228 4833 10240
rect 2850 10176 3101 10184
rect 3153 10176 3167 10184
rect 3219 10176 3655 10184
rect 3707 10176 3721 10184
rect 3773 10176 4209 10184
rect 4261 10176 4275 10184
rect 4327 10176 4763 10184
rect 4815 10176 4829 10228
rect 4889 10184 4915 10240
rect 4971 10184 4997 10240
rect 5053 10184 5079 10240
rect 5135 10184 5161 10240
rect 5217 10184 5243 10240
rect 5299 10228 7651 10240
rect 5299 10184 5317 10228
rect 4881 10176 5317 10184
rect 5369 10176 5383 10228
rect 5435 10176 5871 10228
rect 5923 10176 5937 10228
rect 5989 10176 6425 10228
rect 6477 10176 6491 10228
rect 6543 10176 6979 10228
rect 7031 10176 7045 10228
rect 7097 10176 7533 10228
rect 7585 10176 7599 10228
rect 2850 10160 7651 10176
rect 2850 10104 2859 10160
rect 2915 10104 2942 10160
rect 2998 10104 3025 10160
rect 3081 10158 3108 10160
rect 3164 10158 3191 10160
rect 3081 10106 3101 10158
rect 3164 10106 3167 10158
rect 3081 10104 3108 10106
rect 3164 10104 3191 10106
rect 3247 10104 3274 10160
rect 3330 10104 3357 10160
rect 3413 10104 3439 10160
rect 3495 10104 3521 10160
rect 3577 10104 3603 10160
rect 3659 10158 3685 10160
rect 3741 10158 3767 10160
rect 3659 10104 3685 10106
rect 3741 10104 3767 10106
rect 3823 10104 3849 10160
rect 3905 10104 3931 10160
rect 3987 10104 4013 10160
rect 4069 10104 4095 10160
rect 4151 10104 4177 10160
rect 4233 10158 4259 10160
rect 4315 10158 4341 10160
rect 4327 10106 4341 10158
rect 4233 10104 4259 10106
rect 4315 10104 4341 10106
rect 4397 10104 4423 10160
rect 4479 10104 4505 10160
rect 4561 10104 4587 10160
rect 4643 10104 4669 10160
rect 4725 10104 4751 10160
rect 4807 10158 4833 10160
rect 4815 10106 4829 10158
rect 4807 10104 4833 10106
rect 4889 10104 4915 10160
rect 4971 10104 4997 10160
rect 5053 10104 5079 10160
rect 5135 10104 5161 10160
rect 5217 10104 5243 10160
rect 5299 10158 7651 10160
rect 5299 10106 5317 10158
rect 5369 10106 5383 10158
rect 5435 10106 5871 10158
rect 5923 10106 5937 10158
rect 5989 10106 6425 10158
rect 6477 10106 6491 10158
rect 6543 10106 6979 10158
rect 7031 10106 7045 10158
rect 7097 10106 7533 10158
rect 7585 10106 7599 10158
rect 5299 10104 7651 10106
rect 2850 10100 7651 10104
rect 2528 10060 2712 10074
rect 2528 10008 2580 10060
rect 2632 10008 2660 10060
rect 2528 9851 2712 10008
tri 2712 9851 2792 9931 sw
rect 2528 9827 2792 9851
tri 2528 9563 2792 9827 ne
tri 2792 9602 3041 9851 sw
rect 2468 9298 2474 9350
rect 2526 9298 2539 9350
rect 2591 9298 2604 9350
rect 2656 9298 2662 9350
rect 2468 7549 2662 9298
rect 2468 7497 2474 7549
rect 2526 7497 2539 7549
rect 2591 7497 2604 7549
rect 2656 7497 2662 7549
rect 2468 5654 2662 7497
rect 2468 5602 2474 5654
rect 2526 5602 2539 5654
rect 2591 5602 2604 5654
rect 2656 5602 2662 5654
tri 2454 2717 2468 2731 se
rect 2468 2717 2662 5602
tri 2402 2665 2454 2717 se
rect 2454 2665 2662 2717
tri 2386 2649 2402 2665 se
rect 2402 2649 2662 2665
tri 2334 2597 2386 2649 se
rect 2386 2597 2662 2649
tri 2318 2581 2334 2597 se
rect 2334 2595 2662 2597
rect 2334 2581 2648 2595
tri 2648 2581 2662 2595 nw
rect 2792 5557 3041 9602
rect 5198 9458 5617 9460
rect 5673 9458 5698 9460
rect 5754 9458 5779 9460
rect 5835 9458 5860 9460
rect 5916 9458 5941 9460
rect 5997 9458 6022 9460
rect 6078 9458 6103 9460
rect 6159 9458 6184 9460
rect 6240 9458 6265 9460
rect 6321 9458 6346 9460
rect 6402 9458 6427 9460
rect 6483 9458 6508 9460
rect 6564 9458 6589 9460
rect 6645 9458 6669 9460
rect 6725 9458 6749 9460
rect 6805 9458 6829 9460
rect 6885 9458 6909 9460
rect 6965 9458 6989 9460
rect 7045 9458 7069 9460
rect 7125 9458 7149 9460
rect 7205 9458 7229 9460
rect 7285 9458 7309 9460
rect 7365 9458 7374 9460
rect 5198 9406 5204 9458
rect 5256 9406 5268 9458
rect 5320 9406 5332 9458
rect 5384 9406 5396 9458
rect 5448 9406 5460 9458
rect 5512 9406 5524 9458
rect 5576 9406 5588 9458
rect 5768 9406 5779 9458
rect 5835 9406 5844 9458
rect 6088 9406 6100 9458
rect 6159 9406 6164 9458
rect 6344 9406 6346 9458
rect 6408 9406 6420 9458
rect 6483 9406 6484 9458
rect 6664 9406 6669 9458
rect 6728 9406 6740 9458
rect 6984 9406 6989 9458
rect 7048 9406 7060 9458
rect 7304 9406 7309 9458
rect 7368 9406 7374 9458
rect 5198 9404 5617 9406
rect 5673 9404 5698 9406
rect 5754 9404 5779 9406
rect 5835 9404 5860 9406
rect 5916 9404 5941 9406
rect 5997 9404 6022 9406
rect 6078 9404 6103 9406
rect 6159 9404 6184 9406
rect 6240 9404 6265 9406
rect 6321 9404 6346 9406
rect 6402 9404 6427 9406
rect 6483 9404 6508 9406
rect 6564 9404 6589 9406
rect 6645 9404 6669 9406
rect 6725 9404 6749 9406
rect 6805 9404 6829 9406
rect 6885 9404 6909 9406
rect 6965 9404 6989 9406
rect 7045 9404 7069 9406
rect 7125 9404 7149 9406
rect 7205 9404 7229 9406
rect 7285 9404 7309 9406
rect 7365 9404 7374 9406
rect 5198 8727 7374 8728
rect 5198 7843 5204 8727
rect 7368 7843 7374 8727
rect 5198 7842 7374 7843
rect 5198 7690 5617 7692
rect 5673 7690 5698 7692
rect 5754 7690 5779 7692
rect 5835 7690 5860 7692
rect 5916 7690 5941 7692
rect 5997 7690 6022 7692
rect 6078 7690 6103 7692
rect 6159 7690 6184 7692
rect 6240 7690 6265 7692
rect 6321 7690 6346 7692
rect 6402 7690 6427 7692
rect 6483 7690 6508 7692
rect 6564 7690 6589 7692
rect 6645 7690 6669 7692
rect 6725 7690 6749 7692
rect 6805 7690 6829 7692
rect 6885 7690 6909 7692
rect 6965 7690 6989 7692
rect 7045 7690 7069 7692
rect 7125 7690 7149 7692
rect 7205 7690 7229 7692
rect 7285 7690 7309 7692
rect 7365 7690 7374 7692
rect 5198 7638 5204 7690
rect 5256 7638 5268 7690
rect 5320 7638 5332 7690
rect 5384 7638 5396 7690
rect 5448 7638 5460 7690
rect 5512 7638 5524 7690
rect 5576 7638 5588 7690
rect 5768 7638 5779 7690
rect 5835 7638 5844 7690
rect 6088 7638 6100 7690
rect 6159 7638 6164 7690
rect 6344 7638 6346 7690
rect 6408 7638 6420 7690
rect 6483 7638 6484 7690
rect 6664 7638 6669 7690
rect 6728 7638 6740 7690
rect 6984 7638 6989 7690
rect 7048 7638 7060 7690
rect 7304 7638 7309 7690
rect 7368 7638 7374 7690
rect 5198 7636 5617 7638
rect 5673 7636 5698 7638
rect 5754 7636 5779 7638
rect 5835 7636 5860 7638
rect 5916 7636 5941 7638
rect 5997 7636 6022 7638
rect 6078 7636 6103 7638
rect 6159 7636 6184 7638
rect 6240 7636 6265 7638
rect 6321 7636 6346 7638
rect 6402 7636 6427 7638
rect 6483 7636 6508 7638
rect 6564 7636 6589 7638
rect 6645 7636 6669 7638
rect 6725 7636 6749 7638
rect 6805 7636 6829 7638
rect 6885 7636 6909 7638
rect 6965 7636 6989 7638
rect 7045 7636 7069 7638
rect 7125 7636 7149 7638
rect 7205 7636 7229 7638
rect 7285 7636 7309 7638
rect 7365 7636 7374 7638
rect 5198 6927 7374 6928
rect 5198 6043 5204 6927
rect 7368 6043 7374 6927
rect 5198 6042 7374 6043
rect 5198 5850 5617 5852
rect 5673 5850 5698 5852
rect 5754 5850 5779 5852
rect 5835 5850 5860 5852
rect 5916 5850 5941 5852
rect 5997 5850 6022 5852
rect 6078 5850 6103 5852
rect 6159 5850 6184 5852
rect 6240 5850 6265 5852
rect 6321 5850 6346 5852
rect 6402 5850 6427 5852
rect 6483 5850 6508 5852
rect 6564 5850 6589 5852
rect 6645 5850 6669 5852
rect 6725 5850 6749 5852
rect 6805 5850 6829 5852
rect 6885 5850 6909 5852
rect 6965 5850 6989 5852
rect 7045 5850 7069 5852
rect 7125 5850 7149 5852
rect 7205 5850 7229 5852
rect 7285 5850 7309 5852
rect 7365 5850 7374 5852
rect 5198 5798 5204 5850
rect 5256 5798 5268 5850
rect 5320 5798 5332 5850
rect 5384 5798 5396 5850
rect 5448 5798 5460 5850
rect 5512 5798 5524 5850
rect 5576 5798 5588 5850
rect 5768 5798 5779 5850
rect 5835 5798 5844 5850
rect 6088 5798 6100 5850
rect 6159 5798 6164 5850
rect 6344 5798 6346 5850
rect 6408 5798 6420 5850
rect 6483 5798 6484 5850
rect 6664 5798 6669 5850
rect 6728 5798 6740 5850
rect 6984 5798 6989 5850
rect 7048 5798 7060 5850
rect 7304 5798 7309 5850
rect 7368 5798 7374 5850
rect 5198 5796 5617 5798
rect 5673 5796 5698 5798
rect 5754 5796 5779 5798
rect 5835 5796 5860 5798
rect 5916 5796 5941 5798
rect 5997 5796 6022 5798
rect 6078 5796 6103 5798
rect 6159 5796 6184 5798
rect 6240 5796 6265 5798
rect 6321 5796 6346 5798
rect 6402 5796 6427 5798
rect 6483 5796 6508 5798
rect 6564 5796 6589 5798
rect 6645 5796 6669 5798
rect 6725 5796 6749 5798
rect 6805 5796 6829 5798
rect 6885 5796 6909 5798
rect 6965 5796 6989 5798
rect 7045 5796 7069 5798
rect 7125 5796 7149 5798
rect 7205 5796 7229 5798
rect 7285 5796 7309 5798
rect 7365 5796 7374 5798
rect 2792 5505 2798 5557
rect 2850 5505 2891 5557
rect 2943 5505 2983 5557
rect 3035 5505 3041 5557
rect 2792 5479 3041 5505
rect 2792 5427 2798 5479
rect 2850 5427 2891 5479
rect 2943 5427 2983 5479
rect 3035 5427 3041 5479
tri 2266 2529 2318 2581 se
rect 2318 2529 2596 2581
tri 2596 2529 2648 2581 nw
tri 2250 2513 2266 2529 se
rect 2266 2513 2580 2529
tri 2580 2513 2596 2529 nw
tri 2198 2461 2250 2513 se
rect 2250 2461 2528 2513
tri 2528 2461 2580 2513 nw
tri 2138 2401 2198 2461 se
rect 2198 2401 2468 2461
tri 2468 2401 2528 2461 nw
tri 2000 2263 2138 2401 se
rect 2138 2263 2330 2401
tri 2330 2263 2468 2401 nw
tri 1971 2234 2000 2263 se
rect 2000 2234 2278 2263
rect 1971 2211 2278 2234
tri 2278 2211 2330 2263 nw
rect 1971 2197 2264 2211
tri 2264 2197 2278 2211 nw
rect 1971 2150 2212 2197
rect 1971 2098 1977 2150
rect 2029 2098 2042 2150
rect 2094 2098 2107 2150
rect 2159 2145 2212 2150
tri 2212 2145 2264 2197 nw
rect 2159 2131 2198 2145
tri 2198 2131 2212 2145 nw
rect 2159 2098 2165 2131
tri 2165 2098 2198 2131 nw
rect 2792 1834 3041 5427
rect 5198 4743 7374 4747
rect 5198 4691 5204 4743
rect 5256 4691 5336 4743
rect 5388 4691 5468 4743
rect 5520 4691 5600 4743
rect 5652 4741 5732 4743
rect 5784 4741 5864 4743
rect 5916 4741 5996 4743
rect 6048 4741 6128 4743
rect 6180 4741 6260 4743
rect 6312 4741 6392 4743
rect 6444 4741 6524 4743
rect 6576 4741 6656 4743
rect 6708 4741 6788 4743
rect 6840 4741 6920 4743
rect 6972 4741 7052 4743
rect 7104 4741 7184 4743
rect 7236 4741 7316 4743
rect 5198 4685 5623 4691
rect 5679 4685 5704 4741
rect 5784 4691 5785 4741
rect 5760 4685 5785 4691
rect 5841 4691 5864 4741
rect 5841 4685 5866 4691
rect 5922 4685 5947 4741
rect 6003 4685 6027 4691
rect 6083 4685 6107 4741
rect 6180 4691 6187 4741
rect 6163 4685 6187 4691
rect 6243 4691 6260 4741
rect 6243 4685 6267 4691
rect 6323 4685 6347 4741
rect 6403 4685 6427 4691
rect 6483 4685 6507 4741
rect 6576 4691 6587 4741
rect 6563 4685 6587 4691
rect 6643 4691 6656 4741
rect 6643 4685 6667 4691
rect 6723 4685 6747 4741
rect 6803 4685 6827 4691
rect 6883 4685 6907 4741
rect 6972 4691 6987 4741
rect 6963 4685 6987 4691
rect 7043 4691 7052 4741
rect 7043 4685 7067 4691
rect 7123 4685 7147 4741
rect 7203 4685 7227 4691
rect 7283 4685 7307 4741
rect 7368 4691 7374 4743
rect 7363 4685 7374 4691
rect 5198 4653 7374 4685
rect 5198 4635 5623 4653
rect 5198 4583 5204 4635
rect 5256 4583 5336 4635
rect 5388 4583 5468 4635
rect 5520 4583 5600 4635
rect 5679 4597 5704 4653
rect 5760 4635 5785 4653
rect 5784 4597 5785 4635
rect 5841 4635 5866 4653
rect 5841 4597 5864 4635
rect 5922 4597 5947 4653
rect 6003 4635 6027 4653
rect 6083 4597 6107 4653
rect 6163 4635 6187 4653
rect 6180 4597 6187 4635
rect 6243 4635 6267 4653
rect 6243 4597 6260 4635
rect 6323 4597 6347 4653
rect 6403 4635 6427 4653
rect 6483 4597 6507 4653
rect 6563 4635 6587 4653
rect 6576 4597 6587 4635
rect 6643 4635 6667 4653
rect 6643 4597 6656 4635
rect 6723 4597 6747 4653
rect 6803 4635 6827 4653
rect 6883 4597 6907 4653
rect 6963 4635 6987 4653
rect 6972 4597 6987 4635
rect 7043 4635 7067 4653
rect 7043 4597 7052 4635
rect 7123 4597 7147 4653
rect 7203 4635 7227 4653
rect 7283 4597 7307 4653
rect 7363 4635 7374 4653
rect 5652 4583 5732 4597
rect 5784 4583 5864 4597
rect 5916 4583 5996 4597
rect 6048 4583 6128 4597
rect 6180 4583 6260 4597
rect 6312 4583 6392 4597
rect 6444 4583 6524 4597
rect 6576 4583 6656 4597
rect 6708 4583 6788 4597
rect 6840 4583 6920 4597
rect 6972 4583 7052 4597
rect 7104 4583 7184 4597
rect 7236 4583 7316 4597
rect 7368 4583 7374 4635
rect 5198 4565 7374 4583
rect 5198 4527 5623 4565
rect 5198 4475 5204 4527
rect 5256 4475 5336 4527
rect 5388 4475 5468 4527
rect 5520 4475 5600 4527
rect 5679 4509 5704 4565
rect 5760 4527 5785 4565
rect 5784 4509 5785 4527
rect 5841 4527 5866 4565
rect 5841 4509 5864 4527
rect 5922 4509 5947 4565
rect 6003 4527 6027 4565
rect 6083 4509 6107 4565
rect 6163 4527 6187 4565
rect 6180 4509 6187 4527
rect 6243 4527 6267 4565
rect 6243 4509 6260 4527
rect 6323 4509 6347 4565
rect 6403 4527 6427 4565
rect 6483 4509 6507 4565
rect 6563 4527 6587 4565
rect 6576 4509 6587 4527
rect 6643 4527 6667 4565
rect 6643 4509 6656 4527
rect 6723 4509 6747 4565
rect 6803 4527 6827 4565
rect 6883 4509 6907 4565
rect 6963 4527 6987 4565
rect 6972 4509 6987 4527
rect 7043 4527 7067 4565
rect 7043 4509 7052 4527
rect 7123 4509 7147 4565
rect 7203 4527 7227 4565
rect 7283 4509 7307 4565
rect 7363 4527 7374 4565
rect 5652 4477 5732 4509
rect 5784 4477 5864 4509
rect 5916 4477 5996 4509
rect 6048 4477 6128 4509
rect 6180 4477 6260 4509
rect 6312 4477 6392 4509
rect 6444 4477 6524 4509
rect 6576 4477 6656 4509
rect 6708 4477 6788 4509
rect 6840 4477 6920 4509
rect 6972 4477 7052 4509
rect 7104 4477 7184 4509
rect 7236 4477 7316 4509
rect 5198 4421 5623 4475
rect 5679 4421 5704 4477
rect 5784 4475 5785 4477
rect 5760 4421 5785 4475
rect 5841 4475 5864 4477
rect 5841 4421 5866 4475
rect 5922 4421 5947 4477
rect 6003 4421 6027 4475
rect 6083 4421 6107 4477
rect 6180 4475 6187 4477
rect 6163 4421 6187 4475
rect 6243 4475 6260 4477
rect 6243 4421 6267 4475
rect 6323 4421 6347 4477
rect 6403 4421 6427 4475
rect 6483 4421 6507 4477
rect 6576 4475 6587 4477
rect 6563 4421 6587 4475
rect 6643 4475 6656 4477
rect 6643 4421 6667 4475
rect 6723 4421 6747 4477
rect 6803 4421 6827 4475
rect 6883 4421 6907 4477
rect 6972 4475 6987 4477
rect 6963 4421 6987 4475
rect 7043 4475 7052 4477
rect 7043 4421 7067 4475
rect 7123 4421 7147 4477
rect 7203 4421 7227 4475
rect 7283 4421 7307 4477
rect 7368 4475 7374 4527
rect 7363 4421 7374 4475
rect 5198 4419 7374 4421
rect 5198 4367 5204 4419
rect 5256 4367 5336 4419
rect 5388 4367 5468 4419
rect 5520 4367 5600 4419
rect 5652 4389 5732 4419
rect 5784 4389 5864 4419
rect 5916 4389 5996 4419
rect 6048 4389 6128 4419
rect 6180 4389 6260 4419
rect 6312 4389 6392 4419
rect 6444 4389 6524 4419
rect 6576 4389 6656 4419
rect 6708 4389 6788 4419
rect 6840 4389 6920 4419
rect 6972 4389 7052 4419
rect 7104 4389 7184 4419
rect 7236 4389 7316 4419
rect 5198 4333 5623 4367
rect 5679 4333 5704 4389
rect 5784 4367 5785 4389
rect 5760 4333 5785 4367
rect 5841 4367 5864 4389
rect 5841 4333 5866 4367
rect 5922 4333 5947 4389
rect 6003 4333 6027 4367
rect 6083 4333 6107 4389
rect 6180 4367 6187 4389
rect 6163 4333 6187 4367
rect 6243 4367 6260 4389
rect 6243 4333 6267 4367
rect 6323 4333 6347 4389
rect 6403 4333 6427 4367
rect 6483 4333 6507 4389
rect 6576 4367 6587 4389
rect 6563 4333 6587 4367
rect 6643 4367 6656 4389
rect 6643 4333 6667 4367
rect 6723 4333 6747 4389
rect 6803 4333 6827 4367
rect 6883 4333 6907 4389
rect 6972 4367 6987 4389
rect 6963 4333 6987 4367
rect 7043 4367 7052 4389
rect 7043 4333 7067 4367
rect 7123 4333 7147 4389
rect 7203 4333 7227 4367
rect 7283 4333 7307 4389
rect 7368 4367 7374 4419
rect 7363 4333 7374 4367
rect 5198 4311 7374 4333
rect 5198 4259 5204 4311
rect 5256 4259 5336 4311
rect 5388 4259 5468 4311
rect 5520 4259 5600 4311
rect 5652 4301 5732 4311
rect 5784 4301 5864 4311
rect 5916 4301 5996 4311
rect 6048 4301 6128 4311
rect 6180 4301 6260 4311
rect 6312 4301 6392 4311
rect 6444 4301 6524 4311
rect 6576 4301 6656 4311
rect 6708 4301 6788 4311
rect 6840 4301 6920 4311
rect 6972 4301 7052 4311
rect 7104 4301 7184 4311
rect 7236 4301 7316 4311
rect 5198 4245 5623 4259
rect 5679 4245 5704 4301
rect 5784 4259 5785 4301
rect 5760 4245 5785 4259
rect 5841 4259 5864 4301
rect 5841 4245 5866 4259
rect 5922 4245 5947 4301
rect 6003 4245 6027 4259
rect 6083 4245 6107 4301
rect 6180 4259 6187 4301
rect 6163 4245 6187 4259
rect 6243 4259 6260 4301
rect 6243 4245 6267 4259
rect 6323 4245 6347 4301
rect 6403 4245 6427 4259
rect 6483 4245 6507 4301
rect 6576 4259 6587 4301
rect 6563 4245 6587 4259
rect 6643 4259 6656 4301
rect 6643 4245 6667 4259
rect 6723 4245 6747 4301
rect 6803 4245 6827 4259
rect 6883 4245 6907 4301
rect 6972 4259 6987 4301
rect 6963 4245 6987 4259
rect 7043 4259 7052 4301
rect 7043 4245 7067 4259
rect 7123 4245 7147 4301
rect 7203 4245 7227 4259
rect 7283 4245 7307 4301
rect 7368 4259 7374 4311
rect 7363 4245 7374 4259
rect 5198 4213 7374 4245
rect 5198 4203 5623 4213
rect 5198 4151 5204 4203
rect 5256 4151 5336 4203
rect 5388 4151 5468 4203
rect 5520 4151 5600 4203
rect 5679 4157 5704 4213
rect 5760 4203 5785 4213
rect 5784 4157 5785 4203
rect 5841 4203 5866 4213
rect 5841 4157 5864 4203
rect 5922 4157 5947 4213
rect 6003 4203 6027 4213
rect 6083 4157 6107 4213
rect 6163 4203 6187 4213
rect 6180 4157 6187 4203
rect 6243 4203 6267 4213
rect 6243 4157 6260 4203
rect 6323 4157 6347 4213
rect 6403 4203 6427 4213
rect 6483 4157 6507 4213
rect 6563 4203 6587 4213
rect 6576 4157 6587 4203
rect 6643 4203 6667 4213
rect 6643 4157 6656 4203
rect 6723 4157 6747 4213
rect 6803 4203 6827 4213
rect 6883 4157 6907 4213
rect 6963 4203 6987 4213
rect 6972 4157 6987 4203
rect 7043 4203 7067 4213
rect 7043 4157 7052 4203
rect 7123 4157 7147 4213
rect 7203 4203 7227 4213
rect 7283 4157 7307 4213
rect 7363 4203 7374 4213
rect 5652 4151 5732 4157
rect 5784 4151 5864 4157
rect 5916 4151 5996 4157
rect 6048 4151 6128 4157
rect 6180 4151 6260 4157
rect 6312 4151 6392 4157
rect 6444 4151 6524 4157
rect 6576 4151 6656 4157
rect 6708 4151 6788 4157
rect 6840 4151 6920 4157
rect 6972 4151 7052 4157
rect 7104 4151 7184 4157
rect 7236 4151 7316 4157
rect 7368 4151 7374 4203
rect 5198 4147 7374 4151
rect 5198 3897 5204 3949
rect 5256 3897 5339 3949
rect 5391 3897 5474 3949
rect 5526 3897 5609 3949
rect 5661 3918 5744 3949
rect 5796 3918 5879 3949
rect 5931 3918 6014 3949
rect 6066 3918 6149 3949
rect 6201 3918 6284 3949
rect 6336 3918 6419 3949
rect 6471 3918 6553 3949
rect 6605 3918 6687 3949
rect 6739 3918 6821 3949
rect 6873 3918 6955 3949
rect 7007 3918 7089 3949
rect 7141 3918 7223 3949
rect 7275 3918 7374 3949
rect 5198 3883 5617 3897
rect 5198 3831 5204 3883
rect 5256 3831 5339 3883
rect 5391 3831 5474 3883
rect 5526 3831 5609 3883
rect 5673 3862 5698 3918
rect 5754 3883 5779 3897
rect 5835 3862 5860 3918
rect 5931 3897 5941 3918
rect 5916 3883 5941 3897
rect 5931 3862 5941 3883
rect 5997 3897 6014 3918
rect 5997 3883 6022 3897
rect 5997 3862 6014 3883
rect 6078 3862 6103 3918
rect 6159 3883 6184 3897
rect 6240 3862 6265 3918
rect 6336 3897 6346 3918
rect 6321 3883 6346 3897
rect 6336 3862 6346 3883
rect 6402 3897 6419 3918
rect 6402 3883 6427 3897
rect 6402 3862 6419 3883
rect 6483 3862 6508 3918
rect 6564 3883 6589 3897
rect 6645 3862 6669 3918
rect 6739 3897 6749 3918
rect 6725 3883 6749 3897
rect 6739 3862 6749 3883
rect 6805 3897 6821 3918
rect 6805 3883 6829 3897
rect 6805 3862 6821 3883
rect 6885 3862 6909 3918
rect 6965 3883 6989 3897
rect 7045 3862 7069 3918
rect 7141 3897 7149 3918
rect 7125 3883 7149 3897
rect 7141 3862 7149 3883
rect 7205 3897 7223 3918
rect 7205 3883 7229 3897
rect 7205 3862 7223 3883
rect 7285 3862 7309 3918
rect 7365 3862 7374 3918
rect 5661 3831 5744 3862
rect 5796 3831 5879 3862
rect 5931 3831 6014 3862
rect 6066 3831 6149 3862
rect 6201 3831 6284 3862
rect 6336 3831 6419 3862
rect 6471 3831 6553 3862
rect 6605 3831 6687 3862
rect 6739 3831 6821 3862
rect 6873 3831 6955 3862
rect 7007 3831 7089 3862
rect 7141 3831 7223 3862
rect 7275 3831 7374 3862
rect 5198 3057 7542 3058
rect 5198 3005 5204 3057
rect 5256 3005 5270 3057
rect 5322 3005 5336 3057
rect 5388 3005 5402 3057
rect 5454 3005 5468 3057
rect 5520 3005 5534 3057
rect 5586 3005 5599 3057
rect 5846 3005 5859 3057
rect 5916 3005 5924 3057
rect 6171 3005 6184 3057
rect 6240 3005 6249 3057
rect 6496 3005 6508 3057
rect 6564 3005 6574 3057
rect 6821 3005 6832 3057
rect 6888 3005 6899 3057
rect 7146 3005 7156 3057
rect 7212 3005 7224 3057
rect 7471 3005 7477 3057
rect 7536 3005 7542 3057
rect 5198 3001 5617 3005
rect 5673 3001 5698 3005
rect 5754 3001 5779 3005
rect 5835 3001 5860 3005
rect 5916 3001 5941 3005
rect 5997 3001 6022 3005
rect 6078 3001 6103 3005
rect 6159 3001 6184 3005
rect 6240 3001 6265 3005
rect 6321 3001 6346 3005
rect 6402 3001 6427 3005
rect 6483 3001 6508 3005
rect 6564 3001 6589 3005
rect 6645 3001 6670 3005
rect 6726 3001 6751 3005
rect 6807 3001 6832 3005
rect 6888 3001 6913 3005
rect 6969 3001 6994 3005
rect 7050 3001 7075 3005
rect 7131 3001 7156 3005
rect 7212 3001 7237 3005
rect 7293 3001 7317 3005
rect 7373 3001 7397 3005
rect 7453 3001 7477 3005
rect 7533 3001 7542 3005
rect 5198 2989 7542 3001
rect 5198 2937 5204 2989
rect 5256 2937 5270 2989
rect 5322 2937 5336 2989
rect 5388 2937 5402 2989
rect 5454 2937 5468 2989
rect 5520 2937 5534 2989
rect 5586 2937 5599 2989
rect 5651 2967 5664 2989
rect 5716 2967 5729 2989
rect 5781 2967 5794 2989
rect 5846 2937 5859 2989
rect 5911 2967 5924 2989
rect 5976 2967 5989 2989
rect 6041 2967 6054 2989
rect 6106 2967 6119 2989
rect 5916 2937 5924 2967
rect 6171 2937 6184 2989
rect 6236 2967 6249 2989
rect 6301 2967 6314 2989
rect 6366 2967 6379 2989
rect 6431 2967 6444 2989
rect 6496 2967 6509 2989
rect 6561 2967 6574 2989
rect 6626 2967 6639 2989
rect 6691 2967 6704 2989
rect 6756 2967 6769 2989
rect 6821 2967 6834 2989
rect 6886 2967 6899 2989
rect 6951 2967 6964 2989
rect 7016 2967 7029 2989
rect 7081 2967 7094 2989
rect 7146 2967 7159 2989
rect 7211 2967 7224 2989
rect 7276 2967 7289 2989
rect 7341 2967 7354 2989
rect 7406 2967 7419 2989
rect 7471 2967 7484 2989
rect 6240 2937 6249 2967
rect 6496 2937 6508 2967
rect 6564 2937 6574 2967
rect 6821 2937 6832 2967
rect 6888 2937 6899 2967
rect 7146 2937 7156 2967
rect 7212 2937 7224 2967
rect 7471 2937 7477 2967
rect 7536 2937 7542 2989
rect 5198 2921 5617 2937
rect 5673 2921 5698 2937
rect 5754 2921 5779 2937
rect 5835 2921 5860 2937
rect 5916 2921 5941 2937
rect 5997 2921 6022 2937
rect 6078 2921 6103 2937
rect 6159 2921 6184 2937
rect 6240 2921 6265 2937
rect 6321 2921 6346 2937
rect 6402 2921 6427 2937
rect 6483 2921 6508 2937
rect 6564 2921 6589 2937
rect 6645 2921 6670 2937
rect 6726 2921 6751 2937
rect 6807 2921 6832 2937
rect 6888 2921 6913 2937
rect 6969 2921 6994 2937
rect 7050 2921 7075 2937
rect 7131 2921 7156 2937
rect 7212 2921 7237 2937
rect 7293 2921 7317 2937
rect 7373 2921 7397 2937
rect 7453 2921 7477 2937
rect 7533 2921 7542 2937
rect 5198 2869 5204 2921
rect 5256 2869 5270 2921
rect 5322 2869 5336 2921
rect 5388 2869 5402 2921
rect 5454 2869 5468 2921
rect 5520 2869 5534 2921
rect 5586 2869 5599 2921
rect 5651 2877 5664 2911
rect 5716 2877 5729 2911
rect 5781 2877 5794 2911
rect 5846 2869 5859 2921
rect 5916 2911 5924 2921
rect 5911 2877 5924 2911
rect 5976 2877 5989 2911
rect 6041 2877 6054 2911
rect 6106 2877 6119 2911
rect 5916 2869 5924 2877
rect 6171 2869 6184 2921
rect 6240 2911 6249 2921
rect 6496 2911 6508 2921
rect 6564 2911 6574 2921
rect 6821 2911 6832 2921
rect 6888 2911 6899 2921
rect 7146 2911 7156 2921
rect 7212 2911 7224 2921
rect 7471 2911 7477 2921
rect 6236 2877 6249 2911
rect 6301 2877 6314 2911
rect 6366 2877 6379 2911
rect 6431 2877 6444 2911
rect 6496 2877 6509 2911
rect 6561 2877 6574 2911
rect 6626 2877 6639 2911
rect 6691 2877 6704 2911
rect 6756 2877 6769 2911
rect 6821 2877 6834 2911
rect 6886 2877 6899 2911
rect 6951 2877 6964 2911
rect 7016 2877 7029 2911
rect 7081 2877 7094 2911
rect 7146 2877 7159 2911
rect 7211 2877 7224 2911
rect 7276 2877 7289 2911
rect 7341 2877 7354 2911
rect 7406 2877 7419 2911
rect 7471 2877 7484 2911
rect 6240 2869 6249 2877
rect 6496 2869 6508 2877
rect 6564 2869 6574 2877
rect 6821 2869 6832 2877
rect 6888 2869 6899 2877
rect 7146 2869 7156 2877
rect 7212 2869 7224 2877
rect 7471 2869 7477 2877
rect 7536 2869 7542 2921
rect 5198 2853 5617 2869
rect 5673 2853 5698 2869
rect 5754 2853 5779 2869
rect 5835 2853 5860 2869
rect 5916 2853 5941 2869
rect 5997 2853 6022 2869
rect 6078 2853 6103 2869
rect 6159 2853 6184 2869
rect 6240 2853 6265 2869
rect 6321 2853 6346 2869
rect 6402 2853 6427 2869
rect 6483 2853 6508 2869
rect 6564 2853 6589 2869
rect 6645 2853 6670 2869
rect 6726 2853 6751 2869
rect 6807 2853 6832 2869
rect 6888 2853 6913 2869
rect 6969 2853 6994 2869
rect 7050 2853 7075 2869
rect 7131 2853 7156 2869
rect 7212 2853 7237 2869
rect 7293 2853 7317 2869
rect 7373 2853 7397 2869
rect 7453 2853 7477 2869
rect 7533 2853 7542 2869
rect 5198 2801 5204 2853
rect 5256 2801 5270 2853
rect 5322 2801 5336 2853
rect 5388 2801 5402 2853
rect 5454 2801 5468 2853
rect 5520 2801 5534 2853
rect 5586 2801 5599 2853
rect 5651 2801 5664 2821
rect 5716 2801 5729 2821
rect 5781 2801 5794 2821
rect 5846 2801 5859 2853
rect 5916 2821 5924 2853
rect 5911 2801 5924 2821
rect 5976 2801 5989 2821
rect 6041 2801 6054 2821
rect 6106 2801 6119 2821
rect 6171 2801 6184 2853
rect 6240 2821 6249 2853
rect 6496 2821 6508 2853
rect 6564 2821 6574 2853
rect 6821 2821 6832 2853
rect 6888 2821 6899 2853
rect 7146 2821 7156 2853
rect 7212 2821 7224 2853
rect 7471 2821 7477 2853
rect 6236 2801 6249 2821
rect 6301 2801 6314 2821
rect 6366 2801 6379 2821
rect 6431 2801 6444 2821
rect 6496 2801 6509 2821
rect 6561 2801 6574 2821
rect 6626 2801 6639 2821
rect 6691 2801 6704 2821
rect 6756 2801 6769 2821
rect 6821 2801 6834 2821
rect 6886 2801 6899 2821
rect 6951 2801 6964 2821
rect 7016 2801 7029 2821
rect 7081 2801 7094 2821
rect 7146 2801 7159 2821
rect 7211 2801 7224 2821
rect 7276 2801 7289 2821
rect 7341 2801 7354 2821
rect 7406 2801 7419 2821
rect 7471 2801 7484 2821
rect 7536 2801 7542 2853
rect 5198 2787 7542 2801
rect 5198 2785 5617 2787
rect 5673 2785 5698 2787
rect 5754 2785 5779 2787
rect 5835 2785 5860 2787
rect 5916 2785 5941 2787
rect 5997 2785 6022 2787
rect 6078 2785 6103 2787
rect 6159 2785 6184 2787
rect 6240 2785 6265 2787
rect 6321 2785 6346 2787
rect 6402 2785 6427 2787
rect 6483 2785 6508 2787
rect 6564 2785 6589 2787
rect 6645 2785 6670 2787
rect 6726 2785 6751 2787
rect 6807 2785 6832 2787
rect 6888 2785 6913 2787
rect 6969 2785 6994 2787
rect 7050 2785 7075 2787
rect 7131 2785 7156 2787
rect 7212 2785 7237 2787
rect 7293 2785 7317 2787
rect 7373 2785 7397 2787
rect 7453 2785 7477 2787
rect 7533 2785 7542 2787
rect 5198 2733 5204 2785
rect 5256 2733 5270 2785
rect 5322 2733 5336 2785
rect 5388 2733 5402 2785
rect 5454 2733 5468 2785
rect 5520 2733 5534 2785
rect 5586 2733 5599 2785
rect 5846 2733 5859 2785
rect 5916 2733 5924 2785
rect 6171 2733 6184 2785
rect 6240 2733 6249 2785
rect 6496 2733 6508 2785
rect 6564 2733 6574 2785
rect 6821 2733 6832 2785
rect 6888 2733 6899 2785
rect 7146 2733 7156 2785
rect 7212 2733 7224 2785
rect 7471 2733 7477 2785
rect 7536 2733 7542 2785
rect 5198 2731 5617 2733
rect 5673 2731 5698 2733
rect 5754 2731 5779 2733
rect 5835 2731 5860 2733
rect 5916 2731 5941 2733
rect 5997 2731 6022 2733
rect 6078 2731 6103 2733
rect 6159 2731 6184 2733
rect 6240 2731 6265 2733
rect 6321 2731 6346 2733
rect 6402 2731 6427 2733
rect 6483 2731 6508 2733
rect 6564 2731 6589 2733
rect 6645 2731 6670 2733
rect 6726 2731 6751 2733
rect 6807 2731 6832 2733
rect 6888 2731 6913 2733
rect 6969 2731 6994 2733
rect 7050 2731 7075 2733
rect 7131 2731 7156 2733
rect 7212 2731 7237 2733
rect 7293 2731 7317 2733
rect 7373 2731 7397 2733
rect 7453 2731 7477 2733
rect 7533 2731 7542 2733
rect 5198 2717 7542 2731
rect 5198 2665 5204 2717
rect 5256 2665 5270 2717
rect 5322 2665 5336 2717
rect 5388 2665 5402 2717
rect 5454 2665 5468 2717
rect 5520 2665 5534 2717
rect 5586 2665 5599 2717
rect 5651 2697 5664 2717
rect 5716 2697 5729 2717
rect 5781 2697 5794 2717
rect 5846 2665 5859 2717
rect 5911 2697 5924 2717
rect 5976 2697 5989 2717
rect 6041 2697 6054 2717
rect 6106 2697 6119 2717
rect 5916 2665 5924 2697
rect 6171 2665 6184 2717
rect 6236 2697 6249 2717
rect 6301 2697 6314 2717
rect 6366 2697 6379 2717
rect 6431 2697 6444 2717
rect 6496 2697 6509 2717
rect 6561 2697 6574 2717
rect 6626 2697 6639 2717
rect 6691 2697 6704 2717
rect 6756 2697 6769 2717
rect 6821 2697 6834 2717
rect 6886 2697 6899 2717
rect 6951 2697 6964 2717
rect 7016 2697 7029 2717
rect 7081 2697 7094 2717
rect 7146 2697 7159 2717
rect 7211 2697 7224 2717
rect 7276 2697 7289 2717
rect 7341 2697 7354 2717
rect 7406 2697 7419 2717
rect 7471 2697 7484 2717
rect 6240 2665 6249 2697
rect 6496 2665 6508 2697
rect 6564 2665 6574 2697
rect 6821 2665 6832 2697
rect 6888 2665 6899 2697
rect 7146 2665 7156 2697
rect 7212 2665 7224 2697
rect 7471 2665 7477 2697
rect 7536 2665 7542 2717
rect 5198 2649 5617 2665
rect 5673 2649 5698 2665
rect 5754 2649 5779 2665
rect 5835 2649 5860 2665
rect 5916 2649 5941 2665
rect 5997 2649 6022 2665
rect 6078 2649 6103 2665
rect 6159 2649 6184 2665
rect 6240 2649 6265 2665
rect 6321 2649 6346 2665
rect 6402 2649 6427 2665
rect 6483 2649 6508 2665
rect 6564 2649 6589 2665
rect 6645 2649 6670 2665
rect 6726 2649 6751 2665
rect 6807 2649 6832 2665
rect 6888 2649 6913 2665
rect 6969 2649 6994 2665
rect 7050 2649 7075 2665
rect 7131 2649 7156 2665
rect 7212 2649 7237 2665
rect 7293 2649 7317 2665
rect 7373 2649 7397 2665
rect 7453 2649 7477 2665
rect 7533 2649 7542 2665
rect 5198 2597 5204 2649
rect 5256 2597 5270 2649
rect 5322 2597 5336 2649
rect 5388 2597 5402 2649
rect 5454 2597 5468 2649
rect 5520 2597 5534 2649
rect 5586 2597 5599 2649
rect 5651 2607 5664 2641
rect 5716 2607 5729 2641
rect 5781 2607 5794 2641
rect 5846 2597 5859 2649
rect 5916 2641 5924 2649
rect 5911 2607 5924 2641
rect 5976 2607 5989 2641
rect 6041 2607 6054 2641
rect 6106 2607 6119 2641
rect 5916 2597 5924 2607
rect 6171 2597 6184 2649
rect 6240 2641 6249 2649
rect 6496 2641 6508 2649
rect 6564 2641 6574 2649
rect 6821 2641 6832 2649
rect 6888 2641 6899 2649
rect 7146 2641 7156 2649
rect 7212 2641 7224 2649
rect 7471 2641 7477 2649
rect 6236 2607 6249 2641
rect 6301 2607 6314 2641
rect 6366 2607 6379 2641
rect 6431 2607 6444 2641
rect 6496 2607 6509 2641
rect 6561 2607 6574 2641
rect 6626 2607 6639 2641
rect 6691 2607 6704 2641
rect 6756 2607 6769 2641
rect 6821 2607 6834 2641
rect 6886 2607 6899 2641
rect 6951 2607 6964 2641
rect 7016 2607 7029 2641
rect 7081 2607 7094 2641
rect 7146 2607 7159 2641
rect 7211 2607 7224 2641
rect 7276 2607 7289 2641
rect 7341 2607 7354 2641
rect 7406 2607 7419 2641
rect 7471 2607 7484 2641
rect 6240 2597 6249 2607
rect 6496 2597 6508 2607
rect 6564 2597 6574 2607
rect 6821 2597 6832 2607
rect 6888 2597 6899 2607
rect 7146 2597 7156 2607
rect 7212 2597 7224 2607
rect 7471 2597 7477 2607
rect 7536 2597 7542 2649
rect 5198 2581 5617 2597
rect 5673 2581 5698 2597
rect 5754 2581 5779 2597
rect 5835 2581 5860 2597
rect 5916 2581 5941 2597
rect 5997 2581 6022 2597
rect 6078 2581 6103 2597
rect 6159 2581 6184 2597
rect 6240 2581 6265 2597
rect 6321 2581 6346 2597
rect 6402 2581 6427 2597
rect 6483 2581 6508 2597
rect 6564 2581 6589 2597
rect 6645 2581 6670 2597
rect 6726 2581 6751 2597
rect 6807 2581 6832 2597
rect 6888 2581 6913 2597
rect 6969 2581 6994 2597
rect 7050 2581 7075 2597
rect 7131 2581 7156 2597
rect 7212 2581 7237 2597
rect 7293 2581 7317 2597
rect 7373 2581 7397 2597
rect 7453 2581 7477 2597
rect 7533 2581 7542 2597
rect 5198 2529 5204 2581
rect 5256 2529 5270 2581
rect 5322 2529 5336 2581
rect 5388 2529 5402 2581
rect 5454 2529 5468 2581
rect 5520 2529 5534 2581
rect 5586 2529 5599 2581
rect 5651 2529 5664 2551
rect 5716 2529 5729 2551
rect 5781 2529 5794 2551
rect 5846 2529 5859 2581
rect 5916 2551 5924 2581
rect 5911 2529 5924 2551
rect 5976 2529 5989 2551
rect 6041 2529 6054 2551
rect 6106 2529 6119 2551
rect 6171 2529 6184 2581
rect 6240 2551 6249 2581
rect 6496 2551 6508 2581
rect 6564 2551 6574 2581
rect 6821 2551 6832 2581
rect 6888 2551 6899 2581
rect 7146 2551 7156 2581
rect 7212 2551 7224 2581
rect 7471 2551 7477 2581
rect 6236 2529 6249 2551
rect 6301 2529 6314 2551
rect 6366 2529 6379 2551
rect 6431 2529 6444 2551
rect 6496 2529 6509 2551
rect 6561 2529 6574 2551
rect 6626 2529 6639 2551
rect 6691 2529 6704 2551
rect 6756 2529 6769 2551
rect 6821 2529 6834 2551
rect 6886 2529 6899 2551
rect 6951 2529 6964 2551
rect 7016 2529 7029 2551
rect 7081 2529 7094 2551
rect 7146 2529 7159 2551
rect 7211 2529 7224 2551
rect 7276 2529 7289 2551
rect 7341 2529 7354 2551
rect 7406 2529 7419 2551
rect 7471 2529 7484 2551
rect 7536 2529 7542 2581
rect 5198 2517 7542 2529
rect 5198 2513 5617 2517
rect 5673 2513 5698 2517
rect 5754 2513 5779 2517
rect 5835 2513 5860 2517
rect 5916 2513 5941 2517
rect 5997 2513 6022 2517
rect 6078 2513 6103 2517
rect 6159 2513 6184 2517
rect 6240 2513 6265 2517
rect 6321 2513 6346 2517
rect 6402 2513 6427 2517
rect 6483 2513 6508 2517
rect 6564 2513 6589 2517
rect 6645 2513 6670 2517
rect 6726 2513 6751 2517
rect 6807 2513 6832 2517
rect 6888 2513 6913 2517
rect 6969 2513 6994 2517
rect 7050 2513 7075 2517
rect 7131 2513 7156 2517
rect 7212 2513 7237 2517
rect 7293 2513 7317 2517
rect 7373 2513 7397 2517
rect 7453 2513 7477 2517
rect 7533 2513 7542 2517
rect 5198 2461 5204 2513
rect 5256 2461 5270 2513
rect 5322 2461 5336 2513
rect 5388 2461 5402 2513
rect 5454 2461 5468 2513
rect 5520 2461 5534 2513
rect 5586 2461 5599 2513
rect 5846 2461 5859 2513
rect 5916 2461 5924 2513
rect 6171 2461 6184 2513
rect 6240 2461 6249 2513
rect 6496 2461 6508 2513
rect 6564 2461 6574 2513
rect 6821 2461 6832 2513
rect 6888 2461 6899 2513
rect 7146 2461 7156 2513
rect 7212 2461 7224 2513
rect 7471 2461 7477 2513
rect 7536 2461 7542 2513
rect 5198 2460 7542 2461
rect 3186 2264 5307 2267
rect 3186 2263 3195 2264
rect 3251 2263 3277 2264
rect 3333 2263 3359 2264
rect 3415 2263 3441 2264
rect 3497 2263 3523 2264
rect 3579 2263 3605 2264
rect 3661 2263 3687 2264
rect 3743 2263 3769 2264
rect 3825 2263 3851 2264
rect 3907 2263 3933 2264
rect 3989 2263 4015 2264
rect 4071 2263 4097 2264
rect 4153 2263 4179 2264
rect 4235 2263 4261 2264
rect 4317 2263 4343 2264
rect 4399 2263 4425 2264
rect 4481 2263 4507 2264
rect 4563 2263 4589 2264
rect 4645 2263 4671 2264
rect 4727 2263 4753 2264
rect 4809 2263 4835 2264
rect 4891 2263 4917 2264
rect 3186 2211 3192 2263
rect 3251 2211 3258 2263
rect 3508 2211 3522 2263
rect 3579 2211 3588 2263
rect 3838 2211 3851 2263
rect 3907 2211 3918 2263
rect 4168 2211 4179 2263
rect 4235 2211 4248 2263
rect 4498 2211 4507 2263
rect 4564 2211 4578 2263
rect 4828 2211 4835 2263
rect 4893 2211 4917 2263
rect 3186 2208 3195 2211
rect 3251 2208 3277 2211
rect 3333 2208 3359 2211
rect 3415 2208 3441 2211
rect 3497 2208 3523 2211
rect 3579 2208 3605 2211
rect 3661 2208 3687 2211
rect 3743 2208 3769 2211
rect 3825 2208 3851 2211
rect 3907 2208 3933 2211
rect 3989 2208 4015 2211
rect 4071 2208 4097 2211
rect 4153 2208 4179 2211
rect 4235 2208 4261 2211
rect 4317 2208 4343 2211
rect 4399 2208 4425 2211
rect 4481 2208 4507 2211
rect 4563 2208 4589 2211
rect 4645 2208 4671 2211
rect 4727 2208 4753 2211
rect 4809 2208 4835 2211
rect 4891 2208 4917 2211
rect 4973 2208 4999 2264
rect 5055 2208 5080 2264
rect 5136 2208 5161 2264
rect 5217 2208 5242 2264
rect 5298 2208 5307 2264
rect 6608 2242 7366 2248
rect 3186 2197 5307 2208
rect 3186 2145 3192 2197
rect 3244 2182 3258 2197
rect 3310 2182 3324 2197
rect 3376 2182 3390 2197
rect 3442 2182 3456 2197
rect 3251 2145 3258 2182
rect 3508 2145 3522 2197
rect 3574 2182 3588 2197
rect 3640 2182 3654 2197
rect 3706 2182 3720 2197
rect 3772 2182 3786 2197
rect 3838 2182 3852 2197
rect 3904 2182 3918 2197
rect 3970 2182 3984 2197
rect 4036 2182 4050 2197
rect 4102 2182 4116 2197
rect 4168 2182 4182 2197
rect 4234 2182 4248 2197
rect 4300 2182 4314 2197
rect 4366 2182 4380 2197
rect 4432 2182 4446 2197
rect 4498 2182 4512 2197
rect 3579 2145 3588 2182
rect 3838 2145 3851 2182
rect 3907 2145 3918 2182
rect 4168 2145 4179 2182
rect 4235 2145 4248 2182
rect 4498 2145 4507 2182
rect 4564 2145 4578 2197
rect 4630 2182 4644 2197
rect 4696 2182 4710 2197
rect 4762 2182 4776 2197
rect 4828 2182 4841 2197
rect 4893 2182 5307 2197
rect 4828 2145 4835 2182
rect 4893 2145 4917 2182
rect 3186 2131 3195 2145
rect 3251 2131 3277 2145
rect 3333 2131 3359 2145
rect 3415 2131 3441 2145
rect 3497 2131 3523 2145
rect 3579 2131 3605 2145
rect 3661 2131 3687 2145
rect 3743 2131 3769 2145
rect 3825 2131 3851 2145
rect 3907 2131 3933 2145
rect 3989 2131 4015 2145
rect 4071 2131 4097 2145
rect 4153 2131 4179 2145
rect 4235 2131 4261 2145
rect 4317 2131 4343 2145
rect 4399 2131 4425 2145
rect 4481 2131 4507 2145
rect 4563 2131 4589 2145
rect 4645 2131 4671 2145
rect 4727 2131 4753 2145
rect 4809 2131 4835 2145
rect 4891 2131 4917 2145
rect 3186 2079 3192 2131
rect 3251 2126 3258 2131
rect 3244 2100 3258 2126
rect 3310 2100 3324 2126
rect 3376 2100 3390 2126
rect 3442 2100 3456 2126
rect 3251 2079 3258 2100
rect 3508 2079 3522 2131
rect 3579 2126 3588 2131
rect 3838 2126 3851 2131
rect 3907 2126 3918 2131
rect 4168 2126 4179 2131
rect 4235 2126 4248 2131
rect 4498 2126 4507 2131
rect 3574 2100 3588 2126
rect 3640 2100 3654 2126
rect 3706 2100 3720 2126
rect 3772 2100 3786 2126
rect 3838 2100 3852 2126
rect 3904 2100 3918 2126
rect 3970 2100 3984 2126
rect 4036 2100 4050 2126
rect 4102 2100 4116 2126
rect 4168 2100 4182 2126
rect 4234 2100 4248 2126
rect 4300 2100 4314 2126
rect 4366 2100 4380 2126
rect 4432 2100 4446 2126
rect 4498 2100 4512 2126
rect 3579 2079 3588 2100
rect 3838 2079 3851 2100
rect 3907 2079 3918 2100
rect 4168 2079 4179 2100
rect 4235 2079 4248 2100
rect 4498 2079 4507 2100
rect 4564 2079 4578 2131
rect 4828 2126 4835 2131
rect 4893 2126 4917 2131
rect 4973 2126 4999 2182
rect 5055 2126 5080 2182
rect 5136 2126 5161 2182
rect 5217 2126 5242 2182
rect 5298 2126 5307 2182
rect 4630 2100 4644 2126
rect 4696 2100 4710 2126
rect 4762 2100 4776 2126
rect 4828 2100 4841 2126
rect 4893 2100 5307 2126
rect 4828 2079 4835 2100
rect 4893 2079 4917 2100
rect 3186 2065 3195 2079
rect 3251 2065 3277 2079
rect 3333 2065 3359 2079
rect 3415 2065 3441 2079
rect 3497 2065 3523 2079
rect 3579 2065 3605 2079
rect 3661 2065 3687 2079
rect 3743 2065 3769 2079
rect 3825 2065 3851 2079
rect 3907 2065 3933 2079
rect 3989 2065 4015 2079
rect 4071 2065 4097 2079
rect 4153 2065 4179 2079
rect 4235 2065 4261 2079
rect 4317 2065 4343 2079
rect 4399 2065 4425 2079
rect 4481 2065 4507 2079
rect 4563 2065 4589 2079
rect 4645 2065 4671 2079
rect 4727 2065 4753 2079
rect 4809 2065 4835 2079
rect 4891 2065 4917 2079
rect 3186 2013 3192 2065
rect 3251 2044 3258 2065
rect 3244 2018 3258 2044
rect 3310 2018 3324 2044
rect 3376 2018 3390 2044
rect 3442 2018 3456 2044
rect 3251 2013 3258 2018
rect 3508 2013 3522 2065
rect 3579 2044 3588 2065
rect 3838 2044 3851 2065
rect 3907 2044 3918 2065
rect 4168 2044 4179 2065
rect 4235 2044 4248 2065
rect 4498 2044 4507 2065
rect 3574 2018 3588 2044
rect 3640 2018 3654 2044
rect 3706 2018 3720 2044
rect 3772 2018 3786 2044
rect 3838 2018 3852 2044
rect 3904 2018 3918 2044
rect 3970 2018 3984 2044
rect 4036 2018 4050 2044
rect 4102 2018 4116 2044
rect 4168 2018 4182 2044
rect 4234 2018 4248 2044
rect 4300 2018 4314 2044
rect 4366 2018 4380 2044
rect 4432 2018 4446 2044
rect 4498 2018 4512 2044
rect 3579 2013 3588 2018
rect 3838 2013 3851 2018
rect 3907 2013 3918 2018
rect 4168 2013 4179 2018
rect 4235 2013 4248 2018
rect 4498 2013 4507 2018
rect 4564 2013 4578 2065
rect 4828 2044 4835 2065
rect 4893 2044 4917 2065
rect 4973 2044 4999 2100
rect 5055 2044 5080 2100
rect 5136 2044 5161 2100
rect 5217 2044 5242 2100
rect 5298 2044 5307 2100
rect 4630 2018 4644 2044
rect 4696 2018 4710 2044
rect 4762 2018 4776 2044
rect 4828 2018 4841 2044
rect 4893 2018 5307 2044
rect 4828 2013 4835 2018
rect 4893 2013 4917 2018
rect 3186 1999 3195 2013
rect 3251 1999 3277 2013
rect 3333 1999 3359 2013
rect 3415 1999 3441 2013
rect 3497 1999 3523 2013
rect 3579 1999 3605 2013
rect 3661 1999 3687 2013
rect 3743 1999 3769 2013
rect 3825 1999 3851 2013
rect 3907 1999 3933 2013
rect 3989 1999 4015 2013
rect 4071 1999 4097 2013
rect 4153 1999 4179 2013
rect 4235 1999 4261 2013
rect 4317 1999 4343 2013
rect 4399 1999 4425 2013
rect 4481 1999 4507 2013
rect 4563 1999 4589 2013
rect 4645 1999 4671 2013
rect 4727 1999 4753 2013
rect 4809 1999 4835 2013
rect 4891 1999 4917 2013
rect 3186 1947 3192 1999
rect 3251 1962 3258 1999
rect 3244 1947 3258 1962
rect 3310 1947 3324 1962
rect 3376 1947 3390 1962
rect 3442 1947 3456 1962
rect 3508 1947 3522 1999
rect 3579 1962 3588 1999
rect 3838 1962 3851 1999
rect 3907 1962 3918 1999
rect 4168 1962 4179 1999
rect 4235 1962 4248 1999
rect 4498 1962 4507 1999
rect 3574 1947 3588 1962
rect 3640 1947 3654 1962
rect 3706 1947 3720 1962
rect 3772 1947 3786 1962
rect 3838 1947 3852 1962
rect 3904 1947 3918 1962
rect 3970 1947 3984 1962
rect 4036 1947 4050 1962
rect 4102 1947 4116 1962
rect 4168 1947 4182 1962
rect 4234 1947 4248 1962
rect 4300 1947 4314 1962
rect 4366 1947 4380 1962
rect 4432 1947 4446 1962
rect 4498 1947 4512 1962
rect 4564 1947 4578 1999
rect 4828 1962 4835 1999
rect 4893 1962 4917 1999
rect 4973 1962 4999 2018
rect 5055 1962 5080 2018
rect 5136 1962 5161 2018
rect 5217 1962 5242 2018
rect 5298 1962 5307 2018
rect 4630 1947 4644 1962
rect 4696 1947 4710 1962
rect 4762 1947 4776 1962
rect 4828 1947 4841 1962
rect 4893 1947 5307 1962
rect 3186 1936 5307 1947
rect 3186 1933 3195 1936
rect 3251 1933 3277 1936
rect 3333 1933 3359 1936
rect 3415 1933 3441 1936
rect 3497 1933 3523 1936
rect 3579 1933 3605 1936
rect 3661 1933 3687 1936
rect 3743 1933 3769 1936
rect 3825 1933 3851 1936
rect 3907 1933 3933 1936
rect 3989 1933 4015 1936
rect 4071 1933 4097 1936
rect 4153 1933 4179 1936
rect 4235 1933 4261 1936
rect 4317 1933 4343 1936
rect 4399 1933 4425 1936
rect 4481 1933 4507 1936
rect 4563 1933 4589 1936
rect 4645 1933 4671 1936
rect 4727 1933 4753 1936
rect 4809 1933 4835 1936
rect 4891 1933 4917 1936
rect 3186 1881 3192 1933
rect 3251 1881 3258 1933
rect 3508 1881 3522 1933
rect 3579 1881 3588 1933
rect 3838 1881 3851 1933
rect 3907 1881 3918 1933
rect 4168 1881 4179 1933
rect 4235 1881 4248 1933
rect 4498 1881 4507 1933
rect 4564 1881 4578 1933
rect 4828 1881 4835 1933
rect 4893 1881 4917 1933
rect 3186 1880 3195 1881
rect 3251 1880 3277 1881
rect 3333 1880 3359 1881
rect 3415 1880 3441 1881
rect 3497 1880 3523 1881
rect 3579 1880 3605 1881
rect 3661 1880 3687 1881
rect 3743 1880 3769 1881
rect 3825 1880 3851 1881
rect 3907 1880 3933 1881
rect 3989 1880 4015 1881
rect 4071 1880 4097 1881
rect 4153 1880 4179 1881
rect 4235 1880 4261 1881
rect 4317 1880 4343 1881
rect 4399 1880 4425 1881
rect 4481 1880 4507 1881
rect 4563 1880 4589 1881
rect 4645 1880 4671 1881
rect 4727 1880 4753 1881
rect 4809 1880 4835 1881
rect 4891 1880 4917 1881
rect 4973 1880 4999 1936
rect 5055 1880 5080 1936
rect 5136 1880 5161 1936
rect 5217 1880 5242 1936
rect 5298 1880 5307 1936
rect 3186 1877 5307 1880
rect 5624 2228 6320 2234
rect 5624 2225 5628 2228
rect 5624 2143 5628 2169
rect 5624 2061 5628 2087
rect 5624 1979 5628 2005
rect 5624 1897 5628 1923
rect 2792 1782 2798 1834
rect 2850 1782 2891 1834
rect 2943 1782 2983 1834
rect 3035 1782 3041 1834
rect 2792 1650 3041 1782
rect 2792 1598 2798 1650
rect 2850 1598 2891 1650
rect 2943 1598 2983 1650
rect 3035 1598 3041 1650
rect 2792 1467 3041 1598
rect 2792 1415 2798 1467
rect 2850 1415 2891 1467
rect 2943 1415 2983 1467
rect 3035 1415 3041 1467
rect 2792 1282 3041 1415
rect 2792 1230 2798 1282
rect 2850 1230 2891 1282
rect 2943 1230 2983 1282
rect 3035 1230 3041 1282
rect 2792 1098 3041 1230
rect 2792 1046 2798 1098
rect 2850 1046 2891 1098
rect 2943 1046 2983 1098
rect 3035 1046 3041 1098
rect 5624 1815 5628 1841
rect 5624 1733 5628 1759
rect 5624 1651 5628 1677
rect 5624 1569 5628 1595
rect 5624 1487 5628 1513
rect 5624 1405 5628 1431
rect 5624 1323 5628 1349
rect 5624 1241 5628 1267
rect 5624 1159 5628 1185
rect 5680 1139 5704 1152
rect 5760 1139 5784 1152
rect 5840 1139 5864 1152
rect 5920 1139 5944 1152
rect 6000 1139 6024 1152
rect 6080 1139 6104 1152
rect 6160 1139 6184 1152
rect 6240 1139 6264 1152
rect 5624 1087 5628 1103
rect 5680 1087 5692 1139
rect 5936 1103 5944 1139
rect 5744 1087 5756 1103
rect 5808 1087 5820 1103
rect 5872 1087 5884 1103
rect 5936 1087 5948 1103
rect 6000 1087 6012 1139
rect 6256 1103 6264 1139
rect 6064 1087 6076 1103
rect 6128 1087 6140 1103
rect 6192 1087 6204 1103
rect 6256 1087 6268 1103
rect 5624 1077 6320 1087
rect 5680 1074 5704 1077
rect 5760 1074 5784 1077
rect 5840 1074 5864 1077
rect 5920 1074 5944 1077
rect 6000 1074 6024 1077
rect 6080 1074 6104 1077
rect 6160 1074 6184 1077
rect 6240 1074 6264 1077
rect 5680 1022 5692 1074
rect 5936 1022 5944 1074
rect 6000 1022 6012 1074
rect 6256 1022 6264 1074
rect 5680 1021 5704 1022
rect 5760 1021 5784 1022
rect 5840 1021 5864 1022
rect 5920 1021 5944 1022
rect 6000 1021 6024 1022
rect 6080 1021 6104 1022
rect 6160 1021 6184 1022
rect 6240 1021 6264 1022
rect 5624 1009 6320 1021
rect 5624 994 5628 1009
rect 5680 957 5692 1009
rect 5744 994 5756 1009
rect 5808 994 5820 1009
rect 5872 994 5884 1009
rect 5936 994 5948 1009
rect 5936 957 5944 994
rect 6000 957 6012 1009
rect 6064 994 6076 1009
rect 6128 994 6140 1009
rect 6192 994 6204 1009
rect 6256 994 6268 1009
rect 6256 957 6264 994
rect 5680 944 5704 957
rect 5760 944 5784 957
rect 5840 944 5864 957
rect 5920 944 5944 957
rect 6000 944 6024 957
rect 6080 944 6104 957
rect 6160 944 6184 957
rect 6240 944 6264 957
rect 5624 911 5628 938
rect 5680 892 5692 944
rect 5936 938 5944 944
rect 5744 911 5756 938
rect 5808 911 5820 938
rect 5872 911 5884 938
rect 5936 911 5948 938
rect 5936 892 5944 911
rect 6000 892 6012 944
rect 6256 938 6264 944
rect 6064 911 6076 938
rect 6128 911 6140 938
rect 6192 911 6204 938
rect 6256 911 6268 938
rect 6256 892 6264 911
rect 5680 879 5704 892
rect 5760 879 5784 892
rect 5840 879 5864 892
rect 5920 879 5944 892
rect 6000 879 6024 892
rect 6080 879 6104 892
rect 6160 879 6184 892
rect 6240 879 6264 892
rect 5624 828 5628 855
rect 5680 827 5692 879
rect 5936 855 5944 879
rect 5744 828 5756 855
rect 5808 828 5820 855
rect 5872 828 5884 855
rect 5936 828 5948 855
rect 5936 827 5944 828
rect 6000 827 6012 879
rect 6256 855 6264 879
rect 6064 828 6076 855
rect 6128 828 6140 855
rect 6192 828 6204 855
rect 6256 828 6268 855
rect 6256 827 6264 828
rect 5680 814 5704 827
rect 5760 814 5784 827
rect 5840 814 5864 827
rect 5920 814 5944 827
rect 6000 814 6024 827
rect 6080 814 6104 827
rect 6160 814 6184 827
rect 6240 814 6264 827
rect 5624 762 5628 772
rect 5680 762 5692 814
rect 5936 772 5944 814
rect 5744 762 5756 772
rect 5808 762 5820 772
rect 5872 762 5884 772
rect 5936 762 5948 772
rect 6000 762 6012 814
rect 6256 772 6264 814
rect 6064 762 6076 772
rect 6128 762 6140 772
rect 6192 762 6204 772
rect 6256 762 6268 772
rect 5624 749 6320 762
rect 5624 745 5628 749
rect 5680 697 5692 749
rect 5744 745 5756 749
rect 5808 745 5820 749
rect 5872 745 5884 749
rect 5936 745 5948 749
rect 5936 697 5944 745
rect 6000 697 6012 749
rect 6064 745 6076 749
rect 6128 745 6140 749
rect 6192 745 6204 749
rect 6256 745 6268 749
rect 6256 697 6264 745
rect 5680 689 5704 697
rect 5760 689 5784 697
rect 5840 689 5864 697
rect 5920 689 5944 697
rect 6000 689 6024 697
rect 6080 689 6104 697
rect 6160 689 6184 697
rect 6240 689 6264 697
rect 5624 684 6320 689
rect 5624 662 5628 684
rect 5680 632 5692 684
rect 5744 662 5756 684
rect 5808 662 5820 684
rect 5872 662 5884 684
rect 5936 662 5948 684
rect 5936 632 5944 662
rect 6000 632 6012 684
rect 6064 662 6076 684
rect 6128 662 6140 684
rect 6192 662 6204 684
rect 6256 662 6268 684
rect 6256 632 6264 662
rect 5680 619 5704 632
rect 5760 619 5784 632
rect 5840 619 5864 632
rect 5920 619 5944 632
rect 6000 619 6024 632
rect 6080 619 6104 632
rect 6160 619 6184 632
rect 6240 619 6264 632
rect 5624 579 5628 606
rect 5680 567 5692 619
rect 5936 606 5944 619
rect 5744 579 5756 606
rect 5808 579 5820 606
rect 5872 579 5884 606
rect 5936 579 5948 606
rect 5936 567 5944 579
rect 6000 567 6012 619
rect 6256 606 6264 619
rect 6064 579 6076 606
rect 6128 579 6140 606
rect 6192 579 6204 606
rect 6256 579 6268 606
rect 6256 567 6264 579
rect 5680 554 5704 567
rect 5760 554 5784 567
rect 5840 554 5864 567
rect 5920 554 5944 567
rect 6000 554 6024 567
rect 6080 554 6104 567
rect 6160 554 6184 567
rect 6240 554 6264 567
rect 5624 502 5628 523
rect 5680 502 5692 554
rect 5936 523 5944 554
rect 5744 502 5756 523
rect 5808 502 5820 523
rect 5872 502 5884 523
rect 5936 502 5948 523
rect 6000 502 6012 554
rect 6256 523 6264 554
rect 6064 502 6076 523
rect 6128 502 6140 523
rect 6192 502 6204 523
rect 6256 502 6268 523
rect 5624 496 6320 502
rect 5680 489 5704 496
rect 5760 489 5784 496
rect 5840 489 5864 496
rect 5920 489 5944 496
rect 6000 489 6024 496
rect 6080 489 6104 496
rect 6160 489 6184 496
rect 6240 489 6264 496
rect 5624 437 5628 440
rect 5680 437 5692 489
rect 5936 440 5944 489
rect 5744 437 5756 440
rect 5808 437 5820 440
rect 5872 437 5884 440
rect 5936 437 5948 440
rect 6000 437 6012 489
rect 6256 440 6264 489
rect 6064 437 6076 440
rect 6128 437 6140 440
rect 6192 437 6204 440
rect 6256 437 6268 440
rect 5624 431 6320 437
rect 6608 2190 6611 2242
rect 6663 2239 6711 2242
rect 6763 2239 6811 2242
rect 6863 2239 6911 2242
rect 6963 2239 7011 2242
rect 7063 2239 7111 2242
rect 7163 2239 7211 2242
rect 7263 2239 7311 2242
rect 6608 2183 6615 2190
rect 6671 2183 6701 2239
rect 6763 2190 6787 2239
rect 6863 2190 6873 2239
rect 7101 2190 7111 2239
rect 7187 2190 7211 2239
rect 6757 2183 6787 2190
rect 6843 2183 6873 2190
rect 6929 2183 6959 2190
rect 7015 2183 7045 2190
rect 7101 2183 7131 2190
rect 7187 2183 7217 2190
rect 7273 2183 7303 2239
rect 7363 2190 7366 2242
rect 7359 2183 7366 2190
rect 6608 2157 7366 2183
rect 6608 2108 6615 2157
rect 6608 2056 6611 2108
rect 6671 2101 6701 2157
rect 6757 2108 6787 2157
rect 6843 2108 6873 2157
rect 6929 2108 6959 2157
rect 7015 2108 7045 2157
rect 7101 2108 7131 2157
rect 7187 2108 7217 2157
rect 6763 2101 6787 2108
rect 6863 2101 6873 2108
rect 7101 2101 7111 2108
rect 7187 2101 7211 2108
rect 7273 2101 7303 2157
rect 7359 2108 7366 2157
rect 6663 2075 6711 2101
rect 6763 2075 6811 2101
rect 6863 2075 6911 2101
rect 6963 2075 7011 2101
rect 7063 2075 7111 2101
rect 7163 2075 7211 2101
rect 7263 2075 7311 2101
rect 6608 2019 6615 2056
rect 6671 2019 6701 2075
rect 6763 2056 6787 2075
rect 6863 2056 6873 2075
rect 7101 2056 7111 2075
rect 7187 2056 7211 2075
rect 6757 2019 6787 2056
rect 6843 2019 6873 2056
rect 6929 2019 6959 2056
rect 7015 2019 7045 2056
rect 7101 2019 7131 2056
rect 7187 2019 7217 2056
rect 7273 2019 7303 2075
rect 7363 2056 7366 2108
rect 7359 2019 7366 2056
rect 6608 1993 7366 2019
rect 6608 1973 6615 1993
rect 6608 1921 6611 1973
rect 6671 1937 6701 1993
rect 6757 1973 6787 1993
rect 6843 1973 6873 1993
rect 6929 1973 6959 1993
rect 7015 1973 7045 1993
rect 7101 1973 7131 1993
rect 7187 1973 7217 1993
rect 6763 1937 6787 1973
rect 6863 1937 6873 1973
rect 7101 1937 7111 1973
rect 7187 1937 7211 1973
rect 7273 1937 7303 1993
rect 7359 1973 7366 1993
rect 6663 1921 6711 1937
rect 6763 1921 6811 1937
rect 6863 1921 6911 1937
rect 6963 1921 7011 1937
rect 7063 1921 7111 1937
rect 7163 1921 7211 1937
rect 7263 1921 7311 1937
rect 7363 1921 7366 1973
rect 6608 1911 7366 1921
rect 6608 1855 6615 1911
rect 6671 1855 6701 1911
rect 6757 1855 6787 1911
rect 6843 1855 6873 1911
rect 6929 1855 6959 1911
rect 7015 1855 7045 1911
rect 7101 1855 7131 1911
rect 7187 1855 7217 1911
rect 7273 1855 7303 1911
rect 7359 1855 7366 1911
rect 6608 1838 7366 1855
rect 6608 1786 6611 1838
rect 6663 1828 6711 1838
rect 6763 1828 6811 1838
rect 6863 1828 6911 1838
rect 6963 1828 7011 1838
rect 7063 1828 7111 1838
rect 7163 1828 7211 1838
rect 7263 1828 7311 1838
rect 6608 1772 6615 1786
rect 6671 1772 6701 1828
rect 6763 1786 6787 1828
rect 6863 1786 6873 1828
rect 7101 1786 7111 1828
rect 7187 1786 7211 1828
rect 6757 1772 6787 1786
rect 6843 1772 6873 1786
rect 6929 1772 6959 1786
rect 7015 1772 7045 1786
rect 7101 1772 7131 1786
rect 7187 1772 7217 1786
rect 7273 1772 7303 1828
rect 7363 1786 7366 1838
rect 7359 1772 7366 1786
rect 6608 1745 7366 1772
rect 6608 1703 6615 1745
rect 6608 1651 6611 1703
rect 6671 1689 6701 1745
rect 6757 1703 6787 1745
rect 6843 1703 6873 1745
rect 6929 1703 6959 1745
rect 7015 1703 7045 1745
rect 7101 1703 7131 1745
rect 7187 1703 7217 1745
rect 6763 1689 6787 1703
rect 6863 1689 6873 1703
rect 7101 1689 7111 1703
rect 7187 1689 7211 1703
rect 7273 1689 7303 1745
rect 7359 1703 7366 1745
rect 6663 1662 6711 1689
rect 6763 1662 6811 1689
rect 6863 1662 6911 1689
rect 6963 1662 7011 1689
rect 7063 1662 7111 1689
rect 7163 1662 7211 1689
rect 7263 1662 7311 1689
rect 6608 1606 6615 1651
rect 6671 1606 6701 1662
rect 6763 1651 6787 1662
rect 6863 1651 6873 1662
rect 7101 1651 7111 1662
rect 7187 1651 7211 1662
rect 6757 1606 6787 1651
rect 6843 1606 6873 1651
rect 6929 1606 6959 1651
rect 7015 1606 7045 1651
rect 7101 1606 7131 1651
rect 7187 1606 7217 1651
rect 7273 1606 7303 1662
rect 7363 1651 7366 1703
rect 7359 1606 7366 1651
rect 6608 1579 7366 1606
rect 6608 1568 6615 1579
rect 6608 1516 6611 1568
rect 6671 1523 6701 1579
rect 6757 1568 6787 1579
rect 6843 1568 6873 1579
rect 6929 1568 6959 1579
rect 7015 1568 7045 1579
rect 7101 1568 7131 1579
rect 7187 1568 7217 1579
rect 6763 1523 6787 1568
rect 6863 1523 6873 1568
rect 7101 1523 7111 1568
rect 7187 1523 7211 1568
rect 7273 1523 7303 1579
rect 7359 1568 7366 1579
rect 6663 1516 6711 1523
rect 6763 1516 6811 1523
rect 6863 1516 6911 1523
rect 6963 1516 7011 1523
rect 7063 1516 7111 1523
rect 7163 1516 7211 1523
rect 7263 1516 7311 1523
rect 7363 1516 7366 1568
rect 6608 1496 7366 1516
rect 6608 1440 6615 1496
rect 6671 1440 6701 1496
rect 6757 1440 6787 1496
rect 6843 1440 6873 1496
rect 6929 1440 6959 1496
rect 7015 1440 7045 1496
rect 7101 1440 7131 1496
rect 7187 1440 7217 1496
rect 7273 1440 7303 1496
rect 7359 1440 7366 1496
rect 6608 1433 7366 1440
rect 6608 1381 6611 1433
rect 6663 1413 6711 1433
rect 6763 1413 6811 1433
rect 6863 1413 6911 1433
rect 6963 1413 7011 1433
rect 7063 1413 7111 1433
rect 7163 1413 7211 1433
rect 7263 1413 7311 1433
rect 6608 1357 6615 1381
rect 6671 1357 6701 1413
rect 6763 1381 6787 1413
rect 6863 1381 6873 1413
rect 7101 1381 7111 1413
rect 7187 1381 7211 1413
rect 6757 1357 6787 1381
rect 6843 1357 6873 1381
rect 6929 1357 6959 1381
rect 7015 1357 7045 1381
rect 7101 1357 7131 1381
rect 7187 1357 7217 1381
rect 7273 1357 7303 1413
rect 7363 1381 7366 1433
rect 7359 1357 7366 1381
rect 6608 1330 7366 1357
rect 6608 1298 6615 1330
rect 6608 1246 6611 1298
rect 6671 1274 6701 1330
rect 6757 1298 6787 1330
rect 6843 1298 6873 1330
rect 6929 1298 6959 1330
rect 7015 1298 7045 1330
rect 7101 1298 7131 1330
rect 7187 1298 7217 1330
rect 6763 1274 6787 1298
rect 6863 1274 6873 1298
rect 7101 1274 7111 1298
rect 7187 1274 7211 1298
rect 7273 1274 7303 1330
rect 7359 1298 7366 1330
rect 6663 1247 6711 1274
rect 6763 1247 6811 1274
rect 6863 1247 6911 1274
rect 6963 1247 7011 1274
rect 7063 1247 7111 1274
rect 7163 1247 7211 1274
rect 7263 1247 7311 1274
rect 6608 1191 6615 1246
rect 6671 1191 6701 1247
rect 6763 1246 6787 1247
rect 6863 1246 6873 1247
rect 7101 1246 7111 1247
rect 7187 1246 7211 1247
rect 6757 1191 6787 1246
rect 6843 1191 6873 1246
rect 6929 1191 6959 1246
rect 7015 1191 7045 1246
rect 7101 1191 7131 1246
rect 7187 1191 7217 1246
rect 7273 1191 7303 1247
rect 7363 1246 7366 1298
rect 7359 1191 7366 1246
rect 6608 1164 7366 1191
rect 6608 1163 6615 1164
rect 6608 1111 6611 1163
rect 6608 1108 6615 1111
rect 6671 1108 6701 1164
rect 6757 1163 6787 1164
rect 6843 1163 6873 1164
rect 6929 1163 6959 1164
rect 7015 1163 7045 1164
rect 7101 1163 7131 1164
rect 7187 1163 7217 1164
rect 6763 1111 6787 1163
rect 6863 1111 6873 1163
rect 7101 1111 7111 1163
rect 7187 1111 7211 1163
rect 6757 1108 6787 1111
rect 6843 1108 6873 1111
rect 6929 1108 6959 1111
rect 7015 1108 7045 1111
rect 7101 1108 7131 1111
rect 7187 1108 7217 1111
rect 7273 1108 7303 1164
rect 7359 1163 7366 1164
rect 7363 1111 7366 1163
rect 7359 1108 7366 1111
rect 6608 1081 7366 1108
rect 6608 1028 6615 1081
rect 6608 976 6611 1028
rect 6671 1025 6701 1081
rect 6757 1028 6787 1081
rect 6843 1028 6873 1081
rect 6929 1028 6959 1081
rect 7015 1028 7045 1081
rect 7101 1028 7131 1081
rect 7187 1028 7217 1081
rect 6763 1025 6787 1028
rect 6863 1025 6873 1028
rect 7101 1025 7111 1028
rect 7187 1025 7211 1028
rect 7273 1025 7303 1081
rect 7359 1028 7366 1081
rect 6663 998 6711 1025
rect 6763 998 6811 1025
rect 6863 998 6911 1025
rect 6963 998 7011 1025
rect 7063 998 7111 1025
rect 7163 998 7211 1025
rect 7263 998 7311 1025
rect 6608 942 6615 976
rect 6671 942 6701 998
rect 6763 976 6787 998
rect 6863 976 6873 998
rect 7101 976 7111 998
rect 7187 976 7211 998
rect 6757 942 6787 976
rect 6843 942 6873 976
rect 6929 942 6959 976
rect 7015 942 7045 976
rect 7101 942 7131 976
rect 7187 942 7217 976
rect 7273 942 7303 998
rect 7363 976 7366 1028
rect 7359 942 7366 976
rect 6608 915 7366 942
rect 6608 893 6615 915
rect 6608 841 6611 893
rect 6671 859 6701 915
rect 6757 893 6787 915
rect 6843 893 6873 915
rect 6929 893 6959 915
rect 7015 893 7045 915
rect 7101 893 7131 915
rect 7187 893 7217 915
rect 6763 859 6787 893
rect 6863 859 6873 893
rect 7101 859 7111 893
rect 7187 859 7211 893
rect 7273 859 7303 915
rect 7359 893 7366 915
rect 6663 841 6711 859
rect 6763 841 6811 859
rect 6863 841 6911 859
rect 6963 841 7011 859
rect 7063 841 7111 859
rect 7163 841 7211 859
rect 7263 841 7311 859
rect 7363 841 7366 893
rect 6608 832 7366 841
rect 6608 776 6615 832
rect 6671 776 6701 832
rect 6757 776 6787 832
rect 6843 776 6873 832
rect 6929 776 6959 832
rect 7015 776 7045 832
rect 7101 776 7131 832
rect 7187 776 7217 832
rect 7273 776 7303 832
rect 7359 776 7366 832
rect 6608 758 7366 776
rect 6608 706 6611 758
rect 6663 749 6711 758
rect 6763 749 6811 758
rect 6863 749 6911 758
rect 6963 749 7011 758
rect 7063 749 7111 758
rect 7163 749 7211 758
rect 7263 749 7311 758
rect 6608 693 6615 706
rect 6671 693 6701 749
rect 6763 706 6787 749
rect 6863 706 6873 749
rect 7101 706 7111 749
rect 7187 706 7211 749
rect 6757 693 6787 706
rect 6843 693 6873 706
rect 6929 693 6959 706
rect 7015 693 7045 706
rect 7101 693 7131 706
rect 7187 693 7217 706
rect 7273 693 7303 749
rect 7363 706 7366 758
rect 7359 693 7366 706
rect 6608 666 7366 693
rect 6608 623 6615 666
rect 6608 571 6611 623
rect 6671 610 6701 666
rect 6757 623 6787 666
rect 6843 623 6873 666
rect 6929 623 6959 666
rect 7015 623 7045 666
rect 7101 623 7131 666
rect 7187 623 7217 666
rect 6763 610 6787 623
rect 6863 610 6873 623
rect 7101 610 7111 623
rect 7187 610 7211 623
rect 7273 610 7303 666
rect 7359 623 7366 666
rect 6663 583 6711 610
rect 6763 583 6811 610
rect 6863 583 6911 610
rect 6963 583 7011 610
rect 7063 583 7111 610
rect 7163 583 7211 610
rect 7263 583 7311 610
rect 6608 527 6615 571
rect 6671 527 6701 583
rect 6763 571 6787 583
rect 6863 571 6873 583
rect 7101 571 7111 583
rect 7187 571 7211 583
rect 6757 527 6787 571
rect 6843 527 6873 571
rect 6929 527 6959 571
rect 7015 527 7045 571
rect 7101 527 7131 571
rect 7187 527 7217 571
rect 7273 527 7303 583
rect 7363 571 7366 623
rect 7359 527 7366 571
rect 6608 500 7366 527
rect 6608 488 6615 500
rect 6608 436 6611 488
rect 6671 444 6701 500
rect 6757 488 6787 500
rect 6843 488 6873 500
rect 6929 488 6959 500
rect 7015 488 7045 500
rect 7101 488 7131 500
rect 7187 488 7217 500
rect 6763 444 6787 488
rect 6863 444 6873 488
rect 7101 444 7111 488
rect 7187 444 7211 488
rect 7273 444 7303 500
rect 7359 488 7366 500
rect 6663 436 6711 444
rect 6763 436 6811 444
rect 6863 436 6911 444
rect 6963 436 7011 444
rect 7063 436 7111 444
rect 7163 436 7211 444
rect 7263 436 7311 444
rect 7363 436 7366 488
rect 6608 430 7366 436
<< via2 >>
rect 5613 38720 5669 38724
rect 5696 38720 5752 38724
rect 5613 38668 5646 38720
rect 5646 38668 5660 38720
rect 5660 38668 5669 38720
rect 5696 38668 5712 38720
rect 5712 38668 5752 38720
rect 5779 38668 5835 38724
rect 5861 38668 5917 38724
rect 5943 38668 5999 38724
rect 6025 38668 6081 38724
rect 6107 38720 6163 38724
rect 6189 38720 6245 38724
rect 6107 38668 6148 38720
rect 6148 38668 6163 38720
rect 6189 38668 6200 38720
rect 6200 38668 6214 38720
rect 6214 38668 6245 38720
rect 6271 38668 6327 38724
rect 6353 38668 6409 38724
rect 6435 38668 6491 38724
rect 6517 38668 6573 38724
rect 6599 38668 6655 38724
rect 6681 38720 6737 38724
rect 6763 38720 6819 38724
rect 6681 38668 6702 38720
rect 6702 38668 6737 38720
rect 6763 38668 6768 38720
rect 6768 38668 6819 38720
rect 6845 38668 6901 38724
rect 6927 38668 6983 38724
rect 7009 38668 7065 38724
rect 7091 38668 7147 38724
rect 7173 38668 7229 38724
rect 7255 38720 7311 38724
rect 7337 38720 7393 38724
rect 7255 38668 7256 38720
rect 7256 38668 7308 38720
rect 7308 38668 7311 38720
rect 7337 38668 7374 38720
rect 7374 38668 7393 38720
rect 7419 38668 7475 38724
rect 7501 38668 7557 38724
rect 7583 38668 7639 38724
rect 7665 38668 7721 38724
rect 7747 38668 7803 38724
rect 7829 38720 7885 38724
rect 7911 38720 7967 38724
rect 7829 38668 7862 38720
rect 7862 38668 7876 38720
rect 7876 38668 7885 38720
rect 7911 38668 7928 38720
rect 7928 38668 7967 38720
rect 7993 38672 8047 38724
rect 8047 38672 8049 38724
rect 8075 38672 8099 38724
rect 8099 38672 8131 38724
rect 7993 38668 8049 38672
rect 8075 38668 8131 38672
rect 8157 38672 8169 38724
rect 8169 38672 8213 38724
rect 8157 38668 8213 38672
rect 5613 38599 5646 38644
rect 5646 38599 5660 38644
rect 5660 38599 5669 38644
rect 5696 38599 5712 38644
rect 5712 38599 5752 38644
rect 5613 38588 5669 38599
rect 5696 38588 5752 38599
rect 5779 38588 5835 38644
rect 5861 38588 5917 38644
rect 5943 38588 5999 38644
rect 6025 38588 6081 38644
rect 6107 38599 6148 38644
rect 6148 38599 6163 38644
rect 6189 38599 6200 38644
rect 6200 38599 6214 38644
rect 6214 38599 6245 38644
rect 6107 38588 6163 38599
rect 6189 38588 6245 38599
rect 6271 38588 6327 38644
rect 6353 38588 6409 38644
rect 6435 38588 6491 38644
rect 6517 38588 6573 38644
rect 6599 38588 6655 38644
rect 6681 38599 6702 38644
rect 6702 38599 6737 38644
rect 6763 38599 6768 38644
rect 6768 38599 6819 38644
rect 6681 38588 6737 38599
rect 6763 38588 6819 38599
rect 6845 38588 6901 38644
rect 6927 38588 6983 38644
rect 7009 38588 7065 38644
rect 7091 38588 7147 38644
rect 7173 38588 7229 38644
rect 7255 38599 7256 38644
rect 7256 38599 7308 38644
rect 7308 38599 7311 38644
rect 7337 38599 7374 38644
rect 7374 38599 7393 38644
rect 7255 38588 7311 38599
rect 7337 38588 7393 38599
rect 7419 38588 7475 38644
rect 7501 38588 7557 38644
rect 7583 38588 7639 38644
rect 7665 38588 7721 38644
rect 7747 38588 7803 38644
rect 7829 38599 7862 38644
rect 7862 38599 7876 38644
rect 7876 38599 7885 38644
rect 7911 38599 7928 38644
rect 7928 38599 7967 38644
rect 7829 38588 7885 38599
rect 7911 38588 7967 38599
rect 7993 38603 8047 38644
rect 8047 38603 8049 38644
rect 8075 38603 8099 38644
rect 8099 38603 8131 38644
rect 7993 38588 8049 38603
rect 8075 38588 8131 38603
rect 8157 38603 8169 38644
rect 8169 38603 8213 38644
rect 8157 38588 8213 38603
rect 5613 38530 5646 38564
rect 5646 38530 5660 38564
rect 5660 38530 5669 38564
rect 5696 38530 5712 38564
rect 5712 38530 5752 38564
rect 5613 38513 5669 38530
rect 5696 38513 5752 38530
rect 5613 38508 5646 38513
rect 5646 38508 5660 38513
rect 5660 38508 5669 38513
rect 5696 38508 5712 38513
rect 5712 38508 5752 38513
rect 5779 38508 5835 38564
rect 5861 38508 5917 38564
rect 5943 38508 5999 38564
rect 6025 38508 6081 38564
rect 6107 38530 6148 38564
rect 6148 38530 6163 38564
rect 6189 38530 6200 38564
rect 6200 38530 6214 38564
rect 6214 38530 6245 38564
rect 6107 38513 6163 38530
rect 6189 38513 6245 38530
rect 6107 38508 6148 38513
rect 6148 38508 6163 38513
rect 6189 38508 6200 38513
rect 6200 38508 6214 38513
rect 6214 38508 6245 38513
rect 6271 38508 6327 38564
rect 6353 38508 6409 38564
rect 6435 38508 6491 38564
rect 6517 38508 6573 38564
rect 6599 38508 6655 38564
rect 6681 38530 6702 38564
rect 6702 38530 6737 38564
rect 6763 38530 6768 38564
rect 6768 38530 6819 38564
rect 6681 38513 6737 38530
rect 6763 38513 6819 38530
rect 6681 38508 6702 38513
rect 6702 38508 6737 38513
rect 6763 38508 6768 38513
rect 6768 38508 6819 38513
rect 6845 38508 6901 38564
rect 6927 38508 6983 38564
rect 7009 38508 7065 38564
rect 7091 38508 7147 38564
rect 7173 38508 7229 38564
rect 7255 38530 7256 38564
rect 7256 38530 7308 38564
rect 7308 38530 7311 38564
rect 7337 38530 7374 38564
rect 7374 38530 7393 38564
rect 7255 38513 7311 38530
rect 7337 38513 7393 38530
rect 7255 38508 7256 38513
rect 7256 38508 7308 38513
rect 7308 38508 7311 38513
rect 7337 38508 7374 38513
rect 7374 38508 7393 38513
rect 7419 38508 7475 38564
rect 7501 38508 7557 38564
rect 7583 38508 7639 38564
rect 7665 38508 7721 38564
rect 7747 38508 7803 38564
rect 7829 38530 7862 38564
rect 7862 38530 7876 38564
rect 7876 38530 7885 38564
rect 7911 38530 7928 38564
rect 7928 38530 7967 38564
rect 7829 38513 7885 38530
rect 7911 38513 7967 38530
rect 7829 38508 7862 38513
rect 7862 38508 7876 38513
rect 7876 38508 7885 38513
rect 7911 38508 7928 38513
rect 7928 38508 7967 38513
rect 7993 38534 8047 38564
rect 8047 38534 8049 38564
rect 8075 38534 8099 38564
rect 8099 38534 8131 38564
rect 7993 38517 8049 38534
rect 8075 38517 8131 38534
rect 7993 38508 8047 38517
rect 8047 38508 8049 38517
rect 8075 38508 8099 38517
rect 8099 38508 8131 38517
rect 8157 38534 8169 38564
rect 8169 38534 8213 38564
rect 8157 38517 8213 38534
rect 8157 38508 8169 38517
rect 8169 38508 8213 38517
rect 5613 38461 5646 38484
rect 5646 38461 5660 38484
rect 5660 38461 5669 38484
rect 5696 38461 5712 38484
rect 5712 38461 5752 38484
rect 5613 38444 5669 38461
rect 5696 38444 5752 38461
rect 5613 38428 5646 38444
rect 5646 38428 5660 38444
rect 5660 38428 5669 38444
rect 5696 38428 5712 38444
rect 5712 38428 5752 38444
rect 5779 38428 5835 38484
rect 5861 38428 5917 38484
rect 5943 38428 5999 38484
rect 6025 38428 6081 38484
rect 6107 38461 6148 38484
rect 6148 38461 6163 38484
rect 6189 38461 6200 38484
rect 6200 38461 6214 38484
rect 6214 38461 6245 38484
rect 6107 38444 6163 38461
rect 6189 38444 6245 38461
rect 6107 38428 6148 38444
rect 6148 38428 6163 38444
rect 6189 38428 6200 38444
rect 6200 38428 6214 38444
rect 6214 38428 6245 38444
rect 6271 38428 6327 38484
rect 6353 38428 6409 38484
rect 6435 38428 6491 38484
rect 6517 38428 6573 38484
rect 6599 38428 6655 38484
rect 6681 38461 6702 38484
rect 6702 38461 6737 38484
rect 6763 38461 6768 38484
rect 6768 38461 6819 38484
rect 6681 38444 6737 38461
rect 6763 38444 6819 38461
rect 6681 38428 6702 38444
rect 6702 38428 6737 38444
rect 6763 38428 6768 38444
rect 6768 38428 6819 38444
rect 6845 38428 6901 38484
rect 6927 38428 6983 38484
rect 7009 38428 7065 38484
rect 7091 38428 7147 38484
rect 7173 38428 7229 38484
rect 7255 38461 7256 38484
rect 7256 38461 7308 38484
rect 7308 38461 7311 38484
rect 7337 38461 7374 38484
rect 7374 38461 7393 38484
rect 7255 38444 7311 38461
rect 7337 38444 7393 38461
rect 7255 38428 7256 38444
rect 7256 38428 7308 38444
rect 7308 38428 7311 38444
rect 7337 38428 7374 38444
rect 7374 38428 7393 38444
rect 7419 38428 7475 38484
rect 7501 38428 7557 38484
rect 7583 38428 7639 38484
rect 7665 38428 7721 38484
rect 7747 38428 7803 38484
rect 7829 38461 7862 38484
rect 7862 38461 7876 38484
rect 7876 38461 7885 38484
rect 7911 38461 7928 38484
rect 7928 38461 7967 38484
rect 7829 38444 7885 38461
rect 7911 38444 7967 38461
rect 7829 38428 7862 38444
rect 7862 38428 7876 38444
rect 7876 38428 7885 38444
rect 7911 38428 7928 38444
rect 7928 38428 7967 38444
rect 7993 38465 8047 38484
rect 8047 38465 8049 38484
rect 8075 38465 8099 38484
rect 8099 38465 8131 38484
rect 7993 38448 8049 38465
rect 8075 38448 8131 38465
rect 7993 38428 8047 38448
rect 8047 38428 8049 38448
rect 8075 38428 8099 38448
rect 8099 38428 8131 38448
rect 8157 38465 8169 38484
rect 8169 38465 8213 38484
rect 8157 38448 8213 38465
rect 8157 38428 8169 38448
rect 8169 38428 8213 38448
rect 5613 38392 5646 38404
rect 5646 38392 5660 38404
rect 5660 38392 5669 38404
rect 5696 38392 5712 38404
rect 5712 38392 5752 38404
rect 5613 38375 5669 38392
rect 5696 38375 5752 38392
rect 5613 38348 5646 38375
rect 5646 38348 5660 38375
rect 5660 38348 5669 38375
rect 5696 38348 5712 38375
rect 5712 38348 5752 38375
rect 5779 38348 5835 38404
rect 5861 38348 5917 38404
rect 5943 38348 5999 38404
rect 6025 38348 6081 38404
rect 6107 38392 6148 38404
rect 6148 38392 6163 38404
rect 6189 38392 6200 38404
rect 6200 38392 6214 38404
rect 6214 38392 6245 38404
rect 6107 38375 6163 38392
rect 6189 38375 6245 38392
rect 6107 38348 6148 38375
rect 6148 38348 6163 38375
rect 6189 38348 6200 38375
rect 6200 38348 6214 38375
rect 6214 38348 6245 38375
rect 6271 38348 6327 38404
rect 6353 38348 6409 38404
rect 6435 38348 6491 38404
rect 6517 38348 6573 38404
rect 6599 38348 6655 38404
rect 6681 38392 6702 38404
rect 6702 38392 6737 38404
rect 6763 38392 6768 38404
rect 6768 38392 6819 38404
rect 6681 38375 6737 38392
rect 6763 38375 6819 38392
rect 6681 38348 6702 38375
rect 6702 38348 6737 38375
rect 6763 38348 6768 38375
rect 6768 38348 6819 38375
rect 6845 38348 6901 38404
rect 6927 38348 6983 38404
rect 7009 38348 7065 38404
rect 7091 38348 7147 38404
rect 7173 38348 7229 38404
rect 7255 38392 7256 38404
rect 7256 38392 7308 38404
rect 7308 38392 7311 38404
rect 7337 38392 7374 38404
rect 7374 38392 7393 38404
rect 7255 38375 7311 38392
rect 7337 38375 7393 38392
rect 7255 38348 7256 38375
rect 7256 38348 7308 38375
rect 7308 38348 7311 38375
rect 7337 38348 7374 38375
rect 7374 38348 7393 38375
rect 7419 38348 7475 38404
rect 7501 38348 7557 38404
rect 7583 38348 7639 38404
rect 7665 38348 7721 38404
rect 7747 38348 7803 38404
rect 7829 38392 7862 38404
rect 7862 38392 7876 38404
rect 7876 38392 7885 38404
rect 7911 38392 7928 38404
rect 7928 38392 7967 38404
rect 7829 38375 7885 38392
rect 7911 38375 7967 38392
rect 7829 38348 7862 38375
rect 7862 38348 7876 38375
rect 7876 38348 7885 38375
rect 7911 38348 7928 38375
rect 7928 38348 7967 38375
rect 7993 38396 8047 38404
rect 8047 38396 8049 38404
rect 8075 38396 8099 38404
rect 8099 38396 8131 38404
rect 7993 38378 8049 38396
rect 8075 38378 8131 38396
rect 7993 38348 8047 38378
rect 8047 38348 8049 38378
rect 8075 38348 8099 38378
rect 8099 38348 8131 38378
rect 8157 38396 8169 38404
rect 8169 38396 8213 38404
rect 8157 38378 8213 38396
rect 8157 38348 8169 38378
rect 8169 38348 8213 38378
rect 5613 38323 5646 38324
rect 5646 38323 5660 38324
rect 5660 38323 5669 38324
rect 5696 38323 5712 38324
rect 5712 38323 5752 38324
rect 5613 38306 5669 38323
rect 5696 38306 5752 38323
rect 5613 38268 5646 38306
rect 5646 38268 5660 38306
rect 5660 38268 5669 38306
rect 5696 38268 5712 38306
rect 5712 38268 5752 38306
rect 5779 38268 5835 38324
rect 5861 38268 5917 38324
rect 5943 38268 5999 38324
rect 6025 38268 6081 38324
rect 6107 38323 6148 38324
rect 6148 38323 6163 38324
rect 6189 38323 6200 38324
rect 6200 38323 6214 38324
rect 6214 38323 6245 38324
rect 6107 38306 6163 38323
rect 6189 38306 6245 38323
rect 6107 38268 6148 38306
rect 6148 38268 6163 38306
rect 6189 38268 6200 38306
rect 6200 38268 6214 38306
rect 6214 38268 6245 38306
rect 6271 38268 6327 38324
rect 6353 38268 6409 38324
rect 6435 38268 6491 38324
rect 6517 38268 6573 38324
rect 6599 38268 6655 38324
rect 6681 38323 6702 38324
rect 6702 38323 6737 38324
rect 6763 38323 6768 38324
rect 6768 38323 6819 38324
rect 6681 38306 6737 38323
rect 6763 38306 6819 38323
rect 6681 38268 6702 38306
rect 6702 38268 6737 38306
rect 6763 38268 6768 38306
rect 6768 38268 6819 38306
rect 6845 38268 6901 38324
rect 6927 38268 6983 38324
rect 7009 38268 7065 38324
rect 7091 38268 7147 38324
rect 7173 38268 7229 38324
rect 7255 38323 7256 38324
rect 7256 38323 7308 38324
rect 7308 38323 7311 38324
rect 7337 38323 7374 38324
rect 7374 38323 7393 38324
rect 7255 38306 7311 38323
rect 7337 38306 7393 38323
rect 7255 38268 7256 38306
rect 7256 38268 7308 38306
rect 7308 38268 7311 38306
rect 7337 38268 7374 38306
rect 7374 38268 7393 38306
rect 7419 38268 7475 38324
rect 7501 38268 7557 38324
rect 7583 38268 7639 38324
rect 7665 38268 7721 38324
rect 7747 38268 7803 38324
rect 7829 38323 7862 38324
rect 7862 38323 7876 38324
rect 7876 38323 7885 38324
rect 7911 38323 7928 38324
rect 7928 38323 7967 38324
rect 7829 38306 7885 38323
rect 7911 38306 7967 38323
rect 7829 38268 7862 38306
rect 7862 38268 7876 38306
rect 7876 38268 7885 38306
rect 7911 38268 7928 38306
rect 7928 38268 7967 38306
rect 7993 38308 8049 38324
rect 8075 38308 8131 38324
rect 7993 38268 8047 38308
rect 8047 38268 8049 38308
rect 8075 38268 8099 38308
rect 8099 38268 8131 38308
rect 8157 38308 8213 38324
rect 8157 38268 8169 38308
rect 8169 38268 8213 38308
rect 5613 38236 5669 38244
rect 5696 38236 5752 38244
rect 5613 38188 5646 38236
rect 5646 38188 5660 38236
rect 5660 38188 5669 38236
rect 5696 38188 5712 38236
rect 5712 38188 5752 38236
rect 5779 38188 5835 38244
rect 5861 38188 5917 38244
rect 5943 38188 5999 38244
rect 6025 38188 6081 38244
rect 6107 38236 6163 38244
rect 6189 38236 6245 38244
rect 6107 38188 6148 38236
rect 6148 38188 6163 38236
rect 6189 38188 6200 38236
rect 6200 38188 6214 38236
rect 6214 38188 6245 38236
rect 6271 38188 6327 38244
rect 6353 38188 6409 38244
rect 6435 38188 6491 38244
rect 6517 38188 6573 38244
rect 6599 38188 6655 38244
rect 6681 38236 6737 38244
rect 6763 38236 6819 38244
rect 6681 38188 6702 38236
rect 6702 38188 6737 38236
rect 6763 38188 6768 38236
rect 6768 38188 6819 38236
rect 6845 38188 6901 38244
rect 6927 38188 6983 38244
rect 7009 38188 7065 38244
rect 7091 38188 7147 38244
rect 7173 38188 7229 38244
rect 7255 38236 7311 38244
rect 7337 38236 7393 38244
rect 7255 38188 7256 38236
rect 7256 38188 7308 38236
rect 7308 38188 7311 38236
rect 7337 38188 7374 38236
rect 7374 38188 7393 38236
rect 7419 38188 7475 38244
rect 7501 38188 7557 38244
rect 7583 38188 7639 38244
rect 7665 38188 7721 38244
rect 7747 38188 7803 38244
rect 7829 38236 7885 38244
rect 7911 38236 7967 38244
rect 7829 38188 7862 38236
rect 7862 38188 7876 38236
rect 7876 38188 7885 38236
rect 7911 38188 7928 38236
rect 7928 38188 7967 38236
rect 7993 38238 8049 38244
rect 8075 38238 8131 38244
rect 7993 38188 8047 38238
rect 8047 38188 8049 38238
rect 8075 38188 8099 38238
rect 8099 38188 8131 38238
rect 8157 38238 8213 38244
rect 8157 38188 8169 38238
rect 8169 38188 8213 38238
rect 5613 38114 5646 38164
rect 5646 38114 5660 38164
rect 5660 38114 5669 38164
rect 5696 38114 5712 38164
rect 5712 38114 5752 38164
rect 5613 38108 5669 38114
rect 5696 38108 5752 38114
rect 5779 38108 5835 38164
rect 5861 38108 5917 38164
rect 5943 38108 5999 38164
rect 6025 38108 6081 38164
rect 6107 38114 6148 38164
rect 6148 38114 6163 38164
rect 6189 38114 6200 38164
rect 6200 38114 6214 38164
rect 6214 38114 6245 38164
rect 6107 38108 6163 38114
rect 6189 38108 6245 38114
rect 6271 38108 6327 38164
rect 6353 38108 6409 38164
rect 6435 38108 6491 38164
rect 6517 38108 6573 38164
rect 6599 38108 6655 38164
rect 6681 38114 6702 38164
rect 6702 38114 6737 38164
rect 6763 38114 6768 38164
rect 6768 38114 6819 38164
rect 6681 38108 6737 38114
rect 6763 38108 6819 38114
rect 6845 38108 6901 38164
rect 6927 38108 6983 38164
rect 7009 38108 7065 38164
rect 7091 38108 7147 38164
rect 7173 38108 7229 38164
rect 7255 38114 7256 38164
rect 7256 38114 7308 38164
rect 7308 38114 7311 38164
rect 7337 38114 7374 38164
rect 7374 38114 7393 38164
rect 7255 38108 7311 38114
rect 7337 38108 7393 38114
rect 7419 38108 7475 38164
rect 7501 38108 7557 38164
rect 7583 38108 7639 38164
rect 7665 38108 7721 38164
rect 7747 38108 7803 38164
rect 7829 38114 7862 38164
rect 7862 38114 7876 38164
rect 7876 38114 7885 38164
rect 7911 38114 7928 38164
rect 7928 38114 7967 38164
rect 7829 38108 7885 38114
rect 7911 38108 7967 38114
rect 7993 38116 8047 38164
rect 8047 38116 8049 38164
rect 8075 38116 8099 38164
rect 8099 38116 8131 38164
rect 7993 38108 8049 38116
rect 8075 38108 8131 38116
rect 8157 38116 8169 38164
rect 8169 38116 8213 38164
rect 8157 38108 8213 38116
rect 2738 37931 2794 37987
rect 2819 37931 2875 37987
rect 2900 37931 2956 37987
rect 2981 37931 3037 37987
rect 3062 37982 3118 37987
rect 3143 37982 3199 37987
rect 3062 37931 3101 37982
rect 3101 37931 3118 37982
rect 3143 37931 3153 37982
rect 3153 37931 3167 37982
rect 3167 37931 3199 37982
rect 3224 37931 3280 37987
rect 3305 37931 3361 37987
rect 3386 37931 3442 37987
rect 3467 37931 3523 37987
rect 3548 37931 3604 37987
rect 3629 37982 3685 37987
rect 3710 37982 3766 37987
rect 3629 37931 3655 37982
rect 3655 37931 3685 37982
rect 3710 37931 3721 37982
rect 3721 37931 3766 37982
rect 3791 37931 3847 37987
rect 3872 37931 3928 37987
rect 3953 37931 4009 37987
rect 4034 37931 4090 37987
rect 4115 37931 4171 37987
rect 4196 37982 4252 37987
rect 4277 37982 4333 37987
rect 4196 37931 4209 37982
rect 4209 37931 4252 37982
rect 4277 37931 4327 37982
rect 4327 37931 4333 37982
rect 4358 37931 4414 37987
rect 4439 37931 4495 37987
rect 4520 37931 4576 37987
rect 4601 37931 4657 37987
rect 4682 37931 4738 37987
rect 4763 37982 5299 37987
rect 4763 37930 4815 37982
rect 4815 37930 4829 37982
rect 4829 37930 4881 37982
rect 4881 37930 5299 37982
rect 4763 37913 5299 37930
rect 2738 37851 2794 37907
rect 2819 37851 2875 37907
rect 2900 37851 2956 37907
rect 2981 37851 3037 37907
rect 3062 37861 3101 37907
rect 3101 37861 3118 37907
rect 3143 37861 3153 37907
rect 3153 37861 3167 37907
rect 3167 37861 3199 37907
rect 3062 37851 3118 37861
rect 3143 37851 3199 37861
rect 3224 37851 3280 37907
rect 3305 37851 3361 37907
rect 3386 37851 3442 37907
rect 3467 37851 3523 37907
rect 3548 37851 3604 37907
rect 3629 37861 3655 37907
rect 3655 37861 3685 37907
rect 3710 37861 3721 37907
rect 3721 37861 3766 37907
rect 3629 37851 3685 37861
rect 3710 37851 3766 37861
rect 3791 37851 3847 37907
rect 3872 37851 3928 37907
rect 3953 37851 4009 37907
rect 4034 37851 4090 37907
rect 4115 37851 4171 37907
rect 4196 37861 4209 37907
rect 4209 37861 4252 37907
rect 4277 37861 4327 37907
rect 4327 37861 4333 37907
rect 4196 37851 4252 37861
rect 4277 37851 4333 37861
rect 4358 37851 4414 37907
rect 4439 37851 4495 37907
rect 4520 37851 4576 37907
rect 4601 37851 4657 37907
rect 4682 37851 4738 37907
rect 4763 37861 4815 37913
rect 4815 37861 4829 37913
rect 4829 37861 4881 37913
rect 4881 37861 5299 37913
rect 4763 37844 5299 37861
rect 2738 37771 2794 37827
rect 2819 37771 2875 37827
rect 2900 37771 2956 37827
rect 2981 37771 3037 37827
rect 3062 37792 3101 37827
rect 3101 37792 3118 37827
rect 3143 37792 3153 37827
rect 3153 37792 3167 37827
rect 3167 37792 3199 37827
rect 3062 37775 3118 37792
rect 3143 37775 3199 37792
rect 3062 37771 3101 37775
rect 3101 37771 3118 37775
rect 3143 37771 3153 37775
rect 3153 37771 3167 37775
rect 3167 37771 3199 37775
rect 3224 37771 3280 37827
rect 3305 37771 3361 37827
rect 3386 37771 3442 37827
rect 3467 37771 3523 37827
rect 3548 37771 3604 37827
rect 3629 37792 3655 37827
rect 3655 37792 3685 37827
rect 3710 37792 3721 37827
rect 3721 37792 3766 37827
rect 3629 37775 3685 37792
rect 3710 37775 3766 37792
rect 3629 37771 3655 37775
rect 3655 37771 3685 37775
rect 3710 37771 3721 37775
rect 3721 37771 3766 37775
rect 3791 37771 3847 37827
rect 3872 37771 3928 37827
rect 3953 37771 4009 37827
rect 4034 37771 4090 37827
rect 4115 37771 4171 37827
rect 4196 37792 4209 37827
rect 4209 37792 4252 37827
rect 4277 37792 4327 37827
rect 4327 37792 4333 37827
rect 4196 37775 4252 37792
rect 4277 37775 4333 37792
rect 4196 37771 4209 37775
rect 4209 37771 4252 37775
rect 2738 37691 2794 37747
rect 2819 37691 2875 37747
rect 2900 37691 2956 37747
rect 2981 37691 3037 37747
rect 3062 37723 3101 37747
rect 3101 37723 3118 37747
rect 3143 37723 3153 37747
rect 3153 37723 3167 37747
rect 3167 37723 3199 37747
rect 3062 37706 3118 37723
rect 3143 37706 3199 37723
rect 3062 37691 3101 37706
rect 3101 37691 3118 37706
rect 3143 37691 3153 37706
rect 3153 37691 3167 37706
rect 3167 37691 3199 37706
rect 3224 37691 3280 37747
rect 3305 37691 3361 37747
rect 3386 37691 3442 37747
rect 3467 37691 3523 37747
rect 3548 37691 3604 37747
rect 3629 37723 3655 37747
rect 3655 37723 3685 37747
rect 3710 37723 3721 37747
rect 3721 37723 3766 37747
rect 3629 37706 3685 37723
rect 3710 37706 3766 37723
rect 3629 37691 3655 37706
rect 3655 37691 3685 37706
rect 3710 37691 3721 37706
rect 3721 37691 3766 37706
rect 3791 37691 3847 37747
rect 3872 37691 3928 37747
rect 3953 37691 4009 37747
rect 4034 37691 4090 37747
rect 4115 37691 4171 37747
rect 4196 37723 4209 37747
rect 4209 37723 4252 37747
rect 4277 37771 4327 37775
rect 4327 37771 4333 37775
rect 4358 37771 4414 37827
rect 4439 37771 4495 37827
rect 4520 37771 4576 37827
rect 4601 37771 4657 37827
rect 4682 37771 4738 37827
rect 4763 37792 4815 37844
rect 4815 37792 4829 37844
rect 4829 37792 4881 37844
rect 4881 37792 5299 37844
rect 4763 37775 5299 37792
rect 4277 37723 4327 37747
rect 4327 37723 4333 37747
rect 4196 37706 4252 37723
rect 4277 37706 4333 37723
rect 4196 37691 4209 37706
rect 4209 37691 4252 37706
rect 2738 37611 2794 37667
rect 2819 37611 2875 37667
rect 2900 37611 2956 37667
rect 2981 37611 3037 37667
rect 3062 37654 3101 37667
rect 3101 37654 3118 37667
rect 3143 37654 3153 37667
rect 3153 37654 3167 37667
rect 3167 37654 3199 37667
rect 3062 37636 3118 37654
rect 3143 37636 3199 37654
rect 3062 37611 3101 37636
rect 3101 37611 3118 37636
rect 3143 37611 3153 37636
rect 3153 37611 3167 37636
rect 3167 37611 3199 37636
rect 3224 37611 3280 37667
rect 3305 37611 3361 37667
rect 3386 37611 3442 37667
rect 3467 37611 3523 37667
rect 3548 37611 3604 37667
rect 3629 37654 3655 37667
rect 3655 37654 3685 37667
rect 3710 37654 3721 37667
rect 3721 37654 3766 37667
rect 3629 37636 3685 37654
rect 3710 37636 3766 37654
rect 3629 37611 3655 37636
rect 3655 37611 3685 37636
rect 3710 37611 3721 37636
rect 3721 37611 3766 37636
rect 3791 37611 3847 37667
rect 3872 37611 3928 37667
rect 3953 37611 4009 37667
rect 4034 37611 4090 37667
rect 4115 37611 4171 37667
rect 4196 37654 4209 37667
rect 4209 37654 4252 37667
rect 4277 37691 4327 37706
rect 4327 37691 4333 37706
rect 4358 37691 4414 37747
rect 4439 37691 4495 37747
rect 4520 37691 4576 37747
rect 4601 37691 4657 37747
rect 4682 37691 4738 37747
rect 4763 37723 4815 37775
rect 4815 37723 4829 37775
rect 4829 37723 4881 37775
rect 4881 37723 5299 37775
rect 4763 37706 5299 37723
rect 4277 37654 4327 37667
rect 4327 37654 4333 37667
rect 4196 37636 4252 37654
rect 4277 37636 4333 37654
rect 4196 37611 4209 37636
rect 4209 37611 4252 37636
rect 2738 37531 2794 37587
rect 2819 37531 2875 37587
rect 2900 37531 2956 37587
rect 2981 37531 3037 37587
rect 3062 37584 3101 37587
rect 3101 37584 3118 37587
rect 3143 37584 3153 37587
rect 3153 37584 3167 37587
rect 3167 37584 3199 37587
rect 3062 37566 3118 37584
rect 3143 37566 3199 37584
rect 3062 37531 3101 37566
rect 3101 37531 3118 37566
rect 3143 37531 3153 37566
rect 3153 37531 3167 37566
rect 3167 37531 3199 37566
rect 3224 37531 3280 37587
rect 3305 37531 3361 37587
rect 3386 37531 3442 37587
rect 3467 37531 3523 37587
rect 3548 37531 3604 37587
rect 3629 37584 3655 37587
rect 3655 37584 3685 37587
rect 3710 37584 3721 37587
rect 3721 37584 3766 37587
rect 3629 37566 3685 37584
rect 3710 37566 3766 37584
rect 3629 37531 3655 37566
rect 3655 37531 3685 37566
rect 3710 37531 3721 37566
rect 3721 37531 3766 37566
rect 3791 37531 3847 37587
rect 3872 37531 3928 37587
rect 3953 37531 4009 37587
rect 4034 37531 4090 37587
rect 4115 37531 4171 37587
rect 4196 37584 4209 37587
rect 4209 37584 4252 37587
rect 4277 37611 4327 37636
rect 4327 37611 4333 37636
rect 4358 37611 4414 37667
rect 4439 37611 4495 37667
rect 4520 37611 4576 37667
rect 4601 37611 4657 37667
rect 4682 37611 4738 37667
rect 4763 37654 4815 37706
rect 4815 37654 4829 37706
rect 4829 37654 4881 37706
rect 4881 37654 5299 37706
rect 4763 37636 5299 37654
rect 4277 37584 4327 37587
rect 4327 37584 4333 37587
rect 4196 37566 4252 37584
rect 4277 37566 4333 37584
rect 4196 37531 4209 37566
rect 4209 37531 4252 37566
rect 4277 37531 4327 37566
rect 4327 37531 4333 37566
rect 4358 37531 4414 37587
rect 4439 37531 4495 37587
rect 4520 37531 4576 37587
rect 4601 37531 4657 37587
rect 4682 37531 4738 37587
rect 4763 37584 4815 37636
rect 4815 37584 4829 37636
rect 4829 37584 4881 37636
rect 4881 37584 5299 37636
rect 4763 37566 5299 37584
rect 4763 37514 4815 37566
rect 4815 37514 4829 37566
rect 4829 37514 4881 37566
rect 4881 37514 5299 37566
rect 2738 37451 2794 37507
rect 2819 37451 2875 37507
rect 2900 37451 2956 37507
rect 2981 37451 3037 37507
rect 3062 37496 3118 37507
rect 3143 37496 3199 37507
rect 3062 37451 3101 37496
rect 3101 37451 3118 37496
rect 3143 37451 3153 37496
rect 3153 37451 3167 37496
rect 3167 37451 3199 37496
rect 3224 37451 3280 37507
rect 3305 37451 3361 37507
rect 3386 37451 3442 37507
rect 3467 37451 3523 37507
rect 3548 37451 3604 37507
rect 3629 37496 3685 37507
rect 3710 37496 3766 37507
rect 3629 37451 3655 37496
rect 3655 37451 3685 37496
rect 3710 37451 3721 37496
rect 3721 37451 3766 37496
rect 3791 37451 3847 37507
rect 3872 37451 3928 37507
rect 3953 37451 4009 37507
rect 4034 37451 4090 37507
rect 4115 37451 4171 37507
rect 4196 37496 4252 37507
rect 4277 37496 4333 37507
rect 4196 37451 4209 37496
rect 4209 37451 4252 37496
rect 4277 37451 4327 37496
rect 4327 37451 4333 37496
rect 4358 37451 4414 37507
rect 4439 37451 4495 37507
rect 4520 37451 4576 37507
rect 4601 37451 4657 37507
rect 4682 37451 4738 37507
rect 4763 37496 5299 37514
rect 4763 37444 4815 37496
rect 4815 37444 4829 37496
rect 4829 37444 4881 37496
rect 4881 37444 5299 37496
rect 2738 37371 2794 37427
rect 2819 37371 2875 37427
rect 2900 37371 2956 37427
rect 2981 37371 3037 37427
rect 3062 37426 3118 37427
rect 3143 37426 3199 37427
rect 3062 37374 3101 37426
rect 3101 37374 3118 37426
rect 3143 37374 3153 37426
rect 3153 37374 3167 37426
rect 3167 37374 3199 37426
rect 3062 37371 3118 37374
rect 3143 37371 3199 37374
rect 3224 37371 3280 37427
rect 3305 37371 3361 37427
rect 3386 37371 3442 37427
rect 3467 37371 3523 37427
rect 3548 37371 3604 37427
rect 3629 37426 3685 37427
rect 3710 37426 3766 37427
rect 3629 37374 3655 37426
rect 3655 37374 3685 37426
rect 3710 37374 3721 37426
rect 3721 37374 3766 37426
rect 3629 37371 3685 37374
rect 3710 37371 3766 37374
rect 3791 37371 3847 37427
rect 3872 37371 3928 37427
rect 3953 37371 4009 37427
rect 4034 37371 4090 37427
rect 4115 37371 4171 37427
rect 4196 37426 4252 37427
rect 4277 37426 4333 37427
rect 4196 37374 4209 37426
rect 4209 37374 4252 37426
rect 4277 37374 4327 37426
rect 4327 37374 4333 37426
rect 4196 37371 4252 37374
rect 4277 37371 4333 37374
rect 4358 37371 4414 37427
rect 4439 37371 4495 37427
rect 4520 37371 4576 37427
rect 4601 37371 4657 37427
rect 4682 37371 4738 37427
rect 4763 37426 5299 37444
rect 4763 37374 4815 37426
rect 4815 37374 4829 37426
rect 4829 37374 4881 37426
rect 4881 37374 5299 37426
rect 4763 37371 5299 37374
rect 5613 36720 5669 36724
rect 5696 36720 5752 36724
rect 5613 36668 5646 36720
rect 5646 36668 5660 36720
rect 5660 36668 5669 36720
rect 5696 36668 5712 36720
rect 5712 36668 5752 36720
rect 5778 36668 5834 36724
rect 5860 36668 5916 36724
rect 5942 36668 5998 36724
rect 6024 36668 6080 36724
rect 6106 36720 6162 36724
rect 6188 36720 6244 36724
rect 6106 36668 6148 36720
rect 6148 36668 6162 36720
rect 6188 36668 6200 36720
rect 6200 36668 6214 36720
rect 6214 36668 6244 36720
rect 6270 36668 6326 36724
rect 6352 36668 6408 36724
rect 6434 36668 6490 36724
rect 6516 36668 6572 36724
rect 6598 36668 6654 36724
rect 6680 36720 6736 36724
rect 6762 36720 6818 36724
rect 6680 36668 6702 36720
rect 6702 36668 6736 36720
rect 6762 36668 6768 36720
rect 6768 36668 6818 36720
rect 6844 36668 6900 36724
rect 6926 36668 6982 36724
rect 7008 36668 7064 36724
rect 7090 36668 7146 36724
rect 7172 36668 7228 36724
rect 7254 36720 7310 36724
rect 7336 36720 7392 36724
rect 7254 36668 7256 36720
rect 7256 36668 7308 36720
rect 7308 36668 7310 36720
rect 7336 36668 7374 36720
rect 7374 36668 7392 36720
rect 7418 36668 7474 36724
rect 7500 36668 7556 36724
rect 7582 36668 7638 36724
rect 7664 36668 7720 36724
rect 7746 36668 7802 36724
rect 7828 36720 7884 36724
rect 7910 36720 7966 36724
rect 7828 36668 7862 36720
rect 7862 36668 7876 36720
rect 7876 36668 7884 36720
rect 7910 36668 7928 36720
rect 7928 36668 7966 36720
rect 7992 36672 8047 36724
rect 8047 36672 8048 36724
rect 8074 36672 8099 36724
rect 8099 36672 8130 36724
rect 7992 36668 8048 36672
rect 8074 36668 8130 36672
rect 8156 36672 8169 36724
rect 8169 36672 8212 36724
rect 8156 36668 8212 36672
rect 5613 36599 5646 36644
rect 5646 36599 5660 36644
rect 5660 36599 5669 36644
rect 5696 36599 5712 36644
rect 5712 36599 5752 36644
rect 5613 36588 5669 36599
rect 5696 36588 5752 36599
rect 5778 36588 5834 36644
rect 5860 36588 5916 36644
rect 5942 36588 5998 36644
rect 6024 36588 6080 36644
rect 6106 36599 6148 36644
rect 6148 36599 6162 36644
rect 6188 36599 6200 36644
rect 6200 36599 6214 36644
rect 6214 36599 6244 36644
rect 6106 36588 6162 36599
rect 6188 36588 6244 36599
rect 6270 36588 6326 36644
rect 6352 36588 6408 36644
rect 6434 36588 6490 36644
rect 6516 36588 6572 36644
rect 6598 36588 6654 36644
rect 6680 36599 6702 36644
rect 6702 36599 6736 36644
rect 6762 36599 6768 36644
rect 6768 36599 6818 36644
rect 6680 36588 6736 36599
rect 6762 36588 6818 36599
rect 6844 36588 6900 36644
rect 6926 36588 6982 36644
rect 7008 36588 7064 36644
rect 7090 36588 7146 36644
rect 7172 36588 7228 36644
rect 7254 36599 7256 36644
rect 7256 36599 7308 36644
rect 7308 36599 7310 36644
rect 7336 36599 7374 36644
rect 7374 36599 7392 36644
rect 7254 36588 7310 36599
rect 7336 36588 7392 36599
rect 7418 36588 7474 36644
rect 7500 36588 7556 36644
rect 7582 36588 7638 36644
rect 7664 36588 7720 36644
rect 7746 36588 7802 36644
rect 7828 36599 7862 36644
rect 7862 36599 7876 36644
rect 7876 36599 7884 36644
rect 7910 36599 7928 36644
rect 7928 36599 7966 36644
rect 7828 36588 7884 36599
rect 7910 36588 7966 36599
rect 7992 36603 8047 36644
rect 8047 36603 8048 36644
rect 8074 36603 8099 36644
rect 8099 36603 8130 36644
rect 7992 36588 8048 36603
rect 8074 36588 8130 36603
rect 8156 36603 8169 36644
rect 8169 36603 8212 36644
rect 8156 36588 8212 36603
rect 5613 36530 5646 36564
rect 5646 36530 5660 36564
rect 5660 36530 5669 36564
rect 5696 36530 5712 36564
rect 5712 36530 5752 36564
rect 5613 36513 5669 36530
rect 5696 36513 5752 36530
rect 5613 36508 5646 36513
rect 5646 36508 5660 36513
rect 5660 36508 5669 36513
rect 5696 36508 5712 36513
rect 5712 36508 5752 36513
rect 5778 36508 5834 36564
rect 5860 36508 5916 36564
rect 5942 36508 5998 36564
rect 6024 36508 6080 36564
rect 6106 36530 6148 36564
rect 6148 36530 6162 36564
rect 6188 36530 6200 36564
rect 6200 36530 6214 36564
rect 6214 36530 6244 36564
rect 6106 36513 6162 36530
rect 6188 36513 6244 36530
rect 6106 36508 6148 36513
rect 6148 36508 6162 36513
rect 6188 36508 6200 36513
rect 6200 36508 6214 36513
rect 6214 36508 6244 36513
rect 6270 36508 6326 36564
rect 6352 36508 6408 36564
rect 6434 36508 6490 36564
rect 6516 36508 6572 36564
rect 6598 36508 6654 36564
rect 6680 36530 6702 36564
rect 6702 36530 6736 36564
rect 6762 36530 6768 36564
rect 6768 36530 6818 36564
rect 6680 36513 6736 36530
rect 6762 36513 6818 36530
rect 6680 36508 6702 36513
rect 6702 36508 6736 36513
rect 6762 36508 6768 36513
rect 6768 36508 6818 36513
rect 6844 36508 6900 36564
rect 6926 36508 6982 36564
rect 7008 36508 7064 36564
rect 7090 36508 7146 36564
rect 7172 36508 7228 36564
rect 7254 36530 7256 36564
rect 7256 36530 7308 36564
rect 7308 36530 7310 36564
rect 7336 36530 7374 36564
rect 7374 36530 7392 36564
rect 7254 36513 7310 36530
rect 7336 36513 7392 36530
rect 7254 36508 7256 36513
rect 7256 36508 7308 36513
rect 7308 36508 7310 36513
rect 7336 36508 7374 36513
rect 7374 36508 7392 36513
rect 7418 36508 7474 36564
rect 7500 36508 7556 36564
rect 7582 36508 7638 36564
rect 7664 36508 7720 36564
rect 7746 36508 7802 36564
rect 7828 36530 7862 36564
rect 7862 36530 7876 36564
rect 7876 36530 7884 36564
rect 7910 36530 7928 36564
rect 7928 36530 7966 36564
rect 7828 36513 7884 36530
rect 7910 36513 7966 36530
rect 7828 36508 7862 36513
rect 7862 36508 7876 36513
rect 7876 36508 7884 36513
rect 7910 36508 7928 36513
rect 7928 36508 7966 36513
rect 7992 36534 8047 36564
rect 8047 36534 8048 36564
rect 8074 36534 8099 36564
rect 8099 36534 8130 36564
rect 7992 36517 8048 36534
rect 8074 36517 8130 36534
rect 7992 36508 8047 36517
rect 8047 36508 8048 36517
rect 8074 36508 8099 36517
rect 8099 36508 8130 36517
rect 8156 36534 8169 36564
rect 8169 36534 8212 36564
rect 8156 36517 8212 36534
rect 8156 36508 8169 36517
rect 8169 36508 8212 36517
rect 5613 36461 5646 36484
rect 5646 36461 5660 36484
rect 5660 36461 5669 36484
rect 5696 36461 5712 36484
rect 5712 36461 5752 36484
rect 5613 36444 5669 36461
rect 5696 36444 5752 36461
rect 5613 36428 5646 36444
rect 5646 36428 5660 36444
rect 5660 36428 5669 36444
rect 5696 36428 5712 36444
rect 5712 36428 5752 36444
rect 5778 36428 5834 36484
rect 5860 36428 5916 36484
rect 5942 36428 5998 36484
rect 6024 36428 6080 36484
rect 6106 36461 6148 36484
rect 6148 36461 6162 36484
rect 6188 36461 6200 36484
rect 6200 36461 6214 36484
rect 6214 36461 6244 36484
rect 6106 36444 6162 36461
rect 6188 36444 6244 36461
rect 6106 36428 6148 36444
rect 6148 36428 6162 36444
rect 6188 36428 6200 36444
rect 6200 36428 6214 36444
rect 6214 36428 6244 36444
rect 6270 36428 6326 36484
rect 6352 36428 6408 36484
rect 6434 36428 6490 36484
rect 6516 36428 6572 36484
rect 6598 36428 6654 36484
rect 6680 36461 6702 36484
rect 6702 36461 6736 36484
rect 6762 36461 6768 36484
rect 6768 36461 6818 36484
rect 6680 36444 6736 36461
rect 6762 36444 6818 36461
rect 6680 36428 6702 36444
rect 6702 36428 6736 36444
rect 6762 36428 6768 36444
rect 6768 36428 6818 36444
rect 6844 36428 6900 36484
rect 6926 36428 6982 36484
rect 7008 36428 7064 36484
rect 7090 36428 7146 36484
rect 7172 36428 7228 36484
rect 7254 36461 7256 36484
rect 7256 36461 7308 36484
rect 7308 36461 7310 36484
rect 7336 36461 7374 36484
rect 7374 36461 7392 36484
rect 7254 36444 7310 36461
rect 7336 36444 7392 36461
rect 7254 36428 7256 36444
rect 7256 36428 7308 36444
rect 7308 36428 7310 36444
rect 7336 36428 7374 36444
rect 7374 36428 7392 36444
rect 7418 36428 7474 36484
rect 7500 36428 7556 36484
rect 7582 36428 7638 36484
rect 7664 36428 7720 36484
rect 7746 36428 7802 36484
rect 7828 36461 7862 36484
rect 7862 36461 7876 36484
rect 7876 36461 7884 36484
rect 7910 36461 7928 36484
rect 7928 36461 7966 36484
rect 7828 36444 7884 36461
rect 7910 36444 7966 36461
rect 7828 36428 7862 36444
rect 7862 36428 7876 36444
rect 7876 36428 7884 36444
rect 7910 36428 7928 36444
rect 7928 36428 7966 36444
rect 7992 36465 8047 36484
rect 8047 36465 8048 36484
rect 8074 36465 8099 36484
rect 8099 36465 8130 36484
rect 7992 36448 8048 36465
rect 8074 36448 8130 36465
rect 7992 36428 8047 36448
rect 8047 36428 8048 36448
rect 8074 36428 8099 36448
rect 8099 36428 8130 36448
rect 8156 36465 8169 36484
rect 8169 36465 8212 36484
rect 8156 36448 8212 36465
rect 8156 36428 8169 36448
rect 8169 36428 8212 36448
rect 5613 36392 5646 36404
rect 5646 36392 5660 36404
rect 5660 36392 5669 36404
rect 5696 36392 5712 36404
rect 5712 36392 5752 36404
rect 5613 36375 5669 36392
rect 5696 36375 5752 36392
rect 5613 36348 5646 36375
rect 5646 36348 5660 36375
rect 5660 36348 5669 36375
rect 5696 36348 5712 36375
rect 5712 36348 5752 36375
rect 5778 36348 5834 36404
rect 5860 36348 5916 36404
rect 5942 36348 5998 36404
rect 6024 36348 6080 36404
rect 6106 36392 6148 36404
rect 6148 36392 6162 36404
rect 6188 36392 6200 36404
rect 6200 36392 6214 36404
rect 6214 36392 6244 36404
rect 6106 36375 6162 36392
rect 6188 36375 6244 36392
rect 6106 36348 6148 36375
rect 6148 36348 6162 36375
rect 6188 36348 6200 36375
rect 6200 36348 6214 36375
rect 6214 36348 6244 36375
rect 6270 36348 6326 36404
rect 6352 36348 6408 36404
rect 6434 36348 6490 36404
rect 6516 36348 6572 36404
rect 6598 36348 6654 36404
rect 6680 36392 6702 36404
rect 6702 36392 6736 36404
rect 6762 36392 6768 36404
rect 6768 36392 6818 36404
rect 6680 36375 6736 36392
rect 6762 36375 6818 36392
rect 6680 36348 6702 36375
rect 6702 36348 6736 36375
rect 6762 36348 6768 36375
rect 6768 36348 6818 36375
rect 6844 36348 6900 36404
rect 6926 36348 6982 36404
rect 7008 36348 7064 36404
rect 7090 36348 7146 36404
rect 7172 36348 7228 36404
rect 7254 36392 7256 36404
rect 7256 36392 7308 36404
rect 7308 36392 7310 36404
rect 7336 36392 7374 36404
rect 7374 36392 7392 36404
rect 7254 36375 7310 36392
rect 7336 36375 7392 36392
rect 7254 36348 7256 36375
rect 7256 36348 7308 36375
rect 7308 36348 7310 36375
rect 7336 36348 7374 36375
rect 7374 36348 7392 36375
rect 7418 36348 7474 36404
rect 7500 36348 7556 36404
rect 7582 36348 7638 36404
rect 7664 36348 7720 36404
rect 7746 36348 7802 36404
rect 7828 36392 7862 36404
rect 7862 36392 7876 36404
rect 7876 36392 7884 36404
rect 7910 36392 7928 36404
rect 7928 36392 7966 36404
rect 7828 36375 7884 36392
rect 7910 36375 7966 36392
rect 7828 36348 7862 36375
rect 7862 36348 7876 36375
rect 7876 36348 7884 36375
rect 7910 36348 7928 36375
rect 7928 36348 7966 36375
rect 7992 36396 8047 36404
rect 8047 36396 8048 36404
rect 8074 36396 8099 36404
rect 8099 36396 8130 36404
rect 7992 36378 8048 36396
rect 8074 36378 8130 36396
rect 7992 36348 8047 36378
rect 8047 36348 8048 36378
rect 8074 36348 8099 36378
rect 8099 36348 8130 36378
rect 8156 36396 8169 36404
rect 8169 36396 8212 36404
rect 8156 36378 8212 36396
rect 8156 36348 8169 36378
rect 8169 36348 8212 36378
rect 5613 36323 5646 36324
rect 5646 36323 5660 36324
rect 5660 36323 5669 36324
rect 5696 36323 5712 36324
rect 5712 36323 5752 36324
rect 5613 36306 5669 36323
rect 5696 36306 5752 36323
rect 5613 36268 5646 36306
rect 5646 36268 5660 36306
rect 5660 36268 5669 36306
rect 5696 36268 5712 36306
rect 5712 36268 5752 36306
rect 5778 36268 5834 36324
rect 5860 36268 5916 36324
rect 5942 36268 5998 36324
rect 6024 36268 6080 36324
rect 6106 36323 6148 36324
rect 6148 36323 6162 36324
rect 6188 36323 6200 36324
rect 6200 36323 6214 36324
rect 6214 36323 6244 36324
rect 6106 36306 6162 36323
rect 6188 36306 6244 36323
rect 6106 36268 6148 36306
rect 6148 36268 6162 36306
rect 6188 36268 6200 36306
rect 6200 36268 6214 36306
rect 6214 36268 6244 36306
rect 6270 36268 6326 36324
rect 6352 36268 6408 36324
rect 6434 36268 6490 36324
rect 6516 36268 6572 36324
rect 6598 36268 6654 36324
rect 6680 36323 6702 36324
rect 6702 36323 6736 36324
rect 6762 36323 6768 36324
rect 6768 36323 6818 36324
rect 6680 36306 6736 36323
rect 6762 36306 6818 36323
rect 6680 36268 6702 36306
rect 6702 36268 6736 36306
rect 6762 36268 6768 36306
rect 6768 36268 6818 36306
rect 6844 36268 6900 36324
rect 6926 36268 6982 36324
rect 7008 36268 7064 36324
rect 7090 36268 7146 36324
rect 7172 36268 7228 36324
rect 7254 36323 7256 36324
rect 7256 36323 7308 36324
rect 7308 36323 7310 36324
rect 7336 36323 7374 36324
rect 7374 36323 7392 36324
rect 7254 36306 7310 36323
rect 7336 36306 7392 36323
rect 7254 36268 7256 36306
rect 7256 36268 7308 36306
rect 7308 36268 7310 36306
rect 7336 36268 7374 36306
rect 7374 36268 7392 36306
rect 7418 36268 7474 36324
rect 7500 36268 7556 36324
rect 7582 36268 7638 36324
rect 7664 36268 7720 36324
rect 7746 36268 7802 36324
rect 7828 36323 7862 36324
rect 7862 36323 7876 36324
rect 7876 36323 7884 36324
rect 7910 36323 7928 36324
rect 7928 36323 7966 36324
rect 7828 36306 7884 36323
rect 7910 36306 7966 36323
rect 7828 36268 7862 36306
rect 7862 36268 7876 36306
rect 7876 36268 7884 36306
rect 7910 36268 7928 36306
rect 7928 36268 7966 36306
rect 7992 36308 8048 36324
rect 8074 36308 8130 36324
rect 7992 36268 8047 36308
rect 8047 36268 8048 36308
rect 8074 36268 8099 36308
rect 8099 36268 8130 36308
rect 8156 36308 8212 36324
rect 8156 36268 8169 36308
rect 8169 36268 8212 36308
rect 5613 36236 5669 36244
rect 5696 36236 5752 36244
rect 5613 36188 5646 36236
rect 5646 36188 5660 36236
rect 5660 36188 5669 36236
rect 5696 36188 5712 36236
rect 5712 36188 5752 36236
rect 5778 36188 5834 36244
rect 5860 36188 5916 36244
rect 5942 36188 5998 36244
rect 6024 36188 6080 36244
rect 6106 36236 6162 36244
rect 6188 36236 6244 36244
rect 6106 36188 6148 36236
rect 6148 36188 6162 36236
rect 6188 36188 6200 36236
rect 6200 36188 6214 36236
rect 6214 36188 6244 36236
rect 6270 36188 6326 36244
rect 6352 36188 6408 36244
rect 6434 36188 6490 36244
rect 6516 36188 6572 36244
rect 6598 36188 6654 36244
rect 6680 36236 6736 36244
rect 6762 36236 6818 36244
rect 6680 36188 6702 36236
rect 6702 36188 6736 36236
rect 6762 36188 6768 36236
rect 6768 36188 6818 36236
rect 6844 36188 6900 36244
rect 6926 36188 6982 36244
rect 7008 36188 7064 36244
rect 7090 36188 7146 36244
rect 7172 36188 7228 36244
rect 7254 36236 7310 36244
rect 7336 36236 7392 36244
rect 7254 36188 7256 36236
rect 7256 36188 7308 36236
rect 7308 36188 7310 36236
rect 7336 36188 7374 36236
rect 7374 36188 7392 36236
rect 7418 36188 7474 36244
rect 7500 36188 7556 36244
rect 7582 36188 7638 36244
rect 7664 36188 7720 36244
rect 7746 36188 7802 36244
rect 7828 36236 7884 36244
rect 7910 36236 7966 36244
rect 7828 36188 7862 36236
rect 7862 36188 7876 36236
rect 7876 36188 7884 36236
rect 7910 36188 7928 36236
rect 7928 36188 7966 36236
rect 7992 36238 8048 36244
rect 8074 36238 8130 36244
rect 7992 36188 8047 36238
rect 8047 36188 8048 36238
rect 8074 36188 8099 36238
rect 8099 36188 8130 36238
rect 8156 36238 8212 36244
rect 8156 36188 8169 36238
rect 8169 36188 8212 36238
rect 5613 36114 5646 36164
rect 5646 36114 5660 36164
rect 5660 36114 5669 36164
rect 5696 36114 5712 36164
rect 5712 36114 5752 36164
rect 5613 36108 5669 36114
rect 5696 36108 5752 36114
rect 5778 36108 5834 36164
rect 5860 36108 5916 36164
rect 5942 36108 5998 36164
rect 6024 36108 6080 36164
rect 6106 36114 6148 36164
rect 6148 36114 6162 36164
rect 6188 36114 6200 36164
rect 6200 36114 6214 36164
rect 6214 36114 6244 36164
rect 6106 36108 6162 36114
rect 6188 36108 6244 36114
rect 6270 36108 6326 36164
rect 6352 36108 6408 36164
rect 6434 36108 6490 36164
rect 6516 36108 6572 36164
rect 6598 36108 6654 36164
rect 6680 36114 6702 36164
rect 6702 36114 6736 36164
rect 6762 36114 6768 36164
rect 6768 36114 6818 36164
rect 6680 36108 6736 36114
rect 6762 36108 6818 36114
rect 6844 36108 6900 36164
rect 6926 36108 6982 36164
rect 7008 36108 7064 36164
rect 7090 36108 7146 36164
rect 7172 36108 7228 36164
rect 7254 36114 7256 36164
rect 7256 36114 7308 36164
rect 7308 36114 7310 36164
rect 7336 36114 7374 36164
rect 7374 36114 7392 36164
rect 7254 36108 7310 36114
rect 7336 36108 7392 36114
rect 7418 36108 7474 36164
rect 7500 36108 7556 36164
rect 7582 36108 7638 36164
rect 7664 36108 7720 36164
rect 7746 36108 7802 36164
rect 7828 36114 7862 36164
rect 7862 36114 7876 36164
rect 7876 36114 7884 36164
rect 7910 36114 7928 36164
rect 7928 36114 7966 36164
rect 7828 36108 7884 36114
rect 7910 36108 7966 36114
rect 7992 36116 8047 36164
rect 8047 36116 8048 36164
rect 8074 36116 8099 36164
rect 8099 36116 8130 36164
rect 7992 36108 8048 36116
rect 8074 36108 8130 36116
rect 8156 36116 8169 36164
rect 8169 36116 8212 36164
rect 8156 36108 8212 36116
rect 2733 35931 2789 35987
rect 2814 35931 2870 35987
rect 2895 35931 2951 35987
rect 2976 35931 3032 35987
rect 3057 35982 3113 35987
rect 3138 35982 3194 35987
rect 3057 35931 3101 35982
rect 3101 35931 3113 35982
rect 3138 35931 3153 35982
rect 3153 35931 3167 35982
rect 3167 35931 3194 35982
rect 3219 35931 3275 35987
rect 3300 35931 3356 35987
rect 3381 35931 3437 35987
rect 3462 35931 3518 35987
rect 3543 35931 3599 35987
rect 3624 35982 3680 35987
rect 3705 35982 3761 35987
rect 3624 35931 3655 35982
rect 3655 35931 3680 35982
rect 3705 35931 3707 35982
rect 3707 35931 3721 35982
rect 3721 35931 3761 35982
rect 3786 35931 3842 35987
rect 3867 35931 3923 35987
rect 3948 35931 4004 35987
rect 4029 35931 4085 35987
rect 4110 35931 4166 35987
rect 4191 35982 4247 35987
rect 4272 35982 4328 35987
rect 4191 35931 4209 35982
rect 4209 35931 4247 35982
rect 4272 35931 4275 35982
rect 4275 35931 4327 35982
rect 4327 35931 4328 35982
rect 4353 35931 4409 35987
rect 4434 35931 4490 35987
rect 4515 35931 4571 35987
rect 4596 35931 4652 35987
rect 4677 35931 4733 35987
rect 4758 35982 4814 35987
rect 4839 35982 4895 35987
rect 4758 35931 4763 35982
rect 4763 35931 4814 35982
rect 4839 35931 4881 35982
rect 4881 35931 4895 35982
rect 4920 35931 4976 35987
rect 5001 35931 5057 35987
rect 5082 35931 5138 35987
rect 2733 35851 2789 35907
rect 2814 35851 2870 35907
rect 2895 35851 2951 35907
rect 2976 35851 3032 35907
rect 3057 35861 3101 35907
rect 3101 35861 3113 35907
rect 3138 35861 3153 35907
rect 3153 35861 3167 35907
rect 3167 35861 3194 35907
rect 3057 35851 3113 35861
rect 3138 35851 3194 35861
rect 3219 35851 3275 35907
rect 3300 35851 3356 35907
rect 3381 35851 3437 35907
rect 3462 35851 3518 35907
rect 3543 35851 3599 35907
rect 3624 35861 3655 35907
rect 3655 35861 3680 35907
rect 3705 35861 3707 35907
rect 3707 35861 3721 35907
rect 3721 35861 3761 35907
rect 3624 35851 3680 35861
rect 3705 35851 3761 35861
rect 3786 35851 3842 35907
rect 3867 35851 3923 35907
rect 3948 35851 4004 35907
rect 4029 35851 4085 35907
rect 4110 35851 4166 35907
rect 4191 35861 4209 35907
rect 4209 35861 4247 35907
rect 4272 35861 4275 35907
rect 4275 35861 4327 35907
rect 4327 35861 4328 35907
rect 4191 35851 4247 35861
rect 4272 35851 4328 35861
rect 4353 35851 4409 35907
rect 4434 35851 4490 35907
rect 4515 35851 4571 35907
rect 4596 35851 4652 35907
rect 4677 35851 4733 35907
rect 4758 35861 4763 35907
rect 4763 35861 4814 35907
rect 4839 35861 4881 35907
rect 4881 35861 4895 35907
rect 4758 35851 4814 35861
rect 4839 35851 4895 35861
rect 4920 35851 4976 35907
rect 5001 35851 5057 35907
rect 5082 35851 5138 35907
rect 2733 35771 2789 35827
rect 2814 35771 2870 35827
rect 2895 35771 2951 35827
rect 2976 35771 3032 35827
rect 3057 35792 3101 35827
rect 3101 35792 3113 35827
rect 3138 35792 3153 35827
rect 3153 35792 3167 35827
rect 3167 35792 3194 35827
rect 3057 35775 3113 35792
rect 3138 35775 3194 35792
rect 3057 35771 3101 35775
rect 3101 35771 3113 35775
rect 3138 35771 3153 35775
rect 3153 35771 3167 35775
rect 3167 35771 3194 35775
rect 3219 35771 3275 35827
rect 3300 35771 3356 35827
rect 3381 35771 3437 35827
rect 3462 35771 3518 35827
rect 3543 35771 3599 35827
rect 3624 35792 3655 35827
rect 3655 35792 3680 35827
rect 3705 35792 3707 35827
rect 3707 35792 3721 35827
rect 3721 35792 3761 35827
rect 3624 35775 3680 35792
rect 3705 35775 3761 35792
rect 3624 35771 3655 35775
rect 3655 35771 3680 35775
rect 3705 35771 3707 35775
rect 3707 35771 3721 35775
rect 3721 35771 3761 35775
rect 3786 35771 3842 35827
rect 3867 35771 3923 35827
rect 3948 35771 4004 35827
rect 4029 35771 4085 35827
rect 4110 35771 4166 35827
rect 4191 35792 4209 35827
rect 4209 35792 4247 35827
rect 4272 35792 4275 35827
rect 4275 35792 4327 35827
rect 4327 35792 4328 35827
rect 4191 35775 4247 35792
rect 4272 35775 4328 35792
rect 4191 35771 4209 35775
rect 4209 35771 4247 35775
rect 4272 35771 4275 35775
rect 4275 35771 4327 35775
rect 4327 35771 4328 35775
rect 4353 35771 4409 35827
rect 4434 35771 4490 35827
rect 4515 35771 4571 35827
rect 4596 35771 4652 35827
rect 4677 35771 4733 35827
rect 4758 35792 4763 35827
rect 4763 35792 4814 35827
rect 4839 35792 4881 35827
rect 4881 35792 4895 35827
rect 4758 35775 4814 35792
rect 4839 35775 4895 35792
rect 4758 35771 4763 35775
rect 4763 35771 4814 35775
rect 2733 35691 2789 35747
rect 2814 35691 2870 35747
rect 2895 35691 2951 35747
rect 2976 35691 3032 35747
rect 3057 35723 3101 35747
rect 3101 35723 3113 35747
rect 3138 35723 3153 35747
rect 3153 35723 3167 35747
rect 3167 35723 3194 35747
rect 3057 35706 3113 35723
rect 3138 35706 3194 35723
rect 3057 35691 3101 35706
rect 3101 35691 3113 35706
rect 3138 35691 3153 35706
rect 3153 35691 3167 35706
rect 3167 35691 3194 35706
rect 3219 35691 3275 35747
rect 3300 35691 3356 35747
rect 3381 35691 3437 35747
rect 3462 35691 3518 35747
rect 3543 35691 3599 35747
rect 3624 35723 3655 35747
rect 3655 35723 3680 35747
rect 3705 35723 3707 35747
rect 3707 35723 3721 35747
rect 3721 35723 3761 35747
rect 3624 35706 3680 35723
rect 3705 35706 3761 35723
rect 3624 35691 3655 35706
rect 3655 35691 3680 35706
rect 3705 35691 3707 35706
rect 3707 35691 3721 35706
rect 3721 35691 3761 35706
rect 3786 35691 3842 35747
rect 3867 35691 3923 35747
rect 3948 35691 4004 35747
rect 4029 35691 4085 35747
rect 4110 35691 4166 35747
rect 4191 35723 4209 35747
rect 4209 35723 4247 35747
rect 4272 35723 4275 35747
rect 4275 35723 4327 35747
rect 4327 35723 4328 35747
rect 4191 35706 4247 35723
rect 4272 35706 4328 35723
rect 4191 35691 4209 35706
rect 4209 35691 4247 35706
rect 4272 35691 4275 35706
rect 4275 35691 4327 35706
rect 4327 35691 4328 35706
rect 4353 35691 4409 35747
rect 4434 35691 4490 35747
rect 4515 35691 4571 35747
rect 4596 35691 4652 35747
rect 4677 35691 4733 35747
rect 4758 35723 4763 35747
rect 4763 35723 4814 35747
rect 4839 35771 4881 35775
rect 4881 35771 4895 35775
rect 4920 35771 4976 35827
rect 5001 35771 5057 35827
rect 5082 35771 5138 35827
rect 4839 35723 4881 35747
rect 4881 35723 4895 35747
rect 4758 35706 4814 35723
rect 4839 35706 4895 35723
rect 4758 35691 4763 35706
rect 4763 35691 4814 35706
rect 2733 35611 2789 35667
rect 2814 35611 2870 35667
rect 2895 35611 2951 35667
rect 2976 35611 3032 35667
rect 3057 35654 3101 35667
rect 3101 35654 3113 35667
rect 3138 35654 3153 35667
rect 3153 35654 3167 35667
rect 3167 35654 3194 35667
rect 3057 35636 3113 35654
rect 3138 35636 3194 35654
rect 3057 35611 3101 35636
rect 3101 35611 3113 35636
rect 3138 35611 3153 35636
rect 3153 35611 3167 35636
rect 3167 35611 3194 35636
rect 3219 35611 3275 35667
rect 3300 35611 3356 35667
rect 3381 35611 3437 35667
rect 3462 35611 3518 35667
rect 3543 35611 3599 35667
rect 3624 35654 3655 35667
rect 3655 35654 3680 35667
rect 3705 35654 3707 35667
rect 3707 35654 3721 35667
rect 3721 35654 3761 35667
rect 3624 35636 3680 35654
rect 3705 35636 3761 35654
rect 3624 35611 3655 35636
rect 3655 35611 3680 35636
rect 3705 35611 3707 35636
rect 3707 35611 3721 35636
rect 3721 35611 3761 35636
rect 3786 35611 3842 35667
rect 3867 35611 3923 35667
rect 3948 35611 4004 35667
rect 4029 35611 4085 35667
rect 4110 35611 4166 35667
rect 4191 35654 4209 35667
rect 4209 35654 4247 35667
rect 4272 35654 4275 35667
rect 4275 35654 4327 35667
rect 4327 35654 4328 35667
rect 4191 35636 4247 35654
rect 4272 35636 4328 35654
rect 4191 35611 4209 35636
rect 4209 35611 4247 35636
rect 4272 35611 4275 35636
rect 4275 35611 4327 35636
rect 4327 35611 4328 35636
rect 4353 35611 4409 35667
rect 4434 35611 4490 35667
rect 4515 35611 4571 35667
rect 4596 35611 4652 35667
rect 4677 35611 4733 35667
rect 4758 35654 4763 35667
rect 4763 35654 4814 35667
rect 4839 35691 4881 35706
rect 4881 35691 4895 35706
rect 4920 35691 4976 35747
rect 5001 35691 5057 35747
rect 5082 35691 5138 35747
rect 4839 35654 4881 35667
rect 4881 35654 4895 35667
rect 4758 35636 4814 35654
rect 4839 35636 4895 35654
rect 4758 35611 4763 35636
rect 4763 35611 4814 35636
rect 2733 35531 2789 35587
rect 2814 35531 2870 35587
rect 2895 35531 2951 35587
rect 2976 35531 3032 35587
rect 3057 35584 3101 35587
rect 3101 35584 3113 35587
rect 3138 35584 3153 35587
rect 3153 35584 3167 35587
rect 3167 35584 3194 35587
rect 3057 35566 3113 35584
rect 3138 35566 3194 35584
rect 3057 35531 3101 35566
rect 3101 35531 3113 35566
rect 3138 35531 3153 35566
rect 3153 35531 3167 35566
rect 3167 35531 3194 35566
rect 3219 35531 3275 35587
rect 3300 35531 3356 35587
rect 3381 35531 3437 35587
rect 3462 35531 3518 35587
rect 3543 35531 3599 35587
rect 3624 35584 3655 35587
rect 3655 35584 3680 35587
rect 3705 35584 3707 35587
rect 3707 35584 3721 35587
rect 3721 35584 3761 35587
rect 3624 35566 3680 35584
rect 3705 35566 3761 35584
rect 3624 35531 3655 35566
rect 3655 35531 3680 35566
rect 3705 35531 3707 35566
rect 3707 35531 3721 35566
rect 3721 35531 3761 35566
rect 3786 35531 3842 35587
rect 3867 35531 3923 35587
rect 3948 35531 4004 35587
rect 4029 35531 4085 35587
rect 4110 35531 4166 35587
rect 4191 35584 4209 35587
rect 4209 35584 4247 35587
rect 4272 35584 4275 35587
rect 4275 35584 4327 35587
rect 4327 35584 4328 35587
rect 4191 35566 4247 35584
rect 4272 35566 4328 35584
rect 4191 35531 4209 35566
rect 4209 35531 4247 35566
rect 4272 35531 4275 35566
rect 4275 35531 4327 35566
rect 4327 35531 4328 35566
rect 4353 35531 4409 35587
rect 4434 35531 4490 35587
rect 4515 35531 4571 35587
rect 4596 35531 4652 35587
rect 4677 35531 4733 35587
rect 4758 35584 4763 35587
rect 4763 35584 4814 35587
rect 4839 35611 4881 35636
rect 4881 35611 4895 35636
rect 4920 35611 4976 35667
rect 5001 35611 5057 35667
rect 5082 35611 5138 35667
rect 4839 35584 4881 35587
rect 4881 35584 4895 35587
rect 4758 35566 4814 35584
rect 4839 35566 4895 35584
rect 4758 35531 4763 35566
rect 4763 35531 4814 35566
rect 4839 35531 4881 35566
rect 4881 35531 4895 35566
rect 4920 35531 4976 35587
rect 5001 35531 5057 35587
rect 5082 35531 5138 35587
rect 2733 35451 2789 35507
rect 2814 35451 2870 35507
rect 2895 35451 2951 35507
rect 2976 35451 3032 35507
rect 3057 35496 3113 35507
rect 3138 35496 3194 35507
rect 3057 35451 3101 35496
rect 3101 35451 3113 35496
rect 3138 35451 3153 35496
rect 3153 35451 3167 35496
rect 3167 35451 3194 35496
rect 3219 35451 3275 35507
rect 3300 35451 3356 35507
rect 3381 35451 3437 35507
rect 3462 35451 3518 35507
rect 3543 35451 3599 35507
rect 3624 35496 3680 35507
rect 3705 35496 3761 35507
rect 3624 35451 3655 35496
rect 3655 35451 3680 35496
rect 3705 35451 3707 35496
rect 3707 35451 3721 35496
rect 3721 35451 3761 35496
rect 3786 35451 3842 35507
rect 3867 35451 3923 35507
rect 3948 35451 4004 35507
rect 4029 35451 4085 35507
rect 4110 35451 4166 35507
rect 4191 35496 4247 35507
rect 4272 35496 4328 35507
rect 4191 35451 4209 35496
rect 4209 35451 4247 35496
rect 4272 35451 4275 35496
rect 4275 35451 4327 35496
rect 4327 35451 4328 35496
rect 4353 35451 4409 35507
rect 4434 35451 4490 35507
rect 4515 35451 4571 35507
rect 4596 35451 4652 35507
rect 4677 35451 4733 35507
rect 4758 35496 4814 35507
rect 4839 35496 4895 35507
rect 4758 35451 4763 35496
rect 4763 35451 4814 35496
rect 4839 35451 4881 35496
rect 4881 35451 4895 35496
rect 4920 35451 4976 35507
rect 5001 35451 5057 35507
rect 5082 35451 5138 35507
rect 2733 35371 2789 35427
rect 2814 35371 2870 35427
rect 2895 35371 2951 35427
rect 2976 35371 3032 35427
rect 3057 35426 3113 35427
rect 3138 35426 3194 35427
rect 3057 35374 3101 35426
rect 3101 35374 3113 35426
rect 3138 35374 3153 35426
rect 3153 35374 3167 35426
rect 3167 35374 3194 35426
rect 3057 35371 3113 35374
rect 3138 35371 3194 35374
rect 3219 35371 3275 35427
rect 3300 35371 3356 35427
rect 3381 35371 3437 35427
rect 3462 35371 3518 35427
rect 3543 35371 3599 35427
rect 3624 35426 3680 35427
rect 3705 35426 3761 35427
rect 3624 35374 3655 35426
rect 3655 35374 3680 35426
rect 3705 35374 3707 35426
rect 3707 35374 3721 35426
rect 3721 35374 3761 35426
rect 3624 35371 3680 35374
rect 3705 35371 3761 35374
rect 3786 35371 3842 35427
rect 3867 35371 3923 35427
rect 3948 35371 4004 35427
rect 4029 35371 4085 35427
rect 4110 35371 4166 35427
rect 4191 35426 4247 35427
rect 4272 35426 4328 35427
rect 4191 35374 4209 35426
rect 4209 35374 4247 35426
rect 4272 35374 4275 35426
rect 4275 35374 4327 35426
rect 4327 35374 4328 35426
rect 4191 35371 4247 35374
rect 4272 35371 4328 35374
rect 4353 35371 4409 35427
rect 4434 35371 4490 35427
rect 4515 35371 4571 35427
rect 4596 35371 4652 35427
rect 4677 35371 4733 35427
rect 4758 35426 4814 35427
rect 4839 35426 4895 35427
rect 4758 35374 4763 35426
rect 4763 35374 4814 35426
rect 4839 35374 4881 35426
rect 4881 35374 4895 35426
rect 4758 35371 4814 35374
rect 4839 35371 4895 35374
rect 4920 35371 4976 35427
rect 5001 35371 5057 35427
rect 5082 35371 5138 35427
rect 5163 35371 5299 35987
rect 5613 34720 5669 34724
rect 5696 34720 5752 34724
rect 5613 34668 5646 34720
rect 5646 34668 5660 34720
rect 5660 34668 5669 34720
rect 5696 34668 5712 34720
rect 5712 34668 5752 34720
rect 5779 34668 5835 34724
rect 5861 34668 5917 34724
rect 5943 34668 5999 34724
rect 6025 34668 6081 34724
rect 6107 34720 6163 34724
rect 6189 34720 6245 34724
rect 6107 34668 6148 34720
rect 6148 34668 6163 34720
rect 6189 34668 6200 34720
rect 6200 34668 6214 34720
rect 6214 34668 6245 34720
rect 6271 34668 6327 34724
rect 6353 34668 6409 34724
rect 6435 34668 6491 34724
rect 6517 34668 6573 34724
rect 6599 34668 6655 34724
rect 6681 34720 6737 34724
rect 6763 34720 6819 34724
rect 6681 34668 6702 34720
rect 6702 34668 6737 34720
rect 6763 34668 6768 34720
rect 6768 34668 6819 34720
rect 6845 34668 6901 34724
rect 6927 34668 6983 34724
rect 7009 34668 7065 34724
rect 7091 34668 7147 34724
rect 7173 34668 7229 34724
rect 7255 34720 7311 34724
rect 7337 34720 7393 34724
rect 7255 34668 7256 34720
rect 7256 34668 7308 34720
rect 7308 34668 7311 34720
rect 7337 34668 7374 34720
rect 7374 34668 7393 34720
rect 7419 34668 7475 34724
rect 7501 34668 7557 34724
rect 7583 34668 7639 34724
rect 7665 34668 7721 34724
rect 7747 34668 7803 34724
rect 7829 34720 7885 34724
rect 7911 34720 7967 34724
rect 7829 34668 7862 34720
rect 7862 34668 7876 34720
rect 7876 34668 7885 34720
rect 7911 34668 7928 34720
rect 7928 34668 7967 34720
rect 7993 34672 8047 34724
rect 8047 34672 8049 34724
rect 8075 34672 8099 34724
rect 8099 34672 8131 34724
rect 7993 34668 8049 34672
rect 8075 34668 8131 34672
rect 8157 34672 8169 34724
rect 8169 34672 8213 34724
rect 8157 34668 8213 34672
rect 5613 34599 5646 34644
rect 5646 34599 5660 34644
rect 5660 34599 5669 34644
rect 5696 34599 5712 34644
rect 5712 34599 5752 34644
rect 5613 34588 5669 34599
rect 5696 34588 5752 34599
rect 5779 34588 5835 34644
rect 5861 34588 5917 34644
rect 5943 34588 5999 34644
rect 6025 34588 6081 34644
rect 6107 34599 6148 34644
rect 6148 34599 6163 34644
rect 6189 34599 6200 34644
rect 6200 34599 6214 34644
rect 6214 34599 6245 34644
rect 6107 34588 6163 34599
rect 6189 34588 6245 34599
rect 6271 34588 6327 34644
rect 6353 34588 6409 34644
rect 6435 34588 6491 34644
rect 6517 34588 6573 34644
rect 6599 34588 6655 34644
rect 6681 34599 6702 34644
rect 6702 34599 6737 34644
rect 6763 34599 6768 34644
rect 6768 34599 6819 34644
rect 6681 34588 6737 34599
rect 6763 34588 6819 34599
rect 6845 34588 6901 34644
rect 6927 34588 6983 34644
rect 7009 34588 7065 34644
rect 7091 34588 7147 34644
rect 7173 34588 7229 34644
rect 7255 34599 7256 34644
rect 7256 34599 7308 34644
rect 7308 34599 7311 34644
rect 7337 34599 7374 34644
rect 7374 34599 7393 34644
rect 7255 34588 7311 34599
rect 7337 34588 7393 34599
rect 7419 34588 7475 34644
rect 7501 34588 7557 34644
rect 7583 34588 7639 34644
rect 7665 34588 7721 34644
rect 7747 34588 7803 34644
rect 7829 34599 7862 34644
rect 7862 34599 7876 34644
rect 7876 34599 7885 34644
rect 7911 34599 7928 34644
rect 7928 34599 7967 34644
rect 7829 34588 7885 34599
rect 7911 34588 7967 34599
rect 7993 34603 8047 34644
rect 8047 34603 8049 34644
rect 8075 34603 8099 34644
rect 8099 34603 8131 34644
rect 7993 34588 8049 34603
rect 8075 34588 8131 34603
rect 8157 34603 8169 34644
rect 8169 34603 8213 34644
rect 8157 34588 8213 34603
rect 5613 34530 5646 34564
rect 5646 34530 5660 34564
rect 5660 34530 5669 34564
rect 5696 34530 5712 34564
rect 5712 34530 5752 34564
rect 5613 34513 5669 34530
rect 5696 34513 5752 34530
rect 5613 34508 5646 34513
rect 5646 34508 5660 34513
rect 5660 34508 5669 34513
rect 5696 34508 5712 34513
rect 5712 34508 5752 34513
rect 5779 34508 5835 34564
rect 5861 34508 5917 34564
rect 5943 34508 5999 34564
rect 6025 34508 6081 34564
rect 6107 34530 6148 34564
rect 6148 34530 6163 34564
rect 6189 34530 6200 34564
rect 6200 34530 6214 34564
rect 6214 34530 6245 34564
rect 6107 34513 6163 34530
rect 6189 34513 6245 34530
rect 6107 34508 6148 34513
rect 6148 34508 6163 34513
rect 6189 34508 6200 34513
rect 6200 34508 6214 34513
rect 6214 34508 6245 34513
rect 6271 34508 6327 34564
rect 6353 34508 6409 34564
rect 6435 34508 6491 34564
rect 6517 34508 6573 34564
rect 6599 34508 6655 34564
rect 6681 34530 6702 34564
rect 6702 34530 6737 34564
rect 6763 34530 6768 34564
rect 6768 34530 6819 34564
rect 6681 34513 6737 34530
rect 6763 34513 6819 34530
rect 6681 34508 6702 34513
rect 6702 34508 6737 34513
rect 6763 34508 6768 34513
rect 6768 34508 6819 34513
rect 6845 34508 6901 34564
rect 6927 34508 6983 34564
rect 7009 34508 7065 34564
rect 7091 34508 7147 34564
rect 7173 34508 7229 34564
rect 7255 34530 7256 34564
rect 7256 34530 7308 34564
rect 7308 34530 7311 34564
rect 7337 34530 7374 34564
rect 7374 34530 7393 34564
rect 7255 34513 7311 34530
rect 7337 34513 7393 34530
rect 7255 34508 7256 34513
rect 7256 34508 7308 34513
rect 7308 34508 7311 34513
rect 7337 34508 7374 34513
rect 7374 34508 7393 34513
rect 7419 34508 7475 34564
rect 7501 34508 7557 34564
rect 7583 34508 7639 34564
rect 7665 34508 7721 34564
rect 7747 34508 7803 34564
rect 7829 34530 7862 34564
rect 7862 34530 7876 34564
rect 7876 34530 7885 34564
rect 7911 34530 7928 34564
rect 7928 34530 7967 34564
rect 7829 34513 7885 34530
rect 7911 34513 7967 34530
rect 7829 34508 7862 34513
rect 7862 34508 7876 34513
rect 7876 34508 7885 34513
rect 7911 34508 7928 34513
rect 7928 34508 7967 34513
rect 7993 34534 8047 34564
rect 8047 34534 8049 34564
rect 8075 34534 8099 34564
rect 8099 34534 8131 34564
rect 7993 34517 8049 34534
rect 8075 34517 8131 34534
rect 7993 34508 8047 34517
rect 8047 34508 8049 34517
rect 8075 34508 8099 34517
rect 8099 34508 8131 34517
rect 8157 34534 8169 34564
rect 8169 34534 8213 34564
rect 8157 34517 8213 34534
rect 8157 34508 8169 34517
rect 8169 34508 8213 34517
rect 5613 34461 5646 34484
rect 5646 34461 5660 34484
rect 5660 34461 5669 34484
rect 5696 34461 5712 34484
rect 5712 34461 5752 34484
rect 5613 34444 5669 34461
rect 5696 34444 5752 34461
rect 5613 34428 5646 34444
rect 5646 34428 5660 34444
rect 5660 34428 5669 34444
rect 5696 34428 5712 34444
rect 5712 34428 5752 34444
rect 5779 34428 5835 34484
rect 5861 34428 5917 34484
rect 5943 34428 5999 34484
rect 6025 34428 6081 34484
rect 6107 34461 6148 34484
rect 6148 34461 6163 34484
rect 6189 34461 6200 34484
rect 6200 34461 6214 34484
rect 6214 34461 6245 34484
rect 6107 34444 6163 34461
rect 6189 34444 6245 34461
rect 6107 34428 6148 34444
rect 6148 34428 6163 34444
rect 6189 34428 6200 34444
rect 6200 34428 6214 34444
rect 6214 34428 6245 34444
rect 6271 34428 6327 34484
rect 6353 34428 6409 34484
rect 6435 34428 6491 34484
rect 6517 34428 6573 34484
rect 6599 34428 6655 34484
rect 6681 34461 6702 34484
rect 6702 34461 6737 34484
rect 6763 34461 6768 34484
rect 6768 34461 6819 34484
rect 6681 34444 6737 34461
rect 6763 34444 6819 34461
rect 6681 34428 6702 34444
rect 6702 34428 6737 34444
rect 6763 34428 6768 34444
rect 6768 34428 6819 34444
rect 6845 34428 6901 34484
rect 6927 34428 6983 34484
rect 7009 34428 7065 34484
rect 7091 34428 7147 34484
rect 7173 34428 7229 34484
rect 7255 34461 7256 34484
rect 7256 34461 7308 34484
rect 7308 34461 7311 34484
rect 7337 34461 7374 34484
rect 7374 34461 7393 34484
rect 7255 34444 7311 34461
rect 7337 34444 7393 34461
rect 7255 34428 7256 34444
rect 7256 34428 7308 34444
rect 7308 34428 7311 34444
rect 7337 34428 7374 34444
rect 7374 34428 7393 34444
rect 7419 34428 7475 34484
rect 7501 34428 7557 34484
rect 7583 34428 7639 34484
rect 7665 34428 7721 34484
rect 7747 34428 7803 34484
rect 7829 34461 7862 34484
rect 7862 34461 7876 34484
rect 7876 34461 7885 34484
rect 7911 34461 7928 34484
rect 7928 34461 7967 34484
rect 7829 34444 7885 34461
rect 7911 34444 7967 34461
rect 7829 34428 7862 34444
rect 7862 34428 7876 34444
rect 7876 34428 7885 34444
rect 7911 34428 7928 34444
rect 7928 34428 7967 34444
rect 7993 34465 8047 34484
rect 8047 34465 8049 34484
rect 8075 34465 8099 34484
rect 8099 34465 8131 34484
rect 7993 34448 8049 34465
rect 8075 34448 8131 34465
rect 7993 34428 8047 34448
rect 8047 34428 8049 34448
rect 8075 34428 8099 34448
rect 8099 34428 8131 34448
rect 8157 34465 8169 34484
rect 8169 34465 8213 34484
rect 8157 34448 8213 34465
rect 8157 34428 8169 34448
rect 8169 34428 8213 34448
rect 5613 34392 5646 34404
rect 5646 34392 5660 34404
rect 5660 34392 5669 34404
rect 5696 34392 5712 34404
rect 5712 34392 5752 34404
rect 5613 34375 5669 34392
rect 5696 34375 5752 34392
rect 5613 34348 5646 34375
rect 5646 34348 5660 34375
rect 5660 34348 5669 34375
rect 5696 34348 5712 34375
rect 5712 34348 5752 34375
rect 5779 34348 5835 34404
rect 5861 34348 5917 34404
rect 5943 34348 5999 34404
rect 6025 34348 6081 34404
rect 6107 34392 6148 34404
rect 6148 34392 6163 34404
rect 6189 34392 6200 34404
rect 6200 34392 6214 34404
rect 6214 34392 6245 34404
rect 6107 34375 6163 34392
rect 6189 34375 6245 34392
rect 6107 34348 6148 34375
rect 6148 34348 6163 34375
rect 6189 34348 6200 34375
rect 6200 34348 6214 34375
rect 6214 34348 6245 34375
rect 6271 34348 6327 34404
rect 6353 34348 6409 34404
rect 6435 34348 6491 34404
rect 6517 34348 6573 34404
rect 6599 34348 6655 34404
rect 6681 34392 6702 34404
rect 6702 34392 6737 34404
rect 6763 34392 6768 34404
rect 6768 34392 6819 34404
rect 6681 34375 6737 34392
rect 6763 34375 6819 34392
rect 6681 34348 6702 34375
rect 6702 34348 6737 34375
rect 6763 34348 6768 34375
rect 6768 34348 6819 34375
rect 6845 34348 6901 34404
rect 6927 34348 6983 34404
rect 7009 34348 7065 34404
rect 7091 34348 7147 34404
rect 7173 34348 7229 34404
rect 7255 34392 7256 34404
rect 7256 34392 7308 34404
rect 7308 34392 7311 34404
rect 7337 34392 7374 34404
rect 7374 34392 7393 34404
rect 7255 34375 7311 34392
rect 7337 34375 7393 34392
rect 7255 34348 7256 34375
rect 7256 34348 7308 34375
rect 7308 34348 7311 34375
rect 7337 34348 7374 34375
rect 7374 34348 7393 34375
rect 7419 34348 7475 34404
rect 7501 34348 7557 34404
rect 7583 34348 7639 34404
rect 7665 34348 7721 34404
rect 7747 34348 7803 34404
rect 7829 34392 7862 34404
rect 7862 34392 7876 34404
rect 7876 34392 7885 34404
rect 7911 34392 7928 34404
rect 7928 34392 7967 34404
rect 7829 34375 7885 34392
rect 7911 34375 7967 34392
rect 7829 34348 7862 34375
rect 7862 34348 7876 34375
rect 7876 34348 7885 34375
rect 7911 34348 7928 34375
rect 7928 34348 7967 34375
rect 7993 34396 8047 34404
rect 8047 34396 8049 34404
rect 8075 34396 8099 34404
rect 8099 34396 8131 34404
rect 7993 34378 8049 34396
rect 8075 34378 8131 34396
rect 7993 34348 8047 34378
rect 8047 34348 8049 34378
rect 8075 34348 8099 34378
rect 8099 34348 8131 34378
rect 8157 34396 8169 34404
rect 8169 34396 8213 34404
rect 8157 34378 8213 34396
rect 8157 34348 8169 34378
rect 8169 34348 8213 34378
rect 5613 34323 5646 34324
rect 5646 34323 5660 34324
rect 5660 34323 5669 34324
rect 5696 34323 5712 34324
rect 5712 34323 5752 34324
rect 5613 34306 5669 34323
rect 5696 34306 5752 34323
rect 5613 34268 5646 34306
rect 5646 34268 5660 34306
rect 5660 34268 5669 34306
rect 5696 34268 5712 34306
rect 5712 34268 5752 34306
rect 5779 34268 5835 34324
rect 5861 34268 5917 34324
rect 5943 34268 5999 34324
rect 6025 34268 6081 34324
rect 6107 34323 6148 34324
rect 6148 34323 6163 34324
rect 6189 34323 6200 34324
rect 6200 34323 6214 34324
rect 6214 34323 6245 34324
rect 6107 34306 6163 34323
rect 6189 34306 6245 34323
rect 6107 34268 6148 34306
rect 6148 34268 6163 34306
rect 6189 34268 6200 34306
rect 6200 34268 6214 34306
rect 6214 34268 6245 34306
rect 6271 34268 6327 34324
rect 6353 34268 6409 34324
rect 6435 34268 6491 34324
rect 6517 34268 6573 34324
rect 6599 34268 6655 34324
rect 6681 34323 6702 34324
rect 6702 34323 6737 34324
rect 6763 34323 6768 34324
rect 6768 34323 6819 34324
rect 6681 34306 6737 34323
rect 6763 34306 6819 34323
rect 6681 34268 6702 34306
rect 6702 34268 6737 34306
rect 6763 34268 6768 34306
rect 6768 34268 6819 34306
rect 6845 34268 6901 34324
rect 6927 34268 6983 34324
rect 7009 34268 7065 34324
rect 7091 34268 7147 34324
rect 7173 34268 7229 34324
rect 7255 34323 7256 34324
rect 7256 34323 7308 34324
rect 7308 34323 7311 34324
rect 7337 34323 7374 34324
rect 7374 34323 7393 34324
rect 7255 34306 7311 34323
rect 7337 34306 7393 34323
rect 7255 34268 7256 34306
rect 7256 34268 7308 34306
rect 7308 34268 7311 34306
rect 7337 34268 7374 34306
rect 7374 34268 7393 34306
rect 7419 34268 7475 34324
rect 7501 34268 7557 34324
rect 7583 34268 7639 34324
rect 7665 34268 7721 34324
rect 7747 34268 7803 34324
rect 7829 34323 7862 34324
rect 7862 34323 7876 34324
rect 7876 34323 7885 34324
rect 7911 34323 7928 34324
rect 7928 34323 7967 34324
rect 7829 34306 7885 34323
rect 7911 34306 7967 34323
rect 7829 34268 7862 34306
rect 7862 34268 7876 34306
rect 7876 34268 7885 34306
rect 7911 34268 7928 34306
rect 7928 34268 7967 34306
rect 7993 34308 8049 34324
rect 8075 34308 8131 34324
rect 7993 34268 8047 34308
rect 8047 34268 8049 34308
rect 8075 34268 8099 34308
rect 8099 34268 8131 34308
rect 8157 34308 8213 34324
rect 8157 34268 8169 34308
rect 8169 34268 8213 34308
rect 5613 34236 5669 34244
rect 5696 34236 5752 34244
rect 5613 34188 5646 34236
rect 5646 34188 5660 34236
rect 5660 34188 5669 34236
rect 5696 34188 5712 34236
rect 5712 34188 5752 34236
rect 5779 34188 5835 34244
rect 5861 34188 5917 34244
rect 5943 34188 5999 34244
rect 6025 34188 6081 34244
rect 6107 34236 6163 34244
rect 6189 34236 6245 34244
rect 6107 34188 6148 34236
rect 6148 34188 6163 34236
rect 6189 34188 6200 34236
rect 6200 34188 6214 34236
rect 6214 34188 6245 34236
rect 6271 34188 6327 34244
rect 6353 34188 6409 34244
rect 6435 34188 6491 34244
rect 6517 34188 6573 34244
rect 6599 34188 6655 34244
rect 6681 34236 6737 34244
rect 6763 34236 6819 34244
rect 6681 34188 6702 34236
rect 6702 34188 6737 34236
rect 6763 34188 6768 34236
rect 6768 34188 6819 34236
rect 6845 34188 6901 34244
rect 6927 34188 6983 34244
rect 7009 34188 7065 34244
rect 7091 34188 7147 34244
rect 7173 34188 7229 34244
rect 7255 34236 7311 34244
rect 7337 34236 7393 34244
rect 7255 34188 7256 34236
rect 7256 34188 7308 34236
rect 7308 34188 7311 34236
rect 7337 34188 7374 34236
rect 7374 34188 7393 34236
rect 7419 34188 7475 34244
rect 7501 34188 7557 34244
rect 7583 34188 7639 34244
rect 7665 34188 7721 34244
rect 7747 34188 7803 34244
rect 7829 34236 7885 34244
rect 7911 34236 7967 34244
rect 7829 34188 7862 34236
rect 7862 34188 7876 34236
rect 7876 34188 7885 34236
rect 7911 34188 7928 34236
rect 7928 34188 7967 34236
rect 7993 34238 8049 34244
rect 8075 34238 8131 34244
rect 7993 34188 8047 34238
rect 8047 34188 8049 34238
rect 8075 34188 8099 34238
rect 8099 34188 8131 34238
rect 8157 34238 8213 34244
rect 8157 34188 8169 34238
rect 8169 34188 8213 34238
rect 5613 34114 5646 34164
rect 5646 34114 5660 34164
rect 5660 34114 5669 34164
rect 5696 34114 5712 34164
rect 5712 34114 5752 34164
rect 5613 34108 5669 34114
rect 5696 34108 5752 34114
rect 5779 34108 5835 34164
rect 5861 34108 5917 34164
rect 5943 34108 5999 34164
rect 6025 34108 6081 34164
rect 6107 34114 6148 34164
rect 6148 34114 6163 34164
rect 6189 34114 6200 34164
rect 6200 34114 6214 34164
rect 6214 34114 6245 34164
rect 6107 34108 6163 34114
rect 6189 34108 6245 34114
rect 6271 34108 6327 34164
rect 6353 34108 6409 34164
rect 6435 34108 6491 34164
rect 6517 34108 6573 34164
rect 6599 34108 6655 34164
rect 6681 34114 6702 34164
rect 6702 34114 6737 34164
rect 6763 34114 6768 34164
rect 6768 34114 6819 34164
rect 6681 34108 6737 34114
rect 6763 34108 6819 34114
rect 6845 34108 6901 34164
rect 6927 34108 6983 34164
rect 7009 34108 7065 34164
rect 7091 34108 7147 34164
rect 7173 34108 7229 34164
rect 7255 34114 7256 34164
rect 7256 34114 7308 34164
rect 7308 34114 7311 34164
rect 7337 34114 7374 34164
rect 7374 34114 7393 34164
rect 7255 34108 7311 34114
rect 7337 34108 7393 34114
rect 7419 34108 7475 34164
rect 7501 34108 7557 34164
rect 7583 34108 7639 34164
rect 7665 34108 7721 34164
rect 7747 34108 7803 34164
rect 7829 34114 7862 34164
rect 7862 34114 7876 34164
rect 7876 34114 7885 34164
rect 7911 34114 7928 34164
rect 7928 34114 7967 34164
rect 7829 34108 7885 34114
rect 7911 34108 7967 34114
rect 7993 34116 8047 34164
rect 8047 34116 8049 34164
rect 8075 34116 8099 34164
rect 8099 34116 8131 34164
rect 7993 34108 8049 34116
rect 8075 34108 8131 34116
rect 8157 34116 8169 34164
rect 8169 34116 8213 34164
rect 8157 34108 8213 34116
rect 2733 33931 2789 33987
rect 2814 33931 2870 33987
rect 2895 33931 2951 33987
rect 2976 33931 3032 33987
rect 3057 33982 3113 33987
rect 3138 33982 3194 33987
rect 3057 33931 3101 33982
rect 3101 33931 3113 33982
rect 3138 33931 3153 33982
rect 3153 33931 3167 33982
rect 3167 33931 3194 33982
rect 3219 33931 3275 33987
rect 3300 33931 3356 33987
rect 3381 33931 3437 33987
rect 3462 33931 3518 33987
rect 3543 33931 3599 33987
rect 3624 33982 3680 33987
rect 3705 33982 3761 33987
rect 3624 33931 3655 33982
rect 3655 33931 3680 33982
rect 3705 33931 3707 33982
rect 3707 33931 3721 33982
rect 3721 33931 3761 33982
rect 3786 33931 3842 33987
rect 3867 33931 3923 33987
rect 3948 33931 4004 33987
rect 4029 33931 4085 33987
rect 4110 33931 4166 33987
rect 4191 33982 4247 33987
rect 4272 33982 4328 33987
rect 4191 33931 4209 33982
rect 4209 33931 4247 33982
rect 4272 33931 4275 33982
rect 4275 33931 4327 33982
rect 4327 33931 4328 33982
rect 4353 33931 4409 33987
rect 4434 33931 4490 33987
rect 4515 33931 4571 33987
rect 4596 33931 4652 33987
rect 4677 33931 4733 33987
rect 4758 33982 4814 33987
rect 4839 33982 4895 33987
rect 4758 33931 4763 33982
rect 4763 33931 4814 33982
rect 4839 33931 4881 33982
rect 4881 33931 4895 33982
rect 4920 33931 4976 33987
rect 5001 33931 5057 33987
rect 5082 33931 5138 33987
rect 2733 33851 2789 33907
rect 2814 33851 2870 33907
rect 2895 33851 2951 33907
rect 2976 33851 3032 33907
rect 3057 33861 3101 33907
rect 3101 33861 3113 33907
rect 3138 33861 3153 33907
rect 3153 33861 3167 33907
rect 3167 33861 3194 33907
rect 3057 33851 3113 33861
rect 3138 33851 3194 33861
rect 3219 33851 3275 33907
rect 3300 33851 3356 33907
rect 3381 33851 3437 33907
rect 3462 33851 3518 33907
rect 3543 33851 3599 33907
rect 3624 33861 3655 33907
rect 3655 33861 3680 33907
rect 3705 33861 3707 33907
rect 3707 33861 3721 33907
rect 3721 33861 3761 33907
rect 3624 33851 3680 33861
rect 3705 33851 3761 33861
rect 3786 33851 3842 33907
rect 3867 33851 3923 33907
rect 3948 33851 4004 33907
rect 4029 33851 4085 33907
rect 4110 33851 4166 33907
rect 4191 33861 4209 33907
rect 4209 33861 4247 33907
rect 4272 33861 4275 33907
rect 4275 33861 4327 33907
rect 4327 33861 4328 33907
rect 4191 33851 4247 33861
rect 4272 33851 4328 33861
rect 4353 33851 4409 33907
rect 4434 33851 4490 33907
rect 4515 33851 4571 33907
rect 4596 33851 4652 33907
rect 4677 33851 4733 33907
rect 4758 33861 4763 33907
rect 4763 33861 4814 33907
rect 4839 33861 4881 33907
rect 4881 33861 4895 33907
rect 4758 33851 4814 33861
rect 4839 33851 4895 33861
rect 4920 33851 4976 33907
rect 5001 33851 5057 33907
rect 5082 33851 5138 33907
rect 2733 33771 2789 33827
rect 2814 33771 2870 33827
rect 2895 33771 2951 33827
rect 2976 33771 3032 33827
rect 3057 33792 3101 33827
rect 3101 33792 3113 33827
rect 3138 33792 3153 33827
rect 3153 33792 3167 33827
rect 3167 33792 3194 33827
rect 3057 33775 3113 33792
rect 3138 33775 3194 33792
rect 3057 33771 3101 33775
rect 3101 33771 3113 33775
rect 3138 33771 3153 33775
rect 3153 33771 3167 33775
rect 3167 33771 3194 33775
rect 3219 33771 3275 33827
rect 3300 33771 3356 33827
rect 3381 33771 3437 33827
rect 3462 33771 3518 33827
rect 3543 33771 3599 33827
rect 3624 33792 3655 33827
rect 3655 33792 3680 33827
rect 3705 33792 3707 33827
rect 3707 33792 3721 33827
rect 3721 33792 3761 33827
rect 3624 33775 3680 33792
rect 3705 33775 3761 33792
rect 3624 33771 3655 33775
rect 3655 33771 3680 33775
rect 3705 33771 3707 33775
rect 3707 33771 3721 33775
rect 3721 33771 3761 33775
rect 3786 33771 3842 33827
rect 3867 33771 3923 33827
rect 3948 33771 4004 33827
rect 4029 33771 4085 33827
rect 4110 33771 4166 33827
rect 4191 33792 4209 33827
rect 4209 33792 4247 33827
rect 4272 33792 4275 33827
rect 4275 33792 4327 33827
rect 4327 33792 4328 33827
rect 4191 33775 4247 33792
rect 4272 33775 4328 33792
rect 4191 33771 4209 33775
rect 4209 33771 4247 33775
rect 4272 33771 4275 33775
rect 4275 33771 4327 33775
rect 4327 33771 4328 33775
rect 4353 33771 4409 33827
rect 4434 33771 4490 33827
rect 4515 33771 4571 33827
rect 4596 33771 4652 33827
rect 4677 33771 4733 33827
rect 4758 33792 4763 33827
rect 4763 33792 4814 33827
rect 4839 33792 4881 33827
rect 4881 33792 4895 33827
rect 4758 33775 4814 33792
rect 4839 33775 4895 33792
rect 4758 33771 4763 33775
rect 4763 33771 4814 33775
rect 2733 33691 2789 33747
rect 2814 33691 2870 33747
rect 2895 33691 2951 33747
rect 2976 33691 3032 33747
rect 3057 33723 3101 33747
rect 3101 33723 3113 33747
rect 3138 33723 3153 33747
rect 3153 33723 3167 33747
rect 3167 33723 3194 33747
rect 3057 33706 3113 33723
rect 3138 33706 3194 33723
rect 3057 33691 3101 33706
rect 3101 33691 3113 33706
rect 3138 33691 3153 33706
rect 3153 33691 3167 33706
rect 3167 33691 3194 33706
rect 3219 33691 3275 33747
rect 3300 33691 3356 33747
rect 3381 33691 3437 33747
rect 3462 33691 3518 33747
rect 3543 33691 3599 33747
rect 3624 33723 3655 33747
rect 3655 33723 3680 33747
rect 3705 33723 3707 33747
rect 3707 33723 3721 33747
rect 3721 33723 3761 33747
rect 3624 33706 3680 33723
rect 3705 33706 3761 33723
rect 3624 33691 3655 33706
rect 3655 33691 3680 33706
rect 3705 33691 3707 33706
rect 3707 33691 3721 33706
rect 3721 33691 3761 33706
rect 3786 33691 3842 33747
rect 3867 33691 3923 33747
rect 3948 33691 4004 33747
rect 4029 33691 4085 33747
rect 4110 33691 4166 33747
rect 4191 33723 4209 33747
rect 4209 33723 4247 33747
rect 4272 33723 4275 33747
rect 4275 33723 4327 33747
rect 4327 33723 4328 33747
rect 4191 33706 4247 33723
rect 4272 33706 4328 33723
rect 4191 33691 4209 33706
rect 4209 33691 4247 33706
rect 4272 33691 4275 33706
rect 4275 33691 4327 33706
rect 4327 33691 4328 33706
rect 4353 33691 4409 33747
rect 4434 33691 4490 33747
rect 4515 33691 4571 33747
rect 4596 33691 4652 33747
rect 4677 33691 4733 33747
rect 4758 33723 4763 33747
rect 4763 33723 4814 33747
rect 4839 33771 4881 33775
rect 4881 33771 4895 33775
rect 4920 33771 4976 33827
rect 5001 33771 5057 33827
rect 5082 33771 5138 33827
rect 4839 33723 4881 33747
rect 4881 33723 4895 33747
rect 4758 33706 4814 33723
rect 4839 33706 4895 33723
rect 4758 33691 4763 33706
rect 4763 33691 4814 33706
rect 2733 33611 2789 33667
rect 2814 33611 2870 33667
rect 2895 33611 2951 33667
rect 2976 33611 3032 33667
rect 3057 33654 3101 33667
rect 3101 33654 3113 33667
rect 3138 33654 3153 33667
rect 3153 33654 3167 33667
rect 3167 33654 3194 33667
rect 3057 33636 3113 33654
rect 3138 33636 3194 33654
rect 3057 33611 3101 33636
rect 3101 33611 3113 33636
rect 3138 33611 3153 33636
rect 3153 33611 3167 33636
rect 3167 33611 3194 33636
rect 3219 33611 3275 33667
rect 3300 33611 3356 33667
rect 3381 33611 3437 33667
rect 3462 33611 3518 33667
rect 3543 33611 3599 33667
rect 3624 33654 3655 33667
rect 3655 33654 3680 33667
rect 3705 33654 3707 33667
rect 3707 33654 3721 33667
rect 3721 33654 3761 33667
rect 3624 33636 3680 33654
rect 3705 33636 3761 33654
rect 3624 33611 3655 33636
rect 3655 33611 3680 33636
rect 3705 33611 3707 33636
rect 3707 33611 3721 33636
rect 3721 33611 3761 33636
rect 3786 33611 3842 33667
rect 3867 33611 3923 33667
rect 3948 33611 4004 33667
rect 4029 33611 4085 33667
rect 4110 33611 4166 33667
rect 4191 33654 4209 33667
rect 4209 33654 4247 33667
rect 4272 33654 4275 33667
rect 4275 33654 4327 33667
rect 4327 33654 4328 33667
rect 4191 33636 4247 33654
rect 4272 33636 4328 33654
rect 4191 33611 4209 33636
rect 4209 33611 4247 33636
rect 4272 33611 4275 33636
rect 4275 33611 4327 33636
rect 4327 33611 4328 33636
rect 4353 33611 4409 33667
rect 4434 33611 4490 33667
rect 4515 33611 4571 33667
rect 4596 33611 4652 33667
rect 4677 33611 4733 33667
rect 4758 33654 4763 33667
rect 4763 33654 4814 33667
rect 4839 33691 4881 33706
rect 4881 33691 4895 33706
rect 4920 33691 4976 33747
rect 5001 33691 5057 33747
rect 5082 33691 5138 33747
rect 4839 33654 4881 33667
rect 4881 33654 4895 33667
rect 4758 33636 4814 33654
rect 4839 33636 4895 33654
rect 4758 33611 4763 33636
rect 4763 33611 4814 33636
rect 2733 33531 2789 33587
rect 2814 33531 2870 33587
rect 2895 33531 2951 33587
rect 2976 33531 3032 33587
rect 3057 33584 3101 33587
rect 3101 33584 3113 33587
rect 3138 33584 3153 33587
rect 3153 33584 3167 33587
rect 3167 33584 3194 33587
rect 3057 33566 3113 33584
rect 3138 33566 3194 33584
rect 3057 33531 3101 33566
rect 3101 33531 3113 33566
rect 3138 33531 3153 33566
rect 3153 33531 3167 33566
rect 3167 33531 3194 33566
rect 3219 33531 3275 33587
rect 3300 33531 3356 33587
rect 3381 33531 3437 33587
rect 3462 33531 3518 33587
rect 3543 33531 3599 33587
rect 3624 33584 3655 33587
rect 3655 33584 3680 33587
rect 3705 33584 3707 33587
rect 3707 33584 3721 33587
rect 3721 33584 3761 33587
rect 3624 33566 3680 33584
rect 3705 33566 3761 33584
rect 3624 33531 3655 33566
rect 3655 33531 3680 33566
rect 3705 33531 3707 33566
rect 3707 33531 3721 33566
rect 3721 33531 3761 33566
rect 3786 33531 3842 33587
rect 3867 33531 3923 33587
rect 3948 33531 4004 33587
rect 4029 33531 4085 33587
rect 4110 33531 4166 33587
rect 4191 33584 4209 33587
rect 4209 33584 4247 33587
rect 4272 33584 4275 33587
rect 4275 33584 4327 33587
rect 4327 33584 4328 33587
rect 4191 33566 4247 33584
rect 4272 33566 4328 33584
rect 4191 33531 4209 33566
rect 4209 33531 4247 33566
rect 4272 33531 4275 33566
rect 4275 33531 4327 33566
rect 4327 33531 4328 33566
rect 4353 33531 4409 33587
rect 4434 33531 4490 33587
rect 4515 33531 4571 33587
rect 4596 33531 4652 33587
rect 4677 33531 4733 33587
rect 4758 33584 4763 33587
rect 4763 33584 4814 33587
rect 4839 33611 4881 33636
rect 4881 33611 4895 33636
rect 4920 33611 4976 33667
rect 5001 33611 5057 33667
rect 5082 33611 5138 33667
rect 4839 33584 4881 33587
rect 4881 33584 4895 33587
rect 4758 33566 4814 33584
rect 4839 33566 4895 33584
rect 4758 33531 4763 33566
rect 4763 33531 4814 33566
rect 4839 33531 4881 33566
rect 4881 33531 4895 33566
rect 4920 33531 4976 33587
rect 5001 33531 5057 33587
rect 5082 33531 5138 33587
rect 2733 33451 2789 33507
rect 2814 33451 2870 33507
rect 2895 33451 2951 33507
rect 2976 33451 3032 33507
rect 3057 33496 3113 33507
rect 3138 33496 3194 33507
rect 3057 33451 3101 33496
rect 3101 33451 3113 33496
rect 3138 33451 3153 33496
rect 3153 33451 3167 33496
rect 3167 33451 3194 33496
rect 3219 33451 3275 33507
rect 3300 33451 3356 33507
rect 3381 33451 3437 33507
rect 3462 33451 3518 33507
rect 3543 33451 3599 33507
rect 3624 33496 3680 33507
rect 3705 33496 3761 33507
rect 3624 33451 3655 33496
rect 3655 33451 3680 33496
rect 3705 33451 3707 33496
rect 3707 33451 3721 33496
rect 3721 33451 3761 33496
rect 3786 33451 3842 33507
rect 3867 33451 3923 33507
rect 3948 33451 4004 33507
rect 4029 33451 4085 33507
rect 4110 33451 4166 33507
rect 4191 33496 4247 33507
rect 4272 33496 4328 33507
rect 4191 33451 4209 33496
rect 4209 33451 4247 33496
rect 4272 33451 4275 33496
rect 4275 33451 4327 33496
rect 4327 33451 4328 33496
rect 4353 33451 4409 33507
rect 4434 33451 4490 33507
rect 4515 33451 4571 33507
rect 4596 33451 4652 33507
rect 4677 33451 4733 33507
rect 4758 33496 4814 33507
rect 4839 33496 4895 33507
rect 4758 33451 4763 33496
rect 4763 33451 4814 33496
rect 4839 33451 4881 33496
rect 4881 33451 4895 33496
rect 4920 33451 4976 33507
rect 5001 33451 5057 33507
rect 5082 33451 5138 33507
rect 2733 33371 2789 33427
rect 2814 33371 2870 33427
rect 2895 33371 2951 33427
rect 2976 33371 3032 33427
rect 3057 33426 3113 33427
rect 3138 33426 3194 33427
rect 3057 33374 3101 33426
rect 3101 33374 3113 33426
rect 3138 33374 3153 33426
rect 3153 33374 3167 33426
rect 3167 33374 3194 33426
rect 3057 33371 3113 33374
rect 3138 33371 3194 33374
rect 3219 33371 3275 33427
rect 3300 33371 3356 33427
rect 3381 33371 3437 33427
rect 3462 33371 3518 33427
rect 3543 33371 3599 33427
rect 3624 33426 3680 33427
rect 3705 33426 3761 33427
rect 3624 33374 3655 33426
rect 3655 33374 3680 33426
rect 3705 33374 3707 33426
rect 3707 33374 3721 33426
rect 3721 33374 3761 33426
rect 3624 33371 3680 33374
rect 3705 33371 3761 33374
rect 3786 33371 3842 33427
rect 3867 33371 3923 33427
rect 3948 33371 4004 33427
rect 4029 33371 4085 33427
rect 4110 33371 4166 33427
rect 4191 33426 4247 33427
rect 4272 33426 4328 33427
rect 4191 33374 4209 33426
rect 4209 33374 4247 33426
rect 4272 33374 4275 33426
rect 4275 33374 4327 33426
rect 4327 33374 4328 33426
rect 4191 33371 4247 33374
rect 4272 33371 4328 33374
rect 4353 33371 4409 33427
rect 4434 33371 4490 33427
rect 4515 33371 4571 33427
rect 4596 33371 4652 33427
rect 4677 33371 4733 33427
rect 4758 33426 4814 33427
rect 4839 33426 4895 33427
rect 4758 33374 4763 33426
rect 4763 33374 4814 33426
rect 4839 33374 4881 33426
rect 4881 33374 4895 33426
rect 4758 33371 4814 33374
rect 4839 33371 4895 33374
rect 4920 33371 4976 33427
rect 5001 33371 5057 33427
rect 5082 33371 5138 33427
rect 5163 33371 5299 33987
rect 5613 32720 5669 32724
rect 5696 32720 5752 32724
rect 5613 32668 5646 32720
rect 5646 32668 5660 32720
rect 5660 32668 5669 32720
rect 5696 32668 5712 32720
rect 5712 32668 5752 32720
rect 5779 32668 5835 32724
rect 5861 32668 5917 32724
rect 5943 32668 5999 32724
rect 6025 32668 6081 32724
rect 6107 32720 6163 32724
rect 6189 32720 6245 32724
rect 6107 32668 6148 32720
rect 6148 32668 6163 32720
rect 6189 32668 6200 32720
rect 6200 32668 6214 32720
rect 6214 32668 6245 32720
rect 6271 32668 6327 32724
rect 6353 32668 6409 32724
rect 6435 32668 6491 32724
rect 6517 32668 6573 32724
rect 6599 32668 6655 32724
rect 6681 32720 6737 32724
rect 6763 32720 6819 32724
rect 6681 32668 6702 32720
rect 6702 32668 6737 32720
rect 6763 32668 6768 32720
rect 6768 32668 6819 32720
rect 6845 32668 6901 32724
rect 6927 32668 6983 32724
rect 7009 32668 7065 32724
rect 7091 32668 7147 32724
rect 7173 32668 7229 32724
rect 7255 32720 7311 32724
rect 7337 32720 7393 32724
rect 7255 32668 7256 32720
rect 7256 32668 7308 32720
rect 7308 32668 7311 32720
rect 7337 32668 7374 32720
rect 7374 32668 7393 32720
rect 7419 32668 7475 32724
rect 7501 32668 7557 32724
rect 7583 32668 7639 32724
rect 7665 32668 7721 32724
rect 7747 32668 7803 32724
rect 7829 32720 7885 32724
rect 7911 32720 7967 32724
rect 7829 32668 7862 32720
rect 7862 32668 7876 32720
rect 7876 32668 7885 32720
rect 7911 32668 7928 32720
rect 7928 32668 7967 32720
rect 7993 32672 8047 32724
rect 8047 32672 8049 32724
rect 8075 32672 8099 32724
rect 8099 32672 8131 32724
rect 7993 32668 8049 32672
rect 8075 32668 8131 32672
rect 8157 32672 8169 32724
rect 8169 32672 8213 32724
rect 8157 32668 8213 32672
rect 5613 32599 5646 32644
rect 5646 32599 5660 32644
rect 5660 32599 5669 32644
rect 5696 32599 5712 32644
rect 5712 32599 5752 32644
rect 5613 32588 5669 32599
rect 5696 32588 5752 32599
rect 5779 32588 5835 32644
rect 5861 32588 5917 32644
rect 5943 32588 5999 32644
rect 6025 32588 6081 32644
rect 6107 32599 6148 32644
rect 6148 32599 6163 32644
rect 6189 32599 6200 32644
rect 6200 32599 6214 32644
rect 6214 32599 6245 32644
rect 6107 32588 6163 32599
rect 6189 32588 6245 32599
rect 6271 32588 6327 32644
rect 6353 32588 6409 32644
rect 6435 32588 6491 32644
rect 6517 32588 6573 32644
rect 6599 32588 6655 32644
rect 6681 32599 6702 32644
rect 6702 32599 6737 32644
rect 6763 32599 6768 32644
rect 6768 32599 6819 32644
rect 6681 32588 6737 32599
rect 6763 32588 6819 32599
rect 6845 32588 6901 32644
rect 6927 32588 6983 32644
rect 7009 32588 7065 32644
rect 7091 32588 7147 32644
rect 7173 32588 7229 32644
rect 7255 32599 7256 32644
rect 7256 32599 7308 32644
rect 7308 32599 7311 32644
rect 7337 32599 7374 32644
rect 7374 32599 7393 32644
rect 7255 32588 7311 32599
rect 7337 32588 7393 32599
rect 7419 32588 7475 32644
rect 7501 32588 7557 32644
rect 7583 32588 7639 32644
rect 7665 32588 7721 32644
rect 7747 32588 7803 32644
rect 7829 32599 7862 32644
rect 7862 32599 7876 32644
rect 7876 32599 7885 32644
rect 7911 32599 7928 32644
rect 7928 32599 7967 32644
rect 7829 32588 7885 32599
rect 7911 32588 7967 32599
rect 7993 32603 8047 32644
rect 8047 32603 8049 32644
rect 8075 32603 8099 32644
rect 8099 32603 8131 32644
rect 7993 32588 8049 32603
rect 8075 32588 8131 32603
rect 8157 32603 8169 32644
rect 8169 32603 8213 32644
rect 8157 32588 8213 32603
rect 5613 32530 5646 32564
rect 5646 32530 5660 32564
rect 5660 32530 5669 32564
rect 5696 32530 5712 32564
rect 5712 32530 5752 32564
rect 5613 32513 5669 32530
rect 5696 32513 5752 32530
rect 5613 32508 5646 32513
rect 5646 32508 5660 32513
rect 5660 32508 5669 32513
rect 5696 32508 5712 32513
rect 5712 32508 5752 32513
rect 5779 32508 5835 32564
rect 5861 32508 5917 32564
rect 5943 32508 5999 32564
rect 6025 32508 6081 32564
rect 6107 32530 6148 32564
rect 6148 32530 6163 32564
rect 6189 32530 6200 32564
rect 6200 32530 6214 32564
rect 6214 32530 6245 32564
rect 6107 32513 6163 32530
rect 6189 32513 6245 32530
rect 6107 32508 6148 32513
rect 6148 32508 6163 32513
rect 6189 32508 6200 32513
rect 6200 32508 6214 32513
rect 6214 32508 6245 32513
rect 6271 32508 6327 32564
rect 6353 32508 6409 32564
rect 6435 32508 6491 32564
rect 6517 32508 6573 32564
rect 6599 32508 6655 32564
rect 6681 32530 6702 32564
rect 6702 32530 6737 32564
rect 6763 32530 6768 32564
rect 6768 32530 6819 32564
rect 6681 32513 6737 32530
rect 6763 32513 6819 32530
rect 6681 32508 6702 32513
rect 6702 32508 6737 32513
rect 6763 32508 6768 32513
rect 6768 32508 6819 32513
rect 6845 32508 6901 32564
rect 6927 32508 6983 32564
rect 7009 32508 7065 32564
rect 7091 32508 7147 32564
rect 7173 32508 7229 32564
rect 7255 32530 7256 32564
rect 7256 32530 7308 32564
rect 7308 32530 7311 32564
rect 7337 32530 7374 32564
rect 7374 32530 7393 32564
rect 7255 32513 7311 32530
rect 7337 32513 7393 32530
rect 7255 32508 7256 32513
rect 7256 32508 7308 32513
rect 7308 32508 7311 32513
rect 7337 32508 7374 32513
rect 7374 32508 7393 32513
rect 7419 32508 7475 32564
rect 7501 32508 7557 32564
rect 7583 32508 7639 32564
rect 7665 32508 7721 32564
rect 7747 32508 7803 32564
rect 7829 32530 7862 32564
rect 7862 32530 7876 32564
rect 7876 32530 7885 32564
rect 7911 32530 7928 32564
rect 7928 32530 7967 32564
rect 7829 32513 7885 32530
rect 7911 32513 7967 32530
rect 7829 32508 7862 32513
rect 7862 32508 7876 32513
rect 7876 32508 7885 32513
rect 7911 32508 7928 32513
rect 7928 32508 7967 32513
rect 7993 32534 8047 32564
rect 8047 32534 8049 32564
rect 8075 32534 8099 32564
rect 8099 32534 8131 32564
rect 7993 32517 8049 32534
rect 8075 32517 8131 32534
rect 7993 32508 8047 32517
rect 8047 32508 8049 32517
rect 8075 32508 8099 32517
rect 8099 32508 8131 32517
rect 8157 32534 8169 32564
rect 8169 32534 8213 32564
rect 8157 32517 8213 32534
rect 8157 32508 8169 32517
rect 8169 32508 8213 32517
rect 5613 32461 5646 32484
rect 5646 32461 5660 32484
rect 5660 32461 5669 32484
rect 5696 32461 5712 32484
rect 5712 32461 5752 32484
rect 5613 32444 5669 32461
rect 5696 32444 5752 32461
rect 5613 32428 5646 32444
rect 5646 32428 5660 32444
rect 5660 32428 5669 32444
rect 5696 32428 5712 32444
rect 5712 32428 5752 32444
rect 5779 32428 5835 32484
rect 5861 32428 5917 32484
rect 5943 32428 5999 32484
rect 6025 32428 6081 32484
rect 6107 32461 6148 32484
rect 6148 32461 6163 32484
rect 6189 32461 6200 32484
rect 6200 32461 6214 32484
rect 6214 32461 6245 32484
rect 6107 32444 6163 32461
rect 6189 32444 6245 32461
rect 6107 32428 6148 32444
rect 6148 32428 6163 32444
rect 6189 32428 6200 32444
rect 6200 32428 6214 32444
rect 6214 32428 6245 32444
rect 6271 32428 6327 32484
rect 6353 32428 6409 32484
rect 6435 32428 6491 32484
rect 6517 32428 6573 32484
rect 6599 32428 6655 32484
rect 6681 32461 6702 32484
rect 6702 32461 6737 32484
rect 6763 32461 6768 32484
rect 6768 32461 6819 32484
rect 6681 32444 6737 32461
rect 6763 32444 6819 32461
rect 6681 32428 6702 32444
rect 6702 32428 6737 32444
rect 6763 32428 6768 32444
rect 6768 32428 6819 32444
rect 6845 32428 6901 32484
rect 6927 32428 6983 32484
rect 7009 32428 7065 32484
rect 7091 32428 7147 32484
rect 7173 32428 7229 32484
rect 7255 32461 7256 32484
rect 7256 32461 7308 32484
rect 7308 32461 7311 32484
rect 7337 32461 7374 32484
rect 7374 32461 7393 32484
rect 7255 32444 7311 32461
rect 7337 32444 7393 32461
rect 7255 32428 7256 32444
rect 7256 32428 7308 32444
rect 7308 32428 7311 32444
rect 7337 32428 7374 32444
rect 7374 32428 7393 32444
rect 7419 32428 7475 32484
rect 7501 32428 7557 32484
rect 7583 32428 7639 32484
rect 7665 32428 7721 32484
rect 7747 32428 7803 32484
rect 7829 32461 7862 32484
rect 7862 32461 7876 32484
rect 7876 32461 7885 32484
rect 7911 32461 7928 32484
rect 7928 32461 7967 32484
rect 7829 32444 7885 32461
rect 7911 32444 7967 32461
rect 7829 32428 7862 32444
rect 7862 32428 7876 32444
rect 7876 32428 7885 32444
rect 7911 32428 7928 32444
rect 7928 32428 7967 32444
rect 7993 32465 8047 32484
rect 8047 32465 8049 32484
rect 8075 32465 8099 32484
rect 8099 32465 8131 32484
rect 7993 32448 8049 32465
rect 8075 32448 8131 32465
rect 7993 32428 8047 32448
rect 8047 32428 8049 32448
rect 8075 32428 8099 32448
rect 8099 32428 8131 32448
rect 8157 32465 8169 32484
rect 8169 32465 8213 32484
rect 8157 32448 8213 32465
rect 8157 32428 8169 32448
rect 8169 32428 8213 32448
rect 5613 32392 5646 32404
rect 5646 32392 5660 32404
rect 5660 32392 5669 32404
rect 5696 32392 5712 32404
rect 5712 32392 5752 32404
rect 5613 32375 5669 32392
rect 5696 32375 5752 32392
rect 5613 32348 5646 32375
rect 5646 32348 5660 32375
rect 5660 32348 5669 32375
rect 5696 32348 5712 32375
rect 5712 32348 5752 32375
rect 5779 32348 5835 32404
rect 5861 32348 5917 32404
rect 5943 32348 5999 32404
rect 6025 32348 6081 32404
rect 6107 32392 6148 32404
rect 6148 32392 6163 32404
rect 6189 32392 6200 32404
rect 6200 32392 6214 32404
rect 6214 32392 6245 32404
rect 6107 32375 6163 32392
rect 6189 32375 6245 32392
rect 6107 32348 6148 32375
rect 6148 32348 6163 32375
rect 6189 32348 6200 32375
rect 6200 32348 6214 32375
rect 6214 32348 6245 32375
rect 6271 32348 6327 32404
rect 6353 32348 6409 32404
rect 6435 32348 6491 32404
rect 6517 32348 6573 32404
rect 6599 32348 6655 32404
rect 6681 32392 6702 32404
rect 6702 32392 6737 32404
rect 6763 32392 6768 32404
rect 6768 32392 6819 32404
rect 6681 32375 6737 32392
rect 6763 32375 6819 32392
rect 6681 32348 6702 32375
rect 6702 32348 6737 32375
rect 6763 32348 6768 32375
rect 6768 32348 6819 32375
rect 6845 32348 6901 32404
rect 6927 32348 6983 32404
rect 7009 32348 7065 32404
rect 7091 32348 7147 32404
rect 7173 32348 7229 32404
rect 7255 32392 7256 32404
rect 7256 32392 7308 32404
rect 7308 32392 7311 32404
rect 7337 32392 7374 32404
rect 7374 32392 7393 32404
rect 7255 32375 7311 32392
rect 7337 32375 7393 32392
rect 7255 32348 7256 32375
rect 7256 32348 7308 32375
rect 7308 32348 7311 32375
rect 7337 32348 7374 32375
rect 7374 32348 7393 32375
rect 7419 32348 7475 32404
rect 7501 32348 7557 32404
rect 7583 32348 7639 32404
rect 7665 32348 7721 32404
rect 7747 32348 7803 32404
rect 7829 32392 7862 32404
rect 7862 32392 7876 32404
rect 7876 32392 7885 32404
rect 7911 32392 7928 32404
rect 7928 32392 7967 32404
rect 7829 32375 7885 32392
rect 7911 32375 7967 32392
rect 7829 32348 7862 32375
rect 7862 32348 7876 32375
rect 7876 32348 7885 32375
rect 7911 32348 7928 32375
rect 7928 32348 7967 32375
rect 7993 32396 8047 32404
rect 8047 32396 8049 32404
rect 8075 32396 8099 32404
rect 8099 32396 8131 32404
rect 7993 32378 8049 32396
rect 8075 32378 8131 32396
rect 7993 32348 8047 32378
rect 8047 32348 8049 32378
rect 8075 32348 8099 32378
rect 8099 32348 8131 32378
rect 8157 32396 8169 32404
rect 8169 32396 8213 32404
rect 8157 32378 8213 32396
rect 8157 32348 8169 32378
rect 8169 32348 8213 32378
rect 5613 32323 5646 32324
rect 5646 32323 5660 32324
rect 5660 32323 5669 32324
rect 5696 32323 5712 32324
rect 5712 32323 5752 32324
rect 5613 32306 5669 32323
rect 5696 32306 5752 32323
rect 5613 32268 5646 32306
rect 5646 32268 5660 32306
rect 5660 32268 5669 32306
rect 5696 32268 5712 32306
rect 5712 32268 5752 32306
rect 5779 32268 5835 32324
rect 5861 32268 5917 32324
rect 5943 32268 5999 32324
rect 6025 32268 6081 32324
rect 6107 32323 6148 32324
rect 6148 32323 6163 32324
rect 6189 32323 6200 32324
rect 6200 32323 6214 32324
rect 6214 32323 6245 32324
rect 6107 32306 6163 32323
rect 6189 32306 6245 32323
rect 6107 32268 6148 32306
rect 6148 32268 6163 32306
rect 6189 32268 6200 32306
rect 6200 32268 6214 32306
rect 6214 32268 6245 32306
rect 6271 32268 6327 32324
rect 6353 32268 6409 32324
rect 6435 32268 6491 32324
rect 6517 32268 6573 32324
rect 6599 32268 6655 32324
rect 6681 32323 6702 32324
rect 6702 32323 6737 32324
rect 6763 32323 6768 32324
rect 6768 32323 6819 32324
rect 6681 32306 6737 32323
rect 6763 32306 6819 32323
rect 6681 32268 6702 32306
rect 6702 32268 6737 32306
rect 6763 32268 6768 32306
rect 6768 32268 6819 32306
rect 6845 32268 6901 32324
rect 6927 32268 6983 32324
rect 7009 32268 7065 32324
rect 7091 32268 7147 32324
rect 7173 32268 7229 32324
rect 7255 32323 7256 32324
rect 7256 32323 7308 32324
rect 7308 32323 7311 32324
rect 7337 32323 7374 32324
rect 7374 32323 7393 32324
rect 7255 32306 7311 32323
rect 7337 32306 7393 32323
rect 7255 32268 7256 32306
rect 7256 32268 7308 32306
rect 7308 32268 7311 32306
rect 7337 32268 7374 32306
rect 7374 32268 7393 32306
rect 7419 32268 7475 32324
rect 7501 32268 7557 32324
rect 7583 32268 7639 32324
rect 7665 32268 7721 32324
rect 7747 32268 7803 32324
rect 7829 32323 7862 32324
rect 7862 32323 7876 32324
rect 7876 32323 7885 32324
rect 7911 32323 7928 32324
rect 7928 32323 7967 32324
rect 7829 32306 7885 32323
rect 7911 32306 7967 32323
rect 7829 32268 7862 32306
rect 7862 32268 7876 32306
rect 7876 32268 7885 32306
rect 7911 32268 7928 32306
rect 7928 32268 7967 32306
rect 7993 32308 8049 32324
rect 8075 32308 8131 32324
rect 7993 32268 8047 32308
rect 8047 32268 8049 32308
rect 8075 32268 8099 32308
rect 8099 32268 8131 32308
rect 8157 32308 8213 32324
rect 8157 32268 8169 32308
rect 8169 32268 8213 32308
rect 5613 32236 5669 32244
rect 5696 32236 5752 32244
rect 5613 32188 5646 32236
rect 5646 32188 5660 32236
rect 5660 32188 5669 32236
rect 5696 32188 5712 32236
rect 5712 32188 5752 32236
rect 5779 32188 5835 32244
rect 5861 32188 5917 32244
rect 5943 32188 5999 32244
rect 6025 32188 6081 32244
rect 6107 32236 6163 32244
rect 6189 32236 6245 32244
rect 6107 32188 6148 32236
rect 6148 32188 6163 32236
rect 6189 32188 6200 32236
rect 6200 32188 6214 32236
rect 6214 32188 6245 32236
rect 6271 32188 6327 32244
rect 6353 32188 6409 32244
rect 6435 32188 6491 32244
rect 6517 32188 6573 32244
rect 6599 32188 6655 32244
rect 6681 32236 6737 32244
rect 6763 32236 6819 32244
rect 6681 32188 6702 32236
rect 6702 32188 6737 32236
rect 6763 32188 6768 32236
rect 6768 32188 6819 32236
rect 6845 32188 6901 32244
rect 6927 32188 6983 32244
rect 7009 32188 7065 32244
rect 7091 32188 7147 32244
rect 7173 32188 7229 32244
rect 7255 32236 7311 32244
rect 7337 32236 7393 32244
rect 7255 32188 7256 32236
rect 7256 32188 7308 32236
rect 7308 32188 7311 32236
rect 7337 32188 7374 32236
rect 7374 32188 7393 32236
rect 7419 32188 7475 32244
rect 7501 32188 7557 32244
rect 7583 32188 7639 32244
rect 7665 32188 7721 32244
rect 7747 32188 7803 32244
rect 7829 32236 7885 32244
rect 7911 32236 7967 32244
rect 7829 32188 7862 32236
rect 7862 32188 7876 32236
rect 7876 32188 7885 32236
rect 7911 32188 7928 32236
rect 7928 32188 7967 32236
rect 7993 32238 8049 32244
rect 8075 32238 8131 32244
rect 7993 32188 8047 32238
rect 8047 32188 8049 32238
rect 8075 32188 8099 32238
rect 8099 32188 8131 32238
rect 8157 32238 8213 32244
rect 8157 32188 8169 32238
rect 8169 32188 8213 32238
rect 5613 32114 5646 32164
rect 5646 32114 5660 32164
rect 5660 32114 5669 32164
rect 5696 32114 5712 32164
rect 5712 32114 5752 32164
rect 5613 32108 5669 32114
rect 5696 32108 5752 32114
rect 5779 32108 5835 32164
rect 5861 32108 5917 32164
rect 5943 32108 5999 32164
rect 6025 32108 6081 32164
rect 6107 32114 6148 32164
rect 6148 32114 6163 32164
rect 6189 32114 6200 32164
rect 6200 32114 6214 32164
rect 6214 32114 6245 32164
rect 6107 32108 6163 32114
rect 6189 32108 6245 32114
rect 6271 32108 6327 32164
rect 6353 32108 6409 32164
rect 6435 32108 6491 32164
rect 6517 32108 6573 32164
rect 6599 32108 6655 32164
rect 6681 32114 6702 32164
rect 6702 32114 6737 32164
rect 6763 32114 6768 32164
rect 6768 32114 6819 32164
rect 6681 32108 6737 32114
rect 6763 32108 6819 32114
rect 6845 32108 6901 32164
rect 6927 32108 6983 32164
rect 7009 32108 7065 32164
rect 7091 32108 7147 32164
rect 7173 32108 7229 32164
rect 7255 32114 7256 32164
rect 7256 32114 7308 32164
rect 7308 32114 7311 32164
rect 7337 32114 7374 32164
rect 7374 32114 7393 32164
rect 7255 32108 7311 32114
rect 7337 32108 7393 32114
rect 7419 32108 7475 32164
rect 7501 32108 7557 32164
rect 7583 32108 7639 32164
rect 7665 32108 7721 32164
rect 7747 32108 7803 32164
rect 7829 32114 7862 32164
rect 7862 32114 7876 32164
rect 7876 32114 7885 32164
rect 7911 32114 7928 32164
rect 7928 32114 7967 32164
rect 7829 32108 7885 32114
rect 7911 32108 7967 32114
rect 7993 32116 8047 32164
rect 8047 32116 8049 32164
rect 8075 32116 8099 32164
rect 8099 32116 8131 32164
rect 7993 32108 8049 32116
rect 8075 32108 8131 32116
rect 8157 32116 8169 32164
rect 8169 32116 8213 32164
rect 8157 32108 8213 32116
rect 2733 31931 2789 31987
rect 2814 31931 2870 31987
rect 2895 31931 2951 31987
rect 2976 31931 3032 31987
rect 3057 31982 3113 31987
rect 3138 31982 3194 31987
rect 3057 31931 3101 31982
rect 3101 31931 3113 31982
rect 3138 31931 3153 31982
rect 3153 31931 3167 31982
rect 3167 31931 3194 31982
rect 3219 31931 3275 31987
rect 3300 31931 3356 31987
rect 3381 31931 3437 31987
rect 3462 31931 3518 31987
rect 3543 31931 3599 31987
rect 3624 31982 3680 31987
rect 3705 31982 3761 31987
rect 3624 31931 3655 31982
rect 3655 31931 3680 31982
rect 3705 31931 3707 31982
rect 3707 31931 3721 31982
rect 3721 31931 3761 31982
rect 3786 31931 3842 31987
rect 3867 31931 3923 31987
rect 3948 31931 4004 31987
rect 4029 31931 4085 31987
rect 4110 31931 4166 31987
rect 4191 31982 4247 31987
rect 4272 31982 4328 31987
rect 4191 31931 4209 31982
rect 4209 31931 4247 31982
rect 4272 31931 4275 31982
rect 4275 31931 4327 31982
rect 4327 31931 4328 31982
rect 4353 31931 4409 31987
rect 4434 31931 4490 31987
rect 4515 31931 4571 31987
rect 4596 31931 4652 31987
rect 4677 31931 4733 31987
rect 4758 31982 4814 31987
rect 4839 31982 4895 31987
rect 4758 31931 4763 31982
rect 4763 31931 4814 31982
rect 4839 31931 4881 31982
rect 4881 31931 4895 31982
rect 4920 31931 4976 31987
rect 5001 31931 5057 31987
rect 5082 31931 5138 31987
rect 2733 31851 2789 31907
rect 2814 31851 2870 31907
rect 2895 31851 2951 31907
rect 2976 31851 3032 31907
rect 3057 31861 3101 31907
rect 3101 31861 3113 31907
rect 3138 31861 3153 31907
rect 3153 31861 3167 31907
rect 3167 31861 3194 31907
rect 3057 31851 3113 31861
rect 3138 31851 3194 31861
rect 3219 31851 3275 31907
rect 3300 31851 3356 31907
rect 3381 31851 3437 31907
rect 3462 31851 3518 31907
rect 3543 31851 3599 31907
rect 3624 31861 3655 31907
rect 3655 31861 3680 31907
rect 3705 31861 3707 31907
rect 3707 31861 3721 31907
rect 3721 31861 3761 31907
rect 3624 31851 3680 31861
rect 3705 31851 3761 31861
rect 3786 31851 3842 31907
rect 3867 31851 3923 31907
rect 3948 31851 4004 31907
rect 4029 31851 4085 31907
rect 4110 31851 4166 31907
rect 4191 31861 4209 31907
rect 4209 31861 4247 31907
rect 4272 31861 4275 31907
rect 4275 31861 4327 31907
rect 4327 31861 4328 31907
rect 4191 31851 4247 31861
rect 4272 31851 4328 31861
rect 4353 31851 4409 31907
rect 4434 31851 4490 31907
rect 4515 31851 4571 31907
rect 4596 31851 4652 31907
rect 4677 31851 4733 31907
rect 4758 31861 4763 31907
rect 4763 31861 4814 31907
rect 4839 31861 4881 31907
rect 4881 31861 4895 31907
rect 4758 31851 4814 31861
rect 4839 31851 4895 31861
rect 4920 31851 4976 31907
rect 5001 31851 5057 31907
rect 5082 31851 5138 31907
rect 2733 31771 2789 31827
rect 2814 31771 2870 31827
rect 2895 31771 2951 31827
rect 2976 31771 3032 31827
rect 3057 31792 3101 31827
rect 3101 31792 3113 31827
rect 3138 31792 3153 31827
rect 3153 31792 3167 31827
rect 3167 31792 3194 31827
rect 3057 31775 3113 31792
rect 3138 31775 3194 31792
rect 3057 31771 3101 31775
rect 3101 31771 3113 31775
rect 3138 31771 3153 31775
rect 3153 31771 3167 31775
rect 3167 31771 3194 31775
rect 3219 31771 3275 31827
rect 3300 31771 3356 31827
rect 3381 31771 3437 31827
rect 3462 31771 3518 31827
rect 3543 31771 3599 31827
rect 3624 31792 3655 31827
rect 3655 31792 3680 31827
rect 3705 31792 3707 31827
rect 3707 31792 3721 31827
rect 3721 31792 3761 31827
rect 3624 31775 3680 31792
rect 3705 31775 3761 31792
rect 3624 31771 3655 31775
rect 3655 31771 3680 31775
rect 3705 31771 3707 31775
rect 3707 31771 3721 31775
rect 3721 31771 3761 31775
rect 3786 31771 3842 31827
rect 3867 31771 3923 31827
rect 3948 31771 4004 31827
rect 4029 31771 4085 31827
rect 4110 31771 4166 31827
rect 4191 31792 4209 31827
rect 4209 31792 4247 31827
rect 4272 31792 4275 31827
rect 4275 31792 4327 31827
rect 4327 31792 4328 31827
rect 4191 31775 4247 31792
rect 4272 31775 4328 31792
rect 4191 31771 4209 31775
rect 4209 31771 4247 31775
rect 4272 31771 4275 31775
rect 4275 31771 4327 31775
rect 4327 31771 4328 31775
rect 4353 31771 4409 31827
rect 4434 31771 4490 31827
rect 4515 31771 4571 31827
rect 4596 31771 4652 31827
rect 4677 31771 4733 31827
rect 4758 31792 4763 31827
rect 4763 31792 4814 31827
rect 4839 31792 4881 31827
rect 4881 31792 4895 31827
rect 4758 31775 4814 31792
rect 4839 31775 4895 31792
rect 4758 31771 4763 31775
rect 4763 31771 4814 31775
rect 2733 31691 2789 31747
rect 2814 31691 2870 31747
rect 2895 31691 2951 31747
rect 2976 31691 3032 31747
rect 3057 31723 3101 31747
rect 3101 31723 3113 31747
rect 3138 31723 3153 31747
rect 3153 31723 3167 31747
rect 3167 31723 3194 31747
rect 3057 31706 3113 31723
rect 3138 31706 3194 31723
rect 3057 31691 3101 31706
rect 3101 31691 3113 31706
rect 3138 31691 3153 31706
rect 3153 31691 3167 31706
rect 3167 31691 3194 31706
rect 3219 31691 3275 31747
rect 3300 31691 3356 31747
rect 3381 31691 3437 31747
rect 3462 31691 3518 31747
rect 3543 31691 3599 31747
rect 3624 31723 3655 31747
rect 3655 31723 3680 31747
rect 3705 31723 3707 31747
rect 3707 31723 3721 31747
rect 3721 31723 3761 31747
rect 3624 31706 3680 31723
rect 3705 31706 3761 31723
rect 3624 31691 3655 31706
rect 3655 31691 3680 31706
rect 3705 31691 3707 31706
rect 3707 31691 3721 31706
rect 3721 31691 3761 31706
rect 3786 31691 3842 31747
rect 3867 31691 3923 31747
rect 3948 31691 4004 31747
rect 4029 31691 4085 31747
rect 4110 31691 4166 31747
rect 4191 31723 4209 31747
rect 4209 31723 4247 31747
rect 4272 31723 4275 31747
rect 4275 31723 4327 31747
rect 4327 31723 4328 31747
rect 4191 31706 4247 31723
rect 4272 31706 4328 31723
rect 4191 31691 4209 31706
rect 4209 31691 4247 31706
rect 4272 31691 4275 31706
rect 4275 31691 4327 31706
rect 4327 31691 4328 31706
rect 4353 31691 4409 31747
rect 4434 31691 4490 31747
rect 4515 31691 4571 31747
rect 4596 31691 4652 31747
rect 4677 31691 4733 31747
rect 4758 31723 4763 31747
rect 4763 31723 4814 31747
rect 4839 31771 4881 31775
rect 4881 31771 4895 31775
rect 4920 31771 4976 31827
rect 5001 31771 5057 31827
rect 5082 31771 5138 31827
rect 4839 31723 4881 31747
rect 4881 31723 4895 31747
rect 4758 31706 4814 31723
rect 4839 31706 4895 31723
rect 4758 31691 4763 31706
rect 4763 31691 4814 31706
rect 2733 31611 2789 31667
rect 2814 31611 2870 31667
rect 2895 31611 2951 31667
rect 2976 31611 3032 31667
rect 3057 31654 3101 31667
rect 3101 31654 3113 31667
rect 3138 31654 3153 31667
rect 3153 31654 3167 31667
rect 3167 31654 3194 31667
rect 3057 31636 3113 31654
rect 3138 31636 3194 31654
rect 3057 31611 3101 31636
rect 3101 31611 3113 31636
rect 3138 31611 3153 31636
rect 3153 31611 3167 31636
rect 3167 31611 3194 31636
rect 3219 31611 3275 31667
rect 3300 31611 3356 31667
rect 3381 31611 3437 31667
rect 3462 31611 3518 31667
rect 3543 31611 3599 31667
rect 3624 31654 3655 31667
rect 3655 31654 3680 31667
rect 3705 31654 3707 31667
rect 3707 31654 3721 31667
rect 3721 31654 3761 31667
rect 3624 31636 3680 31654
rect 3705 31636 3761 31654
rect 3624 31611 3655 31636
rect 3655 31611 3680 31636
rect 3705 31611 3707 31636
rect 3707 31611 3721 31636
rect 3721 31611 3761 31636
rect 3786 31611 3842 31667
rect 3867 31611 3923 31667
rect 3948 31611 4004 31667
rect 4029 31611 4085 31667
rect 4110 31611 4166 31667
rect 4191 31654 4209 31667
rect 4209 31654 4247 31667
rect 4272 31654 4275 31667
rect 4275 31654 4327 31667
rect 4327 31654 4328 31667
rect 4191 31636 4247 31654
rect 4272 31636 4328 31654
rect 4191 31611 4209 31636
rect 4209 31611 4247 31636
rect 4272 31611 4275 31636
rect 4275 31611 4327 31636
rect 4327 31611 4328 31636
rect 4353 31611 4409 31667
rect 4434 31611 4490 31667
rect 4515 31611 4571 31667
rect 4596 31611 4652 31667
rect 4677 31611 4733 31667
rect 4758 31654 4763 31667
rect 4763 31654 4814 31667
rect 4839 31691 4881 31706
rect 4881 31691 4895 31706
rect 4920 31691 4976 31747
rect 5001 31691 5057 31747
rect 5082 31691 5138 31747
rect 4839 31654 4881 31667
rect 4881 31654 4895 31667
rect 4758 31636 4814 31654
rect 4839 31636 4895 31654
rect 4758 31611 4763 31636
rect 4763 31611 4814 31636
rect 2733 31531 2789 31587
rect 2814 31531 2870 31587
rect 2895 31531 2951 31587
rect 2976 31531 3032 31587
rect 3057 31584 3101 31587
rect 3101 31584 3113 31587
rect 3138 31584 3153 31587
rect 3153 31584 3167 31587
rect 3167 31584 3194 31587
rect 3057 31566 3113 31584
rect 3138 31566 3194 31584
rect 3057 31531 3101 31566
rect 3101 31531 3113 31566
rect 3138 31531 3153 31566
rect 3153 31531 3167 31566
rect 3167 31531 3194 31566
rect 3219 31531 3275 31587
rect 3300 31531 3356 31587
rect 3381 31531 3437 31587
rect 3462 31531 3518 31587
rect 3543 31531 3599 31587
rect 3624 31584 3655 31587
rect 3655 31584 3680 31587
rect 3705 31584 3707 31587
rect 3707 31584 3721 31587
rect 3721 31584 3761 31587
rect 3624 31566 3680 31584
rect 3705 31566 3761 31584
rect 3624 31531 3655 31566
rect 3655 31531 3680 31566
rect 3705 31531 3707 31566
rect 3707 31531 3721 31566
rect 3721 31531 3761 31566
rect 3786 31531 3842 31587
rect 3867 31531 3923 31587
rect 3948 31531 4004 31587
rect 4029 31531 4085 31587
rect 4110 31531 4166 31587
rect 4191 31584 4209 31587
rect 4209 31584 4247 31587
rect 4272 31584 4275 31587
rect 4275 31584 4327 31587
rect 4327 31584 4328 31587
rect 4191 31566 4247 31584
rect 4272 31566 4328 31584
rect 4191 31531 4209 31566
rect 4209 31531 4247 31566
rect 4272 31531 4275 31566
rect 4275 31531 4327 31566
rect 4327 31531 4328 31566
rect 4353 31531 4409 31587
rect 4434 31531 4490 31587
rect 4515 31531 4571 31587
rect 4596 31531 4652 31587
rect 4677 31531 4733 31587
rect 4758 31584 4763 31587
rect 4763 31584 4814 31587
rect 4839 31611 4881 31636
rect 4881 31611 4895 31636
rect 4920 31611 4976 31667
rect 5001 31611 5057 31667
rect 5082 31611 5138 31667
rect 4839 31584 4881 31587
rect 4881 31584 4895 31587
rect 4758 31566 4814 31584
rect 4839 31566 4895 31584
rect 4758 31531 4763 31566
rect 4763 31531 4814 31566
rect 4839 31531 4881 31566
rect 4881 31531 4895 31566
rect 4920 31531 4976 31587
rect 5001 31531 5057 31587
rect 5082 31531 5138 31587
rect 2733 31451 2789 31507
rect 2814 31451 2870 31507
rect 2895 31451 2951 31507
rect 2976 31451 3032 31507
rect 3057 31496 3113 31507
rect 3138 31496 3194 31507
rect 3057 31451 3101 31496
rect 3101 31451 3113 31496
rect 3138 31451 3153 31496
rect 3153 31451 3167 31496
rect 3167 31451 3194 31496
rect 3219 31451 3275 31507
rect 3300 31451 3356 31507
rect 3381 31451 3437 31507
rect 3462 31451 3518 31507
rect 3543 31451 3599 31507
rect 3624 31496 3680 31507
rect 3705 31496 3761 31507
rect 3624 31451 3655 31496
rect 3655 31451 3680 31496
rect 3705 31451 3707 31496
rect 3707 31451 3721 31496
rect 3721 31451 3761 31496
rect 3786 31451 3842 31507
rect 3867 31451 3923 31507
rect 3948 31451 4004 31507
rect 4029 31451 4085 31507
rect 4110 31451 4166 31507
rect 4191 31496 4247 31507
rect 4272 31496 4328 31507
rect 4191 31451 4209 31496
rect 4209 31451 4247 31496
rect 4272 31451 4275 31496
rect 4275 31451 4327 31496
rect 4327 31451 4328 31496
rect 4353 31451 4409 31507
rect 4434 31451 4490 31507
rect 4515 31451 4571 31507
rect 4596 31451 4652 31507
rect 4677 31451 4733 31507
rect 4758 31496 4814 31507
rect 4839 31496 4895 31507
rect 4758 31451 4763 31496
rect 4763 31451 4814 31496
rect 4839 31451 4881 31496
rect 4881 31451 4895 31496
rect 4920 31451 4976 31507
rect 5001 31451 5057 31507
rect 5082 31451 5138 31507
rect 2733 31371 2789 31427
rect 2814 31371 2870 31427
rect 2895 31371 2951 31427
rect 2976 31371 3032 31427
rect 3057 31426 3113 31427
rect 3138 31426 3194 31427
rect 3057 31374 3101 31426
rect 3101 31374 3113 31426
rect 3138 31374 3153 31426
rect 3153 31374 3167 31426
rect 3167 31374 3194 31426
rect 3057 31371 3113 31374
rect 3138 31371 3194 31374
rect 3219 31371 3275 31427
rect 3300 31371 3356 31427
rect 3381 31371 3437 31427
rect 3462 31371 3518 31427
rect 3543 31371 3599 31427
rect 3624 31426 3680 31427
rect 3705 31426 3761 31427
rect 3624 31374 3655 31426
rect 3655 31374 3680 31426
rect 3705 31374 3707 31426
rect 3707 31374 3721 31426
rect 3721 31374 3761 31426
rect 3624 31371 3680 31374
rect 3705 31371 3761 31374
rect 3786 31371 3842 31427
rect 3867 31371 3923 31427
rect 3948 31371 4004 31427
rect 4029 31371 4085 31427
rect 4110 31371 4166 31427
rect 4191 31426 4247 31427
rect 4272 31426 4328 31427
rect 4191 31374 4209 31426
rect 4209 31374 4247 31426
rect 4272 31374 4275 31426
rect 4275 31374 4327 31426
rect 4327 31374 4328 31426
rect 4191 31371 4247 31374
rect 4272 31371 4328 31374
rect 4353 31371 4409 31427
rect 4434 31371 4490 31427
rect 4515 31371 4571 31427
rect 4596 31371 4652 31427
rect 4677 31371 4733 31427
rect 4758 31426 4814 31427
rect 4839 31426 4895 31427
rect 4758 31374 4763 31426
rect 4763 31374 4814 31426
rect 4839 31374 4881 31426
rect 4881 31374 4895 31426
rect 4758 31371 4814 31374
rect 4839 31371 4895 31374
rect 4920 31371 4976 31427
rect 5001 31371 5057 31427
rect 5082 31371 5138 31427
rect 5163 31371 5299 31987
rect 5613 30720 5669 30724
rect 5696 30720 5752 30724
rect 5613 30668 5646 30720
rect 5646 30668 5660 30720
rect 5660 30668 5669 30720
rect 5696 30668 5712 30720
rect 5712 30668 5752 30720
rect 5779 30668 5835 30724
rect 5861 30668 5917 30724
rect 5943 30668 5999 30724
rect 6025 30668 6081 30724
rect 6107 30720 6163 30724
rect 6189 30720 6245 30724
rect 6107 30668 6148 30720
rect 6148 30668 6163 30720
rect 6189 30668 6200 30720
rect 6200 30668 6214 30720
rect 6214 30668 6245 30720
rect 6271 30668 6327 30724
rect 6353 30668 6409 30724
rect 6435 30668 6491 30724
rect 6517 30668 6573 30724
rect 6599 30668 6655 30724
rect 6681 30720 6737 30724
rect 6763 30720 6819 30724
rect 6681 30668 6702 30720
rect 6702 30668 6737 30720
rect 6763 30668 6768 30720
rect 6768 30668 6819 30720
rect 6845 30668 6901 30724
rect 6927 30668 6983 30724
rect 7009 30668 7065 30724
rect 7091 30668 7147 30724
rect 7173 30668 7229 30724
rect 7255 30720 7311 30724
rect 7337 30720 7393 30724
rect 7255 30668 7256 30720
rect 7256 30668 7308 30720
rect 7308 30668 7311 30720
rect 7337 30668 7374 30720
rect 7374 30668 7393 30720
rect 7419 30668 7475 30724
rect 7501 30668 7557 30724
rect 7583 30668 7639 30724
rect 7665 30668 7721 30724
rect 7747 30668 7803 30724
rect 7829 30720 7885 30724
rect 7911 30720 7967 30724
rect 7829 30668 7862 30720
rect 7862 30668 7876 30720
rect 7876 30668 7885 30720
rect 7911 30668 7928 30720
rect 7928 30668 7967 30720
rect 7993 30672 8047 30724
rect 8047 30672 8049 30724
rect 8075 30672 8099 30724
rect 8099 30672 8131 30724
rect 7993 30668 8049 30672
rect 8075 30668 8131 30672
rect 8157 30672 8169 30724
rect 8169 30672 8213 30724
rect 8157 30668 8213 30672
rect 5613 30599 5646 30644
rect 5646 30599 5660 30644
rect 5660 30599 5669 30644
rect 5696 30599 5712 30644
rect 5712 30599 5752 30644
rect 5613 30588 5669 30599
rect 5696 30588 5752 30599
rect 5779 30588 5835 30644
rect 5861 30588 5917 30644
rect 5943 30588 5999 30644
rect 6025 30588 6081 30644
rect 6107 30599 6148 30644
rect 6148 30599 6163 30644
rect 6189 30599 6200 30644
rect 6200 30599 6214 30644
rect 6214 30599 6245 30644
rect 6107 30588 6163 30599
rect 6189 30588 6245 30599
rect 6271 30588 6327 30644
rect 6353 30588 6409 30644
rect 6435 30588 6491 30644
rect 6517 30588 6573 30644
rect 6599 30588 6655 30644
rect 6681 30599 6702 30644
rect 6702 30599 6737 30644
rect 6763 30599 6768 30644
rect 6768 30599 6819 30644
rect 6681 30588 6737 30599
rect 6763 30588 6819 30599
rect 6845 30588 6901 30644
rect 6927 30588 6983 30644
rect 7009 30588 7065 30644
rect 7091 30588 7147 30644
rect 7173 30588 7229 30644
rect 7255 30599 7256 30644
rect 7256 30599 7308 30644
rect 7308 30599 7311 30644
rect 7337 30599 7374 30644
rect 7374 30599 7393 30644
rect 7255 30588 7311 30599
rect 7337 30588 7393 30599
rect 7419 30588 7475 30644
rect 7501 30588 7557 30644
rect 7583 30588 7639 30644
rect 7665 30588 7721 30644
rect 7747 30588 7803 30644
rect 7829 30599 7862 30644
rect 7862 30599 7876 30644
rect 7876 30599 7885 30644
rect 7911 30599 7928 30644
rect 7928 30599 7967 30644
rect 7829 30588 7885 30599
rect 7911 30588 7967 30599
rect 7993 30603 8047 30644
rect 8047 30603 8049 30644
rect 8075 30603 8099 30644
rect 8099 30603 8131 30644
rect 7993 30588 8049 30603
rect 8075 30588 8131 30603
rect 8157 30603 8169 30644
rect 8169 30603 8213 30644
rect 8157 30588 8213 30603
rect 5613 30530 5646 30564
rect 5646 30530 5660 30564
rect 5660 30530 5669 30564
rect 5696 30530 5712 30564
rect 5712 30530 5752 30564
rect 5613 30513 5669 30530
rect 5696 30513 5752 30530
rect 5613 30508 5646 30513
rect 5646 30508 5660 30513
rect 5660 30508 5669 30513
rect 5696 30508 5712 30513
rect 5712 30508 5752 30513
rect 5779 30508 5835 30564
rect 5861 30508 5917 30564
rect 5943 30508 5999 30564
rect 6025 30508 6081 30564
rect 6107 30530 6148 30564
rect 6148 30530 6163 30564
rect 6189 30530 6200 30564
rect 6200 30530 6214 30564
rect 6214 30530 6245 30564
rect 6107 30513 6163 30530
rect 6189 30513 6245 30530
rect 6107 30508 6148 30513
rect 6148 30508 6163 30513
rect 6189 30508 6200 30513
rect 6200 30508 6214 30513
rect 6214 30508 6245 30513
rect 6271 30508 6327 30564
rect 6353 30508 6409 30564
rect 6435 30508 6491 30564
rect 6517 30508 6573 30564
rect 6599 30508 6655 30564
rect 6681 30530 6702 30564
rect 6702 30530 6737 30564
rect 6763 30530 6768 30564
rect 6768 30530 6819 30564
rect 6681 30513 6737 30530
rect 6763 30513 6819 30530
rect 6681 30508 6702 30513
rect 6702 30508 6737 30513
rect 6763 30508 6768 30513
rect 6768 30508 6819 30513
rect 6845 30508 6901 30564
rect 6927 30508 6983 30564
rect 7009 30508 7065 30564
rect 7091 30508 7147 30564
rect 7173 30508 7229 30564
rect 7255 30530 7256 30564
rect 7256 30530 7308 30564
rect 7308 30530 7311 30564
rect 7337 30530 7374 30564
rect 7374 30530 7393 30564
rect 7255 30513 7311 30530
rect 7337 30513 7393 30530
rect 7255 30508 7256 30513
rect 7256 30508 7308 30513
rect 7308 30508 7311 30513
rect 7337 30508 7374 30513
rect 7374 30508 7393 30513
rect 7419 30508 7475 30564
rect 7501 30508 7557 30564
rect 7583 30508 7639 30564
rect 7665 30508 7721 30564
rect 7747 30508 7803 30564
rect 7829 30530 7862 30564
rect 7862 30530 7876 30564
rect 7876 30530 7885 30564
rect 7911 30530 7928 30564
rect 7928 30530 7967 30564
rect 7829 30513 7885 30530
rect 7911 30513 7967 30530
rect 7829 30508 7862 30513
rect 7862 30508 7876 30513
rect 7876 30508 7885 30513
rect 7911 30508 7928 30513
rect 7928 30508 7967 30513
rect 7993 30534 8047 30564
rect 8047 30534 8049 30564
rect 8075 30534 8099 30564
rect 8099 30534 8131 30564
rect 7993 30517 8049 30534
rect 8075 30517 8131 30534
rect 7993 30508 8047 30517
rect 8047 30508 8049 30517
rect 8075 30508 8099 30517
rect 8099 30508 8131 30517
rect 8157 30534 8169 30564
rect 8169 30534 8213 30564
rect 8157 30517 8213 30534
rect 8157 30508 8169 30517
rect 8169 30508 8213 30517
rect 5613 30461 5646 30484
rect 5646 30461 5660 30484
rect 5660 30461 5669 30484
rect 5696 30461 5712 30484
rect 5712 30461 5752 30484
rect 5613 30444 5669 30461
rect 5696 30444 5752 30461
rect 5613 30428 5646 30444
rect 5646 30428 5660 30444
rect 5660 30428 5669 30444
rect 5696 30428 5712 30444
rect 5712 30428 5752 30444
rect 5779 30428 5835 30484
rect 5861 30428 5917 30484
rect 5943 30428 5999 30484
rect 6025 30428 6081 30484
rect 6107 30461 6148 30484
rect 6148 30461 6163 30484
rect 6189 30461 6200 30484
rect 6200 30461 6214 30484
rect 6214 30461 6245 30484
rect 6107 30444 6163 30461
rect 6189 30444 6245 30461
rect 6107 30428 6148 30444
rect 6148 30428 6163 30444
rect 6189 30428 6200 30444
rect 6200 30428 6214 30444
rect 6214 30428 6245 30444
rect 6271 30428 6327 30484
rect 6353 30428 6409 30484
rect 6435 30428 6491 30484
rect 6517 30428 6573 30484
rect 6599 30428 6655 30484
rect 6681 30461 6702 30484
rect 6702 30461 6737 30484
rect 6763 30461 6768 30484
rect 6768 30461 6819 30484
rect 6681 30444 6737 30461
rect 6763 30444 6819 30461
rect 6681 30428 6702 30444
rect 6702 30428 6737 30444
rect 6763 30428 6768 30444
rect 6768 30428 6819 30444
rect 6845 30428 6901 30484
rect 6927 30428 6983 30484
rect 7009 30428 7065 30484
rect 7091 30428 7147 30484
rect 7173 30428 7229 30484
rect 7255 30461 7256 30484
rect 7256 30461 7308 30484
rect 7308 30461 7311 30484
rect 7337 30461 7374 30484
rect 7374 30461 7393 30484
rect 7255 30444 7311 30461
rect 7337 30444 7393 30461
rect 7255 30428 7256 30444
rect 7256 30428 7308 30444
rect 7308 30428 7311 30444
rect 7337 30428 7374 30444
rect 7374 30428 7393 30444
rect 7419 30428 7475 30484
rect 7501 30428 7557 30484
rect 7583 30428 7639 30484
rect 7665 30428 7721 30484
rect 7747 30428 7803 30484
rect 7829 30461 7862 30484
rect 7862 30461 7876 30484
rect 7876 30461 7885 30484
rect 7911 30461 7928 30484
rect 7928 30461 7967 30484
rect 7829 30444 7885 30461
rect 7911 30444 7967 30461
rect 7829 30428 7862 30444
rect 7862 30428 7876 30444
rect 7876 30428 7885 30444
rect 7911 30428 7928 30444
rect 7928 30428 7967 30444
rect 7993 30465 8047 30484
rect 8047 30465 8049 30484
rect 8075 30465 8099 30484
rect 8099 30465 8131 30484
rect 7993 30448 8049 30465
rect 8075 30448 8131 30465
rect 7993 30428 8047 30448
rect 8047 30428 8049 30448
rect 8075 30428 8099 30448
rect 8099 30428 8131 30448
rect 8157 30465 8169 30484
rect 8169 30465 8213 30484
rect 8157 30448 8213 30465
rect 8157 30428 8169 30448
rect 8169 30428 8213 30448
rect 5613 30392 5646 30404
rect 5646 30392 5660 30404
rect 5660 30392 5669 30404
rect 5696 30392 5712 30404
rect 5712 30392 5752 30404
rect 5613 30375 5669 30392
rect 5696 30375 5752 30392
rect 5613 30348 5646 30375
rect 5646 30348 5660 30375
rect 5660 30348 5669 30375
rect 5696 30348 5712 30375
rect 5712 30348 5752 30375
rect 5779 30348 5835 30404
rect 5861 30348 5917 30404
rect 5943 30348 5999 30404
rect 6025 30348 6081 30404
rect 6107 30392 6148 30404
rect 6148 30392 6163 30404
rect 6189 30392 6200 30404
rect 6200 30392 6214 30404
rect 6214 30392 6245 30404
rect 6107 30375 6163 30392
rect 6189 30375 6245 30392
rect 6107 30348 6148 30375
rect 6148 30348 6163 30375
rect 6189 30348 6200 30375
rect 6200 30348 6214 30375
rect 6214 30348 6245 30375
rect 6271 30348 6327 30404
rect 6353 30348 6409 30404
rect 6435 30348 6491 30404
rect 6517 30348 6573 30404
rect 6599 30348 6655 30404
rect 6681 30392 6702 30404
rect 6702 30392 6737 30404
rect 6763 30392 6768 30404
rect 6768 30392 6819 30404
rect 6681 30375 6737 30392
rect 6763 30375 6819 30392
rect 6681 30348 6702 30375
rect 6702 30348 6737 30375
rect 6763 30348 6768 30375
rect 6768 30348 6819 30375
rect 6845 30348 6901 30404
rect 6927 30348 6983 30404
rect 7009 30348 7065 30404
rect 7091 30348 7147 30404
rect 7173 30348 7229 30404
rect 7255 30392 7256 30404
rect 7256 30392 7308 30404
rect 7308 30392 7311 30404
rect 7337 30392 7374 30404
rect 7374 30392 7393 30404
rect 7255 30375 7311 30392
rect 7337 30375 7393 30392
rect 7255 30348 7256 30375
rect 7256 30348 7308 30375
rect 7308 30348 7311 30375
rect 7337 30348 7374 30375
rect 7374 30348 7393 30375
rect 7419 30348 7475 30404
rect 7501 30348 7557 30404
rect 7583 30348 7639 30404
rect 7665 30348 7721 30404
rect 7747 30348 7803 30404
rect 7829 30392 7862 30404
rect 7862 30392 7876 30404
rect 7876 30392 7885 30404
rect 7911 30392 7928 30404
rect 7928 30392 7967 30404
rect 7829 30375 7885 30392
rect 7911 30375 7967 30392
rect 7829 30348 7862 30375
rect 7862 30348 7876 30375
rect 7876 30348 7885 30375
rect 7911 30348 7928 30375
rect 7928 30348 7967 30375
rect 7993 30396 8047 30404
rect 8047 30396 8049 30404
rect 8075 30396 8099 30404
rect 8099 30396 8131 30404
rect 7993 30378 8049 30396
rect 8075 30378 8131 30396
rect 7993 30348 8047 30378
rect 8047 30348 8049 30378
rect 8075 30348 8099 30378
rect 8099 30348 8131 30378
rect 8157 30396 8169 30404
rect 8169 30396 8213 30404
rect 8157 30378 8213 30396
rect 8157 30348 8169 30378
rect 8169 30348 8213 30378
rect 5613 30323 5646 30324
rect 5646 30323 5660 30324
rect 5660 30323 5669 30324
rect 5696 30323 5712 30324
rect 5712 30323 5752 30324
rect 5613 30306 5669 30323
rect 5696 30306 5752 30323
rect 5613 30268 5646 30306
rect 5646 30268 5660 30306
rect 5660 30268 5669 30306
rect 5696 30268 5712 30306
rect 5712 30268 5752 30306
rect 5779 30268 5835 30324
rect 5861 30268 5917 30324
rect 5943 30268 5999 30324
rect 6025 30268 6081 30324
rect 6107 30323 6148 30324
rect 6148 30323 6163 30324
rect 6189 30323 6200 30324
rect 6200 30323 6214 30324
rect 6214 30323 6245 30324
rect 6107 30306 6163 30323
rect 6189 30306 6245 30323
rect 6107 30268 6148 30306
rect 6148 30268 6163 30306
rect 6189 30268 6200 30306
rect 6200 30268 6214 30306
rect 6214 30268 6245 30306
rect 6271 30268 6327 30324
rect 6353 30268 6409 30324
rect 6435 30268 6491 30324
rect 6517 30268 6573 30324
rect 6599 30268 6655 30324
rect 6681 30323 6702 30324
rect 6702 30323 6737 30324
rect 6763 30323 6768 30324
rect 6768 30323 6819 30324
rect 6681 30306 6737 30323
rect 6763 30306 6819 30323
rect 6681 30268 6702 30306
rect 6702 30268 6737 30306
rect 6763 30268 6768 30306
rect 6768 30268 6819 30306
rect 6845 30268 6901 30324
rect 6927 30268 6983 30324
rect 7009 30268 7065 30324
rect 7091 30268 7147 30324
rect 7173 30268 7229 30324
rect 7255 30323 7256 30324
rect 7256 30323 7308 30324
rect 7308 30323 7311 30324
rect 7337 30323 7374 30324
rect 7374 30323 7393 30324
rect 7255 30306 7311 30323
rect 7337 30306 7393 30323
rect 7255 30268 7256 30306
rect 7256 30268 7308 30306
rect 7308 30268 7311 30306
rect 7337 30268 7374 30306
rect 7374 30268 7393 30306
rect 7419 30268 7475 30324
rect 7501 30268 7557 30324
rect 7583 30268 7639 30324
rect 7665 30268 7721 30324
rect 7747 30268 7803 30324
rect 7829 30323 7862 30324
rect 7862 30323 7876 30324
rect 7876 30323 7885 30324
rect 7911 30323 7928 30324
rect 7928 30323 7967 30324
rect 7829 30306 7885 30323
rect 7911 30306 7967 30323
rect 7829 30268 7862 30306
rect 7862 30268 7876 30306
rect 7876 30268 7885 30306
rect 7911 30268 7928 30306
rect 7928 30268 7967 30306
rect 7993 30308 8049 30324
rect 8075 30308 8131 30324
rect 7993 30268 8047 30308
rect 8047 30268 8049 30308
rect 8075 30268 8099 30308
rect 8099 30268 8131 30308
rect 8157 30308 8213 30324
rect 8157 30268 8169 30308
rect 8169 30268 8213 30308
rect 5613 30236 5669 30244
rect 5696 30236 5752 30244
rect 5613 30188 5646 30236
rect 5646 30188 5660 30236
rect 5660 30188 5669 30236
rect 5696 30188 5712 30236
rect 5712 30188 5752 30236
rect 5779 30188 5835 30244
rect 5861 30188 5917 30244
rect 5943 30188 5999 30244
rect 6025 30188 6081 30244
rect 6107 30236 6163 30244
rect 6189 30236 6245 30244
rect 6107 30188 6148 30236
rect 6148 30188 6163 30236
rect 6189 30188 6200 30236
rect 6200 30188 6214 30236
rect 6214 30188 6245 30236
rect 6271 30188 6327 30244
rect 6353 30188 6409 30244
rect 6435 30188 6491 30244
rect 6517 30188 6573 30244
rect 6599 30188 6655 30244
rect 6681 30236 6737 30244
rect 6763 30236 6819 30244
rect 6681 30188 6702 30236
rect 6702 30188 6737 30236
rect 6763 30188 6768 30236
rect 6768 30188 6819 30236
rect 6845 30188 6901 30244
rect 6927 30188 6983 30244
rect 7009 30188 7065 30244
rect 7091 30188 7147 30244
rect 7173 30188 7229 30244
rect 7255 30236 7311 30244
rect 7337 30236 7393 30244
rect 7255 30188 7256 30236
rect 7256 30188 7308 30236
rect 7308 30188 7311 30236
rect 7337 30188 7374 30236
rect 7374 30188 7393 30236
rect 7419 30188 7475 30244
rect 7501 30188 7557 30244
rect 7583 30188 7639 30244
rect 7665 30188 7721 30244
rect 7747 30188 7803 30244
rect 7829 30236 7885 30244
rect 7911 30236 7967 30244
rect 7829 30188 7862 30236
rect 7862 30188 7876 30236
rect 7876 30188 7885 30236
rect 7911 30188 7928 30236
rect 7928 30188 7967 30236
rect 7993 30238 8049 30244
rect 8075 30238 8131 30244
rect 7993 30188 8047 30238
rect 8047 30188 8049 30238
rect 8075 30188 8099 30238
rect 8099 30188 8131 30238
rect 8157 30238 8213 30244
rect 8157 30188 8169 30238
rect 8169 30188 8213 30238
rect 5613 30114 5646 30164
rect 5646 30114 5660 30164
rect 5660 30114 5669 30164
rect 5696 30114 5712 30164
rect 5712 30114 5752 30164
rect 5613 30108 5669 30114
rect 5696 30108 5752 30114
rect 5779 30108 5835 30164
rect 5861 30108 5917 30164
rect 5943 30108 5999 30164
rect 6025 30108 6081 30164
rect 6107 30114 6148 30164
rect 6148 30114 6163 30164
rect 6189 30114 6200 30164
rect 6200 30114 6214 30164
rect 6214 30114 6245 30164
rect 6107 30108 6163 30114
rect 6189 30108 6245 30114
rect 6271 30108 6327 30164
rect 6353 30108 6409 30164
rect 6435 30108 6491 30164
rect 6517 30108 6573 30164
rect 6599 30108 6655 30164
rect 6681 30114 6702 30164
rect 6702 30114 6737 30164
rect 6763 30114 6768 30164
rect 6768 30114 6819 30164
rect 6681 30108 6737 30114
rect 6763 30108 6819 30114
rect 6845 30108 6901 30164
rect 6927 30108 6983 30164
rect 7009 30108 7065 30164
rect 7091 30108 7147 30164
rect 7173 30108 7229 30164
rect 7255 30114 7256 30164
rect 7256 30114 7308 30164
rect 7308 30114 7311 30164
rect 7337 30114 7374 30164
rect 7374 30114 7393 30164
rect 7255 30108 7311 30114
rect 7337 30108 7393 30114
rect 7419 30108 7475 30164
rect 7501 30108 7557 30164
rect 7583 30108 7639 30164
rect 7665 30108 7721 30164
rect 7747 30108 7803 30164
rect 7829 30114 7862 30164
rect 7862 30114 7876 30164
rect 7876 30114 7885 30164
rect 7911 30114 7928 30164
rect 7928 30114 7967 30164
rect 7829 30108 7885 30114
rect 7911 30108 7967 30114
rect 7993 30116 8047 30164
rect 8047 30116 8049 30164
rect 8075 30116 8099 30164
rect 8099 30116 8131 30164
rect 7993 30108 8049 30116
rect 8075 30108 8131 30116
rect 8157 30116 8169 30164
rect 8169 30116 8213 30164
rect 8157 30108 8213 30116
rect 2733 29931 2789 29987
rect 2814 29931 2870 29987
rect 2895 29931 2951 29987
rect 2976 29931 3032 29987
rect 3057 29982 3113 29987
rect 3138 29982 3194 29987
rect 3057 29931 3101 29982
rect 3101 29931 3113 29982
rect 3138 29931 3153 29982
rect 3153 29931 3167 29982
rect 3167 29931 3194 29982
rect 3219 29931 3275 29987
rect 3300 29931 3356 29987
rect 3381 29931 3437 29987
rect 3462 29931 3518 29987
rect 3543 29931 3599 29987
rect 3624 29982 3680 29987
rect 3705 29982 3761 29987
rect 3624 29931 3655 29982
rect 3655 29931 3680 29982
rect 3705 29931 3707 29982
rect 3707 29931 3721 29982
rect 3721 29931 3761 29982
rect 3786 29931 3842 29987
rect 3867 29931 3923 29987
rect 3948 29931 4004 29987
rect 4029 29931 4085 29987
rect 4110 29931 4166 29987
rect 4191 29982 4247 29987
rect 4272 29982 4328 29987
rect 4191 29931 4209 29982
rect 4209 29931 4247 29982
rect 4272 29931 4275 29982
rect 4275 29931 4327 29982
rect 4327 29931 4328 29982
rect 4353 29931 4409 29987
rect 4434 29931 4490 29987
rect 4515 29931 4571 29987
rect 4596 29931 4652 29987
rect 4677 29931 4733 29987
rect 4758 29982 4814 29987
rect 4839 29982 4895 29987
rect 4758 29931 4763 29982
rect 4763 29931 4814 29982
rect 4839 29931 4881 29982
rect 4881 29931 4895 29982
rect 4920 29931 4976 29987
rect 5001 29931 5057 29987
rect 5082 29931 5138 29987
rect 2733 29851 2789 29907
rect 2814 29851 2870 29907
rect 2895 29851 2951 29907
rect 2976 29851 3032 29907
rect 3057 29861 3101 29907
rect 3101 29861 3113 29907
rect 3138 29861 3153 29907
rect 3153 29861 3167 29907
rect 3167 29861 3194 29907
rect 3057 29851 3113 29861
rect 3138 29851 3194 29861
rect 3219 29851 3275 29907
rect 3300 29851 3356 29907
rect 3381 29851 3437 29907
rect 3462 29851 3518 29907
rect 3543 29851 3599 29907
rect 3624 29861 3655 29907
rect 3655 29861 3680 29907
rect 3705 29861 3707 29907
rect 3707 29861 3721 29907
rect 3721 29861 3761 29907
rect 3624 29851 3680 29861
rect 3705 29851 3761 29861
rect 3786 29851 3842 29907
rect 3867 29851 3923 29907
rect 3948 29851 4004 29907
rect 4029 29851 4085 29907
rect 4110 29851 4166 29907
rect 4191 29861 4209 29907
rect 4209 29861 4247 29907
rect 4272 29861 4275 29907
rect 4275 29861 4327 29907
rect 4327 29861 4328 29907
rect 4191 29851 4247 29861
rect 4272 29851 4328 29861
rect 4353 29851 4409 29907
rect 4434 29851 4490 29907
rect 4515 29851 4571 29907
rect 4596 29851 4652 29907
rect 4677 29851 4733 29907
rect 4758 29861 4763 29907
rect 4763 29861 4814 29907
rect 4839 29861 4881 29907
rect 4881 29861 4895 29907
rect 4758 29851 4814 29861
rect 4839 29851 4895 29861
rect 4920 29851 4976 29907
rect 5001 29851 5057 29907
rect 5082 29851 5138 29907
rect 2733 29771 2789 29827
rect 2814 29771 2870 29827
rect 2895 29771 2951 29827
rect 2976 29771 3032 29827
rect 3057 29792 3101 29827
rect 3101 29792 3113 29827
rect 3138 29792 3153 29827
rect 3153 29792 3167 29827
rect 3167 29792 3194 29827
rect 3057 29775 3113 29792
rect 3138 29775 3194 29792
rect 3057 29771 3101 29775
rect 3101 29771 3113 29775
rect 3138 29771 3153 29775
rect 3153 29771 3167 29775
rect 3167 29771 3194 29775
rect 3219 29771 3275 29827
rect 3300 29771 3356 29827
rect 3381 29771 3437 29827
rect 3462 29771 3518 29827
rect 3543 29771 3599 29827
rect 3624 29792 3655 29827
rect 3655 29792 3680 29827
rect 3705 29792 3707 29827
rect 3707 29792 3721 29827
rect 3721 29792 3761 29827
rect 3624 29775 3680 29792
rect 3705 29775 3761 29792
rect 3624 29771 3655 29775
rect 3655 29771 3680 29775
rect 3705 29771 3707 29775
rect 3707 29771 3721 29775
rect 3721 29771 3761 29775
rect 3786 29771 3842 29827
rect 3867 29771 3923 29827
rect 3948 29771 4004 29827
rect 4029 29771 4085 29827
rect 4110 29771 4166 29827
rect 4191 29792 4209 29827
rect 4209 29792 4247 29827
rect 4272 29792 4275 29827
rect 4275 29792 4327 29827
rect 4327 29792 4328 29827
rect 4191 29775 4247 29792
rect 4272 29775 4328 29792
rect 4191 29771 4209 29775
rect 4209 29771 4247 29775
rect 4272 29771 4275 29775
rect 4275 29771 4327 29775
rect 4327 29771 4328 29775
rect 4353 29771 4409 29827
rect 4434 29771 4490 29827
rect 4515 29771 4571 29827
rect 4596 29771 4652 29827
rect 4677 29771 4733 29827
rect 4758 29792 4763 29827
rect 4763 29792 4814 29827
rect 4839 29792 4881 29827
rect 4881 29792 4895 29827
rect 4758 29775 4814 29792
rect 4839 29775 4895 29792
rect 4758 29771 4763 29775
rect 4763 29771 4814 29775
rect 2733 29691 2789 29747
rect 2814 29691 2870 29747
rect 2895 29691 2951 29747
rect 2976 29691 3032 29747
rect 3057 29723 3101 29747
rect 3101 29723 3113 29747
rect 3138 29723 3153 29747
rect 3153 29723 3167 29747
rect 3167 29723 3194 29747
rect 3057 29706 3113 29723
rect 3138 29706 3194 29723
rect 3057 29691 3101 29706
rect 3101 29691 3113 29706
rect 3138 29691 3153 29706
rect 3153 29691 3167 29706
rect 3167 29691 3194 29706
rect 3219 29691 3275 29747
rect 3300 29691 3356 29747
rect 3381 29691 3437 29747
rect 3462 29691 3518 29747
rect 3543 29691 3599 29747
rect 3624 29723 3655 29747
rect 3655 29723 3680 29747
rect 3705 29723 3707 29747
rect 3707 29723 3721 29747
rect 3721 29723 3761 29747
rect 3624 29706 3680 29723
rect 3705 29706 3761 29723
rect 3624 29691 3655 29706
rect 3655 29691 3680 29706
rect 3705 29691 3707 29706
rect 3707 29691 3721 29706
rect 3721 29691 3761 29706
rect 3786 29691 3842 29747
rect 3867 29691 3923 29747
rect 3948 29691 4004 29747
rect 4029 29691 4085 29747
rect 4110 29691 4166 29747
rect 4191 29723 4209 29747
rect 4209 29723 4247 29747
rect 4272 29723 4275 29747
rect 4275 29723 4327 29747
rect 4327 29723 4328 29747
rect 4191 29706 4247 29723
rect 4272 29706 4328 29723
rect 4191 29691 4209 29706
rect 4209 29691 4247 29706
rect 4272 29691 4275 29706
rect 4275 29691 4327 29706
rect 4327 29691 4328 29706
rect 4353 29691 4409 29747
rect 4434 29691 4490 29747
rect 4515 29691 4571 29747
rect 4596 29691 4652 29747
rect 4677 29691 4733 29747
rect 4758 29723 4763 29747
rect 4763 29723 4814 29747
rect 4839 29771 4881 29775
rect 4881 29771 4895 29775
rect 4920 29771 4976 29827
rect 5001 29771 5057 29827
rect 5082 29771 5138 29827
rect 4839 29723 4881 29747
rect 4881 29723 4895 29747
rect 4758 29706 4814 29723
rect 4839 29706 4895 29723
rect 4758 29691 4763 29706
rect 4763 29691 4814 29706
rect 2733 29611 2789 29667
rect 2814 29611 2870 29667
rect 2895 29611 2951 29667
rect 2976 29611 3032 29667
rect 3057 29654 3101 29667
rect 3101 29654 3113 29667
rect 3138 29654 3153 29667
rect 3153 29654 3167 29667
rect 3167 29654 3194 29667
rect 3057 29636 3113 29654
rect 3138 29636 3194 29654
rect 3057 29611 3101 29636
rect 3101 29611 3113 29636
rect 3138 29611 3153 29636
rect 3153 29611 3167 29636
rect 3167 29611 3194 29636
rect 3219 29611 3275 29667
rect 3300 29611 3356 29667
rect 3381 29611 3437 29667
rect 3462 29611 3518 29667
rect 3543 29611 3599 29667
rect 3624 29654 3655 29667
rect 3655 29654 3680 29667
rect 3705 29654 3707 29667
rect 3707 29654 3721 29667
rect 3721 29654 3761 29667
rect 3624 29636 3680 29654
rect 3705 29636 3761 29654
rect 3624 29611 3655 29636
rect 3655 29611 3680 29636
rect 3705 29611 3707 29636
rect 3707 29611 3721 29636
rect 3721 29611 3761 29636
rect 3786 29611 3842 29667
rect 3867 29611 3923 29667
rect 3948 29611 4004 29667
rect 4029 29611 4085 29667
rect 4110 29611 4166 29667
rect 4191 29654 4209 29667
rect 4209 29654 4247 29667
rect 4272 29654 4275 29667
rect 4275 29654 4327 29667
rect 4327 29654 4328 29667
rect 4191 29636 4247 29654
rect 4272 29636 4328 29654
rect 4191 29611 4209 29636
rect 4209 29611 4247 29636
rect 4272 29611 4275 29636
rect 4275 29611 4327 29636
rect 4327 29611 4328 29636
rect 4353 29611 4409 29667
rect 4434 29611 4490 29667
rect 4515 29611 4571 29667
rect 4596 29611 4652 29667
rect 4677 29611 4733 29667
rect 4758 29654 4763 29667
rect 4763 29654 4814 29667
rect 4839 29691 4881 29706
rect 4881 29691 4895 29706
rect 4920 29691 4976 29747
rect 5001 29691 5057 29747
rect 5082 29691 5138 29747
rect 4839 29654 4881 29667
rect 4881 29654 4895 29667
rect 4758 29636 4814 29654
rect 4839 29636 4895 29654
rect 4758 29611 4763 29636
rect 4763 29611 4814 29636
rect 2733 29531 2789 29587
rect 2814 29531 2870 29587
rect 2895 29531 2951 29587
rect 2976 29531 3032 29587
rect 3057 29584 3101 29587
rect 3101 29584 3113 29587
rect 3138 29584 3153 29587
rect 3153 29584 3167 29587
rect 3167 29584 3194 29587
rect 3057 29566 3113 29584
rect 3138 29566 3194 29584
rect 3057 29531 3101 29566
rect 3101 29531 3113 29566
rect 3138 29531 3153 29566
rect 3153 29531 3167 29566
rect 3167 29531 3194 29566
rect 3219 29531 3275 29587
rect 3300 29531 3356 29587
rect 3381 29531 3437 29587
rect 3462 29531 3518 29587
rect 3543 29531 3599 29587
rect 3624 29584 3655 29587
rect 3655 29584 3680 29587
rect 3705 29584 3707 29587
rect 3707 29584 3721 29587
rect 3721 29584 3761 29587
rect 3624 29566 3680 29584
rect 3705 29566 3761 29584
rect 3624 29531 3655 29566
rect 3655 29531 3680 29566
rect 3705 29531 3707 29566
rect 3707 29531 3721 29566
rect 3721 29531 3761 29566
rect 3786 29531 3842 29587
rect 3867 29531 3923 29587
rect 3948 29531 4004 29587
rect 4029 29531 4085 29587
rect 4110 29531 4166 29587
rect 4191 29584 4209 29587
rect 4209 29584 4247 29587
rect 4272 29584 4275 29587
rect 4275 29584 4327 29587
rect 4327 29584 4328 29587
rect 4191 29566 4247 29584
rect 4272 29566 4328 29584
rect 4191 29531 4209 29566
rect 4209 29531 4247 29566
rect 4272 29531 4275 29566
rect 4275 29531 4327 29566
rect 4327 29531 4328 29566
rect 4353 29531 4409 29587
rect 4434 29531 4490 29587
rect 4515 29531 4571 29587
rect 4596 29531 4652 29587
rect 4677 29531 4733 29587
rect 4758 29584 4763 29587
rect 4763 29584 4814 29587
rect 4839 29611 4881 29636
rect 4881 29611 4895 29636
rect 4920 29611 4976 29667
rect 5001 29611 5057 29667
rect 5082 29611 5138 29667
rect 4839 29584 4881 29587
rect 4881 29584 4895 29587
rect 4758 29566 4814 29584
rect 4839 29566 4895 29584
rect 4758 29531 4763 29566
rect 4763 29531 4814 29566
rect 4839 29531 4881 29566
rect 4881 29531 4895 29566
rect 4920 29531 4976 29587
rect 5001 29531 5057 29587
rect 5082 29531 5138 29587
rect 2733 29451 2789 29507
rect 2814 29451 2870 29507
rect 2895 29451 2951 29507
rect 2976 29451 3032 29507
rect 3057 29496 3113 29507
rect 3138 29496 3194 29507
rect 3057 29451 3101 29496
rect 3101 29451 3113 29496
rect 3138 29451 3153 29496
rect 3153 29451 3167 29496
rect 3167 29451 3194 29496
rect 3219 29451 3275 29507
rect 3300 29451 3356 29507
rect 3381 29451 3437 29507
rect 3462 29451 3518 29507
rect 3543 29451 3599 29507
rect 3624 29496 3680 29507
rect 3705 29496 3761 29507
rect 3624 29451 3655 29496
rect 3655 29451 3680 29496
rect 3705 29451 3707 29496
rect 3707 29451 3721 29496
rect 3721 29451 3761 29496
rect 3786 29451 3842 29507
rect 3867 29451 3923 29507
rect 3948 29451 4004 29507
rect 4029 29451 4085 29507
rect 4110 29451 4166 29507
rect 4191 29496 4247 29507
rect 4272 29496 4328 29507
rect 4191 29451 4209 29496
rect 4209 29451 4247 29496
rect 4272 29451 4275 29496
rect 4275 29451 4327 29496
rect 4327 29451 4328 29496
rect 4353 29451 4409 29507
rect 4434 29451 4490 29507
rect 4515 29451 4571 29507
rect 4596 29451 4652 29507
rect 4677 29451 4733 29507
rect 4758 29496 4814 29507
rect 4839 29496 4895 29507
rect 4758 29451 4763 29496
rect 4763 29451 4814 29496
rect 4839 29451 4881 29496
rect 4881 29451 4895 29496
rect 4920 29451 4976 29507
rect 5001 29451 5057 29507
rect 5082 29451 5138 29507
rect 2733 29371 2789 29427
rect 2814 29371 2870 29427
rect 2895 29371 2951 29427
rect 2976 29371 3032 29427
rect 3057 29426 3113 29427
rect 3138 29426 3194 29427
rect 3057 29374 3101 29426
rect 3101 29374 3113 29426
rect 3138 29374 3153 29426
rect 3153 29374 3167 29426
rect 3167 29374 3194 29426
rect 3057 29371 3113 29374
rect 3138 29371 3194 29374
rect 3219 29371 3275 29427
rect 3300 29371 3356 29427
rect 3381 29371 3437 29427
rect 3462 29371 3518 29427
rect 3543 29371 3599 29427
rect 3624 29426 3680 29427
rect 3705 29426 3761 29427
rect 3624 29374 3655 29426
rect 3655 29374 3680 29426
rect 3705 29374 3707 29426
rect 3707 29374 3721 29426
rect 3721 29374 3761 29426
rect 3624 29371 3680 29374
rect 3705 29371 3761 29374
rect 3786 29371 3842 29427
rect 3867 29371 3923 29427
rect 3948 29371 4004 29427
rect 4029 29371 4085 29427
rect 4110 29371 4166 29427
rect 4191 29426 4247 29427
rect 4272 29426 4328 29427
rect 4191 29374 4209 29426
rect 4209 29374 4247 29426
rect 4272 29374 4275 29426
rect 4275 29374 4327 29426
rect 4327 29374 4328 29426
rect 4191 29371 4247 29374
rect 4272 29371 4328 29374
rect 4353 29371 4409 29427
rect 4434 29371 4490 29427
rect 4515 29371 4571 29427
rect 4596 29371 4652 29427
rect 4677 29371 4733 29427
rect 4758 29426 4814 29427
rect 4839 29426 4895 29427
rect 4758 29374 4763 29426
rect 4763 29374 4814 29426
rect 4839 29374 4881 29426
rect 4881 29374 4895 29426
rect 4758 29371 4814 29374
rect 4839 29371 4895 29374
rect 4920 29371 4976 29427
rect 5001 29371 5057 29427
rect 5082 29371 5138 29427
rect 5163 29371 5299 29987
rect 5613 28720 5669 28724
rect 5696 28720 5752 28724
rect 5613 28668 5646 28720
rect 5646 28668 5660 28720
rect 5660 28668 5669 28720
rect 5696 28668 5712 28720
rect 5712 28668 5752 28720
rect 5779 28668 5835 28724
rect 5861 28668 5917 28724
rect 5943 28668 5999 28724
rect 6025 28668 6081 28724
rect 6107 28720 6163 28724
rect 6189 28720 6245 28724
rect 6107 28668 6148 28720
rect 6148 28668 6163 28720
rect 6189 28668 6200 28720
rect 6200 28668 6214 28720
rect 6214 28668 6245 28720
rect 6271 28668 6327 28724
rect 6353 28668 6409 28724
rect 6435 28668 6491 28724
rect 6517 28668 6573 28724
rect 6599 28668 6655 28724
rect 6681 28720 6737 28724
rect 6763 28720 6819 28724
rect 6681 28668 6702 28720
rect 6702 28668 6737 28720
rect 6763 28668 6768 28720
rect 6768 28668 6819 28720
rect 6845 28668 6901 28724
rect 6927 28668 6983 28724
rect 7009 28668 7065 28724
rect 7091 28668 7147 28724
rect 7173 28668 7229 28724
rect 7255 28720 7311 28724
rect 7337 28720 7393 28724
rect 7255 28668 7256 28720
rect 7256 28668 7308 28720
rect 7308 28668 7311 28720
rect 7337 28668 7374 28720
rect 7374 28668 7393 28720
rect 7419 28668 7475 28724
rect 7501 28668 7557 28724
rect 7583 28668 7639 28724
rect 7665 28668 7721 28724
rect 7747 28668 7803 28724
rect 7829 28720 7885 28724
rect 7911 28720 7967 28724
rect 7829 28668 7862 28720
rect 7862 28668 7876 28720
rect 7876 28668 7885 28720
rect 7911 28668 7928 28720
rect 7928 28668 7967 28720
rect 7993 28672 8047 28724
rect 8047 28672 8049 28724
rect 8075 28672 8099 28724
rect 8099 28672 8131 28724
rect 7993 28668 8049 28672
rect 8075 28668 8131 28672
rect 8157 28672 8169 28724
rect 8169 28672 8213 28724
rect 8157 28668 8213 28672
rect 5613 28599 5646 28644
rect 5646 28599 5660 28644
rect 5660 28599 5669 28644
rect 5696 28599 5712 28644
rect 5712 28599 5752 28644
rect 5613 28588 5669 28599
rect 5696 28588 5752 28599
rect 5779 28588 5835 28644
rect 5861 28588 5917 28644
rect 5943 28588 5999 28644
rect 6025 28588 6081 28644
rect 6107 28599 6148 28644
rect 6148 28599 6163 28644
rect 6189 28599 6200 28644
rect 6200 28599 6214 28644
rect 6214 28599 6245 28644
rect 6107 28588 6163 28599
rect 6189 28588 6245 28599
rect 6271 28588 6327 28644
rect 6353 28588 6409 28644
rect 6435 28588 6491 28644
rect 6517 28588 6573 28644
rect 6599 28588 6655 28644
rect 6681 28599 6702 28644
rect 6702 28599 6737 28644
rect 6763 28599 6768 28644
rect 6768 28599 6819 28644
rect 6681 28588 6737 28599
rect 6763 28588 6819 28599
rect 6845 28588 6901 28644
rect 6927 28588 6983 28644
rect 7009 28588 7065 28644
rect 7091 28588 7147 28644
rect 7173 28588 7229 28644
rect 7255 28599 7256 28644
rect 7256 28599 7308 28644
rect 7308 28599 7311 28644
rect 7337 28599 7374 28644
rect 7374 28599 7393 28644
rect 7255 28588 7311 28599
rect 7337 28588 7393 28599
rect 7419 28588 7475 28644
rect 7501 28588 7557 28644
rect 7583 28588 7639 28644
rect 7665 28588 7721 28644
rect 7747 28588 7803 28644
rect 7829 28599 7862 28644
rect 7862 28599 7876 28644
rect 7876 28599 7885 28644
rect 7911 28599 7928 28644
rect 7928 28599 7967 28644
rect 7829 28588 7885 28599
rect 7911 28588 7967 28599
rect 7993 28603 8047 28644
rect 8047 28603 8049 28644
rect 8075 28603 8099 28644
rect 8099 28603 8131 28644
rect 7993 28588 8049 28603
rect 8075 28588 8131 28603
rect 8157 28603 8169 28644
rect 8169 28603 8213 28644
rect 8157 28588 8213 28603
rect 5613 28530 5646 28564
rect 5646 28530 5660 28564
rect 5660 28530 5669 28564
rect 5696 28530 5712 28564
rect 5712 28530 5752 28564
rect 5613 28513 5669 28530
rect 5696 28513 5752 28530
rect 5613 28508 5646 28513
rect 5646 28508 5660 28513
rect 5660 28508 5669 28513
rect 5696 28508 5712 28513
rect 5712 28508 5752 28513
rect 5779 28508 5835 28564
rect 5861 28508 5917 28564
rect 5943 28508 5999 28564
rect 6025 28508 6081 28564
rect 6107 28530 6148 28564
rect 6148 28530 6163 28564
rect 6189 28530 6200 28564
rect 6200 28530 6214 28564
rect 6214 28530 6245 28564
rect 6107 28513 6163 28530
rect 6189 28513 6245 28530
rect 6107 28508 6148 28513
rect 6148 28508 6163 28513
rect 6189 28508 6200 28513
rect 6200 28508 6214 28513
rect 6214 28508 6245 28513
rect 6271 28508 6327 28564
rect 6353 28508 6409 28564
rect 6435 28508 6491 28564
rect 6517 28508 6573 28564
rect 6599 28508 6655 28564
rect 6681 28530 6702 28564
rect 6702 28530 6737 28564
rect 6763 28530 6768 28564
rect 6768 28530 6819 28564
rect 6681 28513 6737 28530
rect 6763 28513 6819 28530
rect 6681 28508 6702 28513
rect 6702 28508 6737 28513
rect 6763 28508 6768 28513
rect 6768 28508 6819 28513
rect 6845 28508 6901 28564
rect 6927 28508 6983 28564
rect 7009 28508 7065 28564
rect 7091 28508 7147 28564
rect 7173 28508 7229 28564
rect 7255 28530 7256 28564
rect 7256 28530 7308 28564
rect 7308 28530 7311 28564
rect 7337 28530 7374 28564
rect 7374 28530 7393 28564
rect 7255 28513 7311 28530
rect 7337 28513 7393 28530
rect 7255 28508 7256 28513
rect 7256 28508 7308 28513
rect 7308 28508 7311 28513
rect 7337 28508 7374 28513
rect 7374 28508 7393 28513
rect 7419 28508 7475 28564
rect 7501 28508 7557 28564
rect 7583 28508 7639 28564
rect 7665 28508 7721 28564
rect 7747 28508 7803 28564
rect 7829 28530 7862 28564
rect 7862 28530 7876 28564
rect 7876 28530 7885 28564
rect 7911 28530 7928 28564
rect 7928 28530 7967 28564
rect 7829 28513 7885 28530
rect 7911 28513 7967 28530
rect 7829 28508 7862 28513
rect 7862 28508 7876 28513
rect 7876 28508 7885 28513
rect 7911 28508 7928 28513
rect 7928 28508 7967 28513
rect 7993 28534 8047 28564
rect 8047 28534 8049 28564
rect 8075 28534 8099 28564
rect 8099 28534 8131 28564
rect 7993 28517 8049 28534
rect 8075 28517 8131 28534
rect 7993 28508 8047 28517
rect 8047 28508 8049 28517
rect 8075 28508 8099 28517
rect 8099 28508 8131 28517
rect 8157 28534 8169 28564
rect 8169 28534 8213 28564
rect 8157 28517 8213 28534
rect 8157 28508 8169 28517
rect 8169 28508 8213 28517
rect 5613 28461 5646 28484
rect 5646 28461 5660 28484
rect 5660 28461 5669 28484
rect 5696 28461 5712 28484
rect 5712 28461 5752 28484
rect 5613 28444 5669 28461
rect 5696 28444 5752 28461
rect 5613 28428 5646 28444
rect 5646 28428 5660 28444
rect 5660 28428 5669 28444
rect 5696 28428 5712 28444
rect 5712 28428 5752 28444
rect 5779 28428 5835 28484
rect 5861 28428 5917 28484
rect 5943 28428 5999 28484
rect 6025 28428 6081 28484
rect 6107 28461 6148 28484
rect 6148 28461 6163 28484
rect 6189 28461 6200 28484
rect 6200 28461 6214 28484
rect 6214 28461 6245 28484
rect 6107 28444 6163 28461
rect 6189 28444 6245 28461
rect 6107 28428 6148 28444
rect 6148 28428 6163 28444
rect 6189 28428 6200 28444
rect 6200 28428 6214 28444
rect 6214 28428 6245 28444
rect 6271 28428 6327 28484
rect 6353 28428 6409 28484
rect 6435 28428 6491 28484
rect 6517 28428 6573 28484
rect 6599 28428 6655 28484
rect 6681 28461 6702 28484
rect 6702 28461 6737 28484
rect 6763 28461 6768 28484
rect 6768 28461 6819 28484
rect 6681 28444 6737 28461
rect 6763 28444 6819 28461
rect 6681 28428 6702 28444
rect 6702 28428 6737 28444
rect 6763 28428 6768 28444
rect 6768 28428 6819 28444
rect 6845 28428 6901 28484
rect 6927 28428 6983 28484
rect 7009 28428 7065 28484
rect 7091 28428 7147 28484
rect 7173 28428 7229 28484
rect 7255 28461 7256 28484
rect 7256 28461 7308 28484
rect 7308 28461 7311 28484
rect 7337 28461 7374 28484
rect 7374 28461 7393 28484
rect 7255 28444 7311 28461
rect 7337 28444 7393 28461
rect 7255 28428 7256 28444
rect 7256 28428 7308 28444
rect 7308 28428 7311 28444
rect 7337 28428 7374 28444
rect 7374 28428 7393 28444
rect 7419 28428 7475 28484
rect 7501 28428 7557 28484
rect 7583 28428 7639 28484
rect 7665 28428 7721 28484
rect 7747 28428 7803 28484
rect 7829 28461 7862 28484
rect 7862 28461 7876 28484
rect 7876 28461 7885 28484
rect 7911 28461 7928 28484
rect 7928 28461 7967 28484
rect 7829 28444 7885 28461
rect 7911 28444 7967 28461
rect 7829 28428 7862 28444
rect 7862 28428 7876 28444
rect 7876 28428 7885 28444
rect 7911 28428 7928 28444
rect 7928 28428 7967 28444
rect 7993 28465 8047 28484
rect 8047 28465 8049 28484
rect 8075 28465 8099 28484
rect 8099 28465 8131 28484
rect 7993 28448 8049 28465
rect 8075 28448 8131 28465
rect 7993 28428 8047 28448
rect 8047 28428 8049 28448
rect 8075 28428 8099 28448
rect 8099 28428 8131 28448
rect 8157 28465 8169 28484
rect 8169 28465 8213 28484
rect 8157 28448 8213 28465
rect 8157 28428 8169 28448
rect 8169 28428 8213 28448
rect 5613 28392 5646 28404
rect 5646 28392 5660 28404
rect 5660 28392 5669 28404
rect 5696 28392 5712 28404
rect 5712 28392 5752 28404
rect 5613 28375 5669 28392
rect 5696 28375 5752 28392
rect 5613 28348 5646 28375
rect 5646 28348 5660 28375
rect 5660 28348 5669 28375
rect 5696 28348 5712 28375
rect 5712 28348 5752 28375
rect 5779 28348 5835 28404
rect 5861 28348 5917 28404
rect 5943 28348 5999 28404
rect 6025 28348 6081 28404
rect 6107 28392 6148 28404
rect 6148 28392 6163 28404
rect 6189 28392 6200 28404
rect 6200 28392 6214 28404
rect 6214 28392 6245 28404
rect 6107 28375 6163 28392
rect 6189 28375 6245 28392
rect 6107 28348 6148 28375
rect 6148 28348 6163 28375
rect 6189 28348 6200 28375
rect 6200 28348 6214 28375
rect 6214 28348 6245 28375
rect 6271 28348 6327 28404
rect 6353 28348 6409 28404
rect 6435 28348 6491 28404
rect 6517 28348 6573 28404
rect 6599 28348 6655 28404
rect 6681 28392 6702 28404
rect 6702 28392 6737 28404
rect 6763 28392 6768 28404
rect 6768 28392 6819 28404
rect 6681 28375 6737 28392
rect 6763 28375 6819 28392
rect 6681 28348 6702 28375
rect 6702 28348 6737 28375
rect 6763 28348 6768 28375
rect 6768 28348 6819 28375
rect 6845 28348 6901 28404
rect 6927 28348 6983 28404
rect 7009 28348 7065 28404
rect 7091 28348 7147 28404
rect 7173 28348 7229 28404
rect 7255 28392 7256 28404
rect 7256 28392 7308 28404
rect 7308 28392 7311 28404
rect 7337 28392 7374 28404
rect 7374 28392 7393 28404
rect 7255 28375 7311 28392
rect 7337 28375 7393 28392
rect 7255 28348 7256 28375
rect 7256 28348 7308 28375
rect 7308 28348 7311 28375
rect 7337 28348 7374 28375
rect 7374 28348 7393 28375
rect 7419 28348 7475 28404
rect 7501 28348 7557 28404
rect 7583 28348 7639 28404
rect 7665 28348 7721 28404
rect 7747 28348 7803 28404
rect 7829 28392 7862 28404
rect 7862 28392 7876 28404
rect 7876 28392 7885 28404
rect 7911 28392 7928 28404
rect 7928 28392 7967 28404
rect 7829 28375 7885 28392
rect 7911 28375 7967 28392
rect 7829 28348 7862 28375
rect 7862 28348 7876 28375
rect 7876 28348 7885 28375
rect 7911 28348 7928 28375
rect 7928 28348 7967 28375
rect 7993 28396 8047 28404
rect 8047 28396 8049 28404
rect 8075 28396 8099 28404
rect 8099 28396 8131 28404
rect 7993 28378 8049 28396
rect 8075 28378 8131 28396
rect 7993 28348 8047 28378
rect 8047 28348 8049 28378
rect 8075 28348 8099 28378
rect 8099 28348 8131 28378
rect 8157 28396 8169 28404
rect 8169 28396 8213 28404
rect 8157 28378 8213 28396
rect 8157 28348 8169 28378
rect 8169 28348 8213 28378
rect 5613 28323 5646 28324
rect 5646 28323 5660 28324
rect 5660 28323 5669 28324
rect 5696 28323 5712 28324
rect 5712 28323 5752 28324
rect 5613 28306 5669 28323
rect 5696 28306 5752 28323
rect 5613 28268 5646 28306
rect 5646 28268 5660 28306
rect 5660 28268 5669 28306
rect 5696 28268 5712 28306
rect 5712 28268 5752 28306
rect 5779 28268 5835 28324
rect 5861 28268 5917 28324
rect 5943 28268 5999 28324
rect 6025 28268 6081 28324
rect 6107 28323 6148 28324
rect 6148 28323 6163 28324
rect 6189 28323 6200 28324
rect 6200 28323 6214 28324
rect 6214 28323 6245 28324
rect 6107 28306 6163 28323
rect 6189 28306 6245 28323
rect 6107 28268 6148 28306
rect 6148 28268 6163 28306
rect 6189 28268 6200 28306
rect 6200 28268 6214 28306
rect 6214 28268 6245 28306
rect 6271 28268 6327 28324
rect 6353 28268 6409 28324
rect 6435 28268 6491 28324
rect 6517 28268 6573 28324
rect 6599 28268 6655 28324
rect 6681 28323 6702 28324
rect 6702 28323 6737 28324
rect 6763 28323 6768 28324
rect 6768 28323 6819 28324
rect 6681 28306 6737 28323
rect 6763 28306 6819 28323
rect 6681 28268 6702 28306
rect 6702 28268 6737 28306
rect 6763 28268 6768 28306
rect 6768 28268 6819 28306
rect 6845 28268 6901 28324
rect 6927 28268 6983 28324
rect 7009 28268 7065 28324
rect 7091 28268 7147 28324
rect 7173 28268 7229 28324
rect 7255 28323 7256 28324
rect 7256 28323 7308 28324
rect 7308 28323 7311 28324
rect 7337 28323 7374 28324
rect 7374 28323 7393 28324
rect 7255 28306 7311 28323
rect 7337 28306 7393 28323
rect 7255 28268 7256 28306
rect 7256 28268 7308 28306
rect 7308 28268 7311 28306
rect 7337 28268 7374 28306
rect 7374 28268 7393 28306
rect 7419 28268 7475 28324
rect 7501 28268 7557 28324
rect 7583 28268 7639 28324
rect 7665 28268 7721 28324
rect 7747 28268 7803 28324
rect 7829 28323 7862 28324
rect 7862 28323 7876 28324
rect 7876 28323 7885 28324
rect 7911 28323 7928 28324
rect 7928 28323 7967 28324
rect 7829 28306 7885 28323
rect 7911 28306 7967 28323
rect 7829 28268 7862 28306
rect 7862 28268 7876 28306
rect 7876 28268 7885 28306
rect 7911 28268 7928 28306
rect 7928 28268 7967 28306
rect 7993 28308 8049 28324
rect 8075 28308 8131 28324
rect 7993 28268 8047 28308
rect 8047 28268 8049 28308
rect 8075 28268 8099 28308
rect 8099 28268 8131 28308
rect 8157 28308 8213 28324
rect 8157 28268 8169 28308
rect 8169 28268 8213 28308
rect 5613 28236 5669 28244
rect 5696 28236 5752 28244
rect 5613 28188 5646 28236
rect 5646 28188 5660 28236
rect 5660 28188 5669 28236
rect 5696 28188 5712 28236
rect 5712 28188 5752 28236
rect 5779 28188 5835 28244
rect 5861 28188 5917 28244
rect 5943 28188 5999 28244
rect 6025 28188 6081 28244
rect 6107 28236 6163 28244
rect 6189 28236 6245 28244
rect 6107 28188 6148 28236
rect 6148 28188 6163 28236
rect 6189 28188 6200 28236
rect 6200 28188 6214 28236
rect 6214 28188 6245 28236
rect 6271 28188 6327 28244
rect 6353 28188 6409 28244
rect 6435 28188 6491 28244
rect 6517 28188 6573 28244
rect 6599 28188 6655 28244
rect 6681 28236 6737 28244
rect 6763 28236 6819 28244
rect 6681 28188 6702 28236
rect 6702 28188 6737 28236
rect 6763 28188 6768 28236
rect 6768 28188 6819 28236
rect 6845 28188 6901 28244
rect 6927 28188 6983 28244
rect 7009 28188 7065 28244
rect 7091 28188 7147 28244
rect 7173 28188 7229 28244
rect 7255 28236 7311 28244
rect 7337 28236 7393 28244
rect 7255 28188 7256 28236
rect 7256 28188 7308 28236
rect 7308 28188 7311 28236
rect 7337 28188 7374 28236
rect 7374 28188 7393 28236
rect 7419 28188 7475 28244
rect 7501 28188 7557 28244
rect 7583 28188 7639 28244
rect 7665 28188 7721 28244
rect 7747 28188 7803 28244
rect 7829 28236 7885 28244
rect 7911 28236 7967 28244
rect 7829 28188 7862 28236
rect 7862 28188 7876 28236
rect 7876 28188 7885 28236
rect 7911 28188 7928 28236
rect 7928 28188 7967 28236
rect 7993 28238 8049 28244
rect 8075 28238 8131 28244
rect 7993 28188 8047 28238
rect 8047 28188 8049 28238
rect 8075 28188 8099 28238
rect 8099 28188 8131 28238
rect 8157 28238 8213 28244
rect 8157 28188 8169 28238
rect 8169 28188 8213 28238
rect 5613 28114 5646 28164
rect 5646 28114 5660 28164
rect 5660 28114 5669 28164
rect 5696 28114 5712 28164
rect 5712 28114 5752 28164
rect 5613 28108 5669 28114
rect 5696 28108 5752 28114
rect 5779 28108 5835 28164
rect 5861 28108 5917 28164
rect 5943 28108 5999 28164
rect 6025 28108 6081 28164
rect 6107 28114 6148 28164
rect 6148 28114 6163 28164
rect 6189 28114 6200 28164
rect 6200 28114 6214 28164
rect 6214 28114 6245 28164
rect 6107 28108 6163 28114
rect 6189 28108 6245 28114
rect 6271 28108 6327 28164
rect 6353 28108 6409 28164
rect 6435 28108 6491 28164
rect 6517 28108 6573 28164
rect 6599 28108 6655 28164
rect 6681 28114 6702 28164
rect 6702 28114 6737 28164
rect 6763 28114 6768 28164
rect 6768 28114 6819 28164
rect 6681 28108 6737 28114
rect 6763 28108 6819 28114
rect 6845 28108 6901 28164
rect 6927 28108 6983 28164
rect 7009 28108 7065 28164
rect 7091 28108 7147 28164
rect 7173 28108 7229 28164
rect 7255 28114 7256 28164
rect 7256 28114 7308 28164
rect 7308 28114 7311 28164
rect 7337 28114 7374 28164
rect 7374 28114 7393 28164
rect 7255 28108 7311 28114
rect 7337 28108 7393 28114
rect 7419 28108 7475 28164
rect 7501 28108 7557 28164
rect 7583 28108 7639 28164
rect 7665 28108 7721 28164
rect 7747 28108 7803 28164
rect 7829 28114 7862 28164
rect 7862 28114 7876 28164
rect 7876 28114 7885 28164
rect 7911 28114 7928 28164
rect 7928 28114 7967 28164
rect 7829 28108 7885 28114
rect 7911 28108 7967 28114
rect 7993 28116 8047 28164
rect 8047 28116 8049 28164
rect 8075 28116 8099 28164
rect 8099 28116 8131 28164
rect 7993 28108 8049 28116
rect 8075 28108 8131 28116
rect 8157 28116 8169 28164
rect 8169 28116 8213 28164
rect 8157 28108 8213 28116
rect 2733 27931 2789 27987
rect 2814 27931 2870 27987
rect 2895 27931 2951 27987
rect 2976 27931 3032 27987
rect 3057 27931 3113 27987
rect 3138 27931 3194 27987
rect 3219 27931 3275 27987
rect 3300 27931 3356 27987
rect 3381 27931 3437 27987
rect 3462 27931 3518 27987
rect 3543 27931 3599 27987
rect 3624 27931 3680 27987
rect 3705 27931 3761 27987
rect 3786 27931 3842 27987
rect 3867 27931 3923 27987
rect 3948 27931 4004 27987
rect 4029 27931 4085 27987
rect 4110 27931 4166 27987
rect 4191 27931 4247 27987
rect 4272 27931 4328 27987
rect 4353 27931 4409 27987
rect 4434 27931 4490 27987
rect 4515 27931 4571 27987
rect 4596 27931 4652 27987
rect 4677 27931 4733 27987
rect 4758 27931 4814 27987
rect 4839 27931 4895 27987
rect 4920 27931 4976 27987
rect 5001 27931 5057 27987
rect 5082 27931 5138 27987
rect 2733 27851 2789 27907
rect 2814 27851 2870 27907
rect 2895 27851 2951 27907
rect 2976 27851 3032 27907
rect 3057 27851 3113 27907
rect 3138 27851 3194 27907
rect 3219 27851 3275 27907
rect 3300 27851 3356 27907
rect 3381 27851 3437 27907
rect 3462 27851 3518 27907
rect 3543 27851 3599 27907
rect 3624 27851 3680 27907
rect 3705 27851 3761 27907
rect 3786 27851 3842 27907
rect 3867 27851 3923 27907
rect 3948 27851 4004 27907
rect 4029 27851 4085 27907
rect 4110 27851 4166 27907
rect 4191 27851 4247 27907
rect 4272 27851 4328 27907
rect 4353 27851 4409 27907
rect 4434 27851 4490 27907
rect 4515 27851 4571 27907
rect 4596 27851 4652 27907
rect 4677 27851 4733 27907
rect 4758 27851 4814 27907
rect 4839 27851 4895 27907
rect 4920 27851 4976 27907
rect 5001 27851 5057 27907
rect 5082 27851 5138 27907
rect 2733 27771 2789 27827
rect 2814 27771 2870 27827
rect 2895 27771 2951 27827
rect 2976 27771 3032 27827
rect 3057 27771 3113 27827
rect 3138 27771 3194 27827
rect 3219 27771 3275 27827
rect 3300 27771 3356 27827
rect 3381 27771 3437 27827
rect 3462 27771 3518 27827
rect 3543 27771 3599 27827
rect 3624 27771 3680 27827
rect 3705 27771 3761 27827
rect 3786 27771 3842 27827
rect 3867 27771 3923 27827
rect 3948 27771 4004 27827
rect 4029 27771 4085 27827
rect 4110 27771 4166 27827
rect 4191 27771 4247 27827
rect 4272 27771 4328 27827
rect 4353 27771 4409 27827
rect 4434 27771 4490 27827
rect 4515 27771 4571 27827
rect 4596 27771 4652 27827
rect 4677 27771 4733 27827
rect 4758 27771 4814 27827
rect 4839 27771 4895 27827
rect 4920 27771 4976 27827
rect 5001 27771 5057 27827
rect 5082 27771 5138 27827
rect 2733 27691 2789 27747
rect 2814 27691 2870 27747
rect 2895 27691 2951 27747
rect 2976 27691 3032 27747
rect 3057 27691 3113 27747
rect 3138 27691 3194 27747
rect 3219 27691 3275 27747
rect 3300 27691 3356 27747
rect 3381 27691 3437 27747
rect 3462 27691 3518 27747
rect 3543 27691 3599 27747
rect 3624 27691 3680 27747
rect 3705 27691 3761 27747
rect 3786 27691 3842 27747
rect 3867 27691 3923 27747
rect 3948 27691 4004 27747
rect 4029 27691 4085 27747
rect 4110 27691 4166 27747
rect 4191 27691 4247 27747
rect 4272 27691 4328 27747
rect 4353 27691 4409 27747
rect 4434 27691 4490 27747
rect 4515 27691 4571 27747
rect 4596 27691 4652 27747
rect 4677 27691 4733 27747
rect 4758 27691 4814 27747
rect 4839 27691 4895 27747
rect 4920 27691 4976 27747
rect 5001 27691 5057 27747
rect 5082 27691 5138 27747
rect 2733 27611 2789 27667
rect 2814 27611 2870 27667
rect 2895 27611 2951 27667
rect 2976 27611 3032 27667
rect 3057 27611 3113 27667
rect 3138 27611 3194 27667
rect 3219 27611 3275 27667
rect 3300 27611 3356 27667
rect 3381 27611 3437 27667
rect 3462 27611 3518 27667
rect 3543 27611 3599 27667
rect 3624 27611 3680 27667
rect 3705 27611 3761 27667
rect 3786 27611 3842 27667
rect 3867 27611 3923 27667
rect 3948 27611 4004 27667
rect 4029 27611 4085 27667
rect 4110 27611 4166 27667
rect 4191 27611 4247 27667
rect 4272 27611 4328 27667
rect 4353 27611 4409 27667
rect 4434 27611 4490 27667
rect 4515 27611 4571 27667
rect 4596 27611 4652 27667
rect 4677 27611 4733 27667
rect 4758 27611 4814 27667
rect 4839 27611 4895 27667
rect 4920 27611 4976 27667
rect 5001 27611 5057 27667
rect 5082 27611 5138 27667
rect 2733 27531 2789 27587
rect 2814 27531 2870 27587
rect 2895 27531 2951 27587
rect 2976 27531 3032 27587
rect 3057 27531 3113 27587
rect 3138 27531 3194 27587
rect 3219 27531 3275 27587
rect 3300 27531 3356 27587
rect 3381 27531 3437 27587
rect 3462 27531 3518 27587
rect 3543 27531 3599 27587
rect 3624 27531 3680 27587
rect 3705 27531 3761 27587
rect 3786 27531 3842 27587
rect 3867 27531 3923 27587
rect 3948 27531 4004 27587
rect 4029 27531 4085 27587
rect 4110 27531 4166 27587
rect 4191 27531 4247 27587
rect 4272 27531 4328 27587
rect 4353 27531 4409 27587
rect 4434 27531 4490 27587
rect 4515 27531 4571 27587
rect 4596 27531 4652 27587
rect 4677 27531 4733 27587
rect 4758 27531 4814 27587
rect 4839 27531 4895 27587
rect 4920 27531 4976 27587
rect 5001 27531 5057 27587
rect 5082 27531 5138 27587
rect 2733 27451 2789 27507
rect 2814 27451 2870 27507
rect 2895 27451 2951 27507
rect 2976 27451 3032 27507
rect 3057 27451 3113 27507
rect 3138 27451 3194 27507
rect 3219 27451 3275 27507
rect 3300 27451 3356 27507
rect 3381 27451 3437 27507
rect 3462 27451 3518 27507
rect 3543 27451 3599 27507
rect 3624 27451 3680 27507
rect 3705 27451 3761 27507
rect 3786 27451 3842 27507
rect 3867 27451 3923 27507
rect 3948 27451 4004 27507
rect 4029 27451 4085 27507
rect 4110 27451 4166 27507
rect 4191 27451 4247 27507
rect 4272 27451 4328 27507
rect 4353 27451 4409 27507
rect 4434 27451 4490 27507
rect 4515 27451 4571 27507
rect 4596 27451 4652 27507
rect 4677 27451 4733 27507
rect 4758 27451 4814 27507
rect 4839 27451 4895 27507
rect 4920 27451 4976 27507
rect 5001 27451 5057 27507
rect 5082 27451 5138 27507
rect 2733 27371 2789 27427
rect 2814 27371 2870 27427
rect 2895 27371 2951 27427
rect 2976 27371 3032 27427
rect 3057 27371 3113 27427
rect 3138 27371 3194 27427
rect 3219 27371 3275 27427
rect 3300 27371 3356 27427
rect 3381 27371 3437 27427
rect 3462 27371 3518 27427
rect 3543 27371 3599 27427
rect 3624 27371 3680 27427
rect 3705 27371 3761 27427
rect 3786 27371 3842 27427
rect 3867 27371 3923 27427
rect 3948 27371 4004 27427
rect 4029 27371 4085 27427
rect 4110 27371 4166 27427
rect 4191 27371 4247 27427
rect 4272 27371 4328 27427
rect 4353 27371 4409 27427
rect 4434 27371 4490 27427
rect 4515 27371 4571 27427
rect 4596 27371 4652 27427
rect 4677 27371 4733 27427
rect 4758 27371 4814 27427
rect 4839 27371 4895 27427
rect 4920 27371 4976 27427
rect 5001 27371 5057 27427
rect 5082 27371 5138 27427
rect 5163 27371 5299 27987
rect 5613 26720 5669 26724
rect 5696 26720 5752 26724
rect 5613 26668 5646 26720
rect 5646 26668 5660 26720
rect 5660 26668 5669 26720
rect 5696 26668 5712 26720
rect 5712 26668 5752 26720
rect 5779 26668 5835 26724
rect 5861 26668 5917 26724
rect 5943 26668 5999 26724
rect 6025 26668 6081 26724
rect 6107 26720 6163 26724
rect 6189 26720 6245 26724
rect 6107 26668 6148 26720
rect 6148 26668 6163 26720
rect 6189 26668 6200 26720
rect 6200 26668 6214 26720
rect 6214 26668 6245 26720
rect 6271 26668 6327 26724
rect 6353 26668 6409 26724
rect 6435 26668 6491 26724
rect 6517 26668 6573 26724
rect 6599 26668 6655 26724
rect 6681 26720 6737 26724
rect 6763 26720 6819 26724
rect 6681 26668 6702 26720
rect 6702 26668 6737 26720
rect 6763 26668 6768 26720
rect 6768 26668 6819 26720
rect 6845 26668 6901 26724
rect 6927 26668 6983 26724
rect 7009 26668 7065 26724
rect 7091 26668 7147 26724
rect 7173 26668 7229 26724
rect 7255 26720 7311 26724
rect 7337 26720 7393 26724
rect 7255 26668 7256 26720
rect 7256 26668 7308 26720
rect 7308 26668 7311 26720
rect 7337 26668 7374 26720
rect 7374 26668 7393 26720
rect 7419 26668 7475 26724
rect 7501 26668 7557 26724
rect 7583 26668 7639 26724
rect 7665 26668 7721 26724
rect 7747 26668 7803 26724
rect 7829 26720 7885 26724
rect 7911 26720 7967 26724
rect 7829 26668 7862 26720
rect 7862 26668 7876 26720
rect 7876 26668 7885 26720
rect 7911 26668 7928 26720
rect 7928 26668 7967 26720
rect 7993 26672 8047 26724
rect 8047 26672 8049 26724
rect 8075 26672 8099 26724
rect 8099 26672 8131 26724
rect 7993 26668 8049 26672
rect 8075 26668 8131 26672
rect 8157 26672 8169 26724
rect 8169 26672 8213 26724
rect 8157 26668 8213 26672
rect 5613 26599 5646 26644
rect 5646 26599 5660 26644
rect 5660 26599 5669 26644
rect 5696 26599 5712 26644
rect 5712 26599 5752 26644
rect 5613 26588 5669 26599
rect 5696 26588 5752 26599
rect 5779 26588 5835 26644
rect 5861 26588 5917 26644
rect 5943 26588 5999 26644
rect 6025 26588 6081 26644
rect 6107 26599 6148 26644
rect 6148 26599 6163 26644
rect 6189 26599 6200 26644
rect 6200 26599 6214 26644
rect 6214 26599 6245 26644
rect 6107 26588 6163 26599
rect 6189 26588 6245 26599
rect 6271 26588 6327 26644
rect 6353 26588 6409 26644
rect 6435 26588 6491 26644
rect 6517 26588 6573 26644
rect 6599 26588 6655 26644
rect 6681 26599 6702 26644
rect 6702 26599 6737 26644
rect 6763 26599 6768 26644
rect 6768 26599 6819 26644
rect 6681 26588 6737 26599
rect 6763 26588 6819 26599
rect 6845 26588 6901 26644
rect 6927 26588 6983 26644
rect 7009 26588 7065 26644
rect 7091 26588 7147 26644
rect 7173 26588 7229 26644
rect 7255 26599 7256 26644
rect 7256 26599 7308 26644
rect 7308 26599 7311 26644
rect 7337 26599 7374 26644
rect 7374 26599 7393 26644
rect 7255 26588 7311 26599
rect 7337 26588 7393 26599
rect 7419 26588 7475 26644
rect 7501 26588 7557 26644
rect 7583 26588 7639 26644
rect 7665 26588 7721 26644
rect 7747 26588 7803 26644
rect 7829 26599 7862 26644
rect 7862 26599 7876 26644
rect 7876 26599 7885 26644
rect 7911 26599 7928 26644
rect 7928 26599 7967 26644
rect 7829 26588 7885 26599
rect 7911 26588 7967 26599
rect 7993 26603 8047 26644
rect 8047 26603 8049 26644
rect 8075 26603 8099 26644
rect 8099 26603 8131 26644
rect 7993 26588 8049 26603
rect 8075 26588 8131 26603
rect 8157 26603 8169 26644
rect 8169 26603 8213 26644
rect 8157 26588 8213 26603
rect 5613 26530 5646 26564
rect 5646 26530 5660 26564
rect 5660 26530 5669 26564
rect 5696 26530 5712 26564
rect 5712 26530 5752 26564
rect 5613 26513 5669 26530
rect 5696 26513 5752 26530
rect 5613 26508 5646 26513
rect 5646 26508 5660 26513
rect 5660 26508 5669 26513
rect 5696 26508 5712 26513
rect 5712 26508 5752 26513
rect 5779 26508 5835 26564
rect 5861 26508 5917 26564
rect 5943 26508 5999 26564
rect 6025 26508 6081 26564
rect 6107 26530 6148 26564
rect 6148 26530 6163 26564
rect 6189 26530 6200 26564
rect 6200 26530 6214 26564
rect 6214 26530 6245 26564
rect 6107 26513 6163 26530
rect 6189 26513 6245 26530
rect 6107 26508 6148 26513
rect 6148 26508 6163 26513
rect 6189 26508 6200 26513
rect 6200 26508 6214 26513
rect 6214 26508 6245 26513
rect 6271 26508 6327 26564
rect 6353 26508 6409 26564
rect 6435 26508 6491 26564
rect 6517 26508 6573 26564
rect 6599 26508 6655 26564
rect 6681 26530 6702 26564
rect 6702 26530 6737 26564
rect 6763 26530 6768 26564
rect 6768 26530 6819 26564
rect 6681 26513 6737 26530
rect 6763 26513 6819 26530
rect 6681 26508 6702 26513
rect 6702 26508 6737 26513
rect 6763 26508 6768 26513
rect 6768 26508 6819 26513
rect 6845 26508 6901 26564
rect 6927 26508 6983 26564
rect 7009 26508 7065 26564
rect 7091 26508 7147 26564
rect 7173 26508 7229 26564
rect 7255 26530 7256 26564
rect 7256 26530 7308 26564
rect 7308 26530 7311 26564
rect 7337 26530 7374 26564
rect 7374 26530 7393 26564
rect 7255 26513 7311 26530
rect 7337 26513 7393 26530
rect 7255 26508 7256 26513
rect 7256 26508 7308 26513
rect 7308 26508 7311 26513
rect 7337 26508 7374 26513
rect 7374 26508 7393 26513
rect 7419 26508 7475 26564
rect 7501 26508 7557 26564
rect 7583 26508 7639 26564
rect 7665 26508 7721 26564
rect 7747 26508 7803 26564
rect 7829 26530 7862 26564
rect 7862 26530 7876 26564
rect 7876 26530 7885 26564
rect 7911 26530 7928 26564
rect 7928 26530 7967 26564
rect 7829 26513 7885 26530
rect 7911 26513 7967 26530
rect 7829 26508 7862 26513
rect 7862 26508 7876 26513
rect 7876 26508 7885 26513
rect 7911 26508 7928 26513
rect 7928 26508 7967 26513
rect 7993 26534 8047 26564
rect 8047 26534 8049 26564
rect 8075 26534 8099 26564
rect 8099 26534 8131 26564
rect 7993 26517 8049 26534
rect 8075 26517 8131 26534
rect 7993 26508 8047 26517
rect 8047 26508 8049 26517
rect 8075 26508 8099 26517
rect 8099 26508 8131 26517
rect 8157 26534 8169 26564
rect 8169 26534 8213 26564
rect 8157 26517 8213 26534
rect 8157 26508 8169 26517
rect 8169 26508 8213 26517
rect 5613 26461 5646 26484
rect 5646 26461 5660 26484
rect 5660 26461 5669 26484
rect 5696 26461 5712 26484
rect 5712 26461 5752 26484
rect 5613 26444 5669 26461
rect 5696 26444 5752 26461
rect 5613 26428 5646 26444
rect 5646 26428 5660 26444
rect 5660 26428 5669 26444
rect 5696 26428 5712 26444
rect 5712 26428 5752 26444
rect 5779 26428 5835 26484
rect 5861 26428 5917 26484
rect 5943 26428 5999 26484
rect 6025 26428 6081 26484
rect 6107 26461 6148 26484
rect 6148 26461 6163 26484
rect 6189 26461 6200 26484
rect 6200 26461 6214 26484
rect 6214 26461 6245 26484
rect 6107 26444 6163 26461
rect 6189 26444 6245 26461
rect 6107 26428 6148 26444
rect 6148 26428 6163 26444
rect 6189 26428 6200 26444
rect 6200 26428 6214 26444
rect 6214 26428 6245 26444
rect 6271 26428 6327 26484
rect 6353 26428 6409 26484
rect 6435 26428 6491 26484
rect 6517 26428 6573 26484
rect 6599 26428 6655 26484
rect 6681 26461 6702 26484
rect 6702 26461 6737 26484
rect 6763 26461 6768 26484
rect 6768 26461 6819 26484
rect 6681 26444 6737 26461
rect 6763 26444 6819 26461
rect 6681 26428 6702 26444
rect 6702 26428 6737 26444
rect 6763 26428 6768 26444
rect 6768 26428 6819 26444
rect 6845 26428 6901 26484
rect 6927 26428 6983 26484
rect 7009 26428 7065 26484
rect 7091 26428 7147 26484
rect 7173 26428 7229 26484
rect 7255 26461 7256 26484
rect 7256 26461 7308 26484
rect 7308 26461 7311 26484
rect 7337 26461 7374 26484
rect 7374 26461 7393 26484
rect 7255 26444 7311 26461
rect 7337 26444 7393 26461
rect 7255 26428 7256 26444
rect 7256 26428 7308 26444
rect 7308 26428 7311 26444
rect 7337 26428 7374 26444
rect 7374 26428 7393 26444
rect 7419 26428 7475 26484
rect 7501 26428 7557 26484
rect 7583 26428 7639 26484
rect 7665 26428 7721 26484
rect 7747 26428 7803 26484
rect 7829 26461 7862 26484
rect 7862 26461 7876 26484
rect 7876 26461 7885 26484
rect 7911 26461 7928 26484
rect 7928 26461 7967 26484
rect 7829 26444 7885 26461
rect 7911 26444 7967 26461
rect 7829 26428 7862 26444
rect 7862 26428 7876 26444
rect 7876 26428 7885 26444
rect 7911 26428 7928 26444
rect 7928 26428 7967 26444
rect 7993 26465 8047 26484
rect 8047 26465 8049 26484
rect 8075 26465 8099 26484
rect 8099 26465 8131 26484
rect 7993 26448 8049 26465
rect 8075 26448 8131 26465
rect 7993 26428 8047 26448
rect 8047 26428 8049 26448
rect 8075 26428 8099 26448
rect 8099 26428 8131 26448
rect 8157 26465 8169 26484
rect 8169 26465 8213 26484
rect 8157 26448 8213 26465
rect 8157 26428 8169 26448
rect 8169 26428 8213 26448
rect 5613 26392 5646 26404
rect 5646 26392 5660 26404
rect 5660 26392 5669 26404
rect 5696 26392 5712 26404
rect 5712 26392 5752 26404
rect 5613 26375 5669 26392
rect 5696 26375 5752 26392
rect 5613 26348 5646 26375
rect 5646 26348 5660 26375
rect 5660 26348 5669 26375
rect 5696 26348 5712 26375
rect 5712 26348 5752 26375
rect 5779 26348 5835 26404
rect 5861 26348 5917 26404
rect 5943 26348 5999 26404
rect 6025 26348 6081 26404
rect 6107 26392 6148 26404
rect 6148 26392 6163 26404
rect 6189 26392 6200 26404
rect 6200 26392 6214 26404
rect 6214 26392 6245 26404
rect 6107 26375 6163 26392
rect 6189 26375 6245 26392
rect 6107 26348 6148 26375
rect 6148 26348 6163 26375
rect 6189 26348 6200 26375
rect 6200 26348 6214 26375
rect 6214 26348 6245 26375
rect 6271 26348 6327 26404
rect 6353 26348 6409 26404
rect 6435 26348 6491 26404
rect 6517 26348 6573 26404
rect 6599 26348 6655 26404
rect 6681 26392 6702 26404
rect 6702 26392 6737 26404
rect 6763 26392 6768 26404
rect 6768 26392 6819 26404
rect 6681 26375 6737 26392
rect 6763 26375 6819 26392
rect 6681 26348 6702 26375
rect 6702 26348 6737 26375
rect 6763 26348 6768 26375
rect 6768 26348 6819 26375
rect 6845 26348 6901 26404
rect 6927 26348 6983 26404
rect 7009 26348 7065 26404
rect 7091 26348 7147 26404
rect 7173 26348 7229 26404
rect 7255 26392 7256 26404
rect 7256 26392 7308 26404
rect 7308 26392 7311 26404
rect 7337 26392 7374 26404
rect 7374 26392 7393 26404
rect 7255 26375 7311 26392
rect 7337 26375 7393 26392
rect 7255 26348 7256 26375
rect 7256 26348 7308 26375
rect 7308 26348 7311 26375
rect 7337 26348 7374 26375
rect 7374 26348 7393 26375
rect 7419 26348 7475 26404
rect 7501 26348 7557 26404
rect 7583 26348 7639 26404
rect 7665 26348 7721 26404
rect 7747 26348 7803 26404
rect 7829 26392 7862 26404
rect 7862 26392 7876 26404
rect 7876 26392 7885 26404
rect 7911 26392 7928 26404
rect 7928 26392 7967 26404
rect 7829 26375 7885 26392
rect 7911 26375 7967 26392
rect 7829 26348 7862 26375
rect 7862 26348 7876 26375
rect 7876 26348 7885 26375
rect 7911 26348 7928 26375
rect 7928 26348 7967 26375
rect 7993 26396 8047 26404
rect 8047 26396 8049 26404
rect 8075 26396 8099 26404
rect 8099 26396 8131 26404
rect 7993 26378 8049 26396
rect 8075 26378 8131 26396
rect 7993 26348 8047 26378
rect 8047 26348 8049 26378
rect 8075 26348 8099 26378
rect 8099 26348 8131 26378
rect 8157 26396 8169 26404
rect 8169 26396 8213 26404
rect 8157 26378 8213 26396
rect 8157 26348 8169 26378
rect 8169 26348 8213 26378
rect 5613 26323 5646 26324
rect 5646 26323 5660 26324
rect 5660 26323 5669 26324
rect 5696 26323 5712 26324
rect 5712 26323 5752 26324
rect 5613 26306 5669 26323
rect 5696 26306 5752 26323
rect 5613 26268 5646 26306
rect 5646 26268 5660 26306
rect 5660 26268 5669 26306
rect 5696 26268 5712 26306
rect 5712 26268 5752 26306
rect 5779 26268 5835 26324
rect 5861 26268 5917 26324
rect 5943 26268 5999 26324
rect 6025 26268 6081 26324
rect 6107 26323 6148 26324
rect 6148 26323 6163 26324
rect 6189 26323 6200 26324
rect 6200 26323 6214 26324
rect 6214 26323 6245 26324
rect 6107 26306 6163 26323
rect 6189 26306 6245 26323
rect 6107 26268 6148 26306
rect 6148 26268 6163 26306
rect 6189 26268 6200 26306
rect 6200 26268 6214 26306
rect 6214 26268 6245 26306
rect 6271 26268 6327 26324
rect 6353 26268 6409 26324
rect 6435 26268 6491 26324
rect 6517 26268 6573 26324
rect 6599 26268 6655 26324
rect 6681 26323 6702 26324
rect 6702 26323 6737 26324
rect 6763 26323 6768 26324
rect 6768 26323 6819 26324
rect 6681 26306 6737 26323
rect 6763 26306 6819 26323
rect 6681 26268 6702 26306
rect 6702 26268 6737 26306
rect 6763 26268 6768 26306
rect 6768 26268 6819 26306
rect 6845 26268 6901 26324
rect 6927 26268 6983 26324
rect 7009 26268 7065 26324
rect 7091 26268 7147 26324
rect 7173 26268 7229 26324
rect 7255 26323 7256 26324
rect 7256 26323 7308 26324
rect 7308 26323 7311 26324
rect 7337 26323 7374 26324
rect 7374 26323 7393 26324
rect 7255 26306 7311 26323
rect 7337 26306 7393 26323
rect 7255 26268 7256 26306
rect 7256 26268 7308 26306
rect 7308 26268 7311 26306
rect 7337 26268 7374 26306
rect 7374 26268 7393 26306
rect 7419 26268 7475 26324
rect 7501 26268 7557 26324
rect 7583 26268 7639 26324
rect 7665 26268 7721 26324
rect 7747 26268 7803 26324
rect 7829 26323 7862 26324
rect 7862 26323 7876 26324
rect 7876 26323 7885 26324
rect 7911 26323 7928 26324
rect 7928 26323 7967 26324
rect 7829 26306 7885 26323
rect 7911 26306 7967 26323
rect 7829 26268 7862 26306
rect 7862 26268 7876 26306
rect 7876 26268 7885 26306
rect 7911 26268 7928 26306
rect 7928 26268 7967 26306
rect 7993 26308 8049 26324
rect 8075 26308 8131 26324
rect 7993 26268 8047 26308
rect 8047 26268 8049 26308
rect 8075 26268 8099 26308
rect 8099 26268 8131 26308
rect 8157 26308 8213 26324
rect 8157 26268 8169 26308
rect 8169 26268 8213 26308
rect 5613 26236 5669 26244
rect 5696 26236 5752 26244
rect 5613 26188 5646 26236
rect 5646 26188 5660 26236
rect 5660 26188 5669 26236
rect 5696 26188 5712 26236
rect 5712 26188 5752 26236
rect 5779 26188 5835 26244
rect 5861 26188 5917 26244
rect 5943 26188 5999 26244
rect 6025 26188 6081 26244
rect 6107 26236 6163 26244
rect 6189 26236 6245 26244
rect 6107 26188 6148 26236
rect 6148 26188 6163 26236
rect 6189 26188 6200 26236
rect 6200 26188 6214 26236
rect 6214 26188 6245 26236
rect 6271 26188 6327 26244
rect 6353 26188 6409 26244
rect 6435 26188 6491 26244
rect 6517 26188 6573 26244
rect 6599 26188 6655 26244
rect 6681 26236 6737 26244
rect 6763 26236 6819 26244
rect 6681 26188 6702 26236
rect 6702 26188 6737 26236
rect 6763 26188 6768 26236
rect 6768 26188 6819 26236
rect 6845 26188 6901 26244
rect 6927 26188 6983 26244
rect 7009 26188 7065 26244
rect 7091 26188 7147 26244
rect 7173 26188 7229 26244
rect 7255 26236 7311 26244
rect 7337 26236 7393 26244
rect 7255 26188 7256 26236
rect 7256 26188 7308 26236
rect 7308 26188 7311 26236
rect 7337 26188 7374 26236
rect 7374 26188 7393 26236
rect 7419 26188 7475 26244
rect 7501 26188 7557 26244
rect 7583 26188 7639 26244
rect 7665 26188 7721 26244
rect 7747 26188 7803 26244
rect 7829 26236 7885 26244
rect 7911 26236 7967 26244
rect 7829 26188 7862 26236
rect 7862 26188 7876 26236
rect 7876 26188 7885 26236
rect 7911 26188 7928 26236
rect 7928 26188 7967 26236
rect 7993 26238 8049 26244
rect 8075 26238 8131 26244
rect 7993 26188 8047 26238
rect 8047 26188 8049 26238
rect 8075 26188 8099 26238
rect 8099 26188 8131 26238
rect 8157 26238 8213 26244
rect 8157 26188 8169 26238
rect 8169 26188 8213 26238
rect 5613 26114 5646 26164
rect 5646 26114 5660 26164
rect 5660 26114 5669 26164
rect 5696 26114 5712 26164
rect 5712 26114 5752 26164
rect 5613 26108 5669 26114
rect 5696 26108 5752 26114
rect 5779 26108 5835 26164
rect 5861 26108 5917 26164
rect 5943 26108 5999 26164
rect 6025 26108 6081 26164
rect 6107 26114 6148 26164
rect 6148 26114 6163 26164
rect 6189 26114 6200 26164
rect 6200 26114 6214 26164
rect 6214 26114 6245 26164
rect 6107 26108 6163 26114
rect 6189 26108 6245 26114
rect 6271 26108 6327 26164
rect 6353 26108 6409 26164
rect 6435 26108 6491 26164
rect 6517 26108 6573 26164
rect 6599 26108 6655 26164
rect 6681 26114 6702 26164
rect 6702 26114 6737 26164
rect 6763 26114 6768 26164
rect 6768 26114 6819 26164
rect 6681 26108 6737 26114
rect 6763 26108 6819 26114
rect 6845 26108 6901 26164
rect 6927 26108 6983 26164
rect 7009 26108 7065 26164
rect 7091 26108 7147 26164
rect 7173 26108 7229 26164
rect 7255 26114 7256 26164
rect 7256 26114 7308 26164
rect 7308 26114 7311 26164
rect 7337 26114 7374 26164
rect 7374 26114 7393 26164
rect 7255 26108 7311 26114
rect 7337 26108 7393 26114
rect 7419 26108 7475 26164
rect 7501 26108 7557 26164
rect 7583 26108 7639 26164
rect 7665 26108 7721 26164
rect 7747 26108 7803 26164
rect 7829 26114 7862 26164
rect 7862 26114 7876 26164
rect 7876 26114 7885 26164
rect 7911 26114 7928 26164
rect 7928 26114 7967 26164
rect 7829 26108 7885 26114
rect 7911 26108 7967 26114
rect 7993 26116 8047 26164
rect 8047 26116 8049 26164
rect 8075 26116 8099 26164
rect 8099 26116 8131 26164
rect 7993 26108 8049 26116
rect 8075 26108 8131 26116
rect 8157 26116 8169 26164
rect 8169 26116 8213 26164
rect 8157 26108 8213 26116
rect 2733 25931 2789 25987
rect 2814 25931 2870 25987
rect 2895 25931 2951 25987
rect 2976 25931 3032 25987
rect 3057 25931 3113 25987
rect 3138 25931 3194 25987
rect 3219 25931 3275 25987
rect 3300 25931 3356 25987
rect 3381 25931 3437 25987
rect 3462 25931 3518 25987
rect 3543 25931 3599 25987
rect 3624 25931 3680 25987
rect 3705 25931 3761 25987
rect 3786 25931 3842 25987
rect 3867 25931 3923 25987
rect 3948 25931 4004 25987
rect 4029 25931 4085 25987
rect 4110 25931 4166 25987
rect 4191 25931 4247 25987
rect 4272 25931 4328 25987
rect 4353 25931 4409 25987
rect 4434 25931 4490 25987
rect 4515 25931 4571 25987
rect 4596 25931 4652 25987
rect 4677 25931 4733 25987
rect 4758 25931 4814 25987
rect 4839 25931 4895 25987
rect 4920 25931 4976 25987
rect 5001 25931 5057 25987
rect 5082 25931 5138 25987
rect 2733 25851 2789 25907
rect 2814 25851 2870 25907
rect 2895 25851 2951 25907
rect 2976 25851 3032 25907
rect 3057 25851 3113 25907
rect 3138 25851 3194 25907
rect 3219 25851 3275 25907
rect 3300 25851 3356 25907
rect 3381 25851 3437 25907
rect 3462 25851 3518 25907
rect 3543 25851 3599 25907
rect 3624 25851 3680 25907
rect 3705 25851 3761 25907
rect 3786 25851 3842 25907
rect 3867 25851 3923 25907
rect 3948 25851 4004 25907
rect 4029 25851 4085 25907
rect 4110 25851 4166 25907
rect 4191 25851 4247 25907
rect 4272 25851 4328 25907
rect 4353 25851 4409 25907
rect 4434 25851 4490 25907
rect 4515 25851 4571 25907
rect 4596 25851 4652 25907
rect 4677 25851 4733 25907
rect 4758 25851 4814 25907
rect 4839 25851 4895 25907
rect 4920 25851 4976 25907
rect 5001 25851 5057 25907
rect 5082 25851 5138 25907
rect 2733 25771 2789 25827
rect 2814 25771 2870 25827
rect 2895 25771 2951 25827
rect 2976 25771 3032 25827
rect 3057 25771 3113 25827
rect 3138 25771 3194 25827
rect 3219 25771 3275 25827
rect 3300 25771 3356 25827
rect 3381 25771 3437 25827
rect 3462 25771 3518 25827
rect 3543 25771 3599 25827
rect 3624 25771 3680 25827
rect 3705 25771 3761 25827
rect 3786 25771 3842 25827
rect 3867 25771 3923 25827
rect 3948 25771 4004 25827
rect 4029 25771 4085 25827
rect 4110 25771 4166 25827
rect 4191 25771 4247 25827
rect 4272 25771 4328 25827
rect 4353 25771 4409 25827
rect 4434 25771 4490 25827
rect 4515 25771 4571 25827
rect 4596 25771 4652 25827
rect 4677 25771 4733 25827
rect 4758 25771 4814 25827
rect 4839 25771 4895 25827
rect 4920 25771 4976 25827
rect 5001 25771 5057 25827
rect 5082 25771 5138 25827
rect 2733 25691 2789 25747
rect 2814 25691 2870 25747
rect 2895 25691 2951 25747
rect 2976 25691 3032 25747
rect 3057 25691 3113 25747
rect 3138 25691 3194 25747
rect 3219 25691 3275 25747
rect 3300 25691 3356 25747
rect 3381 25691 3437 25747
rect 3462 25691 3518 25747
rect 3543 25691 3599 25747
rect 3624 25691 3680 25747
rect 3705 25691 3761 25747
rect 3786 25691 3842 25747
rect 3867 25691 3923 25747
rect 3948 25691 4004 25747
rect 4029 25691 4085 25747
rect 4110 25691 4166 25747
rect 4191 25691 4247 25747
rect 4272 25691 4328 25747
rect 4353 25691 4409 25747
rect 4434 25691 4490 25747
rect 4515 25691 4571 25747
rect 4596 25691 4652 25747
rect 4677 25691 4733 25747
rect 4758 25691 4814 25747
rect 4839 25691 4895 25747
rect 4920 25691 4976 25747
rect 5001 25691 5057 25747
rect 5082 25691 5138 25747
rect 2733 25611 2789 25667
rect 2814 25611 2870 25667
rect 2895 25611 2951 25667
rect 2976 25611 3032 25667
rect 3057 25611 3113 25667
rect 3138 25611 3194 25667
rect 3219 25611 3275 25667
rect 3300 25611 3356 25667
rect 3381 25611 3437 25667
rect 3462 25611 3518 25667
rect 3543 25611 3599 25667
rect 3624 25611 3680 25667
rect 3705 25611 3761 25667
rect 3786 25611 3842 25667
rect 3867 25611 3923 25667
rect 3948 25611 4004 25667
rect 4029 25611 4085 25667
rect 4110 25611 4166 25667
rect 4191 25611 4247 25667
rect 4272 25611 4328 25667
rect 4353 25611 4409 25667
rect 4434 25611 4490 25667
rect 4515 25611 4571 25667
rect 4596 25611 4652 25667
rect 4677 25611 4733 25667
rect 4758 25611 4814 25667
rect 4839 25611 4895 25667
rect 4920 25611 4976 25667
rect 5001 25611 5057 25667
rect 5082 25611 5138 25667
rect 2733 25531 2789 25587
rect 2814 25531 2870 25587
rect 2895 25531 2951 25587
rect 2976 25531 3032 25587
rect 3057 25531 3113 25587
rect 3138 25531 3194 25587
rect 3219 25531 3275 25587
rect 3300 25531 3356 25587
rect 3381 25531 3437 25587
rect 3462 25531 3518 25587
rect 3543 25531 3599 25587
rect 3624 25531 3680 25587
rect 3705 25531 3761 25587
rect 3786 25531 3842 25587
rect 3867 25531 3923 25587
rect 3948 25531 4004 25587
rect 4029 25531 4085 25587
rect 4110 25531 4166 25587
rect 4191 25531 4247 25587
rect 4272 25531 4328 25587
rect 4353 25531 4409 25587
rect 4434 25531 4490 25587
rect 4515 25531 4571 25587
rect 4596 25531 4652 25587
rect 4677 25531 4733 25587
rect 4758 25531 4814 25587
rect 4839 25531 4895 25587
rect 4920 25531 4976 25587
rect 5001 25531 5057 25587
rect 5082 25531 5138 25587
rect 2733 25451 2789 25507
rect 2814 25451 2870 25507
rect 2895 25451 2951 25507
rect 2976 25451 3032 25507
rect 3057 25451 3113 25507
rect 3138 25451 3194 25507
rect 3219 25451 3275 25507
rect 3300 25451 3356 25507
rect 3381 25451 3437 25507
rect 3462 25451 3518 25507
rect 3543 25451 3599 25507
rect 3624 25451 3680 25507
rect 3705 25451 3761 25507
rect 3786 25451 3842 25507
rect 3867 25451 3923 25507
rect 3948 25451 4004 25507
rect 4029 25451 4085 25507
rect 4110 25451 4166 25507
rect 4191 25451 4247 25507
rect 4272 25451 4328 25507
rect 4353 25451 4409 25507
rect 4434 25451 4490 25507
rect 4515 25451 4571 25507
rect 4596 25451 4652 25507
rect 4677 25451 4733 25507
rect 4758 25451 4814 25507
rect 4839 25451 4895 25507
rect 4920 25451 4976 25507
rect 5001 25451 5057 25507
rect 5082 25451 5138 25507
rect 2733 25371 2789 25427
rect 2814 25371 2870 25427
rect 2895 25371 2951 25427
rect 2976 25371 3032 25427
rect 3057 25371 3113 25427
rect 3138 25371 3194 25427
rect 3219 25371 3275 25427
rect 3300 25371 3356 25427
rect 3381 25371 3437 25427
rect 3462 25371 3518 25427
rect 3543 25371 3599 25427
rect 3624 25371 3680 25427
rect 3705 25371 3761 25427
rect 3786 25371 3842 25427
rect 3867 25371 3923 25427
rect 3948 25371 4004 25427
rect 4029 25371 4085 25427
rect 4110 25371 4166 25427
rect 4191 25371 4247 25427
rect 4272 25371 4328 25427
rect 4353 25371 4409 25427
rect 4434 25371 4490 25427
rect 4515 25371 4571 25427
rect 4596 25371 4652 25427
rect 4677 25371 4733 25427
rect 4758 25371 4814 25427
rect 4839 25371 4895 25427
rect 4920 25371 4976 25427
rect 5001 25371 5057 25427
rect 5082 25371 5138 25427
rect 5163 25371 5299 25987
rect 5613 24720 5669 24724
rect 5696 24720 5752 24724
rect 5613 24668 5646 24720
rect 5646 24668 5660 24720
rect 5660 24668 5669 24720
rect 5696 24668 5712 24720
rect 5712 24668 5752 24720
rect 5779 24668 5835 24724
rect 5861 24668 5917 24724
rect 5943 24668 5999 24724
rect 6025 24668 6081 24724
rect 6107 24720 6163 24724
rect 6189 24720 6245 24724
rect 6107 24668 6148 24720
rect 6148 24668 6163 24720
rect 6189 24668 6200 24720
rect 6200 24668 6214 24720
rect 6214 24668 6245 24720
rect 6271 24668 6327 24724
rect 6353 24668 6409 24724
rect 6435 24668 6491 24724
rect 6517 24668 6573 24724
rect 6599 24668 6655 24724
rect 6681 24720 6737 24724
rect 6763 24720 6819 24724
rect 6681 24668 6702 24720
rect 6702 24668 6737 24720
rect 6763 24668 6768 24720
rect 6768 24668 6819 24720
rect 6845 24668 6901 24724
rect 6927 24668 6983 24724
rect 7009 24668 7065 24724
rect 7091 24668 7147 24724
rect 7173 24668 7229 24724
rect 7255 24720 7311 24724
rect 7337 24720 7393 24724
rect 7255 24668 7256 24720
rect 7256 24668 7308 24720
rect 7308 24668 7311 24720
rect 7337 24668 7374 24720
rect 7374 24668 7393 24720
rect 7419 24668 7475 24724
rect 7501 24668 7557 24724
rect 7583 24668 7639 24724
rect 7665 24668 7721 24724
rect 7747 24668 7803 24724
rect 7829 24720 7885 24724
rect 7911 24720 7967 24724
rect 7829 24668 7862 24720
rect 7862 24668 7876 24720
rect 7876 24668 7885 24720
rect 7911 24668 7928 24720
rect 7928 24668 7967 24720
rect 7993 24672 8047 24724
rect 8047 24672 8049 24724
rect 8075 24672 8099 24724
rect 8099 24672 8131 24724
rect 7993 24668 8049 24672
rect 8075 24668 8131 24672
rect 8157 24672 8169 24724
rect 8169 24672 8213 24724
rect 8157 24668 8213 24672
rect 5613 24599 5646 24644
rect 5646 24599 5660 24644
rect 5660 24599 5669 24644
rect 5696 24599 5712 24644
rect 5712 24599 5752 24644
rect 5613 24588 5669 24599
rect 5696 24588 5752 24599
rect 5779 24588 5835 24644
rect 5861 24588 5917 24644
rect 5943 24588 5999 24644
rect 6025 24588 6081 24644
rect 6107 24599 6148 24644
rect 6148 24599 6163 24644
rect 6189 24599 6200 24644
rect 6200 24599 6214 24644
rect 6214 24599 6245 24644
rect 6107 24588 6163 24599
rect 6189 24588 6245 24599
rect 6271 24588 6327 24644
rect 6353 24588 6409 24644
rect 6435 24588 6491 24644
rect 6517 24588 6573 24644
rect 6599 24588 6655 24644
rect 6681 24599 6702 24644
rect 6702 24599 6737 24644
rect 6763 24599 6768 24644
rect 6768 24599 6819 24644
rect 6681 24588 6737 24599
rect 6763 24588 6819 24599
rect 6845 24588 6901 24644
rect 6927 24588 6983 24644
rect 7009 24588 7065 24644
rect 7091 24588 7147 24644
rect 7173 24588 7229 24644
rect 7255 24599 7256 24644
rect 7256 24599 7308 24644
rect 7308 24599 7311 24644
rect 7337 24599 7374 24644
rect 7374 24599 7393 24644
rect 7255 24588 7311 24599
rect 7337 24588 7393 24599
rect 7419 24588 7475 24644
rect 7501 24588 7557 24644
rect 7583 24588 7639 24644
rect 7665 24588 7721 24644
rect 7747 24588 7803 24644
rect 7829 24599 7862 24644
rect 7862 24599 7876 24644
rect 7876 24599 7885 24644
rect 7911 24599 7928 24644
rect 7928 24599 7967 24644
rect 7829 24588 7885 24599
rect 7911 24588 7967 24599
rect 7993 24603 8047 24644
rect 8047 24603 8049 24644
rect 8075 24603 8099 24644
rect 8099 24603 8131 24644
rect 7993 24588 8049 24603
rect 8075 24588 8131 24603
rect 8157 24603 8169 24644
rect 8169 24603 8213 24644
rect 8157 24588 8213 24603
rect 5613 24530 5646 24564
rect 5646 24530 5660 24564
rect 5660 24530 5669 24564
rect 5696 24530 5712 24564
rect 5712 24530 5752 24564
rect 5613 24513 5669 24530
rect 5696 24513 5752 24530
rect 5613 24508 5646 24513
rect 5646 24508 5660 24513
rect 5660 24508 5669 24513
rect 5696 24508 5712 24513
rect 5712 24508 5752 24513
rect 5779 24508 5835 24564
rect 5861 24508 5917 24564
rect 5943 24508 5999 24564
rect 6025 24508 6081 24564
rect 6107 24530 6148 24564
rect 6148 24530 6163 24564
rect 6189 24530 6200 24564
rect 6200 24530 6214 24564
rect 6214 24530 6245 24564
rect 6107 24513 6163 24530
rect 6189 24513 6245 24530
rect 6107 24508 6148 24513
rect 6148 24508 6163 24513
rect 6189 24508 6200 24513
rect 6200 24508 6214 24513
rect 6214 24508 6245 24513
rect 6271 24508 6327 24564
rect 6353 24508 6409 24564
rect 6435 24508 6491 24564
rect 6517 24508 6573 24564
rect 6599 24508 6655 24564
rect 6681 24530 6702 24564
rect 6702 24530 6737 24564
rect 6763 24530 6768 24564
rect 6768 24530 6819 24564
rect 6681 24513 6737 24530
rect 6763 24513 6819 24530
rect 6681 24508 6702 24513
rect 6702 24508 6737 24513
rect 6763 24508 6768 24513
rect 6768 24508 6819 24513
rect 6845 24508 6901 24564
rect 6927 24508 6983 24564
rect 7009 24508 7065 24564
rect 7091 24508 7147 24564
rect 7173 24508 7229 24564
rect 7255 24530 7256 24564
rect 7256 24530 7308 24564
rect 7308 24530 7311 24564
rect 7337 24530 7374 24564
rect 7374 24530 7393 24564
rect 7255 24513 7311 24530
rect 7337 24513 7393 24530
rect 7255 24508 7256 24513
rect 7256 24508 7308 24513
rect 7308 24508 7311 24513
rect 7337 24508 7374 24513
rect 7374 24508 7393 24513
rect 7419 24508 7475 24564
rect 7501 24508 7557 24564
rect 7583 24508 7639 24564
rect 7665 24508 7721 24564
rect 7747 24508 7803 24564
rect 7829 24530 7862 24564
rect 7862 24530 7876 24564
rect 7876 24530 7885 24564
rect 7911 24530 7928 24564
rect 7928 24530 7967 24564
rect 7829 24513 7885 24530
rect 7911 24513 7967 24530
rect 7829 24508 7862 24513
rect 7862 24508 7876 24513
rect 7876 24508 7885 24513
rect 7911 24508 7928 24513
rect 7928 24508 7967 24513
rect 7993 24534 8047 24564
rect 8047 24534 8049 24564
rect 8075 24534 8099 24564
rect 8099 24534 8131 24564
rect 7993 24517 8049 24534
rect 8075 24517 8131 24534
rect 7993 24508 8047 24517
rect 8047 24508 8049 24517
rect 8075 24508 8099 24517
rect 8099 24508 8131 24517
rect 8157 24534 8169 24564
rect 8169 24534 8213 24564
rect 8157 24517 8213 24534
rect 8157 24508 8169 24517
rect 8169 24508 8213 24517
rect 5613 24461 5646 24484
rect 5646 24461 5660 24484
rect 5660 24461 5669 24484
rect 5696 24461 5712 24484
rect 5712 24461 5752 24484
rect 5613 24444 5669 24461
rect 5696 24444 5752 24461
rect 5613 24428 5646 24444
rect 5646 24428 5660 24444
rect 5660 24428 5669 24444
rect 5696 24428 5712 24444
rect 5712 24428 5752 24444
rect 5779 24428 5835 24484
rect 5861 24428 5917 24484
rect 5943 24428 5999 24484
rect 6025 24428 6081 24484
rect 6107 24461 6148 24484
rect 6148 24461 6163 24484
rect 6189 24461 6200 24484
rect 6200 24461 6214 24484
rect 6214 24461 6245 24484
rect 6107 24444 6163 24461
rect 6189 24444 6245 24461
rect 6107 24428 6148 24444
rect 6148 24428 6163 24444
rect 6189 24428 6200 24444
rect 6200 24428 6214 24444
rect 6214 24428 6245 24444
rect 6271 24428 6327 24484
rect 6353 24428 6409 24484
rect 6435 24428 6491 24484
rect 6517 24428 6573 24484
rect 6599 24428 6655 24484
rect 6681 24461 6702 24484
rect 6702 24461 6737 24484
rect 6763 24461 6768 24484
rect 6768 24461 6819 24484
rect 6681 24444 6737 24461
rect 6763 24444 6819 24461
rect 6681 24428 6702 24444
rect 6702 24428 6737 24444
rect 6763 24428 6768 24444
rect 6768 24428 6819 24444
rect 6845 24428 6901 24484
rect 6927 24428 6983 24484
rect 7009 24428 7065 24484
rect 7091 24428 7147 24484
rect 7173 24428 7229 24484
rect 7255 24461 7256 24484
rect 7256 24461 7308 24484
rect 7308 24461 7311 24484
rect 7337 24461 7374 24484
rect 7374 24461 7393 24484
rect 7255 24444 7311 24461
rect 7337 24444 7393 24461
rect 7255 24428 7256 24444
rect 7256 24428 7308 24444
rect 7308 24428 7311 24444
rect 7337 24428 7374 24444
rect 7374 24428 7393 24444
rect 7419 24428 7475 24484
rect 7501 24428 7557 24484
rect 7583 24428 7639 24484
rect 7665 24428 7721 24484
rect 7747 24428 7803 24484
rect 7829 24461 7862 24484
rect 7862 24461 7876 24484
rect 7876 24461 7885 24484
rect 7911 24461 7928 24484
rect 7928 24461 7967 24484
rect 7829 24444 7885 24461
rect 7911 24444 7967 24461
rect 7829 24428 7862 24444
rect 7862 24428 7876 24444
rect 7876 24428 7885 24444
rect 7911 24428 7928 24444
rect 7928 24428 7967 24444
rect 7993 24465 8047 24484
rect 8047 24465 8049 24484
rect 8075 24465 8099 24484
rect 8099 24465 8131 24484
rect 7993 24448 8049 24465
rect 8075 24448 8131 24465
rect 7993 24428 8047 24448
rect 8047 24428 8049 24448
rect 8075 24428 8099 24448
rect 8099 24428 8131 24448
rect 8157 24465 8169 24484
rect 8169 24465 8213 24484
rect 8157 24448 8213 24465
rect 8157 24428 8169 24448
rect 8169 24428 8213 24448
rect 5613 24392 5646 24404
rect 5646 24392 5660 24404
rect 5660 24392 5669 24404
rect 5696 24392 5712 24404
rect 5712 24392 5752 24404
rect 5613 24375 5669 24392
rect 5696 24375 5752 24392
rect 5613 24348 5646 24375
rect 5646 24348 5660 24375
rect 5660 24348 5669 24375
rect 5696 24348 5712 24375
rect 5712 24348 5752 24375
rect 5779 24348 5835 24404
rect 5861 24348 5917 24404
rect 5943 24348 5999 24404
rect 6025 24348 6081 24404
rect 6107 24392 6148 24404
rect 6148 24392 6163 24404
rect 6189 24392 6200 24404
rect 6200 24392 6214 24404
rect 6214 24392 6245 24404
rect 6107 24375 6163 24392
rect 6189 24375 6245 24392
rect 6107 24348 6148 24375
rect 6148 24348 6163 24375
rect 6189 24348 6200 24375
rect 6200 24348 6214 24375
rect 6214 24348 6245 24375
rect 6271 24348 6327 24404
rect 6353 24348 6409 24404
rect 6435 24348 6491 24404
rect 6517 24348 6573 24404
rect 6599 24348 6655 24404
rect 6681 24392 6702 24404
rect 6702 24392 6737 24404
rect 6763 24392 6768 24404
rect 6768 24392 6819 24404
rect 6681 24375 6737 24392
rect 6763 24375 6819 24392
rect 6681 24348 6702 24375
rect 6702 24348 6737 24375
rect 6763 24348 6768 24375
rect 6768 24348 6819 24375
rect 6845 24348 6901 24404
rect 6927 24348 6983 24404
rect 7009 24348 7065 24404
rect 7091 24348 7147 24404
rect 7173 24348 7229 24404
rect 7255 24392 7256 24404
rect 7256 24392 7308 24404
rect 7308 24392 7311 24404
rect 7337 24392 7374 24404
rect 7374 24392 7393 24404
rect 7255 24375 7311 24392
rect 7337 24375 7393 24392
rect 7255 24348 7256 24375
rect 7256 24348 7308 24375
rect 7308 24348 7311 24375
rect 7337 24348 7374 24375
rect 7374 24348 7393 24375
rect 7419 24348 7475 24404
rect 7501 24348 7557 24404
rect 7583 24348 7639 24404
rect 7665 24348 7721 24404
rect 7747 24348 7803 24404
rect 7829 24392 7862 24404
rect 7862 24392 7876 24404
rect 7876 24392 7885 24404
rect 7911 24392 7928 24404
rect 7928 24392 7967 24404
rect 7829 24375 7885 24392
rect 7911 24375 7967 24392
rect 7829 24348 7862 24375
rect 7862 24348 7876 24375
rect 7876 24348 7885 24375
rect 7911 24348 7928 24375
rect 7928 24348 7967 24375
rect 7993 24396 8047 24404
rect 8047 24396 8049 24404
rect 8075 24396 8099 24404
rect 8099 24396 8131 24404
rect 7993 24378 8049 24396
rect 8075 24378 8131 24396
rect 7993 24348 8047 24378
rect 8047 24348 8049 24378
rect 8075 24348 8099 24378
rect 8099 24348 8131 24378
rect 8157 24396 8169 24404
rect 8169 24396 8213 24404
rect 8157 24378 8213 24396
rect 8157 24348 8169 24378
rect 8169 24348 8213 24378
rect 5613 24323 5646 24324
rect 5646 24323 5660 24324
rect 5660 24323 5669 24324
rect 5696 24323 5712 24324
rect 5712 24323 5752 24324
rect 5613 24306 5669 24323
rect 5696 24306 5752 24323
rect 5613 24268 5646 24306
rect 5646 24268 5660 24306
rect 5660 24268 5669 24306
rect 5696 24268 5712 24306
rect 5712 24268 5752 24306
rect 5779 24268 5835 24324
rect 5861 24268 5917 24324
rect 5943 24268 5999 24324
rect 6025 24268 6081 24324
rect 6107 24323 6148 24324
rect 6148 24323 6163 24324
rect 6189 24323 6200 24324
rect 6200 24323 6214 24324
rect 6214 24323 6245 24324
rect 6107 24306 6163 24323
rect 6189 24306 6245 24323
rect 6107 24268 6148 24306
rect 6148 24268 6163 24306
rect 6189 24268 6200 24306
rect 6200 24268 6214 24306
rect 6214 24268 6245 24306
rect 6271 24268 6327 24324
rect 6353 24268 6409 24324
rect 6435 24268 6491 24324
rect 6517 24268 6573 24324
rect 6599 24268 6655 24324
rect 6681 24323 6702 24324
rect 6702 24323 6737 24324
rect 6763 24323 6768 24324
rect 6768 24323 6819 24324
rect 6681 24306 6737 24323
rect 6763 24306 6819 24323
rect 6681 24268 6702 24306
rect 6702 24268 6737 24306
rect 6763 24268 6768 24306
rect 6768 24268 6819 24306
rect 6845 24268 6901 24324
rect 6927 24268 6983 24324
rect 7009 24268 7065 24324
rect 7091 24268 7147 24324
rect 7173 24268 7229 24324
rect 7255 24323 7256 24324
rect 7256 24323 7308 24324
rect 7308 24323 7311 24324
rect 7337 24323 7374 24324
rect 7374 24323 7393 24324
rect 7255 24306 7311 24323
rect 7337 24306 7393 24323
rect 7255 24268 7256 24306
rect 7256 24268 7308 24306
rect 7308 24268 7311 24306
rect 7337 24268 7374 24306
rect 7374 24268 7393 24306
rect 7419 24268 7475 24324
rect 7501 24268 7557 24324
rect 7583 24268 7639 24324
rect 7665 24268 7721 24324
rect 7747 24268 7803 24324
rect 7829 24323 7862 24324
rect 7862 24323 7876 24324
rect 7876 24323 7885 24324
rect 7911 24323 7928 24324
rect 7928 24323 7967 24324
rect 7829 24306 7885 24323
rect 7911 24306 7967 24323
rect 7829 24268 7862 24306
rect 7862 24268 7876 24306
rect 7876 24268 7885 24306
rect 7911 24268 7928 24306
rect 7928 24268 7967 24306
rect 7993 24308 8049 24324
rect 8075 24308 8131 24324
rect 7993 24268 8047 24308
rect 8047 24268 8049 24308
rect 8075 24268 8099 24308
rect 8099 24268 8131 24308
rect 8157 24308 8213 24324
rect 8157 24268 8169 24308
rect 8169 24268 8213 24308
rect 5613 24236 5669 24244
rect 5696 24236 5752 24244
rect 5613 24188 5646 24236
rect 5646 24188 5660 24236
rect 5660 24188 5669 24236
rect 5696 24188 5712 24236
rect 5712 24188 5752 24236
rect 5779 24188 5835 24244
rect 5861 24188 5917 24244
rect 5943 24188 5999 24244
rect 6025 24188 6081 24244
rect 6107 24236 6163 24244
rect 6189 24236 6245 24244
rect 6107 24188 6148 24236
rect 6148 24188 6163 24236
rect 6189 24188 6200 24236
rect 6200 24188 6214 24236
rect 6214 24188 6245 24236
rect 6271 24188 6327 24244
rect 6353 24188 6409 24244
rect 6435 24188 6491 24244
rect 6517 24188 6573 24244
rect 6599 24188 6655 24244
rect 6681 24236 6737 24244
rect 6763 24236 6819 24244
rect 6681 24188 6702 24236
rect 6702 24188 6737 24236
rect 6763 24188 6768 24236
rect 6768 24188 6819 24236
rect 6845 24188 6901 24244
rect 6927 24188 6983 24244
rect 7009 24188 7065 24244
rect 7091 24188 7147 24244
rect 7173 24188 7229 24244
rect 7255 24236 7311 24244
rect 7337 24236 7393 24244
rect 7255 24188 7256 24236
rect 7256 24188 7308 24236
rect 7308 24188 7311 24236
rect 7337 24188 7374 24236
rect 7374 24188 7393 24236
rect 7419 24188 7475 24244
rect 7501 24188 7557 24244
rect 7583 24188 7639 24244
rect 7665 24188 7721 24244
rect 7747 24188 7803 24244
rect 7829 24236 7885 24244
rect 7911 24236 7967 24244
rect 7829 24188 7862 24236
rect 7862 24188 7876 24236
rect 7876 24188 7885 24236
rect 7911 24188 7928 24236
rect 7928 24188 7967 24236
rect 7993 24238 8049 24244
rect 8075 24238 8131 24244
rect 7993 24188 8047 24238
rect 8047 24188 8049 24238
rect 8075 24188 8099 24238
rect 8099 24188 8131 24238
rect 8157 24238 8213 24244
rect 8157 24188 8169 24238
rect 8169 24188 8213 24238
rect 5613 24114 5646 24164
rect 5646 24114 5660 24164
rect 5660 24114 5669 24164
rect 5696 24114 5712 24164
rect 5712 24114 5752 24164
rect 5613 24108 5669 24114
rect 5696 24108 5752 24114
rect 5779 24108 5835 24164
rect 5861 24108 5917 24164
rect 5943 24108 5999 24164
rect 6025 24108 6081 24164
rect 6107 24114 6148 24164
rect 6148 24114 6163 24164
rect 6189 24114 6200 24164
rect 6200 24114 6214 24164
rect 6214 24114 6245 24164
rect 6107 24108 6163 24114
rect 6189 24108 6245 24114
rect 6271 24108 6327 24164
rect 6353 24108 6409 24164
rect 6435 24108 6491 24164
rect 6517 24108 6573 24164
rect 6599 24108 6655 24164
rect 6681 24114 6702 24164
rect 6702 24114 6737 24164
rect 6763 24114 6768 24164
rect 6768 24114 6819 24164
rect 6681 24108 6737 24114
rect 6763 24108 6819 24114
rect 6845 24108 6901 24164
rect 6927 24108 6983 24164
rect 7009 24108 7065 24164
rect 7091 24108 7147 24164
rect 7173 24108 7229 24164
rect 7255 24114 7256 24164
rect 7256 24114 7308 24164
rect 7308 24114 7311 24164
rect 7337 24114 7374 24164
rect 7374 24114 7393 24164
rect 7255 24108 7311 24114
rect 7337 24108 7393 24114
rect 7419 24108 7475 24164
rect 7501 24108 7557 24164
rect 7583 24108 7639 24164
rect 7665 24108 7721 24164
rect 7747 24108 7803 24164
rect 7829 24114 7862 24164
rect 7862 24114 7876 24164
rect 7876 24114 7885 24164
rect 7911 24114 7928 24164
rect 7928 24114 7967 24164
rect 7829 24108 7885 24114
rect 7911 24108 7967 24114
rect 7993 24116 8047 24164
rect 8047 24116 8049 24164
rect 8075 24116 8099 24164
rect 8099 24116 8131 24164
rect 7993 24108 8049 24116
rect 8075 24108 8131 24116
rect 8157 24116 8169 24164
rect 8169 24116 8213 24164
rect 8157 24108 8213 24116
rect 2733 23931 2789 23987
rect 2814 23931 2870 23987
rect 2895 23931 2951 23987
rect 2976 23931 3032 23987
rect 3057 23931 3113 23987
rect 3138 23931 3194 23987
rect 3219 23931 3275 23987
rect 3300 23931 3356 23987
rect 3381 23931 3437 23987
rect 3462 23931 3518 23987
rect 3543 23931 3599 23987
rect 3624 23931 3680 23987
rect 3705 23931 3761 23987
rect 3786 23931 3842 23987
rect 3867 23931 3923 23987
rect 3948 23931 4004 23987
rect 4029 23931 4085 23987
rect 4110 23931 4166 23987
rect 4191 23931 4247 23987
rect 4272 23931 4328 23987
rect 4353 23931 4409 23987
rect 4434 23931 4490 23987
rect 4515 23931 4571 23987
rect 4596 23931 4652 23987
rect 4677 23931 4733 23987
rect 4758 23931 4814 23987
rect 4839 23931 4895 23987
rect 4920 23931 4976 23987
rect 5001 23931 5057 23987
rect 5082 23931 5138 23987
rect 2733 23851 2789 23907
rect 2814 23851 2870 23907
rect 2895 23851 2951 23907
rect 2976 23851 3032 23907
rect 3057 23851 3113 23907
rect 3138 23851 3194 23907
rect 3219 23851 3275 23907
rect 3300 23851 3356 23907
rect 3381 23851 3437 23907
rect 3462 23851 3518 23907
rect 3543 23851 3599 23907
rect 3624 23851 3680 23907
rect 3705 23851 3761 23907
rect 3786 23851 3842 23907
rect 3867 23851 3923 23907
rect 3948 23851 4004 23907
rect 4029 23851 4085 23907
rect 4110 23851 4166 23907
rect 4191 23851 4247 23907
rect 4272 23851 4328 23907
rect 4353 23851 4409 23907
rect 4434 23851 4490 23907
rect 4515 23851 4571 23907
rect 4596 23851 4652 23907
rect 4677 23851 4733 23907
rect 4758 23851 4814 23907
rect 4839 23851 4895 23907
rect 4920 23851 4976 23907
rect 5001 23851 5057 23907
rect 5082 23851 5138 23907
rect 2733 23771 2789 23827
rect 2814 23771 2870 23827
rect 2895 23771 2951 23827
rect 2976 23771 3032 23827
rect 3057 23771 3113 23827
rect 3138 23771 3194 23827
rect 3219 23771 3275 23827
rect 3300 23771 3356 23827
rect 3381 23771 3437 23827
rect 3462 23771 3518 23827
rect 3543 23771 3599 23827
rect 3624 23771 3680 23827
rect 3705 23771 3761 23827
rect 3786 23771 3842 23827
rect 3867 23771 3923 23827
rect 3948 23771 4004 23827
rect 4029 23771 4085 23827
rect 4110 23771 4166 23827
rect 4191 23771 4247 23827
rect 4272 23771 4328 23827
rect 4353 23771 4409 23827
rect 4434 23771 4490 23827
rect 4515 23771 4571 23827
rect 4596 23771 4652 23827
rect 4677 23771 4733 23827
rect 4758 23771 4814 23827
rect 4839 23771 4895 23827
rect 4920 23771 4976 23827
rect 5001 23771 5057 23827
rect 5082 23771 5138 23827
rect 2733 23691 2789 23747
rect 2814 23691 2870 23747
rect 2895 23691 2951 23747
rect 2976 23691 3032 23747
rect 3057 23691 3113 23747
rect 3138 23691 3194 23747
rect 3219 23691 3275 23747
rect 3300 23691 3356 23747
rect 3381 23691 3437 23747
rect 3462 23691 3518 23747
rect 3543 23691 3599 23747
rect 3624 23691 3680 23747
rect 3705 23691 3761 23747
rect 3786 23691 3842 23747
rect 3867 23691 3923 23747
rect 3948 23691 4004 23747
rect 4029 23691 4085 23747
rect 4110 23691 4166 23747
rect 4191 23691 4247 23747
rect 4272 23691 4328 23747
rect 4353 23691 4409 23747
rect 4434 23691 4490 23747
rect 4515 23691 4571 23747
rect 4596 23691 4652 23747
rect 4677 23691 4733 23747
rect 4758 23691 4814 23747
rect 4839 23691 4895 23747
rect 4920 23691 4976 23747
rect 5001 23691 5057 23747
rect 5082 23691 5138 23747
rect 2733 23611 2789 23667
rect 2814 23611 2870 23667
rect 2895 23611 2951 23667
rect 2976 23611 3032 23667
rect 3057 23611 3113 23667
rect 3138 23611 3194 23667
rect 3219 23611 3275 23667
rect 3300 23611 3356 23667
rect 3381 23611 3437 23667
rect 3462 23611 3518 23667
rect 3543 23611 3599 23667
rect 3624 23611 3680 23667
rect 3705 23611 3761 23667
rect 3786 23611 3842 23667
rect 3867 23611 3923 23667
rect 3948 23611 4004 23667
rect 4029 23611 4085 23667
rect 4110 23611 4166 23667
rect 4191 23611 4247 23667
rect 4272 23611 4328 23667
rect 4353 23611 4409 23667
rect 4434 23611 4490 23667
rect 4515 23611 4571 23667
rect 4596 23611 4652 23667
rect 4677 23611 4733 23667
rect 4758 23611 4814 23667
rect 4839 23611 4895 23667
rect 4920 23611 4976 23667
rect 5001 23611 5057 23667
rect 5082 23611 5138 23667
rect 2733 23531 2789 23587
rect 2814 23531 2870 23587
rect 2895 23531 2951 23587
rect 2976 23531 3032 23587
rect 3057 23531 3113 23587
rect 3138 23531 3194 23587
rect 3219 23531 3275 23587
rect 3300 23531 3356 23587
rect 3381 23531 3437 23587
rect 3462 23531 3518 23587
rect 3543 23531 3599 23587
rect 3624 23531 3680 23587
rect 3705 23531 3761 23587
rect 3786 23531 3842 23587
rect 3867 23531 3923 23587
rect 3948 23531 4004 23587
rect 4029 23531 4085 23587
rect 4110 23531 4166 23587
rect 4191 23531 4247 23587
rect 4272 23531 4328 23587
rect 4353 23531 4409 23587
rect 4434 23531 4490 23587
rect 4515 23531 4571 23587
rect 4596 23531 4652 23587
rect 4677 23531 4733 23587
rect 4758 23531 4814 23587
rect 4839 23531 4895 23587
rect 4920 23531 4976 23587
rect 5001 23531 5057 23587
rect 5082 23531 5138 23587
rect 2733 23451 2789 23507
rect 2814 23451 2870 23507
rect 2895 23451 2951 23507
rect 2976 23451 3032 23507
rect 3057 23451 3113 23507
rect 3138 23451 3194 23507
rect 3219 23451 3275 23507
rect 3300 23451 3356 23507
rect 3381 23451 3437 23507
rect 3462 23451 3518 23507
rect 3543 23451 3599 23507
rect 3624 23451 3680 23507
rect 3705 23451 3761 23507
rect 3786 23451 3842 23507
rect 3867 23451 3923 23507
rect 3948 23451 4004 23507
rect 4029 23451 4085 23507
rect 4110 23451 4166 23507
rect 4191 23451 4247 23507
rect 4272 23451 4328 23507
rect 4353 23451 4409 23507
rect 4434 23451 4490 23507
rect 4515 23451 4571 23507
rect 4596 23451 4652 23507
rect 4677 23451 4733 23507
rect 4758 23451 4814 23507
rect 4839 23451 4895 23507
rect 4920 23451 4976 23507
rect 5001 23451 5057 23507
rect 5082 23451 5138 23507
rect 2733 23371 2789 23427
rect 2814 23371 2870 23427
rect 2895 23371 2951 23427
rect 2976 23371 3032 23427
rect 3057 23371 3113 23427
rect 3138 23371 3194 23427
rect 3219 23371 3275 23427
rect 3300 23371 3356 23427
rect 3381 23371 3437 23427
rect 3462 23371 3518 23427
rect 3543 23371 3599 23427
rect 3624 23371 3680 23427
rect 3705 23371 3761 23427
rect 3786 23371 3842 23427
rect 3867 23371 3923 23427
rect 3948 23371 4004 23427
rect 4029 23371 4085 23427
rect 4110 23371 4166 23427
rect 4191 23371 4247 23427
rect 4272 23371 4328 23427
rect 4353 23371 4409 23427
rect 4434 23371 4490 23427
rect 4515 23371 4571 23427
rect 4596 23371 4652 23427
rect 4677 23371 4733 23427
rect 4758 23371 4814 23427
rect 4839 23371 4895 23427
rect 4920 23371 4976 23427
rect 5001 23371 5057 23427
rect 5082 23371 5138 23427
rect 5163 23371 5299 23987
rect 5613 22720 5669 22724
rect 5696 22720 5752 22724
rect 5613 22668 5646 22720
rect 5646 22668 5660 22720
rect 5660 22668 5669 22720
rect 5696 22668 5712 22720
rect 5712 22668 5752 22720
rect 5779 22668 5835 22724
rect 5861 22668 5917 22724
rect 5943 22668 5999 22724
rect 6025 22668 6081 22724
rect 6107 22720 6163 22724
rect 6189 22720 6245 22724
rect 6107 22668 6148 22720
rect 6148 22668 6163 22720
rect 6189 22668 6200 22720
rect 6200 22668 6214 22720
rect 6214 22668 6245 22720
rect 6271 22668 6327 22724
rect 6353 22668 6409 22724
rect 6435 22668 6491 22724
rect 6517 22668 6573 22724
rect 6599 22668 6655 22724
rect 6681 22720 6737 22724
rect 6763 22720 6819 22724
rect 6681 22668 6702 22720
rect 6702 22668 6737 22720
rect 6763 22668 6768 22720
rect 6768 22668 6819 22720
rect 6845 22668 6901 22724
rect 6927 22668 6983 22724
rect 7009 22668 7065 22724
rect 7091 22668 7147 22724
rect 7173 22668 7229 22724
rect 7255 22720 7311 22724
rect 7337 22720 7393 22724
rect 7255 22668 7256 22720
rect 7256 22668 7308 22720
rect 7308 22668 7311 22720
rect 7337 22668 7374 22720
rect 7374 22668 7393 22720
rect 7419 22668 7475 22724
rect 7501 22668 7557 22724
rect 7583 22668 7639 22724
rect 7665 22668 7721 22724
rect 7747 22668 7803 22724
rect 7829 22720 7885 22724
rect 7911 22720 7967 22724
rect 7829 22668 7862 22720
rect 7862 22668 7876 22720
rect 7876 22668 7885 22720
rect 7911 22668 7928 22720
rect 7928 22668 7967 22720
rect 7993 22672 8047 22724
rect 8047 22672 8049 22724
rect 8075 22672 8099 22724
rect 8099 22672 8131 22724
rect 7993 22668 8049 22672
rect 8075 22668 8131 22672
rect 8157 22672 8169 22724
rect 8169 22672 8213 22724
rect 8157 22668 8213 22672
rect 5613 22599 5646 22644
rect 5646 22599 5660 22644
rect 5660 22599 5669 22644
rect 5696 22599 5712 22644
rect 5712 22599 5752 22644
rect 5613 22588 5669 22599
rect 5696 22588 5752 22599
rect 5779 22588 5835 22644
rect 5861 22588 5917 22644
rect 5943 22588 5999 22644
rect 6025 22588 6081 22644
rect 6107 22599 6148 22644
rect 6148 22599 6163 22644
rect 6189 22599 6200 22644
rect 6200 22599 6214 22644
rect 6214 22599 6245 22644
rect 6107 22588 6163 22599
rect 6189 22588 6245 22599
rect 6271 22588 6327 22644
rect 6353 22588 6409 22644
rect 6435 22588 6491 22644
rect 6517 22588 6573 22644
rect 6599 22588 6655 22644
rect 6681 22599 6702 22644
rect 6702 22599 6737 22644
rect 6763 22599 6768 22644
rect 6768 22599 6819 22644
rect 6681 22588 6737 22599
rect 6763 22588 6819 22599
rect 6845 22588 6901 22644
rect 6927 22588 6983 22644
rect 7009 22588 7065 22644
rect 7091 22588 7147 22644
rect 7173 22588 7229 22644
rect 7255 22599 7256 22644
rect 7256 22599 7308 22644
rect 7308 22599 7311 22644
rect 7337 22599 7374 22644
rect 7374 22599 7393 22644
rect 7255 22588 7311 22599
rect 7337 22588 7393 22599
rect 7419 22588 7475 22644
rect 7501 22588 7557 22644
rect 7583 22588 7639 22644
rect 7665 22588 7721 22644
rect 7747 22588 7803 22644
rect 7829 22599 7862 22644
rect 7862 22599 7876 22644
rect 7876 22599 7885 22644
rect 7911 22599 7928 22644
rect 7928 22599 7967 22644
rect 7829 22588 7885 22599
rect 7911 22588 7967 22599
rect 7993 22603 8047 22644
rect 8047 22603 8049 22644
rect 8075 22603 8099 22644
rect 8099 22603 8131 22644
rect 7993 22588 8049 22603
rect 8075 22588 8131 22603
rect 8157 22603 8169 22644
rect 8169 22603 8213 22644
rect 8157 22588 8213 22603
rect 5613 22530 5646 22564
rect 5646 22530 5660 22564
rect 5660 22530 5669 22564
rect 5696 22530 5712 22564
rect 5712 22530 5752 22564
rect 5613 22513 5669 22530
rect 5696 22513 5752 22530
rect 5613 22508 5646 22513
rect 5646 22508 5660 22513
rect 5660 22508 5669 22513
rect 5696 22508 5712 22513
rect 5712 22508 5752 22513
rect 5779 22508 5835 22564
rect 5861 22508 5917 22564
rect 5943 22508 5999 22564
rect 6025 22508 6081 22564
rect 6107 22530 6148 22564
rect 6148 22530 6163 22564
rect 6189 22530 6200 22564
rect 6200 22530 6214 22564
rect 6214 22530 6245 22564
rect 6107 22513 6163 22530
rect 6189 22513 6245 22530
rect 6107 22508 6148 22513
rect 6148 22508 6163 22513
rect 6189 22508 6200 22513
rect 6200 22508 6214 22513
rect 6214 22508 6245 22513
rect 6271 22508 6327 22564
rect 6353 22508 6409 22564
rect 6435 22508 6491 22564
rect 6517 22508 6573 22564
rect 6599 22508 6655 22564
rect 6681 22530 6702 22564
rect 6702 22530 6737 22564
rect 6763 22530 6768 22564
rect 6768 22530 6819 22564
rect 6681 22513 6737 22530
rect 6763 22513 6819 22530
rect 6681 22508 6702 22513
rect 6702 22508 6737 22513
rect 6763 22508 6768 22513
rect 6768 22508 6819 22513
rect 6845 22508 6901 22564
rect 6927 22508 6983 22564
rect 7009 22508 7065 22564
rect 7091 22508 7147 22564
rect 7173 22508 7229 22564
rect 7255 22530 7256 22564
rect 7256 22530 7308 22564
rect 7308 22530 7311 22564
rect 7337 22530 7374 22564
rect 7374 22530 7393 22564
rect 7255 22513 7311 22530
rect 7337 22513 7393 22530
rect 7255 22508 7256 22513
rect 7256 22508 7308 22513
rect 7308 22508 7311 22513
rect 7337 22508 7374 22513
rect 7374 22508 7393 22513
rect 7419 22508 7475 22564
rect 7501 22508 7557 22564
rect 7583 22508 7639 22564
rect 7665 22508 7721 22564
rect 7747 22508 7803 22564
rect 7829 22530 7862 22564
rect 7862 22530 7876 22564
rect 7876 22530 7885 22564
rect 7911 22530 7928 22564
rect 7928 22530 7967 22564
rect 7829 22513 7885 22530
rect 7911 22513 7967 22530
rect 7829 22508 7862 22513
rect 7862 22508 7876 22513
rect 7876 22508 7885 22513
rect 7911 22508 7928 22513
rect 7928 22508 7967 22513
rect 7993 22534 8047 22564
rect 8047 22534 8049 22564
rect 8075 22534 8099 22564
rect 8099 22534 8131 22564
rect 7993 22517 8049 22534
rect 8075 22517 8131 22534
rect 7993 22508 8047 22517
rect 8047 22508 8049 22517
rect 8075 22508 8099 22517
rect 8099 22508 8131 22517
rect 8157 22534 8169 22564
rect 8169 22534 8213 22564
rect 8157 22517 8213 22534
rect 8157 22508 8169 22517
rect 8169 22508 8213 22517
rect 5613 22461 5646 22484
rect 5646 22461 5660 22484
rect 5660 22461 5669 22484
rect 5696 22461 5712 22484
rect 5712 22461 5752 22484
rect 5613 22444 5669 22461
rect 5696 22444 5752 22461
rect 5613 22428 5646 22444
rect 5646 22428 5660 22444
rect 5660 22428 5669 22444
rect 5696 22428 5712 22444
rect 5712 22428 5752 22444
rect 5779 22428 5835 22484
rect 5861 22428 5917 22484
rect 5943 22428 5999 22484
rect 6025 22428 6081 22484
rect 6107 22461 6148 22484
rect 6148 22461 6163 22484
rect 6189 22461 6200 22484
rect 6200 22461 6214 22484
rect 6214 22461 6245 22484
rect 6107 22444 6163 22461
rect 6189 22444 6245 22461
rect 6107 22428 6148 22444
rect 6148 22428 6163 22444
rect 6189 22428 6200 22444
rect 6200 22428 6214 22444
rect 6214 22428 6245 22444
rect 6271 22428 6327 22484
rect 6353 22428 6409 22484
rect 6435 22428 6491 22484
rect 6517 22428 6573 22484
rect 6599 22428 6655 22484
rect 6681 22461 6702 22484
rect 6702 22461 6737 22484
rect 6763 22461 6768 22484
rect 6768 22461 6819 22484
rect 6681 22444 6737 22461
rect 6763 22444 6819 22461
rect 6681 22428 6702 22444
rect 6702 22428 6737 22444
rect 6763 22428 6768 22444
rect 6768 22428 6819 22444
rect 6845 22428 6901 22484
rect 6927 22428 6983 22484
rect 7009 22428 7065 22484
rect 7091 22428 7147 22484
rect 7173 22428 7229 22484
rect 7255 22461 7256 22484
rect 7256 22461 7308 22484
rect 7308 22461 7311 22484
rect 7337 22461 7374 22484
rect 7374 22461 7393 22484
rect 7255 22444 7311 22461
rect 7337 22444 7393 22461
rect 7255 22428 7256 22444
rect 7256 22428 7308 22444
rect 7308 22428 7311 22444
rect 7337 22428 7374 22444
rect 7374 22428 7393 22444
rect 7419 22428 7475 22484
rect 7501 22428 7557 22484
rect 7583 22428 7639 22484
rect 7665 22428 7721 22484
rect 7747 22428 7803 22484
rect 7829 22461 7862 22484
rect 7862 22461 7876 22484
rect 7876 22461 7885 22484
rect 7911 22461 7928 22484
rect 7928 22461 7967 22484
rect 7829 22444 7885 22461
rect 7911 22444 7967 22461
rect 7829 22428 7862 22444
rect 7862 22428 7876 22444
rect 7876 22428 7885 22444
rect 7911 22428 7928 22444
rect 7928 22428 7967 22444
rect 7993 22465 8047 22484
rect 8047 22465 8049 22484
rect 8075 22465 8099 22484
rect 8099 22465 8131 22484
rect 7993 22448 8049 22465
rect 8075 22448 8131 22465
rect 7993 22428 8047 22448
rect 8047 22428 8049 22448
rect 8075 22428 8099 22448
rect 8099 22428 8131 22448
rect 8157 22465 8169 22484
rect 8169 22465 8213 22484
rect 8157 22448 8213 22465
rect 8157 22428 8169 22448
rect 8169 22428 8213 22448
rect 5613 22392 5646 22404
rect 5646 22392 5660 22404
rect 5660 22392 5669 22404
rect 5696 22392 5712 22404
rect 5712 22392 5752 22404
rect 5613 22375 5669 22392
rect 5696 22375 5752 22392
rect 5613 22348 5646 22375
rect 5646 22348 5660 22375
rect 5660 22348 5669 22375
rect 5696 22348 5712 22375
rect 5712 22348 5752 22375
rect 5779 22348 5835 22404
rect 5861 22348 5917 22404
rect 5943 22348 5999 22404
rect 6025 22348 6081 22404
rect 6107 22392 6148 22404
rect 6148 22392 6163 22404
rect 6189 22392 6200 22404
rect 6200 22392 6214 22404
rect 6214 22392 6245 22404
rect 6107 22375 6163 22392
rect 6189 22375 6245 22392
rect 6107 22348 6148 22375
rect 6148 22348 6163 22375
rect 6189 22348 6200 22375
rect 6200 22348 6214 22375
rect 6214 22348 6245 22375
rect 6271 22348 6327 22404
rect 6353 22348 6409 22404
rect 6435 22348 6491 22404
rect 6517 22348 6573 22404
rect 6599 22348 6655 22404
rect 6681 22392 6702 22404
rect 6702 22392 6737 22404
rect 6763 22392 6768 22404
rect 6768 22392 6819 22404
rect 6681 22375 6737 22392
rect 6763 22375 6819 22392
rect 6681 22348 6702 22375
rect 6702 22348 6737 22375
rect 6763 22348 6768 22375
rect 6768 22348 6819 22375
rect 6845 22348 6901 22404
rect 6927 22348 6983 22404
rect 7009 22348 7065 22404
rect 7091 22348 7147 22404
rect 7173 22348 7229 22404
rect 7255 22392 7256 22404
rect 7256 22392 7308 22404
rect 7308 22392 7311 22404
rect 7337 22392 7374 22404
rect 7374 22392 7393 22404
rect 7255 22375 7311 22392
rect 7337 22375 7393 22392
rect 7255 22348 7256 22375
rect 7256 22348 7308 22375
rect 7308 22348 7311 22375
rect 7337 22348 7374 22375
rect 7374 22348 7393 22375
rect 7419 22348 7475 22404
rect 7501 22348 7557 22404
rect 7583 22348 7639 22404
rect 7665 22348 7721 22404
rect 7747 22348 7803 22404
rect 7829 22392 7862 22404
rect 7862 22392 7876 22404
rect 7876 22392 7885 22404
rect 7911 22392 7928 22404
rect 7928 22392 7967 22404
rect 7829 22375 7885 22392
rect 7911 22375 7967 22392
rect 7829 22348 7862 22375
rect 7862 22348 7876 22375
rect 7876 22348 7885 22375
rect 7911 22348 7928 22375
rect 7928 22348 7967 22375
rect 7993 22396 8047 22404
rect 8047 22396 8049 22404
rect 8075 22396 8099 22404
rect 8099 22396 8131 22404
rect 7993 22378 8049 22396
rect 8075 22378 8131 22396
rect 7993 22348 8047 22378
rect 8047 22348 8049 22378
rect 8075 22348 8099 22378
rect 8099 22348 8131 22378
rect 8157 22396 8169 22404
rect 8169 22396 8213 22404
rect 8157 22378 8213 22396
rect 8157 22348 8169 22378
rect 8169 22348 8213 22378
rect 5613 22323 5646 22324
rect 5646 22323 5660 22324
rect 5660 22323 5669 22324
rect 5696 22323 5712 22324
rect 5712 22323 5752 22324
rect 5613 22306 5669 22323
rect 5696 22306 5752 22323
rect 5613 22268 5646 22306
rect 5646 22268 5660 22306
rect 5660 22268 5669 22306
rect 5696 22268 5712 22306
rect 5712 22268 5752 22306
rect 5779 22268 5835 22324
rect 5861 22268 5917 22324
rect 5943 22268 5999 22324
rect 6025 22268 6081 22324
rect 6107 22323 6148 22324
rect 6148 22323 6163 22324
rect 6189 22323 6200 22324
rect 6200 22323 6214 22324
rect 6214 22323 6245 22324
rect 6107 22306 6163 22323
rect 6189 22306 6245 22323
rect 6107 22268 6148 22306
rect 6148 22268 6163 22306
rect 6189 22268 6200 22306
rect 6200 22268 6214 22306
rect 6214 22268 6245 22306
rect 6271 22268 6327 22324
rect 6353 22268 6409 22324
rect 6435 22268 6491 22324
rect 6517 22268 6573 22324
rect 6599 22268 6655 22324
rect 6681 22323 6702 22324
rect 6702 22323 6737 22324
rect 6763 22323 6768 22324
rect 6768 22323 6819 22324
rect 6681 22306 6737 22323
rect 6763 22306 6819 22323
rect 6681 22268 6702 22306
rect 6702 22268 6737 22306
rect 6763 22268 6768 22306
rect 6768 22268 6819 22306
rect 6845 22268 6901 22324
rect 6927 22268 6983 22324
rect 7009 22268 7065 22324
rect 7091 22268 7147 22324
rect 7173 22268 7229 22324
rect 7255 22323 7256 22324
rect 7256 22323 7308 22324
rect 7308 22323 7311 22324
rect 7337 22323 7374 22324
rect 7374 22323 7393 22324
rect 7255 22306 7311 22323
rect 7337 22306 7393 22323
rect 7255 22268 7256 22306
rect 7256 22268 7308 22306
rect 7308 22268 7311 22306
rect 7337 22268 7374 22306
rect 7374 22268 7393 22306
rect 7419 22268 7475 22324
rect 7501 22268 7557 22324
rect 7583 22268 7639 22324
rect 7665 22268 7721 22324
rect 7747 22268 7803 22324
rect 7829 22323 7862 22324
rect 7862 22323 7876 22324
rect 7876 22323 7885 22324
rect 7911 22323 7928 22324
rect 7928 22323 7967 22324
rect 7829 22306 7885 22323
rect 7911 22306 7967 22323
rect 7829 22268 7862 22306
rect 7862 22268 7876 22306
rect 7876 22268 7885 22306
rect 7911 22268 7928 22306
rect 7928 22268 7967 22306
rect 7993 22308 8049 22324
rect 8075 22308 8131 22324
rect 7993 22268 8047 22308
rect 8047 22268 8049 22308
rect 8075 22268 8099 22308
rect 8099 22268 8131 22308
rect 8157 22308 8213 22324
rect 8157 22268 8169 22308
rect 8169 22268 8213 22308
rect 5613 22236 5669 22244
rect 5696 22236 5752 22244
rect 5613 22188 5646 22236
rect 5646 22188 5660 22236
rect 5660 22188 5669 22236
rect 5696 22188 5712 22236
rect 5712 22188 5752 22236
rect 5779 22188 5835 22244
rect 5861 22188 5917 22244
rect 5943 22188 5999 22244
rect 6025 22188 6081 22244
rect 6107 22236 6163 22244
rect 6189 22236 6245 22244
rect 6107 22188 6148 22236
rect 6148 22188 6163 22236
rect 6189 22188 6200 22236
rect 6200 22188 6214 22236
rect 6214 22188 6245 22236
rect 6271 22188 6327 22244
rect 6353 22188 6409 22244
rect 6435 22188 6491 22244
rect 6517 22188 6573 22244
rect 6599 22188 6655 22244
rect 6681 22236 6737 22244
rect 6763 22236 6819 22244
rect 6681 22188 6702 22236
rect 6702 22188 6737 22236
rect 6763 22188 6768 22236
rect 6768 22188 6819 22236
rect 6845 22188 6901 22244
rect 6927 22188 6983 22244
rect 7009 22188 7065 22244
rect 7091 22188 7147 22244
rect 7173 22188 7229 22244
rect 7255 22236 7311 22244
rect 7337 22236 7393 22244
rect 7255 22188 7256 22236
rect 7256 22188 7308 22236
rect 7308 22188 7311 22236
rect 7337 22188 7374 22236
rect 7374 22188 7393 22236
rect 7419 22188 7475 22244
rect 7501 22188 7557 22244
rect 7583 22188 7639 22244
rect 7665 22188 7721 22244
rect 7747 22188 7803 22244
rect 7829 22236 7885 22244
rect 7911 22236 7967 22244
rect 7829 22188 7862 22236
rect 7862 22188 7876 22236
rect 7876 22188 7885 22236
rect 7911 22188 7928 22236
rect 7928 22188 7967 22236
rect 7993 22238 8049 22244
rect 8075 22238 8131 22244
rect 7993 22188 8047 22238
rect 8047 22188 8049 22238
rect 8075 22188 8099 22238
rect 8099 22188 8131 22238
rect 8157 22238 8213 22244
rect 8157 22188 8169 22238
rect 8169 22188 8213 22238
rect 5613 22114 5646 22164
rect 5646 22114 5660 22164
rect 5660 22114 5669 22164
rect 5696 22114 5712 22164
rect 5712 22114 5752 22164
rect 5613 22108 5669 22114
rect 5696 22108 5752 22114
rect 5779 22108 5835 22164
rect 5861 22108 5917 22164
rect 5943 22108 5999 22164
rect 6025 22108 6081 22164
rect 6107 22114 6148 22164
rect 6148 22114 6163 22164
rect 6189 22114 6200 22164
rect 6200 22114 6214 22164
rect 6214 22114 6245 22164
rect 6107 22108 6163 22114
rect 6189 22108 6245 22114
rect 6271 22108 6327 22164
rect 6353 22108 6409 22164
rect 6435 22108 6491 22164
rect 6517 22108 6573 22164
rect 6599 22108 6655 22164
rect 6681 22114 6702 22164
rect 6702 22114 6737 22164
rect 6763 22114 6768 22164
rect 6768 22114 6819 22164
rect 6681 22108 6737 22114
rect 6763 22108 6819 22114
rect 6845 22108 6901 22164
rect 6927 22108 6983 22164
rect 7009 22108 7065 22164
rect 7091 22108 7147 22164
rect 7173 22108 7229 22164
rect 7255 22114 7256 22164
rect 7256 22114 7308 22164
rect 7308 22114 7311 22164
rect 7337 22114 7374 22164
rect 7374 22114 7393 22164
rect 7255 22108 7311 22114
rect 7337 22108 7393 22114
rect 7419 22108 7475 22164
rect 7501 22108 7557 22164
rect 7583 22108 7639 22164
rect 7665 22108 7721 22164
rect 7747 22108 7803 22164
rect 7829 22114 7862 22164
rect 7862 22114 7876 22164
rect 7876 22114 7885 22164
rect 7911 22114 7928 22164
rect 7928 22114 7967 22164
rect 7829 22108 7885 22114
rect 7911 22108 7967 22114
rect 7993 22116 8047 22164
rect 8047 22116 8049 22164
rect 8075 22116 8099 22164
rect 8099 22116 8131 22164
rect 7993 22108 8049 22116
rect 8075 22108 8131 22116
rect 8157 22116 8169 22164
rect 8169 22116 8213 22164
rect 8157 22108 8213 22116
rect 2733 21931 2789 21987
rect 2814 21931 2870 21987
rect 2895 21931 2951 21987
rect 2976 21931 3032 21987
rect 3057 21931 3113 21987
rect 3138 21931 3194 21987
rect 3219 21931 3275 21987
rect 3300 21931 3356 21987
rect 3381 21931 3437 21987
rect 3462 21931 3518 21987
rect 3543 21931 3599 21987
rect 3624 21931 3680 21987
rect 3705 21931 3761 21987
rect 3786 21931 3842 21987
rect 3867 21931 3923 21987
rect 3948 21931 4004 21987
rect 4029 21931 4085 21987
rect 4110 21931 4166 21987
rect 4191 21931 4247 21987
rect 4272 21931 4328 21987
rect 4353 21931 4409 21987
rect 4434 21931 4490 21987
rect 4515 21931 4571 21987
rect 4596 21931 4652 21987
rect 4677 21931 4733 21987
rect 4758 21931 4814 21987
rect 4839 21931 4895 21987
rect 4920 21931 4976 21987
rect 5001 21931 5057 21987
rect 5082 21931 5138 21987
rect 2733 21851 2789 21907
rect 2814 21851 2870 21907
rect 2895 21851 2951 21907
rect 2976 21851 3032 21907
rect 3057 21851 3113 21907
rect 3138 21851 3194 21907
rect 3219 21851 3275 21907
rect 3300 21851 3356 21907
rect 3381 21851 3437 21907
rect 3462 21851 3518 21907
rect 3543 21851 3599 21907
rect 3624 21851 3680 21907
rect 3705 21851 3761 21907
rect 3786 21851 3842 21907
rect 3867 21851 3923 21907
rect 3948 21851 4004 21907
rect 4029 21851 4085 21907
rect 4110 21851 4166 21907
rect 4191 21851 4247 21907
rect 4272 21851 4328 21907
rect 4353 21851 4409 21907
rect 4434 21851 4490 21907
rect 4515 21851 4571 21907
rect 4596 21851 4652 21907
rect 4677 21851 4733 21907
rect 4758 21851 4814 21907
rect 4839 21851 4895 21907
rect 4920 21851 4976 21907
rect 5001 21851 5057 21907
rect 5082 21851 5138 21907
rect 2733 21771 2789 21827
rect 2814 21771 2870 21827
rect 2895 21771 2951 21827
rect 2976 21771 3032 21827
rect 3057 21771 3113 21827
rect 3138 21771 3194 21827
rect 3219 21771 3275 21827
rect 3300 21771 3356 21827
rect 3381 21771 3437 21827
rect 3462 21771 3518 21827
rect 3543 21771 3599 21827
rect 3624 21771 3680 21827
rect 3705 21771 3761 21827
rect 3786 21771 3842 21827
rect 3867 21771 3923 21827
rect 3948 21771 4004 21827
rect 4029 21771 4085 21827
rect 4110 21771 4166 21827
rect 4191 21771 4247 21827
rect 4272 21771 4328 21827
rect 4353 21771 4409 21827
rect 4434 21771 4490 21827
rect 4515 21771 4571 21827
rect 4596 21771 4652 21827
rect 4677 21771 4733 21827
rect 4758 21771 4814 21827
rect 4839 21771 4895 21827
rect 4920 21771 4976 21827
rect 5001 21771 5057 21827
rect 5082 21771 5138 21827
rect 2733 21691 2789 21747
rect 2814 21691 2870 21747
rect 2895 21691 2951 21747
rect 2976 21691 3032 21747
rect 3057 21691 3113 21747
rect 3138 21691 3194 21747
rect 3219 21691 3275 21747
rect 3300 21691 3356 21747
rect 3381 21691 3437 21747
rect 3462 21691 3518 21747
rect 3543 21691 3599 21747
rect 3624 21691 3680 21747
rect 3705 21691 3761 21747
rect 3786 21691 3842 21747
rect 3867 21691 3923 21747
rect 3948 21691 4004 21747
rect 4029 21691 4085 21747
rect 4110 21691 4166 21747
rect 4191 21691 4247 21747
rect 4272 21691 4328 21747
rect 4353 21691 4409 21747
rect 4434 21691 4490 21747
rect 4515 21691 4571 21747
rect 4596 21691 4652 21747
rect 4677 21691 4733 21747
rect 4758 21691 4814 21747
rect 4839 21691 4895 21747
rect 4920 21691 4976 21747
rect 5001 21691 5057 21747
rect 5082 21691 5138 21747
rect 2733 21611 2789 21667
rect 2814 21611 2870 21667
rect 2895 21611 2951 21667
rect 2976 21611 3032 21667
rect 3057 21611 3113 21667
rect 3138 21611 3194 21667
rect 3219 21611 3275 21667
rect 3300 21611 3356 21667
rect 3381 21611 3437 21667
rect 3462 21611 3518 21667
rect 3543 21611 3599 21667
rect 3624 21611 3680 21667
rect 3705 21611 3761 21667
rect 3786 21611 3842 21667
rect 3867 21611 3923 21667
rect 3948 21611 4004 21667
rect 4029 21611 4085 21667
rect 4110 21611 4166 21667
rect 4191 21611 4247 21667
rect 4272 21611 4328 21667
rect 4353 21611 4409 21667
rect 4434 21611 4490 21667
rect 4515 21611 4571 21667
rect 4596 21611 4652 21667
rect 4677 21611 4733 21667
rect 4758 21611 4814 21667
rect 4839 21611 4895 21667
rect 4920 21611 4976 21667
rect 5001 21611 5057 21667
rect 5082 21611 5138 21667
rect 2733 21531 2789 21587
rect 2814 21531 2870 21587
rect 2895 21531 2951 21587
rect 2976 21531 3032 21587
rect 3057 21531 3113 21587
rect 3138 21531 3194 21587
rect 3219 21531 3275 21587
rect 3300 21531 3356 21587
rect 3381 21531 3437 21587
rect 3462 21531 3518 21587
rect 3543 21531 3599 21587
rect 3624 21531 3680 21587
rect 3705 21531 3761 21587
rect 3786 21531 3842 21587
rect 3867 21531 3923 21587
rect 3948 21531 4004 21587
rect 4029 21531 4085 21587
rect 4110 21531 4166 21587
rect 4191 21531 4247 21587
rect 4272 21531 4328 21587
rect 4353 21531 4409 21587
rect 4434 21531 4490 21587
rect 4515 21531 4571 21587
rect 4596 21531 4652 21587
rect 4677 21531 4733 21587
rect 4758 21531 4814 21587
rect 4839 21531 4895 21587
rect 4920 21531 4976 21587
rect 5001 21531 5057 21587
rect 5082 21531 5138 21587
rect 2733 21451 2789 21507
rect 2814 21451 2870 21507
rect 2895 21451 2951 21507
rect 2976 21451 3032 21507
rect 3057 21451 3113 21507
rect 3138 21451 3194 21507
rect 3219 21451 3275 21507
rect 3300 21451 3356 21507
rect 3381 21451 3437 21507
rect 3462 21451 3518 21507
rect 3543 21451 3599 21507
rect 3624 21451 3680 21507
rect 3705 21451 3761 21507
rect 3786 21451 3842 21507
rect 3867 21451 3923 21507
rect 3948 21451 4004 21507
rect 4029 21451 4085 21507
rect 4110 21451 4166 21507
rect 4191 21451 4247 21507
rect 4272 21451 4328 21507
rect 4353 21451 4409 21507
rect 4434 21451 4490 21507
rect 4515 21451 4571 21507
rect 4596 21451 4652 21507
rect 4677 21451 4733 21507
rect 4758 21451 4814 21507
rect 4839 21451 4895 21507
rect 4920 21451 4976 21507
rect 5001 21451 5057 21507
rect 5082 21451 5138 21507
rect 2733 21371 2789 21427
rect 2814 21371 2870 21427
rect 2895 21371 2951 21427
rect 2976 21371 3032 21427
rect 3057 21371 3113 21427
rect 3138 21371 3194 21427
rect 3219 21371 3275 21427
rect 3300 21371 3356 21427
rect 3381 21371 3437 21427
rect 3462 21371 3518 21427
rect 3543 21371 3599 21427
rect 3624 21371 3680 21427
rect 3705 21371 3761 21427
rect 3786 21371 3842 21427
rect 3867 21371 3923 21427
rect 3948 21371 4004 21427
rect 4029 21371 4085 21427
rect 4110 21371 4166 21427
rect 4191 21371 4247 21427
rect 4272 21371 4328 21427
rect 4353 21371 4409 21427
rect 4434 21371 4490 21427
rect 4515 21371 4571 21427
rect 4596 21371 4652 21427
rect 4677 21371 4733 21427
rect 4758 21371 4814 21427
rect 4839 21371 4895 21427
rect 4920 21371 4976 21427
rect 5001 21371 5057 21427
rect 5082 21371 5138 21427
rect 5163 21371 5299 21987
rect 5613 20720 5669 20724
rect 5696 20720 5752 20724
rect 5613 20668 5646 20720
rect 5646 20668 5660 20720
rect 5660 20668 5669 20720
rect 5696 20668 5712 20720
rect 5712 20668 5752 20720
rect 5779 20668 5835 20724
rect 5861 20668 5917 20724
rect 5943 20668 5999 20724
rect 6025 20668 6081 20724
rect 6107 20720 6163 20724
rect 6189 20720 6245 20724
rect 6107 20668 6148 20720
rect 6148 20668 6163 20720
rect 6189 20668 6200 20720
rect 6200 20668 6214 20720
rect 6214 20668 6245 20720
rect 6271 20668 6327 20724
rect 6353 20668 6409 20724
rect 6435 20668 6491 20724
rect 6517 20668 6573 20724
rect 6599 20668 6655 20724
rect 6681 20720 6737 20724
rect 6763 20720 6819 20724
rect 6681 20668 6702 20720
rect 6702 20668 6737 20720
rect 6763 20668 6768 20720
rect 6768 20668 6819 20720
rect 6845 20668 6901 20724
rect 6927 20668 6983 20724
rect 7009 20668 7065 20724
rect 7091 20668 7147 20724
rect 7173 20668 7229 20724
rect 7255 20720 7311 20724
rect 7337 20720 7393 20724
rect 7255 20668 7256 20720
rect 7256 20668 7308 20720
rect 7308 20668 7311 20720
rect 7337 20668 7374 20720
rect 7374 20668 7393 20720
rect 7419 20668 7475 20724
rect 7501 20668 7557 20724
rect 7583 20668 7639 20724
rect 7665 20668 7721 20724
rect 7747 20668 7803 20724
rect 7829 20720 7885 20724
rect 7911 20720 7967 20724
rect 7829 20668 7862 20720
rect 7862 20668 7876 20720
rect 7876 20668 7885 20720
rect 7911 20668 7928 20720
rect 7928 20668 7967 20720
rect 7993 20672 8047 20724
rect 8047 20672 8049 20724
rect 8075 20672 8099 20724
rect 8099 20672 8131 20724
rect 7993 20668 8049 20672
rect 8075 20668 8131 20672
rect 8157 20672 8169 20724
rect 8169 20672 8213 20724
rect 8157 20668 8213 20672
rect 5613 20599 5646 20644
rect 5646 20599 5660 20644
rect 5660 20599 5669 20644
rect 5696 20599 5712 20644
rect 5712 20599 5752 20644
rect 5613 20588 5669 20599
rect 5696 20588 5752 20599
rect 5779 20588 5835 20644
rect 5861 20588 5917 20644
rect 5943 20588 5999 20644
rect 6025 20588 6081 20644
rect 6107 20599 6148 20644
rect 6148 20599 6163 20644
rect 6189 20599 6200 20644
rect 6200 20599 6214 20644
rect 6214 20599 6245 20644
rect 6107 20588 6163 20599
rect 6189 20588 6245 20599
rect 6271 20588 6327 20644
rect 6353 20588 6409 20644
rect 6435 20588 6491 20644
rect 6517 20588 6573 20644
rect 6599 20588 6655 20644
rect 6681 20599 6702 20644
rect 6702 20599 6737 20644
rect 6763 20599 6768 20644
rect 6768 20599 6819 20644
rect 6681 20588 6737 20599
rect 6763 20588 6819 20599
rect 6845 20588 6901 20644
rect 6927 20588 6983 20644
rect 7009 20588 7065 20644
rect 7091 20588 7147 20644
rect 7173 20588 7229 20644
rect 7255 20599 7256 20644
rect 7256 20599 7308 20644
rect 7308 20599 7311 20644
rect 7337 20599 7374 20644
rect 7374 20599 7393 20644
rect 7255 20588 7311 20599
rect 7337 20588 7393 20599
rect 7419 20588 7475 20644
rect 7501 20588 7557 20644
rect 7583 20588 7639 20644
rect 7665 20588 7721 20644
rect 7747 20588 7803 20644
rect 7829 20599 7862 20644
rect 7862 20599 7876 20644
rect 7876 20599 7885 20644
rect 7911 20599 7928 20644
rect 7928 20599 7967 20644
rect 7829 20588 7885 20599
rect 7911 20588 7967 20599
rect 7993 20603 8047 20644
rect 8047 20603 8049 20644
rect 8075 20603 8099 20644
rect 8099 20603 8131 20644
rect 7993 20588 8049 20603
rect 8075 20588 8131 20603
rect 8157 20603 8169 20644
rect 8169 20603 8213 20644
rect 8157 20588 8213 20603
rect 5613 20530 5646 20564
rect 5646 20530 5660 20564
rect 5660 20530 5669 20564
rect 5696 20530 5712 20564
rect 5712 20530 5752 20564
rect 5613 20513 5669 20530
rect 5696 20513 5752 20530
rect 5613 20508 5646 20513
rect 5646 20508 5660 20513
rect 5660 20508 5669 20513
rect 5696 20508 5712 20513
rect 5712 20508 5752 20513
rect 5779 20508 5835 20564
rect 5861 20508 5917 20564
rect 5943 20508 5999 20564
rect 6025 20508 6081 20564
rect 6107 20530 6148 20564
rect 6148 20530 6163 20564
rect 6189 20530 6200 20564
rect 6200 20530 6214 20564
rect 6214 20530 6245 20564
rect 6107 20513 6163 20530
rect 6189 20513 6245 20530
rect 6107 20508 6148 20513
rect 6148 20508 6163 20513
rect 6189 20508 6200 20513
rect 6200 20508 6214 20513
rect 6214 20508 6245 20513
rect 6271 20508 6327 20564
rect 6353 20508 6409 20564
rect 6435 20508 6491 20564
rect 6517 20508 6573 20564
rect 6599 20508 6655 20564
rect 6681 20530 6702 20564
rect 6702 20530 6737 20564
rect 6763 20530 6768 20564
rect 6768 20530 6819 20564
rect 6681 20513 6737 20530
rect 6763 20513 6819 20530
rect 6681 20508 6702 20513
rect 6702 20508 6737 20513
rect 6763 20508 6768 20513
rect 6768 20508 6819 20513
rect 6845 20508 6901 20564
rect 6927 20508 6983 20564
rect 7009 20508 7065 20564
rect 7091 20508 7147 20564
rect 7173 20508 7229 20564
rect 7255 20530 7256 20564
rect 7256 20530 7308 20564
rect 7308 20530 7311 20564
rect 7337 20530 7374 20564
rect 7374 20530 7393 20564
rect 7255 20513 7311 20530
rect 7337 20513 7393 20530
rect 7255 20508 7256 20513
rect 7256 20508 7308 20513
rect 7308 20508 7311 20513
rect 7337 20508 7374 20513
rect 7374 20508 7393 20513
rect 7419 20508 7475 20564
rect 7501 20508 7557 20564
rect 7583 20508 7639 20564
rect 7665 20508 7721 20564
rect 7747 20508 7803 20564
rect 7829 20530 7862 20564
rect 7862 20530 7876 20564
rect 7876 20530 7885 20564
rect 7911 20530 7928 20564
rect 7928 20530 7967 20564
rect 7829 20513 7885 20530
rect 7911 20513 7967 20530
rect 7829 20508 7862 20513
rect 7862 20508 7876 20513
rect 7876 20508 7885 20513
rect 7911 20508 7928 20513
rect 7928 20508 7967 20513
rect 7993 20534 8047 20564
rect 8047 20534 8049 20564
rect 8075 20534 8099 20564
rect 8099 20534 8131 20564
rect 7993 20517 8049 20534
rect 8075 20517 8131 20534
rect 7993 20508 8047 20517
rect 8047 20508 8049 20517
rect 8075 20508 8099 20517
rect 8099 20508 8131 20517
rect 8157 20534 8169 20564
rect 8169 20534 8213 20564
rect 8157 20517 8213 20534
rect 8157 20508 8169 20517
rect 8169 20508 8213 20517
rect 5613 20461 5646 20484
rect 5646 20461 5660 20484
rect 5660 20461 5669 20484
rect 5696 20461 5712 20484
rect 5712 20461 5752 20484
rect 5613 20444 5669 20461
rect 5696 20444 5752 20461
rect 5613 20428 5646 20444
rect 5646 20428 5660 20444
rect 5660 20428 5669 20444
rect 5696 20428 5712 20444
rect 5712 20428 5752 20444
rect 5779 20428 5835 20484
rect 5861 20428 5917 20484
rect 5943 20428 5999 20484
rect 6025 20428 6081 20484
rect 6107 20461 6148 20484
rect 6148 20461 6163 20484
rect 6189 20461 6200 20484
rect 6200 20461 6214 20484
rect 6214 20461 6245 20484
rect 6107 20444 6163 20461
rect 6189 20444 6245 20461
rect 6107 20428 6148 20444
rect 6148 20428 6163 20444
rect 6189 20428 6200 20444
rect 6200 20428 6214 20444
rect 6214 20428 6245 20444
rect 6271 20428 6327 20484
rect 6353 20428 6409 20484
rect 6435 20428 6491 20484
rect 6517 20428 6573 20484
rect 6599 20428 6655 20484
rect 6681 20461 6702 20484
rect 6702 20461 6737 20484
rect 6763 20461 6768 20484
rect 6768 20461 6819 20484
rect 6681 20444 6737 20461
rect 6763 20444 6819 20461
rect 6681 20428 6702 20444
rect 6702 20428 6737 20444
rect 6763 20428 6768 20444
rect 6768 20428 6819 20444
rect 6845 20428 6901 20484
rect 6927 20428 6983 20484
rect 7009 20428 7065 20484
rect 7091 20428 7147 20484
rect 7173 20428 7229 20484
rect 7255 20461 7256 20484
rect 7256 20461 7308 20484
rect 7308 20461 7311 20484
rect 7337 20461 7374 20484
rect 7374 20461 7393 20484
rect 7255 20444 7311 20461
rect 7337 20444 7393 20461
rect 7255 20428 7256 20444
rect 7256 20428 7308 20444
rect 7308 20428 7311 20444
rect 7337 20428 7374 20444
rect 7374 20428 7393 20444
rect 7419 20428 7475 20484
rect 7501 20428 7557 20484
rect 7583 20428 7639 20484
rect 7665 20428 7721 20484
rect 7747 20428 7803 20484
rect 7829 20461 7862 20484
rect 7862 20461 7876 20484
rect 7876 20461 7885 20484
rect 7911 20461 7928 20484
rect 7928 20461 7967 20484
rect 7829 20444 7885 20461
rect 7911 20444 7967 20461
rect 7829 20428 7862 20444
rect 7862 20428 7876 20444
rect 7876 20428 7885 20444
rect 7911 20428 7928 20444
rect 7928 20428 7967 20444
rect 7993 20465 8047 20484
rect 8047 20465 8049 20484
rect 8075 20465 8099 20484
rect 8099 20465 8131 20484
rect 7993 20448 8049 20465
rect 8075 20448 8131 20465
rect 7993 20428 8047 20448
rect 8047 20428 8049 20448
rect 8075 20428 8099 20448
rect 8099 20428 8131 20448
rect 8157 20465 8169 20484
rect 8169 20465 8213 20484
rect 8157 20448 8213 20465
rect 8157 20428 8169 20448
rect 8169 20428 8213 20448
rect 5613 20392 5646 20404
rect 5646 20392 5660 20404
rect 5660 20392 5669 20404
rect 5696 20392 5712 20404
rect 5712 20392 5752 20404
rect 5613 20375 5669 20392
rect 5696 20375 5752 20392
rect 5613 20348 5646 20375
rect 5646 20348 5660 20375
rect 5660 20348 5669 20375
rect 5696 20348 5712 20375
rect 5712 20348 5752 20375
rect 5779 20348 5835 20404
rect 5861 20348 5917 20404
rect 5943 20348 5999 20404
rect 6025 20348 6081 20404
rect 6107 20392 6148 20404
rect 6148 20392 6163 20404
rect 6189 20392 6200 20404
rect 6200 20392 6214 20404
rect 6214 20392 6245 20404
rect 6107 20375 6163 20392
rect 6189 20375 6245 20392
rect 6107 20348 6148 20375
rect 6148 20348 6163 20375
rect 6189 20348 6200 20375
rect 6200 20348 6214 20375
rect 6214 20348 6245 20375
rect 6271 20348 6327 20404
rect 6353 20348 6409 20404
rect 6435 20348 6491 20404
rect 6517 20348 6573 20404
rect 6599 20348 6655 20404
rect 6681 20392 6702 20404
rect 6702 20392 6737 20404
rect 6763 20392 6768 20404
rect 6768 20392 6819 20404
rect 6681 20375 6737 20392
rect 6763 20375 6819 20392
rect 6681 20348 6702 20375
rect 6702 20348 6737 20375
rect 6763 20348 6768 20375
rect 6768 20348 6819 20375
rect 6845 20348 6901 20404
rect 6927 20348 6983 20404
rect 7009 20348 7065 20404
rect 7091 20348 7147 20404
rect 7173 20348 7229 20404
rect 7255 20392 7256 20404
rect 7256 20392 7308 20404
rect 7308 20392 7311 20404
rect 7337 20392 7374 20404
rect 7374 20392 7393 20404
rect 7255 20375 7311 20392
rect 7337 20375 7393 20392
rect 7255 20348 7256 20375
rect 7256 20348 7308 20375
rect 7308 20348 7311 20375
rect 7337 20348 7374 20375
rect 7374 20348 7393 20375
rect 7419 20348 7475 20404
rect 7501 20348 7557 20404
rect 7583 20348 7639 20404
rect 7665 20348 7721 20404
rect 7747 20348 7803 20404
rect 7829 20392 7862 20404
rect 7862 20392 7876 20404
rect 7876 20392 7885 20404
rect 7911 20392 7928 20404
rect 7928 20392 7967 20404
rect 7829 20375 7885 20392
rect 7911 20375 7967 20392
rect 7829 20348 7862 20375
rect 7862 20348 7876 20375
rect 7876 20348 7885 20375
rect 7911 20348 7928 20375
rect 7928 20348 7967 20375
rect 7993 20396 8047 20404
rect 8047 20396 8049 20404
rect 8075 20396 8099 20404
rect 8099 20396 8131 20404
rect 7993 20378 8049 20396
rect 8075 20378 8131 20396
rect 7993 20348 8047 20378
rect 8047 20348 8049 20378
rect 8075 20348 8099 20378
rect 8099 20348 8131 20378
rect 8157 20396 8169 20404
rect 8169 20396 8213 20404
rect 8157 20378 8213 20396
rect 8157 20348 8169 20378
rect 8169 20348 8213 20378
rect 5613 20323 5646 20324
rect 5646 20323 5660 20324
rect 5660 20323 5669 20324
rect 5696 20323 5712 20324
rect 5712 20323 5752 20324
rect 5613 20306 5669 20323
rect 5696 20306 5752 20323
rect 5613 20268 5646 20306
rect 5646 20268 5660 20306
rect 5660 20268 5669 20306
rect 5696 20268 5712 20306
rect 5712 20268 5752 20306
rect 5779 20268 5835 20324
rect 5861 20268 5917 20324
rect 5943 20268 5999 20324
rect 6025 20268 6081 20324
rect 6107 20323 6148 20324
rect 6148 20323 6163 20324
rect 6189 20323 6200 20324
rect 6200 20323 6214 20324
rect 6214 20323 6245 20324
rect 6107 20306 6163 20323
rect 6189 20306 6245 20323
rect 6107 20268 6148 20306
rect 6148 20268 6163 20306
rect 6189 20268 6200 20306
rect 6200 20268 6214 20306
rect 6214 20268 6245 20306
rect 6271 20268 6327 20324
rect 6353 20268 6409 20324
rect 6435 20268 6491 20324
rect 6517 20268 6573 20324
rect 6599 20268 6655 20324
rect 6681 20323 6702 20324
rect 6702 20323 6737 20324
rect 6763 20323 6768 20324
rect 6768 20323 6819 20324
rect 6681 20306 6737 20323
rect 6763 20306 6819 20323
rect 6681 20268 6702 20306
rect 6702 20268 6737 20306
rect 6763 20268 6768 20306
rect 6768 20268 6819 20306
rect 6845 20268 6901 20324
rect 6927 20268 6983 20324
rect 7009 20268 7065 20324
rect 7091 20268 7147 20324
rect 7173 20268 7229 20324
rect 7255 20323 7256 20324
rect 7256 20323 7308 20324
rect 7308 20323 7311 20324
rect 7337 20323 7374 20324
rect 7374 20323 7393 20324
rect 7255 20306 7311 20323
rect 7337 20306 7393 20323
rect 7255 20268 7256 20306
rect 7256 20268 7308 20306
rect 7308 20268 7311 20306
rect 7337 20268 7374 20306
rect 7374 20268 7393 20306
rect 7419 20268 7475 20324
rect 7501 20268 7557 20324
rect 7583 20268 7639 20324
rect 7665 20268 7721 20324
rect 7747 20268 7803 20324
rect 7829 20323 7862 20324
rect 7862 20323 7876 20324
rect 7876 20323 7885 20324
rect 7911 20323 7928 20324
rect 7928 20323 7967 20324
rect 7829 20306 7885 20323
rect 7911 20306 7967 20323
rect 7829 20268 7862 20306
rect 7862 20268 7876 20306
rect 7876 20268 7885 20306
rect 7911 20268 7928 20306
rect 7928 20268 7967 20306
rect 7993 20308 8049 20324
rect 8075 20308 8131 20324
rect 7993 20268 8047 20308
rect 8047 20268 8049 20308
rect 8075 20268 8099 20308
rect 8099 20268 8131 20308
rect 8157 20308 8213 20324
rect 8157 20268 8169 20308
rect 8169 20268 8213 20308
rect 5613 20236 5669 20244
rect 5696 20236 5752 20244
rect 5613 20188 5646 20236
rect 5646 20188 5660 20236
rect 5660 20188 5669 20236
rect 5696 20188 5712 20236
rect 5712 20188 5752 20236
rect 5779 20188 5835 20244
rect 5861 20188 5917 20244
rect 5943 20188 5999 20244
rect 6025 20188 6081 20244
rect 6107 20236 6163 20244
rect 6189 20236 6245 20244
rect 6107 20188 6148 20236
rect 6148 20188 6163 20236
rect 6189 20188 6200 20236
rect 6200 20188 6214 20236
rect 6214 20188 6245 20236
rect 6271 20188 6327 20244
rect 6353 20188 6409 20244
rect 6435 20188 6491 20244
rect 6517 20188 6573 20244
rect 6599 20188 6655 20244
rect 6681 20236 6737 20244
rect 6763 20236 6819 20244
rect 6681 20188 6702 20236
rect 6702 20188 6737 20236
rect 6763 20188 6768 20236
rect 6768 20188 6819 20236
rect 6845 20188 6901 20244
rect 6927 20188 6983 20244
rect 7009 20188 7065 20244
rect 7091 20188 7147 20244
rect 7173 20188 7229 20244
rect 7255 20236 7311 20244
rect 7337 20236 7393 20244
rect 7255 20188 7256 20236
rect 7256 20188 7308 20236
rect 7308 20188 7311 20236
rect 7337 20188 7374 20236
rect 7374 20188 7393 20236
rect 7419 20188 7475 20244
rect 7501 20188 7557 20244
rect 7583 20188 7639 20244
rect 7665 20188 7721 20244
rect 7747 20188 7803 20244
rect 7829 20236 7885 20244
rect 7911 20236 7967 20244
rect 7829 20188 7862 20236
rect 7862 20188 7876 20236
rect 7876 20188 7885 20236
rect 7911 20188 7928 20236
rect 7928 20188 7967 20236
rect 7993 20238 8049 20244
rect 8075 20238 8131 20244
rect 7993 20188 8047 20238
rect 8047 20188 8049 20238
rect 8075 20188 8099 20238
rect 8099 20188 8131 20238
rect 8157 20238 8213 20244
rect 8157 20188 8169 20238
rect 8169 20188 8213 20238
rect 5613 20114 5646 20164
rect 5646 20114 5660 20164
rect 5660 20114 5669 20164
rect 5696 20114 5712 20164
rect 5712 20114 5752 20164
rect 5613 20108 5669 20114
rect 5696 20108 5752 20114
rect 5779 20108 5835 20164
rect 5861 20108 5917 20164
rect 5943 20108 5999 20164
rect 6025 20108 6081 20164
rect 6107 20114 6148 20164
rect 6148 20114 6163 20164
rect 6189 20114 6200 20164
rect 6200 20114 6214 20164
rect 6214 20114 6245 20164
rect 6107 20108 6163 20114
rect 6189 20108 6245 20114
rect 6271 20108 6327 20164
rect 6353 20108 6409 20164
rect 6435 20108 6491 20164
rect 6517 20108 6573 20164
rect 6599 20108 6655 20164
rect 6681 20114 6702 20164
rect 6702 20114 6737 20164
rect 6763 20114 6768 20164
rect 6768 20114 6819 20164
rect 6681 20108 6737 20114
rect 6763 20108 6819 20114
rect 6845 20108 6901 20164
rect 6927 20108 6983 20164
rect 7009 20108 7065 20164
rect 7091 20108 7147 20164
rect 7173 20108 7229 20164
rect 7255 20114 7256 20164
rect 7256 20114 7308 20164
rect 7308 20114 7311 20164
rect 7337 20114 7374 20164
rect 7374 20114 7393 20164
rect 7255 20108 7311 20114
rect 7337 20108 7393 20114
rect 7419 20108 7475 20164
rect 7501 20108 7557 20164
rect 7583 20108 7639 20164
rect 7665 20108 7721 20164
rect 7747 20108 7803 20164
rect 7829 20114 7862 20164
rect 7862 20114 7876 20164
rect 7876 20114 7885 20164
rect 7911 20114 7928 20164
rect 7928 20114 7967 20164
rect 7829 20108 7885 20114
rect 7911 20108 7967 20114
rect 7993 20116 8047 20164
rect 8047 20116 8049 20164
rect 8075 20116 8099 20164
rect 8099 20116 8131 20164
rect 7993 20108 8049 20116
rect 8075 20108 8131 20116
rect 8157 20116 8169 20164
rect 8169 20116 8213 20164
rect 8157 20108 8213 20116
rect 2733 19931 2789 19987
rect 2814 19931 2870 19987
rect 2895 19931 2951 19987
rect 2976 19931 3032 19987
rect 3057 19931 3113 19987
rect 3138 19931 3194 19987
rect 3219 19931 3275 19987
rect 3300 19931 3356 19987
rect 3381 19931 3437 19987
rect 3462 19931 3518 19987
rect 3543 19931 3599 19987
rect 3624 19931 3680 19987
rect 3705 19931 3761 19987
rect 3786 19931 3842 19987
rect 3867 19931 3923 19987
rect 3948 19931 4004 19987
rect 4029 19931 4085 19987
rect 4110 19931 4166 19987
rect 4191 19931 4247 19987
rect 4272 19931 4328 19987
rect 4353 19931 4409 19987
rect 4434 19931 4490 19987
rect 4515 19931 4571 19987
rect 4596 19931 4652 19987
rect 4677 19931 4733 19987
rect 4758 19931 4814 19987
rect 4839 19931 4895 19987
rect 4920 19931 4976 19987
rect 5001 19931 5057 19987
rect 5082 19931 5138 19987
rect 2733 19851 2789 19907
rect 2814 19851 2870 19907
rect 2895 19851 2951 19907
rect 2976 19851 3032 19907
rect 3057 19851 3113 19907
rect 3138 19851 3194 19907
rect 3219 19851 3275 19907
rect 3300 19851 3356 19907
rect 3381 19851 3437 19907
rect 3462 19851 3518 19907
rect 3543 19851 3599 19907
rect 3624 19851 3680 19907
rect 3705 19851 3761 19907
rect 3786 19851 3842 19907
rect 3867 19851 3923 19907
rect 3948 19851 4004 19907
rect 4029 19851 4085 19907
rect 4110 19851 4166 19907
rect 4191 19851 4247 19907
rect 4272 19851 4328 19907
rect 4353 19851 4409 19907
rect 4434 19851 4490 19907
rect 4515 19851 4571 19907
rect 4596 19851 4652 19907
rect 4677 19851 4733 19907
rect 4758 19851 4814 19907
rect 4839 19851 4895 19907
rect 4920 19851 4976 19907
rect 5001 19851 5057 19907
rect 5082 19851 5138 19907
rect 2733 19771 2789 19827
rect 2814 19771 2870 19827
rect 2895 19771 2951 19827
rect 2976 19771 3032 19827
rect 3057 19771 3113 19827
rect 3138 19771 3194 19827
rect 3219 19771 3275 19827
rect 3300 19771 3356 19827
rect 3381 19771 3437 19827
rect 3462 19771 3518 19827
rect 3543 19771 3599 19827
rect 3624 19771 3680 19827
rect 3705 19771 3761 19827
rect 3786 19771 3842 19827
rect 3867 19771 3923 19827
rect 3948 19771 4004 19827
rect 4029 19771 4085 19827
rect 4110 19771 4166 19827
rect 4191 19771 4247 19827
rect 4272 19771 4328 19827
rect 4353 19771 4409 19827
rect 4434 19771 4490 19827
rect 4515 19771 4571 19827
rect 4596 19771 4652 19827
rect 4677 19771 4733 19827
rect 4758 19771 4814 19827
rect 4839 19771 4895 19827
rect 4920 19771 4976 19827
rect 5001 19771 5057 19827
rect 5082 19771 5138 19827
rect 2733 19691 2789 19747
rect 2814 19691 2870 19747
rect 2895 19691 2951 19747
rect 2976 19691 3032 19747
rect 3057 19691 3113 19747
rect 3138 19691 3194 19747
rect 3219 19691 3275 19747
rect 3300 19691 3356 19747
rect 3381 19691 3437 19747
rect 3462 19691 3518 19747
rect 3543 19691 3599 19747
rect 3624 19691 3680 19747
rect 3705 19691 3761 19747
rect 3786 19691 3842 19747
rect 3867 19691 3923 19747
rect 3948 19691 4004 19747
rect 4029 19691 4085 19747
rect 4110 19691 4166 19747
rect 4191 19691 4247 19747
rect 4272 19691 4328 19747
rect 4353 19691 4409 19747
rect 4434 19691 4490 19747
rect 4515 19691 4571 19747
rect 4596 19691 4652 19747
rect 4677 19691 4733 19747
rect 4758 19691 4814 19747
rect 4839 19691 4895 19747
rect 4920 19691 4976 19747
rect 5001 19691 5057 19747
rect 5082 19691 5138 19747
rect 2733 19611 2789 19667
rect 2814 19611 2870 19667
rect 2895 19611 2951 19667
rect 2976 19611 3032 19667
rect 3057 19611 3113 19667
rect 3138 19611 3194 19667
rect 3219 19611 3275 19667
rect 3300 19611 3356 19667
rect 3381 19611 3437 19667
rect 3462 19611 3518 19667
rect 3543 19611 3599 19667
rect 3624 19611 3680 19667
rect 3705 19611 3761 19667
rect 3786 19611 3842 19667
rect 3867 19611 3923 19667
rect 3948 19611 4004 19667
rect 4029 19611 4085 19667
rect 4110 19611 4166 19667
rect 4191 19611 4247 19667
rect 4272 19611 4328 19667
rect 4353 19611 4409 19667
rect 4434 19611 4490 19667
rect 4515 19611 4571 19667
rect 4596 19611 4652 19667
rect 4677 19611 4733 19667
rect 4758 19611 4814 19667
rect 4839 19611 4895 19667
rect 4920 19611 4976 19667
rect 5001 19611 5057 19667
rect 5082 19611 5138 19667
rect 2733 19531 2789 19587
rect 2814 19531 2870 19587
rect 2895 19531 2951 19587
rect 2976 19531 3032 19587
rect 3057 19531 3113 19587
rect 3138 19531 3194 19587
rect 3219 19531 3275 19587
rect 3300 19531 3356 19587
rect 3381 19531 3437 19587
rect 3462 19531 3518 19587
rect 3543 19531 3599 19587
rect 3624 19531 3680 19587
rect 3705 19531 3761 19587
rect 3786 19531 3842 19587
rect 3867 19531 3923 19587
rect 3948 19531 4004 19587
rect 4029 19531 4085 19587
rect 4110 19531 4166 19587
rect 4191 19531 4247 19587
rect 4272 19531 4328 19587
rect 4353 19531 4409 19587
rect 4434 19531 4490 19587
rect 4515 19531 4571 19587
rect 4596 19531 4652 19587
rect 4677 19531 4733 19587
rect 4758 19531 4814 19587
rect 4839 19531 4895 19587
rect 4920 19531 4976 19587
rect 5001 19531 5057 19587
rect 5082 19531 5138 19587
rect 2733 19451 2789 19507
rect 2814 19451 2870 19507
rect 2895 19451 2951 19507
rect 2976 19451 3032 19507
rect 3057 19451 3113 19507
rect 3138 19451 3194 19507
rect 3219 19451 3275 19507
rect 3300 19451 3356 19507
rect 3381 19451 3437 19507
rect 3462 19451 3518 19507
rect 3543 19451 3599 19507
rect 3624 19451 3680 19507
rect 3705 19451 3761 19507
rect 3786 19451 3842 19507
rect 3867 19451 3923 19507
rect 3948 19451 4004 19507
rect 4029 19451 4085 19507
rect 4110 19451 4166 19507
rect 4191 19451 4247 19507
rect 4272 19451 4328 19507
rect 4353 19451 4409 19507
rect 4434 19451 4490 19507
rect 4515 19451 4571 19507
rect 4596 19451 4652 19507
rect 4677 19451 4733 19507
rect 4758 19451 4814 19507
rect 4839 19451 4895 19507
rect 4920 19451 4976 19507
rect 5001 19451 5057 19507
rect 5082 19451 5138 19507
rect 2733 19371 2789 19427
rect 2814 19371 2870 19427
rect 2895 19371 2951 19427
rect 2976 19371 3032 19427
rect 3057 19371 3113 19427
rect 3138 19371 3194 19427
rect 3219 19371 3275 19427
rect 3300 19371 3356 19427
rect 3381 19371 3437 19427
rect 3462 19371 3518 19427
rect 3543 19371 3599 19427
rect 3624 19371 3680 19427
rect 3705 19371 3761 19427
rect 3786 19371 3842 19427
rect 3867 19371 3923 19427
rect 3948 19371 4004 19427
rect 4029 19371 4085 19427
rect 4110 19371 4166 19427
rect 4191 19371 4247 19427
rect 4272 19371 4328 19427
rect 4353 19371 4409 19427
rect 4434 19371 4490 19427
rect 4515 19371 4571 19427
rect 4596 19371 4652 19427
rect 4677 19371 4733 19427
rect 4758 19371 4814 19427
rect 4839 19371 4895 19427
rect 4920 19371 4976 19427
rect 5001 19371 5057 19427
rect 5082 19371 5138 19427
rect 5163 19371 5299 19987
rect 5613 18720 5669 18724
rect 5696 18720 5752 18724
rect 5613 18668 5646 18720
rect 5646 18668 5660 18720
rect 5660 18668 5669 18720
rect 5696 18668 5712 18720
rect 5712 18668 5752 18720
rect 5779 18668 5835 18724
rect 5861 18668 5917 18724
rect 5943 18668 5999 18724
rect 6025 18668 6081 18724
rect 6107 18720 6163 18724
rect 6189 18720 6245 18724
rect 6107 18668 6148 18720
rect 6148 18668 6163 18720
rect 6189 18668 6200 18720
rect 6200 18668 6214 18720
rect 6214 18668 6245 18720
rect 6271 18668 6327 18724
rect 6353 18668 6409 18724
rect 6435 18668 6491 18724
rect 6517 18668 6573 18724
rect 6599 18668 6655 18724
rect 6681 18720 6737 18724
rect 6763 18720 6819 18724
rect 6681 18668 6702 18720
rect 6702 18668 6737 18720
rect 6763 18668 6768 18720
rect 6768 18668 6819 18720
rect 6845 18668 6901 18724
rect 6927 18668 6983 18724
rect 7009 18668 7065 18724
rect 7091 18668 7147 18724
rect 7173 18668 7229 18724
rect 7255 18720 7311 18724
rect 7337 18720 7393 18724
rect 7255 18668 7256 18720
rect 7256 18668 7308 18720
rect 7308 18668 7311 18720
rect 7337 18668 7374 18720
rect 7374 18668 7393 18720
rect 7419 18668 7475 18724
rect 7501 18668 7557 18724
rect 7583 18668 7639 18724
rect 7665 18668 7721 18724
rect 7747 18668 7803 18724
rect 7829 18720 7885 18724
rect 7911 18720 7967 18724
rect 7829 18668 7862 18720
rect 7862 18668 7876 18720
rect 7876 18668 7885 18720
rect 7911 18668 7928 18720
rect 7928 18668 7967 18720
rect 7993 18672 8047 18724
rect 8047 18672 8049 18724
rect 8075 18672 8099 18724
rect 8099 18672 8131 18724
rect 7993 18668 8049 18672
rect 8075 18668 8131 18672
rect 8157 18672 8169 18724
rect 8169 18672 8213 18724
rect 8157 18668 8213 18672
rect 5613 18599 5646 18644
rect 5646 18599 5660 18644
rect 5660 18599 5669 18644
rect 5696 18599 5712 18644
rect 5712 18599 5752 18644
rect 5613 18588 5669 18599
rect 5696 18588 5752 18599
rect 5779 18588 5835 18644
rect 5861 18588 5917 18644
rect 5943 18588 5999 18644
rect 6025 18588 6081 18644
rect 6107 18599 6148 18644
rect 6148 18599 6163 18644
rect 6189 18599 6200 18644
rect 6200 18599 6214 18644
rect 6214 18599 6245 18644
rect 6107 18588 6163 18599
rect 6189 18588 6245 18599
rect 6271 18588 6327 18644
rect 6353 18588 6409 18644
rect 6435 18588 6491 18644
rect 6517 18588 6573 18644
rect 6599 18588 6655 18644
rect 6681 18599 6702 18644
rect 6702 18599 6737 18644
rect 6763 18599 6768 18644
rect 6768 18599 6819 18644
rect 6681 18588 6737 18599
rect 6763 18588 6819 18599
rect 6845 18588 6901 18644
rect 6927 18588 6983 18644
rect 7009 18588 7065 18644
rect 7091 18588 7147 18644
rect 7173 18588 7229 18644
rect 7255 18599 7256 18644
rect 7256 18599 7308 18644
rect 7308 18599 7311 18644
rect 7337 18599 7374 18644
rect 7374 18599 7393 18644
rect 7255 18588 7311 18599
rect 7337 18588 7393 18599
rect 7419 18588 7475 18644
rect 7501 18588 7557 18644
rect 7583 18588 7639 18644
rect 7665 18588 7721 18644
rect 7747 18588 7803 18644
rect 7829 18599 7862 18644
rect 7862 18599 7876 18644
rect 7876 18599 7885 18644
rect 7911 18599 7928 18644
rect 7928 18599 7967 18644
rect 7829 18588 7885 18599
rect 7911 18588 7967 18599
rect 7993 18603 8047 18644
rect 8047 18603 8049 18644
rect 8075 18603 8099 18644
rect 8099 18603 8131 18644
rect 7993 18588 8049 18603
rect 8075 18588 8131 18603
rect 8157 18603 8169 18644
rect 8169 18603 8213 18644
rect 8157 18588 8213 18603
rect 5613 18530 5646 18564
rect 5646 18530 5660 18564
rect 5660 18530 5669 18564
rect 5696 18530 5712 18564
rect 5712 18530 5752 18564
rect 5613 18513 5669 18530
rect 5696 18513 5752 18530
rect 5613 18508 5646 18513
rect 5646 18508 5660 18513
rect 5660 18508 5669 18513
rect 5696 18508 5712 18513
rect 5712 18508 5752 18513
rect 5779 18508 5835 18564
rect 5861 18508 5917 18564
rect 5943 18508 5999 18564
rect 6025 18508 6081 18564
rect 6107 18530 6148 18564
rect 6148 18530 6163 18564
rect 6189 18530 6200 18564
rect 6200 18530 6214 18564
rect 6214 18530 6245 18564
rect 6107 18513 6163 18530
rect 6189 18513 6245 18530
rect 6107 18508 6148 18513
rect 6148 18508 6163 18513
rect 6189 18508 6200 18513
rect 6200 18508 6214 18513
rect 6214 18508 6245 18513
rect 6271 18508 6327 18564
rect 6353 18508 6409 18564
rect 6435 18508 6491 18564
rect 6517 18508 6573 18564
rect 6599 18508 6655 18564
rect 6681 18530 6702 18564
rect 6702 18530 6737 18564
rect 6763 18530 6768 18564
rect 6768 18530 6819 18564
rect 6681 18513 6737 18530
rect 6763 18513 6819 18530
rect 6681 18508 6702 18513
rect 6702 18508 6737 18513
rect 6763 18508 6768 18513
rect 6768 18508 6819 18513
rect 6845 18508 6901 18564
rect 6927 18508 6983 18564
rect 7009 18508 7065 18564
rect 7091 18508 7147 18564
rect 7173 18508 7229 18564
rect 7255 18530 7256 18564
rect 7256 18530 7308 18564
rect 7308 18530 7311 18564
rect 7337 18530 7374 18564
rect 7374 18530 7393 18564
rect 7255 18513 7311 18530
rect 7337 18513 7393 18530
rect 7255 18508 7256 18513
rect 7256 18508 7308 18513
rect 7308 18508 7311 18513
rect 7337 18508 7374 18513
rect 7374 18508 7393 18513
rect 7419 18508 7475 18564
rect 7501 18508 7557 18564
rect 7583 18508 7639 18564
rect 7665 18508 7721 18564
rect 7747 18508 7803 18564
rect 7829 18530 7862 18564
rect 7862 18530 7876 18564
rect 7876 18530 7885 18564
rect 7911 18530 7928 18564
rect 7928 18530 7967 18564
rect 7829 18513 7885 18530
rect 7911 18513 7967 18530
rect 7829 18508 7862 18513
rect 7862 18508 7876 18513
rect 7876 18508 7885 18513
rect 7911 18508 7928 18513
rect 7928 18508 7967 18513
rect 7993 18534 8047 18564
rect 8047 18534 8049 18564
rect 8075 18534 8099 18564
rect 8099 18534 8131 18564
rect 7993 18517 8049 18534
rect 8075 18517 8131 18534
rect 7993 18508 8047 18517
rect 8047 18508 8049 18517
rect 8075 18508 8099 18517
rect 8099 18508 8131 18517
rect 8157 18534 8169 18564
rect 8169 18534 8213 18564
rect 8157 18517 8213 18534
rect 8157 18508 8169 18517
rect 8169 18508 8213 18517
rect 5613 18461 5646 18484
rect 5646 18461 5660 18484
rect 5660 18461 5669 18484
rect 5696 18461 5712 18484
rect 5712 18461 5752 18484
rect 5613 18444 5669 18461
rect 5696 18444 5752 18461
rect 5613 18428 5646 18444
rect 5646 18428 5660 18444
rect 5660 18428 5669 18444
rect 5696 18428 5712 18444
rect 5712 18428 5752 18444
rect 5779 18428 5835 18484
rect 5861 18428 5917 18484
rect 5943 18428 5999 18484
rect 6025 18428 6081 18484
rect 6107 18461 6148 18484
rect 6148 18461 6163 18484
rect 6189 18461 6200 18484
rect 6200 18461 6214 18484
rect 6214 18461 6245 18484
rect 6107 18444 6163 18461
rect 6189 18444 6245 18461
rect 6107 18428 6148 18444
rect 6148 18428 6163 18444
rect 6189 18428 6200 18444
rect 6200 18428 6214 18444
rect 6214 18428 6245 18444
rect 6271 18428 6327 18484
rect 6353 18428 6409 18484
rect 6435 18428 6491 18484
rect 6517 18428 6573 18484
rect 6599 18428 6655 18484
rect 6681 18461 6702 18484
rect 6702 18461 6737 18484
rect 6763 18461 6768 18484
rect 6768 18461 6819 18484
rect 6681 18444 6737 18461
rect 6763 18444 6819 18461
rect 6681 18428 6702 18444
rect 6702 18428 6737 18444
rect 6763 18428 6768 18444
rect 6768 18428 6819 18444
rect 6845 18428 6901 18484
rect 6927 18428 6983 18484
rect 7009 18428 7065 18484
rect 7091 18428 7147 18484
rect 7173 18428 7229 18484
rect 7255 18461 7256 18484
rect 7256 18461 7308 18484
rect 7308 18461 7311 18484
rect 7337 18461 7374 18484
rect 7374 18461 7393 18484
rect 7255 18444 7311 18461
rect 7337 18444 7393 18461
rect 7255 18428 7256 18444
rect 7256 18428 7308 18444
rect 7308 18428 7311 18444
rect 7337 18428 7374 18444
rect 7374 18428 7393 18444
rect 7419 18428 7475 18484
rect 7501 18428 7557 18484
rect 7583 18428 7639 18484
rect 7665 18428 7721 18484
rect 7747 18428 7803 18484
rect 7829 18461 7862 18484
rect 7862 18461 7876 18484
rect 7876 18461 7885 18484
rect 7911 18461 7928 18484
rect 7928 18461 7967 18484
rect 7829 18444 7885 18461
rect 7911 18444 7967 18461
rect 7829 18428 7862 18444
rect 7862 18428 7876 18444
rect 7876 18428 7885 18444
rect 7911 18428 7928 18444
rect 7928 18428 7967 18444
rect 7993 18465 8047 18484
rect 8047 18465 8049 18484
rect 8075 18465 8099 18484
rect 8099 18465 8131 18484
rect 7993 18448 8049 18465
rect 8075 18448 8131 18465
rect 7993 18428 8047 18448
rect 8047 18428 8049 18448
rect 8075 18428 8099 18448
rect 8099 18428 8131 18448
rect 8157 18465 8169 18484
rect 8169 18465 8213 18484
rect 8157 18448 8213 18465
rect 8157 18428 8169 18448
rect 8169 18428 8213 18448
rect 5613 18392 5646 18404
rect 5646 18392 5660 18404
rect 5660 18392 5669 18404
rect 5696 18392 5712 18404
rect 5712 18392 5752 18404
rect 5613 18375 5669 18392
rect 5696 18375 5752 18392
rect 5613 18348 5646 18375
rect 5646 18348 5660 18375
rect 5660 18348 5669 18375
rect 5696 18348 5712 18375
rect 5712 18348 5752 18375
rect 5779 18348 5835 18404
rect 5861 18348 5917 18404
rect 5943 18348 5999 18404
rect 6025 18348 6081 18404
rect 6107 18392 6148 18404
rect 6148 18392 6163 18404
rect 6189 18392 6200 18404
rect 6200 18392 6214 18404
rect 6214 18392 6245 18404
rect 6107 18375 6163 18392
rect 6189 18375 6245 18392
rect 6107 18348 6148 18375
rect 6148 18348 6163 18375
rect 6189 18348 6200 18375
rect 6200 18348 6214 18375
rect 6214 18348 6245 18375
rect 6271 18348 6327 18404
rect 6353 18348 6409 18404
rect 6435 18348 6491 18404
rect 6517 18348 6573 18404
rect 6599 18348 6655 18404
rect 6681 18392 6702 18404
rect 6702 18392 6737 18404
rect 6763 18392 6768 18404
rect 6768 18392 6819 18404
rect 6681 18375 6737 18392
rect 6763 18375 6819 18392
rect 6681 18348 6702 18375
rect 6702 18348 6737 18375
rect 6763 18348 6768 18375
rect 6768 18348 6819 18375
rect 6845 18348 6901 18404
rect 6927 18348 6983 18404
rect 7009 18348 7065 18404
rect 7091 18348 7147 18404
rect 7173 18348 7229 18404
rect 7255 18392 7256 18404
rect 7256 18392 7308 18404
rect 7308 18392 7311 18404
rect 7337 18392 7374 18404
rect 7374 18392 7393 18404
rect 7255 18375 7311 18392
rect 7337 18375 7393 18392
rect 7255 18348 7256 18375
rect 7256 18348 7308 18375
rect 7308 18348 7311 18375
rect 7337 18348 7374 18375
rect 7374 18348 7393 18375
rect 7419 18348 7475 18404
rect 7501 18348 7557 18404
rect 7583 18348 7639 18404
rect 7665 18348 7721 18404
rect 7747 18348 7803 18404
rect 7829 18392 7862 18404
rect 7862 18392 7876 18404
rect 7876 18392 7885 18404
rect 7911 18392 7928 18404
rect 7928 18392 7967 18404
rect 7829 18375 7885 18392
rect 7911 18375 7967 18392
rect 7829 18348 7862 18375
rect 7862 18348 7876 18375
rect 7876 18348 7885 18375
rect 7911 18348 7928 18375
rect 7928 18348 7967 18375
rect 7993 18396 8047 18404
rect 8047 18396 8049 18404
rect 8075 18396 8099 18404
rect 8099 18396 8131 18404
rect 7993 18378 8049 18396
rect 8075 18378 8131 18396
rect 7993 18348 8047 18378
rect 8047 18348 8049 18378
rect 8075 18348 8099 18378
rect 8099 18348 8131 18378
rect 8157 18396 8169 18404
rect 8169 18396 8213 18404
rect 8157 18378 8213 18396
rect 8157 18348 8169 18378
rect 8169 18348 8213 18378
rect 5613 18323 5646 18324
rect 5646 18323 5660 18324
rect 5660 18323 5669 18324
rect 5696 18323 5712 18324
rect 5712 18323 5752 18324
rect 5613 18306 5669 18323
rect 5696 18306 5752 18323
rect 5613 18268 5646 18306
rect 5646 18268 5660 18306
rect 5660 18268 5669 18306
rect 5696 18268 5712 18306
rect 5712 18268 5752 18306
rect 5779 18268 5835 18324
rect 5861 18268 5917 18324
rect 5943 18268 5999 18324
rect 6025 18268 6081 18324
rect 6107 18323 6148 18324
rect 6148 18323 6163 18324
rect 6189 18323 6200 18324
rect 6200 18323 6214 18324
rect 6214 18323 6245 18324
rect 6107 18306 6163 18323
rect 6189 18306 6245 18323
rect 6107 18268 6148 18306
rect 6148 18268 6163 18306
rect 6189 18268 6200 18306
rect 6200 18268 6214 18306
rect 6214 18268 6245 18306
rect 6271 18268 6327 18324
rect 6353 18268 6409 18324
rect 6435 18268 6491 18324
rect 6517 18268 6573 18324
rect 6599 18268 6655 18324
rect 6681 18323 6702 18324
rect 6702 18323 6737 18324
rect 6763 18323 6768 18324
rect 6768 18323 6819 18324
rect 6681 18306 6737 18323
rect 6763 18306 6819 18323
rect 6681 18268 6702 18306
rect 6702 18268 6737 18306
rect 6763 18268 6768 18306
rect 6768 18268 6819 18306
rect 6845 18268 6901 18324
rect 6927 18268 6983 18324
rect 7009 18268 7065 18324
rect 7091 18268 7147 18324
rect 7173 18268 7229 18324
rect 7255 18323 7256 18324
rect 7256 18323 7308 18324
rect 7308 18323 7311 18324
rect 7337 18323 7374 18324
rect 7374 18323 7393 18324
rect 7255 18306 7311 18323
rect 7337 18306 7393 18323
rect 7255 18268 7256 18306
rect 7256 18268 7308 18306
rect 7308 18268 7311 18306
rect 7337 18268 7374 18306
rect 7374 18268 7393 18306
rect 7419 18268 7475 18324
rect 7501 18268 7557 18324
rect 7583 18268 7639 18324
rect 7665 18268 7721 18324
rect 7747 18268 7803 18324
rect 7829 18323 7862 18324
rect 7862 18323 7876 18324
rect 7876 18323 7885 18324
rect 7911 18323 7928 18324
rect 7928 18323 7967 18324
rect 7829 18306 7885 18323
rect 7911 18306 7967 18323
rect 7829 18268 7862 18306
rect 7862 18268 7876 18306
rect 7876 18268 7885 18306
rect 7911 18268 7928 18306
rect 7928 18268 7967 18306
rect 7993 18308 8049 18324
rect 8075 18308 8131 18324
rect 7993 18268 8047 18308
rect 8047 18268 8049 18308
rect 8075 18268 8099 18308
rect 8099 18268 8131 18308
rect 8157 18308 8213 18324
rect 8157 18268 8169 18308
rect 8169 18268 8213 18308
rect 5613 18236 5669 18244
rect 5696 18236 5752 18244
rect 5613 18188 5646 18236
rect 5646 18188 5660 18236
rect 5660 18188 5669 18236
rect 5696 18188 5712 18236
rect 5712 18188 5752 18236
rect 5779 18188 5835 18244
rect 5861 18188 5917 18244
rect 5943 18188 5999 18244
rect 6025 18188 6081 18244
rect 6107 18236 6163 18244
rect 6189 18236 6245 18244
rect 6107 18188 6148 18236
rect 6148 18188 6163 18236
rect 6189 18188 6200 18236
rect 6200 18188 6214 18236
rect 6214 18188 6245 18236
rect 6271 18188 6327 18244
rect 6353 18188 6409 18244
rect 6435 18188 6491 18244
rect 6517 18188 6573 18244
rect 6599 18188 6655 18244
rect 6681 18236 6737 18244
rect 6763 18236 6819 18244
rect 6681 18188 6702 18236
rect 6702 18188 6737 18236
rect 6763 18188 6768 18236
rect 6768 18188 6819 18236
rect 6845 18188 6901 18244
rect 6927 18188 6983 18244
rect 7009 18188 7065 18244
rect 7091 18188 7147 18244
rect 7173 18188 7229 18244
rect 7255 18236 7311 18244
rect 7337 18236 7393 18244
rect 7255 18188 7256 18236
rect 7256 18188 7308 18236
rect 7308 18188 7311 18236
rect 7337 18188 7374 18236
rect 7374 18188 7393 18236
rect 7419 18188 7475 18244
rect 7501 18188 7557 18244
rect 7583 18188 7639 18244
rect 7665 18188 7721 18244
rect 7747 18188 7803 18244
rect 7829 18236 7885 18244
rect 7911 18236 7967 18244
rect 7829 18188 7862 18236
rect 7862 18188 7876 18236
rect 7876 18188 7885 18236
rect 7911 18188 7928 18236
rect 7928 18188 7967 18236
rect 7993 18238 8049 18244
rect 8075 18238 8131 18244
rect 7993 18188 8047 18238
rect 8047 18188 8049 18238
rect 8075 18188 8099 18238
rect 8099 18188 8131 18238
rect 8157 18238 8213 18244
rect 8157 18188 8169 18238
rect 8169 18188 8213 18238
rect 5613 18114 5646 18164
rect 5646 18114 5660 18164
rect 5660 18114 5669 18164
rect 5696 18114 5712 18164
rect 5712 18114 5752 18164
rect 5613 18108 5669 18114
rect 5696 18108 5752 18114
rect 5779 18108 5835 18164
rect 5861 18108 5917 18164
rect 5943 18108 5999 18164
rect 6025 18108 6081 18164
rect 6107 18114 6148 18164
rect 6148 18114 6163 18164
rect 6189 18114 6200 18164
rect 6200 18114 6214 18164
rect 6214 18114 6245 18164
rect 6107 18108 6163 18114
rect 6189 18108 6245 18114
rect 6271 18108 6327 18164
rect 6353 18108 6409 18164
rect 6435 18108 6491 18164
rect 6517 18108 6573 18164
rect 6599 18108 6655 18164
rect 6681 18114 6702 18164
rect 6702 18114 6737 18164
rect 6763 18114 6768 18164
rect 6768 18114 6819 18164
rect 6681 18108 6737 18114
rect 6763 18108 6819 18114
rect 6845 18108 6901 18164
rect 6927 18108 6983 18164
rect 7009 18108 7065 18164
rect 7091 18108 7147 18164
rect 7173 18108 7229 18164
rect 7255 18114 7256 18164
rect 7256 18114 7308 18164
rect 7308 18114 7311 18164
rect 7337 18114 7374 18164
rect 7374 18114 7393 18164
rect 7255 18108 7311 18114
rect 7337 18108 7393 18114
rect 7419 18108 7475 18164
rect 7501 18108 7557 18164
rect 7583 18108 7639 18164
rect 7665 18108 7721 18164
rect 7747 18108 7803 18164
rect 7829 18114 7862 18164
rect 7862 18114 7876 18164
rect 7876 18114 7885 18164
rect 7911 18114 7928 18164
rect 7928 18114 7967 18164
rect 7829 18108 7885 18114
rect 7911 18108 7967 18114
rect 7993 18116 8047 18164
rect 8047 18116 8049 18164
rect 8075 18116 8099 18164
rect 8099 18116 8131 18164
rect 7993 18108 8049 18116
rect 8075 18108 8131 18116
rect 8157 18116 8169 18164
rect 8169 18116 8213 18164
rect 8157 18108 8213 18116
rect 2733 17931 2789 17987
rect 2814 17931 2870 17987
rect 2895 17931 2951 17987
rect 2976 17931 3032 17987
rect 3057 17931 3113 17987
rect 3138 17931 3194 17987
rect 3219 17931 3275 17987
rect 3300 17931 3356 17987
rect 3381 17931 3437 17987
rect 3462 17931 3518 17987
rect 3543 17931 3599 17987
rect 3624 17931 3680 17987
rect 3705 17931 3761 17987
rect 3786 17931 3842 17987
rect 3867 17931 3923 17987
rect 3948 17931 4004 17987
rect 4029 17931 4085 17987
rect 4110 17931 4166 17987
rect 4191 17931 4247 17987
rect 4272 17931 4328 17987
rect 4353 17931 4409 17987
rect 4434 17931 4490 17987
rect 4515 17931 4571 17987
rect 4596 17931 4652 17987
rect 4677 17931 4733 17987
rect 4758 17931 4814 17987
rect 4839 17931 4895 17987
rect 4920 17931 4976 17987
rect 5001 17931 5057 17987
rect 5082 17931 5138 17987
rect 2733 17851 2789 17907
rect 2814 17851 2870 17907
rect 2895 17851 2951 17907
rect 2976 17851 3032 17907
rect 3057 17851 3113 17907
rect 3138 17851 3194 17907
rect 3219 17851 3275 17907
rect 3300 17851 3356 17907
rect 3381 17851 3437 17907
rect 3462 17851 3518 17907
rect 3543 17851 3599 17907
rect 3624 17851 3680 17907
rect 3705 17851 3761 17907
rect 3786 17851 3842 17907
rect 3867 17851 3923 17907
rect 3948 17851 4004 17907
rect 4029 17851 4085 17907
rect 4110 17851 4166 17907
rect 4191 17851 4247 17907
rect 4272 17851 4328 17907
rect 4353 17851 4409 17907
rect 4434 17851 4490 17907
rect 4515 17851 4571 17907
rect 4596 17851 4652 17907
rect 4677 17851 4733 17907
rect 4758 17851 4814 17907
rect 4839 17851 4895 17907
rect 4920 17851 4976 17907
rect 5001 17851 5057 17907
rect 5082 17851 5138 17907
rect 2733 17771 2789 17827
rect 2814 17771 2870 17827
rect 2895 17771 2951 17827
rect 2976 17771 3032 17827
rect 3057 17771 3113 17827
rect 3138 17771 3194 17827
rect 3219 17771 3275 17827
rect 3300 17771 3356 17827
rect 3381 17771 3437 17827
rect 3462 17771 3518 17827
rect 3543 17771 3599 17827
rect 3624 17771 3680 17827
rect 3705 17771 3761 17827
rect 3786 17771 3842 17827
rect 3867 17771 3923 17827
rect 3948 17771 4004 17827
rect 4029 17771 4085 17827
rect 4110 17771 4166 17827
rect 4191 17771 4247 17827
rect 4272 17771 4328 17827
rect 4353 17771 4409 17827
rect 4434 17771 4490 17827
rect 4515 17771 4571 17827
rect 4596 17771 4652 17827
rect 4677 17771 4733 17827
rect 4758 17771 4814 17827
rect 4839 17771 4895 17827
rect 4920 17771 4976 17827
rect 5001 17771 5057 17827
rect 5082 17771 5138 17827
rect 2733 17691 2789 17747
rect 2814 17691 2870 17747
rect 2895 17691 2951 17747
rect 2976 17691 3032 17747
rect 3057 17691 3113 17747
rect 3138 17691 3194 17747
rect 3219 17691 3275 17747
rect 3300 17691 3356 17747
rect 3381 17691 3437 17747
rect 3462 17691 3518 17747
rect 3543 17691 3599 17747
rect 3624 17691 3680 17747
rect 3705 17691 3761 17747
rect 3786 17691 3842 17747
rect 3867 17691 3923 17747
rect 3948 17691 4004 17747
rect 4029 17691 4085 17747
rect 4110 17691 4166 17747
rect 4191 17691 4247 17747
rect 4272 17691 4328 17747
rect 4353 17691 4409 17747
rect 4434 17691 4490 17747
rect 4515 17691 4571 17747
rect 4596 17691 4652 17747
rect 4677 17691 4733 17747
rect 4758 17691 4814 17747
rect 4839 17691 4895 17747
rect 4920 17691 4976 17747
rect 5001 17691 5057 17747
rect 5082 17691 5138 17747
rect 2733 17611 2789 17667
rect 2814 17611 2870 17667
rect 2895 17611 2951 17667
rect 2976 17611 3032 17667
rect 3057 17611 3113 17667
rect 3138 17611 3194 17667
rect 3219 17611 3275 17667
rect 3300 17611 3356 17667
rect 3381 17611 3437 17667
rect 3462 17611 3518 17667
rect 3543 17611 3599 17667
rect 3624 17611 3680 17667
rect 3705 17611 3761 17667
rect 3786 17611 3842 17667
rect 3867 17611 3923 17667
rect 3948 17611 4004 17667
rect 4029 17611 4085 17667
rect 4110 17611 4166 17667
rect 4191 17611 4247 17667
rect 4272 17611 4328 17667
rect 4353 17611 4409 17667
rect 4434 17611 4490 17667
rect 4515 17611 4571 17667
rect 4596 17611 4652 17667
rect 4677 17611 4733 17667
rect 4758 17611 4814 17667
rect 4839 17611 4895 17667
rect 4920 17611 4976 17667
rect 5001 17611 5057 17667
rect 5082 17611 5138 17667
rect 2733 17531 2789 17587
rect 2814 17531 2870 17587
rect 2895 17531 2951 17587
rect 2976 17531 3032 17587
rect 3057 17531 3113 17587
rect 3138 17531 3194 17587
rect 3219 17531 3275 17587
rect 3300 17531 3356 17587
rect 3381 17531 3437 17587
rect 3462 17531 3518 17587
rect 3543 17531 3599 17587
rect 3624 17531 3680 17587
rect 3705 17531 3761 17587
rect 3786 17531 3842 17587
rect 3867 17531 3923 17587
rect 3948 17531 4004 17587
rect 4029 17531 4085 17587
rect 4110 17531 4166 17587
rect 4191 17531 4247 17587
rect 4272 17531 4328 17587
rect 4353 17531 4409 17587
rect 4434 17531 4490 17587
rect 4515 17531 4571 17587
rect 4596 17531 4652 17587
rect 4677 17531 4733 17587
rect 4758 17531 4814 17587
rect 4839 17531 4895 17587
rect 4920 17531 4976 17587
rect 5001 17531 5057 17587
rect 5082 17531 5138 17587
rect 2733 17451 2789 17507
rect 2814 17451 2870 17507
rect 2895 17451 2951 17507
rect 2976 17451 3032 17507
rect 3057 17451 3113 17507
rect 3138 17451 3194 17507
rect 3219 17451 3275 17507
rect 3300 17451 3356 17507
rect 3381 17451 3437 17507
rect 3462 17451 3518 17507
rect 3543 17451 3599 17507
rect 3624 17451 3680 17507
rect 3705 17451 3761 17507
rect 3786 17451 3842 17507
rect 3867 17451 3923 17507
rect 3948 17451 4004 17507
rect 4029 17451 4085 17507
rect 4110 17451 4166 17507
rect 4191 17451 4247 17507
rect 4272 17451 4328 17507
rect 4353 17451 4409 17507
rect 4434 17451 4490 17507
rect 4515 17451 4571 17507
rect 4596 17451 4652 17507
rect 4677 17451 4733 17507
rect 4758 17451 4814 17507
rect 4839 17451 4895 17507
rect 4920 17451 4976 17507
rect 5001 17451 5057 17507
rect 5082 17451 5138 17507
rect 2733 17371 2789 17427
rect 2814 17371 2870 17427
rect 2895 17371 2951 17427
rect 2976 17371 3032 17427
rect 3057 17371 3113 17427
rect 3138 17371 3194 17427
rect 3219 17371 3275 17427
rect 3300 17371 3356 17427
rect 3381 17371 3437 17427
rect 3462 17371 3518 17427
rect 3543 17371 3599 17427
rect 3624 17371 3680 17427
rect 3705 17371 3761 17427
rect 3786 17371 3842 17427
rect 3867 17371 3923 17427
rect 3948 17371 4004 17427
rect 4029 17371 4085 17427
rect 4110 17371 4166 17427
rect 4191 17371 4247 17427
rect 4272 17371 4328 17427
rect 4353 17371 4409 17427
rect 4434 17371 4490 17427
rect 4515 17371 4571 17427
rect 4596 17371 4652 17427
rect 4677 17371 4733 17427
rect 4758 17371 4814 17427
rect 4839 17371 4895 17427
rect 4920 17371 4976 17427
rect 5001 17371 5057 17427
rect 5082 17371 5138 17427
rect 5163 17371 5299 17987
rect 5613 15452 5669 15456
rect 5696 15452 5752 15456
rect 5613 15400 5646 15452
rect 5646 15400 5660 15452
rect 5660 15400 5669 15452
rect 5696 15400 5712 15452
rect 5712 15400 5752 15452
rect 5779 15400 5835 15456
rect 5861 15400 5917 15456
rect 5943 15400 5999 15456
rect 6025 15400 6081 15456
rect 6107 15452 6163 15456
rect 6189 15452 6245 15456
rect 6107 15400 6148 15452
rect 6148 15400 6163 15452
rect 6189 15400 6200 15452
rect 6200 15400 6214 15452
rect 6214 15400 6245 15452
rect 6271 15400 6327 15456
rect 6353 15400 6409 15456
rect 6435 15400 6491 15456
rect 6517 15400 6573 15456
rect 6599 15400 6655 15456
rect 6681 15452 6737 15456
rect 6763 15452 6819 15456
rect 6681 15400 6702 15452
rect 6702 15400 6737 15452
rect 6763 15400 6768 15452
rect 6768 15400 6819 15452
rect 6845 15400 6901 15456
rect 6927 15400 6983 15456
rect 7009 15400 7065 15456
rect 7091 15400 7147 15456
rect 7173 15400 7229 15456
rect 7255 15452 7311 15456
rect 7337 15452 7393 15456
rect 7255 15400 7256 15452
rect 7256 15400 7308 15452
rect 7308 15400 7311 15452
rect 7337 15400 7374 15452
rect 7374 15400 7393 15452
rect 7419 15400 7475 15456
rect 7501 15400 7557 15456
rect 7583 15400 7639 15456
rect 7665 15400 7721 15456
rect 7747 15400 7803 15456
rect 7829 15452 7885 15456
rect 7911 15452 7967 15456
rect 7829 15400 7862 15452
rect 7862 15400 7876 15452
rect 7876 15400 7885 15452
rect 7911 15400 7928 15452
rect 7928 15400 7967 15452
rect 7993 15404 8047 15456
rect 8047 15404 8049 15456
rect 8075 15404 8099 15456
rect 8099 15404 8131 15456
rect 7993 15400 8049 15404
rect 8075 15400 8131 15404
rect 8157 15404 8169 15456
rect 8169 15404 8213 15456
rect 8157 15400 8213 15404
rect 5613 15331 5646 15376
rect 5646 15331 5660 15376
rect 5660 15331 5669 15376
rect 5696 15331 5712 15376
rect 5712 15331 5752 15376
rect 5613 15320 5669 15331
rect 5696 15320 5752 15331
rect 5779 15320 5835 15376
rect 5861 15320 5917 15376
rect 5943 15320 5999 15376
rect 6025 15320 6081 15376
rect 6107 15331 6148 15376
rect 6148 15331 6163 15376
rect 6189 15331 6200 15376
rect 6200 15331 6214 15376
rect 6214 15331 6245 15376
rect 6107 15320 6163 15331
rect 6189 15320 6245 15331
rect 6271 15320 6327 15376
rect 6353 15320 6409 15376
rect 6435 15320 6491 15376
rect 6517 15320 6573 15376
rect 6599 15320 6655 15376
rect 6681 15331 6702 15376
rect 6702 15331 6737 15376
rect 6763 15331 6768 15376
rect 6768 15331 6819 15376
rect 6681 15320 6737 15331
rect 6763 15320 6819 15331
rect 6845 15320 6901 15376
rect 6927 15320 6983 15376
rect 7009 15320 7065 15376
rect 7091 15320 7147 15376
rect 7173 15320 7229 15376
rect 7255 15331 7256 15376
rect 7256 15331 7308 15376
rect 7308 15331 7311 15376
rect 7337 15331 7374 15376
rect 7374 15331 7393 15376
rect 7255 15320 7311 15331
rect 7337 15320 7393 15331
rect 7419 15320 7475 15376
rect 7501 15320 7557 15376
rect 7583 15320 7639 15376
rect 7665 15320 7721 15376
rect 7747 15320 7803 15376
rect 7829 15331 7862 15376
rect 7862 15331 7876 15376
rect 7876 15331 7885 15376
rect 7911 15331 7928 15376
rect 7928 15331 7967 15376
rect 7829 15320 7885 15331
rect 7911 15320 7967 15331
rect 7993 15335 8047 15376
rect 8047 15335 8049 15376
rect 8075 15335 8099 15376
rect 8099 15335 8131 15376
rect 7993 15320 8049 15335
rect 8075 15320 8131 15335
rect 8157 15335 8169 15376
rect 8169 15335 8213 15376
rect 8157 15320 8213 15335
rect 5613 15262 5646 15296
rect 5646 15262 5660 15296
rect 5660 15262 5669 15296
rect 5696 15262 5712 15296
rect 5712 15262 5752 15296
rect 5613 15245 5669 15262
rect 5696 15245 5752 15262
rect 5613 15240 5646 15245
rect 5646 15240 5660 15245
rect 5660 15240 5669 15245
rect 5696 15240 5712 15245
rect 5712 15240 5752 15245
rect 5779 15240 5835 15296
rect 5861 15240 5917 15296
rect 5943 15240 5999 15296
rect 6025 15240 6081 15296
rect 6107 15262 6148 15296
rect 6148 15262 6163 15296
rect 6189 15262 6200 15296
rect 6200 15262 6214 15296
rect 6214 15262 6245 15296
rect 6107 15245 6163 15262
rect 6189 15245 6245 15262
rect 6107 15240 6148 15245
rect 6148 15240 6163 15245
rect 6189 15240 6200 15245
rect 6200 15240 6214 15245
rect 6214 15240 6245 15245
rect 6271 15240 6327 15296
rect 6353 15240 6409 15296
rect 6435 15240 6491 15296
rect 6517 15240 6573 15296
rect 6599 15240 6655 15296
rect 6681 15262 6702 15296
rect 6702 15262 6737 15296
rect 6763 15262 6768 15296
rect 6768 15262 6819 15296
rect 6681 15245 6737 15262
rect 6763 15245 6819 15262
rect 6681 15240 6702 15245
rect 6702 15240 6737 15245
rect 6763 15240 6768 15245
rect 6768 15240 6819 15245
rect 6845 15240 6901 15296
rect 6927 15240 6983 15296
rect 7009 15240 7065 15296
rect 7091 15240 7147 15296
rect 7173 15240 7229 15296
rect 7255 15262 7256 15296
rect 7256 15262 7308 15296
rect 7308 15262 7311 15296
rect 7337 15262 7374 15296
rect 7374 15262 7393 15296
rect 7255 15245 7311 15262
rect 7337 15245 7393 15262
rect 7255 15240 7256 15245
rect 7256 15240 7308 15245
rect 7308 15240 7311 15245
rect 7337 15240 7374 15245
rect 7374 15240 7393 15245
rect 7419 15240 7475 15296
rect 7501 15240 7557 15296
rect 7583 15240 7639 15296
rect 7665 15240 7721 15296
rect 7747 15240 7803 15296
rect 7829 15262 7862 15296
rect 7862 15262 7876 15296
rect 7876 15262 7885 15296
rect 7911 15262 7928 15296
rect 7928 15262 7967 15296
rect 7829 15245 7885 15262
rect 7911 15245 7967 15262
rect 7829 15240 7862 15245
rect 7862 15240 7876 15245
rect 7876 15240 7885 15245
rect 7911 15240 7928 15245
rect 7928 15240 7967 15245
rect 7993 15266 8047 15296
rect 8047 15266 8049 15296
rect 8075 15266 8099 15296
rect 8099 15266 8131 15296
rect 7993 15249 8049 15266
rect 8075 15249 8131 15266
rect 7993 15240 8047 15249
rect 8047 15240 8049 15249
rect 8075 15240 8099 15249
rect 8099 15240 8131 15249
rect 8157 15266 8169 15296
rect 8169 15266 8213 15296
rect 8157 15249 8213 15266
rect 8157 15240 8169 15249
rect 8169 15240 8213 15249
rect 5613 15193 5646 15216
rect 5646 15193 5660 15216
rect 5660 15193 5669 15216
rect 5696 15193 5712 15216
rect 5712 15193 5752 15216
rect 5613 15176 5669 15193
rect 5696 15176 5752 15193
rect 5613 15160 5646 15176
rect 5646 15160 5660 15176
rect 5660 15160 5669 15176
rect 5696 15160 5712 15176
rect 5712 15160 5752 15176
rect 5779 15160 5835 15216
rect 5861 15160 5917 15216
rect 5943 15160 5999 15216
rect 6025 15160 6081 15216
rect 6107 15193 6148 15216
rect 6148 15193 6163 15216
rect 6189 15193 6200 15216
rect 6200 15193 6214 15216
rect 6214 15193 6245 15216
rect 6107 15176 6163 15193
rect 6189 15176 6245 15193
rect 6107 15160 6148 15176
rect 6148 15160 6163 15176
rect 6189 15160 6200 15176
rect 6200 15160 6214 15176
rect 6214 15160 6245 15176
rect 6271 15160 6327 15216
rect 6353 15160 6409 15216
rect 6435 15160 6491 15216
rect 6517 15160 6573 15216
rect 6599 15160 6655 15216
rect 6681 15193 6702 15216
rect 6702 15193 6737 15216
rect 6763 15193 6768 15216
rect 6768 15193 6819 15216
rect 6681 15176 6737 15193
rect 6763 15176 6819 15193
rect 6681 15160 6702 15176
rect 6702 15160 6737 15176
rect 6763 15160 6768 15176
rect 6768 15160 6819 15176
rect 6845 15160 6901 15216
rect 6927 15160 6983 15216
rect 7009 15160 7065 15216
rect 7091 15160 7147 15216
rect 7173 15160 7229 15216
rect 7255 15193 7256 15216
rect 7256 15193 7308 15216
rect 7308 15193 7311 15216
rect 7337 15193 7374 15216
rect 7374 15193 7393 15216
rect 7255 15176 7311 15193
rect 7337 15176 7393 15193
rect 7255 15160 7256 15176
rect 7256 15160 7308 15176
rect 7308 15160 7311 15176
rect 7337 15160 7374 15176
rect 7374 15160 7393 15176
rect 7419 15160 7475 15216
rect 7501 15160 7557 15216
rect 7583 15160 7639 15216
rect 7665 15160 7721 15216
rect 7747 15160 7803 15216
rect 7829 15193 7862 15216
rect 7862 15193 7876 15216
rect 7876 15193 7885 15216
rect 7911 15193 7928 15216
rect 7928 15193 7967 15216
rect 7829 15176 7885 15193
rect 7911 15176 7967 15193
rect 7829 15160 7862 15176
rect 7862 15160 7876 15176
rect 7876 15160 7885 15176
rect 7911 15160 7928 15176
rect 7928 15160 7967 15176
rect 7993 15197 8047 15216
rect 8047 15197 8049 15216
rect 8075 15197 8099 15216
rect 8099 15197 8131 15216
rect 7993 15180 8049 15197
rect 8075 15180 8131 15197
rect 7993 15160 8047 15180
rect 8047 15160 8049 15180
rect 8075 15160 8099 15180
rect 8099 15160 8131 15180
rect 8157 15197 8169 15216
rect 8169 15197 8213 15216
rect 8157 15180 8213 15197
rect 8157 15160 8169 15180
rect 8169 15160 8213 15180
rect 5613 15124 5646 15136
rect 5646 15124 5660 15136
rect 5660 15124 5669 15136
rect 5696 15124 5712 15136
rect 5712 15124 5752 15136
rect 5613 15107 5669 15124
rect 5696 15107 5752 15124
rect 5613 15080 5646 15107
rect 5646 15080 5660 15107
rect 5660 15080 5669 15107
rect 5696 15080 5712 15107
rect 5712 15080 5752 15107
rect 5779 15080 5835 15136
rect 5861 15080 5917 15136
rect 5943 15080 5999 15136
rect 6025 15080 6081 15136
rect 6107 15124 6148 15136
rect 6148 15124 6163 15136
rect 6189 15124 6200 15136
rect 6200 15124 6214 15136
rect 6214 15124 6245 15136
rect 6107 15107 6163 15124
rect 6189 15107 6245 15124
rect 6107 15080 6148 15107
rect 6148 15080 6163 15107
rect 6189 15080 6200 15107
rect 6200 15080 6214 15107
rect 6214 15080 6245 15107
rect 6271 15080 6327 15136
rect 6353 15080 6409 15136
rect 6435 15080 6491 15136
rect 6517 15080 6573 15136
rect 6599 15080 6655 15136
rect 6681 15124 6702 15136
rect 6702 15124 6737 15136
rect 6763 15124 6768 15136
rect 6768 15124 6819 15136
rect 6681 15107 6737 15124
rect 6763 15107 6819 15124
rect 6681 15080 6702 15107
rect 6702 15080 6737 15107
rect 6763 15080 6768 15107
rect 6768 15080 6819 15107
rect 6845 15080 6901 15136
rect 6927 15080 6983 15136
rect 7009 15080 7065 15136
rect 7091 15080 7147 15136
rect 7173 15080 7229 15136
rect 7255 15124 7256 15136
rect 7256 15124 7308 15136
rect 7308 15124 7311 15136
rect 7337 15124 7374 15136
rect 7374 15124 7393 15136
rect 7255 15107 7311 15124
rect 7337 15107 7393 15124
rect 7255 15080 7256 15107
rect 7256 15080 7308 15107
rect 7308 15080 7311 15107
rect 7337 15080 7374 15107
rect 7374 15080 7393 15107
rect 7419 15080 7475 15136
rect 7501 15080 7557 15136
rect 7583 15080 7639 15136
rect 7665 15080 7721 15136
rect 7747 15080 7803 15136
rect 7829 15124 7862 15136
rect 7862 15124 7876 15136
rect 7876 15124 7885 15136
rect 7911 15124 7928 15136
rect 7928 15124 7967 15136
rect 7829 15107 7885 15124
rect 7911 15107 7967 15124
rect 7829 15080 7862 15107
rect 7862 15080 7876 15107
rect 7876 15080 7885 15107
rect 7911 15080 7928 15107
rect 7928 15080 7967 15107
rect 7993 15128 8047 15136
rect 8047 15128 8049 15136
rect 8075 15128 8099 15136
rect 8099 15128 8131 15136
rect 7993 15110 8049 15128
rect 8075 15110 8131 15128
rect 7993 15080 8047 15110
rect 8047 15080 8049 15110
rect 8075 15080 8099 15110
rect 8099 15080 8131 15110
rect 8157 15128 8169 15136
rect 8169 15128 8213 15136
rect 8157 15110 8213 15128
rect 8157 15080 8169 15110
rect 8169 15080 8213 15110
rect 5613 15055 5646 15056
rect 5646 15055 5660 15056
rect 5660 15055 5669 15056
rect 5696 15055 5712 15056
rect 5712 15055 5752 15056
rect 5613 15038 5669 15055
rect 5696 15038 5752 15055
rect 5613 15000 5646 15038
rect 5646 15000 5660 15038
rect 5660 15000 5669 15038
rect 5696 15000 5712 15038
rect 5712 15000 5752 15038
rect 5779 15000 5835 15056
rect 5861 15000 5917 15056
rect 5943 15000 5999 15056
rect 6025 15000 6081 15056
rect 6107 15055 6148 15056
rect 6148 15055 6163 15056
rect 6189 15055 6200 15056
rect 6200 15055 6214 15056
rect 6214 15055 6245 15056
rect 6107 15038 6163 15055
rect 6189 15038 6245 15055
rect 6107 15000 6148 15038
rect 6148 15000 6163 15038
rect 6189 15000 6200 15038
rect 6200 15000 6214 15038
rect 6214 15000 6245 15038
rect 6271 15000 6327 15056
rect 6353 15000 6409 15056
rect 6435 15000 6491 15056
rect 6517 15000 6573 15056
rect 6599 15000 6655 15056
rect 6681 15055 6702 15056
rect 6702 15055 6737 15056
rect 6763 15055 6768 15056
rect 6768 15055 6819 15056
rect 6681 15038 6737 15055
rect 6763 15038 6819 15055
rect 6681 15000 6702 15038
rect 6702 15000 6737 15038
rect 6763 15000 6768 15038
rect 6768 15000 6819 15038
rect 6845 15000 6901 15056
rect 6927 15000 6983 15056
rect 7009 15000 7065 15056
rect 7091 15000 7147 15056
rect 7173 15000 7229 15056
rect 7255 15055 7256 15056
rect 7256 15055 7308 15056
rect 7308 15055 7311 15056
rect 7337 15055 7374 15056
rect 7374 15055 7393 15056
rect 7255 15038 7311 15055
rect 7337 15038 7393 15055
rect 7255 15000 7256 15038
rect 7256 15000 7308 15038
rect 7308 15000 7311 15038
rect 7337 15000 7374 15038
rect 7374 15000 7393 15038
rect 7419 15000 7475 15056
rect 7501 15000 7557 15056
rect 7583 15000 7639 15056
rect 7665 15000 7721 15056
rect 7747 15000 7803 15056
rect 7829 15055 7862 15056
rect 7862 15055 7876 15056
rect 7876 15055 7885 15056
rect 7911 15055 7928 15056
rect 7928 15055 7967 15056
rect 7829 15038 7885 15055
rect 7911 15038 7967 15055
rect 7829 15000 7862 15038
rect 7862 15000 7876 15038
rect 7876 15000 7885 15038
rect 7911 15000 7928 15038
rect 7928 15000 7967 15038
rect 7993 15040 8049 15056
rect 8075 15040 8131 15056
rect 7993 15000 8047 15040
rect 8047 15000 8049 15040
rect 8075 15000 8099 15040
rect 8099 15000 8131 15040
rect 8157 15040 8213 15056
rect 8157 15000 8169 15040
rect 8169 15000 8213 15040
rect 5613 14968 5669 14976
rect 5696 14968 5752 14976
rect 5613 14920 5646 14968
rect 5646 14920 5660 14968
rect 5660 14920 5669 14968
rect 5696 14920 5712 14968
rect 5712 14920 5752 14968
rect 5779 14920 5835 14976
rect 5861 14920 5917 14976
rect 5943 14920 5999 14976
rect 6025 14920 6081 14976
rect 6107 14968 6163 14976
rect 6189 14968 6245 14976
rect 6107 14920 6148 14968
rect 6148 14920 6163 14968
rect 6189 14920 6200 14968
rect 6200 14920 6214 14968
rect 6214 14920 6245 14968
rect 6271 14920 6327 14976
rect 6353 14920 6409 14976
rect 6435 14920 6491 14976
rect 6517 14920 6573 14976
rect 6599 14920 6655 14976
rect 6681 14968 6737 14976
rect 6763 14968 6819 14976
rect 6681 14920 6702 14968
rect 6702 14920 6737 14968
rect 6763 14920 6768 14968
rect 6768 14920 6819 14968
rect 6845 14920 6901 14976
rect 6927 14920 6983 14976
rect 7009 14920 7065 14976
rect 7091 14920 7147 14976
rect 7173 14920 7229 14976
rect 7255 14968 7311 14976
rect 7337 14968 7393 14976
rect 7255 14920 7256 14968
rect 7256 14920 7308 14968
rect 7308 14920 7311 14968
rect 7337 14920 7374 14968
rect 7374 14920 7393 14968
rect 7419 14920 7475 14976
rect 7501 14920 7557 14976
rect 7583 14920 7639 14976
rect 7665 14920 7721 14976
rect 7747 14920 7803 14976
rect 7829 14968 7885 14976
rect 7911 14968 7967 14976
rect 7829 14920 7862 14968
rect 7862 14920 7876 14968
rect 7876 14920 7885 14968
rect 7911 14920 7928 14968
rect 7928 14920 7967 14968
rect 7993 14970 8049 14976
rect 8075 14970 8131 14976
rect 7993 14920 8047 14970
rect 8047 14920 8049 14970
rect 8075 14920 8099 14970
rect 8099 14920 8131 14970
rect 8157 14970 8213 14976
rect 8157 14920 8169 14970
rect 8169 14920 8213 14970
rect 5613 14846 5646 14896
rect 5646 14846 5660 14896
rect 5660 14846 5669 14896
rect 5696 14846 5712 14896
rect 5712 14846 5752 14896
rect 5613 14840 5669 14846
rect 5696 14840 5752 14846
rect 5779 14840 5835 14896
rect 5861 14840 5917 14896
rect 5943 14840 5999 14896
rect 6025 14840 6081 14896
rect 6107 14846 6148 14896
rect 6148 14846 6163 14896
rect 6189 14846 6200 14896
rect 6200 14846 6214 14896
rect 6214 14846 6245 14896
rect 6107 14840 6163 14846
rect 6189 14840 6245 14846
rect 6271 14840 6327 14896
rect 6353 14840 6409 14896
rect 6435 14840 6491 14896
rect 6517 14840 6573 14896
rect 6599 14840 6655 14896
rect 6681 14846 6702 14896
rect 6702 14846 6737 14896
rect 6763 14846 6768 14896
rect 6768 14846 6819 14896
rect 6681 14840 6737 14846
rect 6763 14840 6819 14846
rect 6845 14840 6901 14896
rect 6927 14840 6983 14896
rect 7009 14840 7065 14896
rect 7091 14840 7147 14896
rect 7173 14840 7229 14896
rect 7255 14846 7256 14896
rect 7256 14846 7308 14896
rect 7308 14846 7311 14896
rect 7337 14846 7374 14896
rect 7374 14846 7393 14896
rect 7255 14840 7311 14846
rect 7337 14840 7393 14846
rect 7419 14840 7475 14896
rect 7501 14840 7557 14896
rect 7583 14840 7639 14896
rect 7665 14840 7721 14896
rect 7747 14840 7803 14896
rect 7829 14846 7862 14896
rect 7862 14846 7876 14896
rect 7876 14846 7885 14896
rect 7911 14846 7928 14896
rect 7928 14846 7967 14896
rect 7829 14840 7885 14846
rect 7911 14840 7967 14846
rect 7993 14848 8047 14896
rect 8047 14848 8049 14896
rect 8075 14848 8099 14896
rect 8099 14848 8131 14896
rect 7993 14840 8049 14848
rect 8075 14840 8131 14848
rect 8157 14848 8169 14896
rect 8169 14848 8213 14896
rect 8157 14840 8213 14848
rect 2733 14663 2789 14719
rect 2814 14663 2870 14719
rect 2895 14663 2951 14719
rect 2976 14663 3032 14719
rect 3057 14714 3113 14719
rect 3138 14714 3194 14719
rect 3057 14663 3101 14714
rect 3101 14663 3113 14714
rect 3138 14663 3153 14714
rect 3153 14663 3167 14714
rect 3167 14663 3194 14714
rect 3219 14663 3275 14719
rect 3300 14663 3356 14719
rect 3381 14663 3437 14719
rect 3462 14663 3518 14719
rect 3543 14663 3599 14719
rect 3624 14714 3680 14719
rect 3705 14714 3761 14719
rect 3624 14663 3655 14714
rect 3655 14663 3680 14714
rect 3705 14663 3707 14714
rect 3707 14663 3721 14714
rect 3721 14663 3761 14714
rect 3786 14663 3842 14719
rect 3867 14663 3923 14719
rect 3948 14663 4004 14719
rect 4029 14663 4085 14719
rect 4110 14663 4166 14719
rect 4191 14714 4247 14719
rect 4272 14714 4328 14719
rect 4191 14663 4209 14714
rect 4209 14663 4247 14714
rect 4272 14663 4275 14714
rect 4275 14663 4327 14714
rect 4327 14663 4328 14714
rect 4353 14663 4409 14719
rect 4434 14663 4490 14719
rect 4515 14663 4571 14719
rect 4596 14663 4652 14719
rect 4677 14663 4733 14719
rect 4758 14714 4814 14719
rect 4839 14714 4895 14719
rect 4758 14663 4763 14714
rect 4763 14663 4814 14714
rect 4839 14663 4881 14714
rect 4881 14663 4895 14714
rect 4920 14663 4976 14719
rect 5001 14663 5057 14719
rect 5082 14663 5138 14719
rect 2733 14583 2789 14639
rect 2814 14583 2870 14639
rect 2895 14583 2951 14639
rect 2976 14583 3032 14639
rect 3057 14593 3101 14639
rect 3101 14593 3113 14639
rect 3138 14593 3153 14639
rect 3153 14593 3167 14639
rect 3167 14593 3194 14639
rect 3057 14583 3113 14593
rect 3138 14583 3194 14593
rect 3219 14583 3275 14639
rect 3300 14583 3356 14639
rect 3381 14583 3437 14639
rect 3462 14583 3518 14639
rect 3543 14583 3599 14639
rect 3624 14593 3655 14639
rect 3655 14593 3680 14639
rect 3705 14593 3707 14639
rect 3707 14593 3721 14639
rect 3721 14593 3761 14639
rect 3624 14583 3680 14593
rect 3705 14583 3761 14593
rect 3786 14583 3842 14639
rect 3867 14583 3923 14639
rect 3948 14583 4004 14639
rect 4029 14583 4085 14639
rect 4110 14583 4166 14639
rect 4191 14593 4209 14639
rect 4209 14593 4247 14639
rect 4272 14593 4275 14639
rect 4275 14593 4327 14639
rect 4327 14593 4328 14639
rect 4191 14583 4247 14593
rect 4272 14583 4328 14593
rect 4353 14583 4409 14639
rect 4434 14583 4490 14639
rect 4515 14583 4571 14639
rect 4596 14583 4652 14639
rect 4677 14583 4733 14639
rect 4758 14593 4763 14639
rect 4763 14593 4814 14639
rect 4839 14593 4881 14639
rect 4881 14593 4895 14639
rect 4758 14583 4814 14593
rect 4839 14583 4895 14593
rect 4920 14583 4976 14639
rect 5001 14583 5057 14639
rect 5082 14583 5138 14639
rect 2733 14503 2789 14559
rect 2814 14503 2870 14559
rect 2895 14503 2951 14559
rect 2976 14503 3032 14559
rect 3057 14524 3101 14559
rect 3101 14524 3113 14559
rect 3138 14524 3153 14559
rect 3153 14524 3167 14559
rect 3167 14524 3194 14559
rect 3057 14507 3113 14524
rect 3138 14507 3194 14524
rect 3057 14503 3101 14507
rect 3101 14503 3113 14507
rect 3138 14503 3153 14507
rect 3153 14503 3167 14507
rect 3167 14503 3194 14507
rect 3219 14503 3275 14559
rect 3300 14503 3356 14559
rect 3381 14503 3437 14559
rect 3462 14503 3518 14559
rect 3543 14503 3599 14559
rect 3624 14524 3655 14559
rect 3655 14524 3680 14559
rect 3705 14524 3707 14559
rect 3707 14524 3721 14559
rect 3721 14524 3761 14559
rect 3624 14507 3680 14524
rect 3705 14507 3761 14524
rect 3624 14503 3655 14507
rect 3655 14503 3680 14507
rect 3705 14503 3707 14507
rect 3707 14503 3721 14507
rect 3721 14503 3761 14507
rect 3786 14503 3842 14559
rect 3867 14503 3923 14559
rect 3948 14503 4004 14559
rect 4029 14503 4085 14559
rect 4110 14503 4166 14559
rect 4191 14524 4209 14559
rect 4209 14524 4247 14559
rect 4272 14524 4275 14559
rect 4275 14524 4327 14559
rect 4327 14524 4328 14559
rect 4191 14507 4247 14524
rect 4272 14507 4328 14524
rect 4191 14503 4209 14507
rect 4209 14503 4247 14507
rect 4272 14503 4275 14507
rect 4275 14503 4327 14507
rect 4327 14503 4328 14507
rect 4353 14503 4409 14559
rect 4434 14503 4490 14559
rect 4515 14503 4571 14559
rect 4596 14503 4652 14559
rect 4677 14503 4733 14559
rect 4758 14524 4763 14559
rect 4763 14524 4814 14559
rect 4839 14524 4881 14559
rect 4881 14524 4895 14559
rect 4758 14507 4814 14524
rect 4839 14507 4895 14524
rect 4758 14503 4763 14507
rect 4763 14503 4814 14507
rect 2733 14423 2789 14479
rect 2814 14423 2870 14479
rect 2895 14423 2951 14479
rect 2976 14423 3032 14479
rect 3057 14455 3101 14479
rect 3101 14455 3113 14479
rect 3138 14455 3153 14479
rect 3153 14455 3167 14479
rect 3167 14455 3194 14479
rect 3057 14438 3113 14455
rect 3138 14438 3194 14455
rect 3057 14423 3101 14438
rect 3101 14423 3113 14438
rect 3138 14423 3153 14438
rect 3153 14423 3167 14438
rect 3167 14423 3194 14438
rect 3219 14423 3275 14479
rect 3300 14423 3356 14479
rect 3381 14423 3437 14479
rect 3462 14423 3518 14479
rect 3543 14423 3599 14479
rect 3624 14455 3655 14479
rect 3655 14455 3680 14479
rect 3705 14455 3707 14479
rect 3707 14455 3721 14479
rect 3721 14455 3761 14479
rect 3624 14438 3680 14455
rect 3705 14438 3761 14455
rect 3624 14423 3655 14438
rect 3655 14423 3680 14438
rect 3705 14423 3707 14438
rect 3707 14423 3721 14438
rect 3721 14423 3761 14438
rect 3786 14423 3842 14479
rect 3867 14423 3923 14479
rect 3948 14423 4004 14479
rect 4029 14423 4085 14479
rect 4110 14423 4166 14479
rect 4191 14455 4209 14479
rect 4209 14455 4247 14479
rect 4272 14455 4275 14479
rect 4275 14455 4327 14479
rect 4327 14455 4328 14479
rect 4191 14438 4247 14455
rect 4272 14438 4328 14455
rect 4191 14423 4209 14438
rect 4209 14423 4247 14438
rect 4272 14423 4275 14438
rect 4275 14423 4327 14438
rect 4327 14423 4328 14438
rect 4353 14423 4409 14479
rect 4434 14423 4490 14479
rect 4515 14423 4571 14479
rect 4596 14423 4652 14479
rect 4677 14423 4733 14479
rect 4758 14455 4763 14479
rect 4763 14455 4814 14479
rect 4839 14503 4881 14507
rect 4881 14503 4895 14507
rect 4920 14503 4976 14559
rect 5001 14503 5057 14559
rect 5082 14503 5138 14559
rect 4839 14455 4881 14479
rect 4881 14455 4895 14479
rect 4758 14438 4814 14455
rect 4839 14438 4895 14455
rect 4758 14423 4763 14438
rect 4763 14423 4814 14438
rect 2733 14343 2789 14399
rect 2814 14343 2870 14399
rect 2895 14343 2951 14399
rect 2976 14343 3032 14399
rect 3057 14386 3101 14399
rect 3101 14386 3113 14399
rect 3138 14386 3153 14399
rect 3153 14386 3167 14399
rect 3167 14386 3194 14399
rect 3057 14368 3113 14386
rect 3138 14368 3194 14386
rect 3057 14343 3101 14368
rect 3101 14343 3113 14368
rect 3138 14343 3153 14368
rect 3153 14343 3167 14368
rect 3167 14343 3194 14368
rect 3219 14343 3275 14399
rect 3300 14343 3356 14399
rect 3381 14343 3437 14399
rect 3462 14343 3518 14399
rect 3543 14343 3599 14399
rect 3624 14386 3655 14399
rect 3655 14386 3680 14399
rect 3705 14386 3707 14399
rect 3707 14386 3721 14399
rect 3721 14386 3761 14399
rect 3624 14368 3680 14386
rect 3705 14368 3761 14386
rect 3624 14343 3655 14368
rect 3655 14343 3680 14368
rect 3705 14343 3707 14368
rect 3707 14343 3721 14368
rect 3721 14343 3761 14368
rect 3786 14343 3842 14399
rect 3867 14343 3923 14399
rect 3948 14343 4004 14399
rect 4029 14343 4085 14399
rect 4110 14343 4166 14399
rect 4191 14386 4209 14399
rect 4209 14386 4247 14399
rect 4272 14386 4275 14399
rect 4275 14386 4327 14399
rect 4327 14386 4328 14399
rect 4191 14368 4247 14386
rect 4272 14368 4328 14386
rect 4191 14343 4209 14368
rect 4209 14343 4247 14368
rect 4272 14343 4275 14368
rect 4275 14343 4327 14368
rect 4327 14343 4328 14368
rect 4353 14343 4409 14399
rect 4434 14343 4490 14399
rect 4515 14343 4571 14399
rect 4596 14343 4652 14399
rect 4677 14343 4733 14399
rect 4758 14386 4763 14399
rect 4763 14386 4814 14399
rect 4839 14423 4881 14438
rect 4881 14423 4895 14438
rect 4920 14423 4976 14479
rect 5001 14423 5057 14479
rect 5082 14423 5138 14479
rect 4839 14386 4881 14399
rect 4881 14386 4895 14399
rect 4758 14368 4814 14386
rect 4839 14368 4895 14386
rect 4758 14343 4763 14368
rect 4763 14343 4814 14368
rect 2733 14263 2789 14319
rect 2814 14263 2870 14319
rect 2895 14263 2951 14319
rect 2976 14263 3032 14319
rect 3057 14316 3101 14319
rect 3101 14316 3113 14319
rect 3138 14316 3153 14319
rect 3153 14316 3167 14319
rect 3167 14316 3194 14319
rect 3057 14298 3113 14316
rect 3138 14298 3194 14316
rect 3057 14263 3101 14298
rect 3101 14263 3113 14298
rect 3138 14263 3153 14298
rect 3153 14263 3167 14298
rect 3167 14263 3194 14298
rect 3219 14263 3275 14319
rect 3300 14263 3356 14319
rect 3381 14263 3437 14319
rect 3462 14263 3518 14319
rect 3543 14263 3599 14319
rect 3624 14316 3655 14319
rect 3655 14316 3680 14319
rect 3705 14316 3707 14319
rect 3707 14316 3721 14319
rect 3721 14316 3761 14319
rect 3624 14298 3680 14316
rect 3705 14298 3761 14316
rect 3624 14263 3655 14298
rect 3655 14263 3680 14298
rect 3705 14263 3707 14298
rect 3707 14263 3721 14298
rect 3721 14263 3761 14298
rect 3786 14263 3842 14319
rect 3867 14263 3923 14319
rect 3948 14263 4004 14319
rect 4029 14263 4085 14319
rect 4110 14263 4166 14319
rect 4191 14316 4209 14319
rect 4209 14316 4247 14319
rect 4272 14316 4275 14319
rect 4275 14316 4327 14319
rect 4327 14316 4328 14319
rect 4191 14298 4247 14316
rect 4272 14298 4328 14316
rect 4191 14263 4209 14298
rect 4209 14263 4247 14298
rect 4272 14263 4275 14298
rect 4275 14263 4327 14298
rect 4327 14263 4328 14298
rect 4353 14263 4409 14319
rect 4434 14263 4490 14319
rect 4515 14263 4571 14319
rect 4596 14263 4652 14319
rect 4677 14263 4733 14319
rect 4758 14316 4763 14319
rect 4763 14316 4814 14319
rect 4839 14343 4881 14368
rect 4881 14343 4895 14368
rect 4920 14343 4976 14399
rect 5001 14343 5057 14399
rect 5082 14343 5138 14399
rect 4839 14316 4881 14319
rect 4881 14316 4895 14319
rect 4758 14298 4814 14316
rect 4839 14298 4895 14316
rect 4758 14263 4763 14298
rect 4763 14263 4814 14298
rect 4839 14263 4881 14298
rect 4881 14263 4895 14298
rect 4920 14263 4976 14319
rect 5001 14263 5057 14319
rect 5082 14263 5138 14319
rect 2733 14183 2789 14239
rect 2814 14183 2870 14239
rect 2895 14183 2951 14239
rect 2976 14183 3032 14239
rect 3057 14228 3113 14239
rect 3138 14228 3194 14239
rect 3057 14183 3101 14228
rect 3101 14183 3113 14228
rect 3138 14183 3153 14228
rect 3153 14183 3167 14228
rect 3167 14183 3194 14228
rect 3219 14183 3275 14239
rect 3300 14183 3356 14239
rect 3381 14183 3437 14239
rect 3462 14183 3518 14239
rect 3543 14183 3599 14239
rect 3624 14228 3680 14239
rect 3705 14228 3761 14239
rect 3624 14183 3655 14228
rect 3655 14183 3680 14228
rect 3705 14183 3707 14228
rect 3707 14183 3721 14228
rect 3721 14183 3761 14228
rect 3786 14183 3842 14239
rect 3867 14183 3923 14239
rect 3948 14183 4004 14239
rect 4029 14183 4085 14239
rect 4110 14183 4166 14239
rect 4191 14228 4247 14239
rect 4272 14228 4328 14239
rect 4191 14183 4209 14228
rect 4209 14183 4247 14228
rect 4272 14183 4275 14228
rect 4275 14183 4327 14228
rect 4327 14183 4328 14228
rect 4353 14183 4409 14239
rect 4434 14183 4490 14239
rect 4515 14183 4571 14239
rect 4596 14183 4652 14239
rect 4677 14183 4733 14239
rect 4758 14228 4814 14239
rect 4839 14228 4895 14239
rect 4758 14183 4763 14228
rect 4763 14183 4814 14228
rect 4839 14183 4881 14228
rect 4881 14183 4895 14228
rect 4920 14183 4976 14239
rect 5001 14183 5057 14239
rect 5082 14183 5138 14239
rect 2733 14103 2789 14159
rect 2814 14103 2870 14159
rect 2895 14103 2951 14159
rect 2976 14103 3032 14159
rect 3057 14158 3113 14159
rect 3138 14158 3194 14159
rect 3057 14106 3101 14158
rect 3101 14106 3113 14158
rect 3138 14106 3153 14158
rect 3153 14106 3167 14158
rect 3167 14106 3194 14158
rect 3057 14103 3113 14106
rect 3138 14103 3194 14106
rect 3219 14103 3275 14159
rect 3300 14103 3356 14159
rect 3381 14103 3437 14159
rect 3462 14103 3518 14159
rect 3543 14103 3599 14159
rect 3624 14158 3680 14159
rect 3705 14158 3761 14159
rect 3624 14106 3655 14158
rect 3655 14106 3680 14158
rect 3705 14106 3707 14158
rect 3707 14106 3721 14158
rect 3721 14106 3761 14158
rect 3624 14103 3680 14106
rect 3705 14103 3761 14106
rect 3786 14103 3842 14159
rect 3867 14103 3923 14159
rect 3948 14103 4004 14159
rect 4029 14103 4085 14159
rect 4110 14103 4166 14159
rect 4191 14158 4247 14159
rect 4272 14158 4328 14159
rect 4191 14106 4209 14158
rect 4209 14106 4247 14158
rect 4272 14106 4275 14158
rect 4275 14106 4327 14158
rect 4327 14106 4328 14158
rect 4191 14103 4247 14106
rect 4272 14103 4328 14106
rect 4353 14103 4409 14159
rect 4434 14103 4490 14159
rect 4515 14103 4571 14159
rect 4596 14103 4652 14159
rect 4677 14103 4733 14159
rect 4758 14158 4814 14159
rect 4839 14158 4895 14159
rect 4758 14106 4763 14158
rect 4763 14106 4814 14158
rect 4839 14106 4881 14158
rect 4881 14106 4895 14158
rect 4758 14103 4814 14106
rect 4839 14103 4895 14106
rect 4920 14103 4976 14159
rect 5001 14103 5057 14159
rect 5082 14103 5138 14159
rect 5163 14103 5299 14719
rect 5613 13452 5669 13456
rect 5696 13452 5752 13456
rect 5613 13400 5646 13452
rect 5646 13400 5660 13452
rect 5660 13400 5669 13452
rect 5696 13400 5712 13452
rect 5712 13400 5752 13452
rect 5779 13400 5835 13456
rect 5861 13400 5917 13456
rect 5943 13400 5999 13456
rect 6025 13400 6081 13456
rect 6107 13452 6163 13456
rect 6189 13452 6245 13456
rect 6107 13400 6148 13452
rect 6148 13400 6163 13452
rect 6189 13400 6200 13452
rect 6200 13400 6214 13452
rect 6214 13400 6245 13452
rect 6271 13400 6327 13456
rect 6353 13400 6409 13456
rect 6435 13400 6491 13456
rect 6517 13400 6573 13456
rect 6599 13400 6655 13456
rect 6681 13452 6737 13456
rect 6763 13452 6819 13456
rect 6681 13400 6702 13452
rect 6702 13400 6737 13452
rect 6763 13400 6768 13452
rect 6768 13400 6819 13452
rect 6845 13400 6901 13456
rect 6927 13400 6983 13456
rect 7009 13400 7065 13456
rect 7091 13400 7147 13456
rect 7173 13400 7229 13456
rect 7255 13452 7311 13456
rect 7337 13452 7393 13456
rect 7255 13400 7256 13452
rect 7256 13400 7308 13452
rect 7308 13400 7311 13452
rect 7337 13400 7374 13452
rect 7374 13400 7393 13452
rect 7419 13400 7475 13456
rect 7501 13400 7557 13456
rect 7583 13400 7639 13456
rect 7665 13400 7721 13456
rect 7747 13400 7803 13456
rect 7829 13452 7885 13456
rect 7911 13452 7967 13456
rect 7829 13400 7862 13452
rect 7862 13400 7876 13452
rect 7876 13400 7885 13452
rect 7911 13400 7928 13452
rect 7928 13400 7967 13452
rect 7993 13404 8047 13456
rect 8047 13404 8049 13456
rect 8075 13404 8099 13456
rect 8099 13404 8131 13456
rect 7993 13400 8049 13404
rect 8075 13400 8131 13404
rect 8157 13404 8169 13456
rect 8169 13404 8213 13456
rect 8157 13400 8213 13404
rect 5613 13331 5646 13376
rect 5646 13331 5660 13376
rect 5660 13331 5669 13376
rect 5696 13331 5712 13376
rect 5712 13331 5752 13376
rect 5613 13320 5669 13331
rect 5696 13320 5752 13331
rect 5779 13320 5835 13376
rect 5861 13320 5917 13376
rect 5943 13320 5999 13376
rect 6025 13320 6081 13376
rect 6107 13331 6148 13376
rect 6148 13331 6163 13376
rect 6189 13331 6200 13376
rect 6200 13331 6214 13376
rect 6214 13331 6245 13376
rect 6107 13320 6163 13331
rect 6189 13320 6245 13331
rect 6271 13320 6327 13376
rect 6353 13320 6409 13376
rect 6435 13320 6491 13376
rect 6517 13320 6573 13376
rect 6599 13320 6655 13376
rect 6681 13331 6702 13376
rect 6702 13331 6737 13376
rect 6763 13331 6768 13376
rect 6768 13331 6819 13376
rect 6681 13320 6737 13331
rect 6763 13320 6819 13331
rect 6845 13320 6901 13376
rect 6927 13320 6983 13376
rect 7009 13320 7065 13376
rect 7091 13320 7147 13376
rect 7173 13320 7229 13376
rect 7255 13331 7256 13376
rect 7256 13331 7308 13376
rect 7308 13331 7311 13376
rect 7337 13331 7374 13376
rect 7374 13331 7393 13376
rect 7255 13320 7311 13331
rect 7337 13320 7393 13331
rect 7419 13320 7475 13376
rect 7501 13320 7557 13376
rect 7583 13320 7639 13376
rect 7665 13320 7721 13376
rect 7747 13320 7803 13376
rect 7829 13331 7862 13376
rect 7862 13331 7876 13376
rect 7876 13331 7885 13376
rect 7911 13331 7928 13376
rect 7928 13331 7967 13376
rect 7829 13320 7885 13331
rect 7911 13320 7967 13331
rect 7993 13335 8047 13376
rect 8047 13335 8049 13376
rect 8075 13335 8099 13376
rect 8099 13335 8131 13376
rect 7993 13320 8049 13335
rect 8075 13320 8131 13335
rect 8157 13335 8169 13376
rect 8169 13335 8213 13376
rect 8157 13320 8213 13335
rect 5613 13262 5646 13296
rect 5646 13262 5660 13296
rect 5660 13262 5669 13296
rect 5696 13262 5712 13296
rect 5712 13262 5752 13296
rect 5613 13245 5669 13262
rect 5696 13245 5752 13262
rect 5613 13240 5646 13245
rect 5646 13240 5660 13245
rect 5660 13240 5669 13245
rect 5696 13240 5712 13245
rect 5712 13240 5752 13245
rect 5779 13240 5835 13296
rect 5861 13240 5917 13296
rect 5943 13240 5999 13296
rect 6025 13240 6081 13296
rect 6107 13262 6148 13296
rect 6148 13262 6163 13296
rect 6189 13262 6200 13296
rect 6200 13262 6214 13296
rect 6214 13262 6245 13296
rect 6107 13245 6163 13262
rect 6189 13245 6245 13262
rect 6107 13240 6148 13245
rect 6148 13240 6163 13245
rect 6189 13240 6200 13245
rect 6200 13240 6214 13245
rect 6214 13240 6245 13245
rect 6271 13240 6327 13296
rect 6353 13240 6409 13296
rect 6435 13240 6491 13296
rect 6517 13240 6573 13296
rect 6599 13240 6655 13296
rect 6681 13262 6702 13296
rect 6702 13262 6737 13296
rect 6763 13262 6768 13296
rect 6768 13262 6819 13296
rect 6681 13245 6737 13262
rect 6763 13245 6819 13262
rect 6681 13240 6702 13245
rect 6702 13240 6737 13245
rect 6763 13240 6768 13245
rect 6768 13240 6819 13245
rect 6845 13240 6901 13296
rect 6927 13240 6983 13296
rect 7009 13240 7065 13296
rect 7091 13240 7147 13296
rect 7173 13240 7229 13296
rect 7255 13262 7256 13296
rect 7256 13262 7308 13296
rect 7308 13262 7311 13296
rect 7337 13262 7374 13296
rect 7374 13262 7393 13296
rect 7255 13245 7311 13262
rect 7337 13245 7393 13262
rect 7255 13240 7256 13245
rect 7256 13240 7308 13245
rect 7308 13240 7311 13245
rect 7337 13240 7374 13245
rect 7374 13240 7393 13245
rect 7419 13240 7475 13296
rect 7501 13240 7557 13296
rect 7583 13240 7639 13296
rect 7665 13240 7721 13296
rect 7747 13240 7803 13296
rect 7829 13262 7862 13296
rect 7862 13262 7876 13296
rect 7876 13262 7885 13296
rect 7911 13262 7928 13296
rect 7928 13262 7967 13296
rect 7829 13245 7885 13262
rect 7911 13245 7967 13262
rect 7829 13240 7862 13245
rect 7862 13240 7876 13245
rect 7876 13240 7885 13245
rect 7911 13240 7928 13245
rect 7928 13240 7967 13245
rect 7993 13266 8047 13296
rect 8047 13266 8049 13296
rect 8075 13266 8099 13296
rect 8099 13266 8131 13296
rect 7993 13249 8049 13266
rect 8075 13249 8131 13266
rect 7993 13240 8047 13249
rect 8047 13240 8049 13249
rect 8075 13240 8099 13249
rect 8099 13240 8131 13249
rect 8157 13266 8169 13296
rect 8169 13266 8213 13296
rect 8157 13249 8213 13266
rect 8157 13240 8169 13249
rect 8169 13240 8213 13249
rect 5613 13193 5646 13216
rect 5646 13193 5660 13216
rect 5660 13193 5669 13216
rect 5696 13193 5712 13216
rect 5712 13193 5752 13216
rect 5613 13176 5669 13193
rect 5696 13176 5752 13193
rect 5613 13160 5646 13176
rect 5646 13160 5660 13176
rect 5660 13160 5669 13176
rect 5696 13160 5712 13176
rect 5712 13160 5752 13176
rect 5779 13160 5835 13216
rect 5861 13160 5917 13216
rect 5943 13160 5999 13216
rect 6025 13160 6081 13216
rect 6107 13193 6148 13216
rect 6148 13193 6163 13216
rect 6189 13193 6200 13216
rect 6200 13193 6214 13216
rect 6214 13193 6245 13216
rect 6107 13176 6163 13193
rect 6189 13176 6245 13193
rect 6107 13160 6148 13176
rect 6148 13160 6163 13176
rect 6189 13160 6200 13176
rect 6200 13160 6214 13176
rect 6214 13160 6245 13176
rect 6271 13160 6327 13216
rect 6353 13160 6409 13216
rect 6435 13160 6491 13216
rect 6517 13160 6573 13216
rect 6599 13160 6655 13216
rect 6681 13193 6702 13216
rect 6702 13193 6737 13216
rect 6763 13193 6768 13216
rect 6768 13193 6819 13216
rect 6681 13176 6737 13193
rect 6763 13176 6819 13193
rect 6681 13160 6702 13176
rect 6702 13160 6737 13176
rect 6763 13160 6768 13176
rect 6768 13160 6819 13176
rect 6845 13160 6901 13216
rect 6927 13160 6983 13216
rect 7009 13160 7065 13216
rect 7091 13160 7147 13216
rect 7173 13160 7229 13216
rect 7255 13193 7256 13216
rect 7256 13193 7308 13216
rect 7308 13193 7311 13216
rect 7337 13193 7374 13216
rect 7374 13193 7393 13216
rect 7255 13176 7311 13193
rect 7337 13176 7393 13193
rect 7255 13160 7256 13176
rect 7256 13160 7308 13176
rect 7308 13160 7311 13176
rect 7337 13160 7374 13176
rect 7374 13160 7393 13176
rect 7419 13160 7475 13216
rect 7501 13160 7557 13216
rect 7583 13160 7639 13216
rect 7665 13160 7721 13216
rect 7747 13160 7803 13216
rect 7829 13193 7862 13216
rect 7862 13193 7876 13216
rect 7876 13193 7885 13216
rect 7911 13193 7928 13216
rect 7928 13193 7967 13216
rect 7829 13176 7885 13193
rect 7911 13176 7967 13193
rect 7829 13160 7862 13176
rect 7862 13160 7876 13176
rect 7876 13160 7885 13176
rect 7911 13160 7928 13176
rect 7928 13160 7967 13176
rect 7993 13197 8047 13216
rect 8047 13197 8049 13216
rect 8075 13197 8099 13216
rect 8099 13197 8131 13216
rect 7993 13180 8049 13197
rect 8075 13180 8131 13197
rect 7993 13160 8047 13180
rect 8047 13160 8049 13180
rect 8075 13160 8099 13180
rect 8099 13160 8131 13180
rect 8157 13197 8169 13216
rect 8169 13197 8213 13216
rect 8157 13180 8213 13197
rect 8157 13160 8169 13180
rect 8169 13160 8213 13180
rect 5613 13124 5646 13136
rect 5646 13124 5660 13136
rect 5660 13124 5669 13136
rect 5696 13124 5712 13136
rect 5712 13124 5752 13136
rect 5613 13107 5669 13124
rect 5696 13107 5752 13124
rect 5613 13080 5646 13107
rect 5646 13080 5660 13107
rect 5660 13080 5669 13107
rect 5696 13080 5712 13107
rect 5712 13080 5752 13107
rect 5779 13080 5835 13136
rect 5861 13080 5917 13136
rect 5943 13080 5999 13136
rect 6025 13080 6081 13136
rect 6107 13124 6148 13136
rect 6148 13124 6163 13136
rect 6189 13124 6200 13136
rect 6200 13124 6214 13136
rect 6214 13124 6245 13136
rect 6107 13107 6163 13124
rect 6189 13107 6245 13124
rect 6107 13080 6148 13107
rect 6148 13080 6163 13107
rect 6189 13080 6200 13107
rect 6200 13080 6214 13107
rect 6214 13080 6245 13107
rect 6271 13080 6327 13136
rect 6353 13080 6409 13136
rect 6435 13080 6491 13136
rect 6517 13080 6573 13136
rect 6599 13080 6655 13136
rect 6681 13124 6702 13136
rect 6702 13124 6737 13136
rect 6763 13124 6768 13136
rect 6768 13124 6819 13136
rect 6681 13107 6737 13124
rect 6763 13107 6819 13124
rect 6681 13080 6702 13107
rect 6702 13080 6737 13107
rect 6763 13080 6768 13107
rect 6768 13080 6819 13107
rect 6845 13080 6901 13136
rect 6927 13080 6983 13136
rect 7009 13080 7065 13136
rect 7091 13080 7147 13136
rect 7173 13080 7229 13136
rect 7255 13124 7256 13136
rect 7256 13124 7308 13136
rect 7308 13124 7311 13136
rect 7337 13124 7374 13136
rect 7374 13124 7393 13136
rect 7255 13107 7311 13124
rect 7337 13107 7393 13124
rect 7255 13080 7256 13107
rect 7256 13080 7308 13107
rect 7308 13080 7311 13107
rect 7337 13080 7374 13107
rect 7374 13080 7393 13107
rect 7419 13080 7475 13136
rect 7501 13080 7557 13136
rect 7583 13080 7639 13136
rect 7665 13080 7721 13136
rect 7747 13080 7803 13136
rect 7829 13124 7862 13136
rect 7862 13124 7876 13136
rect 7876 13124 7885 13136
rect 7911 13124 7928 13136
rect 7928 13124 7967 13136
rect 7829 13107 7885 13124
rect 7911 13107 7967 13124
rect 7829 13080 7862 13107
rect 7862 13080 7876 13107
rect 7876 13080 7885 13107
rect 7911 13080 7928 13107
rect 7928 13080 7967 13107
rect 7993 13128 8047 13136
rect 8047 13128 8049 13136
rect 8075 13128 8099 13136
rect 8099 13128 8131 13136
rect 7993 13110 8049 13128
rect 8075 13110 8131 13128
rect 7993 13080 8047 13110
rect 8047 13080 8049 13110
rect 8075 13080 8099 13110
rect 8099 13080 8131 13110
rect 8157 13128 8169 13136
rect 8169 13128 8213 13136
rect 8157 13110 8213 13128
rect 8157 13080 8169 13110
rect 8169 13080 8213 13110
rect 5613 13055 5646 13056
rect 5646 13055 5660 13056
rect 5660 13055 5669 13056
rect 5696 13055 5712 13056
rect 5712 13055 5752 13056
rect 5613 13038 5669 13055
rect 5696 13038 5752 13055
rect 5613 13000 5646 13038
rect 5646 13000 5660 13038
rect 5660 13000 5669 13038
rect 5696 13000 5712 13038
rect 5712 13000 5752 13038
rect 5779 13000 5835 13056
rect 5861 13000 5917 13056
rect 5943 13000 5999 13056
rect 6025 13000 6081 13056
rect 6107 13055 6148 13056
rect 6148 13055 6163 13056
rect 6189 13055 6200 13056
rect 6200 13055 6214 13056
rect 6214 13055 6245 13056
rect 6107 13038 6163 13055
rect 6189 13038 6245 13055
rect 6107 13000 6148 13038
rect 6148 13000 6163 13038
rect 6189 13000 6200 13038
rect 6200 13000 6214 13038
rect 6214 13000 6245 13038
rect 6271 13000 6327 13056
rect 6353 13000 6409 13056
rect 6435 13000 6491 13056
rect 6517 13000 6573 13056
rect 6599 13000 6655 13056
rect 6681 13055 6702 13056
rect 6702 13055 6737 13056
rect 6763 13055 6768 13056
rect 6768 13055 6819 13056
rect 6681 13038 6737 13055
rect 6763 13038 6819 13055
rect 6681 13000 6702 13038
rect 6702 13000 6737 13038
rect 6763 13000 6768 13038
rect 6768 13000 6819 13038
rect 6845 13000 6901 13056
rect 6927 13000 6983 13056
rect 7009 13000 7065 13056
rect 7091 13000 7147 13056
rect 7173 13000 7229 13056
rect 7255 13055 7256 13056
rect 7256 13055 7308 13056
rect 7308 13055 7311 13056
rect 7337 13055 7374 13056
rect 7374 13055 7393 13056
rect 7255 13038 7311 13055
rect 7337 13038 7393 13055
rect 7255 13000 7256 13038
rect 7256 13000 7308 13038
rect 7308 13000 7311 13038
rect 7337 13000 7374 13038
rect 7374 13000 7393 13038
rect 7419 13000 7475 13056
rect 7501 13000 7557 13056
rect 7583 13000 7639 13056
rect 7665 13000 7721 13056
rect 7747 13000 7803 13056
rect 7829 13055 7862 13056
rect 7862 13055 7876 13056
rect 7876 13055 7885 13056
rect 7911 13055 7928 13056
rect 7928 13055 7967 13056
rect 7829 13038 7885 13055
rect 7911 13038 7967 13055
rect 7829 13000 7862 13038
rect 7862 13000 7876 13038
rect 7876 13000 7885 13038
rect 7911 13000 7928 13038
rect 7928 13000 7967 13038
rect 7993 13040 8049 13056
rect 8075 13040 8131 13056
rect 7993 13000 8047 13040
rect 8047 13000 8049 13040
rect 8075 13000 8099 13040
rect 8099 13000 8131 13040
rect 8157 13040 8213 13056
rect 8157 13000 8169 13040
rect 8169 13000 8213 13040
rect 5613 12968 5669 12976
rect 5696 12968 5752 12976
rect 5613 12920 5646 12968
rect 5646 12920 5660 12968
rect 5660 12920 5669 12968
rect 5696 12920 5712 12968
rect 5712 12920 5752 12968
rect 5779 12920 5835 12976
rect 5861 12920 5917 12976
rect 5943 12920 5999 12976
rect 6025 12920 6081 12976
rect 6107 12968 6163 12976
rect 6189 12968 6245 12976
rect 6107 12920 6148 12968
rect 6148 12920 6163 12968
rect 6189 12920 6200 12968
rect 6200 12920 6214 12968
rect 6214 12920 6245 12968
rect 6271 12920 6327 12976
rect 6353 12920 6409 12976
rect 6435 12920 6491 12976
rect 6517 12920 6573 12976
rect 6599 12920 6655 12976
rect 6681 12968 6737 12976
rect 6763 12968 6819 12976
rect 6681 12920 6702 12968
rect 6702 12920 6737 12968
rect 6763 12920 6768 12968
rect 6768 12920 6819 12968
rect 6845 12920 6901 12976
rect 6927 12920 6983 12976
rect 7009 12920 7065 12976
rect 7091 12920 7147 12976
rect 7173 12920 7229 12976
rect 7255 12968 7311 12976
rect 7337 12968 7393 12976
rect 7255 12920 7256 12968
rect 7256 12920 7308 12968
rect 7308 12920 7311 12968
rect 7337 12920 7374 12968
rect 7374 12920 7393 12968
rect 7419 12920 7475 12976
rect 7501 12920 7557 12976
rect 7583 12920 7639 12976
rect 7665 12920 7721 12976
rect 7747 12920 7803 12976
rect 7829 12968 7885 12976
rect 7911 12968 7967 12976
rect 7829 12920 7862 12968
rect 7862 12920 7876 12968
rect 7876 12920 7885 12968
rect 7911 12920 7928 12968
rect 7928 12920 7967 12968
rect 7993 12970 8049 12976
rect 8075 12970 8131 12976
rect 7993 12920 8047 12970
rect 8047 12920 8049 12970
rect 8075 12920 8099 12970
rect 8099 12920 8131 12970
rect 8157 12970 8213 12976
rect 8157 12920 8169 12970
rect 8169 12920 8213 12970
rect 5613 12846 5646 12896
rect 5646 12846 5660 12896
rect 5660 12846 5669 12896
rect 5696 12846 5712 12896
rect 5712 12846 5752 12896
rect 5613 12840 5669 12846
rect 5696 12840 5752 12846
rect 5779 12840 5835 12896
rect 5861 12840 5917 12896
rect 5943 12840 5999 12896
rect 6025 12840 6081 12896
rect 6107 12846 6148 12896
rect 6148 12846 6163 12896
rect 6189 12846 6200 12896
rect 6200 12846 6214 12896
rect 6214 12846 6245 12896
rect 6107 12840 6163 12846
rect 6189 12840 6245 12846
rect 6271 12840 6327 12896
rect 6353 12840 6409 12896
rect 6435 12840 6491 12896
rect 6517 12840 6573 12896
rect 6599 12840 6655 12896
rect 6681 12846 6702 12896
rect 6702 12846 6737 12896
rect 6763 12846 6768 12896
rect 6768 12846 6819 12896
rect 6681 12840 6737 12846
rect 6763 12840 6819 12846
rect 6845 12840 6901 12896
rect 6927 12840 6983 12896
rect 7009 12840 7065 12896
rect 7091 12840 7147 12896
rect 7173 12840 7229 12896
rect 7255 12846 7256 12896
rect 7256 12846 7308 12896
rect 7308 12846 7311 12896
rect 7337 12846 7374 12896
rect 7374 12846 7393 12896
rect 7255 12840 7311 12846
rect 7337 12840 7393 12846
rect 7419 12840 7475 12896
rect 7501 12840 7557 12896
rect 7583 12840 7639 12896
rect 7665 12840 7721 12896
rect 7747 12840 7803 12896
rect 7829 12846 7862 12896
rect 7862 12846 7876 12896
rect 7876 12846 7885 12896
rect 7911 12846 7928 12896
rect 7928 12846 7967 12896
rect 7829 12840 7885 12846
rect 7911 12840 7967 12846
rect 7993 12848 8047 12896
rect 8047 12848 8049 12896
rect 8075 12848 8099 12896
rect 8099 12848 8131 12896
rect 7993 12840 8049 12848
rect 8075 12840 8131 12848
rect 8157 12848 8169 12896
rect 8169 12848 8213 12896
rect 8157 12840 8213 12848
rect 2733 12663 2789 12719
rect 2814 12663 2870 12719
rect 2895 12663 2951 12719
rect 2976 12663 3032 12719
rect 3057 12714 3113 12719
rect 3138 12714 3194 12719
rect 3057 12663 3101 12714
rect 3101 12663 3113 12714
rect 3138 12663 3153 12714
rect 3153 12663 3167 12714
rect 3167 12663 3194 12714
rect 3219 12663 3275 12719
rect 3300 12663 3356 12719
rect 3381 12663 3437 12719
rect 3462 12663 3518 12719
rect 3543 12663 3599 12719
rect 3624 12714 3680 12719
rect 3705 12714 3761 12719
rect 3624 12663 3655 12714
rect 3655 12663 3680 12714
rect 3705 12663 3707 12714
rect 3707 12663 3721 12714
rect 3721 12663 3761 12714
rect 3786 12663 3842 12719
rect 3867 12663 3923 12719
rect 3948 12663 4004 12719
rect 4029 12663 4085 12719
rect 4110 12663 4166 12719
rect 4191 12714 4247 12719
rect 4272 12714 4328 12719
rect 4191 12663 4209 12714
rect 4209 12663 4247 12714
rect 4272 12663 4275 12714
rect 4275 12663 4327 12714
rect 4327 12663 4328 12714
rect 4353 12663 4409 12719
rect 4434 12663 4490 12719
rect 4515 12663 4571 12719
rect 4596 12663 4652 12719
rect 4677 12663 4733 12719
rect 4758 12714 4814 12719
rect 4839 12714 4895 12719
rect 4758 12663 4763 12714
rect 4763 12663 4814 12714
rect 4839 12663 4881 12714
rect 4881 12663 4895 12714
rect 4920 12663 4976 12719
rect 5001 12663 5057 12719
rect 5082 12663 5138 12719
rect 2733 12583 2789 12639
rect 2814 12583 2870 12639
rect 2895 12583 2951 12639
rect 2976 12583 3032 12639
rect 3057 12593 3101 12639
rect 3101 12593 3113 12639
rect 3138 12593 3153 12639
rect 3153 12593 3167 12639
rect 3167 12593 3194 12639
rect 3057 12583 3113 12593
rect 3138 12583 3194 12593
rect 3219 12583 3275 12639
rect 3300 12583 3356 12639
rect 3381 12583 3437 12639
rect 3462 12583 3518 12639
rect 3543 12583 3599 12639
rect 3624 12593 3655 12639
rect 3655 12593 3680 12639
rect 3705 12593 3707 12639
rect 3707 12593 3721 12639
rect 3721 12593 3761 12639
rect 3624 12583 3680 12593
rect 3705 12583 3761 12593
rect 3786 12583 3842 12639
rect 3867 12583 3923 12639
rect 3948 12583 4004 12639
rect 4029 12583 4085 12639
rect 4110 12583 4166 12639
rect 4191 12593 4209 12639
rect 4209 12593 4247 12639
rect 4272 12593 4275 12639
rect 4275 12593 4327 12639
rect 4327 12593 4328 12639
rect 4191 12583 4247 12593
rect 4272 12583 4328 12593
rect 4353 12583 4409 12639
rect 4434 12583 4490 12639
rect 4515 12583 4571 12639
rect 4596 12583 4652 12639
rect 4677 12583 4733 12639
rect 4758 12593 4763 12639
rect 4763 12593 4814 12639
rect 4839 12593 4881 12639
rect 4881 12593 4895 12639
rect 4758 12583 4814 12593
rect 4839 12583 4895 12593
rect 4920 12583 4976 12639
rect 5001 12583 5057 12639
rect 5082 12583 5138 12639
rect 2733 12503 2789 12559
rect 2814 12503 2870 12559
rect 2895 12503 2951 12559
rect 2976 12503 3032 12559
rect 3057 12524 3101 12559
rect 3101 12524 3113 12559
rect 3138 12524 3153 12559
rect 3153 12524 3167 12559
rect 3167 12524 3194 12559
rect 3057 12507 3113 12524
rect 3138 12507 3194 12524
rect 3057 12503 3101 12507
rect 3101 12503 3113 12507
rect 3138 12503 3153 12507
rect 3153 12503 3167 12507
rect 3167 12503 3194 12507
rect 3219 12503 3275 12559
rect 3300 12503 3356 12559
rect 3381 12503 3437 12559
rect 3462 12503 3518 12559
rect 3543 12503 3599 12559
rect 3624 12524 3655 12559
rect 3655 12524 3680 12559
rect 3705 12524 3707 12559
rect 3707 12524 3721 12559
rect 3721 12524 3761 12559
rect 3624 12507 3680 12524
rect 3705 12507 3761 12524
rect 3624 12503 3655 12507
rect 3655 12503 3680 12507
rect 3705 12503 3707 12507
rect 3707 12503 3721 12507
rect 3721 12503 3761 12507
rect 3786 12503 3842 12559
rect 3867 12503 3923 12559
rect 3948 12503 4004 12559
rect 4029 12503 4085 12559
rect 4110 12503 4166 12559
rect 4191 12524 4209 12559
rect 4209 12524 4247 12559
rect 4272 12524 4275 12559
rect 4275 12524 4327 12559
rect 4327 12524 4328 12559
rect 4191 12507 4247 12524
rect 4272 12507 4328 12524
rect 4191 12503 4209 12507
rect 4209 12503 4247 12507
rect 4272 12503 4275 12507
rect 4275 12503 4327 12507
rect 4327 12503 4328 12507
rect 4353 12503 4409 12559
rect 4434 12503 4490 12559
rect 4515 12503 4571 12559
rect 4596 12503 4652 12559
rect 4677 12503 4733 12559
rect 4758 12524 4763 12559
rect 4763 12524 4814 12559
rect 4839 12524 4881 12559
rect 4881 12524 4895 12559
rect 4758 12507 4814 12524
rect 4839 12507 4895 12524
rect 4758 12503 4763 12507
rect 4763 12503 4814 12507
rect 2733 12423 2789 12479
rect 2814 12423 2870 12479
rect 2895 12423 2951 12479
rect 2976 12423 3032 12479
rect 3057 12455 3101 12479
rect 3101 12455 3113 12479
rect 3138 12455 3153 12479
rect 3153 12455 3167 12479
rect 3167 12455 3194 12479
rect 3057 12438 3113 12455
rect 3138 12438 3194 12455
rect 3057 12423 3101 12438
rect 3101 12423 3113 12438
rect 3138 12423 3153 12438
rect 3153 12423 3167 12438
rect 3167 12423 3194 12438
rect 3219 12423 3275 12479
rect 3300 12423 3356 12479
rect 3381 12423 3437 12479
rect 3462 12423 3518 12479
rect 3543 12423 3599 12479
rect 3624 12455 3655 12479
rect 3655 12455 3680 12479
rect 3705 12455 3707 12479
rect 3707 12455 3721 12479
rect 3721 12455 3761 12479
rect 3624 12438 3680 12455
rect 3705 12438 3761 12455
rect 3624 12423 3655 12438
rect 3655 12423 3680 12438
rect 3705 12423 3707 12438
rect 3707 12423 3721 12438
rect 3721 12423 3761 12438
rect 3786 12423 3842 12479
rect 3867 12423 3923 12479
rect 3948 12423 4004 12479
rect 4029 12423 4085 12479
rect 4110 12423 4166 12479
rect 4191 12455 4209 12479
rect 4209 12455 4247 12479
rect 4272 12455 4275 12479
rect 4275 12455 4327 12479
rect 4327 12455 4328 12479
rect 4191 12438 4247 12455
rect 4272 12438 4328 12455
rect 4191 12423 4209 12438
rect 4209 12423 4247 12438
rect 4272 12423 4275 12438
rect 4275 12423 4327 12438
rect 4327 12423 4328 12438
rect 4353 12423 4409 12479
rect 4434 12423 4490 12479
rect 4515 12423 4571 12479
rect 4596 12423 4652 12479
rect 4677 12423 4733 12479
rect 4758 12455 4763 12479
rect 4763 12455 4814 12479
rect 4839 12503 4881 12507
rect 4881 12503 4895 12507
rect 4920 12503 4976 12559
rect 5001 12503 5057 12559
rect 5082 12503 5138 12559
rect 4839 12455 4881 12479
rect 4881 12455 4895 12479
rect 4758 12438 4814 12455
rect 4839 12438 4895 12455
rect 4758 12423 4763 12438
rect 4763 12423 4814 12438
rect 2733 12343 2789 12399
rect 2814 12343 2870 12399
rect 2895 12343 2951 12399
rect 2976 12343 3032 12399
rect 3057 12386 3101 12399
rect 3101 12386 3113 12399
rect 3138 12386 3153 12399
rect 3153 12386 3167 12399
rect 3167 12386 3194 12399
rect 3057 12368 3113 12386
rect 3138 12368 3194 12386
rect 3057 12343 3101 12368
rect 3101 12343 3113 12368
rect 3138 12343 3153 12368
rect 3153 12343 3167 12368
rect 3167 12343 3194 12368
rect 3219 12343 3275 12399
rect 3300 12343 3356 12399
rect 3381 12343 3437 12399
rect 3462 12343 3518 12399
rect 3543 12343 3599 12399
rect 3624 12386 3655 12399
rect 3655 12386 3680 12399
rect 3705 12386 3707 12399
rect 3707 12386 3721 12399
rect 3721 12386 3761 12399
rect 3624 12368 3680 12386
rect 3705 12368 3761 12386
rect 3624 12343 3655 12368
rect 3655 12343 3680 12368
rect 3705 12343 3707 12368
rect 3707 12343 3721 12368
rect 3721 12343 3761 12368
rect 3786 12343 3842 12399
rect 3867 12343 3923 12399
rect 3948 12343 4004 12399
rect 4029 12343 4085 12399
rect 4110 12343 4166 12399
rect 4191 12386 4209 12399
rect 4209 12386 4247 12399
rect 4272 12386 4275 12399
rect 4275 12386 4327 12399
rect 4327 12386 4328 12399
rect 4191 12368 4247 12386
rect 4272 12368 4328 12386
rect 4191 12343 4209 12368
rect 4209 12343 4247 12368
rect 4272 12343 4275 12368
rect 4275 12343 4327 12368
rect 4327 12343 4328 12368
rect 4353 12343 4409 12399
rect 4434 12343 4490 12399
rect 4515 12343 4571 12399
rect 4596 12343 4652 12399
rect 4677 12343 4733 12399
rect 4758 12386 4763 12399
rect 4763 12386 4814 12399
rect 4839 12423 4881 12438
rect 4881 12423 4895 12438
rect 4920 12423 4976 12479
rect 5001 12423 5057 12479
rect 5082 12423 5138 12479
rect 4839 12386 4881 12399
rect 4881 12386 4895 12399
rect 4758 12368 4814 12386
rect 4839 12368 4895 12386
rect 4758 12343 4763 12368
rect 4763 12343 4814 12368
rect 2733 12263 2789 12319
rect 2814 12263 2870 12319
rect 2895 12263 2951 12319
rect 2976 12263 3032 12319
rect 3057 12316 3101 12319
rect 3101 12316 3113 12319
rect 3138 12316 3153 12319
rect 3153 12316 3167 12319
rect 3167 12316 3194 12319
rect 3057 12298 3113 12316
rect 3138 12298 3194 12316
rect 3057 12263 3101 12298
rect 3101 12263 3113 12298
rect 3138 12263 3153 12298
rect 3153 12263 3167 12298
rect 3167 12263 3194 12298
rect 3219 12263 3275 12319
rect 3300 12263 3356 12319
rect 3381 12263 3437 12319
rect 3462 12263 3518 12319
rect 3543 12263 3599 12319
rect 3624 12316 3655 12319
rect 3655 12316 3680 12319
rect 3705 12316 3707 12319
rect 3707 12316 3721 12319
rect 3721 12316 3761 12319
rect 3624 12298 3680 12316
rect 3705 12298 3761 12316
rect 3624 12263 3655 12298
rect 3655 12263 3680 12298
rect 3705 12263 3707 12298
rect 3707 12263 3721 12298
rect 3721 12263 3761 12298
rect 3786 12263 3842 12319
rect 3867 12263 3923 12319
rect 3948 12263 4004 12319
rect 4029 12263 4085 12319
rect 4110 12263 4166 12319
rect 4191 12316 4209 12319
rect 4209 12316 4247 12319
rect 4272 12316 4275 12319
rect 4275 12316 4327 12319
rect 4327 12316 4328 12319
rect 4191 12298 4247 12316
rect 4272 12298 4328 12316
rect 4191 12263 4209 12298
rect 4209 12263 4247 12298
rect 4272 12263 4275 12298
rect 4275 12263 4327 12298
rect 4327 12263 4328 12298
rect 4353 12263 4409 12319
rect 4434 12263 4490 12319
rect 4515 12263 4571 12319
rect 4596 12263 4652 12319
rect 4677 12263 4733 12319
rect 4758 12316 4763 12319
rect 4763 12316 4814 12319
rect 4839 12343 4881 12368
rect 4881 12343 4895 12368
rect 4920 12343 4976 12399
rect 5001 12343 5057 12399
rect 5082 12343 5138 12399
rect 4839 12316 4881 12319
rect 4881 12316 4895 12319
rect 4758 12298 4814 12316
rect 4839 12298 4895 12316
rect 4758 12263 4763 12298
rect 4763 12263 4814 12298
rect 4839 12263 4881 12298
rect 4881 12263 4895 12298
rect 4920 12263 4976 12319
rect 5001 12263 5057 12319
rect 5082 12263 5138 12319
rect 2733 12183 2789 12239
rect 2814 12183 2870 12239
rect 2895 12183 2951 12239
rect 2976 12183 3032 12239
rect 3057 12228 3113 12239
rect 3138 12228 3194 12239
rect 3057 12183 3101 12228
rect 3101 12183 3113 12228
rect 3138 12183 3153 12228
rect 3153 12183 3167 12228
rect 3167 12183 3194 12228
rect 3219 12183 3275 12239
rect 3300 12183 3356 12239
rect 3381 12183 3437 12239
rect 3462 12183 3518 12239
rect 3543 12183 3599 12239
rect 3624 12228 3680 12239
rect 3705 12228 3761 12239
rect 3624 12183 3655 12228
rect 3655 12183 3680 12228
rect 3705 12183 3707 12228
rect 3707 12183 3721 12228
rect 3721 12183 3761 12228
rect 3786 12183 3842 12239
rect 3867 12183 3923 12239
rect 3948 12183 4004 12239
rect 4029 12183 4085 12239
rect 4110 12183 4166 12239
rect 4191 12228 4247 12239
rect 4272 12228 4328 12239
rect 4191 12183 4209 12228
rect 4209 12183 4247 12228
rect 4272 12183 4275 12228
rect 4275 12183 4327 12228
rect 4327 12183 4328 12228
rect 4353 12183 4409 12239
rect 4434 12183 4490 12239
rect 4515 12183 4571 12239
rect 4596 12183 4652 12239
rect 4677 12183 4733 12239
rect 4758 12228 4814 12239
rect 4839 12228 4895 12239
rect 4758 12183 4763 12228
rect 4763 12183 4814 12228
rect 4839 12183 4881 12228
rect 4881 12183 4895 12228
rect 4920 12183 4976 12239
rect 5001 12183 5057 12239
rect 5082 12183 5138 12239
rect 2733 12103 2789 12159
rect 2814 12103 2870 12159
rect 2895 12103 2951 12159
rect 2976 12103 3032 12159
rect 3057 12158 3113 12159
rect 3138 12158 3194 12159
rect 3057 12106 3101 12158
rect 3101 12106 3113 12158
rect 3138 12106 3153 12158
rect 3153 12106 3167 12158
rect 3167 12106 3194 12158
rect 3057 12103 3113 12106
rect 3138 12103 3194 12106
rect 3219 12103 3275 12159
rect 3300 12103 3356 12159
rect 3381 12103 3437 12159
rect 3462 12103 3518 12159
rect 3543 12103 3599 12159
rect 3624 12158 3680 12159
rect 3705 12158 3761 12159
rect 3624 12106 3655 12158
rect 3655 12106 3680 12158
rect 3705 12106 3707 12158
rect 3707 12106 3721 12158
rect 3721 12106 3761 12158
rect 3624 12103 3680 12106
rect 3705 12103 3761 12106
rect 3786 12103 3842 12159
rect 3867 12103 3923 12159
rect 3948 12103 4004 12159
rect 4029 12103 4085 12159
rect 4110 12103 4166 12159
rect 4191 12158 4247 12159
rect 4272 12158 4328 12159
rect 4191 12106 4209 12158
rect 4209 12106 4247 12158
rect 4272 12106 4275 12158
rect 4275 12106 4327 12158
rect 4327 12106 4328 12158
rect 4191 12103 4247 12106
rect 4272 12103 4328 12106
rect 4353 12103 4409 12159
rect 4434 12103 4490 12159
rect 4515 12103 4571 12159
rect 4596 12103 4652 12159
rect 4677 12103 4733 12159
rect 4758 12158 4814 12159
rect 4839 12158 4895 12159
rect 4758 12106 4763 12158
rect 4763 12106 4814 12158
rect 4839 12106 4881 12158
rect 4881 12106 4895 12158
rect 4758 12103 4814 12106
rect 4839 12103 4895 12106
rect 4920 12103 4976 12159
rect 5001 12103 5057 12159
rect 5082 12103 5138 12159
rect 5163 12103 5299 12719
rect 5613 11452 5669 11456
rect 5696 11452 5752 11456
rect 5613 11400 5646 11452
rect 5646 11400 5660 11452
rect 5660 11400 5669 11452
rect 5696 11400 5712 11452
rect 5712 11400 5752 11452
rect 5779 11400 5835 11456
rect 5861 11400 5917 11456
rect 5943 11400 5999 11456
rect 6025 11400 6081 11456
rect 6107 11452 6163 11456
rect 6189 11452 6245 11456
rect 6107 11400 6148 11452
rect 6148 11400 6163 11452
rect 6189 11400 6200 11452
rect 6200 11400 6214 11452
rect 6214 11400 6245 11452
rect 6271 11400 6327 11456
rect 6353 11400 6409 11456
rect 6435 11400 6491 11456
rect 6517 11400 6573 11456
rect 6599 11400 6655 11456
rect 6681 11452 6737 11456
rect 6763 11452 6819 11456
rect 6681 11400 6702 11452
rect 6702 11400 6737 11452
rect 6763 11400 6768 11452
rect 6768 11400 6819 11452
rect 6845 11400 6901 11456
rect 6927 11400 6983 11456
rect 7009 11400 7065 11456
rect 7091 11400 7147 11456
rect 7173 11400 7229 11456
rect 7255 11452 7311 11456
rect 7337 11452 7393 11456
rect 7255 11400 7256 11452
rect 7256 11400 7308 11452
rect 7308 11400 7311 11452
rect 7337 11400 7374 11452
rect 7374 11400 7393 11452
rect 7419 11400 7475 11456
rect 7501 11400 7557 11456
rect 7583 11400 7639 11456
rect 7665 11400 7721 11456
rect 7747 11400 7803 11456
rect 7829 11452 7885 11456
rect 7911 11452 7967 11456
rect 7829 11400 7862 11452
rect 7862 11400 7876 11452
rect 7876 11400 7885 11452
rect 7911 11400 7928 11452
rect 7928 11400 7967 11452
rect 7993 11404 8047 11456
rect 8047 11404 8049 11456
rect 8075 11404 8099 11456
rect 8099 11404 8131 11456
rect 7993 11400 8049 11404
rect 8075 11400 8131 11404
rect 8157 11404 8169 11456
rect 8169 11404 8213 11456
rect 8157 11400 8213 11404
rect 5613 11331 5646 11376
rect 5646 11331 5660 11376
rect 5660 11331 5669 11376
rect 5696 11331 5712 11376
rect 5712 11331 5752 11376
rect 5613 11320 5669 11331
rect 5696 11320 5752 11331
rect 5779 11320 5835 11376
rect 5861 11320 5917 11376
rect 5943 11320 5999 11376
rect 6025 11320 6081 11376
rect 6107 11331 6148 11376
rect 6148 11331 6163 11376
rect 6189 11331 6200 11376
rect 6200 11331 6214 11376
rect 6214 11331 6245 11376
rect 6107 11320 6163 11331
rect 6189 11320 6245 11331
rect 6271 11320 6327 11376
rect 6353 11320 6409 11376
rect 6435 11320 6491 11376
rect 6517 11320 6573 11376
rect 6599 11320 6655 11376
rect 6681 11331 6702 11376
rect 6702 11331 6737 11376
rect 6763 11331 6768 11376
rect 6768 11331 6819 11376
rect 6681 11320 6737 11331
rect 6763 11320 6819 11331
rect 6845 11320 6901 11376
rect 6927 11320 6983 11376
rect 7009 11320 7065 11376
rect 7091 11320 7147 11376
rect 7173 11320 7229 11376
rect 7255 11331 7256 11376
rect 7256 11331 7308 11376
rect 7308 11331 7311 11376
rect 7337 11331 7374 11376
rect 7374 11331 7393 11376
rect 7255 11320 7311 11331
rect 7337 11320 7393 11331
rect 7419 11320 7475 11376
rect 7501 11320 7557 11376
rect 7583 11320 7639 11376
rect 7665 11320 7721 11376
rect 7747 11320 7803 11376
rect 7829 11331 7862 11376
rect 7862 11331 7876 11376
rect 7876 11331 7885 11376
rect 7911 11331 7928 11376
rect 7928 11331 7967 11376
rect 7829 11320 7885 11331
rect 7911 11320 7967 11331
rect 7993 11335 8047 11376
rect 8047 11335 8049 11376
rect 8075 11335 8099 11376
rect 8099 11335 8131 11376
rect 7993 11320 8049 11335
rect 8075 11320 8131 11335
rect 8157 11335 8169 11376
rect 8169 11335 8213 11376
rect 8157 11320 8213 11335
rect 5613 11262 5646 11296
rect 5646 11262 5660 11296
rect 5660 11262 5669 11296
rect 5696 11262 5712 11296
rect 5712 11262 5752 11296
rect 5613 11245 5669 11262
rect 5696 11245 5752 11262
rect 5613 11240 5646 11245
rect 5646 11240 5660 11245
rect 5660 11240 5669 11245
rect 5696 11240 5712 11245
rect 5712 11240 5752 11245
rect 5779 11240 5835 11296
rect 5861 11240 5917 11296
rect 5943 11240 5999 11296
rect 6025 11240 6081 11296
rect 6107 11262 6148 11296
rect 6148 11262 6163 11296
rect 6189 11262 6200 11296
rect 6200 11262 6214 11296
rect 6214 11262 6245 11296
rect 6107 11245 6163 11262
rect 6189 11245 6245 11262
rect 6107 11240 6148 11245
rect 6148 11240 6163 11245
rect 6189 11240 6200 11245
rect 6200 11240 6214 11245
rect 6214 11240 6245 11245
rect 6271 11240 6327 11296
rect 6353 11240 6409 11296
rect 6435 11240 6491 11296
rect 6517 11240 6573 11296
rect 6599 11240 6655 11296
rect 6681 11262 6702 11296
rect 6702 11262 6737 11296
rect 6763 11262 6768 11296
rect 6768 11262 6819 11296
rect 6681 11245 6737 11262
rect 6763 11245 6819 11262
rect 6681 11240 6702 11245
rect 6702 11240 6737 11245
rect 6763 11240 6768 11245
rect 6768 11240 6819 11245
rect 6845 11240 6901 11296
rect 6927 11240 6983 11296
rect 7009 11240 7065 11296
rect 7091 11240 7147 11296
rect 7173 11240 7229 11296
rect 7255 11262 7256 11296
rect 7256 11262 7308 11296
rect 7308 11262 7311 11296
rect 7337 11262 7374 11296
rect 7374 11262 7393 11296
rect 7255 11245 7311 11262
rect 7337 11245 7393 11262
rect 7255 11240 7256 11245
rect 7256 11240 7308 11245
rect 7308 11240 7311 11245
rect 7337 11240 7374 11245
rect 7374 11240 7393 11245
rect 7419 11240 7475 11296
rect 7501 11240 7557 11296
rect 7583 11240 7639 11296
rect 7665 11240 7721 11296
rect 7747 11240 7803 11296
rect 7829 11262 7862 11296
rect 7862 11262 7876 11296
rect 7876 11262 7885 11296
rect 7911 11262 7928 11296
rect 7928 11262 7967 11296
rect 7829 11245 7885 11262
rect 7911 11245 7967 11262
rect 7829 11240 7862 11245
rect 7862 11240 7876 11245
rect 7876 11240 7885 11245
rect 7911 11240 7928 11245
rect 7928 11240 7967 11245
rect 7993 11266 8047 11296
rect 8047 11266 8049 11296
rect 8075 11266 8099 11296
rect 8099 11266 8131 11296
rect 7993 11249 8049 11266
rect 8075 11249 8131 11266
rect 7993 11240 8047 11249
rect 8047 11240 8049 11249
rect 8075 11240 8099 11249
rect 8099 11240 8131 11249
rect 8157 11266 8169 11296
rect 8169 11266 8213 11296
rect 8157 11249 8213 11266
rect 8157 11240 8169 11249
rect 8169 11240 8213 11249
rect 5613 11193 5646 11216
rect 5646 11193 5660 11216
rect 5660 11193 5669 11216
rect 5696 11193 5712 11216
rect 5712 11193 5752 11216
rect 5613 11176 5669 11193
rect 5696 11176 5752 11193
rect 5613 11160 5646 11176
rect 5646 11160 5660 11176
rect 5660 11160 5669 11176
rect 5696 11160 5712 11176
rect 5712 11160 5752 11176
rect 5779 11160 5835 11216
rect 5861 11160 5917 11216
rect 5943 11160 5999 11216
rect 6025 11160 6081 11216
rect 6107 11193 6148 11216
rect 6148 11193 6163 11216
rect 6189 11193 6200 11216
rect 6200 11193 6214 11216
rect 6214 11193 6245 11216
rect 6107 11176 6163 11193
rect 6189 11176 6245 11193
rect 6107 11160 6148 11176
rect 6148 11160 6163 11176
rect 6189 11160 6200 11176
rect 6200 11160 6214 11176
rect 6214 11160 6245 11176
rect 6271 11160 6327 11216
rect 6353 11160 6409 11216
rect 6435 11160 6491 11216
rect 6517 11160 6573 11216
rect 6599 11160 6655 11216
rect 6681 11193 6702 11216
rect 6702 11193 6737 11216
rect 6763 11193 6768 11216
rect 6768 11193 6819 11216
rect 6681 11176 6737 11193
rect 6763 11176 6819 11193
rect 6681 11160 6702 11176
rect 6702 11160 6737 11176
rect 6763 11160 6768 11176
rect 6768 11160 6819 11176
rect 6845 11160 6901 11216
rect 6927 11160 6983 11216
rect 7009 11160 7065 11216
rect 7091 11160 7147 11216
rect 7173 11160 7229 11216
rect 7255 11193 7256 11216
rect 7256 11193 7308 11216
rect 7308 11193 7311 11216
rect 7337 11193 7374 11216
rect 7374 11193 7393 11216
rect 7255 11176 7311 11193
rect 7337 11176 7393 11193
rect 7255 11160 7256 11176
rect 7256 11160 7308 11176
rect 7308 11160 7311 11176
rect 7337 11160 7374 11176
rect 7374 11160 7393 11176
rect 7419 11160 7475 11216
rect 7501 11160 7557 11216
rect 7583 11160 7639 11216
rect 7665 11160 7721 11216
rect 7747 11160 7803 11216
rect 7829 11193 7862 11216
rect 7862 11193 7876 11216
rect 7876 11193 7885 11216
rect 7911 11193 7928 11216
rect 7928 11193 7967 11216
rect 7829 11176 7885 11193
rect 7911 11176 7967 11193
rect 7829 11160 7862 11176
rect 7862 11160 7876 11176
rect 7876 11160 7885 11176
rect 7911 11160 7928 11176
rect 7928 11160 7967 11176
rect 7993 11197 8047 11216
rect 8047 11197 8049 11216
rect 8075 11197 8099 11216
rect 8099 11197 8131 11216
rect 7993 11180 8049 11197
rect 8075 11180 8131 11197
rect 7993 11160 8047 11180
rect 8047 11160 8049 11180
rect 8075 11160 8099 11180
rect 8099 11160 8131 11180
rect 8157 11197 8169 11216
rect 8169 11197 8213 11216
rect 8157 11180 8213 11197
rect 8157 11160 8169 11180
rect 8169 11160 8213 11180
rect 5613 11124 5646 11136
rect 5646 11124 5660 11136
rect 5660 11124 5669 11136
rect 5696 11124 5712 11136
rect 5712 11124 5752 11136
rect 5613 11107 5669 11124
rect 5696 11107 5752 11124
rect 5613 11080 5646 11107
rect 5646 11080 5660 11107
rect 5660 11080 5669 11107
rect 5696 11080 5712 11107
rect 5712 11080 5752 11107
rect 5779 11080 5835 11136
rect 5861 11080 5917 11136
rect 5943 11080 5999 11136
rect 6025 11080 6081 11136
rect 6107 11124 6148 11136
rect 6148 11124 6163 11136
rect 6189 11124 6200 11136
rect 6200 11124 6214 11136
rect 6214 11124 6245 11136
rect 6107 11107 6163 11124
rect 6189 11107 6245 11124
rect 6107 11080 6148 11107
rect 6148 11080 6163 11107
rect 6189 11080 6200 11107
rect 6200 11080 6214 11107
rect 6214 11080 6245 11107
rect 6271 11080 6327 11136
rect 6353 11080 6409 11136
rect 6435 11080 6491 11136
rect 6517 11080 6573 11136
rect 6599 11080 6655 11136
rect 6681 11124 6702 11136
rect 6702 11124 6737 11136
rect 6763 11124 6768 11136
rect 6768 11124 6819 11136
rect 6681 11107 6737 11124
rect 6763 11107 6819 11124
rect 6681 11080 6702 11107
rect 6702 11080 6737 11107
rect 6763 11080 6768 11107
rect 6768 11080 6819 11107
rect 6845 11080 6901 11136
rect 6927 11080 6983 11136
rect 7009 11080 7065 11136
rect 7091 11080 7147 11136
rect 7173 11080 7229 11136
rect 7255 11124 7256 11136
rect 7256 11124 7308 11136
rect 7308 11124 7311 11136
rect 7337 11124 7374 11136
rect 7374 11124 7393 11136
rect 7255 11107 7311 11124
rect 7337 11107 7393 11124
rect 7255 11080 7256 11107
rect 7256 11080 7308 11107
rect 7308 11080 7311 11107
rect 7337 11080 7374 11107
rect 7374 11080 7393 11107
rect 7419 11080 7475 11136
rect 7501 11080 7557 11136
rect 7583 11080 7639 11136
rect 7665 11080 7721 11136
rect 7747 11080 7803 11136
rect 7829 11124 7862 11136
rect 7862 11124 7876 11136
rect 7876 11124 7885 11136
rect 7911 11124 7928 11136
rect 7928 11124 7967 11136
rect 7829 11107 7885 11124
rect 7911 11107 7967 11124
rect 7829 11080 7862 11107
rect 7862 11080 7876 11107
rect 7876 11080 7885 11107
rect 7911 11080 7928 11107
rect 7928 11080 7967 11107
rect 7993 11128 8047 11136
rect 8047 11128 8049 11136
rect 8075 11128 8099 11136
rect 8099 11128 8131 11136
rect 7993 11110 8049 11128
rect 8075 11110 8131 11128
rect 7993 11080 8047 11110
rect 8047 11080 8049 11110
rect 8075 11080 8099 11110
rect 8099 11080 8131 11110
rect 8157 11128 8169 11136
rect 8169 11128 8213 11136
rect 8157 11110 8213 11128
rect 8157 11080 8169 11110
rect 8169 11080 8213 11110
rect 5613 11055 5646 11056
rect 5646 11055 5660 11056
rect 5660 11055 5669 11056
rect 5696 11055 5712 11056
rect 5712 11055 5752 11056
rect 5613 11038 5669 11055
rect 5696 11038 5752 11055
rect 5613 11000 5646 11038
rect 5646 11000 5660 11038
rect 5660 11000 5669 11038
rect 5696 11000 5712 11038
rect 5712 11000 5752 11038
rect 5779 11000 5835 11056
rect 5861 11000 5917 11056
rect 5943 11000 5999 11056
rect 6025 11000 6081 11056
rect 6107 11055 6148 11056
rect 6148 11055 6163 11056
rect 6189 11055 6200 11056
rect 6200 11055 6214 11056
rect 6214 11055 6245 11056
rect 6107 11038 6163 11055
rect 6189 11038 6245 11055
rect 6107 11000 6148 11038
rect 6148 11000 6163 11038
rect 6189 11000 6200 11038
rect 6200 11000 6214 11038
rect 6214 11000 6245 11038
rect 6271 11000 6327 11056
rect 6353 11000 6409 11056
rect 6435 11000 6491 11056
rect 6517 11000 6573 11056
rect 6599 11000 6655 11056
rect 6681 11055 6702 11056
rect 6702 11055 6737 11056
rect 6763 11055 6768 11056
rect 6768 11055 6819 11056
rect 6681 11038 6737 11055
rect 6763 11038 6819 11055
rect 6681 11000 6702 11038
rect 6702 11000 6737 11038
rect 6763 11000 6768 11038
rect 6768 11000 6819 11038
rect 6845 11000 6901 11056
rect 6927 11000 6983 11056
rect 7009 11000 7065 11056
rect 7091 11000 7147 11056
rect 7173 11000 7229 11056
rect 7255 11055 7256 11056
rect 7256 11055 7308 11056
rect 7308 11055 7311 11056
rect 7337 11055 7374 11056
rect 7374 11055 7393 11056
rect 7255 11038 7311 11055
rect 7337 11038 7393 11055
rect 7255 11000 7256 11038
rect 7256 11000 7308 11038
rect 7308 11000 7311 11038
rect 7337 11000 7374 11038
rect 7374 11000 7393 11038
rect 7419 11000 7475 11056
rect 7501 11000 7557 11056
rect 7583 11000 7639 11056
rect 7665 11000 7721 11056
rect 7747 11000 7803 11056
rect 7829 11055 7862 11056
rect 7862 11055 7876 11056
rect 7876 11055 7885 11056
rect 7911 11055 7928 11056
rect 7928 11055 7967 11056
rect 7829 11038 7885 11055
rect 7911 11038 7967 11055
rect 7829 11000 7862 11038
rect 7862 11000 7876 11038
rect 7876 11000 7885 11038
rect 7911 11000 7928 11038
rect 7928 11000 7967 11038
rect 7993 11040 8049 11056
rect 8075 11040 8131 11056
rect 7993 11000 8047 11040
rect 8047 11000 8049 11040
rect 8075 11000 8099 11040
rect 8099 11000 8131 11040
rect 8157 11040 8213 11056
rect 8157 11000 8169 11040
rect 8169 11000 8213 11040
rect 5613 10968 5669 10976
rect 5696 10968 5752 10976
rect 5613 10920 5646 10968
rect 5646 10920 5660 10968
rect 5660 10920 5669 10968
rect 5696 10920 5712 10968
rect 5712 10920 5752 10968
rect 5779 10920 5835 10976
rect 5861 10920 5917 10976
rect 5943 10920 5999 10976
rect 6025 10920 6081 10976
rect 6107 10968 6163 10976
rect 6189 10968 6245 10976
rect 6107 10920 6148 10968
rect 6148 10920 6163 10968
rect 6189 10920 6200 10968
rect 6200 10920 6214 10968
rect 6214 10920 6245 10968
rect 6271 10920 6327 10976
rect 6353 10920 6409 10976
rect 6435 10920 6491 10976
rect 6517 10920 6573 10976
rect 6599 10920 6655 10976
rect 6681 10968 6737 10976
rect 6763 10968 6819 10976
rect 6681 10920 6702 10968
rect 6702 10920 6737 10968
rect 6763 10920 6768 10968
rect 6768 10920 6819 10968
rect 6845 10920 6901 10976
rect 6927 10920 6983 10976
rect 7009 10920 7065 10976
rect 7091 10920 7147 10976
rect 7173 10920 7229 10976
rect 7255 10968 7311 10976
rect 7337 10968 7393 10976
rect 7255 10920 7256 10968
rect 7256 10920 7308 10968
rect 7308 10920 7311 10968
rect 7337 10920 7374 10968
rect 7374 10920 7393 10968
rect 7419 10920 7475 10976
rect 7501 10920 7557 10976
rect 7583 10920 7639 10976
rect 7665 10920 7721 10976
rect 7747 10920 7803 10976
rect 7829 10968 7885 10976
rect 7911 10968 7967 10976
rect 7829 10920 7862 10968
rect 7862 10920 7876 10968
rect 7876 10920 7885 10968
rect 7911 10920 7928 10968
rect 7928 10920 7967 10968
rect 7993 10970 8049 10976
rect 8075 10970 8131 10976
rect 7993 10920 8047 10970
rect 8047 10920 8049 10970
rect 8075 10920 8099 10970
rect 8099 10920 8131 10970
rect 8157 10970 8213 10976
rect 8157 10920 8169 10970
rect 8169 10920 8213 10970
rect 5613 10846 5646 10896
rect 5646 10846 5660 10896
rect 5660 10846 5669 10896
rect 5696 10846 5712 10896
rect 5712 10846 5752 10896
rect 5613 10840 5669 10846
rect 5696 10840 5752 10846
rect 5779 10840 5835 10896
rect 5861 10840 5917 10896
rect 5943 10840 5999 10896
rect 6025 10840 6081 10896
rect 6107 10846 6148 10896
rect 6148 10846 6163 10896
rect 6189 10846 6200 10896
rect 6200 10846 6214 10896
rect 6214 10846 6245 10896
rect 6107 10840 6163 10846
rect 6189 10840 6245 10846
rect 6271 10840 6327 10896
rect 6353 10840 6409 10896
rect 6435 10840 6491 10896
rect 6517 10840 6573 10896
rect 6599 10840 6655 10896
rect 6681 10846 6702 10896
rect 6702 10846 6737 10896
rect 6763 10846 6768 10896
rect 6768 10846 6819 10896
rect 6681 10840 6737 10846
rect 6763 10840 6819 10846
rect 6845 10840 6901 10896
rect 6927 10840 6983 10896
rect 7009 10840 7065 10896
rect 7091 10840 7147 10896
rect 7173 10840 7229 10896
rect 7255 10846 7256 10896
rect 7256 10846 7308 10896
rect 7308 10846 7311 10896
rect 7337 10846 7374 10896
rect 7374 10846 7393 10896
rect 7255 10840 7311 10846
rect 7337 10840 7393 10846
rect 7419 10840 7475 10896
rect 7501 10840 7557 10896
rect 7583 10840 7639 10896
rect 7665 10840 7721 10896
rect 7747 10840 7803 10896
rect 7829 10846 7862 10896
rect 7862 10846 7876 10896
rect 7876 10846 7885 10896
rect 7911 10846 7928 10896
rect 7928 10846 7967 10896
rect 7829 10840 7885 10846
rect 7911 10840 7967 10846
rect 7993 10848 8047 10896
rect 8047 10848 8049 10896
rect 8075 10848 8099 10896
rect 8099 10848 8131 10896
rect 7993 10840 8049 10848
rect 8075 10840 8131 10848
rect 8157 10848 8169 10896
rect 8169 10848 8213 10896
rect 8157 10840 8213 10848
rect 2859 10664 2915 10720
rect 2942 10664 2998 10720
rect 3025 10664 3081 10720
rect 3108 10714 3164 10720
rect 3191 10714 3247 10720
rect 3108 10664 3153 10714
rect 3153 10664 3164 10714
rect 3191 10664 3219 10714
rect 3219 10664 3247 10714
rect 3274 10664 3330 10720
rect 3357 10664 3413 10720
rect 3439 10664 3495 10720
rect 3521 10664 3577 10720
rect 3603 10714 3659 10720
rect 3685 10714 3741 10720
rect 3767 10714 3823 10720
rect 3603 10664 3655 10714
rect 3655 10664 3659 10714
rect 3685 10664 3707 10714
rect 3707 10664 3721 10714
rect 3721 10664 3741 10714
rect 3767 10664 3773 10714
rect 3773 10664 3823 10714
rect 3849 10664 3905 10720
rect 3931 10664 3987 10720
rect 4013 10664 4069 10720
rect 4095 10664 4151 10720
rect 4177 10714 4233 10720
rect 4259 10714 4315 10720
rect 4177 10664 4209 10714
rect 4209 10664 4233 10714
rect 4259 10664 4261 10714
rect 4261 10664 4275 10714
rect 4275 10664 4315 10714
rect 4341 10664 4397 10720
rect 4423 10664 4479 10720
rect 4505 10664 4561 10720
rect 4587 10664 4643 10720
rect 4669 10664 4725 10720
rect 4751 10714 4807 10720
rect 4833 10714 4889 10720
rect 4751 10664 4763 10714
rect 4763 10664 4807 10714
rect 4833 10664 4881 10714
rect 4881 10664 4889 10714
rect 4915 10664 4971 10720
rect 4997 10664 5053 10720
rect 5079 10664 5135 10720
rect 5161 10664 5217 10720
rect 5243 10664 5299 10720
rect 2859 10584 2915 10640
rect 2942 10584 2998 10640
rect 3025 10584 3081 10640
rect 3108 10593 3153 10640
rect 3153 10593 3164 10640
rect 3191 10593 3219 10640
rect 3219 10593 3247 10640
rect 3108 10584 3164 10593
rect 3191 10584 3247 10593
rect 3274 10584 3330 10640
rect 3357 10584 3413 10640
rect 3439 10584 3495 10640
rect 3521 10584 3577 10640
rect 3603 10593 3655 10640
rect 3655 10593 3659 10640
rect 3685 10593 3707 10640
rect 3707 10593 3721 10640
rect 3721 10593 3741 10640
rect 3767 10593 3773 10640
rect 3773 10593 3823 10640
rect 3603 10584 3659 10593
rect 3685 10584 3741 10593
rect 3767 10584 3823 10593
rect 3849 10584 3905 10640
rect 3931 10584 3987 10640
rect 4013 10584 4069 10640
rect 4095 10584 4151 10640
rect 4177 10593 4209 10640
rect 4209 10593 4233 10640
rect 4259 10593 4261 10640
rect 4261 10593 4275 10640
rect 4275 10593 4315 10640
rect 4177 10584 4233 10593
rect 4259 10584 4315 10593
rect 4341 10584 4397 10640
rect 4423 10584 4479 10640
rect 4505 10584 4561 10640
rect 4587 10584 4643 10640
rect 4669 10584 4725 10640
rect 4751 10593 4763 10640
rect 4763 10593 4807 10640
rect 4833 10593 4881 10640
rect 4881 10593 4889 10640
rect 4751 10584 4807 10593
rect 4833 10584 4889 10593
rect 4915 10584 4971 10640
rect 4997 10584 5053 10640
rect 5079 10584 5135 10640
rect 5161 10584 5217 10640
rect 5243 10584 5299 10640
rect 2859 10504 2915 10560
rect 2942 10504 2998 10560
rect 3025 10504 3081 10560
rect 3108 10524 3153 10560
rect 3153 10524 3164 10560
rect 3191 10524 3219 10560
rect 3219 10524 3247 10560
rect 3108 10507 3164 10524
rect 3191 10507 3247 10524
rect 3108 10504 3153 10507
rect 3153 10504 3164 10507
rect 3191 10504 3219 10507
rect 3219 10504 3247 10507
rect 3274 10504 3330 10560
rect 3357 10504 3413 10560
rect 3439 10504 3495 10560
rect 3521 10504 3577 10560
rect 3603 10524 3655 10560
rect 3655 10524 3659 10560
rect 3685 10524 3707 10560
rect 3707 10524 3721 10560
rect 3721 10524 3741 10560
rect 3767 10524 3773 10560
rect 3773 10524 3823 10560
rect 3603 10507 3659 10524
rect 3685 10507 3741 10524
rect 3767 10507 3823 10524
rect 3603 10504 3655 10507
rect 3655 10504 3659 10507
rect 3685 10504 3707 10507
rect 3707 10504 3721 10507
rect 3721 10504 3741 10507
rect 3767 10504 3773 10507
rect 3773 10504 3823 10507
rect 3849 10504 3905 10560
rect 3931 10504 3987 10560
rect 4013 10504 4069 10560
rect 4095 10504 4151 10560
rect 4177 10524 4209 10560
rect 4209 10524 4233 10560
rect 4259 10524 4261 10560
rect 4261 10524 4275 10560
rect 4275 10524 4315 10560
rect 4177 10507 4233 10524
rect 4259 10507 4315 10524
rect 4177 10504 4209 10507
rect 4209 10504 4233 10507
rect 4259 10504 4261 10507
rect 4261 10504 4275 10507
rect 4275 10504 4315 10507
rect 4341 10504 4397 10560
rect 4423 10504 4479 10560
rect 4505 10504 4561 10560
rect 4587 10504 4643 10560
rect 4669 10504 4725 10560
rect 4751 10524 4763 10560
rect 4763 10524 4807 10560
rect 4833 10524 4881 10560
rect 4881 10524 4889 10560
rect 4751 10507 4807 10524
rect 4833 10507 4889 10524
rect 4751 10504 4763 10507
rect 4763 10504 4807 10507
rect 2859 10424 2915 10480
rect 2942 10424 2998 10480
rect 3025 10424 3081 10480
rect 3108 10455 3153 10480
rect 3153 10455 3164 10480
rect 3191 10455 3219 10480
rect 3219 10455 3247 10480
rect 3108 10438 3164 10455
rect 3191 10438 3247 10455
rect 3108 10424 3153 10438
rect 3153 10424 3164 10438
rect 3191 10424 3219 10438
rect 3219 10424 3247 10438
rect 3274 10424 3330 10480
rect 3357 10424 3413 10480
rect 3439 10424 3495 10480
rect 3521 10424 3577 10480
rect 3603 10455 3655 10480
rect 3655 10455 3659 10480
rect 3685 10455 3707 10480
rect 3707 10455 3721 10480
rect 3721 10455 3741 10480
rect 3767 10455 3773 10480
rect 3773 10455 3823 10480
rect 3603 10438 3659 10455
rect 3685 10438 3741 10455
rect 3767 10438 3823 10455
rect 3603 10424 3655 10438
rect 3655 10424 3659 10438
rect 3685 10424 3707 10438
rect 3707 10424 3721 10438
rect 3721 10424 3741 10438
rect 3767 10424 3773 10438
rect 3773 10424 3823 10438
rect 3849 10424 3905 10480
rect 3931 10424 3987 10480
rect 4013 10424 4069 10480
rect 4095 10424 4151 10480
rect 4177 10455 4209 10480
rect 4209 10455 4233 10480
rect 4259 10455 4261 10480
rect 4261 10455 4275 10480
rect 4275 10455 4315 10480
rect 4177 10438 4233 10455
rect 4259 10438 4315 10455
rect 4177 10424 4209 10438
rect 4209 10424 4233 10438
rect 4259 10424 4261 10438
rect 4261 10424 4275 10438
rect 4275 10424 4315 10438
rect 4341 10424 4397 10480
rect 4423 10424 4479 10480
rect 4505 10424 4561 10480
rect 4587 10424 4643 10480
rect 4669 10424 4725 10480
rect 4751 10455 4763 10480
rect 4763 10455 4807 10480
rect 4833 10504 4881 10507
rect 4881 10504 4889 10507
rect 4915 10504 4971 10560
rect 4997 10504 5053 10560
rect 5079 10504 5135 10560
rect 5161 10504 5217 10560
rect 5243 10504 5299 10560
rect 4833 10455 4881 10480
rect 4881 10455 4889 10480
rect 4751 10438 4807 10455
rect 4833 10438 4889 10455
rect 4751 10424 4763 10438
rect 4763 10424 4807 10438
rect 2859 10344 2915 10400
rect 2942 10344 2998 10400
rect 3025 10344 3081 10400
rect 3108 10386 3153 10400
rect 3153 10386 3164 10400
rect 3191 10386 3219 10400
rect 3219 10386 3247 10400
rect 3108 10368 3164 10386
rect 3191 10368 3247 10386
rect 3108 10344 3153 10368
rect 3153 10344 3164 10368
rect 3191 10344 3219 10368
rect 3219 10344 3247 10368
rect 3274 10344 3330 10400
rect 3357 10344 3413 10400
rect 3439 10344 3495 10400
rect 3521 10344 3577 10400
rect 3603 10386 3655 10400
rect 3655 10386 3659 10400
rect 3685 10386 3707 10400
rect 3707 10386 3721 10400
rect 3721 10386 3741 10400
rect 3767 10386 3773 10400
rect 3773 10386 3823 10400
rect 3603 10368 3659 10386
rect 3685 10368 3741 10386
rect 3767 10368 3823 10386
rect 3603 10344 3655 10368
rect 3655 10344 3659 10368
rect 3685 10344 3707 10368
rect 3707 10344 3721 10368
rect 3721 10344 3741 10368
rect 3767 10344 3773 10368
rect 3773 10344 3823 10368
rect 3849 10344 3905 10400
rect 3931 10344 3987 10400
rect 4013 10344 4069 10400
rect 4095 10344 4151 10400
rect 4177 10386 4209 10400
rect 4209 10386 4233 10400
rect 4259 10386 4261 10400
rect 4261 10386 4275 10400
rect 4275 10386 4315 10400
rect 4177 10368 4233 10386
rect 4259 10368 4315 10386
rect 4177 10344 4209 10368
rect 4209 10344 4233 10368
rect 4259 10344 4261 10368
rect 4261 10344 4275 10368
rect 4275 10344 4315 10368
rect 4341 10344 4397 10400
rect 4423 10344 4479 10400
rect 4505 10344 4561 10400
rect 4587 10344 4643 10400
rect 4669 10344 4725 10400
rect 4751 10386 4763 10400
rect 4763 10386 4807 10400
rect 4833 10424 4881 10438
rect 4881 10424 4889 10438
rect 4915 10424 4971 10480
rect 4997 10424 5053 10480
rect 5079 10424 5135 10480
rect 5161 10424 5217 10480
rect 5243 10424 5299 10480
rect 4833 10386 4881 10400
rect 4881 10386 4889 10400
rect 4751 10368 4807 10386
rect 4833 10368 4889 10386
rect 4751 10344 4763 10368
rect 4763 10344 4807 10368
rect 2859 10264 2915 10320
rect 2942 10264 2998 10320
rect 3025 10264 3081 10320
rect 3108 10316 3153 10320
rect 3153 10316 3164 10320
rect 3191 10316 3219 10320
rect 3219 10316 3247 10320
rect 3108 10298 3164 10316
rect 3191 10298 3247 10316
rect 3108 10264 3153 10298
rect 3153 10264 3164 10298
rect 3191 10264 3219 10298
rect 3219 10264 3247 10298
rect 3274 10264 3330 10320
rect 3357 10264 3413 10320
rect 3439 10264 3495 10320
rect 3521 10264 3577 10320
rect 3603 10316 3655 10320
rect 3655 10316 3659 10320
rect 3685 10316 3707 10320
rect 3707 10316 3721 10320
rect 3721 10316 3741 10320
rect 3767 10316 3773 10320
rect 3773 10316 3823 10320
rect 3603 10298 3659 10316
rect 3685 10298 3741 10316
rect 3767 10298 3823 10316
rect 3603 10264 3655 10298
rect 3655 10264 3659 10298
rect 3685 10264 3707 10298
rect 3707 10264 3721 10298
rect 3721 10264 3741 10298
rect 3767 10264 3773 10298
rect 3773 10264 3823 10298
rect 3849 10264 3905 10320
rect 3931 10264 3987 10320
rect 4013 10264 4069 10320
rect 4095 10264 4151 10320
rect 4177 10316 4209 10320
rect 4209 10316 4233 10320
rect 4259 10316 4261 10320
rect 4261 10316 4275 10320
rect 4275 10316 4315 10320
rect 4177 10298 4233 10316
rect 4259 10298 4315 10316
rect 4177 10264 4209 10298
rect 4209 10264 4233 10298
rect 4259 10264 4261 10298
rect 4261 10264 4275 10298
rect 4275 10264 4315 10298
rect 4341 10264 4397 10320
rect 4423 10264 4479 10320
rect 4505 10264 4561 10320
rect 4587 10264 4643 10320
rect 4669 10264 4725 10320
rect 4751 10316 4763 10320
rect 4763 10316 4807 10320
rect 4833 10344 4881 10368
rect 4881 10344 4889 10368
rect 4915 10344 4971 10400
rect 4997 10344 5053 10400
rect 5079 10344 5135 10400
rect 5161 10344 5217 10400
rect 5243 10344 5299 10400
rect 4833 10316 4881 10320
rect 4881 10316 4889 10320
rect 4751 10298 4807 10316
rect 4833 10298 4889 10316
rect 4751 10264 4763 10298
rect 4763 10264 4807 10298
rect 4833 10264 4881 10298
rect 4881 10264 4889 10298
rect 4915 10264 4971 10320
rect 4997 10264 5053 10320
rect 5079 10264 5135 10320
rect 5161 10264 5217 10320
rect 5243 10264 5299 10320
rect 2859 10184 2915 10240
rect 2942 10184 2998 10240
rect 3025 10184 3081 10240
rect 3108 10228 3164 10240
rect 3191 10228 3247 10240
rect 3108 10184 3153 10228
rect 3153 10184 3164 10228
rect 3191 10184 3219 10228
rect 3219 10184 3247 10228
rect 3274 10184 3330 10240
rect 3357 10184 3413 10240
rect 3439 10184 3495 10240
rect 3521 10184 3577 10240
rect 3603 10228 3659 10240
rect 3685 10228 3741 10240
rect 3767 10228 3823 10240
rect 3603 10184 3655 10228
rect 3655 10184 3659 10228
rect 3685 10184 3707 10228
rect 3707 10184 3721 10228
rect 3721 10184 3741 10228
rect 3767 10184 3773 10228
rect 3773 10184 3823 10228
rect 3849 10184 3905 10240
rect 3931 10184 3987 10240
rect 4013 10184 4069 10240
rect 4095 10184 4151 10240
rect 4177 10228 4233 10240
rect 4259 10228 4315 10240
rect 4177 10184 4209 10228
rect 4209 10184 4233 10228
rect 4259 10184 4261 10228
rect 4261 10184 4275 10228
rect 4275 10184 4315 10228
rect 4341 10184 4397 10240
rect 4423 10184 4479 10240
rect 4505 10184 4561 10240
rect 4587 10184 4643 10240
rect 4669 10184 4725 10240
rect 4751 10228 4807 10240
rect 4833 10228 4889 10240
rect 4751 10184 4763 10228
rect 4763 10184 4807 10228
rect 4833 10184 4881 10228
rect 4881 10184 4889 10228
rect 4915 10184 4971 10240
rect 4997 10184 5053 10240
rect 5079 10184 5135 10240
rect 5161 10184 5217 10240
rect 5243 10184 5299 10240
rect 2859 10104 2915 10160
rect 2942 10104 2998 10160
rect 3025 10104 3081 10160
rect 3108 10158 3164 10160
rect 3191 10158 3247 10160
rect 3108 10106 3153 10158
rect 3153 10106 3164 10158
rect 3191 10106 3219 10158
rect 3219 10106 3247 10158
rect 3108 10104 3164 10106
rect 3191 10104 3247 10106
rect 3274 10104 3330 10160
rect 3357 10104 3413 10160
rect 3439 10104 3495 10160
rect 3521 10104 3577 10160
rect 3603 10158 3659 10160
rect 3685 10158 3741 10160
rect 3767 10158 3823 10160
rect 3603 10106 3655 10158
rect 3655 10106 3659 10158
rect 3685 10106 3707 10158
rect 3707 10106 3721 10158
rect 3721 10106 3741 10158
rect 3767 10106 3773 10158
rect 3773 10106 3823 10158
rect 3603 10104 3659 10106
rect 3685 10104 3741 10106
rect 3767 10104 3823 10106
rect 3849 10104 3905 10160
rect 3931 10104 3987 10160
rect 4013 10104 4069 10160
rect 4095 10104 4151 10160
rect 4177 10158 4233 10160
rect 4259 10158 4315 10160
rect 4177 10106 4209 10158
rect 4209 10106 4233 10158
rect 4259 10106 4261 10158
rect 4261 10106 4275 10158
rect 4275 10106 4315 10158
rect 4177 10104 4233 10106
rect 4259 10104 4315 10106
rect 4341 10104 4397 10160
rect 4423 10104 4479 10160
rect 4505 10104 4561 10160
rect 4587 10104 4643 10160
rect 4669 10104 4725 10160
rect 4751 10158 4807 10160
rect 4833 10158 4889 10160
rect 4751 10106 4763 10158
rect 4763 10106 4807 10158
rect 4833 10106 4881 10158
rect 4881 10106 4889 10158
rect 4751 10104 4807 10106
rect 4833 10104 4889 10106
rect 4915 10104 4971 10160
rect 4997 10104 5053 10160
rect 5079 10104 5135 10160
rect 5161 10104 5217 10160
rect 5243 10104 5299 10160
rect 5617 9458 5673 9460
rect 5698 9458 5754 9460
rect 5779 9458 5835 9460
rect 5860 9458 5916 9460
rect 5941 9458 5997 9460
rect 6022 9458 6078 9460
rect 6103 9458 6159 9460
rect 6184 9458 6240 9460
rect 6265 9458 6321 9460
rect 6346 9458 6402 9460
rect 6427 9458 6483 9460
rect 6508 9458 6564 9460
rect 6589 9458 6645 9460
rect 6669 9458 6725 9460
rect 6749 9458 6805 9460
rect 6829 9458 6885 9460
rect 6909 9458 6965 9460
rect 6989 9458 7045 9460
rect 7069 9458 7125 9460
rect 7149 9458 7205 9460
rect 7229 9458 7285 9460
rect 7309 9458 7365 9460
rect 5617 9406 5640 9458
rect 5640 9406 5652 9458
rect 5652 9406 5673 9458
rect 5698 9406 5704 9458
rect 5704 9406 5716 9458
rect 5716 9406 5754 9458
rect 5779 9406 5780 9458
rect 5780 9406 5832 9458
rect 5832 9406 5835 9458
rect 5860 9406 5896 9458
rect 5896 9406 5908 9458
rect 5908 9406 5916 9458
rect 5941 9406 5960 9458
rect 5960 9406 5972 9458
rect 5972 9406 5997 9458
rect 6022 9406 6024 9458
rect 6024 9406 6036 9458
rect 6036 9406 6078 9458
rect 6103 9406 6152 9458
rect 6152 9406 6159 9458
rect 6184 9406 6216 9458
rect 6216 9406 6228 9458
rect 6228 9406 6240 9458
rect 6265 9406 6280 9458
rect 6280 9406 6292 9458
rect 6292 9406 6321 9458
rect 6346 9406 6356 9458
rect 6356 9406 6402 9458
rect 6427 9406 6472 9458
rect 6472 9406 6483 9458
rect 6508 9406 6536 9458
rect 6536 9406 6548 9458
rect 6548 9406 6564 9458
rect 6589 9406 6600 9458
rect 6600 9406 6612 9458
rect 6612 9406 6645 9458
rect 6669 9406 6676 9458
rect 6676 9406 6725 9458
rect 6749 9406 6792 9458
rect 6792 9406 6804 9458
rect 6804 9406 6805 9458
rect 6829 9406 6856 9458
rect 6856 9406 6868 9458
rect 6868 9406 6885 9458
rect 6909 9406 6920 9458
rect 6920 9406 6932 9458
rect 6932 9406 6965 9458
rect 6989 9406 6996 9458
rect 6996 9406 7045 9458
rect 7069 9406 7112 9458
rect 7112 9406 7124 9458
rect 7124 9406 7125 9458
rect 7149 9406 7176 9458
rect 7176 9406 7188 9458
rect 7188 9406 7205 9458
rect 7229 9406 7240 9458
rect 7240 9406 7252 9458
rect 7252 9406 7285 9458
rect 7309 9406 7316 9458
rect 7316 9406 7365 9458
rect 5617 9404 5673 9406
rect 5698 9404 5754 9406
rect 5779 9404 5835 9406
rect 5860 9404 5916 9406
rect 5941 9404 5997 9406
rect 6022 9404 6078 9406
rect 6103 9404 6159 9406
rect 6184 9404 6240 9406
rect 6265 9404 6321 9406
rect 6346 9404 6402 9406
rect 6427 9404 6483 9406
rect 6508 9404 6564 9406
rect 6589 9404 6645 9406
rect 6669 9404 6725 9406
rect 6749 9404 6805 9406
rect 6829 9404 6885 9406
rect 6909 9404 6965 9406
rect 6989 9404 7045 9406
rect 7069 9404 7125 9406
rect 7149 9404 7205 9406
rect 7229 9404 7285 9406
rect 7309 9404 7365 9406
rect 5621 8657 5677 8713
rect 5705 8657 5761 8713
rect 5789 8657 5845 8713
rect 5873 8657 5929 8713
rect 5957 8657 6013 8713
rect 6041 8657 6097 8713
rect 6125 8657 6181 8713
rect 6209 8657 6265 8713
rect 6293 8657 6349 8713
rect 6377 8657 6433 8713
rect 6461 8657 6517 8713
rect 6545 8657 6601 8713
rect 6629 8657 6685 8713
rect 6713 8657 6769 8713
rect 6797 8657 6853 8713
rect 6881 8657 6937 8713
rect 6965 8657 7021 8713
rect 7048 8657 7104 8713
rect 7131 8657 7187 8713
rect 7214 8657 7270 8713
rect 7297 8657 7353 8713
rect 5621 8577 5677 8633
rect 5705 8577 5761 8633
rect 5789 8577 5845 8633
rect 5873 8577 5929 8633
rect 5957 8577 6013 8633
rect 6041 8577 6097 8633
rect 6125 8577 6181 8633
rect 6209 8577 6265 8633
rect 6293 8577 6349 8633
rect 6377 8577 6433 8633
rect 6461 8577 6517 8633
rect 6545 8577 6601 8633
rect 6629 8577 6685 8633
rect 6713 8577 6769 8633
rect 6797 8577 6853 8633
rect 6881 8577 6937 8633
rect 6965 8577 7021 8633
rect 7048 8577 7104 8633
rect 7131 8577 7187 8633
rect 7214 8577 7270 8633
rect 7297 8577 7353 8633
rect 5621 8497 5677 8553
rect 5705 8497 5761 8553
rect 5789 8497 5845 8553
rect 5873 8497 5929 8553
rect 5957 8497 6013 8553
rect 6041 8497 6097 8553
rect 6125 8497 6181 8553
rect 6209 8497 6265 8553
rect 6293 8497 6349 8553
rect 6377 8497 6433 8553
rect 6461 8497 6517 8553
rect 6545 8497 6601 8553
rect 6629 8497 6685 8553
rect 6713 8497 6769 8553
rect 6797 8497 6853 8553
rect 6881 8497 6937 8553
rect 6965 8497 7021 8553
rect 7048 8497 7104 8553
rect 7131 8497 7187 8553
rect 7214 8497 7270 8553
rect 7297 8497 7353 8553
rect 5621 8417 5677 8473
rect 5705 8417 5761 8473
rect 5789 8417 5845 8473
rect 5873 8417 5929 8473
rect 5957 8417 6013 8473
rect 6041 8417 6097 8473
rect 6125 8417 6181 8473
rect 6209 8417 6265 8473
rect 6293 8417 6349 8473
rect 6377 8417 6433 8473
rect 6461 8417 6517 8473
rect 6545 8417 6601 8473
rect 6629 8417 6685 8473
rect 6713 8417 6769 8473
rect 6797 8417 6853 8473
rect 6881 8417 6937 8473
rect 6965 8417 7021 8473
rect 7048 8417 7104 8473
rect 7131 8417 7187 8473
rect 7214 8417 7270 8473
rect 7297 8417 7353 8473
rect 5621 8337 5677 8393
rect 5705 8337 5761 8393
rect 5789 8337 5845 8393
rect 5873 8337 5929 8393
rect 5957 8337 6013 8393
rect 6041 8337 6097 8393
rect 6125 8337 6181 8393
rect 6209 8337 6265 8393
rect 6293 8337 6349 8393
rect 6377 8337 6433 8393
rect 6461 8337 6517 8393
rect 6545 8337 6601 8393
rect 6629 8337 6685 8393
rect 6713 8337 6769 8393
rect 6797 8337 6853 8393
rect 6881 8337 6937 8393
rect 6965 8337 7021 8393
rect 7048 8337 7104 8393
rect 7131 8337 7187 8393
rect 7214 8337 7270 8393
rect 7297 8337 7353 8393
rect 5621 8257 5677 8313
rect 5705 8257 5761 8313
rect 5789 8257 5845 8313
rect 5873 8257 5929 8313
rect 5957 8257 6013 8313
rect 6041 8257 6097 8313
rect 6125 8257 6181 8313
rect 6209 8257 6265 8313
rect 6293 8257 6349 8313
rect 6377 8257 6433 8313
rect 6461 8257 6517 8313
rect 6545 8257 6601 8313
rect 6629 8257 6685 8313
rect 6713 8257 6769 8313
rect 6797 8257 6853 8313
rect 6881 8257 6937 8313
rect 6965 8257 7021 8313
rect 7048 8257 7104 8313
rect 7131 8257 7187 8313
rect 7214 8257 7270 8313
rect 7297 8257 7353 8313
rect 5621 8177 5677 8233
rect 5705 8177 5761 8233
rect 5789 8177 5845 8233
rect 5873 8177 5929 8233
rect 5957 8177 6013 8233
rect 6041 8177 6097 8233
rect 6125 8177 6181 8233
rect 6209 8177 6265 8233
rect 6293 8177 6349 8233
rect 6377 8177 6433 8233
rect 6461 8177 6517 8233
rect 6545 8177 6601 8233
rect 6629 8177 6685 8233
rect 6713 8177 6769 8233
rect 6797 8177 6853 8233
rect 6881 8177 6937 8233
rect 6965 8177 7021 8233
rect 7048 8177 7104 8233
rect 7131 8177 7187 8233
rect 7214 8177 7270 8233
rect 7297 8177 7353 8233
rect 5621 8097 5677 8153
rect 5705 8097 5761 8153
rect 5789 8097 5845 8153
rect 5873 8097 5929 8153
rect 5957 8097 6013 8153
rect 6041 8097 6097 8153
rect 6125 8097 6181 8153
rect 6209 8097 6265 8153
rect 6293 8097 6349 8153
rect 6377 8097 6433 8153
rect 6461 8097 6517 8153
rect 6545 8097 6601 8153
rect 6629 8097 6685 8153
rect 6713 8097 6769 8153
rect 6797 8097 6853 8153
rect 6881 8097 6937 8153
rect 6965 8097 7021 8153
rect 7048 8097 7104 8153
rect 7131 8097 7187 8153
rect 7214 8097 7270 8153
rect 7297 8097 7353 8153
rect 5621 8017 5677 8073
rect 5705 8017 5761 8073
rect 5789 8017 5845 8073
rect 5873 8017 5929 8073
rect 5957 8017 6013 8073
rect 6041 8017 6097 8073
rect 6125 8017 6181 8073
rect 6209 8017 6265 8073
rect 6293 8017 6349 8073
rect 6377 8017 6433 8073
rect 6461 8017 6517 8073
rect 6545 8017 6601 8073
rect 6629 8017 6685 8073
rect 6713 8017 6769 8073
rect 6797 8017 6853 8073
rect 6881 8017 6937 8073
rect 6965 8017 7021 8073
rect 7048 8017 7104 8073
rect 7131 8017 7187 8073
rect 7214 8017 7270 8073
rect 7297 8017 7353 8073
rect 5621 7937 5677 7993
rect 5705 7937 5761 7993
rect 5789 7937 5845 7993
rect 5873 7937 5929 7993
rect 5957 7937 6013 7993
rect 6041 7937 6097 7993
rect 6125 7937 6181 7993
rect 6209 7937 6265 7993
rect 6293 7937 6349 7993
rect 6377 7937 6433 7993
rect 6461 7937 6517 7993
rect 6545 7937 6601 7993
rect 6629 7937 6685 7993
rect 6713 7937 6769 7993
rect 6797 7937 6853 7993
rect 6881 7937 6937 7993
rect 6965 7937 7021 7993
rect 7048 7937 7104 7993
rect 7131 7937 7187 7993
rect 7214 7937 7270 7993
rect 7297 7937 7353 7993
rect 5621 7857 5677 7913
rect 5705 7857 5761 7913
rect 5789 7857 5845 7913
rect 5873 7857 5929 7913
rect 5957 7857 6013 7913
rect 6041 7857 6097 7913
rect 6125 7857 6181 7913
rect 6209 7857 6265 7913
rect 6293 7857 6349 7913
rect 6377 7857 6433 7913
rect 6461 7857 6517 7913
rect 6545 7857 6601 7913
rect 6629 7857 6685 7913
rect 6713 7857 6769 7913
rect 6797 7857 6853 7913
rect 6881 7857 6937 7913
rect 6965 7857 7021 7913
rect 7048 7857 7104 7913
rect 7131 7857 7187 7913
rect 7214 7857 7270 7913
rect 7297 7857 7353 7913
rect 5617 7690 5673 7692
rect 5698 7690 5754 7692
rect 5779 7690 5835 7692
rect 5860 7690 5916 7692
rect 5941 7690 5997 7692
rect 6022 7690 6078 7692
rect 6103 7690 6159 7692
rect 6184 7690 6240 7692
rect 6265 7690 6321 7692
rect 6346 7690 6402 7692
rect 6427 7690 6483 7692
rect 6508 7690 6564 7692
rect 6589 7690 6645 7692
rect 6669 7690 6725 7692
rect 6749 7690 6805 7692
rect 6829 7690 6885 7692
rect 6909 7690 6965 7692
rect 6989 7690 7045 7692
rect 7069 7690 7125 7692
rect 7149 7690 7205 7692
rect 7229 7690 7285 7692
rect 7309 7690 7365 7692
rect 5617 7638 5640 7690
rect 5640 7638 5652 7690
rect 5652 7638 5673 7690
rect 5698 7638 5704 7690
rect 5704 7638 5716 7690
rect 5716 7638 5754 7690
rect 5779 7638 5780 7690
rect 5780 7638 5832 7690
rect 5832 7638 5835 7690
rect 5860 7638 5896 7690
rect 5896 7638 5908 7690
rect 5908 7638 5916 7690
rect 5941 7638 5960 7690
rect 5960 7638 5972 7690
rect 5972 7638 5997 7690
rect 6022 7638 6024 7690
rect 6024 7638 6036 7690
rect 6036 7638 6078 7690
rect 6103 7638 6152 7690
rect 6152 7638 6159 7690
rect 6184 7638 6216 7690
rect 6216 7638 6228 7690
rect 6228 7638 6240 7690
rect 6265 7638 6280 7690
rect 6280 7638 6292 7690
rect 6292 7638 6321 7690
rect 6346 7638 6356 7690
rect 6356 7638 6402 7690
rect 6427 7638 6472 7690
rect 6472 7638 6483 7690
rect 6508 7638 6536 7690
rect 6536 7638 6548 7690
rect 6548 7638 6564 7690
rect 6589 7638 6600 7690
rect 6600 7638 6612 7690
rect 6612 7638 6645 7690
rect 6669 7638 6676 7690
rect 6676 7638 6725 7690
rect 6749 7638 6792 7690
rect 6792 7638 6804 7690
rect 6804 7638 6805 7690
rect 6829 7638 6856 7690
rect 6856 7638 6868 7690
rect 6868 7638 6885 7690
rect 6909 7638 6920 7690
rect 6920 7638 6932 7690
rect 6932 7638 6965 7690
rect 6989 7638 6996 7690
rect 6996 7638 7045 7690
rect 7069 7638 7112 7690
rect 7112 7638 7124 7690
rect 7124 7638 7125 7690
rect 7149 7638 7176 7690
rect 7176 7638 7188 7690
rect 7188 7638 7205 7690
rect 7229 7638 7240 7690
rect 7240 7638 7252 7690
rect 7252 7638 7285 7690
rect 7309 7638 7316 7690
rect 7316 7638 7365 7690
rect 5617 7636 5673 7638
rect 5698 7636 5754 7638
rect 5779 7636 5835 7638
rect 5860 7636 5916 7638
rect 5941 7636 5997 7638
rect 6022 7636 6078 7638
rect 6103 7636 6159 7638
rect 6184 7636 6240 7638
rect 6265 7636 6321 7638
rect 6346 7636 6402 7638
rect 6427 7636 6483 7638
rect 6508 7636 6564 7638
rect 6589 7636 6645 7638
rect 6669 7636 6725 7638
rect 6749 7636 6805 7638
rect 6829 7636 6885 7638
rect 6909 7636 6965 7638
rect 6989 7636 7045 7638
rect 7069 7636 7125 7638
rect 7149 7636 7205 7638
rect 7229 7636 7285 7638
rect 7309 7636 7365 7638
rect 5621 6859 5677 6915
rect 5705 6859 5761 6915
rect 5789 6859 5845 6915
rect 5873 6859 5929 6915
rect 5957 6859 6013 6915
rect 6041 6859 6097 6915
rect 6125 6859 6181 6915
rect 6209 6859 6265 6915
rect 6293 6859 6349 6915
rect 6377 6859 6433 6915
rect 6461 6859 6517 6915
rect 6545 6859 6601 6915
rect 6629 6859 6685 6915
rect 6713 6859 6769 6915
rect 6797 6859 6853 6915
rect 6881 6859 6937 6915
rect 6965 6859 7021 6915
rect 7048 6859 7104 6915
rect 7131 6859 7187 6915
rect 7214 6859 7270 6915
rect 7297 6859 7353 6915
rect 5621 6779 5677 6835
rect 5705 6779 5761 6835
rect 5789 6779 5845 6835
rect 5873 6779 5929 6835
rect 5957 6779 6013 6835
rect 6041 6779 6097 6835
rect 6125 6779 6181 6835
rect 6209 6779 6265 6835
rect 6293 6779 6349 6835
rect 6377 6779 6433 6835
rect 6461 6779 6517 6835
rect 6545 6779 6601 6835
rect 6629 6779 6685 6835
rect 6713 6779 6769 6835
rect 6797 6779 6853 6835
rect 6881 6779 6937 6835
rect 6965 6779 7021 6835
rect 7048 6779 7104 6835
rect 7131 6779 7187 6835
rect 7214 6779 7270 6835
rect 7297 6779 7353 6835
rect 5621 6699 5677 6755
rect 5705 6699 5761 6755
rect 5789 6699 5845 6755
rect 5873 6699 5929 6755
rect 5957 6699 6013 6755
rect 6041 6699 6097 6755
rect 6125 6699 6181 6755
rect 6209 6699 6265 6755
rect 6293 6699 6349 6755
rect 6377 6699 6433 6755
rect 6461 6699 6517 6755
rect 6545 6699 6601 6755
rect 6629 6699 6685 6755
rect 6713 6699 6769 6755
rect 6797 6699 6853 6755
rect 6881 6699 6937 6755
rect 6965 6699 7021 6755
rect 7048 6699 7104 6755
rect 7131 6699 7187 6755
rect 7214 6699 7270 6755
rect 7297 6699 7353 6755
rect 5621 6619 5677 6675
rect 5705 6619 5761 6675
rect 5789 6619 5845 6675
rect 5873 6619 5929 6675
rect 5957 6619 6013 6675
rect 6041 6619 6097 6675
rect 6125 6619 6181 6675
rect 6209 6619 6265 6675
rect 6293 6619 6349 6675
rect 6377 6619 6433 6675
rect 6461 6619 6517 6675
rect 6545 6619 6601 6675
rect 6629 6619 6685 6675
rect 6713 6619 6769 6675
rect 6797 6619 6853 6675
rect 6881 6619 6937 6675
rect 6965 6619 7021 6675
rect 7048 6619 7104 6675
rect 7131 6619 7187 6675
rect 7214 6619 7270 6675
rect 7297 6619 7353 6675
rect 5621 6539 5677 6595
rect 5705 6539 5761 6595
rect 5789 6539 5845 6595
rect 5873 6539 5929 6595
rect 5957 6539 6013 6595
rect 6041 6539 6097 6595
rect 6125 6539 6181 6595
rect 6209 6539 6265 6595
rect 6293 6539 6349 6595
rect 6377 6539 6433 6595
rect 6461 6539 6517 6595
rect 6545 6539 6601 6595
rect 6629 6539 6685 6595
rect 6713 6539 6769 6595
rect 6797 6539 6853 6595
rect 6881 6539 6937 6595
rect 6965 6539 7021 6595
rect 7048 6539 7104 6595
rect 7131 6539 7187 6595
rect 7214 6539 7270 6595
rect 7297 6539 7353 6595
rect 5621 6459 5677 6515
rect 5705 6459 5761 6515
rect 5789 6459 5845 6515
rect 5873 6459 5929 6515
rect 5957 6459 6013 6515
rect 6041 6459 6097 6515
rect 6125 6459 6181 6515
rect 6209 6459 6265 6515
rect 6293 6459 6349 6515
rect 6377 6459 6433 6515
rect 6461 6459 6517 6515
rect 6545 6459 6601 6515
rect 6629 6459 6685 6515
rect 6713 6459 6769 6515
rect 6797 6459 6853 6515
rect 6881 6459 6937 6515
rect 6965 6459 7021 6515
rect 7048 6459 7104 6515
rect 7131 6459 7187 6515
rect 7214 6459 7270 6515
rect 7297 6459 7353 6515
rect 5621 6379 5677 6435
rect 5705 6379 5761 6435
rect 5789 6379 5845 6435
rect 5873 6379 5929 6435
rect 5957 6379 6013 6435
rect 6041 6379 6097 6435
rect 6125 6379 6181 6435
rect 6209 6379 6265 6435
rect 6293 6379 6349 6435
rect 6377 6379 6433 6435
rect 6461 6379 6517 6435
rect 6545 6379 6601 6435
rect 6629 6379 6685 6435
rect 6713 6379 6769 6435
rect 6797 6379 6853 6435
rect 6881 6379 6937 6435
rect 6965 6379 7021 6435
rect 7048 6379 7104 6435
rect 7131 6379 7187 6435
rect 7214 6379 7270 6435
rect 7297 6379 7353 6435
rect 5621 6299 5677 6355
rect 5705 6299 5761 6355
rect 5789 6299 5845 6355
rect 5873 6299 5929 6355
rect 5957 6299 6013 6355
rect 6041 6299 6097 6355
rect 6125 6299 6181 6355
rect 6209 6299 6265 6355
rect 6293 6299 6349 6355
rect 6377 6299 6433 6355
rect 6461 6299 6517 6355
rect 6545 6299 6601 6355
rect 6629 6299 6685 6355
rect 6713 6299 6769 6355
rect 6797 6299 6853 6355
rect 6881 6299 6937 6355
rect 6965 6299 7021 6355
rect 7048 6299 7104 6355
rect 7131 6299 7187 6355
rect 7214 6299 7270 6355
rect 7297 6299 7353 6355
rect 5621 6219 5677 6275
rect 5705 6219 5761 6275
rect 5789 6219 5845 6275
rect 5873 6219 5929 6275
rect 5957 6219 6013 6275
rect 6041 6219 6097 6275
rect 6125 6219 6181 6275
rect 6209 6219 6265 6275
rect 6293 6219 6349 6275
rect 6377 6219 6433 6275
rect 6461 6219 6517 6275
rect 6545 6219 6601 6275
rect 6629 6219 6685 6275
rect 6713 6219 6769 6275
rect 6797 6219 6853 6275
rect 6881 6219 6937 6275
rect 6965 6219 7021 6275
rect 7048 6219 7104 6275
rect 7131 6219 7187 6275
rect 7214 6219 7270 6275
rect 7297 6219 7353 6275
rect 5621 6139 5677 6195
rect 5705 6139 5761 6195
rect 5789 6139 5845 6195
rect 5873 6139 5929 6195
rect 5957 6139 6013 6195
rect 6041 6139 6097 6195
rect 6125 6139 6181 6195
rect 6209 6139 6265 6195
rect 6293 6139 6349 6195
rect 6377 6139 6433 6195
rect 6461 6139 6517 6195
rect 6545 6139 6601 6195
rect 6629 6139 6685 6195
rect 6713 6139 6769 6195
rect 6797 6139 6853 6195
rect 6881 6139 6937 6195
rect 6965 6139 7021 6195
rect 7048 6139 7104 6195
rect 7131 6139 7187 6195
rect 7214 6139 7270 6195
rect 7297 6139 7353 6195
rect 5621 6059 5677 6115
rect 5705 6059 5761 6115
rect 5789 6059 5845 6115
rect 5873 6059 5929 6115
rect 5957 6059 6013 6115
rect 6041 6059 6097 6115
rect 6125 6059 6181 6115
rect 6209 6059 6265 6115
rect 6293 6059 6349 6115
rect 6377 6059 6433 6115
rect 6461 6059 6517 6115
rect 6545 6059 6601 6115
rect 6629 6059 6685 6115
rect 6713 6059 6769 6115
rect 6797 6059 6853 6115
rect 6881 6059 6937 6115
rect 6965 6059 7021 6115
rect 7048 6059 7104 6115
rect 7131 6059 7187 6115
rect 7214 6059 7270 6115
rect 7297 6059 7353 6115
rect 5617 5850 5673 5852
rect 5698 5850 5754 5852
rect 5779 5850 5835 5852
rect 5860 5850 5916 5852
rect 5941 5850 5997 5852
rect 6022 5850 6078 5852
rect 6103 5850 6159 5852
rect 6184 5850 6240 5852
rect 6265 5850 6321 5852
rect 6346 5850 6402 5852
rect 6427 5850 6483 5852
rect 6508 5850 6564 5852
rect 6589 5850 6645 5852
rect 6669 5850 6725 5852
rect 6749 5850 6805 5852
rect 6829 5850 6885 5852
rect 6909 5850 6965 5852
rect 6989 5850 7045 5852
rect 7069 5850 7125 5852
rect 7149 5850 7205 5852
rect 7229 5850 7285 5852
rect 7309 5850 7365 5852
rect 5617 5798 5640 5850
rect 5640 5798 5652 5850
rect 5652 5798 5673 5850
rect 5698 5798 5704 5850
rect 5704 5798 5716 5850
rect 5716 5798 5754 5850
rect 5779 5798 5780 5850
rect 5780 5798 5832 5850
rect 5832 5798 5835 5850
rect 5860 5798 5896 5850
rect 5896 5798 5908 5850
rect 5908 5798 5916 5850
rect 5941 5798 5960 5850
rect 5960 5798 5972 5850
rect 5972 5798 5997 5850
rect 6022 5798 6024 5850
rect 6024 5798 6036 5850
rect 6036 5798 6078 5850
rect 6103 5798 6152 5850
rect 6152 5798 6159 5850
rect 6184 5798 6216 5850
rect 6216 5798 6228 5850
rect 6228 5798 6240 5850
rect 6265 5798 6280 5850
rect 6280 5798 6292 5850
rect 6292 5798 6321 5850
rect 6346 5798 6356 5850
rect 6356 5798 6402 5850
rect 6427 5798 6472 5850
rect 6472 5798 6483 5850
rect 6508 5798 6536 5850
rect 6536 5798 6548 5850
rect 6548 5798 6564 5850
rect 6589 5798 6600 5850
rect 6600 5798 6612 5850
rect 6612 5798 6645 5850
rect 6669 5798 6676 5850
rect 6676 5798 6725 5850
rect 6749 5798 6792 5850
rect 6792 5798 6804 5850
rect 6804 5798 6805 5850
rect 6829 5798 6856 5850
rect 6856 5798 6868 5850
rect 6868 5798 6885 5850
rect 6909 5798 6920 5850
rect 6920 5798 6932 5850
rect 6932 5798 6965 5850
rect 6989 5798 6996 5850
rect 6996 5798 7045 5850
rect 7069 5798 7112 5850
rect 7112 5798 7124 5850
rect 7124 5798 7125 5850
rect 7149 5798 7176 5850
rect 7176 5798 7188 5850
rect 7188 5798 7205 5850
rect 7229 5798 7240 5850
rect 7240 5798 7252 5850
rect 7252 5798 7285 5850
rect 7309 5798 7316 5850
rect 7316 5798 7365 5850
rect 5617 5796 5673 5798
rect 5698 5796 5754 5798
rect 5779 5796 5835 5798
rect 5860 5796 5916 5798
rect 5941 5796 5997 5798
rect 6022 5796 6078 5798
rect 6103 5796 6159 5798
rect 6184 5796 6240 5798
rect 6265 5796 6321 5798
rect 6346 5796 6402 5798
rect 6427 5796 6483 5798
rect 6508 5796 6564 5798
rect 6589 5796 6645 5798
rect 6669 5796 6725 5798
rect 6749 5796 6805 5798
rect 6829 5796 6885 5798
rect 6909 5796 6965 5798
rect 6989 5796 7045 5798
rect 7069 5796 7125 5798
rect 7149 5796 7205 5798
rect 7229 5796 7285 5798
rect 7309 5796 7365 5798
rect 5623 4691 5652 4741
rect 5652 4691 5679 4741
rect 5623 4685 5679 4691
rect 5704 4691 5732 4741
rect 5732 4691 5760 4741
rect 5704 4685 5760 4691
rect 5785 4685 5841 4741
rect 5866 4691 5916 4741
rect 5916 4691 5922 4741
rect 5866 4685 5922 4691
rect 5947 4691 5996 4741
rect 5996 4691 6003 4741
rect 6027 4691 6048 4741
rect 6048 4691 6083 4741
rect 5947 4685 6003 4691
rect 6027 4685 6083 4691
rect 6107 4691 6128 4741
rect 6128 4691 6163 4741
rect 6107 4685 6163 4691
rect 6187 4685 6243 4741
rect 6267 4691 6312 4741
rect 6312 4691 6323 4741
rect 6267 4685 6323 4691
rect 6347 4691 6392 4741
rect 6392 4691 6403 4741
rect 6427 4691 6444 4741
rect 6444 4691 6483 4741
rect 6347 4685 6403 4691
rect 6427 4685 6483 4691
rect 6507 4691 6524 4741
rect 6524 4691 6563 4741
rect 6507 4685 6563 4691
rect 6587 4685 6643 4741
rect 6667 4691 6708 4741
rect 6708 4691 6723 4741
rect 6667 4685 6723 4691
rect 6747 4691 6788 4741
rect 6788 4691 6803 4741
rect 6827 4691 6840 4741
rect 6840 4691 6883 4741
rect 6747 4685 6803 4691
rect 6827 4685 6883 4691
rect 6907 4691 6920 4741
rect 6920 4691 6963 4741
rect 6907 4685 6963 4691
rect 6987 4685 7043 4741
rect 7067 4691 7104 4741
rect 7104 4691 7123 4741
rect 7067 4685 7123 4691
rect 7147 4691 7184 4741
rect 7184 4691 7203 4741
rect 7227 4691 7236 4741
rect 7236 4691 7283 4741
rect 7147 4685 7203 4691
rect 7227 4685 7283 4691
rect 7307 4691 7316 4741
rect 7316 4691 7363 4741
rect 7307 4685 7363 4691
rect 5623 4635 5679 4653
rect 5623 4597 5652 4635
rect 5652 4597 5679 4635
rect 5704 4635 5760 4653
rect 5704 4597 5732 4635
rect 5732 4597 5760 4635
rect 5785 4597 5841 4653
rect 5866 4635 5922 4653
rect 5866 4597 5916 4635
rect 5916 4597 5922 4635
rect 5947 4635 6003 4653
rect 6027 4635 6083 4653
rect 5947 4597 5996 4635
rect 5996 4597 6003 4635
rect 6027 4597 6048 4635
rect 6048 4597 6083 4635
rect 6107 4635 6163 4653
rect 6107 4597 6128 4635
rect 6128 4597 6163 4635
rect 6187 4597 6243 4653
rect 6267 4635 6323 4653
rect 6267 4597 6312 4635
rect 6312 4597 6323 4635
rect 6347 4635 6403 4653
rect 6427 4635 6483 4653
rect 6347 4597 6392 4635
rect 6392 4597 6403 4635
rect 6427 4597 6444 4635
rect 6444 4597 6483 4635
rect 6507 4635 6563 4653
rect 6507 4597 6524 4635
rect 6524 4597 6563 4635
rect 6587 4597 6643 4653
rect 6667 4635 6723 4653
rect 6667 4597 6708 4635
rect 6708 4597 6723 4635
rect 6747 4635 6803 4653
rect 6827 4635 6883 4653
rect 6747 4597 6788 4635
rect 6788 4597 6803 4635
rect 6827 4597 6840 4635
rect 6840 4597 6883 4635
rect 6907 4635 6963 4653
rect 6907 4597 6920 4635
rect 6920 4597 6963 4635
rect 6987 4597 7043 4653
rect 7067 4635 7123 4653
rect 7067 4597 7104 4635
rect 7104 4597 7123 4635
rect 7147 4635 7203 4653
rect 7227 4635 7283 4653
rect 7147 4597 7184 4635
rect 7184 4597 7203 4635
rect 7227 4597 7236 4635
rect 7236 4597 7283 4635
rect 7307 4635 7363 4653
rect 7307 4597 7316 4635
rect 7316 4597 7363 4635
rect 5623 4527 5679 4565
rect 5623 4509 5652 4527
rect 5652 4509 5679 4527
rect 5704 4527 5760 4565
rect 5704 4509 5732 4527
rect 5732 4509 5760 4527
rect 5785 4509 5841 4565
rect 5866 4527 5922 4565
rect 5866 4509 5916 4527
rect 5916 4509 5922 4527
rect 5947 4527 6003 4565
rect 6027 4527 6083 4565
rect 5947 4509 5996 4527
rect 5996 4509 6003 4527
rect 6027 4509 6048 4527
rect 6048 4509 6083 4527
rect 6107 4527 6163 4565
rect 6107 4509 6128 4527
rect 6128 4509 6163 4527
rect 6187 4509 6243 4565
rect 6267 4527 6323 4565
rect 6267 4509 6312 4527
rect 6312 4509 6323 4527
rect 6347 4527 6403 4565
rect 6427 4527 6483 4565
rect 6347 4509 6392 4527
rect 6392 4509 6403 4527
rect 6427 4509 6444 4527
rect 6444 4509 6483 4527
rect 6507 4527 6563 4565
rect 6507 4509 6524 4527
rect 6524 4509 6563 4527
rect 6587 4509 6643 4565
rect 6667 4527 6723 4565
rect 6667 4509 6708 4527
rect 6708 4509 6723 4527
rect 6747 4527 6803 4565
rect 6827 4527 6883 4565
rect 6747 4509 6788 4527
rect 6788 4509 6803 4527
rect 6827 4509 6840 4527
rect 6840 4509 6883 4527
rect 6907 4527 6963 4565
rect 6907 4509 6920 4527
rect 6920 4509 6963 4527
rect 6987 4509 7043 4565
rect 7067 4527 7123 4565
rect 7067 4509 7104 4527
rect 7104 4509 7123 4527
rect 7147 4527 7203 4565
rect 7227 4527 7283 4565
rect 7147 4509 7184 4527
rect 7184 4509 7203 4527
rect 7227 4509 7236 4527
rect 7236 4509 7283 4527
rect 7307 4527 7363 4565
rect 7307 4509 7316 4527
rect 7316 4509 7363 4527
rect 5623 4475 5652 4477
rect 5652 4475 5679 4477
rect 5623 4421 5679 4475
rect 5704 4475 5732 4477
rect 5732 4475 5760 4477
rect 5704 4421 5760 4475
rect 5785 4421 5841 4477
rect 5866 4475 5916 4477
rect 5916 4475 5922 4477
rect 5866 4421 5922 4475
rect 5947 4475 5996 4477
rect 5996 4475 6003 4477
rect 6027 4475 6048 4477
rect 6048 4475 6083 4477
rect 5947 4421 6003 4475
rect 6027 4421 6083 4475
rect 6107 4475 6128 4477
rect 6128 4475 6163 4477
rect 6107 4421 6163 4475
rect 6187 4421 6243 4477
rect 6267 4475 6312 4477
rect 6312 4475 6323 4477
rect 6267 4421 6323 4475
rect 6347 4475 6392 4477
rect 6392 4475 6403 4477
rect 6427 4475 6444 4477
rect 6444 4475 6483 4477
rect 6347 4421 6403 4475
rect 6427 4421 6483 4475
rect 6507 4475 6524 4477
rect 6524 4475 6563 4477
rect 6507 4421 6563 4475
rect 6587 4421 6643 4477
rect 6667 4475 6708 4477
rect 6708 4475 6723 4477
rect 6667 4421 6723 4475
rect 6747 4475 6788 4477
rect 6788 4475 6803 4477
rect 6827 4475 6840 4477
rect 6840 4475 6883 4477
rect 6747 4421 6803 4475
rect 6827 4421 6883 4475
rect 6907 4475 6920 4477
rect 6920 4475 6963 4477
rect 6907 4421 6963 4475
rect 6987 4421 7043 4477
rect 7067 4475 7104 4477
rect 7104 4475 7123 4477
rect 7067 4421 7123 4475
rect 7147 4475 7184 4477
rect 7184 4475 7203 4477
rect 7227 4475 7236 4477
rect 7236 4475 7283 4477
rect 7147 4421 7203 4475
rect 7227 4421 7283 4475
rect 7307 4475 7316 4477
rect 7316 4475 7363 4477
rect 7307 4421 7363 4475
rect 5623 4367 5652 4389
rect 5652 4367 5679 4389
rect 5623 4333 5679 4367
rect 5704 4367 5732 4389
rect 5732 4367 5760 4389
rect 5704 4333 5760 4367
rect 5785 4333 5841 4389
rect 5866 4367 5916 4389
rect 5916 4367 5922 4389
rect 5866 4333 5922 4367
rect 5947 4367 5996 4389
rect 5996 4367 6003 4389
rect 6027 4367 6048 4389
rect 6048 4367 6083 4389
rect 5947 4333 6003 4367
rect 6027 4333 6083 4367
rect 6107 4367 6128 4389
rect 6128 4367 6163 4389
rect 6107 4333 6163 4367
rect 6187 4333 6243 4389
rect 6267 4367 6312 4389
rect 6312 4367 6323 4389
rect 6267 4333 6323 4367
rect 6347 4367 6392 4389
rect 6392 4367 6403 4389
rect 6427 4367 6444 4389
rect 6444 4367 6483 4389
rect 6347 4333 6403 4367
rect 6427 4333 6483 4367
rect 6507 4367 6524 4389
rect 6524 4367 6563 4389
rect 6507 4333 6563 4367
rect 6587 4333 6643 4389
rect 6667 4367 6708 4389
rect 6708 4367 6723 4389
rect 6667 4333 6723 4367
rect 6747 4367 6788 4389
rect 6788 4367 6803 4389
rect 6827 4367 6840 4389
rect 6840 4367 6883 4389
rect 6747 4333 6803 4367
rect 6827 4333 6883 4367
rect 6907 4367 6920 4389
rect 6920 4367 6963 4389
rect 6907 4333 6963 4367
rect 6987 4333 7043 4389
rect 7067 4367 7104 4389
rect 7104 4367 7123 4389
rect 7067 4333 7123 4367
rect 7147 4367 7184 4389
rect 7184 4367 7203 4389
rect 7227 4367 7236 4389
rect 7236 4367 7283 4389
rect 7147 4333 7203 4367
rect 7227 4333 7283 4367
rect 7307 4367 7316 4389
rect 7316 4367 7363 4389
rect 7307 4333 7363 4367
rect 5623 4259 5652 4301
rect 5652 4259 5679 4301
rect 5623 4245 5679 4259
rect 5704 4259 5732 4301
rect 5732 4259 5760 4301
rect 5704 4245 5760 4259
rect 5785 4245 5841 4301
rect 5866 4259 5916 4301
rect 5916 4259 5922 4301
rect 5866 4245 5922 4259
rect 5947 4259 5996 4301
rect 5996 4259 6003 4301
rect 6027 4259 6048 4301
rect 6048 4259 6083 4301
rect 5947 4245 6003 4259
rect 6027 4245 6083 4259
rect 6107 4259 6128 4301
rect 6128 4259 6163 4301
rect 6107 4245 6163 4259
rect 6187 4245 6243 4301
rect 6267 4259 6312 4301
rect 6312 4259 6323 4301
rect 6267 4245 6323 4259
rect 6347 4259 6392 4301
rect 6392 4259 6403 4301
rect 6427 4259 6444 4301
rect 6444 4259 6483 4301
rect 6347 4245 6403 4259
rect 6427 4245 6483 4259
rect 6507 4259 6524 4301
rect 6524 4259 6563 4301
rect 6507 4245 6563 4259
rect 6587 4245 6643 4301
rect 6667 4259 6708 4301
rect 6708 4259 6723 4301
rect 6667 4245 6723 4259
rect 6747 4259 6788 4301
rect 6788 4259 6803 4301
rect 6827 4259 6840 4301
rect 6840 4259 6883 4301
rect 6747 4245 6803 4259
rect 6827 4245 6883 4259
rect 6907 4259 6920 4301
rect 6920 4259 6963 4301
rect 6907 4245 6963 4259
rect 6987 4245 7043 4301
rect 7067 4259 7104 4301
rect 7104 4259 7123 4301
rect 7067 4245 7123 4259
rect 7147 4259 7184 4301
rect 7184 4259 7203 4301
rect 7227 4259 7236 4301
rect 7236 4259 7283 4301
rect 7147 4245 7203 4259
rect 7227 4245 7283 4259
rect 7307 4259 7316 4301
rect 7316 4259 7363 4301
rect 7307 4245 7363 4259
rect 5623 4203 5679 4213
rect 5623 4157 5652 4203
rect 5652 4157 5679 4203
rect 5704 4203 5760 4213
rect 5704 4157 5732 4203
rect 5732 4157 5760 4203
rect 5785 4157 5841 4213
rect 5866 4203 5922 4213
rect 5866 4157 5916 4203
rect 5916 4157 5922 4203
rect 5947 4203 6003 4213
rect 6027 4203 6083 4213
rect 5947 4157 5996 4203
rect 5996 4157 6003 4203
rect 6027 4157 6048 4203
rect 6048 4157 6083 4203
rect 6107 4203 6163 4213
rect 6107 4157 6128 4203
rect 6128 4157 6163 4203
rect 6187 4157 6243 4213
rect 6267 4203 6323 4213
rect 6267 4157 6312 4203
rect 6312 4157 6323 4203
rect 6347 4203 6403 4213
rect 6427 4203 6483 4213
rect 6347 4157 6392 4203
rect 6392 4157 6403 4203
rect 6427 4157 6444 4203
rect 6444 4157 6483 4203
rect 6507 4203 6563 4213
rect 6507 4157 6524 4203
rect 6524 4157 6563 4203
rect 6587 4157 6643 4213
rect 6667 4203 6723 4213
rect 6667 4157 6708 4203
rect 6708 4157 6723 4203
rect 6747 4203 6803 4213
rect 6827 4203 6883 4213
rect 6747 4157 6788 4203
rect 6788 4157 6803 4203
rect 6827 4157 6840 4203
rect 6840 4157 6883 4203
rect 6907 4203 6963 4213
rect 6907 4157 6920 4203
rect 6920 4157 6963 4203
rect 6987 4157 7043 4213
rect 7067 4203 7123 4213
rect 7067 4157 7104 4203
rect 7104 4157 7123 4203
rect 7147 4203 7203 4213
rect 7227 4203 7283 4213
rect 7147 4157 7184 4203
rect 7184 4157 7203 4203
rect 7227 4157 7236 4203
rect 7236 4157 7283 4203
rect 7307 4203 7363 4213
rect 7307 4157 7316 4203
rect 7316 4157 7363 4203
rect 5617 3897 5661 3918
rect 5661 3897 5673 3918
rect 5617 3883 5673 3897
rect 5617 3862 5661 3883
rect 5661 3862 5673 3883
rect 5698 3897 5744 3918
rect 5744 3897 5754 3918
rect 5779 3897 5796 3918
rect 5796 3897 5835 3918
rect 5698 3883 5754 3897
rect 5779 3883 5835 3897
rect 5698 3862 5744 3883
rect 5744 3862 5754 3883
rect 5779 3862 5796 3883
rect 5796 3862 5835 3883
rect 5860 3897 5879 3918
rect 5879 3897 5916 3918
rect 5860 3883 5916 3897
rect 5860 3862 5879 3883
rect 5879 3862 5916 3883
rect 5941 3862 5997 3918
rect 6022 3897 6066 3918
rect 6066 3897 6078 3918
rect 6022 3883 6078 3897
rect 6022 3862 6066 3883
rect 6066 3862 6078 3883
rect 6103 3897 6149 3918
rect 6149 3897 6159 3918
rect 6184 3897 6201 3918
rect 6201 3897 6240 3918
rect 6103 3883 6159 3897
rect 6184 3883 6240 3897
rect 6103 3862 6149 3883
rect 6149 3862 6159 3883
rect 6184 3862 6201 3883
rect 6201 3862 6240 3883
rect 6265 3897 6284 3918
rect 6284 3897 6321 3918
rect 6265 3883 6321 3897
rect 6265 3862 6284 3883
rect 6284 3862 6321 3883
rect 6346 3862 6402 3918
rect 6427 3897 6471 3918
rect 6471 3897 6483 3918
rect 6427 3883 6483 3897
rect 6427 3862 6471 3883
rect 6471 3862 6483 3883
rect 6508 3897 6553 3918
rect 6553 3897 6564 3918
rect 6589 3897 6605 3918
rect 6605 3897 6645 3918
rect 6508 3883 6564 3897
rect 6589 3883 6645 3897
rect 6508 3862 6553 3883
rect 6553 3862 6564 3883
rect 6589 3862 6605 3883
rect 6605 3862 6645 3883
rect 6669 3897 6687 3918
rect 6687 3897 6725 3918
rect 6669 3883 6725 3897
rect 6669 3862 6687 3883
rect 6687 3862 6725 3883
rect 6749 3862 6805 3918
rect 6829 3897 6873 3918
rect 6873 3897 6885 3918
rect 6829 3883 6885 3897
rect 6829 3862 6873 3883
rect 6873 3862 6885 3883
rect 6909 3897 6955 3918
rect 6955 3897 6965 3918
rect 6989 3897 7007 3918
rect 7007 3897 7045 3918
rect 6909 3883 6965 3897
rect 6989 3883 7045 3897
rect 6909 3862 6955 3883
rect 6955 3862 6965 3883
rect 6989 3862 7007 3883
rect 7007 3862 7045 3883
rect 7069 3897 7089 3918
rect 7089 3897 7125 3918
rect 7069 3883 7125 3897
rect 7069 3862 7089 3883
rect 7089 3862 7125 3883
rect 7149 3862 7205 3918
rect 7229 3897 7275 3918
rect 7275 3897 7285 3918
rect 7229 3883 7285 3897
rect 7229 3862 7275 3883
rect 7275 3862 7285 3883
rect 7309 3862 7365 3918
rect 5617 3005 5651 3057
rect 5651 3005 5664 3057
rect 5664 3005 5673 3057
rect 5698 3005 5716 3057
rect 5716 3005 5729 3057
rect 5729 3005 5754 3057
rect 5779 3005 5781 3057
rect 5781 3005 5794 3057
rect 5794 3005 5835 3057
rect 5860 3005 5911 3057
rect 5911 3005 5916 3057
rect 5941 3005 5976 3057
rect 5976 3005 5989 3057
rect 5989 3005 5997 3057
rect 6022 3005 6041 3057
rect 6041 3005 6054 3057
rect 6054 3005 6078 3057
rect 6103 3005 6106 3057
rect 6106 3005 6119 3057
rect 6119 3005 6159 3057
rect 6184 3005 6236 3057
rect 6236 3005 6240 3057
rect 6265 3005 6301 3057
rect 6301 3005 6314 3057
rect 6314 3005 6321 3057
rect 6346 3005 6366 3057
rect 6366 3005 6379 3057
rect 6379 3005 6402 3057
rect 6427 3005 6431 3057
rect 6431 3005 6444 3057
rect 6444 3005 6483 3057
rect 6508 3005 6509 3057
rect 6509 3005 6561 3057
rect 6561 3005 6564 3057
rect 6589 3005 6626 3057
rect 6626 3005 6639 3057
rect 6639 3005 6645 3057
rect 6670 3005 6691 3057
rect 6691 3005 6704 3057
rect 6704 3005 6726 3057
rect 6751 3005 6756 3057
rect 6756 3005 6769 3057
rect 6769 3005 6807 3057
rect 6832 3005 6834 3057
rect 6834 3005 6886 3057
rect 6886 3005 6888 3057
rect 6913 3005 6951 3057
rect 6951 3005 6964 3057
rect 6964 3005 6969 3057
rect 6994 3005 7016 3057
rect 7016 3005 7029 3057
rect 7029 3005 7050 3057
rect 7075 3005 7081 3057
rect 7081 3005 7094 3057
rect 7094 3005 7131 3057
rect 7156 3005 7159 3057
rect 7159 3005 7211 3057
rect 7211 3005 7212 3057
rect 7237 3005 7276 3057
rect 7276 3005 7289 3057
rect 7289 3005 7293 3057
rect 7317 3005 7341 3057
rect 7341 3005 7354 3057
rect 7354 3005 7373 3057
rect 7397 3005 7406 3057
rect 7406 3005 7419 3057
rect 7419 3005 7453 3057
rect 7477 3005 7484 3057
rect 7484 3005 7533 3057
rect 5617 3001 5673 3005
rect 5698 3001 5754 3005
rect 5779 3001 5835 3005
rect 5860 3001 5916 3005
rect 5941 3001 5997 3005
rect 6022 3001 6078 3005
rect 6103 3001 6159 3005
rect 6184 3001 6240 3005
rect 6265 3001 6321 3005
rect 6346 3001 6402 3005
rect 6427 3001 6483 3005
rect 6508 3001 6564 3005
rect 6589 3001 6645 3005
rect 6670 3001 6726 3005
rect 6751 3001 6807 3005
rect 6832 3001 6888 3005
rect 6913 3001 6969 3005
rect 6994 3001 7050 3005
rect 7075 3001 7131 3005
rect 7156 3001 7212 3005
rect 7237 3001 7293 3005
rect 7317 3001 7373 3005
rect 7397 3001 7453 3005
rect 7477 3001 7533 3005
rect 5617 2937 5651 2967
rect 5651 2937 5664 2967
rect 5664 2937 5673 2967
rect 5698 2937 5716 2967
rect 5716 2937 5729 2967
rect 5729 2937 5754 2967
rect 5779 2937 5781 2967
rect 5781 2937 5794 2967
rect 5794 2937 5835 2967
rect 5860 2937 5911 2967
rect 5911 2937 5916 2967
rect 5941 2937 5976 2967
rect 5976 2937 5989 2967
rect 5989 2937 5997 2967
rect 6022 2937 6041 2967
rect 6041 2937 6054 2967
rect 6054 2937 6078 2967
rect 6103 2937 6106 2967
rect 6106 2937 6119 2967
rect 6119 2937 6159 2967
rect 6184 2937 6236 2967
rect 6236 2937 6240 2967
rect 6265 2937 6301 2967
rect 6301 2937 6314 2967
rect 6314 2937 6321 2967
rect 6346 2937 6366 2967
rect 6366 2937 6379 2967
rect 6379 2937 6402 2967
rect 6427 2937 6431 2967
rect 6431 2937 6444 2967
rect 6444 2937 6483 2967
rect 6508 2937 6509 2967
rect 6509 2937 6561 2967
rect 6561 2937 6564 2967
rect 6589 2937 6626 2967
rect 6626 2937 6639 2967
rect 6639 2937 6645 2967
rect 6670 2937 6691 2967
rect 6691 2937 6704 2967
rect 6704 2937 6726 2967
rect 6751 2937 6756 2967
rect 6756 2937 6769 2967
rect 6769 2937 6807 2967
rect 6832 2937 6834 2967
rect 6834 2937 6886 2967
rect 6886 2937 6888 2967
rect 6913 2937 6951 2967
rect 6951 2937 6964 2967
rect 6964 2937 6969 2967
rect 6994 2937 7016 2967
rect 7016 2937 7029 2967
rect 7029 2937 7050 2967
rect 7075 2937 7081 2967
rect 7081 2937 7094 2967
rect 7094 2937 7131 2967
rect 7156 2937 7159 2967
rect 7159 2937 7211 2967
rect 7211 2937 7212 2967
rect 7237 2937 7276 2967
rect 7276 2937 7289 2967
rect 7289 2937 7293 2967
rect 7317 2937 7341 2967
rect 7341 2937 7354 2967
rect 7354 2937 7373 2967
rect 7397 2937 7406 2967
rect 7406 2937 7419 2967
rect 7419 2937 7453 2967
rect 7477 2937 7484 2967
rect 7484 2937 7533 2967
rect 5617 2921 5673 2937
rect 5698 2921 5754 2937
rect 5779 2921 5835 2937
rect 5860 2921 5916 2937
rect 5941 2921 5997 2937
rect 6022 2921 6078 2937
rect 6103 2921 6159 2937
rect 6184 2921 6240 2937
rect 6265 2921 6321 2937
rect 6346 2921 6402 2937
rect 6427 2921 6483 2937
rect 6508 2921 6564 2937
rect 6589 2921 6645 2937
rect 6670 2921 6726 2937
rect 6751 2921 6807 2937
rect 6832 2921 6888 2937
rect 6913 2921 6969 2937
rect 6994 2921 7050 2937
rect 7075 2921 7131 2937
rect 7156 2921 7212 2937
rect 7237 2921 7293 2937
rect 7317 2921 7373 2937
rect 7397 2921 7453 2937
rect 7477 2921 7533 2937
rect 5617 2911 5651 2921
rect 5651 2911 5664 2921
rect 5664 2911 5673 2921
rect 5698 2911 5716 2921
rect 5716 2911 5729 2921
rect 5729 2911 5754 2921
rect 5779 2911 5781 2921
rect 5781 2911 5794 2921
rect 5794 2911 5835 2921
rect 5617 2869 5651 2877
rect 5651 2869 5664 2877
rect 5664 2869 5673 2877
rect 5698 2869 5716 2877
rect 5716 2869 5729 2877
rect 5729 2869 5754 2877
rect 5779 2869 5781 2877
rect 5781 2869 5794 2877
rect 5794 2869 5835 2877
rect 5860 2911 5911 2921
rect 5911 2911 5916 2921
rect 5941 2911 5976 2921
rect 5976 2911 5989 2921
rect 5989 2911 5997 2921
rect 6022 2911 6041 2921
rect 6041 2911 6054 2921
rect 6054 2911 6078 2921
rect 6103 2911 6106 2921
rect 6106 2911 6119 2921
rect 6119 2911 6159 2921
rect 5860 2869 5911 2877
rect 5911 2869 5916 2877
rect 5941 2869 5976 2877
rect 5976 2869 5989 2877
rect 5989 2869 5997 2877
rect 6022 2869 6041 2877
rect 6041 2869 6054 2877
rect 6054 2869 6078 2877
rect 6103 2869 6106 2877
rect 6106 2869 6119 2877
rect 6119 2869 6159 2877
rect 6184 2911 6236 2921
rect 6236 2911 6240 2921
rect 6265 2911 6301 2921
rect 6301 2911 6314 2921
rect 6314 2911 6321 2921
rect 6346 2911 6366 2921
rect 6366 2911 6379 2921
rect 6379 2911 6402 2921
rect 6427 2911 6431 2921
rect 6431 2911 6444 2921
rect 6444 2911 6483 2921
rect 6508 2911 6509 2921
rect 6509 2911 6561 2921
rect 6561 2911 6564 2921
rect 6589 2911 6626 2921
rect 6626 2911 6639 2921
rect 6639 2911 6645 2921
rect 6670 2911 6691 2921
rect 6691 2911 6704 2921
rect 6704 2911 6726 2921
rect 6751 2911 6756 2921
rect 6756 2911 6769 2921
rect 6769 2911 6807 2921
rect 6832 2911 6834 2921
rect 6834 2911 6886 2921
rect 6886 2911 6888 2921
rect 6913 2911 6951 2921
rect 6951 2911 6964 2921
rect 6964 2911 6969 2921
rect 6994 2911 7016 2921
rect 7016 2911 7029 2921
rect 7029 2911 7050 2921
rect 7075 2911 7081 2921
rect 7081 2911 7094 2921
rect 7094 2911 7131 2921
rect 7156 2911 7159 2921
rect 7159 2911 7211 2921
rect 7211 2911 7212 2921
rect 7237 2911 7276 2921
rect 7276 2911 7289 2921
rect 7289 2911 7293 2921
rect 7317 2911 7341 2921
rect 7341 2911 7354 2921
rect 7354 2911 7373 2921
rect 7397 2911 7406 2921
rect 7406 2911 7419 2921
rect 7419 2911 7453 2921
rect 7477 2911 7484 2921
rect 7484 2911 7533 2921
rect 6184 2869 6236 2877
rect 6236 2869 6240 2877
rect 6265 2869 6301 2877
rect 6301 2869 6314 2877
rect 6314 2869 6321 2877
rect 6346 2869 6366 2877
rect 6366 2869 6379 2877
rect 6379 2869 6402 2877
rect 6427 2869 6431 2877
rect 6431 2869 6444 2877
rect 6444 2869 6483 2877
rect 6508 2869 6509 2877
rect 6509 2869 6561 2877
rect 6561 2869 6564 2877
rect 6589 2869 6626 2877
rect 6626 2869 6639 2877
rect 6639 2869 6645 2877
rect 6670 2869 6691 2877
rect 6691 2869 6704 2877
rect 6704 2869 6726 2877
rect 6751 2869 6756 2877
rect 6756 2869 6769 2877
rect 6769 2869 6807 2877
rect 6832 2869 6834 2877
rect 6834 2869 6886 2877
rect 6886 2869 6888 2877
rect 6913 2869 6951 2877
rect 6951 2869 6964 2877
rect 6964 2869 6969 2877
rect 6994 2869 7016 2877
rect 7016 2869 7029 2877
rect 7029 2869 7050 2877
rect 7075 2869 7081 2877
rect 7081 2869 7094 2877
rect 7094 2869 7131 2877
rect 7156 2869 7159 2877
rect 7159 2869 7211 2877
rect 7211 2869 7212 2877
rect 7237 2869 7276 2877
rect 7276 2869 7289 2877
rect 7289 2869 7293 2877
rect 7317 2869 7341 2877
rect 7341 2869 7354 2877
rect 7354 2869 7373 2877
rect 7397 2869 7406 2877
rect 7406 2869 7419 2877
rect 7419 2869 7453 2877
rect 7477 2869 7484 2877
rect 7484 2869 7533 2877
rect 5617 2853 5673 2869
rect 5698 2853 5754 2869
rect 5779 2853 5835 2869
rect 5860 2853 5916 2869
rect 5941 2853 5997 2869
rect 6022 2853 6078 2869
rect 6103 2853 6159 2869
rect 6184 2853 6240 2869
rect 6265 2853 6321 2869
rect 6346 2853 6402 2869
rect 6427 2853 6483 2869
rect 6508 2853 6564 2869
rect 6589 2853 6645 2869
rect 6670 2853 6726 2869
rect 6751 2853 6807 2869
rect 6832 2853 6888 2869
rect 6913 2853 6969 2869
rect 6994 2853 7050 2869
rect 7075 2853 7131 2869
rect 7156 2853 7212 2869
rect 7237 2853 7293 2869
rect 7317 2853 7373 2869
rect 7397 2853 7453 2869
rect 7477 2853 7533 2869
rect 5617 2821 5651 2853
rect 5651 2821 5664 2853
rect 5664 2821 5673 2853
rect 5698 2821 5716 2853
rect 5716 2821 5729 2853
rect 5729 2821 5754 2853
rect 5779 2821 5781 2853
rect 5781 2821 5794 2853
rect 5794 2821 5835 2853
rect 5860 2821 5911 2853
rect 5911 2821 5916 2853
rect 5941 2821 5976 2853
rect 5976 2821 5989 2853
rect 5989 2821 5997 2853
rect 6022 2821 6041 2853
rect 6041 2821 6054 2853
rect 6054 2821 6078 2853
rect 6103 2821 6106 2853
rect 6106 2821 6119 2853
rect 6119 2821 6159 2853
rect 6184 2821 6236 2853
rect 6236 2821 6240 2853
rect 6265 2821 6301 2853
rect 6301 2821 6314 2853
rect 6314 2821 6321 2853
rect 6346 2821 6366 2853
rect 6366 2821 6379 2853
rect 6379 2821 6402 2853
rect 6427 2821 6431 2853
rect 6431 2821 6444 2853
rect 6444 2821 6483 2853
rect 6508 2821 6509 2853
rect 6509 2821 6561 2853
rect 6561 2821 6564 2853
rect 6589 2821 6626 2853
rect 6626 2821 6639 2853
rect 6639 2821 6645 2853
rect 6670 2821 6691 2853
rect 6691 2821 6704 2853
rect 6704 2821 6726 2853
rect 6751 2821 6756 2853
rect 6756 2821 6769 2853
rect 6769 2821 6807 2853
rect 6832 2821 6834 2853
rect 6834 2821 6886 2853
rect 6886 2821 6888 2853
rect 6913 2821 6951 2853
rect 6951 2821 6964 2853
rect 6964 2821 6969 2853
rect 6994 2821 7016 2853
rect 7016 2821 7029 2853
rect 7029 2821 7050 2853
rect 7075 2821 7081 2853
rect 7081 2821 7094 2853
rect 7094 2821 7131 2853
rect 7156 2821 7159 2853
rect 7159 2821 7211 2853
rect 7211 2821 7212 2853
rect 7237 2821 7276 2853
rect 7276 2821 7289 2853
rect 7289 2821 7293 2853
rect 7317 2821 7341 2853
rect 7341 2821 7354 2853
rect 7354 2821 7373 2853
rect 7397 2821 7406 2853
rect 7406 2821 7419 2853
rect 7419 2821 7453 2853
rect 7477 2821 7484 2853
rect 7484 2821 7533 2853
rect 5617 2785 5673 2787
rect 5698 2785 5754 2787
rect 5779 2785 5835 2787
rect 5860 2785 5916 2787
rect 5941 2785 5997 2787
rect 6022 2785 6078 2787
rect 6103 2785 6159 2787
rect 6184 2785 6240 2787
rect 6265 2785 6321 2787
rect 6346 2785 6402 2787
rect 6427 2785 6483 2787
rect 6508 2785 6564 2787
rect 6589 2785 6645 2787
rect 6670 2785 6726 2787
rect 6751 2785 6807 2787
rect 6832 2785 6888 2787
rect 6913 2785 6969 2787
rect 6994 2785 7050 2787
rect 7075 2785 7131 2787
rect 7156 2785 7212 2787
rect 7237 2785 7293 2787
rect 7317 2785 7373 2787
rect 7397 2785 7453 2787
rect 7477 2785 7533 2787
rect 5617 2733 5651 2785
rect 5651 2733 5664 2785
rect 5664 2733 5673 2785
rect 5698 2733 5716 2785
rect 5716 2733 5729 2785
rect 5729 2733 5754 2785
rect 5779 2733 5781 2785
rect 5781 2733 5794 2785
rect 5794 2733 5835 2785
rect 5860 2733 5911 2785
rect 5911 2733 5916 2785
rect 5941 2733 5976 2785
rect 5976 2733 5989 2785
rect 5989 2733 5997 2785
rect 6022 2733 6041 2785
rect 6041 2733 6054 2785
rect 6054 2733 6078 2785
rect 6103 2733 6106 2785
rect 6106 2733 6119 2785
rect 6119 2733 6159 2785
rect 6184 2733 6236 2785
rect 6236 2733 6240 2785
rect 6265 2733 6301 2785
rect 6301 2733 6314 2785
rect 6314 2733 6321 2785
rect 6346 2733 6366 2785
rect 6366 2733 6379 2785
rect 6379 2733 6402 2785
rect 6427 2733 6431 2785
rect 6431 2733 6444 2785
rect 6444 2733 6483 2785
rect 6508 2733 6509 2785
rect 6509 2733 6561 2785
rect 6561 2733 6564 2785
rect 6589 2733 6626 2785
rect 6626 2733 6639 2785
rect 6639 2733 6645 2785
rect 6670 2733 6691 2785
rect 6691 2733 6704 2785
rect 6704 2733 6726 2785
rect 6751 2733 6756 2785
rect 6756 2733 6769 2785
rect 6769 2733 6807 2785
rect 6832 2733 6834 2785
rect 6834 2733 6886 2785
rect 6886 2733 6888 2785
rect 6913 2733 6951 2785
rect 6951 2733 6964 2785
rect 6964 2733 6969 2785
rect 6994 2733 7016 2785
rect 7016 2733 7029 2785
rect 7029 2733 7050 2785
rect 7075 2733 7081 2785
rect 7081 2733 7094 2785
rect 7094 2733 7131 2785
rect 7156 2733 7159 2785
rect 7159 2733 7211 2785
rect 7211 2733 7212 2785
rect 7237 2733 7276 2785
rect 7276 2733 7289 2785
rect 7289 2733 7293 2785
rect 7317 2733 7341 2785
rect 7341 2733 7354 2785
rect 7354 2733 7373 2785
rect 7397 2733 7406 2785
rect 7406 2733 7419 2785
rect 7419 2733 7453 2785
rect 7477 2733 7484 2785
rect 7484 2733 7533 2785
rect 5617 2731 5673 2733
rect 5698 2731 5754 2733
rect 5779 2731 5835 2733
rect 5860 2731 5916 2733
rect 5941 2731 5997 2733
rect 6022 2731 6078 2733
rect 6103 2731 6159 2733
rect 6184 2731 6240 2733
rect 6265 2731 6321 2733
rect 6346 2731 6402 2733
rect 6427 2731 6483 2733
rect 6508 2731 6564 2733
rect 6589 2731 6645 2733
rect 6670 2731 6726 2733
rect 6751 2731 6807 2733
rect 6832 2731 6888 2733
rect 6913 2731 6969 2733
rect 6994 2731 7050 2733
rect 7075 2731 7131 2733
rect 7156 2731 7212 2733
rect 7237 2731 7293 2733
rect 7317 2731 7373 2733
rect 7397 2731 7453 2733
rect 7477 2731 7533 2733
rect 5617 2665 5651 2697
rect 5651 2665 5664 2697
rect 5664 2665 5673 2697
rect 5698 2665 5716 2697
rect 5716 2665 5729 2697
rect 5729 2665 5754 2697
rect 5779 2665 5781 2697
rect 5781 2665 5794 2697
rect 5794 2665 5835 2697
rect 5860 2665 5911 2697
rect 5911 2665 5916 2697
rect 5941 2665 5976 2697
rect 5976 2665 5989 2697
rect 5989 2665 5997 2697
rect 6022 2665 6041 2697
rect 6041 2665 6054 2697
rect 6054 2665 6078 2697
rect 6103 2665 6106 2697
rect 6106 2665 6119 2697
rect 6119 2665 6159 2697
rect 6184 2665 6236 2697
rect 6236 2665 6240 2697
rect 6265 2665 6301 2697
rect 6301 2665 6314 2697
rect 6314 2665 6321 2697
rect 6346 2665 6366 2697
rect 6366 2665 6379 2697
rect 6379 2665 6402 2697
rect 6427 2665 6431 2697
rect 6431 2665 6444 2697
rect 6444 2665 6483 2697
rect 6508 2665 6509 2697
rect 6509 2665 6561 2697
rect 6561 2665 6564 2697
rect 6589 2665 6626 2697
rect 6626 2665 6639 2697
rect 6639 2665 6645 2697
rect 6670 2665 6691 2697
rect 6691 2665 6704 2697
rect 6704 2665 6726 2697
rect 6751 2665 6756 2697
rect 6756 2665 6769 2697
rect 6769 2665 6807 2697
rect 6832 2665 6834 2697
rect 6834 2665 6886 2697
rect 6886 2665 6888 2697
rect 6913 2665 6951 2697
rect 6951 2665 6964 2697
rect 6964 2665 6969 2697
rect 6994 2665 7016 2697
rect 7016 2665 7029 2697
rect 7029 2665 7050 2697
rect 7075 2665 7081 2697
rect 7081 2665 7094 2697
rect 7094 2665 7131 2697
rect 7156 2665 7159 2697
rect 7159 2665 7211 2697
rect 7211 2665 7212 2697
rect 7237 2665 7276 2697
rect 7276 2665 7289 2697
rect 7289 2665 7293 2697
rect 7317 2665 7341 2697
rect 7341 2665 7354 2697
rect 7354 2665 7373 2697
rect 7397 2665 7406 2697
rect 7406 2665 7419 2697
rect 7419 2665 7453 2697
rect 7477 2665 7484 2697
rect 7484 2665 7533 2697
rect 5617 2649 5673 2665
rect 5698 2649 5754 2665
rect 5779 2649 5835 2665
rect 5860 2649 5916 2665
rect 5941 2649 5997 2665
rect 6022 2649 6078 2665
rect 6103 2649 6159 2665
rect 6184 2649 6240 2665
rect 6265 2649 6321 2665
rect 6346 2649 6402 2665
rect 6427 2649 6483 2665
rect 6508 2649 6564 2665
rect 6589 2649 6645 2665
rect 6670 2649 6726 2665
rect 6751 2649 6807 2665
rect 6832 2649 6888 2665
rect 6913 2649 6969 2665
rect 6994 2649 7050 2665
rect 7075 2649 7131 2665
rect 7156 2649 7212 2665
rect 7237 2649 7293 2665
rect 7317 2649 7373 2665
rect 7397 2649 7453 2665
rect 7477 2649 7533 2665
rect 5617 2641 5651 2649
rect 5651 2641 5664 2649
rect 5664 2641 5673 2649
rect 5698 2641 5716 2649
rect 5716 2641 5729 2649
rect 5729 2641 5754 2649
rect 5779 2641 5781 2649
rect 5781 2641 5794 2649
rect 5794 2641 5835 2649
rect 5617 2597 5651 2607
rect 5651 2597 5664 2607
rect 5664 2597 5673 2607
rect 5698 2597 5716 2607
rect 5716 2597 5729 2607
rect 5729 2597 5754 2607
rect 5779 2597 5781 2607
rect 5781 2597 5794 2607
rect 5794 2597 5835 2607
rect 5860 2641 5911 2649
rect 5911 2641 5916 2649
rect 5941 2641 5976 2649
rect 5976 2641 5989 2649
rect 5989 2641 5997 2649
rect 6022 2641 6041 2649
rect 6041 2641 6054 2649
rect 6054 2641 6078 2649
rect 6103 2641 6106 2649
rect 6106 2641 6119 2649
rect 6119 2641 6159 2649
rect 5860 2597 5911 2607
rect 5911 2597 5916 2607
rect 5941 2597 5976 2607
rect 5976 2597 5989 2607
rect 5989 2597 5997 2607
rect 6022 2597 6041 2607
rect 6041 2597 6054 2607
rect 6054 2597 6078 2607
rect 6103 2597 6106 2607
rect 6106 2597 6119 2607
rect 6119 2597 6159 2607
rect 6184 2641 6236 2649
rect 6236 2641 6240 2649
rect 6265 2641 6301 2649
rect 6301 2641 6314 2649
rect 6314 2641 6321 2649
rect 6346 2641 6366 2649
rect 6366 2641 6379 2649
rect 6379 2641 6402 2649
rect 6427 2641 6431 2649
rect 6431 2641 6444 2649
rect 6444 2641 6483 2649
rect 6508 2641 6509 2649
rect 6509 2641 6561 2649
rect 6561 2641 6564 2649
rect 6589 2641 6626 2649
rect 6626 2641 6639 2649
rect 6639 2641 6645 2649
rect 6670 2641 6691 2649
rect 6691 2641 6704 2649
rect 6704 2641 6726 2649
rect 6751 2641 6756 2649
rect 6756 2641 6769 2649
rect 6769 2641 6807 2649
rect 6832 2641 6834 2649
rect 6834 2641 6886 2649
rect 6886 2641 6888 2649
rect 6913 2641 6951 2649
rect 6951 2641 6964 2649
rect 6964 2641 6969 2649
rect 6994 2641 7016 2649
rect 7016 2641 7029 2649
rect 7029 2641 7050 2649
rect 7075 2641 7081 2649
rect 7081 2641 7094 2649
rect 7094 2641 7131 2649
rect 7156 2641 7159 2649
rect 7159 2641 7211 2649
rect 7211 2641 7212 2649
rect 7237 2641 7276 2649
rect 7276 2641 7289 2649
rect 7289 2641 7293 2649
rect 7317 2641 7341 2649
rect 7341 2641 7354 2649
rect 7354 2641 7373 2649
rect 7397 2641 7406 2649
rect 7406 2641 7419 2649
rect 7419 2641 7453 2649
rect 7477 2641 7484 2649
rect 7484 2641 7533 2649
rect 6184 2597 6236 2607
rect 6236 2597 6240 2607
rect 6265 2597 6301 2607
rect 6301 2597 6314 2607
rect 6314 2597 6321 2607
rect 6346 2597 6366 2607
rect 6366 2597 6379 2607
rect 6379 2597 6402 2607
rect 6427 2597 6431 2607
rect 6431 2597 6444 2607
rect 6444 2597 6483 2607
rect 6508 2597 6509 2607
rect 6509 2597 6561 2607
rect 6561 2597 6564 2607
rect 6589 2597 6626 2607
rect 6626 2597 6639 2607
rect 6639 2597 6645 2607
rect 6670 2597 6691 2607
rect 6691 2597 6704 2607
rect 6704 2597 6726 2607
rect 6751 2597 6756 2607
rect 6756 2597 6769 2607
rect 6769 2597 6807 2607
rect 6832 2597 6834 2607
rect 6834 2597 6886 2607
rect 6886 2597 6888 2607
rect 6913 2597 6951 2607
rect 6951 2597 6964 2607
rect 6964 2597 6969 2607
rect 6994 2597 7016 2607
rect 7016 2597 7029 2607
rect 7029 2597 7050 2607
rect 7075 2597 7081 2607
rect 7081 2597 7094 2607
rect 7094 2597 7131 2607
rect 7156 2597 7159 2607
rect 7159 2597 7211 2607
rect 7211 2597 7212 2607
rect 7237 2597 7276 2607
rect 7276 2597 7289 2607
rect 7289 2597 7293 2607
rect 7317 2597 7341 2607
rect 7341 2597 7354 2607
rect 7354 2597 7373 2607
rect 7397 2597 7406 2607
rect 7406 2597 7419 2607
rect 7419 2597 7453 2607
rect 7477 2597 7484 2607
rect 7484 2597 7533 2607
rect 5617 2581 5673 2597
rect 5698 2581 5754 2597
rect 5779 2581 5835 2597
rect 5860 2581 5916 2597
rect 5941 2581 5997 2597
rect 6022 2581 6078 2597
rect 6103 2581 6159 2597
rect 6184 2581 6240 2597
rect 6265 2581 6321 2597
rect 6346 2581 6402 2597
rect 6427 2581 6483 2597
rect 6508 2581 6564 2597
rect 6589 2581 6645 2597
rect 6670 2581 6726 2597
rect 6751 2581 6807 2597
rect 6832 2581 6888 2597
rect 6913 2581 6969 2597
rect 6994 2581 7050 2597
rect 7075 2581 7131 2597
rect 7156 2581 7212 2597
rect 7237 2581 7293 2597
rect 7317 2581 7373 2597
rect 7397 2581 7453 2597
rect 7477 2581 7533 2597
rect 5617 2551 5651 2581
rect 5651 2551 5664 2581
rect 5664 2551 5673 2581
rect 5698 2551 5716 2581
rect 5716 2551 5729 2581
rect 5729 2551 5754 2581
rect 5779 2551 5781 2581
rect 5781 2551 5794 2581
rect 5794 2551 5835 2581
rect 5860 2551 5911 2581
rect 5911 2551 5916 2581
rect 5941 2551 5976 2581
rect 5976 2551 5989 2581
rect 5989 2551 5997 2581
rect 6022 2551 6041 2581
rect 6041 2551 6054 2581
rect 6054 2551 6078 2581
rect 6103 2551 6106 2581
rect 6106 2551 6119 2581
rect 6119 2551 6159 2581
rect 6184 2551 6236 2581
rect 6236 2551 6240 2581
rect 6265 2551 6301 2581
rect 6301 2551 6314 2581
rect 6314 2551 6321 2581
rect 6346 2551 6366 2581
rect 6366 2551 6379 2581
rect 6379 2551 6402 2581
rect 6427 2551 6431 2581
rect 6431 2551 6444 2581
rect 6444 2551 6483 2581
rect 6508 2551 6509 2581
rect 6509 2551 6561 2581
rect 6561 2551 6564 2581
rect 6589 2551 6626 2581
rect 6626 2551 6639 2581
rect 6639 2551 6645 2581
rect 6670 2551 6691 2581
rect 6691 2551 6704 2581
rect 6704 2551 6726 2581
rect 6751 2551 6756 2581
rect 6756 2551 6769 2581
rect 6769 2551 6807 2581
rect 6832 2551 6834 2581
rect 6834 2551 6886 2581
rect 6886 2551 6888 2581
rect 6913 2551 6951 2581
rect 6951 2551 6964 2581
rect 6964 2551 6969 2581
rect 6994 2551 7016 2581
rect 7016 2551 7029 2581
rect 7029 2551 7050 2581
rect 7075 2551 7081 2581
rect 7081 2551 7094 2581
rect 7094 2551 7131 2581
rect 7156 2551 7159 2581
rect 7159 2551 7211 2581
rect 7211 2551 7212 2581
rect 7237 2551 7276 2581
rect 7276 2551 7289 2581
rect 7289 2551 7293 2581
rect 7317 2551 7341 2581
rect 7341 2551 7354 2581
rect 7354 2551 7373 2581
rect 7397 2551 7406 2581
rect 7406 2551 7419 2581
rect 7419 2551 7453 2581
rect 7477 2551 7484 2581
rect 7484 2551 7533 2581
rect 5617 2513 5673 2517
rect 5698 2513 5754 2517
rect 5779 2513 5835 2517
rect 5860 2513 5916 2517
rect 5941 2513 5997 2517
rect 6022 2513 6078 2517
rect 6103 2513 6159 2517
rect 6184 2513 6240 2517
rect 6265 2513 6321 2517
rect 6346 2513 6402 2517
rect 6427 2513 6483 2517
rect 6508 2513 6564 2517
rect 6589 2513 6645 2517
rect 6670 2513 6726 2517
rect 6751 2513 6807 2517
rect 6832 2513 6888 2517
rect 6913 2513 6969 2517
rect 6994 2513 7050 2517
rect 7075 2513 7131 2517
rect 7156 2513 7212 2517
rect 7237 2513 7293 2517
rect 7317 2513 7373 2517
rect 7397 2513 7453 2517
rect 7477 2513 7533 2517
rect 5617 2461 5651 2513
rect 5651 2461 5664 2513
rect 5664 2461 5673 2513
rect 5698 2461 5716 2513
rect 5716 2461 5729 2513
rect 5729 2461 5754 2513
rect 5779 2461 5781 2513
rect 5781 2461 5794 2513
rect 5794 2461 5835 2513
rect 5860 2461 5911 2513
rect 5911 2461 5916 2513
rect 5941 2461 5976 2513
rect 5976 2461 5989 2513
rect 5989 2461 5997 2513
rect 6022 2461 6041 2513
rect 6041 2461 6054 2513
rect 6054 2461 6078 2513
rect 6103 2461 6106 2513
rect 6106 2461 6119 2513
rect 6119 2461 6159 2513
rect 6184 2461 6236 2513
rect 6236 2461 6240 2513
rect 6265 2461 6301 2513
rect 6301 2461 6314 2513
rect 6314 2461 6321 2513
rect 6346 2461 6366 2513
rect 6366 2461 6379 2513
rect 6379 2461 6402 2513
rect 6427 2461 6431 2513
rect 6431 2461 6444 2513
rect 6444 2461 6483 2513
rect 6508 2461 6509 2513
rect 6509 2461 6561 2513
rect 6561 2461 6564 2513
rect 6589 2461 6626 2513
rect 6626 2461 6639 2513
rect 6639 2461 6645 2513
rect 6670 2461 6691 2513
rect 6691 2461 6704 2513
rect 6704 2461 6726 2513
rect 6751 2461 6756 2513
rect 6756 2461 6769 2513
rect 6769 2461 6807 2513
rect 6832 2461 6834 2513
rect 6834 2461 6886 2513
rect 6886 2461 6888 2513
rect 6913 2461 6951 2513
rect 6951 2461 6964 2513
rect 6964 2461 6969 2513
rect 6994 2461 7016 2513
rect 7016 2461 7029 2513
rect 7029 2461 7050 2513
rect 7075 2461 7081 2513
rect 7081 2461 7094 2513
rect 7094 2461 7131 2513
rect 7156 2461 7159 2513
rect 7159 2461 7211 2513
rect 7211 2461 7212 2513
rect 7237 2461 7276 2513
rect 7276 2461 7289 2513
rect 7289 2461 7293 2513
rect 7317 2461 7341 2513
rect 7341 2461 7354 2513
rect 7354 2461 7373 2513
rect 7397 2461 7406 2513
rect 7406 2461 7419 2513
rect 7419 2461 7453 2513
rect 7477 2461 7484 2513
rect 7484 2461 7533 2513
rect 3195 2263 3251 2264
rect 3277 2263 3333 2264
rect 3359 2263 3415 2264
rect 3441 2263 3497 2264
rect 3523 2263 3579 2264
rect 3605 2263 3661 2264
rect 3687 2263 3743 2264
rect 3769 2263 3825 2264
rect 3851 2263 3907 2264
rect 3933 2263 3989 2264
rect 4015 2263 4071 2264
rect 4097 2263 4153 2264
rect 4179 2263 4235 2264
rect 4261 2263 4317 2264
rect 4343 2263 4399 2264
rect 4425 2263 4481 2264
rect 4507 2263 4563 2264
rect 4589 2263 4645 2264
rect 4671 2263 4727 2264
rect 4753 2263 4809 2264
rect 4835 2263 4891 2264
rect 3195 2211 3244 2263
rect 3244 2211 3251 2263
rect 3277 2211 3310 2263
rect 3310 2211 3324 2263
rect 3324 2211 3333 2263
rect 3359 2211 3376 2263
rect 3376 2211 3390 2263
rect 3390 2211 3415 2263
rect 3441 2211 3442 2263
rect 3442 2211 3456 2263
rect 3456 2211 3497 2263
rect 3523 2211 3574 2263
rect 3574 2211 3579 2263
rect 3605 2211 3640 2263
rect 3640 2211 3654 2263
rect 3654 2211 3661 2263
rect 3687 2211 3706 2263
rect 3706 2211 3720 2263
rect 3720 2211 3743 2263
rect 3769 2211 3772 2263
rect 3772 2211 3786 2263
rect 3786 2211 3825 2263
rect 3851 2211 3852 2263
rect 3852 2211 3904 2263
rect 3904 2211 3907 2263
rect 3933 2211 3970 2263
rect 3970 2211 3984 2263
rect 3984 2211 3989 2263
rect 4015 2211 4036 2263
rect 4036 2211 4050 2263
rect 4050 2211 4071 2263
rect 4097 2211 4102 2263
rect 4102 2211 4116 2263
rect 4116 2211 4153 2263
rect 4179 2211 4182 2263
rect 4182 2211 4234 2263
rect 4234 2211 4235 2263
rect 4261 2211 4300 2263
rect 4300 2211 4314 2263
rect 4314 2211 4317 2263
rect 4343 2211 4366 2263
rect 4366 2211 4380 2263
rect 4380 2211 4399 2263
rect 4425 2211 4432 2263
rect 4432 2211 4446 2263
rect 4446 2211 4481 2263
rect 4507 2211 4512 2263
rect 4512 2211 4563 2263
rect 4589 2211 4630 2263
rect 4630 2211 4644 2263
rect 4644 2211 4645 2263
rect 4671 2211 4696 2263
rect 4696 2211 4710 2263
rect 4710 2211 4727 2263
rect 4753 2211 4762 2263
rect 4762 2211 4776 2263
rect 4776 2211 4809 2263
rect 4835 2211 4841 2263
rect 4841 2211 4891 2263
rect 3195 2208 3251 2211
rect 3277 2208 3333 2211
rect 3359 2208 3415 2211
rect 3441 2208 3497 2211
rect 3523 2208 3579 2211
rect 3605 2208 3661 2211
rect 3687 2208 3743 2211
rect 3769 2208 3825 2211
rect 3851 2208 3907 2211
rect 3933 2208 3989 2211
rect 4015 2208 4071 2211
rect 4097 2208 4153 2211
rect 4179 2208 4235 2211
rect 4261 2208 4317 2211
rect 4343 2208 4399 2211
rect 4425 2208 4481 2211
rect 4507 2208 4563 2211
rect 4589 2208 4645 2211
rect 4671 2208 4727 2211
rect 4753 2208 4809 2211
rect 4835 2208 4891 2211
rect 4917 2208 4973 2264
rect 4999 2208 5055 2264
rect 5080 2208 5136 2264
rect 5161 2208 5217 2264
rect 5242 2208 5298 2264
rect 3195 2145 3244 2182
rect 3244 2145 3251 2182
rect 3277 2145 3310 2182
rect 3310 2145 3324 2182
rect 3324 2145 3333 2182
rect 3359 2145 3376 2182
rect 3376 2145 3390 2182
rect 3390 2145 3415 2182
rect 3441 2145 3442 2182
rect 3442 2145 3456 2182
rect 3456 2145 3497 2182
rect 3523 2145 3574 2182
rect 3574 2145 3579 2182
rect 3605 2145 3640 2182
rect 3640 2145 3654 2182
rect 3654 2145 3661 2182
rect 3687 2145 3706 2182
rect 3706 2145 3720 2182
rect 3720 2145 3743 2182
rect 3769 2145 3772 2182
rect 3772 2145 3786 2182
rect 3786 2145 3825 2182
rect 3851 2145 3852 2182
rect 3852 2145 3904 2182
rect 3904 2145 3907 2182
rect 3933 2145 3970 2182
rect 3970 2145 3984 2182
rect 3984 2145 3989 2182
rect 4015 2145 4036 2182
rect 4036 2145 4050 2182
rect 4050 2145 4071 2182
rect 4097 2145 4102 2182
rect 4102 2145 4116 2182
rect 4116 2145 4153 2182
rect 4179 2145 4182 2182
rect 4182 2145 4234 2182
rect 4234 2145 4235 2182
rect 4261 2145 4300 2182
rect 4300 2145 4314 2182
rect 4314 2145 4317 2182
rect 4343 2145 4366 2182
rect 4366 2145 4380 2182
rect 4380 2145 4399 2182
rect 4425 2145 4432 2182
rect 4432 2145 4446 2182
rect 4446 2145 4481 2182
rect 4507 2145 4512 2182
rect 4512 2145 4563 2182
rect 4589 2145 4630 2182
rect 4630 2145 4644 2182
rect 4644 2145 4645 2182
rect 4671 2145 4696 2182
rect 4696 2145 4710 2182
rect 4710 2145 4727 2182
rect 4753 2145 4762 2182
rect 4762 2145 4776 2182
rect 4776 2145 4809 2182
rect 4835 2145 4841 2182
rect 4841 2145 4891 2182
rect 3195 2131 3251 2145
rect 3277 2131 3333 2145
rect 3359 2131 3415 2145
rect 3441 2131 3497 2145
rect 3523 2131 3579 2145
rect 3605 2131 3661 2145
rect 3687 2131 3743 2145
rect 3769 2131 3825 2145
rect 3851 2131 3907 2145
rect 3933 2131 3989 2145
rect 4015 2131 4071 2145
rect 4097 2131 4153 2145
rect 4179 2131 4235 2145
rect 4261 2131 4317 2145
rect 4343 2131 4399 2145
rect 4425 2131 4481 2145
rect 4507 2131 4563 2145
rect 4589 2131 4645 2145
rect 4671 2131 4727 2145
rect 4753 2131 4809 2145
rect 4835 2131 4891 2145
rect 3195 2126 3244 2131
rect 3244 2126 3251 2131
rect 3277 2126 3310 2131
rect 3310 2126 3324 2131
rect 3324 2126 3333 2131
rect 3359 2126 3376 2131
rect 3376 2126 3390 2131
rect 3390 2126 3415 2131
rect 3441 2126 3442 2131
rect 3442 2126 3456 2131
rect 3456 2126 3497 2131
rect 3195 2079 3244 2100
rect 3244 2079 3251 2100
rect 3277 2079 3310 2100
rect 3310 2079 3324 2100
rect 3324 2079 3333 2100
rect 3359 2079 3376 2100
rect 3376 2079 3390 2100
rect 3390 2079 3415 2100
rect 3441 2079 3442 2100
rect 3442 2079 3456 2100
rect 3456 2079 3497 2100
rect 3523 2126 3574 2131
rect 3574 2126 3579 2131
rect 3605 2126 3640 2131
rect 3640 2126 3654 2131
rect 3654 2126 3661 2131
rect 3687 2126 3706 2131
rect 3706 2126 3720 2131
rect 3720 2126 3743 2131
rect 3769 2126 3772 2131
rect 3772 2126 3786 2131
rect 3786 2126 3825 2131
rect 3851 2126 3852 2131
rect 3852 2126 3904 2131
rect 3904 2126 3907 2131
rect 3933 2126 3970 2131
rect 3970 2126 3984 2131
rect 3984 2126 3989 2131
rect 4015 2126 4036 2131
rect 4036 2126 4050 2131
rect 4050 2126 4071 2131
rect 4097 2126 4102 2131
rect 4102 2126 4116 2131
rect 4116 2126 4153 2131
rect 4179 2126 4182 2131
rect 4182 2126 4234 2131
rect 4234 2126 4235 2131
rect 4261 2126 4300 2131
rect 4300 2126 4314 2131
rect 4314 2126 4317 2131
rect 4343 2126 4366 2131
rect 4366 2126 4380 2131
rect 4380 2126 4399 2131
rect 4425 2126 4432 2131
rect 4432 2126 4446 2131
rect 4446 2126 4481 2131
rect 4507 2126 4512 2131
rect 4512 2126 4563 2131
rect 3523 2079 3574 2100
rect 3574 2079 3579 2100
rect 3605 2079 3640 2100
rect 3640 2079 3654 2100
rect 3654 2079 3661 2100
rect 3687 2079 3706 2100
rect 3706 2079 3720 2100
rect 3720 2079 3743 2100
rect 3769 2079 3772 2100
rect 3772 2079 3786 2100
rect 3786 2079 3825 2100
rect 3851 2079 3852 2100
rect 3852 2079 3904 2100
rect 3904 2079 3907 2100
rect 3933 2079 3970 2100
rect 3970 2079 3984 2100
rect 3984 2079 3989 2100
rect 4015 2079 4036 2100
rect 4036 2079 4050 2100
rect 4050 2079 4071 2100
rect 4097 2079 4102 2100
rect 4102 2079 4116 2100
rect 4116 2079 4153 2100
rect 4179 2079 4182 2100
rect 4182 2079 4234 2100
rect 4234 2079 4235 2100
rect 4261 2079 4300 2100
rect 4300 2079 4314 2100
rect 4314 2079 4317 2100
rect 4343 2079 4366 2100
rect 4366 2079 4380 2100
rect 4380 2079 4399 2100
rect 4425 2079 4432 2100
rect 4432 2079 4446 2100
rect 4446 2079 4481 2100
rect 4507 2079 4512 2100
rect 4512 2079 4563 2100
rect 4589 2126 4630 2131
rect 4630 2126 4644 2131
rect 4644 2126 4645 2131
rect 4671 2126 4696 2131
rect 4696 2126 4710 2131
rect 4710 2126 4727 2131
rect 4753 2126 4762 2131
rect 4762 2126 4776 2131
rect 4776 2126 4809 2131
rect 4835 2126 4841 2131
rect 4841 2126 4891 2131
rect 4917 2126 4973 2182
rect 4999 2126 5055 2182
rect 5080 2126 5136 2182
rect 5161 2126 5217 2182
rect 5242 2126 5298 2182
rect 4589 2079 4630 2100
rect 4630 2079 4644 2100
rect 4644 2079 4645 2100
rect 4671 2079 4696 2100
rect 4696 2079 4710 2100
rect 4710 2079 4727 2100
rect 4753 2079 4762 2100
rect 4762 2079 4776 2100
rect 4776 2079 4809 2100
rect 4835 2079 4841 2100
rect 4841 2079 4891 2100
rect 3195 2065 3251 2079
rect 3277 2065 3333 2079
rect 3359 2065 3415 2079
rect 3441 2065 3497 2079
rect 3523 2065 3579 2079
rect 3605 2065 3661 2079
rect 3687 2065 3743 2079
rect 3769 2065 3825 2079
rect 3851 2065 3907 2079
rect 3933 2065 3989 2079
rect 4015 2065 4071 2079
rect 4097 2065 4153 2079
rect 4179 2065 4235 2079
rect 4261 2065 4317 2079
rect 4343 2065 4399 2079
rect 4425 2065 4481 2079
rect 4507 2065 4563 2079
rect 4589 2065 4645 2079
rect 4671 2065 4727 2079
rect 4753 2065 4809 2079
rect 4835 2065 4891 2079
rect 3195 2044 3244 2065
rect 3244 2044 3251 2065
rect 3277 2044 3310 2065
rect 3310 2044 3324 2065
rect 3324 2044 3333 2065
rect 3359 2044 3376 2065
rect 3376 2044 3390 2065
rect 3390 2044 3415 2065
rect 3441 2044 3442 2065
rect 3442 2044 3456 2065
rect 3456 2044 3497 2065
rect 3195 2013 3244 2018
rect 3244 2013 3251 2018
rect 3277 2013 3310 2018
rect 3310 2013 3324 2018
rect 3324 2013 3333 2018
rect 3359 2013 3376 2018
rect 3376 2013 3390 2018
rect 3390 2013 3415 2018
rect 3441 2013 3442 2018
rect 3442 2013 3456 2018
rect 3456 2013 3497 2018
rect 3523 2044 3574 2065
rect 3574 2044 3579 2065
rect 3605 2044 3640 2065
rect 3640 2044 3654 2065
rect 3654 2044 3661 2065
rect 3687 2044 3706 2065
rect 3706 2044 3720 2065
rect 3720 2044 3743 2065
rect 3769 2044 3772 2065
rect 3772 2044 3786 2065
rect 3786 2044 3825 2065
rect 3851 2044 3852 2065
rect 3852 2044 3904 2065
rect 3904 2044 3907 2065
rect 3933 2044 3970 2065
rect 3970 2044 3984 2065
rect 3984 2044 3989 2065
rect 4015 2044 4036 2065
rect 4036 2044 4050 2065
rect 4050 2044 4071 2065
rect 4097 2044 4102 2065
rect 4102 2044 4116 2065
rect 4116 2044 4153 2065
rect 4179 2044 4182 2065
rect 4182 2044 4234 2065
rect 4234 2044 4235 2065
rect 4261 2044 4300 2065
rect 4300 2044 4314 2065
rect 4314 2044 4317 2065
rect 4343 2044 4366 2065
rect 4366 2044 4380 2065
rect 4380 2044 4399 2065
rect 4425 2044 4432 2065
rect 4432 2044 4446 2065
rect 4446 2044 4481 2065
rect 4507 2044 4512 2065
rect 4512 2044 4563 2065
rect 3523 2013 3574 2018
rect 3574 2013 3579 2018
rect 3605 2013 3640 2018
rect 3640 2013 3654 2018
rect 3654 2013 3661 2018
rect 3687 2013 3706 2018
rect 3706 2013 3720 2018
rect 3720 2013 3743 2018
rect 3769 2013 3772 2018
rect 3772 2013 3786 2018
rect 3786 2013 3825 2018
rect 3851 2013 3852 2018
rect 3852 2013 3904 2018
rect 3904 2013 3907 2018
rect 3933 2013 3970 2018
rect 3970 2013 3984 2018
rect 3984 2013 3989 2018
rect 4015 2013 4036 2018
rect 4036 2013 4050 2018
rect 4050 2013 4071 2018
rect 4097 2013 4102 2018
rect 4102 2013 4116 2018
rect 4116 2013 4153 2018
rect 4179 2013 4182 2018
rect 4182 2013 4234 2018
rect 4234 2013 4235 2018
rect 4261 2013 4300 2018
rect 4300 2013 4314 2018
rect 4314 2013 4317 2018
rect 4343 2013 4366 2018
rect 4366 2013 4380 2018
rect 4380 2013 4399 2018
rect 4425 2013 4432 2018
rect 4432 2013 4446 2018
rect 4446 2013 4481 2018
rect 4507 2013 4512 2018
rect 4512 2013 4563 2018
rect 4589 2044 4630 2065
rect 4630 2044 4644 2065
rect 4644 2044 4645 2065
rect 4671 2044 4696 2065
rect 4696 2044 4710 2065
rect 4710 2044 4727 2065
rect 4753 2044 4762 2065
rect 4762 2044 4776 2065
rect 4776 2044 4809 2065
rect 4835 2044 4841 2065
rect 4841 2044 4891 2065
rect 4917 2044 4973 2100
rect 4999 2044 5055 2100
rect 5080 2044 5136 2100
rect 5161 2044 5217 2100
rect 5242 2044 5298 2100
rect 4589 2013 4630 2018
rect 4630 2013 4644 2018
rect 4644 2013 4645 2018
rect 4671 2013 4696 2018
rect 4696 2013 4710 2018
rect 4710 2013 4727 2018
rect 4753 2013 4762 2018
rect 4762 2013 4776 2018
rect 4776 2013 4809 2018
rect 4835 2013 4841 2018
rect 4841 2013 4891 2018
rect 3195 1999 3251 2013
rect 3277 1999 3333 2013
rect 3359 1999 3415 2013
rect 3441 1999 3497 2013
rect 3523 1999 3579 2013
rect 3605 1999 3661 2013
rect 3687 1999 3743 2013
rect 3769 1999 3825 2013
rect 3851 1999 3907 2013
rect 3933 1999 3989 2013
rect 4015 1999 4071 2013
rect 4097 1999 4153 2013
rect 4179 1999 4235 2013
rect 4261 1999 4317 2013
rect 4343 1999 4399 2013
rect 4425 1999 4481 2013
rect 4507 1999 4563 2013
rect 4589 1999 4645 2013
rect 4671 1999 4727 2013
rect 4753 1999 4809 2013
rect 4835 1999 4891 2013
rect 3195 1962 3244 1999
rect 3244 1962 3251 1999
rect 3277 1962 3310 1999
rect 3310 1962 3324 1999
rect 3324 1962 3333 1999
rect 3359 1962 3376 1999
rect 3376 1962 3390 1999
rect 3390 1962 3415 1999
rect 3441 1962 3442 1999
rect 3442 1962 3456 1999
rect 3456 1962 3497 1999
rect 3523 1962 3574 1999
rect 3574 1962 3579 1999
rect 3605 1962 3640 1999
rect 3640 1962 3654 1999
rect 3654 1962 3661 1999
rect 3687 1962 3706 1999
rect 3706 1962 3720 1999
rect 3720 1962 3743 1999
rect 3769 1962 3772 1999
rect 3772 1962 3786 1999
rect 3786 1962 3825 1999
rect 3851 1962 3852 1999
rect 3852 1962 3904 1999
rect 3904 1962 3907 1999
rect 3933 1962 3970 1999
rect 3970 1962 3984 1999
rect 3984 1962 3989 1999
rect 4015 1962 4036 1999
rect 4036 1962 4050 1999
rect 4050 1962 4071 1999
rect 4097 1962 4102 1999
rect 4102 1962 4116 1999
rect 4116 1962 4153 1999
rect 4179 1962 4182 1999
rect 4182 1962 4234 1999
rect 4234 1962 4235 1999
rect 4261 1962 4300 1999
rect 4300 1962 4314 1999
rect 4314 1962 4317 1999
rect 4343 1962 4366 1999
rect 4366 1962 4380 1999
rect 4380 1962 4399 1999
rect 4425 1962 4432 1999
rect 4432 1962 4446 1999
rect 4446 1962 4481 1999
rect 4507 1962 4512 1999
rect 4512 1962 4563 1999
rect 4589 1962 4630 1999
rect 4630 1962 4644 1999
rect 4644 1962 4645 1999
rect 4671 1962 4696 1999
rect 4696 1962 4710 1999
rect 4710 1962 4727 1999
rect 4753 1962 4762 1999
rect 4762 1962 4776 1999
rect 4776 1962 4809 1999
rect 4835 1962 4841 1999
rect 4841 1962 4891 1999
rect 4917 1962 4973 2018
rect 4999 1962 5055 2018
rect 5080 1962 5136 2018
rect 5161 1962 5217 2018
rect 5242 1962 5298 2018
rect 3195 1933 3251 1936
rect 3277 1933 3333 1936
rect 3359 1933 3415 1936
rect 3441 1933 3497 1936
rect 3523 1933 3579 1936
rect 3605 1933 3661 1936
rect 3687 1933 3743 1936
rect 3769 1933 3825 1936
rect 3851 1933 3907 1936
rect 3933 1933 3989 1936
rect 4015 1933 4071 1936
rect 4097 1933 4153 1936
rect 4179 1933 4235 1936
rect 4261 1933 4317 1936
rect 4343 1933 4399 1936
rect 4425 1933 4481 1936
rect 4507 1933 4563 1936
rect 4589 1933 4645 1936
rect 4671 1933 4727 1936
rect 4753 1933 4809 1936
rect 4835 1933 4891 1936
rect 3195 1881 3244 1933
rect 3244 1881 3251 1933
rect 3277 1881 3310 1933
rect 3310 1881 3324 1933
rect 3324 1881 3333 1933
rect 3359 1881 3376 1933
rect 3376 1881 3390 1933
rect 3390 1881 3415 1933
rect 3441 1881 3442 1933
rect 3442 1881 3456 1933
rect 3456 1881 3497 1933
rect 3523 1881 3574 1933
rect 3574 1881 3579 1933
rect 3605 1881 3640 1933
rect 3640 1881 3654 1933
rect 3654 1881 3661 1933
rect 3687 1881 3706 1933
rect 3706 1881 3720 1933
rect 3720 1881 3743 1933
rect 3769 1881 3772 1933
rect 3772 1881 3786 1933
rect 3786 1881 3825 1933
rect 3851 1881 3852 1933
rect 3852 1881 3904 1933
rect 3904 1881 3907 1933
rect 3933 1881 3970 1933
rect 3970 1881 3984 1933
rect 3984 1881 3989 1933
rect 4015 1881 4036 1933
rect 4036 1881 4050 1933
rect 4050 1881 4071 1933
rect 4097 1881 4102 1933
rect 4102 1881 4116 1933
rect 4116 1881 4153 1933
rect 4179 1881 4182 1933
rect 4182 1881 4234 1933
rect 4234 1881 4235 1933
rect 4261 1881 4300 1933
rect 4300 1881 4314 1933
rect 4314 1881 4317 1933
rect 4343 1881 4366 1933
rect 4366 1881 4380 1933
rect 4380 1881 4399 1933
rect 4425 1881 4432 1933
rect 4432 1881 4446 1933
rect 4446 1881 4481 1933
rect 4507 1881 4512 1933
rect 4512 1881 4563 1933
rect 4589 1881 4630 1933
rect 4630 1881 4644 1933
rect 4644 1881 4645 1933
rect 4671 1881 4696 1933
rect 4696 1881 4710 1933
rect 4710 1881 4727 1933
rect 4753 1881 4762 1933
rect 4762 1881 4776 1933
rect 4776 1881 4809 1933
rect 4835 1881 4841 1933
rect 4841 1881 4891 1933
rect 3195 1880 3251 1881
rect 3277 1880 3333 1881
rect 3359 1880 3415 1881
rect 3441 1880 3497 1881
rect 3523 1880 3579 1881
rect 3605 1880 3661 1881
rect 3687 1880 3743 1881
rect 3769 1880 3825 1881
rect 3851 1880 3907 1881
rect 3933 1880 3989 1881
rect 4015 1880 4071 1881
rect 4097 1880 4153 1881
rect 4179 1880 4235 1881
rect 4261 1880 4317 1881
rect 4343 1880 4399 1881
rect 4425 1880 4481 1881
rect 4507 1880 4563 1881
rect 4589 1880 4645 1881
rect 4671 1880 4727 1881
rect 4753 1880 4809 1881
rect 4835 1880 4891 1881
rect 4917 1880 4973 1936
rect 4999 1880 5055 1936
rect 5080 1880 5136 1936
rect 5161 1880 5217 1936
rect 5242 1880 5298 1936
rect 5624 2169 5628 2225
rect 5628 2169 5680 2225
rect 5704 2169 5760 2225
rect 5784 2169 5840 2225
rect 5864 2169 5920 2225
rect 5944 2169 6000 2225
rect 6024 2169 6080 2225
rect 6104 2169 6160 2225
rect 6184 2169 6240 2225
rect 6264 2169 6320 2225
rect 5624 2087 5628 2143
rect 5628 2087 5680 2143
rect 5704 2087 5760 2143
rect 5784 2087 5840 2143
rect 5864 2087 5920 2143
rect 5944 2087 6000 2143
rect 6024 2087 6080 2143
rect 6104 2087 6160 2143
rect 6184 2087 6240 2143
rect 6264 2087 6320 2143
rect 5624 2005 5628 2061
rect 5628 2005 5680 2061
rect 5704 2005 5760 2061
rect 5784 2005 5840 2061
rect 5864 2005 5920 2061
rect 5944 2005 6000 2061
rect 6024 2005 6080 2061
rect 6104 2005 6160 2061
rect 6184 2005 6240 2061
rect 6264 2005 6320 2061
rect 5624 1923 5628 1979
rect 5628 1923 5680 1979
rect 5704 1923 5760 1979
rect 5784 1923 5840 1979
rect 5864 1923 5920 1979
rect 5944 1923 6000 1979
rect 6024 1923 6080 1979
rect 6104 1923 6160 1979
rect 6184 1923 6240 1979
rect 6264 1923 6320 1979
rect 5624 1841 5628 1897
rect 5628 1841 5680 1897
rect 5704 1841 5760 1897
rect 5784 1841 5840 1897
rect 5864 1841 5920 1897
rect 5944 1841 6000 1897
rect 6024 1841 6080 1897
rect 6104 1841 6160 1897
rect 6184 1841 6240 1897
rect 6264 1841 6320 1897
rect 5624 1759 5628 1815
rect 5628 1759 5680 1815
rect 5704 1759 5760 1815
rect 5784 1759 5840 1815
rect 5864 1759 5920 1815
rect 5944 1759 6000 1815
rect 6024 1759 6080 1815
rect 6104 1759 6160 1815
rect 6184 1759 6240 1815
rect 6264 1759 6320 1815
rect 5624 1677 5628 1733
rect 5628 1677 5680 1733
rect 5704 1677 5760 1733
rect 5784 1677 5840 1733
rect 5864 1677 5920 1733
rect 5944 1677 6000 1733
rect 6024 1677 6080 1733
rect 6104 1677 6160 1733
rect 6184 1677 6240 1733
rect 6264 1677 6320 1733
rect 5624 1595 5628 1651
rect 5628 1595 5680 1651
rect 5704 1595 5760 1651
rect 5784 1595 5840 1651
rect 5864 1595 5920 1651
rect 5944 1595 6000 1651
rect 6024 1595 6080 1651
rect 6104 1595 6160 1651
rect 6184 1595 6240 1651
rect 6264 1595 6320 1651
rect 5624 1513 5628 1569
rect 5628 1513 5680 1569
rect 5704 1513 5760 1569
rect 5784 1513 5840 1569
rect 5864 1513 5920 1569
rect 5944 1513 6000 1569
rect 6024 1513 6080 1569
rect 6104 1513 6160 1569
rect 6184 1513 6240 1569
rect 6264 1513 6320 1569
rect 5624 1431 5628 1487
rect 5628 1431 5680 1487
rect 5704 1431 5760 1487
rect 5784 1431 5840 1487
rect 5864 1431 5920 1487
rect 5944 1431 6000 1487
rect 6024 1431 6080 1487
rect 6104 1431 6160 1487
rect 6184 1431 6240 1487
rect 6264 1431 6320 1487
rect 5624 1349 5628 1405
rect 5628 1349 5680 1405
rect 5704 1349 5760 1405
rect 5784 1349 5840 1405
rect 5864 1349 5920 1405
rect 5944 1349 6000 1405
rect 6024 1349 6080 1405
rect 6104 1349 6160 1405
rect 6184 1349 6240 1405
rect 6264 1349 6320 1405
rect 5624 1267 5628 1323
rect 5628 1267 5680 1323
rect 5704 1267 5760 1323
rect 5784 1267 5840 1323
rect 5864 1267 5920 1323
rect 5944 1267 6000 1323
rect 6024 1267 6080 1323
rect 6104 1267 6160 1323
rect 6184 1267 6240 1323
rect 6264 1267 6320 1323
rect 5624 1185 5628 1241
rect 5628 1185 5680 1241
rect 5704 1185 5760 1241
rect 5784 1185 5840 1241
rect 5864 1185 5920 1241
rect 5944 1185 6000 1241
rect 6024 1185 6080 1241
rect 6104 1185 6160 1241
rect 6184 1185 6240 1241
rect 6264 1185 6320 1241
rect 5624 1152 5628 1159
rect 5628 1152 5680 1159
rect 5704 1152 5760 1159
rect 5784 1152 5840 1159
rect 5864 1152 5920 1159
rect 5944 1152 6000 1159
rect 6024 1152 6080 1159
rect 6104 1152 6160 1159
rect 6184 1152 6240 1159
rect 6264 1152 6320 1159
rect 5624 1139 5680 1152
rect 5704 1139 5760 1152
rect 5784 1139 5840 1152
rect 5864 1139 5920 1152
rect 5944 1139 6000 1152
rect 6024 1139 6080 1152
rect 6104 1139 6160 1152
rect 6184 1139 6240 1152
rect 6264 1139 6320 1152
rect 5624 1103 5628 1139
rect 5628 1103 5680 1139
rect 5704 1103 5744 1139
rect 5744 1103 5756 1139
rect 5756 1103 5760 1139
rect 5784 1103 5808 1139
rect 5808 1103 5820 1139
rect 5820 1103 5840 1139
rect 5864 1103 5872 1139
rect 5872 1103 5884 1139
rect 5884 1103 5920 1139
rect 5944 1103 5948 1139
rect 5948 1103 6000 1139
rect 6024 1103 6064 1139
rect 6064 1103 6076 1139
rect 6076 1103 6080 1139
rect 6104 1103 6128 1139
rect 6128 1103 6140 1139
rect 6140 1103 6160 1139
rect 6184 1103 6192 1139
rect 6192 1103 6204 1139
rect 6204 1103 6240 1139
rect 6264 1103 6268 1139
rect 6268 1103 6320 1139
rect 5624 1074 5680 1077
rect 5704 1074 5760 1077
rect 5784 1074 5840 1077
rect 5864 1074 5920 1077
rect 5944 1074 6000 1077
rect 6024 1074 6080 1077
rect 6104 1074 6160 1077
rect 6184 1074 6240 1077
rect 6264 1074 6320 1077
rect 5624 1022 5628 1074
rect 5628 1022 5680 1074
rect 5704 1022 5744 1074
rect 5744 1022 5756 1074
rect 5756 1022 5760 1074
rect 5784 1022 5808 1074
rect 5808 1022 5820 1074
rect 5820 1022 5840 1074
rect 5864 1022 5872 1074
rect 5872 1022 5884 1074
rect 5884 1022 5920 1074
rect 5944 1022 5948 1074
rect 5948 1022 6000 1074
rect 6024 1022 6064 1074
rect 6064 1022 6076 1074
rect 6076 1022 6080 1074
rect 6104 1022 6128 1074
rect 6128 1022 6140 1074
rect 6140 1022 6160 1074
rect 6184 1022 6192 1074
rect 6192 1022 6204 1074
rect 6204 1022 6240 1074
rect 6264 1022 6268 1074
rect 6268 1022 6320 1074
rect 5624 1021 5680 1022
rect 5704 1021 5760 1022
rect 5784 1021 5840 1022
rect 5864 1021 5920 1022
rect 5944 1021 6000 1022
rect 6024 1021 6080 1022
rect 6104 1021 6160 1022
rect 6184 1021 6240 1022
rect 6264 1021 6320 1022
rect 5624 957 5628 994
rect 5628 957 5680 994
rect 5704 957 5744 994
rect 5744 957 5756 994
rect 5756 957 5760 994
rect 5784 957 5808 994
rect 5808 957 5820 994
rect 5820 957 5840 994
rect 5864 957 5872 994
rect 5872 957 5884 994
rect 5884 957 5920 994
rect 5944 957 5948 994
rect 5948 957 6000 994
rect 6024 957 6064 994
rect 6064 957 6076 994
rect 6076 957 6080 994
rect 6104 957 6128 994
rect 6128 957 6140 994
rect 6140 957 6160 994
rect 6184 957 6192 994
rect 6192 957 6204 994
rect 6204 957 6240 994
rect 6264 957 6268 994
rect 6268 957 6320 994
rect 5624 944 5680 957
rect 5704 944 5760 957
rect 5784 944 5840 957
rect 5864 944 5920 957
rect 5944 944 6000 957
rect 6024 944 6080 957
rect 6104 944 6160 957
rect 6184 944 6240 957
rect 6264 944 6320 957
rect 5624 938 5628 944
rect 5628 938 5680 944
rect 5624 892 5628 911
rect 5628 892 5680 911
rect 5704 938 5744 944
rect 5744 938 5756 944
rect 5756 938 5760 944
rect 5784 938 5808 944
rect 5808 938 5820 944
rect 5820 938 5840 944
rect 5864 938 5872 944
rect 5872 938 5884 944
rect 5884 938 5920 944
rect 5944 938 5948 944
rect 5948 938 6000 944
rect 5704 892 5744 911
rect 5744 892 5756 911
rect 5756 892 5760 911
rect 5784 892 5808 911
rect 5808 892 5820 911
rect 5820 892 5840 911
rect 5864 892 5872 911
rect 5872 892 5884 911
rect 5884 892 5920 911
rect 5944 892 5948 911
rect 5948 892 6000 911
rect 6024 938 6064 944
rect 6064 938 6076 944
rect 6076 938 6080 944
rect 6104 938 6128 944
rect 6128 938 6140 944
rect 6140 938 6160 944
rect 6184 938 6192 944
rect 6192 938 6204 944
rect 6204 938 6240 944
rect 6264 938 6268 944
rect 6268 938 6320 944
rect 6024 892 6064 911
rect 6064 892 6076 911
rect 6076 892 6080 911
rect 6104 892 6128 911
rect 6128 892 6140 911
rect 6140 892 6160 911
rect 6184 892 6192 911
rect 6192 892 6204 911
rect 6204 892 6240 911
rect 6264 892 6268 911
rect 6268 892 6320 911
rect 5624 879 5680 892
rect 5704 879 5760 892
rect 5784 879 5840 892
rect 5864 879 5920 892
rect 5944 879 6000 892
rect 6024 879 6080 892
rect 6104 879 6160 892
rect 6184 879 6240 892
rect 6264 879 6320 892
rect 5624 855 5628 879
rect 5628 855 5680 879
rect 5624 827 5628 828
rect 5628 827 5680 828
rect 5704 855 5744 879
rect 5744 855 5756 879
rect 5756 855 5760 879
rect 5784 855 5808 879
rect 5808 855 5820 879
rect 5820 855 5840 879
rect 5864 855 5872 879
rect 5872 855 5884 879
rect 5884 855 5920 879
rect 5944 855 5948 879
rect 5948 855 6000 879
rect 5704 827 5744 828
rect 5744 827 5756 828
rect 5756 827 5760 828
rect 5784 827 5808 828
rect 5808 827 5820 828
rect 5820 827 5840 828
rect 5864 827 5872 828
rect 5872 827 5884 828
rect 5884 827 5920 828
rect 5944 827 5948 828
rect 5948 827 6000 828
rect 6024 855 6064 879
rect 6064 855 6076 879
rect 6076 855 6080 879
rect 6104 855 6128 879
rect 6128 855 6140 879
rect 6140 855 6160 879
rect 6184 855 6192 879
rect 6192 855 6204 879
rect 6204 855 6240 879
rect 6264 855 6268 879
rect 6268 855 6320 879
rect 6024 827 6064 828
rect 6064 827 6076 828
rect 6076 827 6080 828
rect 6104 827 6128 828
rect 6128 827 6140 828
rect 6140 827 6160 828
rect 6184 827 6192 828
rect 6192 827 6204 828
rect 6204 827 6240 828
rect 6264 827 6268 828
rect 6268 827 6320 828
rect 5624 814 5680 827
rect 5704 814 5760 827
rect 5784 814 5840 827
rect 5864 814 5920 827
rect 5944 814 6000 827
rect 6024 814 6080 827
rect 6104 814 6160 827
rect 6184 814 6240 827
rect 6264 814 6320 827
rect 5624 772 5628 814
rect 5628 772 5680 814
rect 5704 772 5744 814
rect 5744 772 5756 814
rect 5756 772 5760 814
rect 5784 772 5808 814
rect 5808 772 5820 814
rect 5820 772 5840 814
rect 5864 772 5872 814
rect 5872 772 5884 814
rect 5884 772 5920 814
rect 5944 772 5948 814
rect 5948 772 6000 814
rect 6024 772 6064 814
rect 6064 772 6076 814
rect 6076 772 6080 814
rect 6104 772 6128 814
rect 6128 772 6140 814
rect 6140 772 6160 814
rect 6184 772 6192 814
rect 6192 772 6204 814
rect 6204 772 6240 814
rect 6264 772 6268 814
rect 6268 772 6320 814
rect 5624 697 5628 745
rect 5628 697 5680 745
rect 5704 697 5744 745
rect 5744 697 5756 745
rect 5756 697 5760 745
rect 5784 697 5808 745
rect 5808 697 5820 745
rect 5820 697 5840 745
rect 5864 697 5872 745
rect 5872 697 5884 745
rect 5884 697 5920 745
rect 5944 697 5948 745
rect 5948 697 6000 745
rect 6024 697 6064 745
rect 6064 697 6076 745
rect 6076 697 6080 745
rect 6104 697 6128 745
rect 6128 697 6140 745
rect 6140 697 6160 745
rect 6184 697 6192 745
rect 6192 697 6204 745
rect 6204 697 6240 745
rect 6264 697 6268 745
rect 6268 697 6320 745
rect 5624 689 5680 697
rect 5704 689 5760 697
rect 5784 689 5840 697
rect 5864 689 5920 697
rect 5944 689 6000 697
rect 6024 689 6080 697
rect 6104 689 6160 697
rect 6184 689 6240 697
rect 6264 689 6320 697
rect 5624 632 5628 662
rect 5628 632 5680 662
rect 5704 632 5744 662
rect 5744 632 5756 662
rect 5756 632 5760 662
rect 5784 632 5808 662
rect 5808 632 5820 662
rect 5820 632 5840 662
rect 5864 632 5872 662
rect 5872 632 5884 662
rect 5884 632 5920 662
rect 5944 632 5948 662
rect 5948 632 6000 662
rect 6024 632 6064 662
rect 6064 632 6076 662
rect 6076 632 6080 662
rect 6104 632 6128 662
rect 6128 632 6140 662
rect 6140 632 6160 662
rect 6184 632 6192 662
rect 6192 632 6204 662
rect 6204 632 6240 662
rect 6264 632 6268 662
rect 6268 632 6320 662
rect 5624 619 5680 632
rect 5704 619 5760 632
rect 5784 619 5840 632
rect 5864 619 5920 632
rect 5944 619 6000 632
rect 6024 619 6080 632
rect 6104 619 6160 632
rect 6184 619 6240 632
rect 6264 619 6320 632
rect 5624 606 5628 619
rect 5628 606 5680 619
rect 5624 567 5628 579
rect 5628 567 5680 579
rect 5704 606 5744 619
rect 5744 606 5756 619
rect 5756 606 5760 619
rect 5784 606 5808 619
rect 5808 606 5820 619
rect 5820 606 5840 619
rect 5864 606 5872 619
rect 5872 606 5884 619
rect 5884 606 5920 619
rect 5944 606 5948 619
rect 5948 606 6000 619
rect 5704 567 5744 579
rect 5744 567 5756 579
rect 5756 567 5760 579
rect 5784 567 5808 579
rect 5808 567 5820 579
rect 5820 567 5840 579
rect 5864 567 5872 579
rect 5872 567 5884 579
rect 5884 567 5920 579
rect 5944 567 5948 579
rect 5948 567 6000 579
rect 6024 606 6064 619
rect 6064 606 6076 619
rect 6076 606 6080 619
rect 6104 606 6128 619
rect 6128 606 6140 619
rect 6140 606 6160 619
rect 6184 606 6192 619
rect 6192 606 6204 619
rect 6204 606 6240 619
rect 6264 606 6268 619
rect 6268 606 6320 619
rect 6024 567 6064 579
rect 6064 567 6076 579
rect 6076 567 6080 579
rect 6104 567 6128 579
rect 6128 567 6140 579
rect 6140 567 6160 579
rect 6184 567 6192 579
rect 6192 567 6204 579
rect 6204 567 6240 579
rect 6264 567 6268 579
rect 6268 567 6320 579
rect 5624 554 5680 567
rect 5704 554 5760 567
rect 5784 554 5840 567
rect 5864 554 5920 567
rect 5944 554 6000 567
rect 6024 554 6080 567
rect 6104 554 6160 567
rect 6184 554 6240 567
rect 6264 554 6320 567
rect 5624 523 5628 554
rect 5628 523 5680 554
rect 5704 523 5744 554
rect 5744 523 5756 554
rect 5756 523 5760 554
rect 5784 523 5808 554
rect 5808 523 5820 554
rect 5820 523 5840 554
rect 5864 523 5872 554
rect 5872 523 5884 554
rect 5884 523 5920 554
rect 5944 523 5948 554
rect 5948 523 6000 554
rect 6024 523 6064 554
rect 6064 523 6076 554
rect 6076 523 6080 554
rect 6104 523 6128 554
rect 6128 523 6140 554
rect 6140 523 6160 554
rect 6184 523 6192 554
rect 6192 523 6204 554
rect 6204 523 6240 554
rect 6264 523 6268 554
rect 6268 523 6320 554
rect 5624 489 5680 496
rect 5704 489 5760 496
rect 5784 489 5840 496
rect 5864 489 5920 496
rect 5944 489 6000 496
rect 6024 489 6080 496
rect 6104 489 6160 496
rect 6184 489 6240 496
rect 6264 489 6320 496
rect 5624 440 5628 489
rect 5628 440 5680 489
rect 5704 440 5744 489
rect 5744 440 5756 489
rect 5756 440 5760 489
rect 5784 440 5808 489
rect 5808 440 5820 489
rect 5820 440 5840 489
rect 5864 440 5872 489
rect 5872 440 5884 489
rect 5884 440 5920 489
rect 5944 440 5948 489
rect 5948 440 6000 489
rect 6024 440 6064 489
rect 6064 440 6076 489
rect 6076 440 6080 489
rect 6104 440 6128 489
rect 6128 440 6140 489
rect 6140 440 6160 489
rect 6184 440 6192 489
rect 6192 440 6204 489
rect 6204 440 6240 489
rect 6264 440 6268 489
rect 6268 440 6320 489
rect 6615 2190 6663 2239
rect 6663 2190 6671 2239
rect 6615 2183 6671 2190
rect 6701 2190 6711 2239
rect 6711 2190 6757 2239
rect 6787 2190 6811 2239
rect 6811 2190 6843 2239
rect 6873 2190 6911 2239
rect 6911 2190 6929 2239
rect 6959 2190 6963 2239
rect 6963 2190 7011 2239
rect 7011 2190 7015 2239
rect 7045 2190 7063 2239
rect 7063 2190 7101 2239
rect 7131 2190 7163 2239
rect 7163 2190 7187 2239
rect 7217 2190 7263 2239
rect 7263 2190 7273 2239
rect 6701 2183 6757 2190
rect 6787 2183 6843 2190
rect 6873 2183 6929 2190
rect 6959 2183 7015 2190
rect 7045 2183 7101 2190
rect 7131 2183 7187 2190
rect 7217 2183 7273 2190
rect 7303 2190 7311 2239
rect 7311 2190 7359 2239
rect 7303 2183 7359 2190
rect 6615 2108 6671 2157
rect 6615 2101 6663 2108
rect 6663 2101 6671 2108
rect 6701 2108 6757 2157
rect 6787 2108 6843 2157
rect 6873 2108 6929 2157
rect 6959 2108 7015 2157
rect 7045 2108 7101 2157
rect 7131 2108 7187 2157
rect 7217 2108 7273 2157
rect 6701 2101 6711 2108
rect 6711 2101 6757 2108
rect 6787 2101 6811 2108
rect 6811 2101 6843 2108
rect 6873 2101 6911 2108
rect 6911 2101 6929 2108
rect 6959 2101 6963 2108
rect 6963 2101 7011 2108
rect 7011 2101 7015 2108
rect 7045 2101 7063 2108
rect 7063 2101 7101 2108
rect 7131 2101 7163 2108
rect 7163 2101 7187 2108
rect 7217 2101 7263 2108
rect 7263 2101 7273 2108
rect 7303 2108 7359 2157
rect 7303 2101 7311 2108
rect 7311 2101 7359 2108
rect 6615 2056 6663 2075
rect 6663 2056 6671 2075
rect 6615 2019 6671 2056
rect 6701 2056 6711 2075
rect 6711 2056 6757 2075
rect 6787 2056 6811 2075
rect 6811 2056 6843 2075
rect 6873 2056 6911 2075
rect 6911 2056 6929 2075
rect 6959 2056 6963 2075
rect 6963 2056 7011 2075
rect 7011 2056 7015 2075
rect 7045 2056 7063 2075
rect 7063 2056 7101 2075
rect 7131 2056 7163 2075
rect 7163 2056 7187 2075
rect 7217 2056 7263 2075
rect 7263 2056 7273 2075
rect 6701 2019 6757 2056
rect 6787 2019 6843 2056
rect 6873 2019 6929 2056
rect 6959 2019 7015 2056
rect 7045 2019 7101 2056
rect 7131 2019 7187 2056
rect 7217 2019 7273 2056
rect 7303 2056 7311 2075
rect 7311 2056 7359 2075
rect 7303 2019 7359 2056
rect 6615 1973 6671 1993
rect 6615 1937 6663 1973
rect 6663 1937 6671 1973
rect 6701 1973 6757 1993
rect 6787 1973 6843 1993
rect 6873 1973 6929 1993
rect 6959 1973 7015 1993
rect 7045 1973 7101 1993
rect 7131 1973 7187 1993
rect 7217 1973 7273 1993
rect 6701 1937 6711 1973
rect 6711 1937 6757 1973
rect 6787 1937 6811 1973
rect 6811 1937 6843 1973
rect 6873 1937 6911 1973
rect 6911 1937 6929 1973
rect 6959 1937 6963 1973
rect 6963 1937 7011 1973
rect 7011 1937 7015 1973
rect 7045 1937 7063 1973
rect 7063 1937 7101 1973
rect 7131 1937 7163 1973
rect 7163 1937 7187 1973
rect 7217 1937 7263 1973
rect 7263 1937 7273 1973
rect 7303 1973 7359 1993
rect 7303 1937 7311 1973
rect 7311 1937 7359 1973
rect 6615 1855 6671 1911
rect 6701 1855 6757 1911
rect 6787 1855 6843 1911
rect 6873 1855 6929 1911
rect 6959 1855 7015 1911
rect 7045 1855 7101 1911
rect 7131 1855 7187 1911
rect 7217 1855 7273 1911
rect 7303 1855 7359 1911
rect 6615 1786 6663 1828
rect 6663 1786 6671 1828
rect 6615 1772 6671 1786
rect 6701 1786 6711 1828
rect 6711 1786 6757 1828
rect 6787 1786 6811 1828
rect 6811 1786 6843 1828
rect 6873 1786 6911 1828
rect 6911 1786 6929 1828
rect 6959 1786 6963 1828
rect 6963 1786 7011 1828
rect 7011 1786 7015 1828
rect 7045 1786 7063 1828
rect 7063 1786 7101 1828
rect 7131 1786 7163 1828
rect 7163 1786 7187 1828
rect 7217 1786 7263 1828
rect 7263 1786 7273 1828
rect 6701 1772 6757 1786
rect 6787 1772 6843 1786
rect 6873 1772 6929 1786
rect 6959 1772 7015 1786
rect 7045 1772 7101 1786
rect 7131 1772 7187 1786
rect 7217 1772 7273 1786
rect 7303 1786 7311 1828
rect 7311 1786 7359 1828
rect 7303 1772 7359 1786
rect 6615 1703 6671 1745
rect 6615 1689 6663 1703
rect 6663 1689 6671 1703
rect 6701 1703 6757 1745
rect 6787 1703 6843 1745
rect 6873 1703 6929 1745
rect 6959 1703 7015 1745
rect 7045 1703 7101 1745
rect 7131 1703 7187 1745
rect 7217 1703 7273 1745
rect 6701 1689 6711 1703
rect 6711 1689 6757 1703
rect 6787 1689 6811 1703
rect 6811 1689 6843 1703
rect 6873 1689 6911 1703
rect 6911 1689 6929 1703
rect 6959 1689 6963 1703
rect 6963 1689 7011 1703
rect 7011 1689 7015 1703
rect 7045 1689 7063 1703
rect 7063 1689 7101 1703
rect 7131 1689 7163 1703
rect 7163 1689 7187 1703
rect 7217 1689 7263 1703
rect 7263 1689 7273 1703
rect 7303 1703 7359 1745
rect 7303 1689 7311 1703
rect 7311 1689 7359 1703
rect 6615 1651 6663 1662
rect 6663 1651 6671 1662
rect 6615 1606 6671 1651
rect 6701 1651 6711 1662
rect 6711 1651 6757 1662
rect 6787 1651 6811 1662
rect 6811 1651 6843 1662
rect 6873 1651 6911 1662
rect 6911 1651 6929 1662
rect 6959 1651 6963 1662
rect 6963 1651 7011 1662
rect 7011 1651 7015 1662
rect 7045 1651 7063 1662
rect 7063 1651 7101 1662
rect 7131 1651 7163 1662
rect 7163 1651 7187 1662
rect 7217 1651 7263 1662
rect 7263 1651 7273 1662
rect 6701 1606 6757 1651
rect 6787 1606 6843 1651
rect 6873 1606 6929 1651
rect 6959 1606 7015 1651
rect 7045 1606 7101 1651
rect 7131 1606 7187 1651
rect 7217 1606 7273 1651
rect 7303 1651 7311 1662
rect 7311 1651 7359 1662
rect 7303 1606 7359 1651
rect 6615 1568 6671 1579
rect 6615 1523 6663 1568
rect 6663 1523 6671 1568
rect 6701 1568 6757 1579
rect 6787 1568 6843 1579
rect 6873 1568 6929 1579
rect 6959 1568 7015 1579
rect 7045 1568 7101 1579
rect 7131 1568 7187 1579
rect 7217 1568 7273 1579
rect 6701 1523 6711 1568
rect 6711 1523 6757 1568
rect 6787 1523 6811 1568
rect 6811 1523 6843 1568
rect 6873 1523 6911 1568
rect 6911 1523 6929 1568
rect 6959 1523 6963 1568
rect 6963 1523 7011 1568
rect 7011 1523 7015 1568
rect 7045 1523 7063 1568
rect 7063 1523 7101 1568
rect 7131 1523 7163 1568
rect 7163 1523 7187 1568
rect 7217 1523 7263 1568
rect 7263 1523 7273 1568
rect 7303 1568 7359 1579
rect 7303 1523 7311 1568
rect 7311 1523 7359 1568
rect 6615 1440 6671 1496
rect 6701 1440 6757 1496
rect 6787 1440 6843 1496
rect 6873 1440 6929 1496
rect 6959 1440 7015 1496
rect 7045 1440 7101 1496
rect 7131 1440 7187 1496
rect 7217 1440 7273 1496
rect 7303 1440 7359 1496
rect 6615 1381 6663 1413
rect 6663 1381 6671 1413
rect 6615 1357 6671 1381
rect 6701 1381 6711 1413
rect 6711 1381 6757 1413
rect 6787 1381 6811 1413
rect 6811 1381 6843 1413
rect 6873 1381 6911 1413
rect 6911 1381 6929 1413
rect 6959 1381 6963 1413
rect 6963 1381 7011 1413
rect 7011 1381 7015 1413
rect 7045 1381 7063 1413
rect 7063 1381 7101 1413
rect 7131 1381 7163 1413
rect 7163 1381 7187 1413
rect 7217 1381 7263 1413
rect 7263 1381 7273 1413
rect 6701 1357 6757 1381
rect 6787 1357 6843 1381
rect 6873 1357 6929 1381
rect 6959 1357 7015 1381
rect 7045 1357 7101 1381
rect 7131 1357 7187 1381
rect 7217 1357 7273 1381
rect 7303 1381 7311 1413
rect 7311 1381 7359 1413
rect 7303 1357 7359 1381
rect 6615 1298 6671 1330
rect 6615 1274 6663 1298
rect 6663 1274 6671 1298
rect 6701 1298 6757 1330
rect 6787 1298 6843 1330
rect 6873 1298 6929 1330
rect 6959 1298 7015 1330
rect 7045 1298 7101 1330
rect 7131 1298 7187 1330
rect 7217 1298 7273 1330
rect 6701 1274 6711 1298
rect 6711 1274 6757 1298
rect 6787 1274 6811 1298
rect 6811 1274 6843 1298
rect 6873 1274 6911 1298
rect 6911 1274 6929 1298
rect 6959 1274 6963 1298
rect 6963 1274 7011 1298
rect 7011 1274 7015 1298
rect 7045 1274 7063 1298
rect 7063 1274 7101 1298
rect 7131 1274 7163 1298
rect 7163 1274 7187 1298
rect 7217 1274 7263 1298
rect 7263 1274 7273 1298
rect 7303 1298 7359 1330
rect 7303 1274 7311 1298
rect 7311 1274 7359 1298
rect 6615 1246 6663 1247
rect 6663 1246 6671 1247
rect 6615 1191 6671 1246
rect 6701 1246 6711 1247
rect 6711 1246 6757 1247
rect 6787 1246 6811 1247
rect 6811 1246 6843 1247
rect 6873 1246 6911 1247
rect 6911 1246 6929 1247
rect 6959 1246 6963 1247
rect 6963 1246 7011 1247
rect 7011 1246 7015 1247
rect 7045 1246 7063 1247
rect 7063 1246 7101 1247
rect 7131 1246 7163 1247
rect 7163 1246 7187 1247
rect 7217 1246 7263 1247
rect 7263 1246 7273 1247
rect 6701 1191 6757 1246
rect 6787 1191 6843 1246
rect 6873 1191 6929 1246
rect 6959 1191 7015 1246
rect 7045 1191 7101 1246
rect 7131 1191 7187 1246
rect 7217 1191 7273 1246
rect 7303 1246 7311 1247
rect 7311 1246 7359 1247
rect 7303 1191 7359 1246
rect 6615 1163 6671 1164
rect 6615 1111 6663 1163
rect 6663 1111 6671 1163
rect 6615 1108 6671 1111
rect 6701 1163 6757 1164
rect 6787 1163 6843 1164
rect 6873 1163 6929 1164
rect 6959 1163 7015 1164
rect 7045 1163 7101 1164
rect 7131 1163 7187 1164
rect 7217 1163 7273 1164
rect 6701 1111 6711 1163
rect 6711 1111 6757 1163
rect 6787 1111 6811 1163
rect 6811 1111 6843 1163
rect 6873 1111 6911 1163
rect 6911 1111 6929 1163
rect 6959 1111 6963 1163
rect 6963 1111 7011 1163
rect 7011 1111 7015 1163
rect 7045 1111 7063 1163
rect 7063 1111 7101 1163
rect 7131 1111 7163 1163
rect 7163 1111 7187 1163
rect 7217 1111 7263 1163
rect 7263 1111 7273 1163
rect 6701 1108 6757 1111
rect 6787 1108 6843 1111
rect 6873 1108 6929 1111
rect 6959 1108 7015 1111
rect 7045 1108 7101 1111
rect 7131 1108 7187 1111
rect 7217 1108 7273 1111
rect 7303 1163 7359 1164
rect 7303 1111 7311 1163
rect 7311 1111 7359 1163
rect 7303 1108 7359 1111
rect 6615 1028 6671 1081
rect 6615 1025 6663 1028
rect 6663 1025 6671 1028
rect 6701 1028 6757 1081
rect 6787 1028 6843 1081
rect 6873 1028 6929 1081
rect 6959 1028 7015 1081
rect 7045 1028 7101 1081
rect 7131 1028 7187 1081
rect 7217 1028 7273 1081
rect 6701 1025 6711 1028
rect 6711 1025 6757 1028
rect 6787 1025 6811 1028
rect 6811 1025 6843 1028
rect 6873 1025 6911 1028
rect 6911 1025 6929 1028
rect 6959 1025 6963 1028
rect 6963 1025 7011 1028
rect 7011 1025 7015 1028
rect 7045 1025 7063 1028
rect 7063 1025 7101 1028
rect 7131 1025 7163 1028
rect 7163 1025 7187 1028
rect 7217 1025 7263 1028
rect 7263 1025 7273 1028
rect 7303 1028 7359 1081
rect 7303 1025 7311 1028
rect 7311 1025 7359 1028
rect 6615 976 6663 998
rect 6663 976 6671 998
rect 6615 942 6671 976
rect 6701 976 6711 998
rect 6711 976 6757 998
rect 6787 976 6811 998
rect 6811 976 6843 998
rect 6873 976 6911 998
rect 6911 976 6929 998
rect 6959 976 6963 998
rect 6963 976 7011 998
rect 7011 976 7015 998
rect 7045 976 7063 998
rect 7063 976 7101 998
rect 7131 976 7163 998
rect 7163 976 7187 998
rect 7217 976 7263 998
rect 7263 976 7273 998
rect 6701 942 6757 976
rect 6787 942 6843 976
rect 6873 942 6929 976
rect 6959 942 7015 976
rect 7045 942 7101 976
rect 7131 942 7187 976
rect 7217 942 7273 976
rect 7303 976 7311 998
rect 7311 976 7359 998
rect 7303 942 7359 976
rect 6615 893 6671 915
rect 6615 859 6663 893
rect 6663 859 6671 893
rect 6701 893 6757 915
rect 6787 893 6843 915
rect 6873 893 6929 915
rect 6959 893 7015 915
rect 7045 893 7101 915
rect 7131 893 7187 915
rect 7217 893 7273 915
rect 6701 859 6711 893
rect 6711 859 6757 893
rect 6787 859 6811 893
rect 6811 859 6843 893
rect 6873 859 6911 893
rect 6911 859 6929 893
rect 6959 859 6963 893
rect 6963 859 7011 893
rect 7011 859 7015 893
rect 7045 859 7063 893
rect 7063 859 7101 893
rect 7131 859 7163 893
rect 7163 859 7187 893
rect 7217 859 7263 893
rect 7263 859 7273 893
rect 7303 893 7359 915
rect 7303 859 7311 893
rect 7311 859 7359 893
rect 6615 776 6671 832
rect 6701 776 6757 832
rect 6787 776 6843 832
rect 6873 776 6929 832
rect 6959 776 7015 832
rect 7045 776 7101 832
rect 7131 776 7187 832
rect 7217 776 7273 832
rect 7303 776 7359 832
rect 6615 706 6663 749
rect 6663 706 6671 749
rect 6615 693 6671 706
rect 6701 706 6711 749
rect 6711 706 6757 749
rect 6787 706 6811 749
rect 6811 706 6843 749
rect 6873 706 6911 749
rect 6911 706 6929 749
rect 6959 706 6963 749
rect 6963 706 7011 749
rect 7011 706 7015 749
rect 7045 706 7063 749
rect 7063 706 7101 749
rect 7131 706 7163 749
rect 7163 706 7187 749
rect 7217 706 7263 749
rect 7263 706 7273 749
rect 6701 693 6757 706
rect 6787 693 6843 706
rect 6873 693 6929 706
rect 6959 693 7015 706
rect 7045 693 7101 706
rect 7131 693 7187 706
rect 7217 693 7273 706
rect 7303 706 7311 749
rect 7311 706 7359 749
rect 7303 693 7359 706
rect 6615 623 6671 666
rect 6615 610 6663 623
rect 6663 610 6671 623
rect 6701 623 6757 666
rect 6787 623 6843 666
rect 6873 623 6929 666
rect 6959 623 7015 666
rect 7045 623 7101 666
rect 7131 623 7187 666
rect 7217 623 7273 666
rect 6701 610 6711 623
rect 6711 610 6757 623
rect 6787 610 6811 623
rect 6811 610 6843 623
rect 6873 610 6911 623
rect 6911 610 6929 623
rect 6959 610 6963 623
rect 6963 610 7011 623
rect 7011 610 7015 623
rect 7045 610 7063 623
rect 7063 610 7101 623
rect 7131 610 7163 623
rect 7163 610 7187 623
rect 7217 610 7263 623
rect 7263 610 7273 623
rect 7303 623 7359 666
rect 7303 610 7311 623
rect 7311 610 7359 623
rect 6615 571 6663 583
rect 6663 571 6671 583
rect 6615 527 6671 571
rect 6701 571 6711 583
rect 6711 571 6757 583
rect 6787 571 6811 583
rect 6811 571 6843 583
rect 6873 571 6911 583
rect 6911 571 6929 583
rect 6959 571 6963 583
rect 6963 571 7011 583
rect 7011 571 7015 583
rect 7045 571 7063 583
rect 7063 571 7101 583
rect 7131 571 7163 583
rect 7163 571 7187 583
rect 7217 571 7263 583
rect 7263 571 7273 583
rect 6701 527 6757 571
rect 6787 527 6843 571
rect 6873 527 6929 571
rect 6959 527 7015 571
rect 7045 527 7101 571
rect 7131 527 7187 571
rect 7217 527 7273 571
rect 7303 571 7311 583
rect 7311 571 7359 583
rect 7303 527 7359 571
rect 6615 488 6671 500
rect 6615 444 6663 488
rect 6663 444 6671 488
rect 6701 488 6757 500
rect 6787 488 6843 500
rect 6873 488 6929 500
rect 6959 488 7015 500
rect 7045 488 7101 500
rect 7131 488 7187 500
rect 7217 488 7273 500
rect 6701 444 6711 488
rect 6711 444 6757 488
rect 6787 444 6811 488
rect 6811 444 6843 488
rect 6873 444 6911 488
rect 6911 444 6929 488
rect 6959 444 6963 488
rect 6963 444 7011 488
rect 7011 444 7015 488
rect 7045 444 7063 488
rect 7063 444 7101 488
rect 7131 444 7163 488
rect 7163 444 7187 488
rect 7217 444 7263 488
rect 7263 444 7273 488
rect 7303 488 7359 500
rect 7303 444 7311 488
rect 7311 444 7359 488
<< metal3 >>
rect 5608 38724 8218 38735
rect 5608 38668 5613 38724
rect 5669 38668 5696 38724
rect 5752 38668 5779 38724
rect 5835 38668 5861 38724
rect 5917 38668 5943 38724
rect 5999 38668 6025 38724
rect 6081 38668 6107 38724
rect 6163 38668 6189 38724
rect 6245 38668 6271 38724
rect 6327 38668 6353 38724
rect 6409 38668 6435 38724
rect 6491 38668 6517 38724
rect 6573 38668 6599 38724
rect 6655 38668 6681 38724
rect 6737 38668 6763 38724
rect 6819 38668 6845 38724
rect 6901 38668 6927 38724
rect 6983 38668 7009 38724
rect 7065 38668 7091 38724
rect 7147 38668 7173 38724
rect 7229 38668 7255 38724
rect 7311 38668 7337 38724
rect 7393 38668 7419 38724
rect 7475 38668 7501 38724
rect 7557 38668 7583 38724
rect 7639 38668 7665 38724
rect 7721 38668 7747 38724
rect 7803 38668 7829 38724
rect 7885 38668 7911 38724
rect 7967 38668 7993 38724
rect 8049 38668 8075 38724
rect 8131 38668 8157 38724
rect 8213 38668 8218 38724
rect 5608 38644 8218 38668
rect 5608 38588 5613 38644
rect 5669 38588 5696 38644
rect 5752 38588 5779 38644
rect 5835 38588 5861 38644
rect 5917 38588 5943 38644
rect 5999 38588 6025 38644
rect 6081 38588 6107 38644
rect 6163 38588 6189 38644
rect 6245 38588 6271 38644
rect 6327 38588 6353 38644
rect 6409 38588 6435 38644
rect 6491 38588 6517 38644
rect 6573 38588 6599 38644
rect 6655 38588 6681 38644
rect 6737 38588 6763 38644
rect 6819 38588 6845 38644
rect 6901 38588 6927 38644
rect 6983 38588 7009 38644
rect 7065 38588 7091 38644
rect 7147 38588 7173 38644
rect 7229 38588 7255 38644
rect 7311 38588 7337 38644
rect 7393 38588 7419 38644
rect 7475 38588 7501 38644
rect 7557 38588 7583 38644
rect 7639 38588 7665 38644
rect 7721 38588 7747 38644
rect 7803 38588 7829 38644
rect 7885 38588 7911 38644
rect 7967 38588 7993 38644
rect 8049 38588 8075 38644
rect 8131 38588 8157 38644
rect 8213 38588 8218 38644
rect 5608 38564 8218 38588
rect 5608 38508 5613 38564
rect 5669 38508 5696 38564
rect 5752 38508 5779 38564
rect 5835 38508 5861 38564
rect 5917 38508 5943 38564
rect 5999 38508 6025 38564
rect 6081 38508 6107 38564
rect 6163 38508 6189 38564
rect 6245 38508 6271 38564
rect 6327 38508 6353 38564
rect 6409 38508 6435 38564
rect 6491 38508 6517 38564
rect 6573 38508 6599 38564
rect 6655 38508 6681 38564
rect 6737 38508 6763 38564
rect 6819 38508 6845 38564
rect 6901 38508 6927 38564
rect 6983 38508 7009 38564
rect 7065 38508 7091 38564
rect 7147 38508 7173 38564
rect 7229 38508 7255 38564
rect 7311 38508 7337 38564
rect 7393 38508 7419 38564
rect 7475 38508 7501 38564
rect 7557 38508 7583 38564
rect 7639 38508 7665 38564
rect 7721 38508 7747 38564
rect 7803 38508 7829 38564
rect 7885 38508 7911 38564
rect 7967 38508 7993 38564
rect 8049 38508 8075 38564
rect 8131 38508 8157 38564
rect 8213 38508 8218 38564
rect 5608 38484 8218 38508
rect 5608 38428 5613 38484
rect 5669 38428 5696 38484
rect 5752 38428 5779 38484
rect 5835 38428 5861 38484
rect 5917 38428 5943 38484
rect 5999 38428 6025 38484
rect 6081 38428 6107 38484
rect 6163 38428 6189 38484
rect 6245 38428 6271 38484
rect 6327 38428 6353 38484
rect 6409 38428 6435 38484
rect 6491 38428 6517 38484
rect 6573 38428 6599 38484
rect 6655 38428 6681 38484
rect 6737 38428 6763 38484
rect 6819 38428 6845 38484
rect 6901 38428 6927 38484
rect 6983 38428 7009 38484
rect 7065 38428 7091 38484
rect 7147 38428 7173 38484
rect 7229 38428 7255 38484
rect 7311 38428 7337 38484
rect 7393 38428 7419 38484
rect 7475 38428 7501 38484
rect 7557 38428 7583 38484
rect 7639 38428 7665 38484
rect 7721 38428 7747 38484
rect 7803 38428 7829 38484
rect 7885 38428 7911 38484
rect 7967 38428 7993 38484
rect 8049 38428 8075 38484
rect 8131 38428 8157 38484
rect 8213 38428 8218 38484
rect 5608 38404 8218 38428
rect 5608 38348 5613 38404
rect 5669 38348 5696 38404
rect 5752 38348 5779 38404
rect 5835 38348 5861 38404
rect 5917 38348 5943 38404
rect 5999 38348 6025 38404
rect 6081 38348 6107 38404
rect 6163 38348 6189 38404
rect 6245 38348 6271 38404
rect 6327 38348 6353 38404
rect 6409 38348 6435 38404
rect 6491 38348 6517 38404
rect 6573 38348 6599 38404
rect 6655 38348 6681 38404
rect 6737 38348 6763 38404
rect 6819 38348 6845 38404
rect 6901 38348 6927 38404
rect 6983 38348 7009 38404
rect 7065 38348 7091 38404
rect 7147 38348 7173 38404
rect 7229 38348 7255 38404
rect 7311 38348 7337 38404
rect 7393 38348 7419 38404
rect 7475 38348 7501 38404
rect 7557 38348 7583 38404
rect 7639 38348 7665 38404
rect 7721 38348 7747 38404
rect 7803 38348 7829 38404
rect 7885 38348 7911 38404
rect 7967 38348 7993 38404
rect 8049 38348 8075 38404
rect 8131 38348 8157 38404
rect 8213 38348 8218 38404
rect 5608 38324 8218 38348
rect 5608 38268 5613 38324
rect 5669 38268 5696 38324
rect 5752 38268 5779 38324
rect 5835 38268 5861 38324
rect 5917 38268 5943 38324
rect 5999 38268 6025 38324
rect 6081 38268 6107 38324
rect 6163 38268 6189 38324
rect 6245 38268 6271 38324
rect 6327 38268 6353 38324
rect 6409 38268 6435 38324
rect 6491 38268 6517 38324
rect 6573 38268 6599 38324
rect 6655 38268 6681 38324
rect 6737 38268 6763 38324
rect 6819 38268 6845 38324
rect 6901 38268 6927 38324
rect 6983 38268 7009 38324
rect 7065 38268 7091 38324
rect 7147 38268 7173 38324
rect 7229 38268 7255 38324
rect 7311 38268 7337 38324
rect 7393 38268 7419 38324
rect 7475 38268 7501 38324
rect 7557 38268 7583 38324
rect 7639 38268 7665 38324
rect 7721 38268 7747 38324
rect 7803 38268 7829 38324
rect 7885 38268 7911 38324
rect 7967 38268 7993 38324
rect 8049 38268 8075 38324
rect 8131 38268 8157 38324
rect 8213 38268 8218 38324
rect 5608 38244 8218 38268
rect 5608 38188 5613 38244
rect 5669 38188 5696 38244
rect 5752 38188 5779 38244
rect 5835 38188 5861 38244
rect 5917 38188 5943 38244
rect 5999 38188 6025 38244
rect 6081 38188 6107 38244
rect 6163 38188 6189 38244
rect 6245 38188 6271 38244
rect 6327 38188 6353 38244
rect 6409 38188 6435 38244
rect 6491 38188 6517 38244
rect 6573 38188 6599 38244
rect 6655 38188 6681 38244
rect 6737 38188 6763 38244
rect 6819 38188 6845 38244
rect 6901 38188 6927 38244
rect 6983 38188 7009 38244
rect 7065 38188 7091 38244
rect 7147 38188 7173 38244
rect 7229 38188 7255 38244
rect 7311 38188 7337 38244
rect 7393 38188 7419 38244
rect 7475 38188 7501 38244
rect 7557 38188 7583 38244
rect 7639 38188 7665 38244
rect 7721 38188 7747 38244
rect 7803 38188 7829 38244
rect 7885 38188 7911 38244
rect 7967 38188 7993 38244
rect 8049 38188 8075 38244
rect 8131 38188 8157 38244
rect 8213 38188 8218 38244
rect 5608 38164 8218 38188
rect 5608 38108 5613 38164
rect 5669 38108 5696 38164
rect 5752 38108 5779 38164
rect 5835 38108 5861 38164
rect 5917 38108 5943 38164
rect 5999 38108 6025 38164
rect 6081 38108 6107 38164
rect 6163 38108 6189 38164
rect 6245 38108 6271 38164
rect 6327 38108 6353 38164
rect 6409 38108 6435 38164
rect 6491 38108 6517 38164
rect 6573 38108 6599 38164
rect 6655 38108 6681 38164
rect 6737 38108 6763 38164
rect 6819 38108 6845 38164
rect 6901 38108 6927 38164
rect 6983 38108 7009 38164
rect 7065 38108 7091 38164
rect 7147 38108 7173 38164
rect 7229 38108 7255 38164
rect 7311 38108 7337 38164
rect 7393 38108 7419 38164
rect 7475 38108 7501 38164
rect 7557 38108 7583 38164
rect 7639 38108 7665 38164
rect 7721 38108 7747 38164
rect 7803 38108 7829 38164
rect 7885 38108 7911 38164
rect 7967 38108 7993 38164
rect 8049 38108 8075 38164
rect 8131 38108 8157 38164
rect 8213 38108 8218 38164
rect 2724 37987 5308 37992
rect 2724 37931 2738 37987
rect 2794 37931 2819 37987
rect 2875 37931 2900 37987
rect 2956 37931 2981 37987
rect 3037 37931 3062 37987
rect 3118 37931 3143 37987
rect 3199 37931 3224 37987
rect 3280 37931 3305 37987
rect 3361 37931 3386 37987
rect 3442 37931 3467 37987
rect 3523 37931 3548 37987
rect 3604 37931 3629 37987
rect 3685 37931 3710 37987
rect 3766 37931 3791 37987
rect 3847 37931 3872 37987
rect 3928 37931 3953 37987
rect 4009 37931 4034 37987
rect 4090 37931 4115 37987
rect 4171 37931 4196 37987
rect 4252 37931 4277 37987
rect 4333 37931 4358 37987
rect 4414 37931 4439 37987
rect 4495 37931 4520 37987
rect 4576 37931 4601 37987
rect 4657 37931 4682 37987
rect 4738 37931 4763 37987
rect 2724 37907 4763 37931
rect 2724 37851 2738 37907
rect 2794 37851 2819 37907
rect 2875 37851 2900 37907
rect 2956 37851 2981 37907
rect 3037 37851 3062 37907
rect 3118 37851 3143 37907
rect 3199 37851 3224 37907
rect 3280 37851 3305 37907
rect 3361 37851 3386 37907
rect 3442 37851 3467 37907
rect 3523 37851 3548 37907
rect 3604 37851 3629 37907
rect 3685 37851 3710 37907
rect 3766 37851 3791 37907
rect 3847 37851 3872 37907
rect 3928 37851 3953 37907
rect 4009 37851 4034 37907
rect 4090 37851 4115 37907
rect 4171 37851 4196 37907
rect 4252 37851 4277 37907
rect 4333 37851 4358 37907
rect 4414 37851 4439 37907
rect 4495 37851 4520 37907
rect 4576 37851 4601 37907
rect 4657 37851 4682 37907
rect 4738 37851 4763 37907
rect 2724 37827 4763 37851
rect 2724 37771 2738 37827
rect 2794 37771 2819 37827
rect 2875 37771 2900 37827
rect 2956 37771 2981 37827
rect 3037 37771 3062 37827
rect 3118 37771 3143 37827
rect 3199 37771 3224 37827
rect 3280 37771 3305 37827
rect 3361 37771 3386 37827
rect 3442 37771 3467 37827
rect 3523 37771 3548 37827
rect 3604 37771 3629 37827
rect 3685 37771 3710 37827
rect 3766 37771 3791 37827
rect 3847 37771 3872 37827
rect 3928 37771 3953 37827
rect 4009 37771 4034 37827
rect 4090 37771 4115 37827
rect 4171 37771 4196 37827
rect 4252 37771 4277 37827
rect 4333 37771 4358 37827
rect 4414 37771 4439 37827
rect 4495 37771 4520 37827
rect 4576 37771 4601 37827
rect 4657 37771 4682 37827
rect 4738 37771 4763 37827
rect 2724 37747 4763 37771
rect 2724 37691 2738 37747
rect 2794 37691 2819 37747
rect 2875 37691 2900 37747
rect 2956 37691 2981 37747
rect 3037 37691 3062 37747
rect 3118 37691 3143 37747
rect 3199 37691 3224 37747
rect 3280 37691 3305 37747
rect 3361 37691 3386 37747
rect 3442 37691 3467 37747
rect 3523 37691 3548 37747
rect 3604 37691 3629 37747
rect 3685 37691 3710 37747
rect 3766 37691 3791 37747
rect 3847 37691 3872 37747
rect 3928 37691 3953 37747
rect 4009 37691 4034 37747
rect 4090 37691 4115 37747
rect 4171 37691 4196 37747
rect 4252 37691 4277 37747
rect 4333 37691 4358 37747
rect 4414 37691 4439 37747
rect 4495 37691 4520 37747
rect 4576 37691 4601 37747
rect 4657 37691 4682 37747
rect 4738 37691 4763 37747
rect 2724 37667 4763 37691
rect 2724 37611 2738 37667
rect 2794 37611 2819 37667
rect 2875 37611 2900 37667
rect 2956 37611 2981 37667
rect 3037 37611 3062 37667
rect 3118 37611 3143 37667
rect 3199 37611 3224 37667
rect 3280 37611 3305 37667
rect 3361 37611 3386 37667
rect 3442 37611 3467 37667
rect 3523 37611 3548 37667
rect 3604 37611 3629 37667
rect 3685 37611 3710 37667
rect 3766 37611 3791 37667
rect 3847 37611 3872 37667
rect 3928 37611 3953 37667
rect 4009 37611 4034 37667
rect 4090 37611 4115 37667
rect 4171 37611 4196 37667
rect 4252 37611 4277 37667
rect 4333 37611 4358 37667
rect 4414 37611 4439 37667
rect 4495 37611 4520 37667
rect 4576 37611 4601 37667
rect 4657 37611 4682 37667
rect 4738 37611 4763 37667
rect 2724 37587 4763 37611
rect 2724 37531 2738 37587
rect 2794 37531 2819 37587
rect 2875 37531 2900 37587
rect 2956 37531 2981 37587
rect 3037 37531 3062 37587
rect 3118 37531 3143 37587
rect 3199 37531 3224 37587
rect 3280 37531 3305 37587
rect 3361 37531 3386 37587
rect 3442 37531 3467 37587
rect 3523 37531 3548 37587
rect 3604 37531 3629 37587
rect 3685 37531 3710 37587
rect 3766 37531 3791 37587
rect 3847 37531 3872 37587
rect 3928 37531 3953 37587
rect 4009 37531 4034 37587
rect 4090 37531 4115 37587
rect 4171 37531 4196 37587
rect 4252 37531 4277 37587
rect 4333 37531 4358 37587
rect 4414 37531 4439 37587
rect 4495 37531 4520 37587
rect 4576 37531 4601 37587
rect 4657 37531 4682 37587
rect 4738 37531 4763 37587
rect 2724 37507 4763 37531
rect 2724 37451 2738 37507
rect 2794 37451 2819 37507
rect 2875 37451 2900 37507
rect 2956 37451 2981 37507
rect 3037 37451 3062 37507
rect 3118 37451 3143 37507
rect 3199 37451 3224 37507
rect 3280 37451 3305 37507
rect 3361 37451 3386 37507
rect 3442 37451 3467 37507
rect 3523 37451 3548 37507
rect 3604 37451 3629 37507
rect 3685 37451 3710 37507
rect 3766 37451 3791 37507
rect 3847 37451 3872 37507
rect 3928 37451 3953 37507
rect 4009 37451 4034 37507
rect 4090 37451 4115 37507
rect 4171 37451 4196 37507
rect 4252 37451 4277 37507
rect 4333 37451 4358 37507
rect 4414 37451 4439 37507
rect 4495 37451 4520 37507
rect 4576 37451 4601 37507
rect 4657 37451 4682 37507
rect 4738 37451 4763 37507
rect 2724 37427 4763 37451
rect 2724 37371 2738 37427
rect 2794 37371 2819 37427
rect 2875 37371 2900 37427
rect 2956 37371 2981 37427
rect 3037 37371 3062 37427
rect 3118 37371 3143 37427
rect 3199 37371 3224 37427
rect 3280 37371 3305 37427
rect 3361 37371 3386 37427
rect 3442 37371 3467 37427
rect 3523 37371 3548 37427
rect 3604 37371 3629 37427
rect 3685 37371 3710 37427
rect 3766 37371 3791 37427
rect 3847 37371 3872 37427
rect 3928 37371 3953 37427
rect 4009 37371 4034 37427
rect 4090 37371 4115 37427
rect 4171 37371 4196 37427
rect 4252 37371 4277 37427
rect 4333 37371 4358 37427
rect 4414 37371 4439 37427
rect 4495 37371 4520 37427
rect 4576 37371 4601 37427
rect 4657 37371 4682 37427
rect 4738 37371 4763 37427
rect 5299 37371 5308 37987
rect 2724 35987 5308 37371
rect 2724 35931 2733 35987
rect 2789 35931 2814 35987
rect 2870 35931 2895 35987
rect 2951 35931 2976 35987
rect 3032 35931 3057 35987
rect 3113 35931 3138 35987
rect 3194 35931 3219 35987
rect 3275 35931 3300 35987
rect 3356 35931 3381 35987
rect 3437 35931 3462 35987
rect 3518 35931 3543 35987
rect 3599 35931 3624 35987
rect 3680 35931 3705 35987
rect 3761 35931 3786 35987
rect 3842 35931 3867 35987
rect 3923 35931 3948 35987
rect 4004 35931 4029 35987
rect 4085 35931 4110 35987
rect 4166 35931 4191 35987
rect 4247 35931 4272 35987
rect 4328 35931 4353 35987
rect 4409 35931 4434 35987
rect 4490 35931 4515 35987
rect 4571 35931 4596 35987
rect 4652 35931 4677 35987
rect 4733 35931 4758 35987
rect 4814 35931 4839 35987
rect 4895 35931 4920 35987
rect 4976 35931 5001 35987
rect 5057 35931 5082 35987
rect 5138 35931 5163 35987
rect 2724 35907 5163 35931
rect 2724 35851 2733 35907
rect 2789 35851 2814 35907
rect 2870 35851 2895 35907
rect 2951 35851 2976 35907
rect 3032 35851 3057 35907
rect 3113 35851 3138 35907
rect 3194 35851 3219 35907
rect 3275 35851 3300 35907
rect 3356 35851 3381 35907
rect 3437 35851 3462 35907
rect 3518 35851 3543 35907
rect 3599 35851 3624 35907
rect 3680 35851 3705 35907
rect 3761 35851 3786 35907
rect 3842 35851 3867 35907
rect 3923 35851 3948 35907
rect 4004 35851 4029 35907
rect 4085 35851 4110 35907
rect 4166 35851 4191 35907
rect 4247 35851 4272 35907
rect 4328 35851 4353 35907
rect 4409 35851 4434 35907
rect 4490 35851 4515 35907
rect 4571 35851 4596 35907
rect 4652 35851 4677 35907
rect 4733 35851 4758 35907
rect 4814 35851 4839 35907
rect 4895 35851 4920 35907
rect 4976 35851 5001 35907
rect 5057 35851 5082 35907
rect 5138 35851 5163 35907
rect 2724 35827 5163 35851
rect 2724 35771 2733 35827
rect 2789 35771 2814 35827
rect 2870 35771 2895 35827
rect 2951 35771 2976 35827
rect 3032 35771 3057 35827
rect 3113 35771 3138 35827
rect 3194 35771 3219 35827
rect 3275 35771 3300 35827
rect 3356 35771 3381 35827
rect 3437 35771 3462 35827
rect 3518 35771 3543 35827
rect 3599 35771 3624 35827
rect 3680 35771 3705 35827
rect 3761 35771 3786 35827
rect 3842 35771 3867 35827
rect 3923 35771 3948 35827
rect 4004 35771 4029 35827
rect 4085 35771 4110 35827
rect 4166 35771 4191 35827
rect 4247 35771 4272 35827
rect 4328 35771 4353 35827
rect 4409 35771 4434 35827
rect 4490 35771 4515 35827
rect 4571 35771 4596 35827
rect 4652 35771 4677 35827
rect 4733 35771 4758 35827
rect 4814 35771 4839 35827
rect 4895 35771 4920 35827
rect 4976 35771 5001 35827
rect 5057 35771 5082 35827
rect 5138 35771 5163 35827
rect 2724 35747 5163 35771
rect 2724 35691 2733 35747
rect 2789 35691 2814 35747
rect 2870 35691 2895 35747
rect 2951 35691 2976 35747
rect 3032 35691 3057 35747
rect 3113 35691 3138 35747
rect 3194 35691 3219 35747
rect 3275 35691 3300 35747
rect 3356 35691 3381 35747
rect 3437 35691 3462 35747
rect 3518 35691 3543 35747
rect 3599 35691 3624 35747
rect 3680 35691 3705 35747
rect 3761 35691 3786 35747
rect 3842 35691 3867 35747
rect 3923 35691 3948 35747
rect 4004 35691 4029 35747
rect 4085 35691 4110 35747
rect 4166 35691 4191 35747
rect 4247 35691 4272 35747
rect 4328 35691 4353 35747
rect 4409 35691 4434 35747
rect 4490 35691 4515 35747
rect 4571 35691 4596 35747
rect 4652 35691 4677 35747
rect 4733 35691 4758 35747
rect 4814 35691 4839 35747
rect 4895 35691 4920 35747
rect 4976 35691 5001 35747
rect 5057 35691 5082 35747
rect 5138 35691 5163 35747
rect 2724 35667 5163 35691
rect 2724 35611 2733 35667
rect 2789 35611 2814 35667
rect 2870 35611 2895 35667
rect 2951 35611 2976 35667
rect 3032 35611 3057 35667
rect 3113 35611 3138 35667
rect 3194 35611 3219 35667
rect 3275 35611 3300 35667
rect 3356 35611 3381 35667
rect 3437 35611 3462 35667
rect 3518 35611 3543 35667
rect 3599 35611 3624 35667
rect 3680 35611 3705 35667
rect 3761 35611 3786 35667
rect 3842 35611 3867 35667
rect 3923 35611 3948 35667
rect 4004 35611 4029 35667
rect 4085 35611 4110 35667
rect 4166 35611 4191 35667
rect 4247 35611 4272 35667
rect 4328 35611 4353 35667
rect 4409 35611 4434 35667
rect 4490 35611 4515 35667
rect 4571 35611 4596 35667
rect 4652 35611 4677 35667
rect 4733 35611 4758 35667
rect 4814 35611 4839 35667
rect 4895 35611 4920 35667
rect 4976 35611 5001 35667
rect 5057 35611 5082 35667
rect 5138 35611 5163 35667
rect 2724 35587 5163 35611
rect 2724 35531 2733 35587
rect 2789 35531 2814 35587
rect 2870 35531 2895 35587
rect 2951 35531 2976 35587
rect 3032 35531 3057 35587
rect 3113 35531 3138 35587
rect 3194 35531 3219 35587
rect 3275 35531 3300 35587
rect 3356 35531 3381 35587
rect 3437 35531 3462 35587
rect 3518 35531 3543 35587
rect 3599 35531 3624 35587
rect 3680 35531 3705 35587
rect 3761 35531 3786 35587
rect 3842 35531 3867 35587
rect 3923 35531 3948 35587
rect 4004 35531 4029 35587
rect 4085 35531 4110 35587
rect 4166 35531 4191 35587
rect 4247 35531 4272 35587
rect 4328 35531 4353 35587
rect 4409 35531 4434 35587
rect 4490 35531 4515 35587
rect 4571 35531 4596 35587
rect 4652 35531 4677 35587
rect 4733 35531 4758 35587
rect 4814 35531 4839 35587
rect 4895 35531 4920 35587
rect 4976 35531 5001 35587
rect 5057 35531 5082 35587
rect 5138 35531 5163 35587
rect 2724 35507 5163 35531
rect 2724 35451 2733 35507
rect 2789 35451 2814 35507
rect 2870 35451 2895 35507
rect 2951 35451 2976 35507
rect 3032 35451 3057 35507
rect 3113 35451 3138 35507
rect 3194 35451 3219 35507
rect 3275 35451 3300 35507
rect 3356 35451 3381 35507
rect 3437 35451 3462 35507
rect 3518 35451 3543 35507
rect 3599 35451 3624 35507
rect 3680 35451 3705 35507
rect 3761 35451 3786 35507
rect 3842 35451 3867 35507
rect 3923 35451 3948 35507
rect 4004 35451 4029 35507
rect 4085 35451 4110 35507
rect 4166 35451 4191 35507
rect 4247 35451 4272 35507
rect 4328 35451 4353 35507
rect 4409 35451 4434 35507
rect 4490 35451 4515 35507
rect 4571 35451 4596 35507
rect 4652 35451 4677 35507
rect 4733 35451 4758 35507
rect 4814 35451 4839 35507
rect 4895 35451 4920 35507
rect 4976 35451 5001 35507
rect 5057 35451 5082 35507
rect 5138 35451 5163 35507
rect 2724 35427 5163 35451
rect 2724 35371 2733 35427
rect 2789 35371 2814 35427
rect 2870 35371 2895 35427
rect 2951 35371 2976 35427
rect 3032 35371 3057 35427
rect 3113 35371 3138 35427
rect 3194 35371 3219 35427
rect 3275 35371 3300 35427
rect 3356 35371 3381 35427
rect 3437 35371 3462 35427
rect 3518 35371 3543 35427
rect 3599 35371 3624 35427
rect 3680 35371 3705 35427
rect 3761 35371 3786 35427
rect 3842 35371 3867 35427
rect 3923 35371 3948 35427
rect 4004 35371 4029 35427
rect 4085 35371 4110 35427
rect 4166 35371 4191 35427
rect 4247 35371 4272 35427
rect 4328 35371 4353 35427
rect 4409 35371 4434 35427
rect 4490 35371 4515 35427
rect 4571 35371 4596 35427
rect 4652 35371 4677 35427
rect 4733 35371 4758 35427
rect 4814 35371 4839 35427
rect 4895 35371 4920 35427
rect 4976 35371 5001 35427
rect 5057 35371 5082 35427
rect 5138 35371 5163 35427
rect 5299 35371 5308 35987
rect 2724 33987 5308 35371
rect 2724 33931 2733 33987
rect 2789 33931 2814 33987
rect 2870 33931 2895 33987
rect 2951 33931 2976 33987
rect 3032 33931 3057 33987
rect 3113 33931 3138 33987
rect 3194 33931 3219 33987
rect 3275 33931 3300 33987
rect 3356 33931 3381 33987
rect 3437 33931 3462 33987
rect 3518 33931 3543 33987
rect 3599 33931 3624 33987
rect 3680 33931 3705 33987
rect 3761 33931 3786 33987
rect 3842 33931 3867 33987
rect 3923 33931 3948 33987
rect 4004 33931 4029 33987
rect 4085 33931 4110 33987
rect 4166 33931 4191 33987
rect 4247 33931 4272 33987
rect 4328 33931 4353 33987
rect 4409 33931 4434 33987
rect 4490 33931 4515 33987
rect 4571 33931 4596 33987
rect 4652 33931 4677 33987
rect 4733 33931 4758 33987
rect 4814 33931 4839 33987
rect 4895 33931 4920 33987
rect 4976 33931 5001 33987
rect 5057 33931 5082 33987
rect 5138 33931 5163 33987
rect 2724 33907 5163 33931
rect 2724 33851 2733 33907
rect 2789 33851 2814 33907
rect 2870 33851 2895 33907
rect 2951 33851 2976 33907
rect 3032 33851 3057 33907
rect 3113 33851 3138 33907
rect 3194 33851 3219 33907
rect 3275 33851 3300 33907
rect 3356 33851 3381 33907
rect 3437 33851 3462 33907
rect 3518 33851 3543 33907
rect 3599 33851 3624 33907
rect 3680 33851 3705 33907
rect 3761 33851 3786 33907
rect 3842 33851 3867 33907
rect 3923 33851 3948 33907
rect 4004 33851 4029 33907
rect 4085 33851 4110 33907
rect 4166 33851 4191 33907
rect 4247 33851 4272 33907
rect 4328 33851 4353 33907
rect 4409 33851 4434 33907
rect 4490 33851 4515 33907
rect 4571 33851 4596 33907
rect 4652 33851 4677 33907
rect 4733 33851 4758 33907
rect 4814 33851 4839 33907
rect 4895 33851 4920 33907
rect 4976 33851 5001 33907
rect 5057 33851 5082 33907
rect 5138 33851 5163 33907
rect 2724 33827 5163 33851
rect 2724 33771 2733 33827
rect 2789 33771 2814 33827
rect 2870 33771 2895 33827
rect 2951 33771 2976 33827
rect 3032 33771 3057 33827
rect 3113 33771 3138 33827
rect 3194 33771 3219 33827
rect 3275 33771 3300 33827
rect 3356 33771 3381 33827
rect 3437 33771 3462 33827
rect 3518 33771 3543 33827
rect 3599 33771 3624 33827
rect 3680 33771 3705 33827
rect 3761 33771 3786 33827
rect 3842 33771 3867 33827
rect 3923 33771 3948 33827
rect 4004 33771 4029 33827
rect 4085 33771 4110 33827
rect 4166 33771 4191 33827
rect 4247 33771 4272 33827
rect 4328 33771 4353 33827
rect 4409 33771 4434 33827
rect 4490 33771 4515 33827
rect 4571 33771 4596 33827
rect 4652 33771 4677 33827
rect 4733 33771 4758 33827
rect 4814 33771 4839 33827
rect 4895 33771 4920 33827
rect 4976 33771 5001 33827
rect 5057 33771 5082 33827
rect 5138 33771 5163 33827
rect 2724 33747 5163 33771
rect 2724 33691 2733 33747
rect 2789 33691 2814 33747
rect 2870 33691 2895 33747
rect 2951 33691 2976 33747
rect 3032 33691 3057 33747
rect 3113 33691 3138 33747
rect 3194 33691 3219 33747
rect 3275 33691 3300 33747
rect 3356 33691 3381 33747
rect 3437 33691 3462 33747
rect 3518 33691 3543 33747
rect 3599 33691 3624 33747
rect 3680 33691 3705 33747
rect 3761 33691 3786 33747
rect 3842 33691 3867 33747
rect 3923 33691 3948 33747
rect 4004 33691 4029 33747
rect 4085 33691 4110 33747
rect 4166 33691 4191 33747
rect 4247 33691 4272 33747
rect 4328 33691 4353 33747
rect 4409 33691 4434 33747
rect 4490 33691 4515 33747
rect 4571 33691 4596 33747
rect 4652 33691 4677 33747
rect 4733 33691 4758 33747
rect 4814 33691 4839 33747
rect 4895 33691 4920 33747
rect 4976 33691 5001 33747
rect 5057 33691 5082 33747
rect 5138 33691 5163 33747
rect 2724 33667 5163 33691
rect 2724 33611 2733 33667
rect 2789 33611 2814 33667
rect 2870 33611 2895 33667
rect 2951 33611 2976 33667
rect 3032 33611 3057 33667
rect 3113 33611 3138 33667
rect 3194 33611 3219 33667
rect 3275 33611 3300 33667
rect 3356 33611 3381 33667
rect 3437 33611 3462 33667
rect 3518 33611 3543 33667
rect 3599 33611 3624 33667
rect 3680 33611 3705 33667
rect 3761 33611 3786 33667
rect 3842 33611 3867 33667
rect 3923 33611 3948 33667
rect 4004 33611 4029 33667
rect 4085 33611 4110 33667
rect 4166 33611 4191 33667
rect 4247 33611 4272 33667
rect 4328 33611 4353 33667
rect 4409 33611 4434 33667
rect 4490 33611 4515 33667
rect 4571 33611 4596 33667
rect 4652 33611 4677 33667
rect 4733 33611 4758 33667
rect 4814 33611 4839 33667
rect 4895 33611 4920 33667
rect 4976 33611 5001 33667
rect 5057 33611 5082 33667
rect 5138 33611 5163 33667
rect 2724 33587 5163 33611
rect 2724 33531 2733 33587
rect 2789 33531 2814 33587
rect 2870 33531 2895 33587
rect 2951 33531 2976 33587
rect 3032 33531 3057 33587
rect 3113 33531 3138 33587
rect 3194 33531 3219 33587
rect 3275 33531 3300 33587
rect 3356 33531 3381 33587
rect 3437 33531 3462 33587
rect 3518 33531 3543 33587
rect 3599 33531 3624 33587
rect 3680 33531 3705 33587
rect 3761 33531 3786 33587
rect 3842 33531 3867 33587
rect 3923 33531 3948 33587
rect 4004 33531 4029 33587
rect 4085 33531 4110 33587
rect 4166 33531 4191 33587
rect 4247 33531 4272 33587
rect 4328 33531 4353 33587
rect 4409 33531 4434 33587
rect 4490 33531 4515 33587
rect 4571 33531 4596 33587
rect 4652 33531 4677 33587
rect 4733 33531 4758 33587
rect 4814 33531 4839 33587
rect 4895 33531 4920 33587
rect 4976 33531 5001 33587
rect 5057 33531 5082 33587
rect 5138 33531 5163 33587
rect 2724 33507 5163 33531
rect 2724 33451 2733 33507
rect 2789 33451 2814 33507
rect 2870 33451 2895 33507
rect 2951 33451 2976 33507
rect 3032 33451 3057 33507
rect 3113 33451 3138 33507
rect 3194 33451 3219 33507
rect 3275 33451 3300 33507
rect 3356 33451 3381 33507
rect 3437 33451 3462 33507
rect 3518 33451 3543 33507
rect 3599 33451 3624 33507
rect 3680 33451 3705 33507
rect 3761 33451 3786 33507
rect 3842 33451 3867 33507
rect 3923 33451 3948 33507
rect 4004 33451 4029 33507
rect 4085 33451 4110 33507
rect 4166 33451 4191 33507
rect 4247 33451 4272 33507
rect 4328 33451 4353 33507
rect 4409 33451 4434 33507
rect 4490 33451 4515 33507
rect 4571 33451 4596 33507
rect 4652 33451 4677 33507
rect 4733 33451 4758 33507
rect 4814 33451 4839 33507
rect 4895 33451 4920 33507
rect 4976 33451 5001 33507
rect 5057 33451 5082 33507
rect 5138 33451 5163 33507
rect 2724 33427 5163 33451
rect 2724 33371 2733 33427
rect 2789 33371 2814 33427
rect 2870 33371 2895 33427
rect 2951 33371 2976 33427
rect 3032 33371 3057 33427
rect 3113 33371 3138 33427
rect 3194 33371 3219 33427
rect 3275 33371 3300 33427
rect 3356 33371 3381 33427
rect 3437 33371 3462 33427
rect 3518 33371 3543 33427
rect 3599 33371 3624 33427
rect 3680 33371 3705 33427
rect 3761 33371 3786 33427
rect 3842 33371 3867 33427
rect 3923 33371 3948 33427
rect 4004 33371 4029 33427
rect 4085 33371 4110 33427
rect 4166 33371 4191 33427
rect 4247 33371 4272 33427
rect 4328 33371 4353 33427
rect 4409 33371 4434 33427
rect 4490 33371 4515 33427
rect 4571 33371 4596 33427
rect 4652 33371 4677 33427
rect 4733 33371 4758 33427
rect 4814 33371 4839 33427
rect 4895 33371 4920 33427
rect 4976 33371 5001 33427
rect 5057 33371 5082 33427
rect 5138 33371 5163 33427
rect 5299 33371 5308 33987
rect 2724 31987 5308 33371
rect 2724 31931 2733 31987
rect 2789 31931 2814 31987
rect 2870 31931 2895 31987
rect 2951 31931 2976 31987
rect 3032 31931 3057 31987
rect 3113 31931 3138 31987
rect 3194 31931 3219 31987
rect 3275 31931 3300 31987
rect 3356 31931 3381 31987
rect 3437 31931 3462 31987
rect 3518 31931 3543 31987
rect 3599 31931 3624 31987
rect 3680 31931 3705 31987
rect 3761 31931 3786 31987
rect 3842 31931 3867 31987
rect 3923 31931 3948 31987
rect 4004 31931 4029 31987
rect 4085 31931 4110 31987
rect 4166 31931 4191 31987
rect 4247 31931 4272 31987
rect 4328 31931 4353 31987
rect 4409 31931 4434 31987
rect 4490 31931 4515 31987
rect 4571 31931 4596 31987
rect 4652 31931 4677 31987
rect 4733 31931 4758 31987
rect 4814 31931 4839 31987
rect 4895 31931 4920 31987
rect 4976 31931 5001 31987
rect 5057 31931 5082 31987
rect 5138 31931 5163 31987
rect 2724 31907 5163 31931
rect 2724 31851 2733 31907
rect 2789 31851 2814 31907
rect 2870 31851 2895 31907
rect 2951 31851 2976 31907
rect 3032 31851 3057 31907
rect 3113 31851 3138 31907
rect 3194 31851 3219 31907
rect 3275 31851 3300 31907
rect 3356 31851 3381 31907
rect 3437 31851 3462 31907
rect 3518 31851 3543 31907
rect 3599 31851 3624 31907
rect 3680 31851 3705 31907
rect 3761 31851 3786 31907
rect 3842 31851 3867 31907
rect 3923 31851 3948 31907
rect 4004 31851 4029 31907
rect 4085 31851 4110 31907
rect 4166 31851 4191 31907
rect 4247 31851 4272 31907
rect 4328 31851 4353 31907
rect 4409 31851 4434 31907
rect 4490 31851 4515 31907
rect 4571 31851 4596 31907
rect 4652 31851 4677 31907
rect 4733 31851 4758 31907
rect 4814 31851 4839 31907
rect 4895 31851 4920 31907
rect 4976 31851 5001 31907
rect 5057 31851 5082 31907
rect 5138 31851 5163 31907
rect 2724 31827 5163 31851
rect 2724 31771 2733 31827
rect 2789 31771 2814 31827
rect 2870 31771 2895 31827
rect 2951 31771 2976 31827
rect 3032 31771 3057 31827
rect 3113 31771 3138 31827
rect 3194 31771 3219 31827
rect 3275 31771 3300 31827
rect 3356 31771 3381 31827
rect 3437 31771 3462 31827
rect 3518 31771 3543 31827
rect 3599 31771 3624 31827
rect 3680 31771 3705 31827
rect 3761 31771 3786 31827
rect 3842 31771 3867 31827
rect 3923 31771 3948 31827
rect 4004 31771 4029 31827
rect 4085 31771 4110 31827
rect 4166 31771 4191 31827
rect 4247 31771 4272 31827
rect 4328 31771 4353 31827
rect 4409 31771 4434 31827
rect 4490 31771 4515 31827
rect 4571 31771 4596 31827
rect 4652 31771 4677 31827
rect 4733 31771 4758 31827
rect 4814 31771 4839 31827
rect 4895 31771 4920 31827
rect 4976 31771 5001 31827
rect 5057 31771 5082 31827
rect 5138 31771 5163 31827
rect 2724 31747 5163 31771
rect 2724 31691 2733 31747
rect 2789 31691 2814 31747
rect 2870 31691 2895 31747
rect 2951 31691 2976 31747
rect 3032 31691 3057 31747
rect 3113 31691 3138 31747
rect 3194 31691 3219 31747
rect 3275 31691 3300 31747
rect 3356 31691 3381 31747
rect 3437 31691 3462 31747
rect 3518 31691 3543 31747
rect 3599 31691 3624 31747
rect 3680 31691 3705 31747
rect 3761 31691 3786 31747
rect 3842 31691 3867 31747
rect 3923 31691 3948 31747
rect 4004 31691 4029 31747
rect 4085 31691 4110 31747
rect 4166 31691 4191 31747
rect 4247 31691 4272 31747
rect 4328 31691 4353 31747
rect 4409 31691 4434 31747
rect 4490 31691 4515 31747
rect 4571 31691 4596 31747
rect 4652 31691 4677 31747
rect 4733 31691 4758 31747
rect 4814 31691 4839 31747
rect 4895 31691 4920 31747
rect 4976 31691 5001 31747
rect 5057 31691 5082 31747
rect 5138 31691 5163 31747
rect 2724 31667 5163 31691
rect 2724 31611 2733 31667
rect 2789 31611 2814 31667
rect 2870 31611 2895 31667
rect 2951 31611 2976 31667
rect 3032 31611 3057 31667
rect 3113 31611 3138 31667
rect 3194 31611 3219 31667
rect 3275 31611 3300 31667
rect 3356 31611 3381 31667
rect 3437 31611 3462 31667
rect 3518 31611 3543 31667
rect 3599 31611 3624 31667
rect 3680 31611 3705 31667
rect 3761 31611 3786 31667
rect 3842 31611 3867 31667
rect 3923 31611 3948 31667
rect 4004 31611 4029 31667
rect 4085 31611 4110 31667
rect 4166 31611 4191 31667
rect 4247 31611 4272 31667
rect 4328 31611 4353 31667
rect 4409 31611 4434 31667
rect 4490 31611 4515 31667
rect 4571 31611 4596 31667
rect 4652 31611 4677 31667
rect 4733 31611 4758 31667
rect 4814 31611 4839 31667
rect 4895 31611 4920 31667
rect 4976 31611 5001 31667
rect 5057 31611 5082 31667
rect 5138 31611 5163 31667
rect 2724 31587 5163 31611
rect 2724 31531 2733 31587
rect 2789 31531 2814 31587
rect 2870 31531 2895 31587
rect 2951 31531 2976 31587
rect 3032 31531 3057 31587
rect 3113 31531 3138 31587
rect 3194 31531 3219 31587
rect 3275 31531 3300 31587
rect 3356 31531 3381 31587
rect 3437 31531 3462 31587
rect 3518 31531 3543 31587
rect 3599 31531 3624 31587
rect 3680 31531 3705 31587
rect 3761 31531 3786 31587
rect 3842 31531 3867 31587
rect 3923 31531 3948 31587
rect 4004 31531 4029 31587
rect 4085 31531 4110 31587
rect 4166 31531 4191 31587
rect 4247 31531 4272 31587
rect 4328 31531 4353 31587
rect 4409 31531 4434 31587
rect 4490 31531 4515 31587
rect 4571 31531 4596 31587
rect 4652 31531 4677 31587
rect 4733 31531 4758 31587
rect 4814 31531 4839 31587
rect 4895 31531 4920 31587
rect 4976 31531 5001 31587
rect 5057 31531 5082 31587
rect 5138 31531 5163 31587
rect 2724 31507 5163 31531
rect 2724 31451 2733 31507
rect 2789 31451 2814 31507
rect 2870 31451 2895 31507
rect 2951 31451 2976 31507
rect 3032 31451 3057 31507
rect 3113 31451 3138 31507
rect 3194 31451 3219 31507
rect 3275 31451 3300 31507
rect 3356 31451 3381 31507
rect 3437 31451 3462 31507
rect 3518 31451 3543 31507
rect 3599 31451 3624 31507
rect 3680 31451 3705 31507
rect 3761 31451 3786 31507
rect 3842 31451 3867 31507
rect 3923 31451 3948 31507
rect 4004 31451 4029 31507
rect 4085 31451 4110 31507
rect 4166 31451 4191 31507
rect 4247 31451 4272 31507
rect 4328 31451 4353 31507
rect 4409 31451 4434 31507
rect 4490 31451 4515 31507
rect 4571 31451 4596 31507
rect 4652 31451 4677 31507
rect 4733 31451 4758 31507
rect 4814 31451 4839 31507
rect 4895 31451 4920 31507
rect 4976 31451 5001 31507
rect 5057 31451 5082 31507
rect 5138 31451 5163 31507
rect 2724 31427 5163 31451
rect 2724 31371 2733 31427
rect 2789 31371 2814 31427
rect 2870 31371 2895 31427
rect 2951 31371 2976 31427
rect 3032 31371 3057 31427
rect 3113 31371 3138 31427
rect 3194 31371 3219 31427
rect 3275 31371 3300 31427
rect 3356 31371 3381 31427
rect 3437 31371 3462 31427
rect 3518 31371 3543 31427
rect 3599 31371 3624 31427
rect 3680 31371 3705 31427
rect 3761 31371 3786 31427
rect 3842 31371 3867 31427
rect 3923 31371 3948 31427
rect 4004 31371 4029 31427
rect 4085 31371 4110 31427
rect 4166 31371 4191 31427
rect 4247 31371 4272 31427
rect 4328 31371 4353 31427
rect 4409 31371 4434 31427
rect 4490 31371 4515 31427
rect 4571 31371 4596 31427
rect 4652 31371 4677 31427
rect 4733 31371 4758 31427
rect 4814 31371 4839 31427
rect 4895 31371 4920 31427
rect 4976 31371 5001 31427
rect 5057 31371 5082 31427
rect 5138 31371 5163 31427
rect 5299 31371 5308 31987
rect 2724 29987 5308 31371
rect 2724 29931 2733 29987
rect 2789 29931 2814 29987
rect 2870 29931 2895 29987
rect 2951 29931 2976 29987
rect 3032 29931 3057 29987
rect 3113 29931 3138 29987
rect 3194 29931 3219 29987
rect 3275 29931 3300 29987
rect 3356 29931 3381 29987
rect 3437 29931 3462 29987
rect 3518 29931 3543 29987
rect 3599 29931 3624 29987
rect 3680 29931 3705 29987
rect 3761 29931 3786 29987
rect 3842 29931 3867 29987
rect 3923 29931 3948 29987
rect 4004 29931 4029 29987
rect 4085 29931 4110 29987
rect 4166 29931 4191 29987
rect 4247 29931 4272 29987
rect 4328 29931 4353 29987
rect 4409 29931 4434 29987
rect 4490 29931 4515 29987
rect 4571 29931 4596 29987
rect 4652 29931 4677 29987
rect 4733 29931 4758 29987
rect 4814 29931 4839 29987
rect 4895 29931 4920 29987
rect 4976 29931 5001 29987
rect 5057 29931 5082 29987
rect 5138 29931 5163 29987
rect 2724 29907 5163 29931
rect 2724 29851 2733 29907
rect 2789 29851 2814 29907
rect 2870 29851 2895 29907
rect 2951 29851 2976 29907
rect 3032 29851 3057 29907
rect 3113 29851 3138 29907
rect 3194 29851 3219 29907
rect 3275 29851 3300 29907
rect 3356 29851 3381 29907
rect 3437 29851 3462 29907
rect 3518 29851 3543 29907
rect 3599 29851 3624 29907
rect 3680 29851 3705 29907
rect 3761 29851 3786 29907
rect 3842 29851 3867 29907
rect 3923 29851 3948 29907
rect 4004 29851 4029 29907
rect 4085 29851 4110 29907
rect 4166 29851 4191 29907
rect 4247 29851 4272 29907
rect 4328 29851 4353 29907
rect 4409 29851 4434 29907
rect 4490 29851 4515 29907
rect 4571 29851 4596 29907
rect 4652 29851 4677 29907
rect 4733 29851 4758 29907
rect 4814 29851 4839 29907
rect 4895 29851 4920 29907
rect 4976 29851 5001 29907
rect 5057 29851 5082 29907
rect 5138 29851 5163 29907
rect 2724 29827 5163 29851
rect 2724 29771 2733 29827
rect 2789 29771 2814 29827
rect 2870 29771 2895 29827
rect 2951 29771 2976 29827
rect 3032 29771 3057 29827
rect 3113 29771 3138 29827
rect 3194 29771 3219 29827
rect 3275 29771 3300 29827
rect 3356 29771 3381 29827
rect 3437 29771 3462 29827
rect 3518 29771 3543 29827
rect 3599 29771 3624 29827
rect 3680 29771 3705 29827
rect 3761 29771 3786 29827
rect 3842 29771 3867 29827
rect 3923 29771 3948 29827
rect 4004 29771 4029 29827
rect 4085 29771 4110 29827
rect 4166 29771 4191 29827
rect 4247 29771 4272 29827
rect 4328 29771 4353 29827
rect 4409 29771 4434 29827
rect 4490 29771 4515 29827
rect 4571 29771 4596 29827
rect 4652 29771 4677 29827
rect 4733 29771 4758 29827
rect 4814 29771 4839 29827
rect 4895 29771 4920 29827
rect 4976 29771 5001 29827
rect 5057 29771 5082 29827
rect 5138 29771 5163 29827
rect 2724 29747 5163 29771
rect 2724 29691 2733 29747
rect 2789 29691 2814 29747
rect 2870 29691 2895 29747
rect 2951 29691 2976 29747
rect 3032 29691 3057 29747
rect 3113 29691 3138 29747
rect 3194 29691 3219 29747
rect 3275 29691 3300 29747
rect 3356 29691 3381 29747
rect 3437 29691 3462 29747
rect 3518 29691 3543 29747
rect 3599 29691 3624 29747
rect 3680 29691 3705 29747
rect 3761 29691 3786 29747
rect 3842 29691 3867 29747
rect 3923 29691 3948 29747
rect 4004 29691 4029 29747
rect 4085 29691 4110 29747
rect 4166 29691 4191 29747
rect 4247 29691 4272 29747
rect 4328 29691 4353 29747
rect 4409 29691 4434 29747
rect 4490 29691 4515 29747
rect 4571 29691 4596 29747
rect 4652 29691 4677 29747
rect 4733 29691 4758 29747
rect 4814 29691 4839 29747
rect 4895 29691 4920 29747
rect 4976 29691 5001 29747
rect 5057 29691 5082 29747
rect 5138 29691 5163 29747
rect 2724 29667 5163 29691
rect 2724 29611 2733 29667
rect 2789 29611 2814 29667
rect 2870 29611 2895 29667
rect 2951 29611 2976 29667
rect 3032 29611 3057 29667
rect 3113 29611 3138 29667
rect 3194 29611 3219 29667
rect 3275 29611 3300 29667
rect 3356 29611 3381 29667
rect 3437 29611 3462 29667
rect 3518 29611 3543 29667
rect 3599 29611 3624 29667
rect 3680 29611 3705 29667
rect 3761 29611 3786 29667
rect 3842 29611 3867 29667
rect 3923 29611 3948 29667
rect 4004 29611 4029 29667
rect 4085 29611 4110 29667
rect 4166 29611 4191 29667
rect 4247 29611 4272 29667
rect 4328 29611 4353 29667
rect 4409 29611 4434 29667
rect 4490 29611 4515 29667
rect 4571 29611 4596 29667
rect 4652 29611 4677 29667
rect 4733 29611 4758 29667
rect 4814 29611 4839 29667
rect 4895 29611 4920 29667
rect 4976 29611 5001 29667
rect 5057 29611 5082 29667
rect 5138 29611 5163 29667
rect 2724 29587 5163 29611
rect 2724 29531 2733 29587
rect 2789 29531 2814 29587
rect 2870 29531 2895 29587
rect 2951 29531 2976 29587
rect 3032 29531 3057 29587
rect 3113 29531 3138 29587
rect 3194 29531 3219 29587
rect 3275 29531 3300 29587
rect 3356 29531 3381 29587
rect 3437 29531 3462 29587
rect 3518 29531 3543 29587
rect 3599 29531 3624 29587
rect 3680 29531 3705 29587
rect 3761 29531 3786 29587
rect 3842 29531 3867 29587
rect 3923 29531 3948 29587
rect 4004 29531 4029 29587
rect 4085 29531 4110 29587
rect 4166 29531 4191 29587
rect 4247 29531 4272 29587
rect 4328 29531 4353 29587
rect 4409 29531 4434 29587
rect 4490 29531 4515 29587
rect 4571 29531 4596 29587
rect 4652 29531 4677 29587
rect 4733 29531 4758 29587
rect 4814 29531 4839 29587
rect 4895 29531 4920 29587
rect 4976 29531 5001 29587
rect 5057 29531 5082 29587
rect 5138 29531 5163 29587
rect 2724 29507 5163 29531
rect 2724 29451 2733 29507
rect 2789 29451 2814 29507
rect 2870 29451 2895 29507
rect 2951 29451 2976 29507
rect 3032 29451 3057 29507
rect 3113 29451 3138 29507
rect 3194 29451 3219 29507
rect 3275 29451 3300 29507
rect 3356 29451 3381 29507
rect 3437 29451 3462 29507
rect 3518 29451 3543 29507
rect 3599 29451 3624 29507
rect 3680 29451 3705 29507
rect 3761 29451 3786 29507
rect 3842 29451 3867 29507
rect 3923 29451 3948 29507
rect 4004 29451 4029 29507
rect 4085 29451 4110 29507
rect 4166 29451 4191 29507
rect 4247 29451 4272 29507
rect 4328 29451 4353 29507
rect 4409 29451 4434 29507
rect 4490 29451 4515 29507
rect 4571 29451 4596 29507
rect 4652 29451 4677 29507
rect 4733 29451 4758 29507
rect 4814 29451 4839 29507
rect 4895 29451 4920 29507
rect 4976 29451 5001 29507
rect 5057 29451 5082 29507
rect 5138 29451 5163 29507
rect 2724 29427 5163 29451
rect 2724 29371 2733 29427
rect 2789 29371 2814 29427
rect 2870 29371 2895 29427
rect 2951 29371 2976 29427
rect 3032 29371 3057 29427
rect 3113 29371 3138 29427
rect 3194 29371 3219 29427
rect 3275 29371 3300 29427
rect 3356 29371 3381 29427
rect 3437 29371 3462 29427
rect 3518 29371 3543 29427
rect 3599 29371 3624 29427
rect 3680 29371 3705 29427
rect 3761 29371 3786 29427
rect 3842 29371 3867 29427
rect 3923 29371 3948 29427
rect 4004 29371 4029 29427
rect 4085 29371 4110 29427
rect 4166 29371 4191 29427
rect 4247 29371 4272 29427
rect 4328 29371 4353 29427
rect 4409 29371 4434 29427
rect 4490 29371 4515 29427
rect 4571 29371 4596 29427
rect 4652 29371 4677 29427
rect 4733 29371 4758 29427
rect 4814 29371 4839 29427
rect 4895 29371 4920 29427
rect 4976 29371 5001 29427
rect 5057 29371 5082 29427
rect 5138 29371 5163 29427
rect 5299 29371 5308 29987
rect 2724 27987 5308 29371
rect 2724 27931 2733 27987
rect 2789 27931 2814 27987
rect 2870 27931 2895 27987
rect 2951 27931 2976 27987
rect 3032 27931 3057 27987
rect 3113 27931 3138 27987
rect 3194 27931 3219 27987
rect 3275 27931 3300 27987
rect 3356 27931 3381 27987
rect 3437 27931 3462 27987
rect 3518 27931 3543 27987
rect 3599 27931 3624 27987
rect 3680 27931 3705 27987
rect 3761 27931 3786 27987
rect 3842 27931 3867 27987
rect 3923 27931 3948 27987
rect 4004 27931 4029 27987
rect 4085 27931 4110 27987
rect 4166 27931 4191 27987
rect 4247 27931 4272 27987
rect 4328 27931 4353 27987
rect 4409 27931 4434 27987
rect 4490 27931 4515 27987
rect 4571 27931 4596 27987
rect 4652 27931 4677 27987
rect 4733 27931 4758 27987
rect 4814 27931 4839 27987
rect 4895 27931 4920 27987
rect 4976 27931 5001 27987
rect 5057 27931 5082 27987
rect 5138 27931 5163 27987
rect 2724 27907 5163 27931
rect 2724 27851 2733 27907
rect 2789 27851 2814 27907
rect 2870 27851 2895 27907
rect 2951 27851 2976 27907
rect 3032 27851 3057 27907
rect 3113 27851 3138 27907
rect 3194 27851 3219 27907
rect 3275 27851 3300 27907
rect 3356 27851 3381 27907
rect 3437 27851 3462 27907
rect 3518 27851 3543 27907
rect 3599 27851 3624 27907
rect 3680 27851 3705 27907
rect 3761 27851 3786 27907
rect 3842 27851 3867 27907
rect 3923 27851 3948 27907
rect 4004 27851 4029 27907
rect 4085 27851 4110 27907
rect 4166 27851 4191 27907
rect 4247 27851 4272 27907
rect 4328 27851 4353 27907
rect 4409 27851 4434 27907
rect 4490 27851 4515 27907
rect 4571 27851 4596 27907
rect 4652 27851 4677 27907
rect 4733 27851 4758 27907
rect 4814 27851 4839 27907
rect 4895 27851 4920 27907
rect 4976 27851 5001 27907
rect 5057 27851 5082 27907
rect 5138 27851 5163 27907
rect 2724 27827 5163 27851
rect 2724 27771 2733 27827
rect 2789 27771 2814 27827
rect 2870 27771 2895 27827
rect 2951 27771 2976 27827
rect 3032 27771 3057 27827
rect 3113 27771 3138 27827
rect 3194 27771 3219 27827
rect 3275 27771 3300 27827
rect 3356 27771 3381 27827
rect 3437 27771 3462 27827
rect 3518 27771 3543 27827
rect 3599 27771 3624 27827
rect 3680 27771 3705 27827
rect 3761 27771 3786 27827
rect 3842 27771 3867 27827
rect 3923 27771 3948 27827
rect 4004 27771 4029 27827
rect 4085 27771 4110 27827
rect 4166 27771 4191 27827
rect 4247 27771 4272 27827
rect 4328 27771 4353 27827
rect 4409 27771 4434 27827
rect 4490 27771 4515 27827
rect 4571 27771 4596 27827
rect 4652 27771 4677 27827
rect 4733 27771 4758 27827
rect 4814 27771 4839 27827
rect 4895 27771 4920 27827
rect 4976 27771 5001 27827
rect 5057 27771 5082 27827
rect 5138 27771 5163 27827
rect 2724 27747 5163 27771
rect 2724 27691 2733 27747
rect 2789 27691 2814 27747
rect 2870 27691 2895 27747
rect 2951 27691 2976 27747
rect 3032 27691 3057 27747
rect 3113 27691 3138 27747
rect 3194 27691 3219 27747
rect 3275 27691 3300 27747
rect 3356 27691 3381 27747
rect 3437 27691 3462 27747
rect 3518 27691 3543 27747
rect 3599 27691 3624 27747
rect 3680 27691 3705 27747
rect 3761 27691 3786 27747
rect 3842 27691 3867 27747
rect 3923 27691 3948 27747
rect 4004 27691 4029 27747
rect 4085 27691 4110 27747
rect 4166 27691 4191 27747
rect 4247 27691 4272 27747
rect 4328 27691 4353 27747
rect 4409 27691 4434 27747
rect 4490 27691 4515 27747
rect 4571 27691 4596 27747
rect 4652 27691 4677 27747
rect 4733 27691 4758 27747
rect 4814 27691 4839 27747
rect 4895 27691 4920 27747
rect 4976 27691 5001 27747
rect 5057 27691 5082 27747
rect 5138 27691 5163 27747
rect 2724 27667 5163 27691
rect 2724 27611 2733 27667
rect 2789 27611 2814 27667
rect 2870 27611 2895 27667
rect 2951 27611 2976 27667
rect 3032 27611 3057 27667
rect 3113 27611 3138 27667
rect 3194 27611 3219 27667
rect 3275 27611 3300 27667
rect 3356 27611 3381 27667
rect 3437 27611 3462 27667
rect 3518 27611 3543 27667
rect 3599 27611 3624 27667
rect 3680 27611 3705 27667
rect 3761 27611 3786 27667
rect 3842 27611 3867 27667
rect 3923 27611 3948 27667
rect 4004 27611 4029 27667
rect 4085 27611 4110 27667
rect 4166 27611 4191 27667
rect 4247 27611 4272 27667
rect 4328 27611 4353 27667
rect 4409 27611 4434 27667
rect 4490 27611 4515 27667
rect 4571 27611 4596 27667
rect 4652 27611 4677 27667
rect 4733 27611 4758 27667
rect 4814 27611 4839 27667
rect 4895 27611 4920 27667
rect 4976 27611 5001 27667
rect 5057 27611 5082 27667
rect 5138 27611 5163 27667
rect 2724 27587 5163 27611
rect 2724 27531 2733 27587
rect 2789 27531 2814 27587
rect 2870 27531 2895 27587
rect 2951 27531 2976 27587
rect 3032 27531 3057 27587
rect 3113 27531 3138 27587
rect 3194 27531 3219 27587
rect 3275 27531 3300 27587
rect 3356 27531 3381 27587
rect 3437 27531 3462 27587
rect 3518 27531 3543 27587
rect 3599 27531 3624 27587
rect 3680 27531 3705 27587
rect 3761 27531 3786 27587
rect 3842 27531 3867 27587
rect 3923 27531 3948 27587
rect 4004 27531 4029 27587
rect 4085 27531 4110 27587
rect 4166 27531 4191 27587
rect 4247 27531 4272 27587
rect 4328 27531 4353 27587
rect 4409 27531 4434 27587
rect 4490 27531 4515 27587
rect 4571 27531 4596 27587
rect 4652 27531 4677 27587
rect 4733 27531 4758 27587
rect 4814 27531 4839 27587
rect 4895 27531 4920 27587
rect 4976 27531 5001 27587
rect 5057 27531 5082 27587
rect 5138 27531 5163 27587
rect 2724 27507 5163 27531
rect 2724 27451 2733 27507
rect 2789 27451 2814 27507
rect 2870 27451 2895 27507
rect 2951 27451 2976 27507
rect 3032 27451 3057 27507
rect 3113 27451 3138 27507
rect 3194 27451 3219 27507
rect 3275 27451 3300 27507
rect 3356 27451 3381 27507
rect 3437 27451 3462 27507
rect 3518 27451 3543 27507
rect 3599 27451 3624 27507
rect 3680 27451 3705 27507
rect 3761 27451 3786 27507
rect 3842 27451 3867 27507
rect 3923 27451 3948 27507
rect 4004 27451 4029 27507
rect 4085 27451 4110 27507
rect 4166 27451 4191 27507
rect 4247 27451 4272 27507
rect 4328 27451 4353 27507
rect 4409 27451 4434 27507
rect 4490 27451 4515 27507
rect 4571 27451 4596 27507
rect 4652 27451 4677 27507
rect 4733 27451 4758 27507
rect 4814 27451 4839 27507
rect 4895 27451 4920 27507
rect 4976 27451 5001 27507
rect 5057 27451 5082 27507
rect 5138 27451 5163 27507
rect 2724 27427 5163 27451
rect 2724 27371 2733 27427
rect 2789 27371 2814 27427
rect 2870 27371 2895 27427
rect 2951 27371 2976 27427
rect 3032 27371 3057 27427
rect 3113 27371 3138 27427
rect 3194 27371 3219 27427
rect 3275 27371 3300 27427
rect 3356 27371 3381 27427
rect 3437 27371 3462 27427
rect 3518 27371 3543 27427
rect 3599 27371 3624 27427
rect 3680 27371 3705 27427
rect 3761 27371 3786 27427
rect 3842 27371 3867 27427
rect 3923 27371 3948 27427
rect 4004 27371 4029 27427
rect 4085 27371 4110 27427
rect 4166 27371 4191 27427
rect 4247 27371 4272 27427
rect 4328 27371 4353 27427
rect 4409 27371 4434 27427
rect 4490 27371 4515 27427
rect 4571 27371 4596 27427
rect 4652 27371 4677 27427
rect 4733 27371 4758 27427
rect 4814 27371 4839 27427
rect 4895 27371 4920 27427
rect 4976 27371 5001 27427
rect 5057 27371 5082 27427
rect 5138 27371 5163 27427
rect 5299 27371 5308 27987
rect 2724 25987 5308 27371
rect 2724 25931 2733 25987
rect 2789 25931 2814 25987
rect 2870 25931 2895 25987
rect 2951 25931 2976 25987
rect 3032 25931 3057 25987
rect 3113 25931 3138 25987
rect 3194 25931 3219 25987
rect 3275 25931 3300 25987
rect 3356 25931 3381 25987
rect 3437 25931 3462 25987
rect 3518 25931 3543 25987
rect 3599 25931 3624 25987
rect 3680 25931 3705 25987
rect 3761 25931 3786 25987
rect 3842 25931 3867 25987
rect 3923 25931 3948 25987
rect 4004 25931 4029 25987
rect 4085 25931 4110 25987
rect 4166 25931 4191 25987
rect 4247 25931 4272 25987
rect 4328 25931 4353 25987
rect 4409 25931 4434 25987
rect 4490 25931 4515 25987
rect 4571 25931 4596 25987
rect 4652 25931 4677 25987
rect 4733 25931 4758 25987
rect 4814 25931 4839 25987
rect 4895 25931 4920 25987
rect 4976 25931 5001 25987
rect 5057 25931 5082 25987
rect 5138 25931 5163 25987
rect 2724 25907 5163 25931
rect 2724 25851 2733 25907
rect 2789 25851 2814 25907
rect 2870 25851 2895 25907
rect 2951 25851 2976 25907
rect 3032 25851 3057 25907
rect 3113 25851 3138 25907
rect 3194 25851 3219 25907
rect 3275 25851 3300 25907
rect 3356 25851 3381 25907
rect 3437 25851 3462 25907
rect 3518 25851 3543 25907
rect 3599 25851 3624 25907
rect 3680 25851 3705 25907
rect 3761 25851 3786 25907
rect 3842 25851 3867 25907
rect 3923 25851 3948 25907
rect 4004 25851 4029 25907
rect 4085 25851 4110 25907
rect 4166 25851 4191 25907
rect 4247 25851 4272 25907
rect 4328 25851 4353 25907
rect 4409 25851 4434 25907
rect 4490 25851 4515 25907
rect 4571 25851 4596 25907
rect 4652 25851 4677 25907
rect 4733 25851 4758 25907
rect 4814 25851 4839 25907
rect 4895 25851 4920 25907
rect 4976 25851 5001 25907
rect 5057 25851 5082 25907
rect 5138 25851 5163 25907
rect 2724 25827 5163 25851
rect 2724 25771 2733 25827
rect 2789 25771 2814 25827
rect 2870 25771 2895 25827
rect 2951 25771 2976 25827
rect 3032 25771 3057 25827
rect 3113 25771 3138 25827
rect 3194 25771 3219 25827
rect 3275 25771 3300 25827
rect 3356 25771 3381 25827
rect 3437 25771 3462 25827
rect 3518 25771 3543 25827
rect 3599 25771 3624 25827
rect 3680 25771 3705 25827
rect 3761 25771 3786 25827
rect 3842 25771 3867 25827
rect 3923 25771 3948 25827
rect 4004 25771 4029 25827
rect 4085 25771 4110 25827
rect 4166 25771 4191 25827
rect 4247 25771 4272 25827
rect 4328 25771 4353 25827
rect 4409 25771 4434 25827
rect 4490 25771 4515 25827
rect 4571 25771 4596 25827
rect 4652 25771 4677 25827
rect 4733 25771 4758 25827
rect 4814 25771 4839 25827
rect 4895 25771 4920 25827
rect 4976 25771 5001 25827
rect 5057 25771 5082 25827
rect 5138 25771 5163 25827
rect 2724 25747 5163 25771
rect 2724 25691 2733 25747
rect 2789 25691 2814 25747
rect 2870 25691 2895 25747
rect 2951 25691 2976 25747
rect 3032 25691 3057 25747
rect 3113 25691 3138 25747
rect 3194 25691 3219 25747
rect 3275 25691 3300 25747
rect 3356 25691 3381 25747
rect 3437 25691 3462 25747
rect 3518 25691 3543 25747
rect 3599 25691 3624 25747
rect 3680 25691 3705 25747
rect 3761 25691 3786 25747
rect 3842 25691 3867 25747
rect 3923 25691 3948 25747
rect 4004 25691 4029 25747
rect 4085 25691 4110 25747
rect 4166 25691 4191 25747
rect 4247 25691 4272 25747
rect 4328 25691 4353 25747
rect 4409 25691 4434 25747
rect 4490 25691 4515 25747
rect 4571 25691 4596 25747
rect 4652 25691 4677 25747
rect 4733 25691 4758 25747
rect 4814 25691 4839 25747
rect 4895 25691 4920 25747
rect 4976 25691 5001 25747
rect 5057 25691 5082 25747
rect 5138 25691 5163 25747
rect 2724 25667 5163 25691
rect 2724 25611 2733 25667
rect 2789 25611 2814 25667
rect 2870 25611 2895 25667
rect 2951 25611 2976 25667
rect 3032 25611 3057 25667
rect 3113 25611 3138 25667
rect 3194 25611 3219 25667
rect 3275 25611 3300 25667
rect 3356 25611 3381 25667
rect 3437 25611 3462 25667
rect 3518 25611 3543 25667
rect 3599 25611 3624 25667
rect 3680 25611 3705 25667
rect 3761 25611 3786 25667
rect 3842 25611 3867 25667
rect 3923 25611 3948 25667
rect 4004 25611 4029 25667
rect 4085 25611 4110 25667
rect 4166 25611 4191 25667
rect 4247 25611 4272 25667
rect 4328 25611 4353 25667
rect 4409 25611 4434 25667
rect 4490 25611 4515 25667
rect 4571 25611 4596 25667
rect 4652 25611 4677 25667
rect 4733 25611 4758 25667
rect 4814 25611 4839 25667
rect 4895 25611 4920 25667
rect 4976 25611 5001 25667
rect 5057 25611 5082 25667
rect 5138 25611 5163 25667
rect 2724 25587 5163 25611
rect 2724 25531 2733 25587
rect 2789 25531 2814 25587
rect 2870 25531 2895 25587
rect 2951 25531 2976 25587
rect 3032 25531 3057 25587
rect 3113 25531 3138 25587
rect 3194 25531 3219 25587
rect 3275 25531 3300 25587
rect 3356 25531 3381 25587
rect 3437 25531 3462 25587
rect 3518 25531 3543 25587
rect 3599 25531 3624 25587
rect 3680 25531 3705 25587
rect 3761 25531 3786 25587
rect 3842 25531 3867 25587
rect 3923 25531 3948 25587
rect 4004 25531 4029 25587
rect 4085 25531 4110 25587
rect 4166 25531 4191 25587
rect 4247 25531 4272 25587
rect 4328 25531 4353 25587
rect 4409 25531 4434 25587
rect 4490 25531 4515 25587
rect 4571 25531 4596 25587
rect 4652 25531 4677 25587
rect 4733 25531 4758 25587
rect 4814 25531 4839 25587
rect 4895 25531 4920 25587
rect 4976 25531 5001 25587
rect 5057 25531 5082 25587
rect 5138 25531 5163 25587
rect 2724 25507 5163 25531
rect 2724 25451 2733 25507
rect 2789 25451 2814 25507
rect 2870 25451 2895 25507
rect 2951 25451 2976 25507
rect 3032 25451 3057 25507
rect 3113 25451 3138 25507
rect 3194 25451 3219 25507
rect 3275 25451 3300 25507
rect 3356 25451 3381 25507
rect 3437 25451 3462 25507
rect 3518 25451 3543 25507
rect 3599 25451 3624 25507
rect 3680 25451 3705 25507
rect 3761 25451 3786 25507
rect 3842 25451 3867 25507
rect 3923 25451 3948 25507
rect 4004 25451 4029 25507
rect 4085 25451 4110 25507
rect 4166 25451 4191 25507
rect 4247 25451 4272 25507
rect 4328 25451 4353 25507
rect 4409 25451 4434 25507
rect 4490 25451 4515 25507
rect 4571 25451 4596 25507
rect 4652 25451 4677 25507
rect 4733 25451 4758 25507
rect 4814 25451 4839 25507
rect 4895 25451 4920 25507
rect 4976 25451 5001 25507
rect 5057 25451 5082 25507
rect 5138 25451 5163 25507
rect 2724 25427 5163 25451
rect 2724 25371 2733 25427
rect 2789 25371 2814 25427
rect 2870 25371 2895 25427
rect 2951 25371 2976 25427
rect 3032 25371 3057 25427
rect 3113 25371 3138 25427
rect 3194 25371 3219 25427
rect 3275 25371 3300 25427
rect 3356 25371 3381 25427
rect 3437 25371 3462 25427
rect 3518 25371 3543 25427
rect 3599 25371 3624 25427
rect 3680 25371 3705 25427
rect 3761 25371 3786 25427
rect 3842 25371 3867 25427
rect 3923 25371 3948 25427
rect 4004 25371 4029 25427
rect 4085 25371 4110 25427
rect 4166 25371 4191 25427
rect 4247 25371 4272 25427
rect 4328 25371 4353 25427
rect 4409 25371 4434 25427
rect 4490 25371 4515 25427
rect 4571 25371 4596 25427
rect 4652 25371 4677 25427
rect 4733 25371 4758 25427
rect 4814 25371 4839 25427
rect 4895 25371 4920 25427
rect 4976 25371 5001 25427
rect 5057 25371 5082 25427
rect 5138 25371 5163 25427
rect 5299 25371 5308 25987
rect 2724 23987 5308 25371
rect 2724 23931 2733 23987
rect 2789 23931 2814 23987
rect 2870 23931 2895 23987
rect 2951 23931 2976 23987
rect 3032 23931 3057 23987
rect 3113 23931 3138 23987
rect 3194 23931 3219 23987
rect 3275 23931 3300 23987
rect 3356 23931 3381 23987
rect 3437 23931 3462 23987
rect 3518 23931 3543 23987
rect 3599 23931 3624 23987
rect 3680 23931 3705 23987
rect 3761 23931 3786 23987
rect 3842 23931 3867 23987
rect 3923 23931 3948 23987
rect 4004 23931 4029 23987
rect 4085 23931 4110 23987
rect 4166 23931 4191 23987
rect 4247 23931 4272 23987
rect 4328 23931 4353 23987
rect 4409 23931 4434 23987
rect 4490 23931 4515 23987
rect 4571 23931 4596 23987
rect 4652 23931 4677 23987
rect 4733 23931 4758 23987
rect 4814 23931 4839 23987
rect 4895 23931 4920 23987
rect 4976 23931 5001 23987
rect 5057 23931 5082 23987
rect 5138 23931 5163 23987
rect 2724 23907 5163 23931
rect 2724 23851 2733 23907
rect 2789 23851 2814 23907
rect 2870 23851 2895 23907
rect 2951 23851 2976 23907
rect 3032 23851 3057 23907
rect 3113 23851 3138 23907
rect 3194 23851 3219 23907
rect 3275 23851 3300 23907
rect 3356 23851 3381 23907
rect 3437 23851 3462 23907
rect 3518 23851 3543 23907
rect 3599 23851 3624 23907
rect 3680 23851 3705 23907
rect 3761 23851 3786 23907
rect 3842 23851 3867 23907
rect 3923 23851 3948 23907
rect 4004 23851 4029 23907
rect 4085 23851 4110 23907
rect 4166 23851 4191 23907
rect 4247 23851 4272 23907
rect 4328 23851 4353 23907
rect 4409 23851 4434 23907
rect 4490 23851 4515 23907
rect 4571 23851 4596 23907
rect 4652 23851 4677 23907
rect 4733 23851 4758 23907
rect 4814 23851 4839 23907
rect 4895 23851 4920 23907
rect 4976 23851 5001 23907
rect 5057 23851 5082 23907
rect 5138 23851 5163 23907
rect 2724 23827 5163 23851
rect 2724 23771 2733 23827
rect 2789 23771 2814 23827
rect 2870 23771 2895 23827
rect 2951 23771 2976 23827
rect 3032 23771 3057 23827
rect 3113 23771 3138 23827
rect 3194 23771 3219 23827
rect 3275 23771 3300 23827
rect 3356 23771 3381 23827
rect 3437 23771 3462 23827
rect 3518 23771 3543 23827
rect 3599 23771 3624 23827
rect 3680 23771 3705 23827
rect 3761 23771 3786 23827
rect 3842 23771 3867 23827
rect 3923 23771 3948 23827
rect 4004 23771 4029 23827
rect 4085 23771 4110 23827
rect 4166 23771 4191 23827
rect 4247 23771 4272 23827
rect 4328 23771 4353 23827
rect 4409 23771 4434 23827
rect 4490 23771 4515 23827
rect 4571 23771 4596 23827
rect 4652 23771 4677 23827
rect 4733 23771 4758 23827
rect 4814 23771 4839 23827
rect 4895 23771 4920 23827
rect 4976 23771 5001 23827
rect 5057 23771 5082 23827
rect 5138 23771 5163 23827
rect 2724 23747 5163 23771
rect 2724 23691 2733 23747
rect 2789 23691 2814 23747
rect 2870 23691 2895 23747
rect 2951 23691 2976 23747
rect 3032 23691 3057 23747
rect 3113 23691 3138 23747
rect 3194 23691 3219 23747
rect 3275 23691 3300 23747
rect 3356 23691 3381 23747
rect 3437 23691 3462 23747
rect 3518 23691 3543 23747
rect 3599 23691 3624 23747
rect 3680 23691 3705 23747
rect 3761 23691 3786 23747
rect 3842 23691 3867 23747
rect 3923 23691 3948 23747
rect 4004 23691 4029 23747
rect 4085 23691 4110 23747
rect 4166 23691 4191 23747
rect 4247 23691 4272 23747
rect 4328 23691 4353 23747
rect 4409 23691 4434 23747
rect 4490 23691 4515 23747
rect 4571 23691 4596 23747
rect 4652 23691 4677 23747
rect 4733 23691 4758 23747
rect 4814 23691 4839 23747
rect 4895 23691 4920 23747
rect 4976 23691 5001 23747
rect 5057 23691 5082 23747
rect 5138 23691 5163 23747
rect 2724 23667 5163 23691
rect 2724 23611 2733 23667
rect 2789 23611 2814 23667
rect 2870 23611 2895 23667
rect 2951 23611 2976 23667
rect 3032 23611 3057 23667
rect 3113 23611 3138 23667
rect 3194 23611 3219 23667
rect 3275 23611 3300 23667
rect 3356 23611 3381 23667
rect 3437 23611 3462 23667
rect 3518 23611 3543 23667
rect 3599 23611 3624 23667
rect 3680 23611 3705 23667
rect 3761 23611 3786 23667
rect 3842 23611 3867 23667
rect 3923 23611 3948 23667
rect 4004 23611 4029 23667
rect 4085 23611 4110 23667
rect 4166 23611 4191 23667
rect 4247 23611 4272 23667
rect 4328 23611 4353 23667
rect 4409 23611 4434 23667
rect 4490 23611 4515 23667
rect 4571 23611 4596 23667
rect 4652 23611 4677 23667
rect 4733 23611 4758 23667
rect 4814 23611 4839 23667
rect 4895 23611 4920 23667
rect 4976 23611 5001 23667
rect 5057 23611 5082 23667
rect 5138 23611 5163 23667
rect 2724 23587 5163 23611
rect 2724 23531 2733 23587
rect 2789 23531 2814 23587
rect 2870 23531 2895 23587
rect 2951 23531 2976 23587
rect 3032 23531 3057 23587
rect 3113 23531 3138 23587
rect 3194 23531 3219 23587
rect 3275 23531 3300 23587
rect 3356 23531 3381 23587
rect 3437 23531 3462 23587
rect 3518 23531 3543 23587
rect 3599 23531 3624 23587
rect 3680 23531 3705 23587
rect 3761 23531 3786 23587
rect 3842 23531 3867 23587
rect 3923 23531 3948 23587
rect 4004 23531 4029 23587
rect 4085 23531 4110 23587
rect 4166 23531 4191 23587
rect 4247 23531 4272 23587
rect 4328 23531 4353 23587
rect 4409 23531 4434 23587
rect 4490 23531 4515 23587
rect 4571 23531 4596 23587
rect 4652 23531 4677 23587
rect 4733 23531 4758 23587
rect 4814 23531 4839 23587
rect 4895 23531 4920 23587
rect 4976 23531 5001 23587
rect 5057 23531 5082 23587
rect 5138 23531 5163 23587
rect 2724 23507 5163 23531
rect 2724 23451 2733 23507
rect 2789 23451 2814 23507
rect 2870 23451 2895 23507
rect 2951 23451 2976 23507
rect 3032 23451 3057 23507
rect 3113 23451 3138 23507
rect 3194 23451 3219 23507
rect 3275 23451 3300 23507
rect 3356 23451 3381 23507
rect 3437 23451 3462 23507
rect 3518 23451 3543 23507
rect 3599 23451 3624 23507
rect 3680 23451 3705 23507
rect 3761 23451 3786 23507
rect 3842 23451 3867 23507
rect 3923 23451 3948 23507
rect 4004 23451 4029 23507
rect 4085 23451 4110 23507
rect 4166 23451 4191 23507
rect 4247 23451 4272 23507
rect 4328 23451 4353 23507
rect 4409 23451 4434 23507
rect 4490 23451 4515 23507
rect 4571 23451 4596 23507
rect 4652 23451 4677 23507
rect 4733 23451 4758 23507
rect 4814 23451 4839 23507
rect 4895 23451 4920 23507
rect 4976 23451 5001 23507
rect 5057 23451 5082 23507
rect 5138 23451 5163 23507
rect 2724 23427 5163 23451
rect 2724 23371 2733 23427
rect 2789 23371 2814 23427
rect 2870 23371 2895 23427
rect 2951 23371 2976 23427
rect 3032 23371 3057 23427
rect 3113 23371 3138 23427
rect 3194 23371 3219 23427
rect 3275 23371 3300 23427
rect 3356 23371 3381 23427
rect 3437 23371 3462 23427
rect 3518 23371 3543 23427
rect 3599 23371 3624 23427
rect 3680 23371 3705 23427
rect 3761 23371 3786 23427
rect 3842 23371 3867 23427
rect 3923 23371 3948 23427
rect 4004 23371 4029 23427
rect 4085 23371 4110 23427
rect 4166 23371 4191 23427
rect 4247 23371 4272 23427
rect 4328 23371 4353 23427
rect 4409 23371 4434 23427
rect 4490 23371 4515 23427
rect 4571 23371 4596 23427
rect 4652 23371 4677 23427
rect 4733 23371 4758 23427
rect 4814 23371 4839 23427
rect 4895 23371 4920 23427
rect 4976 23371 5001 23427
rect 5057 23371 5082 23427
rect 5138 23371 5163 23427
rect 5299 23371 5308 23987
rect 2724 21987 5308 23371
rect 2724 21931 2733 21987
rect 2789 21931 2814 21987
rect 2870 21931 2895 21987
rect 2951 21931 2976 21987
rect 3032 21931 3057 21987
rect 3113 21931 3138 21987
rect 3194 21931 3219 21987
rect 3275 21931 3300 21987
rect 3356 21931 3381 21987
rect 3437 21931 3462 21987
rect 3518 21931 3543 21987
rect 3599 21931 3624 21987
rect 3680 21931 3705 21987
rect 3761 21931 3786 21987
rect 3842 21931 3867 21987
rect 3923 21931 3948 21987
rect 4004 21931 4029 21987
rect 4085 21931 4110 21987
rect 4166 21931 4191 21987
rect 4247 21931 4272 21987
rect 4328 21931 4353 21987
rect 4409 21931 4434 21987
rect 4490 21931 4515 21987
rect 4571 21931 4596 21987
rect 4652 21931 4677 21987
rect 4733 21931 4758 21987
rect 4814 21931 4839 21987
rect 4895 21931 4920 21987
rect 4976 21931 5001 21987
rect 5057 21931 5082 21987
rect 5138 21931 5163 21987
rect 2724 21907 5163 21931
rect 2724 21851 2733 21907
rect 2789 21851 2814 21907
rect 2870 21851 2895 21907
rect 2951 21851 2976 21907
rect 3032 21851 3057 21907
rect 3113 21851 3138 21907
rect 3194 21851 3219 21907
rect 3275 21851 3300 21907
rect 3356 21851 3381 21907
rect 3437 21851 3462 21907
rect 3518 21851 3543 21907
rect 3599 21851 3624 21907
rect 3680 21851 3705 21907
rect 3761 21851 3786 21907
rect 3842 21851 3867 21907
rect 3923 21851 3948 21907
rect 4004 21851 4029 21907
rect 4085 21851 4110 21907
rect 4166 21851 4191 21907
rect 4247 21851 4272 21907
rect 4328 21851 4353 21907
rect 4409 21851 4434 21907
rect 4490 21851 4515 21907
rect 4571 21851 4596 21907
rect 4652 21851 4677 21907
rect 4733 21851 4758 21907
rect 4814 21851 4839 21907
rect 4895 21851 4920 21907
rect 4976 21851 5001 21907
rect 5057 21851 5082 21907
rect 5138 21851 5163 21907
rect 2724 21827 5163 21851
rect 2724 21771 2733 21827
rect 2789 21771 2814 21827
rect 2870 21771 2895 21827
rect 2951 21771 2976 21827
rect 3032 21771 3057 21827
rect 3113 21771 3138 21827
rect 3194 21771 3219 21827
rect 3275 21771 3300 21827
rect 3356 21771 3381 21827
rect 3437 21771 3462 21827
rect 3518 21771 3543 21827
rect 3599 21771 3624 21827
rect 3680 21771 3705 21827
rect 3761 21771 3786 21827
rect 3842 21771 3867 21827
rect 3923 21771 3948 21827
rect 4004 21771 4029 21827
rect 4085 21771 4110 21827
rect 4166 21771 4191 21827
rect 4247 21771 4272 21827
rect 4328 21771 4353 21827
rect 4409 21771 4434 21827
rect 4490 21771 4515 21827
rect 4571 21771 4596 21827
rect 4652 21771 4677 21827
rect 4733 21771 4758 21827
rect 4814 21771 4839 21827
rect 4895 21771 4920 21827
rect 4976 21771 5001 21827
rect 5057 21771 5082 21827
rect 5138 21771 5163 21827
rect 2724 21747 5163 21771
rect 2724 21691 2733 21747
rect 2789 21691 2814 21747
rect 2870 21691 2895 21747
rect 2951 21691 2976 21747
rect 3032 21691 3057 21747
rect 3113 21691 3138 21747
rect 3194 21691 3219 21747
rect 3275 21691 3300 21747
rect 3356 21691 3381 21747
rect 3437 21691 3462 21747
rect 3518 21691 3543 21747
rect 3599 21691 3624 21747
rect 3680 21691 3705 21747
rect 3761 21691 3786 21747
rect 3842 21691 3867 21747
rect 3923 21691 3948 21747
rect 4004 21691 4029 21747
rect 4085 21691 4110 21747
rect 4166 21691 4191 21747
rect 4247 21691 4272 21747
rect 4328 21691 4353 21747
rect 4409 21691 4434 21747
rect 4490 21691 4515 21747
rect 4571 21691 4596 21747
rect 4652 21691 4677 21747
rect 4733 21691 4758 21747
rect 4814 21691 4839 21747
rect 4895 21691 4920 21747
rect 4976 21691 5001 21747
rect 5057 21691 5082 21747
rect 5138 21691 5163 21747
rect 2724 21667 5163 21691
rect 2724 21611 2733 21667
rect 2789 21611 2814 21667
rect 2870 21611 2895 21667
rect 2951 21611 2976 21667
rect 3032 21611 3057 21667
rect 3113 21611 3138 21667
rect 3194 21611 3219 21667
rect 3275 21611 3300 21667
rect 3356 21611 3381 21667
rect 3437 21611 3462 21667
rect 3518 21611 3543 21667
rect 3599 21611 3624 21667
rect 3680 21611 3705 21667
rect 3761 21611 3786 21667
rect 3842 21611 3867 21667
rect 3923 21611 3948 21667
rect 4004 21611 4029 21667
rect 4085 21611 4110 21667
rect 4166 21611 4191 21667
rect 4247 21611 4272 21667
rect 4328 21611 4353 21667
rect 4409 21611 4434 21667
rect 4490 21611 4515 21667
rect 4571 21611 4596 21667
rect 4652 21611 4677 21667
rect 4733 21611 4758 21667
rect 4814 21611 4839 21667
rect 4895 21611 4920 21667
rect 4976 21611 5001 21667
rect 5057 21611 5082 21667
rect 5138 21611 5163 21667
rect 2724 21587 5163 21611
rect 2724 21531 2733 21587
rect 2789 21531 2814 21587
rect 2870 21531 2895 21587
rect 2951 21531 2976 21587
rect 3032 21531 3057 21587
rect 3113 21531 3138 21587
rect 3194 21531 3219 21587
rect 3275 21531 3300 21587
rect 3356 21531 3381 21587
rect 3437 21531 3462 21587
rect 3518 21531 3543 21587
rect 3599 21531 3624 21587
rect 3680 21531 3705 21587
rect 3761 21531 3786 21587
rect 3842 21531 3867 21587
rect 3923 21531 3948 21587
rect 4004 21531 4029 21587
rect 4085 21531 4110 21587
rect 4166 21531 4191 21587
rect 4247 21531 4272 21587
rect 4328 21531 4353 21587
rect 4409 21531 4434 21587
rect 4490 21531 4515 21587
rect 4571 21531 4596 21587
rect 4652 21531 4677 21587
rect 4733 21531 4758 21587
rect 4814 21531 4839 21587
rect 4895 21531 4920 21587
rect 4976 21531 5001 21587
rect 5057 21531 5082 21587
rect 5138 21531 5163 21587
rect 2724 21507 5163 21531
rect 2724 21451 2733 21507
rect 2789 21451 2814 21507
rect 2870 21451 2895 21507
rect 2951 21451 2976 21507
rect 3032 21451 3057 21507
rect 3113 21451 3138 21507
rect 3194 21451 3219 21507
rect 3275 21451 3300 21507
rect 3356 21451 3381 21507
rect 3437 21451 3462 21507
rect 3518 21451 3543 21507
rect 3599 21451 3624 21507
rect 3680 21451 3705 21507
rect 3761 21451 3786 21507
rect 3842 21451 3867 21507
rect 3923 21451 3948 21507
rect 4004 21451 4029 21507
rect 4085 21451 4110 21507
rect 4166 21451 4191 21507
rect 4247 21451 4272 21507
rect 4328 21451 4353 21507
rect 4409 21451 4434 21507
rect 4490 21451 4515 21507
rect 4571 21451 4596 21507
rect 4652 21451 4677 21507
rect 4733 21451 4758 21507
rect 4814 21451 4839 21507
rect 4895 21451 4920 21507
rect 4976 21451 5001 21507
rect 5057 21451 5082 21507
rect 5138 21451 5163 21507
rect 2724 21427 5163 21451
rect 2724 21371 2733 21427
rect 2789 21371 2814 21427
rect 2870 21371 2895 21427
rect 2951 21371 2976 21427
rect 3032 21371 3057 21427
rect 3113 21371 3138 21427
rect 3194 21371 3219 21427
rect 3275 21371 3300 21427
rect 3356 21371 3381 21427
rect 3437 21371 3462 21427
rect 3518 21371 3543 21427
rect 3599 21371 3624 21427
rect 3680 21371 3705 21427
rect 3761 21371 3786 21427
rect 3842 21371 3867 21427
rect 3923 21371 3948 21427
rect 4004 21371 4029 21427
rect 4085 21371 4110 21427
rect 4166 21371 4191 21427
rect 4247 21371 4272 21427
rect 4328 21371 4353 21427
rect 4409 21371 4434 21427
rect 4490 21371 4515 21427
rect 4571 21371 4596 21427
rect 4652 21371 4677 21427
rect 4733 21371 4758 21427
rect 4814 21371 4839 21427
rect 4895 21371 4920 21427
rect 4976 21371 5001 21427
rect 5057 21371 5082 21427
rect 5138 21371 5163 21427
rect 5299 21371 5308 21987
rect 2724 19987 5308 21371
rect 2724 19931 2733 19987
rect 2789 19931 2814 19987
rect 2870 19931 2895 19987
rect 2951 19931 2976 19987
rect 3032 19931 3057 19987
rect 3113 19931 3138 19987
rect 3194 19931 3219 19987
rect 3275 19931 3300 19987
rect 3356 19931 3381 19987
rect 3437 19931 3462 19987
rect 3518 19931 3543 19987
rect 3599 19931 3624 19987
rect 3680 19931 3705 19987
rect 3761 19931 3786 19987
rect 3842 19931 3867 19987
rect 3923 19931 3948 19987
rect 4004 19931 4029 19987
rect 4085 19931 4110 19987
rect 4166 19931 4191 19987
rect 4247 19931 4272 19987
rect 4328 19931 4353 19987
rect 4409 19931 4434 19987
rect 4490 19931 4515 19987
rect 4571 19931 4596 19987
rect 4652 19931 4677 19987
rect 4733 19931 4758 19987
rect 4814 19931 4839 19987
rect 4895 19931 4920 19987
rect 4976 19931 5001 19987
rect 5057 19931 5082 19987
rect 5138 19931 5163 19987
rect 2724 19907 5163 19931
rect 2724 19851 2733 19907
rect 2789 19851 2814 19907
rect 2870 19851 2895 19907
rect 2951 19851 2976 19907
rect 3032 19851 3057 19907
rect 3113 19851 3138 19907
rect 3194 19851 3219 19907
rect 3275 19851 3300 19907
rect 3356 19851 3381 19907
rect 3437 19851 3462 19907
rect 3518 19851 3543 19907
rect 3599 19851 3624 19907
rect 3680 19851 3705 19907
rect 3761 19851 3786 19907
rect 3842 19851 3867 19907
rect 3923 19851 3948 19907
rect 4004 19851 4029 19907
rect 4085 19851 4110 19907
rect 4166 19851 4191 19907
rect 4247 19851 4272 19907
rect 4328 19851 4353 19907
rect 4409 19851 4434 19907
rect 4490 19851 4515 19907
rect 4571 19851 4596 19907
rect 4652 19851 4677 19907
rect 4733 19851 4758 19907
rect 4814 19851 4839 19907
rect 4895 19851 4920 19907
rect 4976 19851 5001 19907
rect 5057 19851 5082 19907
rect 5138 19851 5163 19907
rect 2724 19827 5163 19851
rect 2724 19771 2733 19827
rect 2789 19771 2814 19827
rect 2870 19771 2895 19827
rect 2951 19771 2976 19827
rect 3032 19771 3057 19827
rect 3113 19771 3138 19827
rect 3194 19771 3219 19827
rect 3275 19771 3300 19827
rect 3356 19771 3381 19827
rect 3437 19771 3462 19827
rect 3518 19771 3543 19827
rect 3599 19771 3624 19827
rect 3680 19771 3705 19827
rect 3761 19771 3786 19827
rect 3842 19771 3867 19827
rect 3923 19771 3948 19827
rect 4004 19771 4029 19827
rect 4085 19771 4110 19827
rect 4166 19771 4191 19827
rect 4247 19771 4272 19827
rect 4328 19771 4353 19827
rect 4409 19771 4434 19827
rect 4490 19771 4515 19827
rect 4571 19771 4596 19827
rect 4652 19771 4677 19827
rect 4733 19771 4758 19827
rect 4814 19771 4839 19827
rect 4895 19771 4920 19827
rect 4976 19771 5001 19827
rect 5057 19771 5082 19827
rect 5138 19771 5163 19827
rect 2724 19747 5163 19771
rect 2724 19691 2733 19747
rect 2789 19691 2814 19747
rect 2870 19691 2895 19747
rect 2951 19691 2976 19747
rect 3032 19691 3057 19747
rect 3113 19691 3138 19747
rect 3194 19691 3219 19747
rect 3275 19691 3300 19747
rect 3356 19691 3381 19747
rect 3437 19691 3462 19747
rect 3518 19691 3543 19747
rect 3599 19691 3624 19747
rect 3680 19691 3705 19747
rect 3761 19691 3786 19747
rect 3842 19691 3867 19747
rect 3923 19691 3948 19747
rect 4004 19691 4029 19747
rect 4085 19691 4110 19747
rect 4166 19691 4191 19747
rect 4247 19691 4272 19747
rect 4328 19691 4353 19747
rect 4409 19691 4434 19747
rect 4490 19691 4515 19747
rect 4571 19691 4596 19747
rect 4652 19691 4677 19747
rect 4733 19691 4758 19747
rect 4814 19691 4839 19747
rect 4895 19691 4920 19747
rect 4976 19691 5001 19747
rect 5057 19691 5082 19747
rect 5138 19691 5163 19747
rect 2724 19667 5163 19691
rect 2724 19611 2733 19667
rect 2789 19611 2814 19667
rect 2870 19611 2895 19667
rect 2951 19611 2976 19667
rect 3032 19611 3057 19667
rect 3113 19611 3138 19667
rect 3194 19611 3219 19667
rect 3275 19611 3300 19667
rect 3356 19611 3381 19667
rect 3437 19611 3462 19667
rect 3518 19611 3543 19667
rect 3599 19611 3624 19667
rect 3680 19611 3705 19667
rect 3761 19611 3786 19667
rect 3842 19611 3867 19667
rect 3923 19611 3948 19667
rect 4004 19611 4029 19667
rect 4085 19611 4110 19667
rect 4166 19611 4191 19667
rect 4247 19611 4272 19667
rect 4328 19611 4353 19667
rect 4409 19611 4434 19667
rect 4490 19611 4515 19667
rect 4571 19611 4596 19667
rect 4652 19611 4677 19667
rect 4733 19611 4758 19667
rect 4814 19611 4839 19667
rect 4895 19611 4920 19667
rect 4976 19611 5001 19667
rect 5057 19611 5082 19667
rect 5138 19611 5163 19667
rect 2724 19587 5163 19611
rect 2724 19531 2733 19587
rect 2789 19531 2814 19587
rect 2870 19531 2895 19587
rect 2951 19531 2976 19587
rect 3032 19531 3057 19587
rect 3113 19531 3138 19587
rect 3194 19531 3219 19587
rect 3275 19531 3300 19587
rect 3356 19531 3381 19587
rect 3437 19531 3462 19587
rect 3518 19531 3543 19587
rect 3599 19531 3624 19587
rect 3680 19531 3705 19587
rect 3761 19531 3786 19587
rect 3842 19531 3867 19587
rect 3923 19531 3948 19587
rect 4004 19531 4029 19587
rect 4085 19531 4110 19587
rect 4166 19531 4191 19587
rect 4247 19531 4272 19587
rect 4328 19531 4353 19587
rect 4409 19531 4434 19587
rect 4490 19531 4515 19587
rect 4571 19531 4596 19587
rect 4652 19531 4677 19587
rect 4733 19531 4758 19587
rect 4814 19531 4839 19587
rect 4895 19531 4920 19587
rect 4976 19531 5001 19587
rect 5057 19531 5082 19587
rect 5138 19531 5163 19587
rect 2724 19507 5163 19531
rect 2724 19451 2733 19507
rect 2789 19451 2814 19507
rect 2870 19451 2895 19507
rect 2951 19451 2976 19507
rect 3032 19451 3057 19507
rect 3113 19451 3138 19507
rect 3194 19451 3219 19507
rect 3275 19451 3300 19507
rect 3356 19451 3381 19507
rect 3437 19451 3462 19507
rect 3518 19451 3543 19507
rect 3599 19451 3624 19507
rect 3680 19451 3705 19507
rect 3761 19451 3786 19507
rect 3842 19451 3867 19507
rect 3923 19451 3948 19507
rect 4004 19451 4029 19507
rect 4085 19451 4110 19507
rect 4166 19451 4191 19507
rect 4247 19451 4272 19507
rect 4328 19451 4353 19507
rect 4409 19451 4434 19507
rect 4490 19451 4515 19507
rect 4571 19451 4596 19507
rect 4652 19451 4677 19507
rect 4733 19451 4758 19507
rect 4814 19451 4839 19507
rect 4895 19451 4920 19507
rect 4976 19451 5001 19507
rect 5057 19451 5082 19507
rect 5138 19451 5163 19507
rect 2724 19427 5163 19451
rect 2724 19371 2733 19427
rect 2789 19371 2814 19427
rect 2870 19371 2895 19427
rect 2951 19371 2976 19427
rect 3032 19371 3057 19427
rect 3113 19371 3138 19427
rect 3194 19371 3219 19427
rect 3275 19371 3300 19427
rect 3356 19371 3381 19427
rect 3437 19371 3462 19427
rect 3518 19371 3543 19427
rect 3599 19371 3624 19427
rect 3680 19371 3705 19427
rect 3761 19371 3786 19427
rect 3842 19371 3867 19427
rect 3923 19371 3948 19427
rect 4004 19371 4029 19427
rect 4085 19371 4110 19427
rect 4166 19371 4191 19427
rect 4247 19371 4272 19427
rect 4328 19371 4353 19427
rect 4409 19371 4434 19427
rect 4490 19371 4515 19427
rect 4571 19371 4596 19427
rect 4652 19371 4677 19427
rect 4733 19371 4758 19427
rect 4814 19371 4839 19427
rect 4895 19371 4920 19427
rect 4976 19371 5001 19427
rect 5057 19371 5082 19427
rect 5138 19371 5163 19427
rect 5299 19371 5308 19987
rect 2724 17987 5308 19371
rect 2724 17931 2733 17987
rect 2789 17931 2814 17987
rect 2870 17931 2895 17987
rect 2951 17931 2976 17987
rect 3032 17931 3057 17987
rect 3113 17931 3138 17987
rect 3194 17931 3219 17987
rect 3275 17931 3300 17987
rect 3356 17931 3381 17987
rect 3437 17931 3462 17987
rect 3518 17931 3543 17987
rect 3599 17931 3624 17987
rect 3680 17931 3705 17987
rect 3761 17931 3786 17987
rect 3842 17931 3867 17987
rect 3923 17931 3948 17987
rect 4004 17931 4029 17987
rect 4085 17931 4110 17987
rect 4166 17931 4191 17987
rect 4247 17931 4272 17987
rect 4328 17931 4353 17987
rect 4409 17931 4434 17987
rect 4490 17931 4515 17987
rect 4571 17931 4596 17987
rect 4652 17931 4677 17987
rect 4733 17931 4758 17987
rect 4814 17931 4839 17987
rect 4895 17931 4920 17987
rect 4976 17931 5001 17987
rect 5057 17931 5082 17987
rect 5138 17931 5163 17987
rect 2724 17907 5163 17931
rect 2724 17851 2733 17907
rect 2789 17851 2814 17907
rect 2870 17851 2895 17907
rect 2951 17851 2976 17907
rect 3032 17851 3057 17907
rect 3113 17851 3138 17907
rect 3194 17851 3219 17907
rect 3275 17851 3300 17907
rect 3356 17851 3381 17907
rect 3437 17851 3462 17907
rect 3518 17851 3543 17907
rect 3599 17851 3624 17907
rect 3680 17851 3705 17907
rect 3761 17851 3786 17907
rect 3842 17851 3867 17907
rect 3923 17851 3948 17907
rect 4004 17851 4029 17907
rect 4085 17851 4110 17907
rect 4166 17851 4191 17907
rect 4247 17851 4272 17907
rect 4328 17851 4353 17907
rect 4409 17851 4434 17907
rect 4490 17851 4515 17907
rect 4571 17851 4596 17907
rect 4652 17851 4677 17907
rect 4733 17851 4758 17907
rect 4814 17851 4839 17907
rect 4895 17851 4920 17907
rect 4976 17851 5001 17907
rect 5057 17851 5082 17907
rect 5138 17851 5163 17907
rect 2724 17827 5163 17851
rect 2724 17771 2733 17827
rect 2789 17771 2814 17827
rect 2870 17771 2895 17827
rect 2951 17771 2976 17827
rect 3032 17771 3057 17827
rect 3113 17771 3138 17827
rect 3194 17771 3219 17827
rect 3275 17771 3300 17827
rect 3356 17771 3381 17827
rect 3437 17771 3462 17827
rect 3518 17771 3543 17827
rect 3599 17771 3624 17827
rect 3680 17771 3705 17827
rect 3761 17771 3786 17827
rect 3842 17771 3867 17827
rect 3923 17771 3948 17827
rect 4004 17771 4029 17827
rect 4085 17771 4110 17827
rect 4166 17771 4191 17827
rect 4247 17771 4272 17827
rect 4328 17771 4353 17827
rect 4409 17771 4434 17827
rect 4490 17771 4515 17827
rect 4571 17771 4596 17827
rect 4652 17771 4677 17827
rect 4733 17771 4758 17827
rect 4814 17771 4839 17827
rect 4895 17771 4920 17827
rect 4976 17771 5001 17827
rect 5057 17771 5082 17827
rect 5138 17771 5163 17827
rect 2724 17747 5163 17771
rect 2724 17691 2733 17747
rect 2789 17691 2814 17747
rect 2870 17691 2895 17747
rect 2951 17691 2976 17747
rect 3032 17691 3057 17747
rect 3113 17691 3138 17747
rect 3194 17691 3219 17747
rect 3275 17691 3300 17747
rect 3356 17691 3381 17747
rect 3437 17691 3462 17747
rect 3518 17691 3543 17747
rect 3599 17691 3624 17747
rect 3680 17691 3705 17747
rect 3761 17691 3786 17747
rect 3842 17691 3867 17747
rect 3923 17691 3948 17747
rect 4004 17691 4029 17747
rect 4085 17691 4110 17747
rect 4166 17691 4191 17747
rect 4247 17691 4272 17747
rect 4328 17691 4353 17747
rect 4409 17691 4434 17747
rect 4490 17691 4515 17747
rect 4571 17691 4596 17747
rect 4652 17691 4677 17747
rect 4733 17691 4758 17747
rect 4814 17691 4839 17747
rect 4895 17691 4920 17747
rect 4976 17691 5001 17747
rect 5057 17691 5082 17747
rect 5138 17691 5163 17747
rect 2724 17667 5163 17691
rect 2724 17611 2733 17667
rect 2789 17611 2814 17667
rect 2870 17611 2895 17667
rect 2951 17611 2976 17667
rect 3032 17611 3057 17667
rect 3113 17611 3138 17667
rect 3194 17611 3219 17667
rect 3275 17611 3300 17667
rect 3356 17611 3381 17667
rect 3437 17611 3462 17667
rect 3518 17611 3543 17667
rect 3599 17611 3624 17667
rect 3680 17611 3705 17667
rect 3761 17611 3786 17667
rect 3842 17611 3867 17667
rect 3923 17611 3948 17667
rect 4004 17611 4029 17667
rect 4085 17611 4110 17667
rect 4166 17611 4191 17667
rect 4247 17611 4272 17667
rect 4328 17611 4353 17667
rect 4409 17611 4434 17667
rect 4490 17611 4515 17667
rect 4571 17611 4596 17667
rect 4652 17611 4677 17667
rect 4733 17611 4758 17667
rect 4814 17611 4839 17667
rect 4895 17611 4920 17667
rect 4976 17611 5001 17667
rect 5057 17611 5082 17667
rect 5138 17611 5163 17667
rect 2724 17587 5163 17611
rect 2724 17531 2733 17587
rect 2789 17531 2814 17587
rect 2870 17531 2895 17587
rect 2951 17531 2976 17587
rect 3032 17531 3057 17587
rect 3113 17531 3138 17587
rect 3194 17531 3219 17587
rect 3275 17531 3300 17587
rect 3356 17531 3381 17587
rect 3437 17531 3462 17587
rect 3518 17531 3543 17587
rect 3599 17531 3624 17587
rect 3680 17531 3705 17587
rect 3761 17531 3786 17587
rect 3842 17531 3867 17587
rect 3923 17531 3948 17587
rect 4004 17531 4029 17587
rect 4085 17531 4110 17587
rect 4166 17531 4191 17587
rect 4247 17531 4272 17587
rect 4328 17531 4353 17587
rect 4409 17531 4434 17587
rect 4490 17531 4515 17587
rect 4571 17531 4596 17587
rect 4652 17531 4677 17587
rect 4733 17531 4758 17587
rect 4814 17531 4839 17587
rect 4895 17531 4920 17587
rect 4976 17531 5001 17587
rect 5057 17531 5082 17587
rect 5138 17531 5163 17587
rect 2724 17507 5163 17531
rect 2724 17451 2733 17507
rect 2789 17451 2814 17507
rect 2870 17451 2895 17507
rect 2951 17451 2976 17507
rect 3032 17451 3057 17507
rect 3113 17451 3138 17507
rect 3194 17451 3219 17507
rect 3275 17451 3300 17507
rect 3356 17451 3381 17507
rect 3437 17451 3462 17507
rect 3518 17451 3543 17507
rect 3599 17451 3624 17507
rect 3680 17451 3705 17507
rect 3761 17451 3786 17507
rect 3842 17451 3867 17507
rect 3923 17451 3948 17507
rect 4004 17451 4029 17507
rect 4085 17451 4110 17507
rect 4166 17451 4191 17507
rect 4247 17451 4272 17507
rect 4328 17451 4353 17507
rect 4409 17451 4434 17507
rect 4490 17451 4515 17507
rect 4571 17451 4596 17507
rect 4652 17451 4677 17507
rect 4733 17451 4758 17507
rect 4814 17451 4839 17507
rect 4895 17451 4920 17507
rect 4976 17451 5001 17507
rect 5057 17451 5082 17507
rect 5138 17451 5163 17507
rect 2724 17427 5163 17451
rect 2724 17371 2733 17427
rect 2789 17371 2814 17427
rect 2870 17371 2895 17427
rect 2951 17371 2976 17427
rect 3032 17371 3057 17427
rect 3113 17371 3138 17427
rect 3194 17371 3219 17427
rect 3275 17371 3300 17427
rect 3356 17371 3381 17427
rect 3437 17371 3462 17427
rect 3518 17371 3543 17427
rect 3599 17371 3624 17427
rect 3680 17371 3705 17427
rect 3761 17371 3786 17427
rect 3842 17371 3867 17427
rect 3923 17371 3948 17427
rect 4004 17371 4029 17427
rect 4085 17371 4110 17427
rect 4166 17371 4191 17427
rect 4247 17371 4272 17427
rect 4328 17371 4353 17427
rect 4409 17371 4434 17427
rect 4490 17371 4515 17427
rect 4571 17371 4596 17427
rect 4652 17371 4677 17427
rect 4733 17371 4758 17427
rect 4814 17371 4839 17427
rect 4895 17371 4920 17427
rect 4976 17371 5001 17427
rect 5057 17371 5082 17427
rect 5138 17371 5163 17427
rect 5299 17371 5308 17987
rect 2724 14719 5308 17371
rect 2724 14663 2733 14719
rect 2789 14663 2814 14719
rect 2870 14663 2895 14719
rect 2951 14663 2976 14719
rect 3032 14663 3057 14719
rect 3113 14663 3138 14719
rect 3194 14663 3219 14719
rect 3275 14663 3300 14719
rect 3356 14663 3381 14719
rect 3437 14663 3462 14719
rect 3518 14663 3543 14719
rect 3599 14663 3624 14719
rect 3680 14663 3705 14719
rect 3761 14663 3786 14719
rect 3842 14663 3867 14719
rect 3923 14663 3948 14719
rect 4004 14663 4029 14719
rect 4085 14663 4110 14719
rect 4166 14663 4191 14719
rect 4247 14663 4272 14719
rect 4328 14663 4353 14719
rect 4409 14663 4434 14719
rect 4490 14663 4515 14719
rect 4571 14663 4596 14719
rect 4652 14663 4677 14719
rect 4733 14663 4758 14719
rect 4814 14663 4839 14719
rect 4895 14663 4920 14719
rect 4976 14663 5001 14719
rect 5057 14663 5082 14719
rect 5138 14663 5163 14719
rect 2724 14639 5163 14663
rect 2724 14583 2733 14639
rect 2789 14583 2814 14639
rect 2870 14583 2895 14639
rect 2951 14583 2976 14639
rect 3032 14583 3057 14639
rect 3113 14583 3138 14639
rect 3194 14583 3219 14639
rect 3275 14583 3300 14639
rect 3356 14583 3381 14639
rect 3437 14583 3462 14639
rect 3518 14583 3543 14639
rect 3599 14583 3624 14639
rect 3680 14583 3705 14639
rect 3761 14583 3786 14639
rect 3842 14583 3867 14639
rect 3923 14583 3948 14639
rect 4004 14583 4029 14639
rect 4085 14583 4110 14639
rect 4166 14583 4191 14639
rect 4247 14583 4272 14639
rect 4328 14583 4353 14639
rect 4409 14583 4434 14639
rect 4490 14583 4515 14639
rect 4571 14583 4596 14639
rect 4652 14583 4677 14639
rect 4733 14583 4758 14639
rect 4814 14583 4839 14639
rect 4895 14583 4920 14639
rect 4976 14583 5001 14639
rect 5057 14583 5082 14639
rect 5138 14583 5163 14639
rect 2724 14559 5163 14583
rect 2724 14503 2733 14559
rect 2789 14503 2814 14559
rect 2870 14503 2895 14559
rect 2951 14503 2976 14559
rect 3032 14503 3057 14559
rect 3113 14503 3138 14559
rect 3194 14503 3219 14559
rect 3275 14503 3300 14559
rect 3356 14503 3381 14559
rect 3437 14503 3462 14559
rect 3518 14503 3543 14559
rect 3599 14503 3624 14559
rect 3680 14503 3705 14559
rect 3761 14503 3786 14559
rect 3842 14503 3867 14559
rect 3923 14503 3948 14559
rect 4004 14503 4029 14559
rect 4085 14503 4110 14559
rect 4166 14503 4191 14559
rect 4247 14503 4272 14559
rect 4328 14503 4353 14559
rect 4409 14503 4434 14559
rect 4490 14503 4515 14559
rect 4571 14503 4596 14559
rect 4652 14503 4677 14559
rect 4733 14503 4758 14559
rect 4814 14503 4839 14559
rect 4895 14503 4920 14559
rect 4976 14503 5001 14559
rect 5057 14503 5082 14559
rect 5138 14503 5163 14559
rect 2724 14479 5163 14503
rect 2724 14423 2733 14479
rect 2789 14423 2814 14479
rect 2870 14423 2895 14479
rect 2951 14423 2976 14479
rect 3032 14423 3057 14479
rect 3113 14423 3138 14479
rect 3194 14423 3219 14479
rect 3275 14423 3300 14479
rect 3356 14423 3381 14479
rect 3437 14423 3462 14479
rect 3518 14423 3543 14479
rect 3599 14423 3624 14479
rect 3680 14423 3705 14479
rect 3761 14423 3786 14479
rect 3842 14423 3867 14479
rect 3923 14423 3948 14479
rect 4004 14423 4029 14479
rect 4085 14423 4110 14479
rect 4166 14423 4191 14479
rect 4247 14423 4272 14479
rect 4328 14423 4353 14479
rect 4409 14423 4434 14479
rect 4490 14423 4515 14479
rect 4571 14423 4596 14479
rect 4652 14423 4677 14479
rect 4733 14423 4758 14479
rect 4814 14423 4839 14479
rect 4895 14423 4920 14479
rect 4976 14423 5001 14479
rect 5057 14423 5082 14479
rect 5138 14423 5163 14479
rect 2724 14399 5163 14423
rect 2724 14343 2733 14399
rect 2789 14343 2814 14399
rect 2870 14343 2895 14399
rect 2951 14343 2976 14399
rect 3032 14343 3057 14399
rect 3113 14343 3138 14399
rect 3194 14343 3219 14399
rect 3275 14343 3300 14399
rect 3356 14343 3381 14399
rect 3437 14343 3462 14399
rect 3518 14343 3543 14399
rect 3599 14343 3624 14399
rect 3680 14343 3705 14399
rect 3761 14343 3786 14399
rect 3842 14343 3867 14399
rect 3923 14343 3948 14399
rect 4004 14343 4029 14399
rect 4085 14343 4110 14399
rect 4166 14343 4191 14399
rect 4247 14343 4272 14399
rect 4328 14343 4353 14399
rect 4409 14343 4434 14399
rect 4490 14343 4515 14399
rect 4571 14343 4596 14399
rect 4652 14343 4677 14399
rect 4733 14343 4758 14399
rect 4814 14343 4839 14399
rect 4895 14343 4920 14399
rect 4976 14343 5001 14399
rect 5057 14343 5082 14399
rect 5138 14343 5163 14399
rect 2724 14319 5163 14343
rect 2724 14263 2733 14319
rect 2789 14263 2814 14319
rect 2870 14263 2895 14319
rect 2951 14263 2976 14319
rect 3032 14263 3057 14319
rect 3113 14263 3138 14319
rect 3194 14263 3219 14319
rect 3275 14263 3300 14319
rect 3356 14263 3381 14319
rect 3437 14263 3462 14319
rect 3518 14263 3543 14319
rect 3599 14263 3624 14319
rect 3680 14263 3705 14319
rect 3761 14263 3786 14319
rect 3842 14263 3867 14319
rect 3923 14263 3948 14319
rect 4004 14263 4029 14319
rect 4085 14263 4110 14319
rect 4166 14263 4191 14319
rect 4247 14263 4272 14319
rect 4328 14263 4353 14319
rect 4409 14263 4434 14319
rect 4490 14263 4515 14319
rect 4571 14263 4596 14319
rect 4652 14263 4677 14319
rect 4733 14263 4758 14319
rect 4814 14263 4839 14319
rect 4895 14263 4920 14319
rect 4976 14263 5001 14319
rect 5057 14263 5082 14319
rect 5138 14263 5163 14319
rect 2724 14239 5163 14263
rect 2724 14183 2733 14239
rect 2789 14183 2814 14239
rect 2870 14183 2895 14239
rect 2951 14183 2976 14239
rect 3032 14183 3057 14239
rect 3113 14183 3138 14239
rect 3194 14183 3219 14239
rect 3275 14183 3300 14239
rect 3356 14183 3381 14239
rect 3437 14183 3462 14239
rect 3518 14183 3543 14239
rect 3599 14183 3624 14239
rect 3680 14183 3705 14239
rect 3761 14183 3786 14239
rect 3842 14183 3867 14239
rect 3923 14183 3948 14239
rect 4004 14183 4029 14239
rect 4085 14183 4110 14239
rect 4166 14183 4191 14239
rect 4247 14183 4272 14239
rect 4328 14183 4353 14239
rect 4409 14183 4434 14239
rect 4490 14183 4515 14239
rect 4571 14183 4596 14239
rect 4652 14183 4677 14239
rect 4733 14183 4758 14239
rect 4814 14183 4839 14239
rect 4895 14183 4920 14239
rect 4976 14183 5001 14239
rect 5057 14183 5082 14239
rect 5138 14183 5163 14239
rect 2724 14159 5163 14183
rect 2724 14103 2733 14159
rect 2789 14103 2814 14159
rect 2870 14103 2895 14159
rect 2951 14103 2976 14159
rect 3032 14103 3057 14159
rect 3113 14103 3138 14159
rect 3194 14103 3219 14159
rect 3275 14103 3300 14159
rect 3356 14103 3381 14159
rect 3437 14103 3462 14159
rect 3518 14103 3543 14159
rect 3599 14103 3624 14159
rect 3680 14103 3705 14159
rect 3761 14103 3786 14159
rect 3842 14103 3867 14159
rect 3923 14103 3948 14159
rect 4004 14103 4029 14159
rect 4085 14103 4110 14159
rect 4166 14103 4191 14159
rect 4247 14103 4272 14159
rect 4328 14103 4353 14159
rect 4409 14103 4434 14159
rect 4490 14103 4515 14159
rect 4571 14103 4596 14159
rect 4652 14103 4677 14159
rect 4733 14103 4758 14159
rect 4814 14103 4839 14159
rect 4895 14103 4920 14159
rect 4976 14103 5001 14159
rect 5057 14103 5082 14159
rect 5138 14103 5163 14159
rect 5299 14103 5308 14719
rect 2724 12719 5308 14103
rect 2724 12663 2733 12719
rect 2789 12663 2814 12719
rect 2870 12663 2895 12719
rect 2951 12663 2976 12719
rect 3032 12663 3057 12719
rect 3113 12663 3138 12719
rect 3194 12663 3219 12719
rect 3275 12663 3300 12719
rect 3356 12663 3381 12719
rect 3437 12663 3462 12719
rect 3518 12663 3543 12719
rect 3599 12663 3624 12719
rect 3680 12663 3705 12719
rect 3761 12663 3786 12719
rect 3842 12663 3867 12719
rect 3923 12663 3948 12719
rect 4004 12663 4029 12719
rect 4085 12663 4110 12719
rect 4166 12663 4191 12719
rect 4247 12663 4272 12719
rect 4328 12663 4353 12719
rect 4409 12663 4434 12719
rect 4490 12663 4515 12719
rect 4571 12663 4596 12719
rect 4652 12663 4677 12719
rect 4733 12663 4758 12719
rect 4814 12663 4839 12719
rect 4895 12663 4920 12719
rect 4976 12663 5001 12719
rect 5057 12663 5082 12719
rect 5138 12663 5163 12719
rect 2724 12639 5163 12663
rect 2724 12583 2733 12639
rect 2789 12583 2814 12639
rect 2870 12583 2895 12639
rect 2951 12583 2976 12639
rect 3032 12583 3057 12639
rect 3113 12583 3138 12639
rect 3194 12583 3219 12639
rect 3275 12583 3300 12639
rect 3356 12583 3381 12639
rect 3437 12583 3462 12639
rect 3518 12583 3543 12639
rect 3599 12583 3624 12639
rect 3680 12583 3705 12639
rect 3761 12583 3786 12639
rect 3842 12583 3867 12639
rect 3923 12583 3948 12639
rect 4004 12583 4029 12639
rect 4085 12583 4110 12639
rect 4166 12583 4191 12639
rect 4247 12583 4272 12639
rect 4328 12583 4353 12639
rect 4409 12583 4434 12639
rect 4490 12583 4515 12639
rect 4571 12583 4596 12639
rect 4652 12583 4677 12639
rect 4733 12583 4758 12639
rect 4814 12583 4839 12639
rect 4895 12583 4920 12639
rect 4976 12583 5001 12639
rect 5057 12583 5082 12639
rect 5138 12583 5163 12639
rect 2724 12559 5163 12583
rect 2724 12503 2733 12559
rect 2789 12503 2814 12559
rect 2870 12503 2895 12559
rect 2951 12503 2976 12559
rect 3032 12503 3057 12559
rect 3113 12503 3138 12559
rect 3194 12503 3219 12559
rect 3275 12503 3300 12559
rect 3356 12503 3381 12559
rect 3437 12503 3462 12559
rect 3518 12503 3543 12559
rect 3599 12503 3624 12559
rect 3680 12503 3705 12559
rect 3761 12503 3786 12559
rect 3842 12503 3867 12559
rect 3923 12503 3948 12559
rect 4004 12503 4029 12559
rect 4085 12503 4110 12559
rect 4166 12503 4191 12559
rect 4247 12503 4272 12559
rect 4328 12503 4353 12559
rect 4409 12503 4434 12559
rect 4490 12503 4515 12559
rect 4571 12503 4596 12559
rect 4652 12503 4677 12559
rect 4733 12503 4758 12559
rect 4814 12503 4839 12559
rect 4895 12503 4920 12559
rect 4976 12503 5001 12559
rect 5057 12503 5082 12559
rect 5138 12503 5163 12559
rect 2724 12479 5163 12503
rect 2724 12423 2733 12479
rect 2789 12423 2814 12479
rect 2870 12423 2895 12479
rect 2951 12423 2976 12479
rect 3032 12423 3057 12479
rect 3113 12423 3138 12479
rect 3194 12423 3219 12479
rect 3275 12423 3300 12479
rect 3356 12423 3381 12479
rect 3437 12423 3462 12479
rect 3518 12423 3543 12479
rect 3599 12423 3624 12479
rect 3680 12423 3705 12479
rect 3761 12423 3786 12479
rect 3842 12423 3867 12479
rect 3923 12423 3948 12479
rect 4004 12423 4029 12479
rect 4085 12423 4110 12479
rect 4166 12423 4191 12479
rect 4247 12423 4272 12479
rect 4328 12423 4353 12479
rect 4409 12423 4434 12479
rect 4490 12423 4515 12479
rect 4571 12423 4596 12479
rect 4652 12423 4677 12479
rect 4733 12423 4758 12479
rect 4814 12423 4839 12479
rect 4895 12423 4920 12479
rect 4976 12423 5001 12479
rect 5057 12423 5082 12479
rect 5138 12423 5163 12479
rect 2724 12399 5163 12423
rect 2724 12343 2733 12399
rect 2789 12343 2814 12399
rect 2870 12343 2895 12399
rect 2951 12343 2976 12399
rect 3032 12343 3057 12399
rect 3113 12343 3138 12399
rect 3194 12343 3219 12399
rect 3275 12343 3300 12399
rect 3356 12343 3381 12399
rect 3437 12343 3462 12399
rect 3518 12343 3543 12399
rect 3599 12343 3624 12399
rect 3680 12343 3705 12399
rect 3761 12343 3786 12399
rect 3842 12343 3867 12399
rect 3923 12343 3948 12399
rect 4004 12343 4029 12399
rect 4085 12343 4110 12399
rect 4166 12343 4191 12399
rect 4247 12343 4272 12399
rect 4328 12343 4353 12399
rect 4409 12343 4434 12399
rect 4490 12343 4515 12399
rect 4571 12343 4596 12399
rect 4652 12343 4677 12399
rect 4733 12343 4758 12399
rect 4814 12343 4839 12399
rect 4895 12343 4920 12399
rect 4976 12343 5001 12399
rect 5057 12343 5082 12399
rect 5138 12343 5163 12399
rect 2724 12319 5163 12343
rect 2724 12263 2733 12319
rect 2789 12263 2814 12319
rect 2870 12263 2895 12319
rect 2951 12263 2976 12319
rect 3032 12263 3057 12319
rect 3113 12263 3138 12319
rect 3194 12263 3219 12319
rect 3275 12263 3300 12319
rect 3356 12263 3381 12319
rect 3437 12263 3462 12319
rect 3518 12263 3543 12319
rect 3599 12263 3624 12319
rect 3680 12263 3705 12319
rect 3761 12263 3786 12319
rect 3842 12263 3867 12319
rect 3923 12263 3948 12319
rect 4004 12263 4029 12319
rect 4085 12263 4110 12319
rect 4166 12263 4191 12319
rect 4247 12263 4272 12319
rect 4328 12263 4353 12319
rect 4409 12263 4434 12319
rect 4490 12263 4515 12319
rect 4571 12263 4596 12319
rect 4652 12263 4677 12319
rect 4733 12263 4758 12319
rect 4814 12263 4839 12319
rect 4895 12263 4920 12319
rect 4976 12263 5001 12319
rect 5057 12263 5082 12319
rect 5138 12263 5163 12319
rect 2724 12239 5163 12263
rect 2724 12183 2733 12239
rect 2789 12183 2814 12239
rect 2870 12183 2895 12239
rect 2951 12183 2976 12239
rect 3032 12183 3057 12239
rect 3113 12183 3138 12239
rect 3194 12183 3219 12239
rect 3275 12183 3300 12239
rect 3356 12183 3381 12239
rect 3437 12183 3462 12239
rect 3518 12183 3543 12239
rect 3599 12183 3624 12239
rect 3680 12183 3705 12239
rect 3761 12183 3786 12239
rect 3842 12183 3867 12239
rect 3923 12183 3948 12239
rect 4004 12183 4029 12239
rect 4085 12183 4110 12239
rect 4166 12183 4191 12239
rect 4247 12183 4272 12239
rect 4328 12183 4353 12239
rect 4409 12183 4434 12239
rect 4490 12183 4515 12239
rect 4571 12183 4596 12239
rect 4652 12183 4677 12239
rect 4733 12183 4758 12239
rect 4814 12183 4839 12239
rect 4895 12183 4920 12239
rect 4976 12183 5001 12239
rect 5057 12183 5082 12239
rect 5138 12183 5163 12239
rect 2724 12159 5163 12183
rect 2724 12103 2733 12159
rect 2789 12103 2814 12159
rect 2870 12103 2895 12159
rect 2951 12103 2976 12159
rect 3032 12103 3057 12159
rect 3113 12103 3138 12159
rect 3194 12103 3219 12159
rect 3275 12103 3300 12159
rect 3356 12103 3381 12159
rect 3437 12103 3462 12159
rect 3518 12103 3543 12159
rect 3599 12103 3624 12159
rect 3680 12103 3705 12159
rect 3761 12103 3786 12159
rect 3842 12103 3867 12159
rect 3923 12103 3948 12159
rect 4004 12103 4029 12159
rect 4085 12103 4110 12159
rect 4166 12103 4191 12159
rect 4247 12103 4272 12159
rect 4328 12103 4353 12159
rect 4409 12103 4434 12159
rect 4490 12103 4515 12159
rect 4571 12103 4596 12159
rect 4652 12103 4677 12159
rect 4733 12103 4758 12159
rect 4814 12103 4839 12159
rect 4895 12103 4920 12159
rect 4976 12103 5001 12159
rect 5057 12103 5082 12159
rect 5138 12103 5163 12159
rect 5299 12103 5308 12719
rect 2724 10720 5308 12103
rect 2724 10664 2859 10720
rect 2915 10664 2942 10720
rect 2998 10664 3025 10720
rect 3081 10664 3108 10720
rect 3164 10664 3191 10720
rect 3247 10664 3274 10720
rect 3330 10664 3357 10720
rect 3413 10664 3439 10720
rect 3495 10664 3521 10720
rect 3577 10664 3603 10720
rect 3659 10664 3685 10720
rect 3741 10664 3767 10720
rect 3823 10664 3849 10720
rect 3905 10664 3931 10720
rect 3987 10664 4013 10720
rect 4069 10664 4095 10720
rect 4151 10664 4177 10720
rect 4233 10664 4259 10720
rect 4315 10664 4341 10720
rect 4397 10664 4423 10720
rect 4479 10664 4505 10720
rect 4561 10664 4587 10720
rect 4643 10664 4669 10720
rect 4725 10664 4751 10720
rect 4807 10664 4833 10720
rect 4889 10664 4915 10720
rect 4971 10664 4997 10720
rect 5053 10664 5079 10720
rect 5135 10664 5161 10720
rect 5217 10664 5243 10720
rect 5299 10664 5308 10720
rect 2724 10640 5308 10664
rect 2724 10584 2859 10640
rect 2915 10584 2942 10640
rect 2998 10584 3025 10640
rect 3081 10584 3108 10640
rect 3164 10584 3191 10640
rect 3247 10584 3274 10640
rect 3330 10584 3357 10640
rect 3413 10584 3439 10640
rect 3495 10584 3521 10640
rect 3577 10584 3603 10640
rect 3659 10584 3685 10640
rect 3741 10584 3767 10640
rect 3823 10584 3849 10640
rect 3905 10584 3931 10640
rect 3987 10584 4013 10640
rect 4069 10584 4095 10640
rect 4151 10584 4177 10640
rect 4233 10584 4259 10640
rect 4315 10584 4341 10640
rect 4397 10584 4423 10640
rect 4479 10584 4505 10640
rect 4561 10584 4587 10640
rect 4643 10584 4669 10640
rect 4725 10584 4751 10640
rect 4807 10584 4833 10640
rect 4889 10584 4915 10640
rect 4971 10584 4997 10640
rect 5053 10584 5079 10640
rect 5135 10584 5161 10640
rect 5217 10584 5243 10640
rect 5299 10584 5308 10640
rect 2724 10560 5308 10584
rect 2724 10504 2859 10560
rect 2915 10504 2942 10560
rect 2998 10504 3025 10560
rect 3081 10504 3108 10560
rect 3164 10504 3191 10560
rect 3247 10504 3274 10560
rect 3330 10504 3357 10560
rect 3413 10504 3439 10560
rect 3495 10504 3521 10560
rect 3577 10504 3603 10560
rect 3659 10504 3685 10560
rect 3741 10504 3767 10560
rect 3823 10504 3849 10560
rect 3905 10504 3931 10560
rect 3987 10504 4013 10560
rect 4069 10504 4095 10560
rect 4151 10504 4177 10560
rect 4233 10504 4259 10560
rect 4315 10504 4341 10560
rect 4397 10504 4423 10560
rect 4479 10504 4505 10560
rect 4561 10504 4587 10560
rect 4643 10504 4669 10560
rect 4725 10504 4751 10560
rect 4807 10504 4833 10560
rect 4889 10504 4915 10560
rect 4971 10504 4997 10560
rect 5053 10504 5079 10560
rect 5135 10504 5161 10560
rect 5217 10504 5243 10560
rect 5299 10504 5308 10560
rect 2724 10480 5308 10504
rect 2724 10424 2859 10480
rect 2915 10424 2942 10480
rect 2998 10424 3025 10480
rect 3081 10424 3108 10480
rect 3164 10424 3191 10480
rect 3247 10424 3274 10480
rect 3330 10424 3357 10480
rect 3413 10424 3439 10480
rect 3495 10424 3521 10480
rect 3577 10424 3603 10480
rect 3659 10424 3685 10480
rect 3741 10424 3767 10480
rect 3823 10424 3849 10480
rect 3905 10424 3931 10480
rect 3987 10424 4013 10480
rect 4069 10424 4095 10480
rect 4151 10424 4177 10480
rect 4233 10424 4259 10480
rect 4315 10424 4341 10480
rect 4397 10424 4423 10480
rect 4479 10424 4505 10480
rect 4561 10424 4587 10480
rect 4643 10424 4669 10480
rect 4725 10424 4751 10480
rect 4807 10424 4833 10480
rect 4889 10424 4915 10480
rect 4971 10424 4997 10480
rect 5053 10424 5079 10480
rect 5135 10424 5161 10480
rect 5217 10424 5243 10480
rect 5299 10424 5308 10480
rect 2724 10400 5308 10424
rect 2724 10344 2859 10400
rect 2915 10344 2942 10400
rect 2998 10344 3025 10400
rect 3081 10344 3108 10400
rect 3164 10344 3191 10400
rect 3247 10344 3274 10400
rect 3330 10344 3357 10400
rect 3413 10344 3439 10400
rect 3495 10344 3521 10400
rect 3577 10344 3603 10400
rect 3659 10344 3685 10400
rect 3741 10344 3767 10400
rect 3823 10344 3849 10400
rect 3905 10344 3931 10400
rect 3987 10344 4013 10400
rect 4069 10344 4095 10400
rect 4151 10344 4177 10400
rect 4233 10344 4259 10400
rect 4315 10344 4341 10400
rect 4397 10344 4423 10400
rect 4479 10344 4505 10400
rect 4561 10344 4587 10400
rect 4643 10344 4669 10400
rect 4725 10344 4751 10400
rect 4807 10344 4833 10400
rect 4889 10344 4915 10400
rect 4971 10344 4997 10400
rect 5053 10344 5079 10400
rect 5135 10344 5161 10400
rect 5217 10344 5243 10400
rect 5299 10344 5308 10400
rect 2724 10320 5308 10344
rect 2724 10264 2859 10320
rect 2915 10264 2942 10320
rect 2998 10264 3025 10320
rect 3081 10264 3108 10320
rect 3164 10264 3191 10320
rect 3247 10264 3274 10320
rect 3330 10264 3357 10320
rect 3413 10264 3439 10320
rect 3495 10264 3521 10320
rect 3577 10264 3603 10320
rect 3659 10264 3685 10320
rect 3741 10264 3767 10320
rect 3823 10264 3849 10320
rect 3905 10264 3931 10320
rect 3987 10264 4013 10320
rect 4069 10264 4095 10320
rect 4151 10264 4177 10320
rect 4233 10264 4259 10320
rect 4315 10264 4341 10320
rect 4397 10264 4423 10320
rect 4479 10264 4505 10320
rect 4561 10264 4587 10320
rect 4643 10264 4669 10320
rect 4725 10264 4751 10320
rect 4807 10264 4833 10320
rect 4889 10264 4915 10320
rect 4971 10264 4997 10320
rect 5053 10264 5079 10320
rect 5135 10264 5161 10320
rect 5217 10264 5243 10320
rect 5299 10264 5308 10320
rect 2724 10240 5308 10264
rect 2724 10184 2859 10240
rect 2915 10184 2942 10240
rect 2998 10184 3025 10240
rect 3081 10184 3108 10240
rect 3164 10184 3191 10240
rect 3247 10184 3274 10240
rect 3330 10184 3357 10240
rect 3413 10184 3439 10240
rect 3495 10184 3521 10240
rect 3577 10184 3603 10240
rect 3659 10184 3685 10240
rect 3741 10184 3767 10240
rect 3823 10184 3849 10240
rect 3905 10184 3931 10240
rect 3987 10184 4013 10240
rect 4069 10184 4095 10240
rect 4151 10184 4177 10240
rect 4233 10184 4259 10240
rect 4315 10184 4341 10240
rect 4397 10184 4423 10240
rect 4479 10184 4505 10240
rect 4561 10184 4587 10240
rect 4643 10184 4669 10240
rect 4725 10184 4751 10240
rect 4807 10184 4833 10240
rect 4889 10184 4915 10240
rect 4971 10184 4997 10240
rect 5053 10184 5079 10240
rect 5135 10184 5161 10240
rect 5217 10184 5243 10240
rect 5299 10184 5308 10240
rect 2724 10160 5308 10184
rect 2724 10104 2859 10160
rect 2915 10104 2942 10160
rect 2998 10104 3025 10160
rect 3081 10104 3108 10160
rect 3164 10104 3191 10160
rect 3247 10104 3274 10160
rect 3330 10104 3357 10160
rect 3413 10104 3439 10160
rect 3495 10104 3521 10160
rect 3577 10104 3603 10160
rect 3659 10104 3685 10160
rect 3741 10104 3767 10160
rect 3823 10104 3849 10160
rect 3905 10104 3931 10160
rect 3987 10104 4013 10160
rect 4069 10104 4095 10160
rect 4151 10104 4177 10160
rect 4233 10104 4259 10160
rect 4315 10104 4341 10160
rect 4397 10104 4423 10160
rect 4479 10104 4505 10160
rect 4561 10104 4587 10160
rect 4643 10104 4669 10160
rect 4725 10104 4751 10160
rect 4807 10104 4833 10160
rect 4889 10104 4915 10160
rect 4971 10104 4997 10160
rect 5053 10104 5079 10160
rect 5135 10104 5161 10160
rect 5217 10104 5243 10160
rect 5299 10104 5308 10160
rect 2724 2264 5308 10104
rect 2724 2208 3195 2264
rect 3251 2208 3277 2264
rect 3333 2208 3359 2264
rect 3415 2208 3441 2264
rect 3497 2208 3523 2264
rect 3579 2208 3605 2264
rect 3661 2208 3687 2264
rect 3743 2208 3769 2264
rect 3825 2208 3851 2264
rect 3907 2208 3933 2264
rect 3989 2208 4015 2264
rect 4071 2208 4097 2264
rect 4153 2208 4179 2264
rect 4235 2208 4261 2264
rect 4317 2208 4343 2264
rect 4399 2208 4425 2264
rect 4481 2208 4507 2264
rect 4563 2208 4589 2264
rect 4645 2208 4671 2264
rect 4727 2208 4753 2264
rect 4809 2208 4835 2264
rect 4891 2208 4917 2264
rect 4973 2208 4999 2264
rect 5055 2208 5080 2264
rect 5136 2208 5161 2264
rect 5217 2208 5242 2264
rect 5298 2208 5308 2264
rect 2724 2182 5308 2208
rect 2724 2126 3195 2182
rect 3251 2126 3277 2182
rect 3333 2126 3359 2182
rect 3415 2126 3441 2182
rect 3497 2126 3523 2182
rect 3579 2126 3605 2182
rect 3661 2126 3687 2182
rect 3743 2126 3769 2182
rect 3825 2126 3851 2182
rect 3907 2126 3933 2182
rect 3989 2126 4015 2182
rect 4071 2126 4097 2182
rect 4153 2126 4179 2182
rect 4235 2126 4261 2182
rect 4317 2126 4343 2182
rect 4399 2126 4425 2182
rect 4481 2126 4507 2182
rect 4563 2126 4589 2182
rect 4645 2126 4671 2182
rect 4727 2126 4753 2182
rect 4809 2126 4835 2182
rect 4891 2126 4917 2182
rect 4973 2126 4999 2182
rect 5055 2126 5080 2182
rect 5136 2126 5161 2182
rect 5217 2126 5242 2182
rect 5298 2126 5308 2182
rect 2724 2100 5308 2126
rect 2724 2044 3195 2100
rect 3251 2044 3277 2100
rect 3333 2044 3359 2100
rect 3415 2044 3441 2100
rect 3497 2044 3523 2100
rect 3579 2044 3605 2100
rect 3661 2044 3687 2100
rect 3743 2044 3769 2100
rect 3825 2044 3851 2100
rect 3907 2044 3933 2100
rect 3989 2044 4015 2100
rect 4071 2044 4097 2100
rect 4153 2044 4179 2100
rect 4235 2044 4261 2100
rect 4317 2044 4343 2100
rect 4399 2044 4425 2100
rect 4481 2044 4507 2100
rect 4563 2044 4589 2100
rect 4645 2044 4671 2100
rect 4727 2044 4753 2100
rect 4809 2044 4835 2100
rect 4891 2044 4917 2100
rect 4973 2044 4999 2100
rect 5055 2044 5080 2100
rect 5136 2044 5161 2100
rect 5217 2044 5242 2100
rect 5298 2044 5308 2100
rect 2724 2018 5308 2044
rect 2724 1962 3195 2018
rect 3251 1962 3277 2018
rect 3333 1962 3359 2018
rect 3415 1962 3441 2018
rect 3497 1962 3523 2018
rect 3579 1962 3605 2018
rect 3661 1962 3687 2018
rect 3743 1962 3769 2018
rect 3825 1962 3851 2018
rect 3907 1962 3933 2018
rect 3989 1962 4015 2018
rect 4071 1962 4097 2018
rect 4153 1962 4179 2018
rect 4235 1962 4261 2018
rect 4317 1962 4343 2018
rect 4399 1962 4425 2018
rect 4481 1962 4507 2018
rect 4563 1962 4589 2018
rect 4645 1962 4671 2018
rect 4727 1962 4753 2018
rect 4809 1962 4835 2018
rect 4891 1962 4917 2018
rect 4973 1962 4999 2018
rect 5055 1962 5080 2018
rect 5136 1962 5161 2018
rect 5217 1962 5242 2018
rect 5298 1962 5308 2018
rect 2724 1936 5308 1962
rect 2724 1880 3195 1936
rect 3251 1880 3277 1936
rect 3333 1880 3359 1936
rect 3415 1880 3441 1936
rect 3497 1880 3523 1936
rect 3579 1880 3605 1936
rect 3661 1880 3687 1936
rect 3743 1880 3769 1936
rect 3825 1880 3851 1936
rect 3907 1880 3933 1936
rect 3989 1880 4015 1936
rect 4071 1880 4097 1936
rect 4153 1880 4179 1936
rect 4235 1880 4261 1936
rect 4317 1880 4343 1936
rect 4399 1880 4425 1936
rect 4481 1880 4507 1936
rect 4563 1880 4589 1936
rect 4645 1880 4671 1936
rect 4727 1880 4753 1936
rect 4809 1880 4835 1936
rect 4891 1880 4917 1936
rect 4973 1880 4999 1936
rect 5055 1880 5080 1936
rect 5136 1880 5161 1936
rect 5217 1880 5242 1936
rect 5298 1880 5308 1936
rect 2724 0 5308 1880
rect 5608 36724 8218 38108
rect 5608 36668 5613 36724
rect 5669 36668 5696 36724
rect 5752 36668 5778 36724
rect 5834 36668 5860 36724
rect 5916 36668 5942 36724
rect 5998 36668 6024 36724
rect 6080 36668 6106 36724
rect 6162 36668 6188 36724
rect 6244 36668 6270 36724
rect 6326 36668 6352 36724
rect 6408 36668 6434 36724
rect 6490 36668 6516 36724
rect 6572 36668 6598 36724
rect 6654 36668 6680 36724
rect 6736 36668 6762 36724
rect 6818 36668 6844 36724
rect 6900 36668 6926 36724
rect 6982 36668 7008 36724
rect 7064 36668 7090 36724
rect 7146 36668 7172 36724
rect 7228 36668 7254 36724
rect 7310 36668 7336 36724
rect 7392 36668 7418 36724
rect 7474 36668 7500 36724
rect 7556 36668 7582 36724
rect 7638 36668 7664 36724
rect 7720 36668 7746 36724
rect 7802 36668 7828 36724
rect 7884 36668 7910 36724
rect 7966 36668 7992 36724
rect 8048 36668 8074 36724
rect 8130 36668 8156 36724
rect 8212 36668 8218 36724
rect 5608 36644 8218 36668
rect 5608 36588 5613 36644
rect 5669 36588 5696 36644
rect 5752 36588 5778 36644
rect 5834 36588 5860 36644
rect 5916 36588 5942 36644
rect 5998 36588 6024 36644
rect 6080 36588 6106 36644
rect 6162 36588 6188 36644
rect 6244 36588 6270 36644
rect 6326 36588 6352 36644
rect 6408 36588 6434 36644
rect 6490 36588 6516 36644
rect 6572 36588 6598 36644
rect 6654 36588 6680 36644
rect 6736 36588 6762 36644
rect 6818 36588 6844 36644
rect 6900 36588 6926 36644
rect 6982 36588 7008 36644
rect 7064 36588 7090 36644
rect 7146 36588 7172 36644
rect 7228 36588 7254 36644
rect 7310 36588 7336 36644
rect 7392 36588 7418 36644
rect 7474 36588 7500 36644
rect 7556 36588 7582 36644
rect 7638 36588 7664 36644
rect 7720 36588 7746 36644
rect 7802 36588 7828 36644
rect 7884 36588 7910 36644
rect 7966 36588 7992 36644
rect 8048 36588 8074 36644
rect 8130 36588 8156 36644
rect 8212 36588 8218 36644
rect 5608 36564 8218 36588
rect 5608 36508 5613 36564
rect 5669 36508 5696 36564
rect 5752 36508 5778 36564
rect 5834 36508 5860 36564
rect 5916 36508 5942 36564
rect 5998 36508 6024 36564
rect 6080 36508 6106 36564
rect 6162 36508 6188 36564
rect 6244 36508 6270 36564
rect 6326 36508 6352 36564
rect 6408 36508 6434 36564
rect 6490 36508 6516 36564
rect 6572 36508 6598 36564
rect 6654 36508 6680 36564
rect 6736 36508 6762 36564
rect 6818 36508 6844 36564
rect 6900 36508 6926 36564
rect 6982 36508 7008 36564
rect 7064 36508 7090 36564
rect 7146 36508 7172 36564
rect 7228 36508 7254 36564
rect 7310 36508 7336 36564
rect 7392 36508 7418 36564
rect 7474 36508 7500 36564
rect 7556 36508 7582 36564
rect 7638 36508 7664 36564
rect 7720 36508 7746 36564
rect 7802 36508 7828 36564
rect 7884 36508 7910 36564
rect 7966 36508 7992 36564
rect 8048 36508 8074 36564
rect 8130 36508 8156 36564
rect 8212 36508 8218 36564
rect 5608 36484 8218 36508
rect 5608 36428 5613 36484
rect 5669 36428 5696 36484
rect 5752 36428 5778 36484
rect 5834 36428 5860 36484
rect 5916 36428 5942 36484
rect 5998 36428 6024 36484
rect 6080 36428 6106 36484
rect 6162 36428 6188 36484
rect 6244 36428 6270 36484
rect 6326 36428 6352 36484
rect 6408 36428 6434 36484
rect 6490 36428 6516 36484
rect 6572 36428 6598 36484
rect 6654 36428 6680 36484
rect 6736 36428 6762 36484
rect 6818 36428 6844 36484
rect 6900 36428 6926 36484
rect 6982 36428 7008 36484
rect 7064 36428 7090 36484
rect 7146 36428 7172 36484
rect 7228 36428 7254 36484
rect 7310 36428 7336 36484
rect 7392 36428 7418 36484
rect 7474 36428 7500 36484
rect 7556 36428 7582 36484
rect 7638 36428 7664 36484
rect 7720 36428 7746 36484
rect 7802 36428 7828 36484
rect 7884 36428 7910 36484
rect 7966 36428 7992 36484
rect 8048 36428 8074 36484
rect 8130 36428 8156 36484
rect 8212 36428 8218 36484
rect 5608 36404 8218 36428
rect 5608 36348 5613 36404
rect 5669 36348 5696 36404
rect 5752 36348 5778 36404
rect 5834 36348 5860 36404
rect 5916 36348 5942 36404
rect 5998 36348 6024 36404
rect 6080 36348 6106 36404
rect 6162 36348 6188 36404
rect 6244 36348 6270 36404
rect 6326 36348 6352 36404
rect 6408 36348 6434 36404
rect 6490 36348 6516 36404
rect 6572 36348 6598 36404
rect 6654 36348 6680 36404
rect 6736 36348 6762 36404
rect 6818 36348 6844 36404
rect 6900 36348 6926 36404
rect 6982 36348 7008 36404
rect 7064 36348 7090 36404
rect 7146 36348 7172 36404
rect 7228 36348 7254 36404
rect 7310 36348 7336 36404
rect 7392 36348 7418 36404
rect 7474 36348 7500 36404
rect 7556 36348 7582 36404
rect 7638 36348 7664 36404
rect 7720 36348 7746 36404
rect 7802 36348 7828 36404
rect 7884 36348 7910 36404
rect 7966 36348 7992 36404
rect 8048 36348 8074 36404
rect 8130 36348 8156 36404
rect 8212 36348 8218 36404
rect 5608 36324 8218 36348
rect 5608 36268 5613 36324
rect 5669 36268 5696 36324
rect 5752 36268 5778 36324
rect 5834 36268 5860 36324
rect 5916 36268 5942 36324
rect 5998 36268 6024 36324
rect 6080 36268 6106 36324
rect 6162 36268 6188 36324
rect 6244 36268 6270 36324
rect 6326 36268 6352 36324
rect 6408 36268 6434 36324
rect 6490 36268 6516 36324
rect 6572 36268 6598 36324
rect 6654 36268 6680 36324
rect 6736 36268 6762 36324
rect 6818 36268 6844 36324
rect 6900 36268 6926 36324
rect 6982 36268 7008 36324
rect 7064 36268 7090 36324
rect 7146 36268 7172 36324
rect 7228 36268 7254 36324
rect 7310 36268 7336 36324
rect 7392 36268 7418 36324
rect 7474 36268 7500 36324
rect 7556 36268 7582 36324
rect 7638 36268 7664 36324
rect 7720 36268 7746 36324
rect 7802 36268 7828 36324
rect 7884 36268 7910 36324
rect 7966 36268 7992 36324
rect 8048 36268 8074 36324
rect 8130 36268 8156 36324
rect 8212 36268 8218 36324
rect 5608 36244 8218 36268
rect 5608 36188 5613 36244
rect 5669 36188 5696 36244
rect 5752 36188 5778 36244
rect 5834 36188 5860 36244
rect 5916 36188 5942 36244
rect 5998 36188 6024 36244
rect 6080 36188 6106 36244
rect 6162 36188 6188 36244
rect 6244 36188 6270 36244
rect 6326 36188 6352 36244
rect 6408 36188 6434 36244
rect 6490 36188 6516 36244
rect 6572 36188 6598 36244
rect 6654 36188 6680 36244
rect 6736 36188 6762 36244
rect 6818 36188 6844 36244
rect 6900 36188 6926 36244
rect 6982 36188 7008 36244
rect 7064 36188 7090 36244
rect 7146 36188 7172 36244
rect 7228 36188 7254 36244
rect 7310 36188 7336 36244
rect 7392 36188 7418 36244
rect 7474 36188 7500 36244
rect 7556 36188 7582 36244
rect 7638 36188 7664 36244
rect 7720 36188 7746 36244
rect 7802 36188 7828 36244
rect 7884 36188 7910 36244
rect 7966 36188 7992 36244
rect 8048 36188 8074 36244
rect 8130 36188 8156 36244
rect 8212 36188 8218 36244
rect 5608 36164 8218 36188
rect 5608 36108 5613 36164
rect 5669 36108 5696 36164
rect 5752 36108 5778 36164
rect 5834 36108 5860 36164
rect 5916 36108 5942 36164
rect 5998 36108 6024 36164
rect 6080 36108 6106 36164
rect 6162 36108 6188 36164
rect 6244 36108 6270 36164
rect 6326 36108 6352 36164
rect 6408 36108 6434 36164
rect 6490 36108 6516 36164
rect 6572 36108 6598 36164
rect 6654 36108 6680 36164
rect 6736 36108 6762 36164
rect 6818 36108 6844 36164
rect 6900 36108 6926 36164
rect 6982 36108 7008 36164
rect 7064 36108 7090 36164
rect 7146 36108 7172 36164
rect 7228 36108 7254 36164
rect 7310 36108 7336 36164
rect 7392 36108 7418 36164
rect 7474 36108 7500 36164
rect 7556 36108 7582 36164
rect 7638 36108 7664 36164
rect 7720 36108 7746 36164
rect 7802 36108 7828 36164
rect 7884 36108 7910 36164
rect 7966 36108 7992 36164
rect 8048 36108 8074 36164
rect 8130 36108 8156 36164
rect 8212 36108 8218 36164
rect 5608 34724 8218 36108
rect 5608 34668 5613 34724
rect 5669 34668 5696 34724
rect 5752 34668 5779 34724
rect 5835 34668 5861 34724
rect 5917 34668 5943 34724
rect 5999 34668 6025 34724
rect 6081 34668 6107 34724
rect 6163 34668 6189 34724
rect 6245 34668 6271 34724
rect 6327 34668 6353 34724
rect 6409 34668 6435 34724
rect 6491 34668 6517 34724
rect 6573 34668 6599 34724
rect 6655 34668 6681 34724
rect 6737 34668 6763 34724
rect 6819 34668 6845 34724
rect 6901 34668 6927 34724
rect 6983 34668 7009 34724
rect 7065 34668 7091 34724
rect 7147 34668 7173 34724
rect 7229 34668 7255 34724
rect 7311 34668 7337 34724
rect 7393 34668 7419 34724
rect 7475 34668 7501 34724
rect 7557 34668 7583 34724
rect 7639 34668 7665 34724
rect 7721 34668 7747 34724
rect 7803 34668 7829 34724
rect 7885 34668 7911 34724
rect 7967 34668 7993 34724
rect 8049 34668 8075 34724
rect 8131 34668 8157 34724
rect 8213 34668 8218 34724
rect 5608 34644 8218 34668
rect 5608 34588 5613 34644
rect 5669 34588 5696 34644
rect 5752 34588 5779 34644
rect 5835 34588 5861 34644
rect 5917 34588 5943 34644
rect 5999 34588 6025 34644
rect 6081 34588 6107 34644
rect 6163 34588 6189 34644
rect 6245 34588 6271 34644
rect 6327 34588 6353 34644
rect 6409 34588 6435 34644
rect 6491 34588 6517 34644
rect 6573 34588 6599 34644
rect 6655 34588 6681 34644
rect 6737 34588 6763 34644
rect 6819 34588 6845 34644
rect 6901 34588 6927 34644
rect 6983 34588 7009 34644
rect 7065 34588 7091 34644
rect 7147 34588 7173 34644
rect 7229 34588 7255 34644
rect 7311 34588 7337 34644
rect 7393 34588 7419 34644
rect 7475 34588 7501 34644
rect 7557 34588 7583 34644
rect 7639 34588 7665 34644
rect 7721 34588 7747 34644
rect 7803 34588 7829 34644
rect 7885 34588 7911 34644
rect 7967 34588 7993 34644
rect 8049 34588 8075 34644
rect 8131 34588 8157 34644
rect 8213 34588 8218 34644
rect 5608 34564 8218 34588
rect 5608 34508 5613 34564
rect 5669 34508 5696 34564
rect 5752 34508 5779 34564
rect 5835 34508 5861 34564
rect 5917 34508 5943 34564
rect 5999 34508 6025 34564
rect 6081 34508 6107 34564
rect 6163 34508 6189 34564
rect 6245 34508 6271 34564
rect 6327 34508 6353 34564
rect 6409 34508 6435 34564
rect 6491 34508 6517 34564
rect 6573 34508 6599 34564
rect 6655 34508 6681 34564
rect 6737 34508 6763 34564
rect 6819 34508 6845 34564
rect 6901 34508 6927 34564
rect 6983 34508 7009 34564
rect 7065 34508 7091 34564
rect 7147 34508 7173 34564
rect 7229 34508 7255 34564
rect 7311 34508 7337 34564
rect 7393 34508 7419 34564
rect 7475 34508 7501 34564
rect 7557 34508 7583 34564
rect 7639 34508 7665 34564
rect 7721 34508 7747 34564
rect 7803 34508 7829 34564
rect 7885 34508 7911 34564
rect 7967 34508 7993 34564
rect 8049 34508 8075 34564
rect 8131 34508 8157 34564
rect 8213 34508 8218 34564
rect 5608 34484 8218 34508
rect 5608 34428 5613 34484
rect 5669 34428 5696 34484
rect 5752 34428 5779 34484
rect 5835 34428 5861 34484
rect 5917 34428 5943 34484
rect 5999 34428 6025 34484
rect 6081 34428 6107 34484
rect 6163 34428 6189 34484
rect 6245 34428 6271 34484
rect 6327 34428 6353 34484
rect 6409 34428 6435 34484
rect 6491 34428 6517 34484
rect 6573 34428 6599 34484
rect 6655 34428 6681 34484
rect 6737 34428 6763 34484
rect 6819 34428 6845 34484
rect 6901 34428 6927 34484
rect 6983 34428 7009 34484
rect 7065 34428 7091 34484
rect 7147 34428 7173 34484
rect 7229 34428 7255 34484
rect 7311 34428 7337 34484
rect 7393 34428 7419 34484
rect 7475 34428 7501 34484
rect 7557 34428 7583 34484
rect 7639 34428 7665 34484
rect 7721 34428 7747 34484
rect 7803 34428 7829 34484
rect 7885 34428 7911 34484
rect 7967 34428 7993 34484
rect 8049 34428 8075 34484
rect 8131 34428 8157 34484
rect 8213 34428 8218 34484
rect 5608 34404 8218 34428
rect 5608 34348 5613 34404
rect 5669 34348 5696 34404
rect 5752 34348 5779 34404
rect 5835 34348 5861 34404
rect 5917 34348 5943 34404
rect 5999 34348 6025 34404
rect 6081 34348 6107 34404
rect 6163 34348 6189 34404
rect 6245 34348 6271 34404
rect 6327 34348 6353 34404
rect 6409 34348 6435 34404
rect 6491 34348 6517 34404
rect 6573 34348 6599 34404
rect 6655 34348 6681 34404
rect 6737 34348 6763 34404
rect 6819 34348 6845 34404
rect 6901 34348 6927 34404
rect 6983 34348 7009 34404
rect 7065 34348 7091 34404
rect 7147 34348 7173 34404
rect 7229 34348 7255 34404
rect 7311 34348 7337 34404
rect 7393 34348 7419 34404
rect 7475 34348 7501 34404
rect 7557 34348 7583 34404
rect 7639 34348 7665 34404
rect 7721 34348 7747 34404
rect 7803 34348 7829 34404
rect 7885 34348 7911 34404
rect 7967 34348 7993 34404
rect 8049 34348 8075 34404
rect 8131 34348 8157 34404
rect 8213 34348 8218 34404
rect 5608 34324 8218 34348
rect 5608 34268 5613 34324
rect 5669 34268 5696 34324
rect 5752 34268 5779 34324
rect 5835 34268 5861 34324
rect 5917 34268 5943 34324
rect 5999 34268 6025 34324
rect 6081 34268 6107 34324
rect 6163 34268 6189 34324
rect 6245 34268 6271 34324
rect 6327 34268 6353 34324
rect 6409 34268 6435 34324
rect 6491 34268 6517 34324
rect 6573 34268 6599 34324
rect 6655 34268 6681 34324
rect 6737 34268 6763 34324
rect 6819 34268 6845 34324
rect 6901 34268 6927 34324
rect 6983 34268 7009 34324
rect 7065 34268 7091 34324
rect 7147 34268 7173 34324
rect 7229 34268 7255 34324
rect 7311 34268 7337 34324
rect 7393 34268 7419 34324
rect 7475 34268 7501 34324
rect 7557 34268 7583 34324
rect 7639 34268 7665 34324
rect 7721 34268 7747 34324
rect 7803 34268 7829 34324
rect 7885 34268 7911 34324
rect 7967 34268 7993 34324
rect 8049 34268 8075 34324
rect 8131 34268 8157 34324
rect 8213 34268 8218 34324
rect 5608 34244 8218 34268
rect 5608 34188 5613 34244
rect 5669 34188 5696 34244
rect 5752 34188 5779 34244
rect 5835 34188 5861 34244
rect 5917 34188 5943 34244
rect 5999 34188 6025 34244
rect 6081 34188 6107 34244
rect 6163 34188 6189 34244
rect 6245 34188 6271 34244
rect 6327 34188 6353 34244
rect 6409 34188 6435 34244
rect 6491 34188 6517 34244
rect 6573 34188 6599 34244
rect 6655 34188 6681 34244
rect 6737 34188 6763 34244
rect 6819 34188 6845 34244
rect 6901 34188 6927 34244
rect 6983 34188 7009 34244
rect 7065 34188 7091 34244
rect 7147 34188 7173 34244
rect 7229 34188 7255 34244
rect 7311 34188 7337 34244
rect 7393 34188 7419 34244
rect 7475 34188 7501 34244
rect 7557 34188 7583 34244
rect 7639 34188 7665 34244
rect 7721 34188 7747 34244
rect 7803 34188 7829 34244
rect 7885 34188 7911 34244
rect 7967 34188 7993 34244
rect 8049 34188 8075 34244
rect 8131 34188 8157 34244
rect 8213 34188 8218 34244
rect 5608 34164 8218 34188
rect 5608 34108 5613 34164
rect 5669 34108 5696 34164
rect 5752 34108 5779 34164
rect 5835 34108 5861 34164
rect 5917 34108 5943 34164
rect 5999 34108 6025 34164
rect 6081 34108 6107 34164
rect 6163 34108 6189 34164
rect 6245 34108 6271 34164
rect 6327 34108 6353 34164
rect 6409 34108 6435 34164
rect 6491 34108 6517 34164
rect 6573 34108 6599 34164
rect 6655 34108 6681 34164
rect 6737 34108 6763 34164
rect 6819 34108 6845 34164
rect 6901 34108 6927 34164
rect 6983 34108 7009 34164
rect 7065 34108 7091 34164
rect 7147 34108 7173 34164
rect 7229 34108 7255 34164
rect 7311 34108 7337 34164
rect 7393 34108 7419 34164
rect 7475 34108 7501 34164
rect 7557 34108 7583 34164
rect 7639 34108 7665 34164
rect 7721 34108 7747 34164
rect 7803 34108 7829 34164
rect 7885 34108 7911 34164
rect 7967 34108 7993 34164
rect 8049 34108 8075 34164
rect 8131 34108 8157 34164
rect 8213 34108 8218 34164
rect 5608 32724 8218 34108
rect 5608 32668 5613 32724
rect 5669 32668 5696 32724
rect 5752 32668 5779 32724
rect 5835 32668 5861 32724
rect 5917 32668 5943 32724
rect 5999 32668 6025 32724
rect 6081 32668 6107 32724
rect 6163 32668 6189 32724
rect 6245 32668 6271 32724
rect 6327 32668 6353 32724
rect 6409 32668 6435 32724
rect 6491 32668 6517 32724
rect 6573 32668 6599 32724
rect 6655 32668 6681 32724
rect 6737 32668 6763 32724
rect 6819 32668 6845 32724
rect 6901 32668 6927 32724
rect 6983 32668 7009 32724
rect 7065 32668 7091 32724
rect 7147 32668 7173 32724
rect 7229 32668 7255 32724
rect 7311 32668 7337 32724
rect 7393 32668 7419 32724
rect 7475 32668 7501 32724
rect 7557 32668 7583 32724
rect 7639 32668 7665 32724
rect 7721 32668 7747 32724
rect 7803 32668 7829 32724
rect 7885 32668 7911 32724
rect 7967 32668 7993 32724
rect 8049 32668 8075 32724
rect 8131 32668 8157 32724
rect 8213 32668 8218 32724
rect 5608 32644 8218 32668
rect 5608 32588 5613 32644
rect 5669 32588 5696 32644
rect 5752 32588 5779 32644
rect 5835 32588 5861 32644
rect 5917 32588 5943 32644
rect 5999 32588 6025 32644
rect 6081 32588 6107 32644
rect 6163 32588 6189 32644
rect 6245 32588 6271 32644
rect 6327 32588 6353 32644
rect 6409 32588 6435 32644
rect 6491 32588 6517 32644
rect 6573 32588 6599 32644
rect 6655 32588 6681 32644
rect 6737 32588 6763 32644
rect 6819 32588 6845 32644
rect 6901 32588 6927 32644
rect 6983 32588 7009 32644
rect 7065 32588 7091 32644
rect 7147 32588 7173 32644
rect 7229 32588 7255 32644
rect 7311 32588 7337 32644
rect 7393 32588 7419 32644
rect 7475 32588 7501 32644
rect 7557 32588 7583 32644
rect 7639 32588 7665 32644
rect 7721 32588 7747 32644
rect 7803 32588 7829 32644
rect 7885 32588 7911 32644
rect 7967 32588 7993 32644
rect 8049 32588 8075 32644
rect 8131 32588 8157 32644
rect 8213 32588 8218 32644
rect 5608 32564 8218 32588
rect 5608 32508 5613 32564
rect 5669 32508 5696 32564
rect 5752 32508 5779 32564
rect 5835 32508 5861 32564
rect 5917 32508 5943 32564
rect 5999 32508 6025 32564
rect 6081 32508 6107 32564
rect 6163 32508 6189 32564
rect 6245 32508 6271 32564
rect 6327 32508 6353 32564
rect 6409 32508 6435 32564
rect 6491 32508 6517 32564
rect 6573 32508 6599 32564
rect 6655 32508 6681 32564
rect 6737 32508 6763 32564
rect 6819 32508 6845 32564
rect 6901 32508 6927 32564
rect 6983 32508 7009 32564
rect 7065 32508 7091 32564
rect 7147 32508 7173 32564
rect 7229 32508 7255 32564
rect 7311 32508 7337 32564
rect 7393 32508 7419 32564
rect 7475 32508 7501 32564
rect 7557 32508 7583 32564
rect 7639 32508 7665 32564
rect 7721 32508 7747 32564
rect 7803 32508 7829 32564
rect 7885 32508 7911 32564
rect 7967 32508 7993 32564
rect 8049 32508 8075 32564
rect 8131 32508 8157 32564
rect 8213 32508 8218 32564
rect 5608 32484 8218 32508
rect 5608 32428 5613 32484
rect 5669 32428 5696 32484
rect 5752 32428 5779 32484
rect 5835 32428 5861 32484
rect 5917 32428 5943 32484
rect 5999 32428 6025 32484
rect 6081 32428 6107 32484
rect 6163 32428 6189 32484
rect 6245 32428 6271 32484
rect 6327 32428 6353 32484
rect 6409 32428 6435 32484
rect 6491 32428 6517 32484
rect 6573 32428 6599 32484
rect 6655 32428 6681 32484
rect 6737 32428 6763 32484
rect 6819 32428 6845 32484
rect 6901 32428 6927 32484
rect 6983 32428 7009 32484
rect 7065 32428 7091 32484
rect 7147 32428 7173 32484
rect 7229 32428 7255 32484
rect 7311 32428 7337 32484
rect 7393 32428 7419 32484
rect 7475 32428 7501 32484
rect 7557 32428 7583 32484
rect 7639 32428 7665 32484
rect 7721 32428 7747 32484
rect 7803 32428 7829 32484
rect 7885 32428 7911 32484
rect 7967 32428 7993 32484
rect 8049 32428 8075 32484
rect 8131 32428 8157 32484
rect 8213 32428 8218 32484
rect 5608 32404 8218 32428
rect 5608 32348 5613 32404
rect 5669 32348 5696 32404
rect 5752 32348 5779 32404
rect 5835 32348 5861 32404
rect 5917 32348 5943 32404
rect 5999 32348 6025 32404
rect 6081 32348 6107 32404
rect 6163 32348 6189 32404
rect 6245 32348 6271 32404
rect 6327 32348 6353 32404
rect 6409 32348 6435 32404
rect 6491 32348 6517 32404
rect 6573 32348 6599 32404
rect 6655 32348 6681 32404
rect 6737 32348 6763 32404
rect 6819 32348 6845 32404
rect 6901 32348 6927 32404
rect 6983 32348 7009 32404
rect 7065 32348 7091 32404
rect 7147 32348 7173 32404
rect 7229 32348 7255 32404
rect 7311 32348 7337 32404
rect 7393 32348 7419 32404
rect 7475 32348 7501 32404
rect 7557 32348 7583 32404
rect 7639 32348 7665 32404
rect 7721 32348 7747 32404
rect 7803 32348 7829 32404
rect 7885 32348 7911 32404
rect 7967 32348 7993 32404
rect 8049 32348 8075 32404
rect 8131 32348 8157 32404
rect 8213 32348 8218 32404
rect 5608 32324 8218 32348
rect 5608 32268 5613 32324
rect 5669 32268 5696 32324
rect 5752 32268 5779 32324
rect 5835 32268 5861 32324
rect 5917 32268 5943 32324
rect 5999 32268 6025 32324
rect 6081 32268 6107 32324
rect 6163 32268 6189 32324
rect 6245 32268 6271 32324
rect 6327 32268 6353 32324
rect 6409 32268 6435 32324
rect 6491 32268 6517 32324
rect 6573 32268 6599 32324
rect 6655 32268 6681 32324
rect 6737 32268 6763 32324
rect 6819 32268 6845 32324
rect 6901 32268 6927 32324
rect 6983 32268 7009 32324
rect 7065 32268 7091 32324
rect 7147 32268 7173 32324
rect 7229 32268 7255 32324
rect 7311 32268 7337 32324
rect 7393 32268 7419 32324
rect 7475 32268 7501 32324
rect 7557 32268 7583 32324
rect 7639 32268 7665 32324
rect 7721 32268 7747 32324
rect 7803 32268 7829 32324
rect 7885 32268 7911 32324
rect 7967 32268 7993 32324
rect 8049 32268 8075 32324
rect 8131 32268 8157 32324
rect 8213 32268 8218 32324
rect 5608 32244 8218 32268
rect 5608 32188 5613 32244
rect 5669 32188 5696 32244
rect 5752 32188 5779 32244
rect 5835 32188 5861 32244
rect 5917 32188 5943 32244
rect 5999 32188 6025 32244
rect 6081 32188 6107 32244
rect 6163 32188 6189 32244
rect 6245 32188 6271 32244
rect 6327 32188 6353 32244
rect 6409 32188 6435 32244
rect 6491 32188 6517 32244
rect 6573 32188 6599 32244
rect 6655 32188 6681 32244
rect 6737 32188 6763 32244
rect 6819 32188 6845 32244
rect 6901 32188 6927 32244
rect 6983 32188 7009 32244
rect 7065 32188 7091 32244
rect 7147 32188 7173 32244
rect 7229 32188 7255 32244
rect 7311 32188 7337 32244
rect 7393 32188 7419 32244
rect 7475 32188 7501 32244
rect 7557 32188 7583 32244
rect 7639 32188 7665 32244
rect 7721 32188 7747 32244
rect 7803 32188 7829 32244
rect 7885 32188 7911 32244
rect 7967 32188 7993 32244
rect 8049 32188 8075 32244
rect 8131 32188 8157 32244
rect 8213 32188 8218 32244
rect 5608 32164 8218 32188
rect 5608 32108 5613 32164
rect 5669 32108 5696 32164
rect 5752 32108 5779 32164
rect 5835 32108 5861 32164
rect 5917 32108 5943 32164
rect 5999 32108 6025 32164
rect 6081 32108 6107 32164
rect 6163 32108 6189 32164
rect 6245 32108 6271 32164
rect 6327 32108 6353 32164
rect 6409 32108 6435 32164
rect 6491 32108 6517 32164
rect 6573 32108 6599 32164
rect 6655 32108 6681 32164
rect 6737 32108 6763 32164
rect 6819 32108 6845 32164
rect 6901 32108 6927 32164
rect 6983 32108 7009 32164
rect 7065 32108 7091 32164
rect 7147 32108 7173 32164
rect 7229 32108 7255 32164
rect 7311 32108 7337 32164
rect 7393 32108 7419 32164
rect 7475 32108 7501 32164
rect 7557 32108 7583 32164
rect 7639 32108 7665 32164
rect 7721 32108 7747 32164
rect 7803 32108 7829 32164
rect 7885 32108 7911 32164
rect 7967 32108 7993 32164
rect 8049 32108 8075 32164
rect 8131 32108 8157 32164
rect 8213 32108 8218 32164
rect 5608 30724 8218 32108
rect 5608 30668 5613 30724
rect 5669 30668 5696 30724
rect 5752 30668 5779 30724
rect 5835 30668 5861 30724
rect 5917 30668 5943 30724
rect 5999 30668 6025 30724
rect 6081 30668 6107 30724
rect 6163 30668 6189 30724
rect 6245 30668 6271 30724
rect 6327 30668 6353 30724
rect 6409 30668 6435 30724
rect 6491 30668 6517 30724
rect 6573 30668 6599 30724
rect 6655 30668 6681 30724
rect 6737 30668 6763 30724
rect 6819 30668 6845 30724
rect 6901 30668 6927 30724
rect 6983 30668 7009 30724
rect 7065 30668 7091 30724
rect 7147 30668 7173 30724
rect 7229 30668 7255 30724
rect 7311 30668 7337 30724
rect 7393 30668 7419 30724
rect 7475 30668 7501 30724
rect 7557 30668 7583 30724
rect 7639 30668 7665 30724
rect 7721 30668 7747 30724
rect 7803 30668 7829 30724
rect 7885 30668 7911 30724
rect 7967 30668 7993 30724
rect 8049 30668 8075 30724
rect 8131 30668 8157 30724
rect 8213 30668 8218 30724
rect 5608 30644 8218 30668
rect 5608 30588 5613 30644
rect 5669 30588 5696 30644
rect 5752 30588 5779 30644
rect 5835 30588 5861 30644
rect 5917 30588 5943 30644
rect 5999 30588 6025 30644
rect 6081 30588 6107 30644
rect 6163 30588 6189 30644
rect 6245 30588 6271 30644
rect 6327 30588 6353 30644
rect 6409 30588 6435 30644
rect 6491 30588 6517 30644
rect 6573 30588 6599 30644
rect 6655 30588 6681 30644
rect 6737 30588 6763 30644
rect 6819 30588 6845 30644
rect 6901 30588 6927 30644
rect 6983 30588 7009 30644
rect 7065 30588 7091 30644
rect 7147 30588 7173 30644
rect 7229 30588 7255 30644
rect 7311 30588 7337 30644
rect 7393 30588 7419 30644
rect 7475 30588 7501 30644
rect 7557 30588 7583 30644
rect 7639 30588 7665 30644
rect 7721 30588 7747 30644
rect 7803 30588 7829 30644
rect 7885 30588 7911 30644
rect 7967 30588 7993 30644
rect 8049 30588 8075 30644
rect 8131 30588 8157 30644
rect 8213 30588 8218 30644
rect 5608 30564 8218 30588
rect 5608 30508 5613 30564
rect 5669 30508 5696 30564
rect 5752 30508 5779 30564
rect 5835 30508 5861 30564
rect 5917 30508 5943 30564
rect 5999 30508 6025 30564
rect 6081 30508 6107 30564
rect 6163 30508 6189 30564
rect 6245 30508 6271 30564
rect 6327 30508 6353 30564
rect 6409 30508 6435 30564
rect 6491 30508 6517 30564
rect 6573 30508 6599 30564
rect 6655 30508 6681 30564
rect 6737 30508 6763 30564
rect 6819 30508 6845 30564
rect 6901 30508 6927 30564
rect 6983 30508 7009 30564
rect 7065 30508 7091 30564
rect 7147 30508 7173 30564
rect 7229 30508 7255 30564
rect 7311 30508 7337 30564
rect 7393 30508 7419 30564
rect 7475 30508 7501 30564
rect 7557 30508 7583 30564
rect 7639 30508 7665 30564
rect 7721 30508 7747 30564
rect 7803 30508 7829 30564
rect 7885 30508 7911 30564
rect 7967 30508 7993 30564
rect 8049 30508 8075 30564
rect 8131 30508 8157 30564
rect 8213 30508 8218 30564
rect 5608 30484 8218 30508
rect 5608 30428 5613 30484
rect 5669 30428 5696 30484
rect 5752 30428 5779 30484
rect 5835 30428 5861 30484
rect 5917 30428 5943 30484
rect 5999 30428 6025 30484
rect 6081 30428 6107 30484
rect 6163 30428 6189 30484
rect 6245 30428 6271 30484
rect 6327 30428 6353 30484
rect 6409 30428 6435 30484
rect 6491 30428 6517 30484
rect 6573 30428 6599 30484
rect 6655 30428 6681 30484
rect 6737 30428 6763 30484
rect 6819 30428 6845 30484
rect 6901 30428 6927 30484
rect 6983 30428 7009 30484
rect 7065 30428 7091 30484
rect 7147 30428 7173 30484
rect 7229 30428 7255 30484
rect 7311 30428 7337 30484
rect 7393 30428 7419 30484
rect 7475 30428 7501 30484
rect 7557 30428 7583 30484
rect 7639 30428 7665 30484
rect 7721 30428 7747 30484
rect 7803 30428 7829 30484
rect 7885 30428 7911 30484
rect 7967 30428 7993 30484
rect 8049 30428 8075 30484
rect 8131 30428 8157 30484
rect 8213 30428 8218 30484
rect 5608 30404 8218 30428
rect 5608 30348 5613 30404
rect 5669 30348 5696 30404
rect 5752 30348 5779 30404
rect 5835 30348 5861 30404
rect 5917 30348 5943 30404
rect 5999 30348 6025 30404
rect 6081 30348 6107 30404
rect 6163 30348 6189 30404
rect 6245 30348 6271 30404
rect 6327 30348 6353 30404
rect 6409 30348 6435 30404
rect 6491 30348 6517 30404
rect 6573 30348 6599 30404
rect 6655 30348 6681 30404
rect 6737 30348 6763 30404
rect 6819 30348 6845 30404
rect 6901 30348 6927 30404
rect 6983 30348 7009 30404
rect 7065 30348 7091 30404
rect 7147 30348 7173 30404
rect 7229 30348 7255 30404
rect 7311 30348 7337 30404
rect 7393 30348 7419 30404
rect 7475 30348 7501 30404
rect 7557 30348 7583 30404
rect 7639 30348 7665 30404
rect 7721 30348 7747 30404
rect 7803 30348 7829 30404
rect 7885 30348 7911 30404
rect 7967 30348 7993 30404
rect 8049 30348 8075 30404
rect 8131 30348 8157 30404
rect 8213 30348 8218 30404
rect 5608 30324 8218 30348
rect 5608 30268 5613 30324
rect 5669 30268 5696 30324
rect 5752 30268 5779 30324
rect 5835 30268 5861 30324
rect 5917 30268 5943 30324
rect 5999 30268 6025 30324
rect 6081 30268 6107 30324
rect 6163 30268 6189 30324
rect 6245 30268 6271 30324
rect 6327 30268 6353 30324
rect 6409 30268 6435 30324
rect 6491 30268 6517 30324
rect 6573 30268 6599 30324
rect 6655 30268 6681 30324
rect 6737 30268 6763 30324
rect 6819 30268 6845 30324
rect 6901 30268 6927 30324
rect 6983 30268 7009 30324
rect 7065 30268 7091 30324
rect 7147 30268 7173 30324
rect 7229 30268 7255 30324
rect 7311 30268 7337 30324
rect 7393 30268 7419 30324
rect 7475 30268 7501 30324
rect 7557 30268 7583 30324
rect 7639 30268 7665 30324
rect 7721 30268 7747 30324
rect 7803 30268 7829 30324
rect 7885 30268 7911 30324
rect 7967 30268 7993 30324
rect 8049 30268 8075 30324
rect 8131 30268 8157 30324
rect 8213 30268 8218 30324
rect 5608 30244 8218 30268
rect 5608 30188 5613 30244
rect 5669 30188 5696 30244
rect 5752 30188 5779 30244
rect 5835 30188 5861 30244
rect 5917 30188 5943 30244
rect 5999 30188 6025 30244
rect 6081 30188 6107 30244
rect 6163 30188 6189 30244
rect 6245 30188 6271 30244
rect 6327 30188 6353 30244
rect 6409 30188 6435 30244
rect 6491 30188 6517 30244
rect 6573 30188 6599 30244
rect 6655 30188 6681 30244
rect 6737 30188 6763 30244
rect 6819 30188 6845 30244
rect 6901 30188 6927 30244
rect 6983 30188 7009 30244
rect 7065 30188 7091 30244
rect 7147 30188 7173 30244
rect 7229 30188 7255 30244
rect 7311 30188 7337 30244
rect 7393 30188 7419 30244
rect 7475 30188 7501 30244
rect 7557 30188 7583 30244
rect 7639 30188 7665 30244
rect 7721 30188 7747 30244
rect 7803 30188 7829 30244
rect 7885 30188 7911 30244
rect 7967 30188 7993 30244
rect 8049 30188 8075 30244
rect 8131 30188 8157 30244
rect 8213 30188 8218 30244
rect 5608 30164 8218 30188
rect 5608 30108 5613 30164
rect 5669 30108 5696 30164
rect 5752 30108 5779 30164
rect 5835 30108 5861 30164
rect 5917 30108 5943 30164
rect 5999 30108 6025 30164
rect 6081 30108 6107 30164
rect 6163 30108 6189 30164
rect 6245 30108 6271 30164
rect 6327 30108 6353 30164
rect 6409 30108 6435 30164
rect 6491 30108 6517 30164
rect 6573 30108 6599 30164
rect 6655 30108 6681 30164
rect 6737 30108 6763 30164
rect 6819 30108 6845 30164
rect 6901 30108 6927 30164
rect 6983 30108 7009 30164
rect 7065 30108 7091 30164
rect 7147 30108 7173 30164
rect 7229 30108 7255 30164
rect 7311 30108 7337 30164
rect 7393 30108 7419 30164
rect 7475 30108 7501 30164
rect 7557 30108 7583 30164
rect 7639 30108 7665 30164
rect 7721 30108 7747 30164
rect 7803 30108 7829 30164
rect 7885 30108 7911 30164
rect 7967 30108 7993 30164
rect 8049 30108 8075 30164
rect 8131 30108 8157 30164
rect 8213 30108 8218 30164
rect 5608 28724 8218 30108
rect 5608 28668 5613 28724
rect 5669 28668 5696 28724
rect 5752 28668 5779 28724
rect 5835 28668 5861 28724
rect 5917 28668 5943 28724
rect 5999 28668 6025 28724
rect 6081 28668 6107 28724
rect 6163 28668 6189 28724
rect 6245 28668 6271 28724
rect 6327 28668 6353 28724
rect 6409 28668 6435 28724
rect 6491 28668 6517 28724
rect 6573 28668 6599 28724
rect 6655 28668 6681 28724
rect 6737 28668 6763 28724
rect 6819 28668 6845 28724
rect 6901 28668 6927 28724
rect 6983 28668 7009 28724
rect 7065 28668 7091 28724
rect 7147 28668 7173 28724
rect 7229 28668 7255 28724
rect 7311 28668 7337 28724
rect 7393 28668 7419 28724
rect 7475 28668 7501 28724
rect 7557 28668 7583 28724
rect 7639 28668 7665 28724
rect 7721 28668 7747 28724
rect 7803 28668 7829 28724
rect 7885 28668 7911 28724
rect 7967 28668 7993 28724
rect 8049 28668 8075 28724
rect 8131 28668 8157 28724
rect 8213 28668 8218 28724
rect 5608 28644 8218 28668
rect 5608 28588 5613 28644
rect 5669 28588 5696 28644
rect 5752 28588 5779 28644
rect 5835 28588 5861 28644
rect 5917 28588 5943 28644
rect 5999 28588 6025 28644
rect 6081 28588 6107 28644
rect 6163 28588 6189 28644
rect 6245 28588 6271 28644
rect 6327 28588 6353 28644
rect 6409 28588 6435 28644
rect 6491 28588 6517 28644
rect 6573 28588 6599 28644
rect 6655 28588 6681 28644
rect 6737 28588 6763 28644
rect 6819 28588 6845 28644
rect 6901 28588 6927 28644
rect 6983 28588 7009 28644
rect 7065 28588 7091 28644
rect 7147 28588 7173 28644
rect 7229 28588 7255 28644
rect 7311 28588 7337 28644
rect 7393 28588 7419 28644
rect 7475 28588 7501 28644
rect 7557 28588 7583 28644
rect 7639 28588 7665 28644
rect 7721 28588 7747 28644
rect 7803 28588 7829 28644
rect 7885 28588 7911 28644
rect 7967 28588 7993 28644
rect 8049 28588 8075 28644
rect 8131 28588 8157 28644
rect 8213 28588 8218 28644
rect 5608 28564 8218 28588
rect 5608 28508 5613 28564
rect 5669 28508 5696 28564
rect 5752 28508 5779 28564
rect 5835 28508 5861 28564
rect 5917 28508 5943 28564
rect 5999 28508 6025 28564
rect 6081 28508 6107 28564
rect 6163 28508 6189 28564
rect 6245 28508 6271 28564
rect 6327 28508 6353 28564
rect 6409 28508 6435 28564
rect 6491 28508 6517 28564
rect 6573 28508 6599 28564
rect 6655 28508 6681 28564
rect 6737 28508 6763 28564
rect 6819 28508 6845 28564
rect 6901 28508 6927 28564
rect 6983 28508 7009 28564
rect 7065 28508 7091 28564
rect 7147 28508 7173 28564
rect 7229 28508 7255 28564
rect 7311 28508 7337 28564
rect 7393 28508 7419 28564
rect 7475 28508 7501 28564
rect 7557 28508 7583 28564
rect 7639 28508 7665 28564
rect 7721 28508 7747 28564
rect 7803 28508 7829 28564
rect 7885 28508 7911 28564
rect 7967 28508 7993 28564
rect 8049 28508 8075 28564
rect 8131 28508 8157 28564
rect 8213 28508 8218 28564
rect 5608 28484 8218 28508
rect 5608 28428 5613 28484
rect 5669 28428 5696 28484
rect 5752 28428 5779 28484
rect 5835 28428 5861 28484
rect 5917 28428 5943 28484
rect 5999 28428 6025 28484
rect 6081 28428 6107 28484
rect 6163 28428 6189 28484
rect 6245 28428 6271 28484
rect 6327 28428 6353 28484
rect 6409 28428 6435 28484
rect 6491 28428 6517 28484
rect 6573 28428 6599 28484
rect 6655 28428 6681 28484
rect 6737 28428 6763 28484
rect 6819 28428 6845 28484
rect 6901 28428 6927 28484
rect 6983 28428 7009 28484
rect 7065 28428 7091 28484
rect 7147 28428 7173 28484
rect 7229 28428 7255 28484
rect 7311 28428 7337 28484
rect 7393 28428 7419 28484
rect 7475 28428 7501 28484
rect 7557 28428 7583 28484
rect 7639 28428 7665 28484
rect 7721 28428 7747 28484
rect 7803 28428 7829 28484
rect 7885 28428 7911 28484
rect 7967 28428 7993 28484
rect 8049 28428 8075 28484
rect 8131 28428 8157 28484
rect 8213 28428 8218 28484
rect 5608 28404 8218 28428
rect 5608 28348 5613 28404
rect 5669 28348 5696 28404
rect 5752 28348 5779 28404
rect 5835 28348 5861 28404
rect 5917 28348 5943 28404
rect 5999 28348 6025 28404
rect 6081 28348 6107 28404
rect 6163 28348 6189 28404
rect 6245 28348 6271 28404
rect 6327 28348 6353 28404
rect 6409 28348 6435 28404
rect 6491 28348 6517 28404
rect 6573 28348 6599 28404
rect 6655 28348 6681 28404
rect 6737 28348 6763 28404
rect 6819 28348 6845 28404
rect 6901 28348 6927 28404
rect 6983 28348 7009 28404
rect 7065 28348 7091 28404
rect 7147 28348 7173 28404
rect 7229 28348 7255 28404
rect 7311 28348 7337 28404
rect 7393 28348 7419 28404
rect 7475 28348 7501 28404
rect 7557 28348 7583 28404
rect 7639 28348 7665 28404
rect 7721 28348 7747 28404
rect 7803 28348 7829 28404
rect 7885 28348 7911 28404
rect 7967 28348 7993 28404
rect 8049 28348 8075 28404
rect 8131 28348 8157 28404
rect 8213 28348 8218 28404
rect 5608 28324 8218 28348
rect 5608 28268 5613 28324
rect 5669 28268 5696 28324
rect 5752 28268 5779 28324
rect 5835 28268 5861 28324
rect 5917 28268 5943 28324
rect 5999 28268 6025 28324
rect 6081 28268 6107 28324
rect 6163 28268 6189 28324
rect 6245 28268 6271 28324
rect 6327 28268 6353 28324
rect 6409 28268 6435 28324
rect 6491 28268 6517 28324
rect 6573 28268 6599 28324
rect 6655 28268 6681 28324
rect 6737 28268 6763 28324
rect 6819 28268 6845 28324
rect 6901 28268 6927 28324
rect 6983 28268 7009 28324
rect 7065 28268 7091 28324
rect 7147 28268 7173 28324
rect 7229 28268 7255 28324
rect 7311 28268 7337 28324
rect 7393 28268 7419 28324
rect 7475 28268 7501 28324
rect 7557 28268 7583 28324
rect 7639 28268 7665 28324
rect 7721 28268 7747 28324
rect 7803 28268 7829 28324
rect 7885 28268 7911 28324
rect 7967 28268 7993 28324
rect 8049 28268 8075 28324
rect 8131 28268 8157 28324
rect 8213 28268 8218 28324
rect 5608 28244 8218 28268
rect 5608 28188 5613 28244
rect 5669 28188 5696 28244
rect 5752 28188 5779 28244
rect 5835 28188 5861 28244
rect 5917 28188 5943 28244
rect 5999 28188 6025 28244
rect 6081 28188 6107 28244
rect 6163 28188 6189 28244
rect 6245 28188 6271 28244
rect 6327 28188 6353 28244
rect 6409 28188 6435 28244
rect 6491 28188 6517 28244
rect 6573 28188 6599 28244
rect 6655 28188 6681 28244
rect 6737 28188 6763 28244
rect 6819 28188 6845 28244
rect 6901 28188 6927 28244
rect 6983 28188 7009 28244
rect 7065 28188 7091 28244
rect 7147 28188 7173 28244
rect 7229 28188 7255 28244
rect 7311 28188 7337 28244
rect 7393 28188 7419 28244
rect 7475 28188 7501 28244
rect 7557 28188 7583 28244
rect 7639 28188 7665 28244
rect 7721 28188 7747 28244
rect 7803 28188 7829 28244
rect 7885 28188 7911 28244
rect 7967 28188 7993 28244
rect 8049 28188 8075 28244
rect 8131 28188 8157 28244
rect 8213 28188 8218 28244
rect 5608 28164 8218 28188
rect 5608 28108 5613 28164
rect 5669 28108 5696 28164
rect 5752 28108 5779 28164
rect 5835 28108 5861 28164
rect 5917 28108 5943 28164
rect 5999 28108 6025 28164
rect 6081 28108 6107 28164
rect 6163 28108 6189 28164
rect 6245 28108 6271 28164
rect 6327 28108 6353 28164
rect 6409 28108 6435 28164
rect 6491 28108 6517 28164
rect 6573 28108 6599 28164
rect 6655 28108 6681 28164
rect 6737 28108 6763 28164
rect 6819 28108 6845 28164
rect 6901 28108 6927 28164
rect 6983 28108 7009 28164
rect 7065 28108 7091 28164
rect 7147 28108 7173 28164
rect 7229 28108 7255 28164
rect 7311 28108 7337 28164
rect 7393 28108 7419 28164
rect 7475 28108 7501 28164
rect 7557 28108 7583 28164
rect 7639 28108 7665 28164
rect 7721 28108 7747 28164
rect 7803 28108 7829 28164
rect 7885 28108 7911 28164
rect 7967 28108 7993 28164
rect 8049 28108 8075 28164
rect 8131 28108 8157 28164
rect 8213 28108 8218 28164
rect 5608 26724 8218 28108
rect 5608 26668 5613 26724
rect 5669 26668 5696 26724
rect 5752 26668 5779 26724
rect 5835 26668 5861 26724
rect 5917 26668 5943 26724
rect 5999 26668 6025 26724
rect 6081 26668 6107 26724
rect 6163 26668 6189 26724
rect 6245 26668 6271 26724
rect 6327 26668 6353 26724
rect 6409 26668 6435 26724
rect 6491 26668 6517 26724
rect 6573 26668 6599 26724
rect 6655 26668 6681 26724
rect 6737 26668 6763 26724
rect 6819 26668 6845 26724
rect 6901 26668 6927 26724
rect 6983 26668 7009 26724
rect 7065 26668 7091 26724
rect 7147 26668 7173 26724
rect 7229 26668 7255 26724
rect 7311 26668 7337 26724
rect 7393 26668 7419 26724
rect 7475 26668 7501 26724
rect 7557 26668 7583 26724
rect 7639 26668 7665 26724
rect 7721 26668 7747 26724
rect 7803 26668 7829 26724
rect 7885 26668 7911 26724
rect 7967 26668 7993 26724
rect 8049 26668 8075 26724
rect 8131 26668 8157 26724
rect 8213 26668 8218 26724
rect 5608 26644 8218 26668
rect 5608 26588 5613 26644
rect 5669 26588 5696 26644
rect 5752 26588 5779 26644
rect 5835 26588 5861 26644
rect 5917 26588 5943 26644
rect 5999 26588 6025 26644
rect 6081 26588 6107 26644
rect 6163 26588 6189 26644
rect 6245 26588 6271 26644
rect 6327 26588 6353 26644
rect 6409 26588 6435 26644
rect 6491 26588 6517 26644
rect 6573 26588 6599 26644
rect 6655 26588 6681 26644
rect 6737 26588 6763 26644
rect 6819 26588 6845 26644
rect 6901 26588 6927 26644
rect 6983 26588 7009 26644
rect 7065 26588 7091 26644
rect 7147 26588 7173 26644
rect 7229 26588 7255 26644
rect 7311 26588 7337 26644
rect 7393 26588 7419 26644
rect 7475 26588 7501 26644
rect 7557 26588 7583 26644
rect 7639 26588 7665 26644
rect 7721 26588 7747 26644
rect 7803 26588 7829 26644
rect 7885 26588 7911 26644
rect 7967 26588 7993 26644
rect 8049 26588 8075 26644
rect 8131 26588 8157 26644
rect 8213 26588 8218 26644
rect 5608 26564 8218 26588
rect 5608 26508 5613 26564
rect 5669 26508 5696 26564
rect 5752 26508 5779 26564
rect 5835 26508 5861 26564
rect 5917 26508 5943 26564
rect 5999 26508 6025 26564
rect 6081 26508 6107 26564
rect 6163 26508 6189 26564
rect 6245 26508 6271 26564
rect 6327 26508 6353 26564
rect 6409 26508 6435 26564
rect 6491 26508 6517 26564
rect 6573 26508 6599 26564
rect 6655 26508 6681 26564
rect 6737 26508 6763 26564
rect 6819 26508 6845 26564
rect 6901 26508 6927 26564
rect 6983 26508 7009 26564
rect 7065 26508 7091 26564
rect 7147 26508 7173 26564
rect 7229 26508 7255 26564
rect 7311 26508 7337 26564
rect 7393 26508 7419 26564
rect 7475 26508 7501 26564
rect 7557 26508 7583 26564
rect 7639 26508 7665 26564
rect 7721 26508 7747 26564
rect 7803 26508 7829 26564
rect 7885 26508 7911 26564
rect 7967 26508 7993 26564
rect 8049 26508 8075 26564
rect 8131 26508 8157 26564
rect 8213 26508 8218 26564
rect 5608 26484 8218 26508
rect 5608 26428 5613 26484
rect 5669 26428 5696 26484
rect 5752 26428 5779 26484
rect 5835 26428 5861 26484
rect 5917 26428 5943 26484
rect 5999 26428 6025 26484
rect 6081 26428 6107 26484
rect 6163 26428 6189 26484
rect 6245 26428 6271 26484
rect 6327 26428 6353 26484
rect 6409 26428 6435 26484
rect 6491 26428 6517 26484
rect 6573 26428 6599 26484
rect 6655 26428 6681 26484
rect 6737 26428 6763 26484
rect 6819 26428 6845 26484
rect 6901 26428 6927 26484
rect 6983 26428 7009 26484
rect 7065 26428 7091 26484
rect 7147 26428 7173 26484
rect 7229 26428 7255 26484
rect 7311 26428 7337 26484
rect 7393 26428 7419 26484
rect 7475 26428 7501 26484
rect 7557 26428 7583 26484
rect 7639 26428 7665 26484
rect 7721 26428 7747 26484
rect 7803 26428 7829 26484
rect 7885 26428 7911 26484
rect 7967 26428 7993 26484
rect 8049 26428 8075 26484
rect 8131 26428 8157 26484
rect 8213 26428 8218 26484
rect 5608 26404 8218 26428
rect 5608 26348 5613 26404
rect 5669 26348 5696 26404
rect 5752 26348 5779 26404
rect 5835 26348 5861 26404
rect 5917 26348 5943 26404
rect 5999 26348 6025 26404
rect 6081 26348 6107 26404
rect 6163 26348 6189 26404
rect 6245 26348 6271 26404
rect 6327 26348 6353 26404
rect 6409 26348 6435 26404
rect 6491 26348 6517 26404
rect 6573 26348 6599 26404
rect 6655 26348 6681 26404
rect 6737 26348 6763 26404
rect 6819 26348 6845 26404
rect 6901 26348 6927 26404
rect 6983 26348 7009 26404
rect 7065 26348 7091 26404
rect 7147 26348 7173 26404
rect 7229 26348 7255 26404
rect 7311 26348 7337 26404
rect 7393 26348 7419 26404
rect 7475 26348 7501 26404
rect 7557 26348 7583 26404
rect 7639 26348 7665 26404
rect 7721 26348 7747 26404
rect 7803 26348 7829 26404
rect 7885 26348 7911 26404
rect 7967 26348 7993 26404
rect 8049 26348 8075 26404
rect 8131 26348 8157 26404
rect 8213 26348 8218 26404
rect 5608 26324 8218 26348
rect 5608 26268 5613 26324
rect 5669 26268 5696 26324
rect 5752 26268 5779 26324
rect 5835 26268 5861 26324
rect 5917 26268 5943 26324
rect 5999 26268 6025 26324
rect 6081 26268 6107 26324
rect 6163 26268 6189 26324
rect 6245 26268 6271 26324
rect 6327 26268 6353 26324
rect 6409 26268 6435 26324
rect 6491 26268 6517 26324
rect 6573 26268 6599 26324
rect 6655 26268 6681 26324
rect 6737 26268 6763 26324
rect 6819 26268 6845 26324
rect 6901 26268 6927 26324
rect 6983 26268 7009 26324
rect 7065 26268 7091 26324
rect 7147 26268 7173 26324
rect 7229 26268 7255 26324
rect 7311 26268 7337 26324
rect 7393 26268 7419 26324
rect 7475 26268 7501 26324
rect 7557 26268 7583 26324
rect 7639 26268 7665 26324
rect 7721 26268 7747 26324
rect 7803 26268 7829 26324
rect 7885 26268 7911 26324
rect 7967 26268 7993 26324
rect 8049 26268 8075 26324
rect 8131 26268 8157 26324
rect 8213 26268 8218 26324
rect 5608 26244 8218 26268
rect 5608 26188 5613 26244
rect 5669 26188 5696 26244
rect 5752 26188 5779 26244
rect 5835 26188 5861 26244
rect 5917 26188 5943 26244
rect 5999 26188 6025 26244
rect 6081 26188 6107 26244
rect 6163 26188 6189 26244
rect 6245 26188 6271 26244
rect 6327 26188 6353 26244
rect 6409 26188 6435 26244
rect 6491 26188 6517 26244
rect 6573 26188 6599 26244
rect 6655 26188 6681 26244
rect 6737 26188 6763 26244
rect 6819 26188 6845 26244
rect 6901 26188 6927 26244
rect 6983 26188 7009 26244
rect 7065 26188 7091 26244
rect 7147 26188 7173 26244
rect 7229 26188 7255 26244
rect 7311 26188 7337 26244
rect 7393 26188 7419 26244
rect 7475 26188 7501 26244
rect 7557 26188 7583 26244
rect 7639 26188 7665 26244
rect 7721 26188 7747 26244
rect 7803 26188 7829 26244
rect 7885 26188 7911 26244
rect 7967 26188 7993 26244
rect 8049 26188 8075 26244
rect 8131 26188 8157 26244
rect 8213 26188 8218 26244
rect 5608 26164 8218 26188
rect 5608 26108 5613 26164
rect 5669 26108 5696 26164
rect 5752 26108 5779 26164
rect 5835 26108 5861 26164
rect 5917 26108 5943 26164
rect 5999 26108 6025 26164
rect 6081 26108 6107 26164
rect 6163 26108 6189 26164
rect 6245 26108 6271 26164
rect 6327 26108 6353 26164
rect 6409 26108 6435 26164
rect 6491 26108 6517 26164
rect 6573 26108 6599 26164
rect 6655 26108 6681 26164
rect 6737 26108 6763 26164
rect 6819 26108 6845 26164
rect 6901 26108 6927 26164
rect 6983 26108 7009 26164
rect 7065 26108 7091 26164
rect 7147 26108 7173 26164
rect 7229 26108 7255 26164
rect 7311 26108 7337 26164
rect 7393 26108 7419 26164
rect 7475 26108 7501 26164
rect 7557 26108 7583 26164
rect 7639 26108 7665 26164
rect 7721 26108 7747 26164
rect 7803 26108 7829 26164
rect 7885 26108 7911 26164
rect 7967 26108 7993 26164
rect 8049 26108 8075 26164
rect 8131 26108 8157 26164
rect 8213 26108 8218 26164
rect 5608 24724 8218 26108
rect 5608 24668 5613 24724
rect 5669 24668 5696 24724
rect 5752 24668 5779 24724
rect 5835 24668 5861 24724
rect 5917 24668 5943 24724
rect 5999 24668 6025 24724
rect 6081 24668 6107 24724
rect 6163 24668 6189 24724
rect 6245 24668 6271 24724
rect 6327 24668 6353 24724
rect 6409 24668 6435 24724
rect 6491 24668 6517 24724
rect 6573 24668 6599 24724
rect 6655 24668 6681 24724
rect 6737 24668 6763 24724
rect 6819 24668 6845 24724
rect 6901 24668 6927 24724
rect 6983 24668 7009 24724
rect 7065 24668 7091 24724
rect 7147 24668 7173 24724
rect 7229 24668 7255 24724
rect 7311 24668 7337 24724
rect 7393 24668 7419 24724
rect 7475 24668 7501 24724
rect 7557 24668 7583 24724
rect 7639 24668 7665 24724
rect 7721 24668 7747 24724
rect 7803 24668 7829 24724
rect 7885 24668 7911 24724
rect 7967 24668 7993 24724
rect 8049 24668 8075 24724
rect 8131 24668 8157 24724
rect 8213 24668 8218 24724
rect 5608 24644 8218 24668
rect 5608 24588 5613 24644
rect 5669 24588 5696 24644
rect 5752 24588 5779 24644
rect 5835 24588 5861 24644
rect 5917 24588 5943 24644
rect 5999 24588 6025 24644
rect 6081 24588 6107 24644
rect 6163 24588 6189 24644
rect 6245 24588 6271 24644
rect 6327 24588 6353 24644
rect 6409 24588 6435 24644
rect 6491 24588 6517 24644
rect 6573 24588 6599 24644
rect 6655 24588 6681 24644
rect 6737 24588 6763 24644
rect 6819 24588 6845 24644
rect 6901 24588 6927 24644
rect 6983 24588 7009 24644
rect 7065 24588 7091 24644
rect 7147 24588 7173 24644
rect 7229 24588 7255 24644
rect 7311 24588 7337 24644
rect 7393 24588 7419 24644
rect 7475 24588 7501 24644
rect 7557 24588 7583 24644
rect 7639 24588 7665 24644
rect 7721 24588 7747 24644
rect 7803 24588 7829 24644
rect 7885 24588 7911 24644
rect 7967 24588 7993 24644
rect 8049 24588 8075 24644
rect 8131 24588 8157 24644
rect 8213 24588 8218 24644
rect 5608 24564 8218 24588
rect 5608 24508 5613 24564
rect 5669 24508 5696 24564
rect 5752 24508 5779 24564
rect 5835 24508 5861 24564
rect 5917 24508 5943 24564
rect 5999 24508 6025 24564
rect 6081 24508 6107 24564
rect 6163 24508 6189 24564
rect 6245 24508 6271 24564
rect 6327 24508 6353 24564
rect 6409 24508 6435 24564
rect 6491 24508 6517 24564
rect 6573 24508 6599 24564
rect 6655 24508 6681 24564
rect 6737 24508 6763 24564
rect 6819 24508 6845 24564
rect 6901 24508 6927 24564
rect 6983 24508 7009 24564
rect 7065 24508 7091 24564
rect 7147 24508 7173 24564
rect 7229 24508 7255 24564
rect 7311 24508 7337 24564
rect 7393 24508 7419 24564
rect 7475 24508 7501 24564
rect 7557 24508 7583 24564
rect 7639 24508 7665 24564
rect 7721 24508 7747 24564
rect 7803 24508 7829 24564
rect 7885 24508 7911 24564
rect 7967 24508 7993 24564
rect 8049 24508 8075 24564
rect 8131 24508 8157 24564
rect 8213 24508 8218 24564
rect 5608 24484 8218 24508
rect 5608 24428 5613 24484
rect 5669 24428 5696 24484
rect 5752 24428 5779 24484
rect 5835 24428 5861 24484
rect 5917 24428 5943 24484
rect 5999 24428 6025 24484
rect 6081 24428 6107 24484
rect 6163 24428 6189 24484
rect 6245 24428 6271 24484
rect 6327 24428 6353 24484
rect 6409 24428 6435 24484
rect 6491 24428 6517 24484
rect 6573 24428 6599 24484
rect 6655 24428 6681 24484
rect 6737 24428 6763 24484
rect 6819 24428 6845 24484
rect 6901 24428 6927 24484
rect 6983 24428 7009 24484
rect 7065 24428 7091 24484
rect 7147 24428 7173 24484
rect 7229 24428 7255 24484
rect 7311 24428 7337 24484
rect 7393 24428 7419 24484
rect 7475 24428 7501 24484
rect 7557 24428 7583 24484
rect 7639 24428 7665 24484
rect 7721 24428 7747 24484
rect 7803 24428 7829 24484
rect 7885 24428 7911 24484
rect 7967 24428 7993 24484
rect 8049 24428 8075 24484
rect 8131 24428 8157 24484
rect 8213 24428 8218 24484
rect 5608 24404 8218 24428
rect 5608 24348 5613 24404
rect 5669 24348 5696 24404
rect 5752 24348 5779 24404
rect 5835 24348 5861 24404
rect 5917 24348 5943 24404
rect 5999 24348 6025 24404
rect 6081 24348 6107 24404
rect 6163 24348 6189 24404
rect 6245 24348 6271 24404
rect 6327 24348 6353 24404
rect 6409 24348 6435 24404
rect 6491 24348 6517 24404
rect 6573 24348 6599 24404
rect 6655 24348 6681 24404
rect 6737 24348 6763 24404
rect 6819 24348 6845 24404
rect 6901 24348 6927 24404
rect 6983 24348 7009 24404
rect 7065 24348 7091 24404
rect 7147 24348 7173 24404
rect 7229 24348 7255 24404
rect 7311 24348 7337 24404
rect 7393 24348 7419 24404
rect 7475 24348 7501 24404
rect 7557 24348 7583 24404
rect 7639 24348 7665 24404
rect 7721 24348 7747 24404
rect 7803 24348 7829 24404
rect 7885 24348 7911 24404
rect 7967 24348 7993 24404
rect 8049 24348 8075 24404
rect 8131 24348 8157 24404
rect 8213 24348 8218 24404
rect 5608 24324 8218 24348
rect 5608 24268 5613 24324
rect 5669 24268 5696 24324
rect 5752 24268 5779 24324
rect 5835 24268 5861 24324
rect 5917 24268 5943 24324
rect 5999 24268 6025 24324
rect 6081 24268 6107 24324
rect 6163 24268 6189 24324
rect 6245 24268 6271 24324
rect 6327 24268 6353 24324
rect 6409 24268 6435 24324
rect 6491 24268 6517 24324
rect 6573 24268 6599 24324
rect 6655 24268 6681 24324
rect 6737 24268 6763 24324
rect 6819 24268 6845 24324
rect 6901 24268 6927 24324
rect 6983 24268 7009 24324
rect 7065 24268 7091 24324
rect 7147 24268 7173 24324
rect 7229 24268 7255 24324
rect 7311 24268 7337 24324
rect 7393 24268 7419 24324
rect 7475 24268 7501 24324
rect 7557 24268 7583 24324
rect 7639 24268 7665 24324
rect 7721 24268 7747 24324
rect 7803 24268 7829 24324
rect 7885 24268 7911 24324
rect 7967 24268 7993 24324
rect 8049 24268 8075 24324
rect 8131 24268 8157 24324
rect 8213 24268 8218 24324
rect 5608 24244 8218 24268
rect 5608 24188 5613 24244
rect 5669 24188 5696 24244
rect 5752 24188 5779 24244
rect 5835 24188 5861 24244
rect 5917 24188 5943 24244
rect 5999 24188 6025 24244
rect 6081 24188 6107 24244
rect 6163 24188 6189 24244
rect 6245 24188 6271 24244
rect 6327 24188 6353 24244
rect 6409 24188 6435 24244
rect 6491 24188 6517 24244
rect 6573 24188 6599 24244
rect 6655 24188 6681 24244
rect 6737 24188 6763 24244
rect 6819 24188 6845 24244
rect 6901 24188 6927 24244
rect 6983 24188 7009 24244
rect 7065 24188 7091 24244
rect 7147 24188 7173 24244
rect 7229 24188 7255 24244
rect 7311 24188 7337 24244
rect 7393 24188 7419 24244
rect 7475 24188 7501 24244
rect 7557 24188 7583 24244
rect 7639 24188 7665 24244
rect 7721 24188 7747 24244
rect 7803 24188 7829 24244
rect 7885 24188 7911 24244
rect 7967 24188 7993 24244
rect 8049 24188 8075 24244
rect 8131 24188 8157 24244
rect 8213 24188 8218 24244
rect 5608 24164 8218 24188
rect 5608 24108 5613 24164
rect 5669 24108 5696 24164
rect 5752 24108 5779 24164
rect 5835 24108 5861 24164
rect 5917 24108 5943 24164
rect 5999 24108 6025 24164
rect 6081 24108 6107 24164
rect 6163 24108 6189 24164
rect 6245 24108 6271 24164
rect 6327 24108 6353 24164
rect 6409 24108 6435 24164
rect 6491 24108 6517 24164
rect 6573 24108 6599 24164
rect 6655 24108 6681 24164
rect 6737 24108 6763 24164
rect 6819 24108 6845 24164
rect 6901 24108 6927 24164
rect 6983 24108 7009 24164
rect 7065 24108 7091 24164
rect 7147 24108 7173 24164
rect 7229 24108 7255 24164
rect 7311 24108 7337 24164
rect 7393 24108 7419 24164
rect 7475 24108 7501 24164
rect 7557 24108 7583 24164
rect 7639 24108 7665 24164
rect 7721 24108 7747 24164
rect 7803 24108 7829 24164
rect 7885 24108 7911 24164
rect 7967 24108 7993 24164
rect 8049 24108 8075 24164
rect 8131 24108 8157 24164
rect 8213 24108 8218 24164
rect 5608 22724 8218 24108
rect 5608 22668 5613 22724
rect 5669 22668 5696 22724
rect 5752 22668 5779 22724
rect 5835 22668 5861 22724
rect 5917 22668 5943 22724
rect 5999 22668 6025 22724
rect 6081 22668 6107 22724
rect 6163 22668 6189 22724
rect 6245 22668 6271 22724
rect 6327 22668 6353 22724
rect 6409 22668 6435 22724
rect 6491 22668 6517 22724
rect 6573 22668 6599 22724
rect 6655 22668 6681 22724
rect 6737 22668 6763 22724
rect 6819 22668 6845 22724
rect 6901 22668 6927 22724
rect 6983 22668 7009 22724
rect 7065 22668 7091 22724
rect 7147 22668 7173 22724
rect 7229 22668 7255 22724
rect 7311 22668 7337 22724
rect 7393 22668 7419 22724
rect 7475 22668 7501 22724
rect 7557 22668 7583 22724
rect 7639 22668 7665 22724
rect 7721 22668 7747 22724
rect 7803 22668 7829 22724
rect 7885 22668 7911 22724
rect 7967 22668 7993 22724
rect 8049 22668 8075 22724
rect 8131 22668 8157 22724
rect 8213 22668 8218 22724
rect 5608 22644 8218 22668
rect 5608 22588 5613 22644
rect 5669 22588 5696 22644
rect 5752 22588 5779 22644
rect 5835 22588 5861 22644
rect 5917 22588 5943 22644
rect 5999 22588 6025 22644
rect 6081 22588 6107 22644
rect 6163 22588 6189 22644
rect 6245 22588 6271 22644
rect 6327 22588 6353 22644
rect 6409 22588 6435 22644
rect 6491 22588 6517 22644
rect 6573 22588 6599 22644
rect 6655 22588 6681 22644
rect 6737 22588 6763 22644
rect 6819 22588 6845 22644
rect 6901 22588 6927 22644
rect 6983 22588 7009 22644
rect 7065 22588 7091 22644
rect 7147 22588 7173 22644
rect 7229 22588 7255 22644
rect 7311 22588 7337 22644
rect 7393 22588 7419 22644
rect 7475 22588 7501 22644
rect 7557 22588 7583 22644
rect 7639 22588 7665 22644
rect 7721 22588 7747 22644
rect 7803 22588 7829 22644
rect 7885 22588 7911 22644
rect 7967 22588 7993 22644
rect 8049 22588 8075 22644
rect 8131 22588 8157 22644
rect 8213 22588 8218 22644
rect 5608 22564 8218 22588
rect 5608 22508 5613 22564
rect 5669 22508 5696 22564
rect 5752 22508 5779 22564
rect 5835 22508 5861 22564
rect 5917 22508 5943 22564
rect 5999 22508 6025 22564
rect 6081 22508 6107 22564
rect 6163 22508 6189 22564
rect 6245 22508 6271 22564
rect 6327 22508 6353 22564
rect 6409 22508 6435 22564
rect 6491 22508 6517 22564
rect 6573 22508 6599 22564
rect 6655 22508 6681 22564
rect 6737 22508 6763 22564
rect 6819 22508 6845 22564
rect 6901 22508 6927 22564
rect 6983 22508 7009 22564
rect 7065 22508 7091 22564
rect 7147 22508 7173 22564
rect 7229 22508 7255 22564
rect 7311 22508 7337 22564
rect 7393 22508 7419 22564
rect 7475 22508 7501 22564
rect 7557 22508 7583 22564
rect 7639 22508 7665 22564
rect 7721 22508 7747 22564
rect 7803 22508 7829 22564
rect 7885 22508 7911 22564
rect 7967 22508 7993 22564
rect 8049 22508 8075 22564
rect 8131 22508 8157 22564
rect 8213 22508 8218 22564
rect 5608 22484 8218 22508
rect 5608 22428 5613 22484
rect 5669 22428 5696 22484
rect 5752 22428 5779 22484
rect 5835 22428 5861 22484
rect 5917 22428 5943 22484
rect 5999 22428 6025 22484
rect 6081 22428 6107 22484
rect 6163 22428 6189 22484
rect 6245 22428 6271 22484
rect 6327 22428 6353 22484
rect 6409 22428 6435 22484
rect 6491 22428 6517 22484
rect 6573 22428 6599 22484
rect 6655 22428 6681 22484
rect 6737 22428 6763 22484
rect 6819 22428 6845 22484
rect 6901 22428 6927 22484
rect 6983 22428 7009 22484
rect 7065 22428 7091 22484
rect 7147 22428 7173 22484
rect 7229 22428 7255 22484
rect 7311 22428 7337 22484
rect 7393 22428 7419 22484
rect 7475 22428 7501 22484
rect 7557 22428 7583 22484
rect 7639 22428 7665 22484
rect 7721 22428 7747 22484
rect 7803 22428 7829 22484
rect 7885 22428 7911 22484
rect 7967 22428 7993 22484
rect 8049 22428 8075 22484
rect 8131 22428 8157 22484
rect 8213 22428 8218 22484
rect 5608 22404 8218 22428
rect 5608 22348 5613 22404
rect 5669 22348 5696 22404
rect 5752 22348 5779 22404
rect 5835 22348 5861 22404
rect 5917 22348 5943 22404
rect 5999 22348 6025 22404
rect 6081 22348 6107 22404
rect 6163 22348 6189 22404
rect 6245 22348 6271 22404
rect 6327 22348 6353 22404
rect 6409 22348 6435 22404
rect 6491 22348 6517 22404
rect 6573 22348 6599 22404
rect 6655 22348 6681 22404
rect 6737 22348 6763 22404
rect 6819 22348 6845 22404
rect 6901 22348 6927 22404
rect 6983 22348 7009 22404
rect 7065 22348 7091 22404
rect 7147 22348 7173 22404
rect 7229 22348 7255 22404
rect 7311 22348 7337 22404
rect 7393 22348 7419 22404
rect 7475 22348 7501 22404
rect 7557 22348 7583 22404
rect 7639 22348 7665 22404
rect 7721 22348 7747 22404
rect 7803 22348 7829 22404
rect 7885 22348 7911 22404
rect 7967 22348 7993 22404
rect 8049 22348 8075 22404
rect 8131 22348 8157 22404
rect 8213 22348 8218 22404
rect 5608 22324 8218 22348
rect 5608 22268 5613 22324
rect 5669 22268 5696 22324
rect 5752 22268 5779 22324
rect 5835 22268 5861 22324
rect 5917 22268 5943 22324
rect 5999 22268 6025 22324
rect 6081 22268 6107 22324
rect 6163 22268 6189 22324
rect 6245 22268 6271 22324
rect 6327 22268 6353 22324
rect 6409 22268 6435 22324
rect 6491 22268 6517 22324
rect 6573 22268 6599 22324
rect 6655 22268 6681 22324
rect 6737 22268 6763 22324
rect 6819 22268 6845 22324
rect 6901 22268 6927 22324
rect 6983 22268 7009 22324
rect 7065 22268 7091 22324
rect 7147 22268 7173 22324
rect 7229 22268 7255 22324
rect 7311 22268 7337 22324
rect 7393 22268 7419 22324
rect 7475 22268 7501 22324
rect 7557 22268 7583 22324
rect 7639 22268 7665 22324
rect 7721 22268 7747 22324
rect 7803 22268 7829 22324
rect 7885 22268 7911 22324
rect 7967 22268 7993 22324
rect 8049 22268 8075 22324
rect 8131 22268 8157 22324
rect 8213 22268 8218 22324
rect 5608 22244 8218 22268
rect 5608 22188 5613 22244
rect 5669 22188 5696 22244
rect 5752 22188 5779 22244
rect 5835 22188 5861 22244
rect 5917 22188 5943 22244
rect 5999 22188 6025 22244
rect 6081 22188 6107 22244
rect 6163 22188 6189 22244
rect 6245 22188 6271 22244
rect 6327 22188 6353 22244
rect 6409 22188 6435 22244
rect 6491 22188 6517 22244
rect 6573 22188 6599 22244
rect 6655 22188 6681 22244
rect 6737 22188 6763 22244
rect 6819 22188 6845 22244
rect 6901 22188 6927 22244
rect 6983 22188 7009 22244
rect 7065 22188 7091 22244
rect 7147 22188 7173 22244
rect 7229 22188 7255 22244
rect 7311 22188 7337 22244
rect 7393 22188 7419 22244
rect 7475 22188 7501 22244
rect 7557 22188 7583 22244
rect 7639 22188 7665 22244
rect 7721 22188 7747 22244
rect 7803 22188 7829 22244
rect 7885 22188 7911 22244
rect 7967 22188 7993 22244
rect 8049 22188 8075 22244
rect 8131 22188 8157 22244
rect 8213 22188 8218 22244
rect 5608 22164 8218 22188
rect 5608 22108 5613 22164
rect 5669 22108 5696 22164
rect 5752 22108 5779 22164
rect 5835 22108 5861 22164
rect 5917 22108 5943 22164
rect 5999 22108 6025 22164
rect 6081 22108 6107 22164
rect 6163 22108 6189 22164
rect 6245 22108 6271 22164
rect 6327 22108 6353 22164
rect 6409 22108 6435 22164
rect 6491 22108 6517 22164
rect 6573 22108 6599 22164
rect 6655 22108 6681 22164
rect 6737 22108 6763 22164
rect 6819 22108 6845 22164
rect 6901 22108 6927 22164
rect 6983 22108 7009 22164
rect 7065 22108 7091 22164
rect 7147 22108 7173 22164
rect 7229 22108 7255 22164
rect 7311 22108 7337 22164
rect 7393 22108 7419 22164
rect 7475 22108 7501 22164
rect 7557 22108 7583 22164
rect 7639 22108 7665 22164
rect 7721 22108 7747 22164
rect 7803 22108 7829 22164
rect 7885 22108 7911 22164
rect 7967 22108 7993 22164
rect 8049 22108 8075 22164
rect 8131 22108 8157 22164
rect 8213 22108 8218 22164
rect 5608 20724 8218 22108
rect 5608 20668 5613 20724
rect 5669 20668 5696 20724
rect 5752 20668 5779 20724
rect 5835 20668 5861 20724
rect 5917 20668 5943 20724
rect 5999 20668 6025 20724
rect 6081 20668 6107 20724
rect 6163 20668 6189 20724
rect 6245 20668 6271 20724
rect 6327 20668 6353 20724
rect 6409 20668 6435 20724
rect 6491 20668 6517 20724
rect 6573 20668 6599 20724
rect 6655 20668 6681 20724
rect 6737 20668 6763 20724
rect 6819 20668 6845 20724
rect 6901 20668 6927 20724
rect 6983 20668 7009 20724
rect 7065 20668 7091 20724
rect 7147 20668 7173 20724
rect 7229 20668 7255 20724
rect 7311 20668 7337 20724
rect 7393 20668 7419 20724
rect 7475 20668 7501 20724
rect 7557 20668 7583 20724
rect 7639 20668 7665 20724
rect 7721 20668 7747 20724
rect 7803 20668 7829 20724
rect 7885 20668 7911 20724
rect 7967 20668 7993 20724
rect 8049 20668 8075 20724
rect 8131 20668 8157 20724
rect 8213 20668 8218 20724
rect 5608 20644 8218 20668
rect 5608 20588 5613 20644
rect 5669 20588 5696 20644
rect 5752 20588 5779 20644
rect 5835 20588 5861 20644
rect 5917 20588 5943 20644
rect 5999 20588 6025 20644
rect 6081 20588 6107 20644
rect 6163 20588 6189 20644
rect 6245 20588 6271 20644
rect 6327 20588 6353 20644
rect 6409 20588 6435 20644
rect 6491 20588 6517 20644
rect 6573 20588 6599 20644
rect 6655 20588 6681 20644
rect 6737 20588 6763 20644
rect 6819 20588 6845 20644
rect 6901 20588 6927 20644
rect 6983 20588 7009 20644
rect 7065 20588 7091 20644
rect 7147 20588 7173 20644
rect 7229 20588 7255 20644
rect 7311 20588 7337 20644
rect 7393 20588 7419 20644
rect 7475 20588 7501 20644
rect 7557 20588 7583 20644
rect 7639 20588 7665 20644
rect 7721 20588 7747 20644
rect 7803 20588 7829 20644
rect 7885 20588 7911 20644
rect 7967 20588 7993 20644
rect 8049 20588 8075 20644
rect 8131 20588 8157 20644
rect 8213 20588 8218 20644
rect 5608 20564 8218 20588
rect 5608 20508 5613 20564
rect 5669 20508 5696 20564
rect 5752 20508 5779 20564
rect 5835 20508 5861 20564
rect 5917 20508 5943 20564
rect 5999 20508 6025 20564
rect 6081 20508 6107 20564
rect 6163 20508 6189 20564
rect 6245 20508 6271 20564
rect 6327 20508 6353 20564
rect 6409 20508 6435 20564
rect 6491 20508 6517 20564
rect 6573 20508 6599 20564
rect 6655 20508 6681 20564
rect 6737 20508 6763 20564
rect 6819 20508 6845 20564
rect 6901 20508 6927 20564
rect 6983 20508 7009 20564
rect 7065 20508 7091 20564
rect 7147 20508 7173 20564
rect 7229 20508 7255 20564
rect 7311 20508 7337 20564
rect 7393 20508 7419 20564
rect 7475 20508 7501 20564
rect 7557 20508 7583 20564
rect 7639 20508 7665 20564
rect 7721 20508 7747 20564
rect 7803 20508 7829 20564
rect 7885 20508 7911 20564
rect 7967 20508 7993 20564
rect 8049 20508 8075 20564
rect 8131 20508 8157 20564
rect 8213 20508 8218 20564
rect 5608 20484 8218 20508
rect 5608 20428 5613 20484
rect 5669 20428 5696 20484
rect 5752 20428 5779 20484
rect 5835 20428 5861 20484
rect 5917 20428 5943 20484
rect 5999 20428 6025 20484
rect 6081 20428 6107 20484
rect 6163 20428 6189 20484
rect 6245 20428 6271 20484
rect 6327 20428 6353 20484
rect 6409 20428 6435 20484
rect 6491 20428 6517 20484
rect 6573 20428 6599 20484
rect 6655 20428 6681 20484
rect 6737 20428 6763 20484
rect 6819 20428 6845 20484
rect 6901 20428 6927 20484
rect 6983 20428 7009 20484
rect 7065 20428 7091 20484
rect 7147 20428 7173 20484
rect 7229 20428 7255 20484
rect 7311 20428 7337 20484
rect 7393 20428 7419 20484
rect 7475 20428 7501 20484
rect 7557 20428 7583 20484
rect 7639 20428 7665 20484
rect 7721 20428 7747 20484
rect 7803 20428 7829 20484
rect 7885 20428 7911 20484
rect 7967 20428 7993 20484
rect 8049 20428 8075 20484
rect 8131 20428 8157 20484
rect 8213 20428 8218 20484
rect 5608 20404 8218 20428
rect 5608 20348 5613 20404
rect 5669 20348 5696 20404
rect 5752 20348 5779 20404
rect 5835 20348 5861 20404
rect 5917 20348 5943 20404
rect 5999 20348 6025 20404
rect 6081 20348 6107 20404
rect 6163 20348 6189 20404
rect 6245 20348 6271 20404
rect 6327 20348 6353 20404
rect 6409 20348 6435 20404
rect 6491 20348 6517 20404
rect 6573 20348 6599 20404
rect 6655 20348 6681 20404
rect 6737 20348 6763 20404
rect 6819 20348 6845 20404
rect 6901 20348 6927 20404
rect 6983 20348 7009 20404
rect 7065 20348 7091 20404
rect 7147 20348 7173 20404
rect 7229 20348 7255 20404
rect 7311 20348 7337 20404
rect 7393 20348 7419 20404
rect 7475 20348 7501 20404
rect 7557 20348 7583 20404
rect 7639 20348 7665 20404
rect 7721 20348 7747 20404
rect 7803 20348 7829 20404
rect 7885 20348 7911 20404
rect 7967 20348 7993 20404
rect 8049 20348 8075 20404
rect 8131 20348 8157 20404
rect 8213 20348 8218 20404
rect 5608 20324 8218 20348
rect 5608 20268 5613 20324
rect 5669 20268 5696 20324
rect 5752 20268 5779 20324
rect 5835 20268 5861 20324
rect 5917 20268 5943 20324
rect 5999 20268 6025 20324
rect 6081 20268 6107 20324
rect 6163 20268 6189 20324
rect 6245 20268 6271 20324
rect 6327 20268 6353 20324
rect 6409 20268 6435 20324
rect 6491 20268 6517 20324
rect 6573 20268 6599 20324
rect 6655 20268 6681 20324
rect 6737 20268 6763 20324
rect 6819 20268 6845 20324
rect 6901 20268 6927 20324
rect 6983 20268 7009 20324
rect 7065 20268 7091 20324
rect 7147 20268 7173 20324
rect 7229 20268 7255 20324
rect 7311 20268 7337 20324
rect 7393 20268 7419 20324
rect 7475 20268 7501 20324
rect 7557 20268 7583 20324
rect 7639 20268 7665 20324
rect 7721 20268 7747 20324
rect 7803 20268 7829 20324
rect 7885 20268 7911 20324
rect 7967 20268 7993 20324
rect 8049 20268 8075 20324
rect 8131 20268 8157 20324
rect 8213 20268 8218 20324
rect 5608 20244 8218 20268
rect 5608 20188 5613 20244
rect 5669 20188 5696 20244
rect 5752 20188 5779 20244
rect 5835 20188 5861 20244
rect 5917 20188 5943 20244
rect 5999 20188 6025 20244
rect 6081 20188 6107 20244
rect 6163 20188 6189 20244
rect 6245 20188 6271 20244
rect 6327 20188 6353 20244
rect 6409 20188 6435 20244
rect 6491 20188 6517 20244
rect 6573 20188 6599 20244
rect 6655 20188 6681 20244
rect 6737 20188 6763 20244
rect 6819 20188 6845 20244
rect 6901 20188 6927 20244
rect 6983 20188 7009 20244
rect 7065 20188 7091 20244
rect 7147 20188 7173 20244
rect 7229 20188 7255 20244
rect 7311 20188 7337 20244
rect 7393 20188 7419 20244
rect 7475 20188 7501 20244
rect 7557 20188 7583 20244
rect 7639 20188 7665 20244
rect 7721 20188 7747 20244
rect 7803 20188 7829 20244
rect 7885 20188 7911 20244
rect 7967 20188 7993 20244
rect 8049 20188 8075 20244
rect 8131 20188 8157 20244
rect 8213 20188 8218 20244
rect 5608 20164 8218 20188
rect 5608 20108 5613 20164
rect 5669 20108 5696 20164
rect 5752 20108 5779 20164
rect 5835 20108 5861 20164
rect 5917 20108 5943 20164
rect 5999 20108 6025 20164
rect 6081 20108 6107 20164
rect 6163 20108 6189 20164
rect 6245 20108 6271 20164
rect 6327 20108 6353 20164
rect 6409 20108 6435 20164
rect 6491 20108 6517 20164
rect 6573 20108 6599 20164
rect 6655 20108 6681 20164
rect 6737 20108 6763 20164
rect 6819 20108 6845 20164
rect 6901 20108 6927 20164
rect 6983 20108 7009 20164
rect 7065 20108 7091 20164
rect 7147 20108 7173 20164
rect 7229 20108 7255 20164
rect 7311 20108 7337 20164
rect 7393 20108 7419 20164
rect 7475 20108 7501 20164
rect 7557 20108 7583 20164
rect 7639 20108 7665 20164
rect 7721 20108 7747 20164
rect 7803 20108 7829 20164
rect 7885 20108 7911 20164
rect 7967 20108 7993 20164
rect 8049 20108 8075 20164
rect 8131 20108 8157 20164
rect 8213 20108 8218 20164
rect 5608 18724 8218 20108
rect 5608 18668 5613 18724
rect 5669 18668 5696 18724
rect 5752 18668 5779 18724
rect 5835 18668 5861 18724
rect 5917 18668 5943 18724
rect 5999 18668 6025 18724
rect 6081 18668 6107 18724
rect 6163 18668 6189 18724
rect 6245 18668 6271 18724
rect 6327 18668 6353 18724
rect 6409 18668 6435 18724
rect 6491 18668 6517 18724
rect 6573 18668 6599 18724
rect 6655 18668 6681 18724
rect 6737 18668 6763 18724
rect 6819 18668 6845 18724
rect 6901 18668 6927 18724
rect 6983 18668 7009 18724
rect 7065 18668 7091 18724
rect 7147 18668 7173 18724
rect 7229 18668 7255 18724
rect 7311 18668 7337 18724
rect 7393 18668 7419 18724
rect 7475 18668 7501 18724
rect 7557 18668 7583 18724
rect 7639 18668 7665 18724
rect 7721 18668 7747 18724
rect 7803 18668 7829 18724
rect 7885 18668 7911 18724
rect 7967 18668 7993 18724
rect 8049 18668 8075 18724
rect 8131 18668 8157 18724
rect 8213 18668 8218 18724
rect 5608 18644 8218 18668
rect 5608 18588 5613 18644
rect 5669 18588 5696 18644
rect 5752 18588 5779 18644
rect 5835 18588 5861 18644
rect 5917 18588 5943 18644
rect 5999 18588 6025 18644
rect 6081 18588 6107 18644
rect 6163 18588 6189 18644
rect 6245 18588 6271 18644
rect 6327 18588 6353 18644
rect 6409 18588 6435 18644
rect 6491 18588 6517 18644
rect 6573 18588 6599 18644
rect 6655 18588 6681 18644
rect 6737 18588 6763 18644
rect 6819 18588 6845 18644
rect 6901 18588 6927 18644
rect 6983 18588 7009 18644
rect 7065 18588 7091 18644
rect 7147 18588 7173 18644
rect 7229 18588 7255 18644
rect 7311 18588 7337 18644
rect 7393 18588 7419 18644
rect 7475 18588 7501 18644
rect 7557 18588 7583 18644
rect 7639 18588 7665 18644
rect 7721 18588 7747 18644
rect 7803 18588 7829 18644
rect 7885 18588 7911 18644
rect 7967 18588 7993 18644
rect 8049 18588 8075 18644
rect 8131 18588 8157 18644
rect 8213 18588 8218 18644
rect 5608 18564 8218 18588
rect 5608 18508 5613 18564
rect 5669 18508 5696 18564
rect 5752 18508 5779 18564
rect 5835 18508 5861 18564
rect 5917 18508 5943 18564
rect 5999 18508 6025 18564
rect 6081 18508 6107 18564
rect 6163 18508 6189 18564
rect 6245 18508 6271 18564
rect 6327 18508 6353 18564
rect 6409 18508 6435 18564
rect 6491 18508 6517 18564
rect 6573 18508 6599 18564
rect 6655 18508 6681 18564
rect 6737 18508 6763 18564
rect 6819 18508 6845 18564
rect 6901 18508 6927 18564
rect 6983 18508 7009 18564
rect 7065 18508 7091 18564
rect 7147 18508 7173 18564
rect 7229 18508 7255 18564
rect 7311 18508 7337 18564
rect 7393 18508 7419 18564
rect 7475 18508 7501 18564
rect 7557 18508 7583 18564
rect 7639 18508 7665 18564
rect 7721 18508 7747 18564
rect 7803 18508 7829 18564
rect 7885 18508 7911 18564
rect 7967 18508 7993 18564
rect 8049 18508 8075 18564
rect 8131 18508 8157 18564
rect 8213 18508 8218 18564
rect 5608 18484 8218 18508
rect 5608 18428 5613 18484
rect 5669 18428 5696 18484
rect 5752 18428 5779 18484
rect 5835 18428 5861 18484
rect 5917 18428 5943 18484
rect 5999 18428 6025 18484
rect 6081 18428 6107 18484
rect 6163 18428 6189 18484
rect 6245 18428 6271 18484
rect 6327 18428 6353 18484
rect 6409 18428 6435 18484
rect 6491 18428 6517 18484
rect 6573 18428 6599 18484
rect 6655 18428 6681 18484
rect 6737 18428 6763 18484
rect 6819 18428 6845 18484
rect 6901 18428 6927 18484
rect 6983 18428 7009 18484
rect 7065 18428 7091 18484
rect 7147 18428 7173 18484
rect 7229 18428 7255 18484
rect 7311 18428 7337 18484
rect 7393 18428 7419 18484
rect 7475 18428 7501 18484
rect 7557 18428 7583 18484
rect 7639 18428 7665 18484
rect 7721 18428 7747 18484
rect 7803 18428 7829 18484
rect 7885 18428 7911 18484
rect 7967 18428 7993 18484
rect 8049 18428 8075 18484
rect 8131 18428 8157 18484
rect 8213 18428 8218 18484
rect 5608 18404 8218 18428
rect 5608 18348 5613 18404
rect 5669 18348 5696 18404
rect 5752 18348 5779 18404
rect 5835 18348 5861 18404
rect 5917 18348 5943 18404
rect 5999 18348 6025 18404
rect 6081 18348 6107 18404
rect 6163 18348 6189 18404
rect 6245 18348 6271 18404
rect 6327 18348 6353 18404
rect 6409 18348 6435 18404
rect 6491 18348 6517 18404
rect 6573 18348 6599 18404
rect 6655 18348 6681 18404
rect 6737 18348 6763 18404
rect 6819 18348 6845 18404
rect 6901 18348 6927 18404
rect 6983 18348 7009 18404
rect 7065 18348 7091 18404
rect 7147 18348 7173 18404
rect 7229 18348 7255 18404
rect 7311 18348 7337 18404
rect 7393 18348 7419 18404
rect 7475 18348 7501 18404
rect 7557 18348 7583 18404
rect 7639 18348 7665 18404
rect 7721 18348 7747 18404
rect 7803 18348 7829 18404
rect 7885 18348 7911 18404
rect 7967 18348 7993 18404
rect 8049 18348 8075 18404
rect 8131 18348 8157 18404
rect 8213 18348 8218 18404
rect 5608 18324 8218 18348
rect 5608 18268 5613 18324
rect 5669 18268 5696 18324
rect 5752 18268 5779 18324
rect 5835 18268 5861 18324
rect 5917 18268 5943 18324
rect 5999 18268 6025 18324
rect 6081 18268 6107 18324
rect 6163 18268 6189 18324
rect 6245 18268 6271 18324
rect 6327 18268 6353 18324
rect 6409 18268 6435 18324
rect 6491 18268 6517 18324
rect 6573 18268 6599 18324
rect 6655 18268 6681 18324
rect 6737 18268 6763 18324
rect 6819 18268 6845 18324
rect 6901 18268 6927 18324
rect 6983 18268 7009 18324
rect 7065 18268 7091 18324
rect 7147 18268 7173 18324
rect 7229 18268 7255 18324
rect 7311 18268 7337 18324
rect 7393 18268 7419 18324
rect 7475 18268 7501 18324
rect 7557 18268 7583 18324
rect 7639 18268 7665 18324
rect 7721 18268 7747 18324
rect 7803 18268 7829 18324
rect 7885 18268 7911 18324
rect 7967 18268 7993 18324
rect 8049 18268 8075 18324
rect 8131 18268 8157 18324
rect 8213 18268 8218 18324
rect 5608 18244 8218 18268
rect 5608 18188 5613 18244
rect 5669 18188 5696 18244
rect 5752 18188 5779 18244
rect 5835 18188 5861 18244
rect 5917 18188 5943 18244
rect 5999 18188 6025 18244
rect 6081 18188 6107 18244
rect 6163 18188 6189 18244
rect 6245 18188 6271 18244
rect 6327 18188 6353 18244
rect 6409 18188 6435 18244
rect 6491 18188 6517 18244
rect 6573 18188 6599 18244
rect 6655 18188 6681 18244
rect 6737 18188 6763 18244
rect 6819 18188 6845 18244
rect 6901 18188 6927 18244
rect 6983 18188 7009 18244
rect 7065 18188 7091 18244
rect 7147 18188 7173 18244
rect 7229 18188 7255 18244
rect 7311 18188 7337 18244
rect 7393 18188 7419 18244
rect 7475 18188 7501 18244
rect 7557 18188 7583 18244
rect 7639 18188 7665 18244
rect 7721 18188 7747 18244
rect 7803 18188 7829 18244
rect 7885 18188 7911 18244
rect 7967 18188 7993 18244
rect 8049 18188 8075 18244
rect 8131 18188 8157 18244
rect 8213 18188 8218 18244
rect 5608 18164 8218 18188
rect 5608 18108 5613 18164
rect 5669 18108 5696 18164
rect 5752 18108 5779 18164
rect 5835 18108 5861 18164
rect 5917 18108 5943 18164
rect 5999 18108 6025 18164
rect 6081 18108 6107 18164
rect 6163 18108 6189 18164
rect 6245 18108 6271 18164
rect 6327 18108 6353 18164
rect 6409 18108 6435 18164
rect 6491 18108 6517 18164
rect 6573 18108 6599 18164
rect 6655 18108 6681 18164
rect 6737 18108 6763 18164
rect 6819 18108 6845 18164
rect 6901 18108 6927 18164
rect 6983 18108 7009 18164
rect 7065 18108 7091 18164
rect 7147 18108 7173 18164
rect 7229 18108 7255 18164
rect 7311 18108 7337 18164
rect 7393 18108 7419 18164
rect 7475 18108 7501 18164
rect 7557 18108 7583 18164
rect 7639 18108 7665 18164
rect 7721 18108 7747 18164
rect 7803 18108 7829 18164
rect 7885 18108 7911 18164
rect 7967 18108 7993 18164
rect 8049 18108 8075 18164
rect 8131 18108 8157 18164
rect 8213 18108 8218 18164
rect 5608 15456 8218 18108
rect 5608 15400 5613 15456
rect 5669 15400 5696 15456
rect 5752 15400 5779 15456
rect 5835 15400 5861 15456
rect 5917 15400 5943 15456
rect 5999 15400 6025 15456
rect 6081 15400 6107 15456
rect 6163 15400 6189 15456
rect 6245 15400 6271 15456
rect 6327 15400 6353 15456
rect 6409 15400 6435 15456
rect 6491 15400 6517 15456
rect 6573 15400 6599 15456
rect 6655 15400 6681 15456
rect 6737 15400 6763 15456
rect 6819 15400 6845 15456
rect 6901 15400 6927 15456
rect 6983 15400 7009 15456
rect 7065 15400 7091 15456
rect 7147 15400 7173 15456
rect 7229 15400 7255 15456
rect 7311 15400 7337 15456
rect 7393 15400 7419 15456
rect 7475 15400 7501 15456
rect 7557 15400 7583 15456
rect 7639 15400 7665 15456
rect 7721 15400 7747 15456
rect 7803 15400 7829 15456
rect 7885 15400 7911 15456
rect 7967 15400 7993 15456
rect 8049 15400 8075 15456
rect 8131 15400 8157 15456
rect 8213 15400 8218 15456
rect 5608 15376 8218 15400
rect 5608 15320 5613 15376
rect 5669 15320 5696 15376
rect 5752 15320 5779 15376
rect 5835 15320 5861 15376
rect 5917 15320 5943 15376
rect 5999 15320 6025 15376
rect 6081 15320 6107 15376
rect 6163 15320 6189 15376
rect 6245 15320 6271 15376
rect 6327 15320 6353 15376
rect 6409 15320 6435 15376
rect 6491 15320 6517 15376
rect 6573 15320 6599 15376
rect 6655 15320 6681 15376
rect 6737 15320 6763 15376
rect 6819 15320 6845 15376
rect 6901 15320 6927 15376
rect 6983 15320 7009 15376
rect 7065 15320 7091 15376
rect 7147 15320 7173 15376
rect 7229 15320 7255 15376
rect 7311 15320 7337 15376
rect 7393 15320 7419 15376
rect 7475 15320 7501 15376
rect 7557 15320 7583 15376
rect 7639 15320 7665 15376
rect 7721 15320 7747 15376
rect 7803 15320 7829 15376
rect 7885 15320 7911 15376
rect 7967 15320 7993 15376
rect 8049 15320 8075 15376
rect 8131 15320 8157 15376
rect 8213 15320 8218 15376
rect 5608 15296 8218 15320
rect 5608 15240 5613 15296
rect 5669 15240 5696 15296
rect 5752 15240 5779 15296
rect 5835 15240 5861 15296
rect 5917 15240 5943 15296
rect 5999 15240 6025 15296
rect 6081 15240 6107 15296
rect 6163 15240 6189 15296
rect 6245 15240 6271 15296
rect 6327 15240 6353 15296
rect 6409 15240 6435 15296
rect 6491 15240 6517 15296
rect 6573 15240 6599 15296
rect 6655 15240 6681 15296
rect 6737 15240 6763 15296
rect 6819 15240 6845 15296
rect 6901 15240 6927 15296
rect 6983 15240 7009 15296
rect 7065 15240 7091 15296
rect 7147 15240 7173 15296
rect 7229 15240 7255 15296
rect 7311 15240 7337 15296
rect 7393 15240 7419 15296
rect 7475 15240 7501 15296
rect 7557 15240 7583 15296
rect 7639 15240 7665 15296
rect 7721 15240 7747 15296
rect 7803 15240 7829 15296
rect 7885 15240 7911 15296
rect 7967 15240 7993 15296
rect 8049 15240 8075 15296
rect 8131 15240 8157 15296
rect 8213 15240 8218 15296
rect 5608 15216 8218 15240
rect 5608 15160 5613 15216
rect 5669 15160 5696 15216
rect 5752 15160 5779 15216
rect 5835 15160 5861 15216
rect 5917 15160 5943 15216
rect 5999 15160 6025 15216
rect 6081 15160 6107 15216
rect 6163 15160 6189 15216
rect 6245 15160 6271 15216
rect 6327 15160 6353 15216
rect 6409 15160 6435 15216
rect 6491 15160 6517 15216
rect 6573 15160 6599 15216
rect 6655 15160 6681 15216
rect 6737 15160 6763 15216
rect 6819 15160 6845 15216
rect 6901 15160 6927 15216
rect 6983 15160 7009 15216
rect 7065 15160 7091 15216
rect 7147 15160 7173 15216
rect 7229 15160 7255 15216
rect 7311 15160 7337 15216
rect 7393 15160 7419 15216
rect 7475 15160 7501 15216
rect 7557 15160 7583 15216
rect 7639 15160 7665 15216
rect 7721 15160 7747 15216
rect 7803 15160 7829 15216
rect 7885 15160 7911 15216
rect 7967 15160 7993 15216
rect 8049 15160 8075 15216
rect 8131 15160 8157 15216
rect 8213 15160 8218 15216
rect 5608 15136 8218 15160
rect 5608 15080 5613 15136
rect 5669 15080 5696 15136
rect 5752 15080 5779 15136
rect 5835 15080 5861 15136
rect 5917 15080 5943 15136
rect 5999 15080 6025 15136
rect 6081 15080 6107 15136
rect 6163 15080 6189 15136
rect 6245 15080 6271 15136
rect 6327 15080 6353 15136
rect 6409 15080 6435 15136
rect 6491 15080 6517 15136
rect 6573 15080 6599 15136
rect 6655 15080 6681 15136
rect 6737 15080 6763 15136
rect 6819 15080 6845 15136
rect 6901 15080 6927 15136
rect 6983 15080 7009 15136
rect 7065 15080 7091 15136
rect 7147 15080 7173 15136
rect 7229 15080 7255 15136
rect 7311 15080 7337 15136
rect 7393 15080 7419 15136
rect 7475 15080 7501 15136
rect 7557 15080 7583 15136
rect 7639 15080 7665 15136
rect 7721 15080 7747 15136
rect 7803 15080 7829 15136
rect 7885 15080 7911 15136
rect 7967 15080 7993 15136
rect 8049 15080 8075 15136
rect 8131 15080 8157 15136
rect 8213 15080 8218 15136
rect 5608 15056 8218 15080
rect 5608 15000 5613 15056
rect 5669 15000 5696 15056
rect 5752 15000 5779 15056
rect 5835 15000 5861 15056
rect 5917 15000 5943 15056
rect 5999 15000 6025 15056
rect 6081 15000 6107 15056
rect 6163 15000 6189 15056
rect 6245 15000 6271 15056
rect 6327 15000 6353 15056
rect 6409 15000 6435 15056
rect 6491 15000 6517 15056
rect 6573 15000 6599 15056
rect 6655 15000 6681 15056
rect 6737 15000 6763 15056
rect 6819 15000 6845 15056
rect 6901 15000 6927 15056
rect 6983 15000 7009 15056
rect 7065 15000 7091 15056
rect 7147 15000 7173 15056
rect 7229 15000 7255 15056
rect 7311 15000 7337 15056
rect 7393 15000 7419 15056
rect 7475 15000 7501 15056
rect 7557 15000 7583 15056
rect 7639 15000 7665 15056
rect 7721 15000 7747 15056
rect 7803 15000 7829 15056
rect 7885 15000 7911 15056
rect 7967 15000 7993 15056
rect 8049 15000 8075 15056
rect 8131 15000 8157 15056
rect 8213 15000 8218 15056
rect 5608 14976 8218 15000
rect 5608 14920 5613 14976
rect 5669 14920 5696 14976
rect 5752 14920 5779 14976
rect 5835 14920 5861 14976
rect 5917 14920 5943 14976
rect 5999 14920 6025 14976
rect 6081 14920 6107 14976
rect 6163 14920 6189 14976
rect 6245 14920 6271 14976
rect 6327 14920 6353 14976
rect 6409 14920 6435 14976
rect 6491 14920 6517 14976
rect 6573 14920 6599 14976
rect 6655 14920 6681 14976
rect 6737 14920 6763 14976
rect 6819 14920 6845 14976
rect 6901 14920 6927 14976
rect 6983 14920 7009 14976
rect 7065 14920 7091 14976
rect 7147 14920 7173 14976
rect 7229 14920 7255 14976
rect 7311 14920 7337 14976
rect 7393 14920 7419 14976
rect 7475 14920 7501 14976
rect 7557 14920 7583 14976
rect 7639 14920 7665 14976
rect 7721 14920 7747 14976
rect 7803 14920 7829 14976
rect 7885 14920 7911 14976
rect 7967 14920 7993 14976
rect 8049 14920 8075 14976
rect 8131 14920 8157 14976
rect 8213 14920 8218 14976
rect 5608 14896 8218 14920
rect 5608 14840 5613 14896
rect 5669 14840 5696 14896
rect 5752 14840 5779 14896
rect 5835 14840 5861 14896
rect 5917 14840 5943 14896
rect 5999 14840 6025 14896
rect 6081 14840 6107 14896
rect 6163 14840 6189 14896
rect 6245 14840 6271 14896
rect 6327 14840 6353 14896
rect 6409 14840 6435 14896
rect 6491 14840 6517 14896
rect 6573 14840 6599 14896
rect 6655 14840 6681 14896
rect 6737 14840 6763 14896
rect 6819 14840 6845 14896
rect 6901 14840 6927 14896
rect 6983 14840 7009 14896
rect 7065 14840 7091 14896
rect 7147 14840 7173 14896
rect 7229 14840 7255 14896
rect 7311 14840 7337 14896
rect 7393 14840 7419 14896
rect 7475 14840 7501 14896
rect 7557 14840 7583 14896
rect 7639 14840 7665 14896
rect 7721 14840 7747 14896
rect 7803 14840 7829 14896
rect 7885 14840 7911 14896
rect 7967 14840 7993 14896
rect 8049 14840 8075 14896
rect 8131 14840 8157 14896
rect 8213 14840 8218 14896
rect 5608 13456 8218 14840
rect 5608 13400 5613 13456
rect 5669 13400 5696 13456
rect 5752 13400 5779 13456
rect 5835 13400 5861 13456
rect 5917 13400 5943 13456
rect 5999 13400 6025 13456
rect 6081 13400 6107 13456
rect 6163 13400 6189 13456
rect 6245 13400 6271 13456
rect 6327 13400 6353 13456
rect 6409 13400 6435 13456
rect 6491 13400 6517 13456
rect 6573 13400 6599 13456
rect 6655 13400 6681 13456
rect 6737 13400 6763 13456
rect 6819 13400 6845 13456
rect 6901 13400 6927 13456
rect 6983 13400 7009 13456
rect 7065 13400 7091 13456
rect 7147 13400 7173 13456
rect 7229 13400 7255 13456
rect 7311 13400 7337 13456
rect 7393 13400 7419 13456
rect 7475 13400 7501 13456
rect 7557 13400 7583 13456
rect 7639 13400 7665 13456
rect 7721 13400 7747 13456
rect 7803 13400 7829 13456
rect 7885 13400 7911 13456
rect 7967 13400 7993 13456
rect 8049 13400 8075 13456
rect 8131 13400 8157 13456
rect 8213 13400 8218 13456
rect 5608 13376 8218 13400
rect 5608 13320 5613 13376
rect 5669 13320 5696 13376
rect 5752 13320 5779 13376
rect 5835 13320 5861 13376
rect 5917 13320 5943 13376
rect 5999 13320 6025 13376
rect 6081 13320 6107 13376
rect 6163 13320 6189 13376
rect 6245 13320 6271 13376
rect 6327 13320 6353 13376
rect 6409 13320 6435 13376
rect 6491 13320 6517 13376
rect 6573 13320 6599 13376
rect 6655 13320 6681 13376
rect 6737 13320 6763 13376
rect 6819 13320 6845 13376
rect 6901 13320 6927 13376
rect 6983 13320 7009 13376
rect 7065 13320 7091 13376
rect 7147 13320 7173 13376
rect 7229 13320 7255 13376
rect 7311 13320 7337 13376
rect 7393 13320 7419 13376
rect 7475 13320 7501 13376
rect 7557 13320 7583 13376
rect 7639 13320 7665 13376
rect 7721 13320 7747 13376
rect 7803 13320 7829 13376
rect 7885 13320 7911 13376
rect 7967 13320 7993 13376
rect 8049 13320 8075 13376
rect 8131 13320 8157 13376
rect 8213 13320 8218 13376
rect 5608 13296 8218 13320
rect 5608 13240 5613 13296
rect 5669 13240 5696 13296
rect 5752 13240 5779 13296
rect 5835 13240 5861 13296
rect 5917 13240 5943 13296
rect 5999 13240 6025 13296
rect 6081 13240 6107 13296
rect 6163 13240 6189 13296
rect 6245 13240 6271 13296
rect 6327 13240 6353 13296
rect 6409 13240 6435 13296
rect 6491 13240 6517 13296
rect 6573 13240 6599 13296
rect 6655 13240 6681 13296
rect 6737 13240 6763 13296
rect 6819 13240 6845 13296
rect 6901 13240 6927 13296
rect 6983 13240 7009 13296
rect 7065 13240 7091 13296
rect 7147 13240 7173 13296
rect 7229 13240 7255 13296
rect 7311 13240 7337 13296
rect 7393 13240 7419 13296
rect 7475 13240 7501 13296
rect 7557 13240 7583 13296
rect 7639 13240 7665 13296
rect 7721 13240 7747 13296
rect 7803 13240 7829 13296
rect 7885 13240 7911 13296
rect 7967 13240 7993 13296
rect 8049 13240 8075 13296
rect 8131 13240 8157 13296
rect 8213 13240 8218 13296
rect 5608 13216 8218 13240
rect 5608 13160 5613 13216
rect 5669 13160 5696 13216
rect 5752 13160 5779 13216
rect 5835 13160 5861 13216
rect 5917 13160 5943 13216
rect 5999 13160 6025 13216
rect 6081 13160 6107 13216
rect 6163 13160 6189 13216
rect 6245 13160 6271 13216
rect 6327 13160 6353 13216
rect 6409 13160 6435 13216
rect 6491 13160 6517 13216
rect 6573 13160 6599 13216
rect 6655 13160 6681 13216
rect 6737 13160 6763 13216
rect 6819 13160 6845 13216
rect 6901 13160 6927 13216
rect 6983 13160 7009 13216
rect 7065 13160 7091 13216
rect 7147 13160 7173 13216
rect 7229 13160 7255 13216
rect 7311 13160 7337 13216
rect 7393 13160 7419 13216
rect 7475 13160 7501 13216
rect 7557 13160 7583 13216
rect 7639 13160 7665 13216
rect 7721 13160 7747 13216
rect 7803 13160 7829 13216
rect 7885 13160 7911 13216
rect 7967 13160 7993 13216
rect 8049 13160 8075 13216
rect 8131 13160 8157 13216
rect 8213 13160 8218 13216
rect 5608 13136 8218 13160
rect 5608 13080 5613 13136
rect 5669 13080 5696 13136
rect 5752 13080 5779 13136
rect 5835 13080 5861 13136
rect 5917 13080 5943 13136
rect 5999 13080 6025 13136
rect 6081 13080 6107 13136
rect 6163 13080 6189 13136
rect 6245 13080 6271 13136
rect 6327 13080 6353 13136
rect 6409 13080 6435 13136
rect 6491 13080 6517 13136
rect 6573 13080 6599 13136
rect 6655 13080 6681 13136
rect 6737 13080 6763 13136
rect 6819 13080 6845 13136
rect 6901 13080 6927 13136
rect 6983 13080 7009 13136
rect 7065 13080 7091 13136
rect 7147 13080 7173 13136
rect 7229 13080 7255 13136
rect 7311 13080 7337 13136
rect 7393 13080 7419 13136
rect 7475 13080 7501 13136
rect 7557 13080 7583 13136
rect 7639 13080 7665 13136
rect 7721 13080 7747 13136
rect 7803 13080 7829 13136
rect 7885 13080 7911 13136
rect 7967 13080 7993 13136
rect 8049 13080 8075 13136
rect 8131 13080 8157 13136
rect 8213 13080 8218 13136
rect 5608 13056 8218 13080
rect 5608 13000 5613 13056
rect 5669 13000 5696 13056
rect 5752 13000 5779 13056
rect 5835 13000 5861 13056
rect 5917 13000 5943 13056
rect 5999 13000 6025 13056
rect 6081 13000 6107 13056
rect 6163 13000 6189 13056
rect 6245 13000 6271 13056
rect 6327 13000 6353 13056
rect 6409 13000 6435 13056
rect 6491 13000 6517 13056
rect 6573 13000 6599 13056
rect 6655 13000 6681 13056
rect 6737 13000 6763 13056
rect 6819 13000 6845 13056
rect 6901 13000 6927 13056
rect 6983 13000 7009 13056
rect 7065 13000 7091 13056
rect 7147 13000 7173 13056
rect 7229 13000 7255 13056
rect 7311 13000 7337 13056
rect 7393 13000 7419 13056
rect 7475 13000 7501 13056
rect 7557 13000 7583 13056
rect 7639 13000 7665 13056
rect 7721 13000 7747 13056
rect 7803 13000 7829 13056
rect 7885 13000 7911 13056
rect 7967 13000 7993 13056
rect 8049 13000 8075 13056
rect 8131 13000 8157 13056
rect 8213 13000 8218 13056
rect 5608 12976 8218 13000
rect 5608 12920 5613 12976
rect 5669 12920 5696 12976
rect 5752 12920 5779 12976
rect 5835 12920 5861 12976
rect 5917 12920 5943 12976
rect 5999 12920 6025 12976
rect 6081 12920 6107 12976
rect 6163 12920 6189 12976
rect 6245 12920 6271 12976
rect 6327 12920 6353 12976
rect 6409 12920 6435 12976
rect 6491 12920 6517 12976
rect 6573 12920 6599 12976
rect 6655 12920 6681 12976
rect 6737 12920 6763 12976
rect 6819 12920 6845 12976
rect 6901 12920 6927 12976
rect 6983 12920 7009 12976
rect 7065 12920 7091 12976
rect 7147 12920 7173 12976
rect 7229 12920 7255 12976
rect 7311 12920 7337 12976
rect 7393 12920 7419 12976
rect 7475 12920 7501 12976
rect 7557 12920 7583 12976
rect 7639 12920 7665 12976
rect 7721 12920 7747 12976
rect 7803 12920 7829 12976
rect 7885 12920 7911 12976
rect 7967 12920 7993 12976
rect 8049 12920 8075 12976
rect 8131 12920 8157 12976
rect 8213 12920 8218 12976
rect 5608 12896 8218 12920
rect 5608 12840 5613 12896
rect 5669 12840 5696 12896
rect 5752 12840 5779 12896
rect 5835 12840 5861 12896
rect 5917 12840 5943 12896
rect 5999 12840 6025 12896
rect 6081 12840 6107 12896
rect 6163 12840 6189 12896
rect 6245 12840 6271 12896
rect 6327 12840 6353 12896
rect 6409 12840 6435 12896
rect 6491 12840 6517 12896
rect 6573 12840 6599 12896
rect 6655 12840 6681 12896
rect 6737 12840 6763 12896
rect 6819 12840 6845 12896
rect 6901 12840 6927 12896
rect 6983 12840 7009 12896
rect 7065 12840 7091 12896
rect 7147 12840 7173 12896
rect 7229 12840 7255 12896
rect 7311 12840 7337 12896
rect 7393 12840 7419 12896
rect 7475 12840 7501 12896
rect 7557 12840 7583 12896
rect 7639 12840 7665 12896
rect 7721 12840 7747 12896
rect 7803 12840 7829 12896
rect 7885 12840 7911 12896
rect 7967 12840 7993 12896
rect 8049 12840 8075 12896
rect 8131 12840 8157 12896
rect 8213 12840 8218 12896
rect 5608 11456 8218 12840
rect 5608 11400 5613 11456
rect 5669 11400 5696 11456
rect 5752 11400 5779 11456
rect 5835 11400 5861 11456
rect 5917 11400 5943 11456
rect 5999 11400 6025 11456
rect 6081 11400 6107 11456
rect 6163 11400 6189 11456
rect 6245 11400 6271 11456
rect 6327 11400 6353 11456
rect 6409 11400 6435 11456
rect 6491 11400 6517 11456
rect 6573 11400 6599 11456
rect 6655 11400 6681 11456
rect 6737 11400 6763 11456
rect 6819 11400 6845 11456
rect 6901 11400 6927 11456
rect 6983 11400 7009 11456
rect 7065 11400 7091 11456
rect 7147 11400 7173 11456
rect 7229 11400 7255 11456
rect 7311 11400 7337 11456
rect 7393 11400 7419 11456
rect 7475 11400 7501 11456
rect 7557 11400 7583 11456
rect 7639 11400 7665 11456
rect 7721 11400 7747 11456
rect 7803 11400 7829 11456
rect 7885 11400 7911 11456
rect 7967 11400 7993 11456
rect 8049 11400 8075 11456
rect 8131 11400 8157 11456
rect 8213 11400 8218 11456
rect 5608 11376 8218 11400
rect 5608 11320 5613 11376
rect 5669 11320 5696 11376
rect 5752 11320 5779 11376
rect 5835 11320 5861 11376
rect 5917 11320 5943 11376
rect 5999 11320 6025 11376
rect 6081 11320 6107 11376
rect 6163 11320 6189 11376
rect 6245 11320 6271 11376
rect 6327 11320 6353 11376
rect 6409 11320 6435 11376
rect 6491 11320 6517 11376
rect 6573 11320 6599 11376
rect 6655 11320 6681 11376
rect 6737 11320 6763 11376
rect 6819 11320 6845 11376
rect 6901 11320 6927 11376
rect 6983 11320 7009 11376
rect 7065 11320 7091 11376
rect 7147 11320 7173 11376
rect 7229 11320 7255 11376
rect 7311 11320 7337 11376
rect 7393 11320 7419 11376
rect 7475 11320 7501 11376
rect 7557 11320 7583 11376
rect 7639 11320 7665 11376
rect 7721 11320 7747 11376
rect 7803 11320 7829 11376
rect 7885 11320 7911 11376
rect 7967 11320 7993 11376
rect 8049 11320 8075 11376
rect 8131 11320 8157 11376
rect 8213 11320 8218 11376
rect 5608 11296 8218 11320
rect 5608 11240 5613 11296
rect 5669 11240 5696 11296
rect 5752 11240 5779 11296
rect 5835 11240 5861 11296
rect 5917 11240 5943 11296
rect 5999 11240 6025 11296
rect 6081 11240 6107 11296
rect 6163 11240 6189 11296
rect 6245 11240 6271 11296
rect 6327 11240 6353 11296
rect 6409 11240 6435 11296
rect 6491 11240 6517 11296
rect 6573 11240 6599 11296
rect 6655 11240 6681 11296
rect 6737 11240 6763 11296
rect 6819 11240 6845 11296
rect 6901 11240 6927 11296
rect 6983 11240 7009 11296
rect 7065 11240 7091 11296
rect 7147 11240 7173 11296
rect 7229 11240 7255 11296
rect 7311 11240 7337 11296
rect 7393 11240 7419 11296
rect 7475 11240 7501 11296
rect 7557 11240 7583 11296
rect 7639 11240 7665 11296
rect 7721 11240 7747 11296
rect 7803 11240 7829 11296
rect 7885 11240 7911 11296
rect 7967 11240 7993 11296
rect 8049 11240 8075 11296
rect 8131 11240 8157 11296
rect 8213 11240 8218 11296
rect 5608 11216 8218 11240
rect 5608 11160 5613 11216
rect 5669 11160 5696 11216
rect 5752 11160 5779 11216
rect 5835 11160 5861 11216
rect 5917 11160 5943 11216
rect 5999 11160 6025 11216
rect 6081 11160 6107 11216
rect 6163 11160 6189 11216
rect 6245 11160 6271 11216
rect 6327 11160 6353 11216
rect 6409 11160 6435 11216
rect 6491 11160 6517 11216
rect 6573 11160 6599 11216
rect 6655 11160 6681 11216
rect 6737 11160 6763 11216
rect 6819 11160 6845 11216
rect 6901 11160 6927 11216
rect 6983 11160 7009 11216
rect 7065 11160 7091 11216
rect 7147 11160 7173 11216
rect 7229 11160 7255 11216
rect 7311 11160 7337 11216
rect 7393 11160 7419 11216
rect 7475 11160 7501 11216
rect 7557 11160 7583 11216
rect 7639 11160 7665 11216
rect 7721 11160 7747 11216
rect 7803 11160 7829 11216
rect 7885 11160 7911 11216
rect 7967 11160 7993 11216
rect 8049 11160 8075 11216
rect 8131 11160 8157 11216
rect 8213 11160 8218 11216
rect 5608 11136 8218 11160
rect 5608 11080 5613 11136
rect 5669 11080 5696 11136
rect 5752 11080 5779 11136
rect 5835 11080 5861 11136
rect 5917 11080 5943 11136
rect 5999 11080 6025 11136
rect 6081 11080 6107 11136
rect 6163 11080 6189 11136
rect 6245 11080 6271 11136
rect 6327 11080 6353 11136
rect 6409 11080 6435 11136
rect 6491 11080 6517 11136
rect 6573 11080 6599 11136
rect 6655 11080 6681 11136
rect 6737 11080 6763 11136
rect 6819 11080 6845 11136
rect 6901 11080 6927 11136
rect 6983 11080 7009 11136
rect 7065 11080 7091 11136
rect 7147 11080 7173 11136
rect 7229 11080 7255 11136
rect 7311 11080 7337 11136
rect 7393 11080 7419 11136
rect 7475 11080 7501 11136
rect 7557 11080 7583 11136
rect 7639 11080 7665 11136
rect 7721 11080 7747 11136
rect 7803 11080 7829 11136
rect 7885 11080 7911 11136
rect 7967 11080 7993 11136
rect 8049 11080 8075 11136
rect 8131 11080 8157 11136
rect 8213 11080 8218 11136
rect 5608 11056 8218 11080
rect 5608 11000 5613 11056
rect 5669 11000 5696 11056
rect 5752 11000 5779 11056
rect 5835 11000 5861 11056
rect 5917 11000 5943 11056
rect 5999 11000 6025 11056
rect 6081 11000 6107 11056
rect 6163 11000 6189 11056
rect 6245 11000 6271 11056
rect 6327 11000 6353 11056
rect 6409 11000 6435 11056
rect 6491 11000 6517 11056
rect 6573 11000 6599 11056
rect 6655 11000 6681 11056
rect 6737 11000 6763 11056
rect 6819 11000 6845 11056
rect 6901 11000 6927 11056
rect 6983 11000 7009 11056
rect 7065 11000 7091 11056
rect 7147 11000 7173 11056
rect 7229 11000 7255 11056
rect 7311 11000 7337 11056
rect 7393 11000 7419 11056
rect 7475 11000 7501 11056
rect 7557 11000 7583 11056
rect 7639 11000 7665 11056
rect 7721 11000 7747 11056
rect 7803 11000 7829 11056
rect 7885 11000 7911 11056
rect 7967 11000 7993 11056
rect 8049 11000 8075 11056
rect 8131 11000 8157 11056
rect 8213 11000 8218 11056
rect 5608 10976 8218 11000
rect 5608 10920 5613 10976
rect 5669 10920 5696 10976
rect 5752 10920 5779 10976
rect 5835 10920 5861 10976
rect 5917 10920 5943 10976
rect 5999 10920 6025 10976
rect 6081 10920 6107 10976
rect 6163 10920 6189 10976
rect 6245 10920 6271 10976
rect 6327 10920 6353 10976
rect 6409 10920 6435 10976
rect 6491 10920 6517 10976
rect 6573 10920 6599 10976
rect 6655 10920 6681 10976
rect 6737 10920 6763 10976
rect 6819 10920 6845 10976
rect 6901 10920 6927 10976
rect 6983 10920 7009 10976
rect 7065 10920 7091 10976
rect 7147 10920 7173 10976
rect 7229 10920 7255 10976
rect 7311 10920 7337 10976
rect 7393 10920 7419 10976
rect 7475 10920 7501 10976
rect 7557 10920 7583 10976
rect 7639 10920 7665 10976
rect 7721 10920 7747 10976
rect 7803 10920 7829 10976
rect 7885 10920 7911 10976
rect 7967 10920 7993 10976
rect 8049 10920 8075 10976
rect 8131 10920 8157 10976
rect 8213 10920 8218 10976
rect 5608 10896 8218 10920
rect 5608 10840 5613 10896
rect 5669 10840 5696 10896
rect 5752 10840 5779 10896
rect 5835 10840 5861 10896
rect 5917 10840 5943 10896
rect 5999 10840 6025 10896
rect 6081 10840 6107 10896
rect 6163 10840 6189 10896
rect 6245 10840 6271 10896
rect 6327 10840 6353 10896
rect 6409 10840 6435 10896
rect 6491 10840 6517 10896
rect 6573 10840 6599 10896
rect 6655 10840 6681 10896
rect 6737 10840 6763 10896
rect 6819 10840 6845 10896
rect 6901 10840 6927 10896
rect 6983 10840 7009 10896
rect 7065 10840 7091 10896
rect 7147 10840 7173 10896
rect 7229 10840 7255 10896
rect 7311 10840 7337 10896
rect 7393 10840 7419 10896
rect 7475 10840 7501 10896
rect 7557 10840 7583 10896
rect 7639 10840 7665 10896
rect 7721 10840 7747 10896
rect 7803 10840 7829 10896
rect 7885 10840 7911 10896
rect 7967 10840 7993 10896
rect 8049 10840 8075 10896
rect 8131 10840 8157 10896
rect 8213 10840 8218 10896
rect 5608 9460 8218 10840
rect 5608 9404 5617 9460
rect 5673 9404 5698 9460
rect 5754 9404 5779 9460
rect 5835 9404 5860 9460
rect 5916 9404 5941 9460
rect 5997 9404 6022 9460
rect 6078 9404 6103 9460
rect 6159 9404 6184 9460
rect 6240 9404 6265 9460
rect 6321 9404 6346 9460
rect 6402 9404 6427 9460
rect 6483 9404 6508 9460
rect 6564 9404 6589 9460
rect 6645 9404 6669 9460
rect 6725 9404 6749 9460
rect 6805 9404 6829 9460
rect 6885 9404 6909 9460
rect 6965 9404 6989 9460
rect 7045 9404 7069 9460
rect 7125 9404 7149 9460
rect 7205 9404 7229 9460
rect 7285 9404 7309 9460
rect 7365 9404 8218 9460
rect 5608 8713 8218 9404
rect 5608 8657 5621 8713
rect 5677 8657 5705 8713
rect 5761 8657 5789 8713
rect 5845 8657 5873 8713
rect 5929 8657 5957 8713
rect 6013 8657 6041 8713
rect 6097 8657 6125 8713
rect 6181 8657 6209 8713
rect 6265 8657 6293 8713
rect 6349 8657 6377 8713
rect 6433 8657 6461 8713
rect 6517 8657 6545 8713
rect 6601 8657 6629 8713
rect 6685 8657 6713 8713
rect 6769 8657 6797 8713
rect 6853 8657 6881 8713
rect 6937 8657 6965 8713
rect 7021 8657 7048 8713
rect 7104 8657 7131 8713
rect 7187 8657 7214 8713
rect 7270 8657 7297 8713
rect 7353 8657 8218 8713
rect 5608 8633 8218 8657
rect 5608 8577 5621 8633
rect 5677 8577 5705 8633
rect 5761 8577 5789 8633
rect 5845 8577 5873 8633
rect 5929 8577 5957 8633
rect 6013 8577 6041 8633
rect 6097 8577 6125 8633
rect 6181 8577 6209 8633
rect 6265 8577 6293 8633
rect 6349 8577 6377 8633
rect 6433 8577 6461 8633
rect 6517 8577 6545 8633
rect 6601 8577 6629 8633
rect 6685 8577 6713 8633
rect 6769 8577 6797 8633
rect 6853 8577 6881 8633
rect 6937 8577 6965 8633
rect 7021 8577 7048 8633
rect 7104 8577 7131 8633
rect 7187 8577 7214 8633
rect 7270 8577 7297 8633
rect 7353 8577 8218 8633
rect 5608 8553 8218 8577
rect 5608 8497 5621 8553
rect 5677 8497 5705 8553
rect 5761 8497 5789 8553
rect 5845 8497 5873 8553
rect 5929 8497 5957 8553
rect 6013 8497 6041 8553
rect 6097 8497 6125 8553
rect 6181 8497 6209 8553
rect 6265 8497 6293 8553
rect 6349 8497 6377 8553
rect 6433 8497 6461 8553
rect 6517 8497 6545 8553
rect 6601 8497 6629 8553
rect 6685 8497 6713 8553
rect 6769 8497 6797 8553
rect 6853 8497 6881 8553
rect 6937 8497 6965 8553
rect 7021 8497 7048 8553
rect 7104 8497 7131 8553
rect 7187 8497 7214 8553
rect 7270 8497 7297 8553
rect 7353 8497 8218 8553
rect 5608 8473 8218 8497
rect 5608 8417 5621 8473
rect 5677 8417 5705 8473
rect 5761 8417 5789 8473
rect 5845 8417 5873 8473
rect 5929 8417 5957 8473
rect 6013 8417 6041 8473
rect 6097 8417 6125 8473
rect 6181 8417 6209 8473
rect 6265 8417 6293 8473
rect 6349 8417 6377 8473
rect 6433 8417 6461 8473
rect 6517 8417 6545 8473
rect 6601 8417 6629 8473
rect 6685 8417 6713 8473
rect 6769 8417 6797 8473
rect 6853 8417 6881 8473
rect 6937 8417 6965 8473
rect 7021 8417 7048 8473
rect 7104 8417 7131 8473
rect 7187 8417 7214 8473
rect 7270 8417 7297 8473
rect 7353 8417 8218 8473
rect 5608 8393 8218 8417
rect 5608 8337 5621 8393
rect 5677 8337 5705 8393
rect 5761 8337 5789 8393
rect 5845 8337 5873 8393
rect 5929 8337 5957 8393
rect 6013 8337 6041 8393
rect 6097 8337 6125 8393
rect 6181 8337 6209 8393
rect 6265 8337 6293 8393
rect 6349 8337 6377 8393
rect 6433 8337 6461 8393
rect 6517 8337 6545 8393
rect 6601 8337 6629 8393
rect 6685 8337 6713 8393
rect 6769 8337 6797 8393
rect 6853 8337 6881 8393
rect 6937 8337 6965 8393
rect 7021 8337 7048 8393
rect 7104 8337 7131 8393
rect 7187 8337 7214 8393
rect 7270 8337 7297 8393
rect 7353 8337 8218 8393
rect 5608 8313 8218 8337
rect 5608 8257 5621 8313
rect 5677 8257 5705 8313
rect 5761 8257 5789 8313
rect 5845 8257 5873 8313
rect 5929 8257 5957 8313
rect 6013 8257 6041 8313
rect 6097 8257 6125 8313
rect 6181 8257 6209 8313
rect 6265 8257 6293 8313
rect 6349 8257 6377 8313
rect 6433 8257 6461 8313
rect 6517 8257 6545 8313
rect 6601 8257 6629 8313
rect 6685 8257 6713 8313
rect 6769 8257 6797 8313
rect 6853 8257 6881 8313
rect 6937 8257 6965 8313
rect 7021 8257 7048 8313
rect 7104 8257 7131 8313
rect 7187 8257 7214 8313
rect 7270 8257 7297 8313
rect 7353 8257 8218 8313
rect 5608 8233 8218 8257
rect 5608 8177 5621 8233
rect 5677 8177 5705 8233
rect 5761 8177 5789 8233
rect 5845 8177 5873 8233
rect 5929 8177 5957 8233
rect 6013 8177 6041 8233
rect 6097 8177 6125 8233
rect 6181 8177 6209 8233
rect 6265 8177 6293 8233
rect 6349 8177 6377 8233
rect 6433 8177 6461 8233
rect 6517 8177 6545 8233
rect 6601 8177 6629 8233
rect 6685 8177 6713 8233
rect 6769 8177 6797 8233
rect 6853 8177 6881 8233
rect 6937 8177 6965 8233
rect 7021 8177 7048 8233
rect 7104 8177 7131 8233
rect 7187 8177 7214 8233
rect 7270 8177 7297 8233
rect 7353 8177 8218 8233
rect 5608 8153 8218 8177
rect 5608 8097 5621 8153
rect 5677 8097 5705 8153
rect 5761 8097 5789 8153
rect 5845 8097 5873 8153
rect 5929 8097 5957 8153
rect 6013 8097 6041 8153
rect 6097 8097 6125 8153
rect 6181 8097 6209 8153
rect 6265 8097 6293 8153
rect 6349 8097 6377 8153
rect 6433 8097 6461 8153
rect 6517 8097 6545 8153
rect 6601 8097 6629 8153
rect 6685 8097 6713 8153
rect 6769 8097 6797 8153
rect 6853 8097 6881 8153
rect 6937 8097 6965 8153
rect 7021 8097 7048 8153
rect 7104 8097 7131 8153
rect 7187 8097 7214 8153
rect 7270 8097 7297 8153
rect 7353 8097 8218 8153
rect 5608 8073 8218 8097
rect 5608 8017 5621 8073
rect 5677 8017 5705 8073
rect 5761 8017 5789 8073
rect 5845 8017 5873 8073
rect 5929 8017 5957 8073
rect 6013 8017 6041 8073
rect 6097 8017 6125 8073
rect 6181 8017 6209 8073
rect 6265 8017 6293 8073
rect 6349 8017 6377 8073
rect 6433 8017 6461 8073
rect 6517 8017 6545 8073
rect 6601 8017 6629 8073
rect 6685 8017 6713 8073
rect 6769 8017 6797 8073
rect 6853 8017 6881 8073
rect 6937 8017 6965 8073
rect 7021 8017 7048 8073
rect 7104 8017 7131 8073
rect 7187 8017 7214 8073
rect 7270 8017 7297 8073
rect 7353 8017 8218 8073
rect 5608 7993 8218 8017
rect 5608 7937 5621 7993
rect 5677 7937 5705 7993
rect 5761 7937 5789 7993
rect 5845 7937 5873 7993
rect 5929 7937 5957 7993
rect 6013 7937 6041 7993
rect 6097 7937 6125 7993
rect 6181 7937 6209 7993
rect 6265 7937 6293 7993
rect 6349 7937 6377 7993
rect 6433 7937 6461 7993
rect 6517 7937 6545 7993
rect 6601 7937 6629 7993
rect 6685 7937 6713 7993
rect 6769 7937 6797 7993
rect 6853 7937 6881 7993
rect 6937 7937 6965 7993
rect 7021 7937 7048 7993
rect 7104 7937 7131 7993
rect 7187 7937 7214 7993
rect 7270 7937 7297 7993
rect 7353 7937 8218 7993
rect 5608 7913 8218 7937
rect 5608 7857 5621 7913
rect 5677 7857 5705 7913
rect 5761 7857 5789 7913
rect 5845 7857 5873 7913
rect 5929 7857 5957 7913
rect 6013 7857 6041 7913
rect 6097 7857 6125 7913
rect 6181 7857 6209 7913
rect 6265 7857 6293 7913
rect 6349 7857 6377 7913
rect 6433 7857 6461 7913
rect 6517 7857 6545 7913
rect 6601 7857 6629 7913
rect 6685 7857 6713 7913
rect 6769 7857 6797 7913
rect 6853 7857 6881 7913
rect 6937 7857 6965 7913
rect 7021 7857 7048 7913
rect 7104 7857 7131 7913
rect 7187 7857 7214 7913
rect 7270 7857 7297 7913
rect 7353 7857 8218 7913
rect 5608 7692 8218 7857
rect 5608 7636 5617 7692
rect 5673 7636 5698 7692
rect 5754 7636 5779 7692
rect 5835 7636 5860 7692
rect 5916 7636 5941 7692
rect 5997 7636 6022 7692
rect 6078 7636 6103 7692
rect 6159 7636 6184 7692
rect 6240 7636 6265 7692
rect 6321 7636 6346 7692
rect 6402 7636 6427 7692
rect 6483 7636 6508 7692
rect 6564 7636 6589 7692
rect 6645 7636 6669 7692
rect 6725 7636 6749 7692
rect 6805 7636 6829 7692
rect 6885 7636 6909 7692
rect 6965 7636 6989 7692
rect 7045 7636 7069 7692
rect 7125 7636 7149 7692
rect 7205 7636 7229 7692
rect 7285 7636 7309 7692
rect 7365 7636 8218 7692
rect 5608 6915 8218 7636
rect 5608 6859 5621 6915
rect 5677 6859 5705 6915
rect 5761 6859 5789 6915
rect 5845 6859 5873 6915
rect 5929 6859 5957 6915
rect 6013 6859 6041 6915
rect 6097 6859 6125 6915
rect 6181 6859 6209 6915
rect 6265 6859 6293 6915
rect 6349 6859 6377 6915
rect 6433 6859 6461 6915
rect 6517 6859 6545 6915
rect 6601 6859 6629 6915
rect 6685 6859 6713 6915
rect 6769 6859 6797 6915
rect 6853 6859 6881 6915
rect 6937 6859 6965 6915
rect 7021 6859 7048 6915
rect 7104 6859 7131 6915
rect 7187 6859 7214 6915
rect 7270 6859 7297 6915
rect 7353 6859 8218 6915
rect 5608 6835 8218 6859
rect 5608 6779 5621 6835
rect 5677 6779 5705 6835
rect 5761 6779 5789 6835
rect 5845 6779 5873 6835
rect 5929 6779 5957 6835
rect 6013 6779 6041 6835
rect 6097 6779 6125 6835
rect 6181 6779 6209 6835
rect 6265 6779 6293 6835
rect 6349 6779 6377 6835
rect 6433 6779 6461 6835
rect 6517 6779 6545 6835
rect 6601 6779 6629 6835
rect 6685 6779 6713 6835
rect 6769 6779 6797 6835
rect 6853 6779 6881 6835
rect 6937 6779 6965 6835
rect 7021 6779 7048 6835
rect 7104 6779 7131 6835
rect 7187 6779 7214 6835
rect 7270 6779 7297 6835
rect 7353 6779 8218 6835
rect 5608 6755 8218 6779
rect 5608 6699 5621 6755
rect 5677 6699 5705 6755
rect 5761 6699 5789 6755
rect 5845 6699 5873 6755
rect 5929 6699 5957 6755
rect 6013 6699 6041 6755
rect 6097 6699 6125 6755
rect 6181 6699 6209 6755
rect 6265 6699 6293 6755
rect 6349 6699 6377 6755
rect 6433 6699 6461 6755
rect 6517 6699 6545 6755
rect 6601 6699 6629 6755
rect 6685 6699 6713 6755
rect 6769 6699 6797 6755
rect 6853 6699 6881 6755
rect 6937 6699 6965 6755
rect 7021 6699 7048 6755
rect 7104 6699 7131 6755
rect 7187 6699 7214 6755
rect 7270 6699 7297 6755
rect 7353 6699 8218 6755
rect 5608 6675 8218 6699
rect 5608 6619 5621 6675
rect 5677 6619 5705 6675
rect 5761 6619 5789 6675
rect 5845 6619 5873 6675
rect 5929 6619 5957 6675
rect 6013 6619 6041 6675
rect 6097 6619 6125 6675
rect 6181 6619 6209 6675
rect 6265 6619 6293 6675
rect 6349 6619 6377 6675
rect 6433 6619 6461 6675
rect 6517 6619 6545 6675
rect 6601 6619 6629 6675
rect 6685 6619 6713 6675
rect 6769 6619 6797 6675
rect 6853 6619 6881 6675
rect 6937 6619 6965 6675
rect 7021 6619 7048 6675
rect 7104 6619 7131 6675
rect 7187 6619 7214 6675
rect 7270 6619 7297 6675
rect 7353 6619 8218 6675
rect 5608 6595 8218 6619
rect 5608 6539 5621 6595
rect 5677 6539 5705 6595
rect 5761 6539 5789 6595
rect 5845 6539 5873 6595
rect 5929 6539 5957 6595
rect 6013 6539 6041 6595
rect 6097 6539 6125 6595
rect 6181 6539 6209 6595
rect 6265 6539 6293 6595
rect 6349 6539 6377 6595
rect 6433 6539 6461 6595
rect 6517 6539 6545 6595
rect 6601 6539 6629 6595
rect 6685 6539 6713 6595
rect 6769 6539 6797 6595
rect 6853 6539 6881 6595
rect 6937 6539 6965 6595
rect 7021 6539 7048 6595
rect 7104 6539 7131 6595
rect 7187 6539 7214 6595
rect 7270 6539 7297 6595
rect 7353 6539 8218 6595
rect 5608 6515 8218 6539
rect 5608 6459 5621 6515
rect 5677 6459 5705 6515
rect 5761 6459 5789 6515
rect 5845 6459 5873 6515
rect 5929 6459 5957 6515
rect 6013 6459 6041 6515
rect 6097 6459 6125 6515
rect 6181 6459 6209 6515
rect 6265 6459 6293 6515
rect 6349 6459 6377 6515
rect 6433 6459 6461 6515
rect 6517 6459 6545 6515
rect 6601 6459 6629 6515
rect 6685 6459 6713 6515
rect 6769 6459 6797 6515
rect 6853 6459 6881 6515
rect 6937 6459 6965 6515
rect 7021 6459 7048 6515
rect 7104 6459 7131 6515
rect 7187 6459 7214 6515
rect 7270 6459 7297 6515
rect 7353 6459 8218 6515
rect 5608 6435 8218 6459
rect 5608 6379 5621 6435
rect 5677 6379 5705 6435
rect 5761 6379 5789 6435
rect 5845 6379 5873 6435
rect 5929 6379 5957 6435
rect 6013 6379 6041 6435
rect 6097 6379 6125 6435
rect 6181 6379 6209 6435
rect 6265 6379 6293 6435
rect 6349 6379 6377 6435
rect 6433 6379 6461 6435
rect 6517 6379 6545 6435
rect 6601 6379 6629 6435
rect 6685 6379 6713 6435
rect 6769 6379 6797 6435
rect 6853 6379 6881 6435
rect 6937 6379 6965 6435
rect 7021 6379 7048 6435
rect 7104 6379 7131 6435
rect 7187 6379 7214 6435
rect 7270 6379 7297 6435
rect 7353 6379 8218 6435
rect 5608 6355 8218 6379
rect 5608 6299 5621 6355
rect 5677 6299 5705 6355
rect 5761 6299 5789 6355
rect 5845 6299 5873 6355
rect 5929 6299 5957 6355
rect 6013 6299 6041 6355
rect 6097 6299 6125 6355
rect 6181 6299 6209 6355
rect 6265 6299 6293 6355
rect 6349 6299 6377 6355
rect 6433 6299 6461 6355
rect 6517 6299 6545 6355
rect 6601 6299 6629 6355
rect 6685 6299 6713 6355
rect 6769 6299 6797 6355
rect 6853 6299 6881 6355
rect 6937 6299 6965 6355
rect 7021 6299 7048 6355
rect 7104 6299 7131 6355
rect 7187 6299 7214 6355
rect 7270 6299 7297 6355
rect 7353 6299 8218 6355
rect 5608 6275 8218 6299
rect 5608 6219 5621 6275
rect 5677 6219 5705 6275
rect 5761 6219 5789 6275
rect 5845 6219 5873 6275
rect 5929 6219 5957 6275
rect 6013 6219 6041 6275
rect 6097 6219 6125 6275
rect 6181 6219 6209 6275
rect 6265 6219 6293 6275
rect 6349 6219 6377 6275
rect 6433 6219 6461 6275
rect 6517 6219 6545 6275
rect 6601 6219 6629 6275
rect 6685 6219 6713 6275
rect 6769 6219 6797 6275
rect 6853 6219 6881 6275
rect 6937 6219 6965 6275
rect 7021 6219 7048 6275
rect 7104 6219 7131 6275
rect 7187 6219 7214 6275
rect 7270 6219 7297 6275
rect 7353 6219 8218 6275
rect 5608 6195 8218 6219
rect 5608 6139 5621 6195
rect 5677 6139 5705 6195
rect 5761 6139 5789 6195
rect 5845 6139 5873 6195
rect 5929 6139 5957 6195
rect 6013 6139 6041 6195
rect 6097 6139 6125 6195
rect 6181 6139 6209 6195
rect 6265 6139 6293 6195
rect 6349 6139 6377 6195
rect 6433 6139 6461 6195
rect 6517 6139 6545 6195
rect 6601 6139 6629 6195
rect 6685 6139 6713 6195
rect 6769 6139 6797 6195
rect 6853 6139 6881 6195
rect 6937 6139 6965 6195
rect 7021 6139 7048 6195
rect 7104 6139 7131 6195
rect 7187 6139 7214 6195
rect 7270 6139 7297 6195
rect 7353 6139 8218 6195
rect 5608 6115 8218 6139
rect 5608 6059 5621 6115
rect 5677 6059 5705 6115
rect 5761 6059 5789 6115
rect 5845 6059 5873 6115
rect 5929 6059 5957 6115
rect 6013 6059 6041 6115
rect 6097 6059 6125 6115
rect 6181 6059 6209 6115
rect 6265 6059 6293 6115
rect 6349 6059 6377 6115
rect 6433 6059 6461 6115
rect 6517 6059 6545 6115
rect 6601 6059 6629 6115
rect 6685 6059 6713 6115
rect 6769 6059 6797 6115
rect 6853 6059 6881 6115
rect 6937 6059 6965 6115
rect 7021 6059 7048 6115
rect 7104 6059 7131 6115
rect 7187 6059 7214 6115
rect 7270 6059 7297 6115
rect 7353 6059 8218 6115
rect 5608 5852 8218 6059
rect 5608 5796 5617 5852
rect 5673 5796 5698 5852
rect 5754 5796 5779 5852
rect 5835 5796 5860 5852
rect 5916 5796 5941 5852
rect 5997 5796 6022 5852
rect 6078 5796 6103 5852
rect 6159 5796 6184 5852
rect 6240 5796 6265 5852
rect 6321 5796 6346 5852
rect 6402 5796 6427 5852
rect 6483 5796 6508 5852
rect 6564 5796 6589 5852
rect 6645 5796 6669 5852
rect 6725 5796 6749 5852
rect 6805 5796 6829 5852
rect 6885 5796 6909 5852
rect 6965 5796 6989 5852
rect 7045 5796 7069 5852
rect 7125 5796 7149 5852
rect 7205 5796 7229 5852
rect 7285 5796 7309 5852
rect 7365 5796 8218 5852
rect 5608 4741 8218 5796
rect 5608 4685 5623 4741
rect 5679 4685 5704 4741
rect 5760 4685 5785 4741
rect 5841 4685 5866 4741
rect 5922 4685 5947 4741
rect 6003 4685 6027 4741
rect 6083 4685 6107 4741
rect 6163 4685 6187 4741
rect 6243 4685 6267 4741
rect 6323 4685 6347 4741
rect 6403 4685 6427 4741
rect 6483 4685 6507 4741
rect 6563 4685 6587 4741
rect 6643 4685 6667 4741
rect 6723 4685 6747 4741
rect 6803 4685 6827 4741
rect 6883 4685 6907 4741
rect 6963 4685 6987 4741
rect 7043 4685 7067 4741
rect 7123 4685 7147 4741
rect 7203 4685 7227 4741
rect 7283 4685 7307 4741
rect 7363 4685 8218 4741
rect 5608 4653 8218 4685
rect 5608 4597 5623 4653
rect 5679 4597 5704 4653
rect 5760 4597 5785 4653
rect 5841 4597 5866 4653
rect 5922 4597 5947 4653
rect 6003 4597 6027 4653
rect 6083 4597 6107 4653
rect 6163 4597 6187 4653
rect 6243 4597 6267 4653
rect 6323 4597 6347 4653
rect 6403 4597 6427 4653
rect 6483 4597 6507 4653
rect 6563 4597 6587 4653
rect 6643 4597 6667 4653
rect 6723 4597 6747 4653
rect 6803 4597 6827 4653
rect 6883 4597 6907 4653
rect 6963 4597 6987 4653
rect 7043 4597 7067 4653
rect 7123 4597 7147 4653
rect 7203 4597 7227 4653
rect 7283 4597 7307 4653
rect 7363 4597 8218 4653
rect 5608 4565 8218 4597
rect 5608 4509 5623 4565
rect 5679 4509 5704 4565
rect 5760 4509 5785 4565
rect 5841 4509 5866 4565
rect 5922 4509 5947 4565
rect 6003 4509 6027 4565
rect 6083 4509 6107 4565
rect 6163 4509 6187 4565
rect 6243 4509 6267 4565
rect 6323 4509 6347 4565
rect 6403 4509 6427 4565
rect 6483 4509 6507 4565
rect 6563 4509 6587 4565
rect 6643 4509 6667 4565
rect 6723 4509 6747 4565
rect 6803 4509 6827 4565
rect 6883 4509 6907 4565
rect 6963 4509 6987 4565
rect 7043 4509 7067 4565
rect 7123 4509 7147 4565
rect 7203 4509 7227 4565
rect 7283 4509 7307 4565
rect 7363 4509 8218 4565
rect 5608 4477 8218 4509
rect 5608 4421 5623 4477
rect 5679 4421 5704 4477
rect 5760 4421 5785 4477
rect 5841 4421 5866 4477
rect 5922 4421 5947 4477
rect 6003 4421 6027 4477
rect 6083 4421 6107 4477
rect 6163 4421 6187 4477
rect 6243 4421 6267 4477
rect 6323 4421 6347 4477
rect 6403 4421 6427 4477
rect 6483 4421 6507 4477
rect 6563 4421 6587 4477
rect 6643 4421 6667 4477
rect 6723 4421 6747 4477
rect 6803 4421 6827 4477
rect 6883 4421 6907 4477
rect 6963 4421 6987 4477
rect 7043 4421 7067 4477
rect 7123 4421 7147 4477
rect 7203 4421 7227 4477
rect 7283 4421 7307 4477
rect 7363 4421 8218 4477
rect 5608 4389 8218 4421
rect 5608 4333 5623 4389
rect 5679 4333 5704 4389
rect 5760 4333 5785 4389
rect 5841 4333 5866 4389
rect 5922 4333 5947 4389
rect 6003 4333 6027 4389
rect 6083 4333 6107 4389
rect 6163 4333 6187 4389
rect 6243 4333 6267 4389
rect 6323 4333 6347 4389
rect 6403 4333 6427 4389
rect 6483 4333 6507 4389
rect 6563 4333 6587 4389
rect 6643 4333 6667 4389
rect 6723 4333 6747 4389
rect 6803 4333 6827 4389
rect 6883 4333 6907 4389
rect 6963 4333 6987 4389
rect 7043 4333 7067 4389
rect 7123 4333 7147 4389
rect 7203 4333 7227 4389
rect 7283 4333 7307 4389
rect 7363 4333 8218 4389
rect 5608 4301 8218 4333
rect 5608 4245 5623 4301
rect 5679 4245 5704 4301
rect 5760 4245 5785 4301
rect 5841 4245 5866 4301
rect 5922 4245 5947 4301
rect 6003 4245 6027 4301
rect 6083 4245 6107 4301
rect 6163 4245 6187 4301
rect 6243 4245 6267 4301
rect 6323 4245 6347 4301
rect 6403 4245 6427 4301
rect 6483 4245 6507 4301
rect 6563 4245 6587 4301
rect 6643 4245 6667 4301
rect 6723 4245 6747 4301
rect 6803 4245 6827 4301
rect 6883 4245 6907 4301
rect 6963 4245 6987 4301
rect 7043 4245 7067 4301
rect 7123 4245 7147 4301
rect 7203 4245 7227 4301
rect 7283 4245 7307 4301
rect 7363 4245 8218 4301
rect 5608 4213 8218 4245
rect 5608 4157 5623 4213
rect 5679 4157 5704 4213
rect 5760 4157 5785 4213
rect 5841 4157 5866 4213
rect 5922 4157 5947 4213
rect 6003 4157 6027 4213
rect 6083 4157 6107 4213
rect 6163 4157 6187 4213
rect 6243 4157 6267 4213
rect 6323 4157 6347 4213
rect 6403 4157 6427 4213
rect 6483 4157 6507 4213
rect 6563 4157 6587 4213
rect 6643 4157 6667 4213
rect 6723 4157 6747 4213
rect 6803 4157 6827 4213
rect 6883 4157 6907 4213
rect 6963 4157 6987 4213
rect 7043 4157 7067 4213
rect 7123 4157 7147 4213
rect 7203 4157 7227 4213
rect 7283 4157 7307 4213
rect 7363 4157 8218 4213
rect 5608 3918 8218 4157
rect 5608 3862 5617 3918
rect 5673 3862 5698 3918
rect 5754 3862 5779 3918
rect 5835 3862 5860 3918
rect 5916 3862 5941 3918
rect 5997 3862 6022 3918
rect 6078 3862 6103 3918
rect 6159 3862 6184 3918
rect 6240 3862 6265 3918
rect 6321 3862 6346 3918
rect 6402 3862 6427 3918
rect 6483 3862 6508 3918
rect 6564 3862 6589 3918
rect 6645 3862 6669 3918
rect 6725 3862 6749 3918
rect 6805 3862 6829 3918
rect 6885 3862 6909 3918
rect 6965 3862 6989 3918
rect 7045 3862 7069 3918
rect 7125 3862 7149 3918
rect 7205 3862 7229 3918
rect 7285 3862 7309 3918
rect 7365 3862 8218 3918
rect 5608 3057 8218 3862
rect 5608 3001 5617 3057
rect 5673 3001 5698 3057
rect 5754 3001 5779 3057
rect 5835 3001 5860 3057
rect 5916 3001 5941 3057
rect 5997 3001 6022 3057
rect 6078 3001 6103 3057
rect 6159 3001 6184 3057
rect 6240 3001 6265 3057
rect 6321 3001 6346 3057
rect 6402 3001 6427 3057
rect 6483 3001 6508 3057
rect 6564 3001 6589 3057
rect 6645 3001 6670 3057
rect 6726 3001 6751 3057
rect 6807 3001 6832 3057
rect 6888 3001 6913 3057
rect 6969 3001 6994 3057
rect 7050 3001 7075 3057
rect 7131 3001 7156 3057
rect 7212 3001 7237 3057
rect 7293 3001 7317 3057
rect 7373 3001 7397 3057
rect 7453 3001 7477 3057
rect 7533 3001 8218 3057
rect 5608 2967 8218 3001
rect 5608 2911 5617 2967
rect 5673 2911 5698 2967
rect 5754 2911 5779 2967
rect 5835 2911 5860 2967
rect 5916 2911 5941 2967
rect 5997 2911 6022 2967
rect 6078 2911 6103 2967
rect 6159 2911 6184 2967
rect 6240 2911 6265 2967
rect 6321 2911 6346 2967
rect 6402 2911 6427 2967
rect 6483 2911 6508 2967
rect 6564 2911 6589 2967
rect 6645 2911 6670 2967
rect 6726 2911 6751 2967
rect 6807 2911 6832 2967
rect 6888 2911 6913 2967
rect 6969 2911 6994 2967
rect 7050 2911 7075 2967
rect 7131 2911 7156 2967
rect 7212 2911 7237 2967
rect 7293 2911 7317 2967
rect 7373 2911 7397 2967
rect 7453 2911 7477 2967
rect 7533 2911 8218 2967
rect 5608 2877 8218 2911
rect 5608 2821 5617 2877
rect 5673 2821 5698 2877
rect 5754 2821 5779 2877
rect 5835 2821 5860 2877
rect 5916 2821 5941 2877
rect 5997 2821 6022 2877
rect 6078 2821 6103 2877
rect 6159 2821 6184 2877
rect 6240 2821 6265 2877
rect 6321 2821 6346 2877
rect 6402 2821 6427 2877
rect 6483 2821 6508 2877
rect 6564 2821 6589 2877
rect 6645 2821 6670 2877
rect 6726 2821 6751 2877
rect 6807 2821 6832 2877
rect 6888 2821 6913 2877
rect 6969 2821 6994 2877
rect 7050 2821 7075 2877
rect 7131 2821 7156 2877
rect 7212 2821 7237 2877
rect 7293 2821 7317 2877
rect 7373 2821 7397 2877
rect 7453 2821 7477 2877
rect 7533 2821 8218 2877
rect 5608 2787 8218 2821
rect 5608 2731 5617 2787
rect 5673 2731 5698 2787
rect 5754 2731 5779 2787
rect 5835 2731 5860 2787
rect 5916 2731 5941 2787
rect 5997 2731 6022 2787
rect 6078 2731 6103 2787
rect 6159 2731 6184 2787
rect 6240 2731 6265 2787
rect 6321 2731 6346 2787
rect 6402 2731 6427 2787
rect 6483 2731 6508 2787
rect 6564 2731 6589 2787
rect 6645 2731 6670 2787
rect 6726 2731 6751 2787
rect 6807 2731 6832 2787
rect 6888 2731 6913 2787
rect 6969 2731 6994 2787
rect 7050 2731 7075 2787
rect 7131 2731 7156 2787
rect 7212 2731 7237 2787
rect 7293 2731 7317 2787
rect 7373 2731 7397 2787
rect 7453 2731 7477 2787
rect 7533 2731 8218 2787
rect 5608 2697 8218 2731
rect 5608 2641 5617 2697
rect 5673 2641 5698 2697
rect 5754 2641 5779 2697
rect 5835 2641 5860 2697
rect 5916 2641 5941 2697
rect 5997 2641 6022 2697
rect 6078 2641 6103 2697
rect 6159 2641 6184 2697
rect 6240 2641 6265 2697
rect 6321 2641 6346 2697
rect 6402 2641 6427 2697
rect 6483 2641 6508 2697
rect 6564 2641 6589 2697
rect 6645 2641 6670 2697
rect 6726 2641 6751 2697
rect 6807 2641 6832 2697
rect 6888 2641 6913 2697
rect 6969 2641 6994 2697
rect 7050 2641 7075 2697
rect 7131 2641 7156 2697
rect 7212 2641 7237 2697
rect 7293 2641 7317 2697
rect 7373 2641 7397 2697
rect 7453 2641 7477 2697
rect 7533 2641 8218 2697
rect 5608 2607 8218 2641
rect 5608 2551 5617 2607
rect 5673 2551 5698 2607
rect 5754 2551 5779 2607
rect 5835 2551 5860 2607
rect 5916 2551 5941 2607
rect 5997 2551 6022 2607
rect 6078 2551 6103 2607
rect 6159 2551 6184 2607
rect 6240 2551 6265 2607
rect 6321 2551 6346 2607
rect 6402 2551 6427 2607
rect 6483 2551 6508 2607
rect 6564 2551 6589 2607
rect 6645 2551 6670 2607
rect 6726 2551 6751 2607
rect 6807 2551 6832 2607
rect 6888 2551 6913 2607
rect 6969 2551 6994 2607
rect 7050 2551 7075 2607
rect 7131 2551 7156 2607
rect 7212 2551 7237 2607
rect 7293 2551 7317 2607
rect 7373 2551 7397 2607
rect 7453 2551 7477 2607
rect 7533 2551 8218 2607
rect 5608 2517 8218 2551
rect 5608 2461 5617 2517
rect 5673 2461 5698 2517
rect 5754 2461 5779 2517
rect 5835 2461 5860 2517
rect 5916 2461 5941 2517
rect 5997 2461 6022 2517
rect 6078 2461 6103 2517
rect 6159 2461 6184 2517
rect 6240 2461 6265 2517
rect 6321 2461 6346 2517
rect 6402 2461 6427 2517
rect 6483 2461 6508 2517
rect 6564 2461 6589 2517
rect 6645 2461 6670 2517
rect 6726 2461 6751 2517
rect 6807 2461 6832 2517
rect 6888 2461 6913 2517
rect 6969 2461 6994 2517
rect 7050 2461 7075 2517
rect 7131 2461 7156 2517
rect 7212 2461 7237 2517
rect 7293 2461 7317 2517
rect 7373 2461 7397 2517
rect 7453 2461 7477 2517
rect 7533 2461 8218 2517
rect 5608 2239 8218 2461
rect 5608 2225 6615 2239
rect 5608 2169 5624 2225
rect 5680 2169 5704 2225
rect 5760 2169 5784 2225
rect 5840 2169 5864 2225
rect 5920 2169 5944 2225
rect 6000 2169 6024 2225
rect 6080 2169 6104 2225
rect 6160 2169 6184 2225
rect 6240 2169 6264 2225
rect 6320 2183 6615 2225
rect 6671 2183 6701 2239
rect 6757 2183 6787 2239
rect 6843 2183 6873 2239
rect 6929 2183 6959 2239
rect 7015 2183 7045 2239
rect 7101 2183 7131 2239
rect 7187 2183 7217 2239
rect 7273 2183 7303 2239
rect 7359 2183 8218 2239
rect 6320 2169 8218 2183
rect 5608 2157 8218 2169
rect 5608 2143 6615 2157
rect 5608 2087 5624 2143
rect 5680 2087 5704 2143
rect 5760 2087 5784 2143
rect 5840 2087 5864 2143
rect 5920 2087 5944 2143
rect 6000 2087 6024 2143
rect 6080 2087 6104 2143
rect 6160 2087 6184 2143
rect 6240 2087 6264 2143
rect 6320 2101 6615 2143
rect 6671 2101 6701 2157
rect 6757 2101 6787 2157
rect 6843 2101 6873 2157
rect 6929 2101 6959 2157
rect 7015 2101 7045 2157
rect 7101 2101 7131 2157
rect 7187 2101 7217 2157
rect 7273 2101 7303 2157
rect 7359 2101 8218 2157
rect 6320 2087 8218 2101
rect 5608 2075 8218 2087
rect 5608 2061 6615 2075
rect 5608 2005 5624 2061
rect 5680 2005 5704 2061
rect 5760 2005 5784 2061
rect 5840 2005 5864 2061
rect 5920 2005 5944 2061
rect 6000 2005 6024 2061
rect 6080 2005 6104 2061
rect 6160 2005 6184 2061
rect 6240 2005 6264 2061
rect 6320 2019 6615 2061
rect 6671 2019 6701 2075
rect 6757 2019 6787 2075
rect 6843 2019 6873 2075
rect 6929 2019 6959 2075
rect 7015 2019 7045 2075
rect 7101 2019 7131 2075
rect 7187 2019 7217 2075
rect 7273 2019 7303 2075
rect 7359 2019 8218 2075
rect 6320 2005 8218 2019
rect 5608 1993 8218 2005
rect 5608 1979 6615 1993
rect 5608 1923 5624 1979
rect 5680 1923 5704 1979
rect 5760 1923 5784 1979
rect 5840 1923 5864 1979
rect 5920 1923 5944 1979
rect 6000 1923 6024 1979
rect 6080 1923 6104 1979
rect 6160 1923 6184 1979
rect 6240 1923 6264 1979
rect 6320 1937 6615 1979
rect 6671 1937 6701 1993
rect 6757 1937 6787 1993
rect 6843 1937 6873 1993
rect 6929 1937 6959 1993
rect 7015 1937 7045 1993
rect 7101 1937 7131 1993
rect 7187 1937 7217 1993
rect 7273 1937 7303 1993
rect 7359 1937 8218 1993
rect 6320 1923 8218 1937
rect 5608 1911 8218 1923
rect 5608 1897 6615 1911
rect 5608 1841 5624 1897
rect 5680 1841 5704 1897
rect 5760 1841 5784 1897
rect 5840 1841 5864 1897
rect 5920 1841 5944 1897
rect 6000 1841 6024 1897
rect 6080 1841 6104 1897
rect 6160 1841 6184 1897
rect 6240 1841 6264 1897
rect 6320 1855 6615 1897
rect 6671 1855 6701 1911
rect 6757 1855 6787 1911
rect 6843 1855 6873 1911
rect 6929 1855 6959 1911
rect 7015 1855 7045 1911
rect 7101 1855 7131 1911
rect 7187 1855 7217 1911
rect 7273 1855 7303 1911
rect 7359 1855 8218 1911
rect 6320 1841 8218 1855
rect 5608 1828 8218 1841
rect 5608 1815 6615 1828
rect 5608 1759 5624 1815
rect 5680 1759 5704 1815
rect 5760 1759 5784 1815
rect 5840 1759 5864 1815
rect 5920 1759 5944 1815
rect 6000 1759 6024 1815
rect 6080 1759 6104 1815
rect 6160 1759 6184 1815
rect 6240 1759 6264 1815
rect 6320 1772 6615 1815
rect 6671 1772 6701 1828
rect 6757 1772 6787 1828
rect 6843 1772 6873 1828
rect 6929 1772 6959 1828
rect 7015 1772 7045 1828
rect 7101 1772 7131 1828
rect 7187 1772 7217 1828
rect 7273 1772 7303 1828
rect 7359 1772 8218 1828
rect 6320 1759 8218 1772
rect 5608 1745 8218 1759
rect 5608 1733 6615 1745
rect 5608 1677 5624 1733
rect 5680 1677 5704 1733
rect 5760 1677 5784 1733
rect 5840 1677 5864 1733
rect 5920 1677 5944 1733
rect 6000 1677 6024 1733
rect 6080 1677 6104 1733
rect 6160 1677 6184 1733
rect 6240 1677 6264 1733
rect 6320 1689 6615 1733
rect 6671 1689 6701 1745
rect 6757 1689 6787 1745
rect 6843 1689 6873 1745
rect 6929 1689 6959 1745
rect 7015 1689 7045 1745
rect 7101 1689 7131 1745
rect 7187 1689 7217 1745
rect 7273 1689 7303 1745
rect 7359 1689 8218 1745
rect 6320 1677 8218 1689
rect 5608 1662 8218 1677
rect 5608 1651 6615 1662
rect 5608 1595 5624 1651
rect 5680 1595 5704 1651
rect 5760 1595 5784 1651
rect 5840 1595 5864 1651
rect 5920 1595 5944 1651
rect 6000 1595 6024 1651
rect 6080 1595 6104 1651
rect 6160 1595 6184 1651
rect 6240 1595 6264 1651
rect 6320 1606 6615 1651
rect 6671 1606 6701 1662
rect 6757 1606 6787 1662
rect 6843 1606 6873 1662
rect 6929 1606 6959 1662
rect 7015 1606 7045 1662
rect 7101 1606 7131 1662
rect 7187 1606 7217 1662
rect 7273 1606 7303 1662
rect 7359 1606 8218 1662
rect 6320 1595 8218 1606
rect 5608 1579 8218 1595
rect 5608 1569 6615 1579
rect 5608 1513 5624 1569
rect 5680 1513 5704 1569
rect 5760 1513 5784 1569
rect 5840 1513 5864 1569
rect 5920 1513 5944 1569
rect 6000 1513 6024 1569
rect 6080 1513 6104 1569
rect 6160 1513 6184 1569
rect 6240 1513 6264 1569
rect 6320 1523 6615 1569
rect 6671 1523 6701 1579
rect 6757 1523 6787 1579
rect 6843 1523 6873 1579
rect 6929 1523 6959 1579
rect 7015 1523 7045 1579
rect 7101 1523 7131 1579
rect 7187 1523 7217 1579
rect 7273 1523 7303 1579
rect 7359 1523 8218 1579
rect 6320 1513 8218 1523
rect 5608 1496 8218 1513
rect 5608 1487 6615 1496
rect 5608 1431 5624 1487
rect 5680 1431 5704 1487
rect 5760 1431 5784 1487
rect 5840 1431 5864 1487
rect 5920 1431 5944 1487
rect 6000 1431 6024 1487
rect 6080 1431 6104 1487
rect 6160 1431 6184 1487
rect 6240 1431 6264 1487
rect 6320 1440 6615 1487
rect 6671 1440 6701 1496
rect 6757 1440 6787 1496
rect 6843 1440 6873 1496
rect 6929 1440 6959 1496
rect 7015 1440 7045 1496
rect 7101 1440 7131 1496
rect 7187 1440 7217 1496
rect 7273 1440 7303 1496
rect 7359 1440 8218 1496
rect 6320 1431 8218 1440
rect 5608 1413 8218 1431
rect 5608 1405 6615 1413
rect 5608 1349 5624 1405
rect 5680 1349 5704 1405
rect 5760 1349 5784 1405
rect 5840 1349 5864 1405
rect 5920 1349 5944 1405
rect 6000 1349 6024 1405
rect 6080 1349 6104 1405
rect 6160 1349 6184 1405
rect 6240 1349 6264 1405
rect 6320 1357 6615 1405
rect 6671 1357 6701 1413
rect 6757 1357 6787 1413
rect 6843 1357 6873 1413
rect 6929 1357 6959 1413
rect 7015 1357 7045 1413
rect 7101 1357 7131 1413
rect 7187 1357 7217 1413
rect 7273 1357 7303 1413
rect 7359 1357 8218 1413
rect 6320 1349 8218 1357
rect 5608 1330 8218 1349
rect 5608 1323 6615 1330
rect 5608 1267 5624 1323
rect 5680 1267 5704 1323
rect 5760 1267 5784 1323
rect 5840 1267 5864 1323
rect 5920 1267 5944 1323
rect 6000 1267 6024 1323
rect 6080 1267 6104 1323
rect 6160 1267 6184 1323
rect 6240 1267 6264 1323
rect 6320 1274 6615 1323
rect 6671 1274 6701 1330
rect 6757 1274 6787 1330
rect 6843 1274 6873 1330
rect 6929 1274 6959 1330
rect 7015 1274 7045 1330
rect 7101 1274 7131 1330
rect 7187 1274 7217 1330
rect 7273 1274 7303 1330
rect 7359 1274 8218 1330
rect 6320 1267 8218 1274
rect 5608 1247 8218 1267
rect 5608 1241 6615 1247
rect 5608 1185 5624 1241
rect 5680 1185 5704 1241
rect 5760 1185 5784 1241
rect 5840 1185 5864 1241
rect 5920 1185 5944 1241
rect 6000 1185 6024 1241
rect 6080 1185 6104 1241
rect 6160 1185 6184 1241
rect 6240 1185 6264 1241
rect 6320 1191 6615 1241
rect 6671 1191 6701 1247
rect 6757 1191 6787 1247
rect 6843 1191 6873 1247
rect 6929 1191 6959 1247
rect 7015 1191 7045 1247
rect 7101 1191 7131 1247
rect 7187 1191 7217 1247
rect 7273 1191 7303 1247
rect 7359 1191 8218 1247
rect 6320 1185 8218 1191
rect 5608 1164 8218 1185
rect 5608 1159 6615 1164
rect 5608 1103 5624 1159
rect 5680 1103 5704 1159
rect 5760 1103 5784 1159
rect 5840 1103 5864 1159
rect 5920 1103 5944 1159
rect 6000 1103 6024 1159
rect 6080 1103 6104 1159
rect 6160 1103 6184 1159
rect 6240 1103 6264 1159
rect 6320 1108 6615 1159
rect 6671 1108 6701 1164
rect 6757 1108 6787 1164
rect 6843 1108 6873 1164
rect 6929 1108 6959 1164
rect 7015 1108 7045 1164
rect 7101 1108 7131 1164
rect 7187 1108 7217 1164
rect 7273 1108 7303 1164
rect 7359 1108 8218 1164
rect 6320 1103 8218 1108
rect 5608 1081 8218 1103
rect 5608 1077 6615 1081
rect 5608 1021 5624 1077
rect 5680 1021 5704 1077
rect 5760 1021 5784 1077
rect 5840 1021 5864 1077
rect 5920 1021 5944 1077
rect 6000 1021 6024 1077
rect 6080 1021 6104 1077
rect 6160 1021 6184 1077
rect 6240 1021 6264 1077
rect 6320 1025 6615 1077
rect 6671 1025 6701 1081
rect 6757 1025 6787 1081
rect 6843 1025 6873 1081
rect 6929 1025 6959 1081
rect 7015 1025 7045 1081
rect 7101 1025 7131 1081
rect 7187 1025 7217 1081
rect 7273 1025 7303 1081
rect 7359 1025 8218 1081
rect 6320 1021 8218 1025
rect 5608 998 8218 1021
rect 5608 994 6615 998
rect 5608 938 5624 994
rect 5680 938 5704 994
rect 5760 938 5784 994
rect 5840 938 5864 994
rect 5920 938 5944 994
rect 6000 938 6024 994
rect 6080 938 6104 994
rect 6160 938 6184 994
rect 6240 938 6264 994
rect 6320 942 6615 994
rect 6671 942 6701 998
rect 6757 942 6787 998
rect 6843 942 6873 998
rect 6929 942 6959 998
rect 7015 942 7045 998
rect 7101 942 7131 998
rect 7187 942 7217 998
rect 7273 942 7303 998
rect 7359 942 8218 998
rect 6320 938 8218 942
rect 5608 915 8218 938
rect 5608 911 6615 915
rect 5608 855 5624 911
rect 5680 855 5704 911
rect 5760 855 5784 911
rect 5840 855 5864 911
rect 5920 855 5944 911
rect 6000 855 6024 911
rect 6080 855 6104 911
rect 6160 855 6184 911
rect 6240 855 6264 911
rect 6320 859 6615 911
rect 6671 859 6701 915
rect 6757 859 6787 915
rect 6843 859 6873 915
rect 6929 859 6959 915
rect 7015 859 7045 915
rect 7101 859 7131 915
rect 7187 859 7217 915
rect 7273 859 7303 915
rect 7359 859 8218 915
rect 6320 855 8218 859
rect 5608 832 8218 855
rect 5608 828 6615 832
rect 5608 772 5624 828
rect 5680 772 5704 828
rect 5760 772 5784 828
rect 5840 772 5864 828
rect 5920 772 5944 828
rect 6000 772 6024 828
rect 6080 772 6104 828
rect 6160 772 6184 828
rect 6240 772 6264 828
rect 6320 776 6615 828
rect 6671 776 6701 832
rect 6757 776 6787 832
rect 6843 776 6873 832
rect 6929 776 6959 832
rect 7015 776 7045 832
rect 7101 776 7131 832
rect 7187 776 7217 832
rect 7273 776 7303 832
rect 7359 776 8218 832
rect 6320 772 8218 776
rect 5608 749 8218 772
rect 5608 745 6615 749
rect 5608 689 5624 745
rect 5680 689 5704 745
rect 5760 689 5784 745
rect 5840 689 5864 745
rect 5920 689 5944 745
rect 6000 689 6024 745
rect 6080 689 6104 745
rect 6160 689 6184 745
rect 6240 689 6264 745
rect 6320 693 6615 745
rect 6671 693 6701 749
rect 6757 693 6787 749
rect 6843 693 6873 749
rect 6929 693 6959 749
rect 7015 693 7045 749
rect 7101 693 7131 749
rect 7187 693 7217 749
rect 7273 693 7303 749
rect 7359 693 8218 749
rect 6320 689 8218 693
rect 5608 666 8218 689
rect 5608 662 6615 666
rect 5608 606 5624 662
rect 5680 606 5704 662
rect 5760 606 5784 662
rect 5840 606 5864 662
rect 5920 606 5944 662
rect 6000 606 6024 662
rect 6080 606 6104 662
rect 6160 606 6184 662
rect 6240 606 6264 662
rect 6320 610 6615 662
rect 6671 610 6701 666
rect 6757 610 6787 666
rect 6843 610 6873 666
rect 6929 610 6959 666
rect 7015 610 7045 666
rect 7101 610 7131 666
rect 7187 610 7217 666
rect 7273 610 7303 666
rect 7359 610 8218 666
rect 6320 606 8218 610
rect 5608 583 8218 606
rect 5608 579 6615 583
rect 5608 523 5624 579
rect 5680 523 5704 579
rect 5760 523 5784 579
rect 5840 523 5864 579
rect 5920 523 5944 579
rect 6000 523 6024 579
rect 6080 523 6104 579
rect 6160 523 6184 579
rect 6240 523 6264 579
rect 6320 527 6615 579
rect 6671 527 6701 583
rect 6757 527 6787 583
rect 6843 527 6873 583
rect 6929 527 6959 583
rect 7015 527 7045 583
rect 7101 527 7131 583
rect 7187 527 7217 583
rect 7273 527 7303 583
rect 7359 527 8218 583
rect 6320 523 8218 527
rect 5608 500 8218 523
rect 5608 496 6615 500
rect 5608 440 5624 496
rect 5680 440 5704 496
rect 5760 440 5784 496
rect 5840 440 5864 496
rect 5920 440 5944 496
rect 6000 440 6024 496
rect 6080 440 6104 496
rect 6160 440 6184 496
rect 6240 440 6264 496
rect 6320 444 6615 496
rect 6671 444 6701 500
rect 6757 444 6787 500
rect 6843 444 6873 500
rect 6929 444 6959 500
rect 7015 444 7045 500
rect 7101 444 7131 500
rect 7187 444 7217 500
rect 7273 444 7303 500
rect 7359 444 8218 500
rect 6320 440 8218 444
rect 5608 0 8218 440
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_0
timestamp 1704896540
transform 1 0 6493 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_1
timestamp 1704896540
transform 1 0 5939 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_2
timestamp 1704896540
transform 1 0 6425 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_3
timestamp 1704896540
transform 1 0 5871 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_4
timestamp 1704896540
transform 1 0 5385 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_5
timestamp 1704896540
transform 1 0 5317 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_6
timestamp 1704896540
transform 1 0 4831 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_7
timestamp 1704896540
transform 1 0 4763 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_8
timestamp 1704896540
transform 1 0 4277 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_9
timestamp 1704896540
transform 1 0 3723 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_10
timestamp 1704896540
transform 1 0 3655 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_11
timestamp 1704896540
transform 1 0 3169 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_12
timestamp 1704896540
transform 1 0 3101 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_13
timestamp 1704896540
transform 1 0 4209 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_14
timestamp 1704896540
transform 1 0 6493 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_15
timestamp 1704896540
transform 1 0 6493 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_16
timestamp 1704896540
transform 1 0 6493 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_17
timestamp 1704896540
transform 1 0 5939 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_18
timestamp 1704896540
transform 1 0 5939 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_19
timestamp 1704896540
transform 1 0 5939 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_20
timestamp 1704896540
transform 1 0 6425 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_21
timestamp 1704896540
transform 1 0 6425 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_22
timestamp 1704896540
transform 1 0 6425 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_23
timestamp 1704896540
transform 1 0 5871 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_24
timestamp 1704896540
transform 1 0 5871 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_25
timestamp 1704896540
transform 1 0 5871 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_26
timestamp 1704896540
transform 1 0 5385 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_27
timestamp 1704896540
transform 1 0 5385 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_28
timestamp 1704896540
transform 1 0 5385 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_29
timestamp 1704896540
transform 1 0 5317 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_30
timestamp 1704896540
transform 1 0 5317 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_31
timestamp 1704896540
transform 1 0 5317 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_32
timestamp 1704896540
transform 1 0 4831 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_33
timestamp 1704896540
transform 1 0 4831 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_34
timestamp 1704896540
transform 1 0 4831 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_35
timestamp 1704896540
transform 1 0 4763 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_36
timestamp 1704896540
transform 1 0 4763 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_37
timestamp 1704896540
transform 1 0 4763 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_38
timestamp 1704896540
transform 1 0 4277 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_39
timestamp 1704896540
transform 1 0 4277 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_40
timestamp 1704896540
transform 1 0 4277 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_41
timestamp 1704896540
transform 1 0 4209 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_42
timestamp 1704896540
transform 1 0 4209 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_43
timestamp 1704896540
transform 1 0 4209 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_44
timestamp 1704896540
transform 1 0 3723 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_45
timestamp 1704896540
transform 1 0 3723 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_46
timestamp 1704896540
transform 1 0 3723 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_47
timestamp 1704896540
transform 1 0 3655 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_48
timestamp 1704896540
transform 1 0 3655 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_49
timestamp 1704896540
transform 1 0 3655 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_50
timestamp 1704896540
transform 1 0 3169 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_51
timestamp 1704896540
transform 1 0 3169 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_52
timestamp 1704896540
transform 1 0 3169 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_53
timestamp 1704896540
transform 1 0 3101 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_54
timestamp 1704896540
transform 1 0 3101 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_55
timestamp 1704896540
transform 1 0 3101 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_56
timestamp 1704896540
transform 1 0 5317 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_57
timestamp 1704896540
transform 1 0 5317 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_58
timestamp 1704896540
transform 1 0 5317 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_59
timestamp 1704896540
transform 1 0 5317 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_60
timestamp 1704896540
transform 1 0 5317 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_61
timestamp 1704896540
transform 1 0 5385 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_62
timestamp 1704896540
transform 1 0 5385 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_63
timestamp 1704896540
transform 1 0 5385 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_64
timestamp 1704896540
transform 1 0 5385 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_65
timestamp 1704896540
transform 1 0 5385 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_66
timestamp 1704896540
transform 1 0 5871 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_67
timestamp 1704896540
transform 1 0 5871 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_68
timestamp 1704896540
transform 1 0 5871 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_69
timestamp 1704896540
transform 1 0 5871 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_70
timestamp 1704896540
transform 1 0 5871 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_71
timestamp 1704896540
transform 1 0 5939 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_72
timestamp 1704896540
transform 1 0 5939 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_73
timestamp 1704896540
transform 1 0 5939 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_74
timestamp 1704896540
transform 1 0 5939 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_75
timestamp 1704896540
transform 1 0 5939 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_76
timestamp 1704896540
transform 1 0 6425 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_77
timestamp 1704896540
transform 1 0 6425 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_78
timestamp 1704896540
transform 1 0 6425 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_79
timestamp 1704896540
transform 1 0 6425 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_80
timestamp 1704896540
transform 1 0 6425 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_81
timestamp 1704896540
transform 1 0 6493 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_82
timestamp 1704896540
transform 1 0 6493 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_83
timestamp 1704896540
transform 1 0 6493 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_84
timestamp 1704896540
transform 1 0 6493 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_85
timestamp 1704896540
transform 1 0 6493 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_86
timestamp 1704896540
transform 1 0 5317 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_87
timestamp 1704896540
transform 1 0 6493 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_88
timestamp 1704896540
transform 1 0 6425 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_89
timestamp 1704896540
transform 1 0 5939 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_90
timestamp 1704896540
transform 1 0 5871 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_91
timestamp 1704896540
transform 1 0 6493 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_92
timestamp 1704896540
transform 1 0 5939 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_93
timestamp 1704896540
transform 1 0 6425 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_94
timestamp 1704896540
transform 1 0 5871 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_95
timestamp 1704896540
transform 1 0 5385 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_96
timestamp 1704896540
transform 1 0 5317 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_97
timestamp 1704896540
transform 1 0 4831 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_98
timestamp 1704896540
transform 1 0 4763 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_99
timestamp 1704896540
transform 1 0 4277 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_100
timestamp 1704896540
transform 1 0 4209 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_101
timestamp 1704896540
transform 1 0 3723 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_102
timestamp 1704896540
transform 1 0 3655 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_103
timestamp 1704896540
transform 1 0 3169 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_104
timestamp 1704896540
transform 1 0 3101 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_105
timestamp 1704896540
transform 1 0 6425 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_106
timestamp 1704896540
transform 1 0 4209 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_107
timestamp 1704896540
transform 1 0 6979 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_108
timestamp 1704896540
transform 1 0 7047 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_109
timestamp 1704896540
transform 1 0 6979 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_110
timestamp 1704896540
transform 1 0 6979 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_111
timestamp 1704896540
transform 1 0 7047 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_112
timestamp 1704896540
transform 1 0 7047 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_113
timestamp 1704896540
transform 1 0 6979 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_114
timestamp 1704896540
transform 1 0 6979 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_115
timestamp 1704896540
transform 1 0 6979 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_116
timestamp 1704896540
transform 1 0 6979 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_117
timestamp 1704896540
transform 1 0 6979 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_118
timestamp 1704896540
transform 1 0 6979 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_119
timestamp 1704896540
transform 1 0 7047 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_120
timestamp 1704896540
transform 1 0 7047 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_121
timestamp 1704896540
transform 1 0 7047 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_122
timestamp 1704896540
transform 1 0 7047 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_123
timestamp 1704896540
transform 1 0 7047 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_124
timestamp 1704896540
transform 1 0 7047 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_125
timestamp 1704896540
transform 1 0 6979 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_126
timestamp 1704896540
transform 1 0 6979 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_127
timestamp 1704896540
transform 1 0 6979 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_128
timestamp 1704896540
transform 1 0 6979 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_129
timestamp 1704896540
transform 1 0 6979 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_130
timestamp 1704896540
transform 1 0 7047 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_131
timestamp 1704896540
transform 1 0 7047 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_132
timestamp 1704896540
transform 1 0 7047 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_133
timestamp 1704896540
transform 1 0 7047 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_134
timestamp 1704896540
transform 1 0 7047 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_135
timestamp 1704896540
transform 1 0 5385 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_136
timestamp 1704896540
transform 1 0 7601 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_137
timestamp 1704896540
transform 1 0 7533 0 -1 11454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_138
timestamp 1704896540
transform 1 0 7601 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_139
timestamp 1704896540
transform 1 0 7533 0 -1 13454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_140
timestamp 1704896540
transform 1 0 7601 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_141
timestamp 1704896540
transform 1 0 7533 0 -1 15454
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_142
timestamp 1704896540
transform 1 0 7601 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_143
timestamp 1704896540
transform 1 0 7533 0 -1 18722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_144
timestamp 1704896540
transform 1 0 7601 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_145
timestamp 1704896540
transform 1 0 7533 0 -1 20722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_146
timestamp 1704896540
transform 1 0 7601 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_147
timestamp 1704896540
transform 1 0 7601 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_148
timestamp 1704896540
transform 1 0 7601 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_149
timestamp 1704896540
transform 1 0 7601 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_150
timestamp 1704896540
transform 1 0 7601 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_151
timestamp 1704896540
transform 1 0 7533 0 -1 22722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_152
timestamp 1704896540
transform 1 0 7533 0 -1 24722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_153
timestamp 1704896540
transform 1 0 7533 0 -1 26722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_154
timestamp 1704896540
transform 1 0 7533 0 -1 28722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_155
timestamp 1704896540
transform 1 0 7533 0 -1 30722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_156
timestamp 1704896540
transform 1 0 7601 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_157
timestamp 1704896540
transform 1 0 7601 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_158
timestamp 1704896540
transform 1 0 7601 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_159
timestamp 1704896540
transform 1 0 7601 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_160
timestamp 1704896540
transform 1 0 7533 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_161
timestamp 1704896540
transform 1 0 7533 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_162
timestamp 1704896540
transform 1 0 7533 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_163
timestamp 1704896540
transform 1 0 7533 0 -1 38722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_164
timestamp 1704896540
transform 1 0 4831 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_165
timestamp 1704896540
transform 1 0 3101 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_166
timestamp 1704896540
transform 1 0 3101 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_167
timestamp 1704896540
transform 1 0 3101 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_168
timestamp 1704896540
transform 1 0 3169 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_169
timestamp 1704896540
transform 1 0 3169 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_170
timestamp 1704896540
transform 1 0 3169 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_171
timestamp 1704896540
transform 1 0 3655 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_172
timestamp 1704896540
transform 1 0 3655 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_173
timestamp 1704896540
transform 1 0 3655 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_174
timestamp 1704896540
transform 1 0 3723 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_175
timestamp 1704896540
transform 1 0 3723 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_176
timestamp 1704896540
transform 1 0 3723 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_177
timestamp 1704896540
transform 1 0 4209 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_178
timestamp 1704896540
transform 1 0 4209 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_179
timestamp 1704896540
transform 1 0 4277 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_180
timestamp 1704896540
transform 1 0 4277 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_181
timestamp 1704896540
transform 1 0 4277 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_182
timestamp 1704896540
transform 1 0 4763 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_183
timestamp 1704896540
transform 1 0 4763 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_184
timestamp 1704896540
transform 1 0 4763 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_185
timestamp 1704896540
transform 1 0 4831 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_186
timestamp 1704896540
transform 1 0 4831 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_187
timestamp 1704896540
transform 1 0 5317 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_188
timestamp 1704896540
transform 1 0 5317 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_189
timestamp 1704896540
transform 1 0 5317 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_190
timestamp 1704896540
transform 1 0 5385 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_191
timestamp 1704896540
transform 1 0 5385 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_192
timestamp 1704896540
transform 1 0 5385 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_193
timestamp 1704896540
transform 1 0 5871 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_194
timestamp 1704896540
transform 1 0 5871 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_195
timestamp 1704896540
transform 1 0 5871 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_196
timestamp 1704896540
transform 1 0 6425 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_197
timestamp 1704896540
transform 1 0 6425 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_198
timestamp 1704896540
transform 1 0 5939 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_199
timestamp 1704896540
transform 1 0 5939 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_200
timestamp 1704896540
transform 1 0 5939 0 -1 36722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_201
timestamp 1704896540
transform 1 0 6493 0 -1 32722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_202
timestamp 1704896540
transform 1 0 6493 0 -1 34722
box -26 -26 76 1376
use DFL1_CDNS_55959141808682  DFL1_CDNS_55959141808682_203
timestamp 1704896540
transform 1 0 6493 0 -1 36722
box -26 -26 76 1376
use nfet_CDNS_55959141808707  nfet_CDNS_55959141808707_0
timestamp 1704896540
transform 1 0 5239 0 1 25372
box -266 -32 2756 1432
use nfet_CDNS_55959141808707  nfet_CDNS_55959141808707_1
timestamp 1704896540
transform 1 0 5239 0 1 23372
box -266 -32 2756 1432
use nfet_CDNS_55959141808707  nfet_CDNS_55959141808707_2
timestamp 1704896540
transform 1 0 5239 0 1 21372
box -266 -32 2756 1432
use nfet_CDNS_55959141808707  nfet_CDNS_55959141808707_3
timestamp 1704896540
transform 1 0 5239 0 1 19372
box -266 -32 2756 1432
use nfet_CDNS_55959141808707  nfet_CDNS_55959141808707_4
timestamp 1704896540
transform 1 0 5239 0 1 17372
box -266 -32 2756 1432
use nfet_CDNS_55959141808707  nfet_CDNS_55959141808707_5
timestamp 1704896540
transform 1 0 5239 0 1 27372
box -266 -32 2756 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_0
timestamp 1704896540
transform 1 0 3023 0 1 29372
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_1
timestamp 1704896540
transform 1 0 3023 0 1 14104
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_2
timestamp 1704896540
transform 1 0 3023 0 1 12104
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_3
timestamp 1704896540
transform 1 0 3023 0 1 10104
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_4
timestamp 1704896540
transform 1 0 3023 0 1 31372
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_5
timestamp 1704896540
transform 1 0 3023 0 1 33372
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_6
timestamp 1704896540
transform 1 0 3023 0 1 35372
box -266 -32 4972 1432
use nfet_CDNS_55959141808708  nfet_CDNS_55959141808708_7
timestamp 1704896540
transform 1 0 3023 0 1 37372
box -266 -32 4972 1432
use nfet_CDNS_55959141808709  nfet_CDNS_55959141808709_0
timestamp 1704896540
transform 1 0 2824 0 1 4163
box -79 -32 4303 1432
use nfet_CDNS_55959141808710  nfet_CDNS_55959141808710_0
timestamp 1704896540
transform 1 0 2468 0 1 6058
box -79 -32 4991 1432
use nfet_CDNS_55959141808710  nfet_CDNS_55959141808710_1
timestamp 1704896540
transform 1 0 2468 0 1 7858
box -79 -32 4991 1432
use nfet_CDNS_55959141808711  nfet_CDNS_55959141808711_0
timestamp 1704896540
transform 1 0 2640 0 1 4163
box -82 -32 210 1432
use pfet_CDNS_55959141808687  pfet_CDNS_55959141808687_0
timestamp 1704896540
transform 0 1 3531 1 0 1008
box -92 -36 956 1436
use pfet_CDNS_55959141808687  pfet_CDNS_55959141808687_1
timestamp 1704896540
transform 0 1 2001 1 0 1008
box -92 -36 956 1436
use PYbentRes_CDNS_55959141808706  PYbentRes_CDNS_55959141808706_0
timestamp 1704896540
transform 0 -1 220 1 0 294
box -50 -1458 38933 66
<< labels >>
flabel comment s 8266 38990 8266 38990 0 FreeSans 600 90 0 0 condiode
flabel comment s 7370 3694 7370 3694 0 FreeSans 600 180 0 0 condiode
flabel metal1 s 7727 0 7877 350 2 FreeSans 1000 90 0 0 ogc_lvc
port 2 nsew power bidirectional
flabel metal3 s 2727 0 5308 925 0 FreeSans 96 0 0 0 drn_lvc
port 3 nsew power bidirectional
flabel metal3 s 5608 0 8218 925 0 FreeSans 96 0 0 0 src_bdy_lvc
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 9579 39600
string GDS_END 6061972
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2770452
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
