magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 372 226
<< mvnmos >>
rect 0 0 120 200
rect 176 0 296 200
<< mvndiff >>
rect -50 0 0 200
rect 296 0 346 200
<< poly >>
rect 0 200 120 226
rect 0 -26 120 0
rect 176 200 296 226
rect 176 -26 296 0
<< metal1 >>
rect -51 -16 -5 186
rect 125 -16 171 186
rect 301 -16 347 186
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_0
timestamp 1704896540
transform 1 0 120 0 1 0
box -26 -26 82 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1704896540
transform 1 0 296 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 148 85 148 85 0 FreeSans 300 0 0 0 D
flabel comment s 324 85 324 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86863750
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86862360
<< end >>
