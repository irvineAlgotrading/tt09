magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -79 -26 535 226
<< mvnmos >>
rect 0 0 200 200
rect 256 0 456 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 200 182 256 200
rect 200 148 211 182
rect 245 148 256 182
rect 200 114 256 148
rect 200 80 211 114
rect 245 80 256 114
rect 200 46 256 80
rect 200 12 211 46
rect 245 12 256 46
rect 200 0 256 12
rect 456 182 509 200
rect 456 148 467 182
rect 501 148 509 182
rect 456 114 509 148
rect 456 80 467 114
rect 501 80 509 114
rect 456 46 509 80
rect 456 12 467 46
rect 501 12 509 46
rect 456 0 509 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 211 148 245 182
rect 211 80 245 114
rect 211 12 245 46
rect 467 148 501 182
rect 467 80 501 114
rect 467 12 501 46
<< poly >>
rect 0 200 200 226
rect 256 200 456 226
rect 0 -26 200 0
rect 256 -26 456 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 211 182 245 198
rect 211 114 245 148
rect 211 46 245 80
rect 211 -4 245 12
rect 467 182 501 198
rect 467 114 501 148
rect 467 46 501 80
rect 467 -4 501 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1704896540
transform 1 0 200 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_1
timestamp 1704896540
transform 1 0 456 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 228 97 228 97 0 FreeSans 300 0 0 0 D
flabel comment s 484 97 484 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 87889456
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87888066
<< end >>
