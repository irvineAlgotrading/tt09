magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 67 0 100
rect -50 33 -34 67
rect -50 0 0 33
rect 2040 67 2090 100
rect 2074 33 2090 67
rect 2040 0 2090 33
<< polycont >>
rect -34 33 0 67
rect 2040 33 2074 67
<< npolyres >>
rect 0 0 2040 100
<< locali >>
rect -34 67 0 83
rect -34 17 0 33
rect 2040 67 2074 83
rect 2040 17 2074 33
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform 1 0 2024 0 1 17
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform 1 0 -50 0 1 17
box 0 0 1 1
<< properties >>
string GDS_END 91719880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91719400
<< end >>
