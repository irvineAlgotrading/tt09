magic
tech sky130B
timestamp 1704896540
<< viali >>
rect 0 0 125 89
<< metal1 >>
rect -6 89 131 92
rect -6 0 0 89
rect 125 0 131 89
rect -6 -3 131 0
<< properties >>
string GDS_END 87590034
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87589134
<< end >>
