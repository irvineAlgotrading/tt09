magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 0 0 832 38350
<< ndiff >>
rect 26 102 39 136
rect 73 102 86 136
rect 26 68 86 102
rect 26 34 39 68
rect 73 34 86 68
rect 26 26 86 34
rect 746 38314 806 38324
rect 746 38280 759 38314
rect 793 38280 806 38314
rect 746 38246 806 38280
rect 746 38212 759 38246
rect 793 38212 806 38246
<< ndiffc >>
rect 39 102 73 136
rect 39 34 73 68
rect 759 38280 793 38314
rect 759 38212 793 38246
<< ndiffres >>
rect 26 38264 206 38324
rect 26 136 86 38264
rect 146 86 206 38264
rect 266 38264 446 38324
rect 266 86 326 38264
rect 146 26 326 86
rect 386 86 446 38264
rect 506 38264 686 38324
rect 506 86 566 38264
rect 386 26 566 86
rect 626 86 686 38264
rect 746 86 806 38212
rect 626 26 806 86
<< locali >>
rect 743 38314 809 38316
rect 743 38280 759 38314
rect 793 38280 809 38314
rect 743 38246 809 38280
rect 743 38212 759 38246
rect 793 38212 809 38246
rect 23 102 39 136
rect 73 102 89 136
rect 23 68 89 102
rect 23 34 39 68
rect 73 34 89 68
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform 0 -1 805 1 0 38204
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 0 -1 805 1 0 38272
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1704896540
transform 0 -1 85 1 0 26
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1704896540
transform 0 -1 85 1 0 94
box 0 0 1 1
<< properties >>
string GDS_END 6673440
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6670996
<< end >>
