magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< obsli1 >>
rect 34 3292 2158 3358
rect 34 100 100 3292
rect 260 3066 1932 3132
rect 260 326 326 3066
rect 662 2664 1530 2730
rect 662 728 728 2664
rect 893 893 1299 2499
rect 1464 728 1530 2664
rect 662 662 1530 728
rect 1866 326 1932 3066
rect 260 260 1932 326
rect 2092 100 2158 3292
rect 34 34 2158 100
<< obsm1 >>
rect 38 3296 2154 3354
rect 38 96 96 3296
rect 264 3070 1928 3128
rect 264 322 322 3070
rect 666 2668 1526 2726
rect 666 724 724 2668
rect 923 911 1269 2481
rect 1468 724 1526 2668
rect 666 666 1526 724
rect 1870 322 1928 3070
rect 264 264 1928 322
rect 2096 96 2154 3296
rect 38 38 2154 96
<< properties >>
string FIXED_BBOX 26 26 2166 3366
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9008578
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8938614
<< end >>
