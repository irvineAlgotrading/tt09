magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_0
timestamp 1704896540
transform 1 0 641 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_1
timestamp 1704896540
transform 1 0 1633 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_2
timestamp 1704896540
transform 1 0 2625 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_3
timestamp 1704896540
transform 1 0 3617 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_4
timestamp 1704896540
transform 1 0 4609 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_5
timestamp 1704896540
transform 1 0 5601 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_6
timestamp 1704896540
transform 1 0 6593 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_7
timestamp 1704896540
transform 1 0 7585 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_8
timestamp 1704896540
transform 1 0 8577 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_9
timestamp 1704896540
transform 1 0 9569 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_10
timestamp 1704896540
transform 1 0 10561 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_11
timestamp 1704896540
transform 1 0 11553 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 17338386
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 17325410
<< end >>
