magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -603 3571 2375 5914
<< pwell >>
rect 2727 43 2813 1121
<< mvpsubdiff >>
rect 2753 1071 2787 1095
rect 2753 999 2787 1037
rect 2753 927 2787 965
rect 2753 855 2787 893
rect 2753 783 2787 821
rect 2753 711 2787 749
rect 2753 638 2787 677
rect 2753 565 2787 604
rect 2753 492 2787 531
rect 2753 419 2787 458
rect 2753 346 2787 385
rect 2753 273 2787 312
rect 2753 200 2787 239
rect 2753 127 2787 166
rect 2753 69 2787 93
<< mvnsubdiff >>
rect -537 5814 2309 5848
rect -537 5780 -503 5814
rect -469 5780 -435 5814
rect -401 5780 -367 5814
rect -333 5780 -263 5814
rect -229 5780 -194 5814
rect -160 5780 -125 5814
rect -91 5780 -56 5814
rect -22 5780 13 5814
rect 47 5780 82 5814
rect 116 5780 151 5814
rect 185 5780 220 5814
rect 254 5780 289 5814
rect 323 5780 358 5814
rect 392 5780 427 5814
rect 461 5780 496 5814
rect 530 5780 565 5814
rect 599 5780 634 5814
rect 668 5780 703 5814
rect 737 5780 772 5814
rect 806 5780 841 5814
rect 875 5780 910 5814
rect 944 5780 979 5814
rect 1013 5780 1048 5814
rect 1082 5780 1117 5814
rect 1151 5780 1186 5814
rect 1220 5780 1255 5814
rect 1289 5780 1324 5814
rect 1358 5780 1393 5814
rect 1427 5780 1462 5814
rect 1496 5780 1531 5814
rect 1565 5780 1600 5814
rect 1634 5780 1669 5814
rect 1703 5780 1738 5814
rect 1772 5780 1807 5814
rect -537 5746 1807 5780
rect -537 5744 -263 5746
rect -537 5710 -503 5744
rect -469 5710 -435 5744
rect -401 5710 -367 5744
rect -333 5712 -263 5744
rect -229 5712 -194 5746
rect -160 5712 -125 5746
rect -91 5712 -56 5746
rect -22 5712 13 5746
rect 47 5712 82 5746
rect 116 5712 151 5746
rect 185 5712 220 5746
rect 254 5712 289 5746
rect 323 5712 358 5746
rect 392 5712 427 5746
rect 461 5712 496 5746
rect 530 5712 565 5746
rect 599 5712 634 5746
rect 668 5712 703 5746
rect 737 5712 772 5746
rect 806 5712 841 5746
rect 875 5712 910 5746
rect 944 5712 979 5746
rect 1013 5712 1048 5746
rect 1082 5712 1117 5746
rect 1151 5712 1186 5746
rect 1220 5712 1255 5746
rect 1289 5712 1324 5746
rect 1358 5712 1393 5746
rect 1427 5712 1462 5746
rect 1496 5712 1531 5746
rect 1565 5712 1600 5746
rect 1634 5712 1669 5746
rect 1703 5712 1738 5746
rect 1772 5712 1807 5746
rect -333 5710 1807 5712
rect -537 5678 1807 5710
rect -537 5674 -263 5678
rect -537 5640 -503 5674
rect -469 5640 -435 5674
rect -401 5640 -367 5674
rect -333 5644 -263 5674
rect -229 5644 -194 5678
rect -160 5644 -125 5678
rect -91 5644 -56 5678
rect -22 5644 13 5678
rect 47 5644 82 5678
rect 116 5644 151 5678
rect 185 5644 220 5678
rect 254 5644 289 5678
rect 323 5644 358 5678
rect 392 5644 427 5678
rect 461 5644 496 5678
rect 530 5644 565 5678
rect 599 5644 634 5678
rect 668 5644 703 5678
rect 737 5644 772 5678
rect 806 5644 841 5678
rect 875 5644 910 5678
rect 944 5644 979 5678
rect 1013 5644 1048 5678
rect 1082 5644 1117 5678
rect 1151 5644 1186 5678
rect 1220 5644 1255 5678
rect 1289 5644 1324 5678
rect 1358 5644 1393 5678
rect 1427 5644 1462 5678
rect 1496 5644 1531 5678
rect 1565 5644 1600 5678
rect 1634 5644 1669 5678
rect 1703 5644 1738 5678
rect 1772 5644 1807 5678
rect 1977 5802 2309 5814
rect 1977 5768 2037 5802
rect 2071 5768 2105 5802
rect 2139 5768 2173 5802
rect 2207 5768 2241 5802
rect 2275 5768 2309 5802
rect 1977 5731 2309 5768
rect 1977 5697 2037 5731
rect 2071 5697 2105 5731
rect 2139 5697 2173 5731
rect 2207 5697 2241 5731
rect 2275 5697 2309 5731
rect 1977 5660 2309 5697
rect 1977 5644 2037 5660
rect -333 5640 2037 5644
rect -537 5626 2037 5640
rect 2071 5626 2105 5660
rect 2139 5626 2173 5660
rect 2207 5626 2241 5660
rect 2275 5626 2309 5660
rect -537 5610 2309 5626
rect -537 5609 -294 5610
rect -537 5604 -299 5609
rect -537 5570 -503 5604
rect -469 5570 -435 5604
rect -401 5570 -367 5604
rect -333 5570 -299 5604
rect -537 5534 -299 5570
rect -537 5500 -503 5534
rect -469 5500 -435 5534
rect -401 5500 -367 5534
rect -333 5500 -299 5534
rect 2003 5589 2309 5610
rect 2003 5555 2037 5589
rect 2071 5555 2105 5589
rect 2139 5555 2173 5589
rect 2207 5555 2241 5589
rect 2275 5555 2309 5589
rect -537 5464 -299 5500
rect 2003 5518 2309 5555
rect 2003 5484 2037 5518
rect 2071 5484 2105 5518
rect 2139 5484 2173 5518
rect 2207 5484 2241 5518
rect 2275 5484 2309 5518
rect -537 5430 -503 5464
rect -469 5430 -435 5464
rect -401 5430 -367 5464
rect -333 5430 -299 5464
rect -537 5394 -299 5430
rect -537 5360 -503 5394
rect -469 5360 -435 5394
rect -401 5360 -367 5394
rect -333 5360 -299 5394
rect -537 5324 -299 5360
rect -537 5290 -503 5324
rect -469 5290 -435 5324
rect -401 5290 -367 5324
rect -333 5290 -299 5324
rect -537 5254 -299 5290
rect -537 5220 -503 5254
rect -469 5220 -435 5254
rect -401 5220 -367 5254
rect -333 5220 -299 5254
rect -537 5184 -299 5220
rect -537 5150 -503 5184
rect -469 5150 -435 5184
rect -401 5150 -367 5184
rect -333 5150 -299 5184
rect -537 5114 -299 5150
rect -537 5080 -503 5114
rect -469 5080 -435 5114
rect -401 5080 -367 5114
rect -333 5080 -299 5114
rect -537 5044 -299 5080
rect -537 5010 -503 5044
rect -469 5010 -435 5044
rect -401 5010 -367 5044
rect -333 5010 -299 5044
rect -537 4974 -299 5010
rect -537 4940 -503 4974
rect -469 4940 -435 4974
rect -401 4940 -367 4974
rect -333 4940 -299 4974
rect -537 4904 -299 4940
rect -537 4870 -503 4904
rect -469 4870 -435 4904
rect -401 4870 -367 4904
rect -333 4870 -299 4904
rect -537 4834 -299 4870
rect -537 4800 -503 4834
rect -469 4800 -435 4834
rect -401 4800 -367 4834
rect -333 4800 -299 4834
rect -537 4764 -299 4800
rect -537 4730 -503 4764
rect -469 4730 -435 4764
rect -401 4730 -367 4764
rect -333 4760 -299 4764
rect 2003 5446 2309 5484
rect 2003 5412 2037 5446
rect 2071 5412 2105 5446
rect 2139 5412 2173 5446
rect 2207 5412 2241 5446
rect 2275 5412 2309 5446
rect 2003 5374 2309 5412
rect 2003 5340 2037 5374
rect 2071 5340 2105 5374
rect 2139 5340 2173 5374
rect 2207 5340 2241 5374
rect 2275 5340 2309 5374
rect 2003 5302 2309 5340
rect 2003 5268 2037 5302
rect 2071 5268 2105 5302
rect 2139 5268 2173 5302
rect 2207 5268 2241 5302
rect 2275 5268 2309 5302
rect 2003 5230 2309 5268
rect 2003 5196 2037 5230
rect 2071 5196 2105 5230
rect 2139 5196 2173 5230
rect 2207 5196 2241 5230
rect 2275 5196 2309 5230
rect 2003 5158 2309 5196
rect 2003 5124 2037 5158
rect 2071 5124 2105 5158
rect 2139 5124 2173 5158
rect 2207 5124 2241 5158
rect 2275 5124 2309 5158
rect 2003 5086 2309 5124
rect 2003 5052 2037 5086
rect 2071 5052 2105 5086
rect 2139 5052 2173 5086
rect 2207 5052 2241 5086
rect 2275 5052 2309 5086
rect 2003 5014 2309 5052
rect 2003 4980 2037 5014
rect 2071 4980 2105 5014
rect 2139 4980 2173 5014
rect 2207 4980 2241 5014
rect 2275 4980 2309 5014
rect 2003 4942 2309 4980
rect 2003 4908 2037 4942
rect 2071 4908 2105 4942
rect 2139 4908 2173 4942
rect 2207 4908 2241 4942
rect 2275 4908 2309 4942
rect 2003 4870 2309 4908
rect 2003 4836 2037 4870
rect 2071 4836 2105 4870
rect 2139 4836 2173 4870
rect 2207 4836 2241 4870
rect 2275 4836 2309 4870
rect 2003 4798 2309 4836
rect 2003 4764 2037 4798
rect 2071 4764 2105 4798
rect 2139 4764 2173 4798
rect 2207 4764 2241 4798
rect 2275 4764 2309 4798
rect 2003 4760 2309 4764
rect -333 4730 2309 4760
rect -537 4726 2309 4730
rect -537 4694 -265 4726
rect -537 4660 -503 4694
rect -469 4660 -435 4694
rect -401 4660 -367 4694
rect -333 4692 -265 4694
rect -231 4692 -196 4726
rect -162 4692 -127 4726
rect -93 4692 -58 4726
rect -24 4692 11 4726
rect 45 4692 80 4726
rect 114 4692 149 4726
rect 183 4692 218 4726
rect 252 4692 287 4726
rect 321 4692 356 4726
rect 390 4692 425 4726
rect 459 4692 494 4726
rect 528 4692 563 4726
rect 597 4692 632 4726
rect 666 4692 701 4726
rect 735 4692 770 4726
rect 804 4692 839 4726
rect 873 4692 908 4726
rect 942 4692 977 4726
rect 1011 4692 1046 4726
rect 1080 4692 1115 4726
rect 1149 4692 1184 4726
rect 1218 4692 1254 4726
rect 1288 4692 1324 4726
rect 1358 4692 1394 4726
rect 1428 4692 1464 4726
rect 1498 4692 1534 4726
rect 1568 4692 1604 4726
rect 1638 4692 1674 4726
rect 1708 4692 1744 4726
rect 1778 4692 1814 4726
rect 1848 4692 1884 4726
rect 1918 4692 1954 4726
rect 1988 4692 2037 4726
rect 2071 4692 2105 4726
rect 2139 4692 2173 4726
rect 2207 4692 2241 4726
rect 2275 4692 2309 4726
rect -333 4660 2309 4692
rect -537 4658 2309 4660
rect -537 4624 -299 4658
rect -537 4590 -503 4624
rect -469 4590 -435 4624
rect -401 4590 -367 4624
rect -333 4590 -299 4624
rect -537 4554 -299 4590
rect -537 4520 -503 4554
rect -469 4520 -435 4554
rect -401 4520 -367 4554
rect -333 4520 -299 4554
rect -537 4484 -299 4520
rect -537 4450 -503 4484
rect -469 4450 -435 4484
rect -401 4450 -367 4484
rect -333 4450 -299 4484
rect -537 4413 -299 4450
rect -537 4379 -503 4413
rect -469 4379 -435 4413
rect -401 4379 -367 4413
rect -333 4379 -299 4413
rect -537 4342 -299 4379
rect 740 4640 842 4658
rect 740 4606 774 4640
rect 808 4606 842 4640
rect 740 4568 842 4606
rect 740 4534 774 4568
rect 808 4534 842 4568
rect 1799 4624 2309 4658
rect 1799 4590 1833 4624
rect 1867 4590 1901 4624
rect 1935 4590 1969 4624
rect 2003 4590 2037 4624
rect 2071 4590 2105 4624
rect 2139 4590 2173 4624
rect 2207 4590 2241 4624
rect 2275 4590 2309 4624
rect 740 4496 842 4534
rect 1799 4554 2309 4590
rect 1799 4520 1833 4554
rect 1867 4520 1901 4554
rect 1935 4520 1969 4554
rect 2003 4520 2037 4554
rect 2071 4520 2105 4554
rect 2139 4520 2173 4554
rect 2207 4520 2241 4554
rect 2275 4520 2309 4554
rect 740 4462 774 4496
rect 808 4462 842 4496
rect 740 4424 842 4462
rect 740 4390 774 4424
rect 808 4390 842 4424
rect -537 4308 -503 4342
rect -469 4308 -435 4342
rect -401 4308 -367 4342
rect -333 4308 -299 4342
rect 740 4352 842 4390
rect 740 4318 774 4352
rect 808 4318 842 4352
rect -537 4271 -299 4308
rect -537 4237 -503 4271
rect -469 4237 -435 4271
rect -401 4237 -367 4271
rect -333 4237 -299 4271
rect -537 4200 -299 4237
rect 740 4280 842 4318
rect 740 4246 774 4280
rect 808 4246 842 4280
rect 740 4208 842 4246
rect -537 4166 -503 4200
rect -469 4166 -435 4200
rect -401 4166 -367 4200
rect -333 4166 -299 4200
rect -537 4129 -299 4166
rect 740 4174 774 4208
rect 808 4174 842 4208
rect 740 4136 842 4174
rect -537 4095 -503 4129
rect -469 4095 -435 4129
rect -401 4095 -367 4129
rect -333 4095 -299 4129
rect -537 4058 -299 4095
rect -537 4024 -503 4058
rect -469 4024 -435 4058
rect -401 4024 -367 4058
rect -333 4024 -299 4058
rect -537 3987 -299 4024
rect -537 3953 -503 3987
rect -469 3953 -435 3987
rect -401 3953 -367 3987
rect -333 3953 -299 3987
rect -537 3916 -299 3953
rect -537 3882 -503 3916
rect -469 3882 -435 3916
rect -401 3882 -367 3916
rect -333 3882 -299 3916
rect -537 3845 -299 3882
rect -537 3811 -503 3845
rect -469 3811 -435 3845
rect -401 3811 -367 3845
rect -333 3811 -299 3845
rect -537 3807 -299 3811
rect 740 4102 774 4136
rect 808 4102 842 4136
rect 740 4064 842 4102
rect 740 4030 774 4064
rect 808 4030 842 4064
rect 740 3991 842 4030
rect 740 3957 774 3991
rect 808 3957 842 3991
rect 740 3918 842 3957
rect 740 3884 774 3918
rect 808 3884 842 3918
rect 740 3845 842 3884
rect 740 3811 774 3845
rect 808 3811 842 3845
rect 740 3807 842 3811
rect 1799 4484 2309 4520
rect 1799 4450 1833 4484
rect 1867 4450 1901 4484
rect 1935 4450 1969 4484
rect 2003 4450 2037 4484
rect 2071 4450 2105 4484
rect 2139 4450 2173 4484
rect 2207 4450 2241 4484
rect 2275 4450 2309 4484
rect 1799 4413 2309 4450
rect 1799 4379 1833 4413
rect 1867 4379 1901 4413
rect 1935 4379 1969 4413
rect 2003 4379 2037 4413
rect 2071 4379 2105 4413
rect 2139 4379 2173 4413
rect 2207 4379 2241 4413
rect 2275 4379 2309 4413
rect 1799 4342 2309 4379
rect 1799 4308 1833 4342
rect 1867 4308 1901 4342
rect 1935 4308 1969 4342
rect 2003 4308 2037 4342
rect 2071 4308 2105 4342
rect 2139 4308 2173 4342
rect 2207 4308 2241 4342
rect 2275 4308 2309 4342
rect 1799 4271 2309 4308
rect 1799 4237 1833 4271
rect 1867 4237 1901 4271
rect 1935 4237 1969 4271
rect 2003 4237 2037 4271
rect 2071 4237 2105 4271
rect 2139 4237 2173 4271
rect 2207 4237 2241 4271
rect 2275 4237 2309 4271
rect 1799 4200 2309 4237
rect 1799 4166 1833 4200
rect 1867 4166 1901 4200
rect 1935 4166 1969 4200
rect 2003 4166 2037 4200
rect 2071 4166 2105 4200
rect 2139 4166 2173 4200
rect 2207 4166 2241 4200
rect 2275 4166 2309 4200
rect 1799 4129 2309 4166
rect 1799 4095 1833 4129
rect 1867 4095 1901 4129
rect 1935 4095 1969 4129
rect 2003 4095 2037 4129
rect 2071 4095 2105 4129
rect 2139 4095 2173 4129
rect 2207 4095 2241 4129
rect 2275 4095 2309 4129
rect 1799 4058 2309 4095
rect 1799 4024 1833 4058
rect 1867 4024 1901 4058
rect 1935 4024 1969 4058
rect 2003 4024 2037 4058
rect 2071 4024 2105 4058
rect 2139 4024 2173 4058
rect 2207 4024 2241 4058
rect 2275 4024 2309 4058
rect 1799 3987 2309 4024
rect 1799 3953 1833 3987
rect 1867 3953 1901 3987
rect 1935 3953 1969 3987
rect 2003 3953 2037 3987
rect 2071 3953 2105 3987
rect 2139 3953 2173 3987
rect 2207 3953 2241 3987
rect 2275 3953 2309 3987
rect 1799 3916 2309 3953
rect 1799 3882 1833 3916
rect 1867 3882 1901 3916
rect 1935 3882 1969 3916
rect 2003 3882 2037 3916
rect 2071 3882 2105 3916
rect 2139 3882 2173 3916
rect 2207 3882 2241 3916
rect 2275 3882 2309 3916
rect 1799 3845 2309 3882
rect 1799 3811 1833 3845
rect 1867 3811 1901 3845
rect 1935 3811 1969 3845
rect 2003 3811 2037 3845
rect 2071 3811 2105 3845
rect 2139 3811 2173 3845
rect 2207 3811 2241 3845
rect 2275 3811 2309 3845
rect 1799 3807 2309 3811
rect -537 3773 2309 3807
rect -537 3671 -503 3773
rect 619 3739 654 3773
rect 688 3739 723 3773
rect 757 3739 792 3773
rect 826 3739 861 3773
rect 895 3739 930 3773
rect 964 3739 999 3773
rect 1033 3739 1068 3773
rect 1102 3739 1137 3773
rect 1171 3739 1206 3773
rect 1240 3739 1275 3773
rect 1309 3739 1344 3773
rect 1378 3739 1413 3773
rect 1447 3739 1482 3773
rect 1516 3739 1551 3773
rect 1585 3739 1620 3773
rect 1654 3739 1689 3773
rect 1723 3739 1758 3773
rect 1792 3739 1827 3773
rect 1861 3739 1896 3773
rect 1930 3739 1965 3773
rect 1999 3739 2034 3773
rect 2068 3739 2103 3773
rect 2137 3739 2172 3773
rect 2206 3739 2241 3773
rect 2275 3739 2309 3773
rect 619 3705 2309 3739
rect 619 3671 654 3705
rect 688 3671 723 3705
rect 757 3671 792 3705
rect 826 3671 861 3705
rect 895 3671 930 3705
rect 964 3671 999 3705
rect 1033 3671 1068 3705
rect 1102 3671 1137 3705
rect 1171 3671 1206 3705
rect 1240 3671 1275 3705
rect 1309 3671 1344 3705
rect 1378 3671 1413 3705
rect 1447 3671 1482 3705
rect 1516 3671 1551 3705
rect 1585 3671 1620 3705
rect 1654 3671 1689 3705
rect 1723 3671 1758 3705
rect 1792 3671 1827 3705
rect 1861 3671 1896 3705
rect 1930 3671 1965 3705
rect 1999 3671 2034 3705
rect 2068 3671 2103 3705
rect 2137 3671 2172 3705
rect 2206 3671 2241 3705
rect 2275 3671 2309 3705
rect -537 3637 2309 3671
<< mvpsubdiffcont >>
rect 2753 1037 2787 1071
rect 2753 965 2787 999
rect 2753 893 2787 927
rect 2753 821 2787 855
rect 2753 749 2787 783
rect 2753 677 2787 711
rect 2753 604 2787 638
rect 2753 531 2787 565
rect 2753 458 2787 492
rect 2753 385 2787 419
rect 2753 312 2787 346
rect 2753 239 2787 273
rect 2753 166 2787 200
rect 2753 93 2787 127
<< mvnsubdiffcont >>
rect -503 5780 -469 5814
rect -435 5780 -401 5814
rect -367 5780 -333 5814
rect -263 5780 -229 5814
rect -194 5780 -160 5814
rect -125 5780 -91 5814
rect -56 5780 -22 5814
rect 13 5780 47 5814
rect 82 5780 116 5814
rect 151 5780 185 5814
rect 220 5780 254 5814
rect 289 5780 323 5814
rect 358 5780 392 5814
rect 427 5780 461 5814
rect 496 5780 530 5814
rect 565 5780 599 5814
rect 634 5780 668 5814
rect 703 5780 737 5814
rect 772 5780 806 5814
rect 841 5780 875 5814
rect 910 5780 944 5814
rect 979 5780 1013 5814
rect 1048 5780 1082 5814
rect 1117 5780 1151 5814
rect 1186 5780 1220 5814
rect 1255 5780 1289 5814
rect 1324 5780 1358 5814
rect 1393 5780 1427 5814
rect 1462 5780 1496 5814
rect 1531 5780 1565 5814
rect 1600 5780 1634 5814
rect 1669 5780 1703 5814
rect 1738 5780 1772 5814
rect -503 5710 -469 5744
rect -435 5710 -401 5744
rect -367 5710 -333 5744
rect -263 5712 -229 5746
rect -194 5712 -160 5746
rect -125 5712 -91 5746
rect -56 5712 -22 5746
rect 13 5712 47 5746
rect 82 5712 116 5746
rect 151 5712 185 5746
rect 220 5712 254 5746
rect 289 5712 323 5746
rect 358 5712 392 5746
rect 427 5712 461 5746
rect 496 5712 530 5746
rect 565 5712 599 5746
rect 634 5712 668 5746
rect 703 5712 737 5746
rect 772 5712 806 5746
rect 841 5712 875 5746
rect 910 5712 944 5746
rect 979 5712 1013 5746
rect 1048 5712 1082 5746
rect 1117 5712 1151 5746
rect 1186 5712 1220 5746
rect 1255 5712 1289 5746
rect 1324 5712 1358 5746
rect 1393 5712 1427 5746
rect 1462 5712 1496 5746
rect 1531 5712 1565 5746
rect 1600 5712 1634 5746
rect 1669 5712 1703 5746
rect 1738 5712 1772 5746
rect -503 5640 -469 5674
rect -435 5640 -401 5674
rect -367 5640 -333 5674
rect -263 5644 -229 5678
rect -194 5644 -160 5678
rect -125 5644 -91 5678
rect -56 5644 -22 5678
rect 13 5644 47 5678
rect 82 5644 116 5678
rect 151 5644 185 5678
rect 220 5644 254 5678
rect 289 5644 323 5678
rect 358 5644 392 5678
rect 427 5644 461 5678
rect 496 5644 530 5678
rect 565 5644 599 5678
rect 634 5644 668 5678
rect 703 5644 737 5678
rect 772 5644 806 5678
rect 841 5644 875 5678
rect 910 5644 944 5678
rect 979 5644 1013 5678
rect 1048 5644 1082 5678
rect 1117 5644 1151 5678
rect 1186 5644 1220 5678
rect 1255 5644 1289 5678
rect 1324 5644 1358 5678
rect 1393 5644 1427 5678
rect 1462 5644 1496 5678
rect 1531 5644 1565 5678
rect 1600 5644 1634 5678
rect 1669 5644 1703 5678
rect 1738 5644 1772 5678
rect 1807 5644 1977 5814
rect 2037 5768 2071 5802
rect 2105 5768 2139 5802
rect 2173 5768 2207 5802
rect 2241 5768 2275 5802
rect 2037 5697 2071 5731
rect 2105 5697 2139 5731
rect 2173 5697 2207 5731
rect 2241 5697 2275 5731
rect 2037 5626 2071 5660
rect 2105 5626 2139 5660
rect 2173 5626 2207 5660
rect 2241 5626 2275 5660
rect -503 5570 -469 5604
rect -435 5570 -401 5604
rect -367 5570 -333 5604
rect -503 5500 -469 5534
rect -435 5500 -401 5534
rect -367 5500 -333 5534
rect 2037 5555 2071 5589
rect 2105 5555 2139 5589
rect 2173 5555 2207 5589
rect 2241 5555 2275 5589
rect 2037 5484 2071 5518
rect 2105 5484 2139 5518
rect 2173 5484 2207 5518
rect 2241 5484 2275 5518
rect -503 5430 -469 5464
rect -435 5430 -401 5464
rect -367 5430 -333 5464
rect -503 5360 -469 5394
rect -435 5360 -401 5394
rect -367 5360 -333 5394
rect -503 5290 -469 5324
rect -435 5290 -401 5324
rect -367 5290 -333 5324
rect -503 5220 -469 5254
rect -435 5220 -401 5254
rect -367 5220 -333 5254
rect -503 5150 -469 5184
rect -435 5150 -401 5184
rect -367 5150 -333 5184
rect -503 5080 -469 5114
rect -435 5080 -401 5114
rect -367 5080 -333 5114
rect -503 5010 -469 5044
rect -435 5010 -401 5044
rect -367 5010 -333 5044
rect -503 4940 -469 4974
rect -435 4940 -401 4974
rect -367 4940 -333 4974
rect -503 4870 -469 4904
rect -435 4870 -401 4904
rect -367 4870 -333 4904
rect -503 4800 -469 4834
rect -435 4800 -401 4834
rect -367 4800 -333 4834
rect -503 4730 -469 4764
rect -435 4730 -401 4764
rect -367 4730 -333 4764
rect 2037 5412 2071 5446
rect 2105 5412 2139 5446
rect 2173 5412 2207 5446
rect 2241 5412 2275 5446
rect 2037 5340 2071 5374
rect 2105 5340 2139 5374
rect 2173 5340 2207 5374
rect 2241 5340 2275 5374
rect 2037 5268 2071 5302
rect 2105 5268 2139 5302
rect 2173 5268 2207 5302
rect 2241 5268 2275 5302
rect 2037 5196 2071 5230
rect 2105 5196 2139 5230
rect 2173 5196 2207 5230
rect 2241 5196 2275 5230
rect 2037 5124 2071 5158
rect 2105 5124 2139 5158
rect 2173 5124 2207 5158
rect 2241 5124 2275 5158
rect 2037 5052 2071 5086
rect 2105 5052 2139 5086
rect 2173 5052 2207 5086
rect 2241 5052 2275 5086
rect 2037 4980 2071 5014
rect 2105 4980 2139 5014
rect 2173 4980 2207 5014
rect 2241 4980 2275 5014
rect 2037 4908 2071 4942
rect 2105 4908 2139 4942
rect 2173 4908 2207 4942
rect 2241 4908 2275 4942
rect 2037 4836 2071 4870
rect 2105 4836 2139 4870
rect 2173 4836 2207 4870
rect 2241 4836 2275 4870
rect 2037 4764 2071 4798
rect 2105 4764 2139 4798
rect 2173 4764 2207 4798
rect 2241 4764 2275 4798
rect -503 4660 -469 4694
rect -435 4660 -401 4694
rect -367 4660 -333 4694
rect -265 4692 -231 4726
rect -196 4692 -162 4726
rect -127 4692 -93 4726
rect -58 4692 -24 4726
rect 11 4692 45 4726
rect 80 4692 114 4726
rect 149 4692 183 4726
rect 218 4692 252 4726
rect 287 4692 321 4726
rect 356 4692 390 4726
rect 425 4692 459 4726
rect 494 4692 528 4726
rect 563 4692 597 4726
rect 632 4692 666 4726
rect 701 4692 735 4726
rect 770 4692 804 4726
rect 839 4692 873 4726
rect 908 4692 942 4726
rect 977 4692 1011 4726
rect 1046 4692 1080 4726
rect 1115 4692 1149 4726
rect 1184 4692 1218 4726
rect 1254 4692 1288 4726
rect 1324 4692 1358 4726
rect 1394 4692 1428 4726
rect 1464 4692 1498 4726
rect 1534 4692 1568 4726
rect 1604 4692 1638 4726
rect 1674 4692 1708 4726
rect 1744 4692 1778 4726
rect 1814 4692 1848 4726
rect 1884 4692 1918 4726
rect 1954 4692 1988 4726
rect 2037 4692 2071 4726
rect 2105 4692 2139 4726
rect 2173 4692 2207 4726
rect 2241 4692 2275 4726
rect -503 4590 -469 4624
rect -435 4590 -401 4624
rect -367 4590 -333 4624
rect -503 4520 -469 4554
rect -435 4520 -401 4554
rect -367 4520 -333 4554
rect -503 4450 -469 4484
rect -435 4450 -401 4484
rect -367 4450 -333 4484
rect -503 4379 -469 4413
rect -435 4379 -401 4413
rect -367 4379 -333 4413
rect 774 4606 808 4640
rect 774 4534 808 4568
rect 1833 4590 1867 4624
rect 1901 4590 1935 4624
rect 1969 4590 2003 4624
rect 2037 4590 2071 4624
rect 2105 4590 2139 4624
rect 2173 4590 2207 4624
rect 2241 4590 2275 4624
rect 1833 4520 1867 4554
rect 1901 4520 1935 4554
rect 1969 4520 2003 4554
rect 2037 4520 2071 4554
rect 2105 4520 2139 4554
rect 2173 4520 2207 4554
rect 2241 4520 2275 4554
rect 774 4462 808 4496
rect 774 4390 808 4424
rect -503 4308 -469 4342
rect -435 4308 -401 4342
rect -367 4308 -333 4342
rect 774 4318 808 4352
rect -503 4237 -469 4271
rect -435 4237 -401 4271
rect -367 4237 -333 4271
rect 774 4246 808 4280
rect -503 4166 -469 4200
rect -435 4166 -401 4200
rect -367 4166 -333 4200
rect 774 4174 808 4208
rect -503 4095 -469 4129
rect -435 4095 -401 4129
rect -367 4095 -333 4129
rect -503 4024 -469 4058
rect -435 4024 -401 4058
rect -367 4024 -333 4058
rect -503 3953 -469 3987
rect -435 3953 -401 3987
rect -367 3953 -333 3987
rect -503 3882 -469 3916
rect -435 3882 -401 3916
rect -367 3882 -333 3916
rect -503 3811 -469 3845
rect -435 3811 -401 3845
rect -367 3811 -333 3845
rect 774 4102 808 4136
rect 774 4030 808 4064
rect 774 3957 808 3991
rect 774 3884 808 3918
rect 774 3811 808 3845
rect 1833 4450 1867 4484
rect 1901 4450 1935 4484
rect 1969 4450 2003 4484
rect 2037 4450 2071 4484
rect 2105 4450 2139 4484
rect 2173 4450 2207 4484
rect 2241 4450 2275 4484
rect 1833 4379 1867 4413
rect 1901 4379 1935 4413
rect 1969 4379 2003 4413
rect 2037 4379 2071 4413
rect 2105 4379 2139 4413
rect 2173 4379 2207 4413
rect 2241 4379 2275 4413
rect 1833 4308 1867 4342
rect 1901 4308 1935 4342
rect 1969 4308 2003 4342
rect 2037 4308 2071 4342
rect 2105 4308 2139 4342
rect 2173 4308 2207 4342
rect 2241 4308 2275 4342
rect 1833 4237 1867 4271
rect 1901 4237 1935 4271
rect 1969 4237 2003 4271
rect 2037 4237 2071 4271
rect 2105 4237 2139 4271
rect 2173 4237 2207 4271
rect 2241 4237 2275 4271
rect 1833 4166 1867 4200
rect 1901 4166 1935 4200
rect 1969 4166 2003 4200
rect 2037 4166 2071 4200
rect 2105 4166 2139 4200
rect 2173 4166 2207 4200
rect 2241 4166 2275 4200
rect 1833 4095 1867 4129
rect 1901 4095 1935 4129
rect 1969 4095 2003 4129
rect 2037 4095 2071 4129
rect 2105 4095 2139 4129
rect 2173 4095 2207 4129
rect 2241 4095 2275 4129
rect 1833 4024 1867 4058
rect 1901 4024 1935 4058
rect 1969 4024 2003 4058
rect 2037 4024 2071 4058
rect 2105 4024 2139 4058
rect 2173 4024 2207 4058
rect 2241 4024 2275 4058
rect 1833 3953 1867 3987
rect 1901 3953 1935 3987
rect 1969 3953 2003 3987
rect 2037 3953 2071 3987
rect 2105 3953 2139 3987
rect 2173 3953 2207 3987
rect 2241 3953 2275 3987
rect 1833 3882 1867 3916
rect 1901 3882 1935 3916
rect 1969 3882 2003 3916
rect 2037 3882 2071 3916
rect 2105 3882 2139 3916
rect 2173 3882 2207 3916
rect 2241 3882 2275 3916
rect 1833 3811 1867 3845
rect 1901 3811 1935 3845
rect 1969 3811 2003 3845
rect 2037 3811 2071 3845
rect 2105 3811 2139 3845
rect 2173 3811 2207 3845
rect 2241 3811 2275 3845
rect -503 3671 619 3773
rect 654 3739 688 3773
rect 723 3739 757 3773
rect 792 3739 826 3773
rect 861 3739 895 3773
rect 930 3739 964 3773
rect 999 3739 1033 3773
rect 1068 3739 1102 3773
rect 1137 3739 1171 3773
rect 1206 3739 1240 3773
rect 1275 3739 1309 3773
rect 1344 3739 1378 3773
rect 1413 3739 1447 3773
rect 1482 3739 1516 3773
rect 1551 3739 1585 3773
rect 1620 3739 1654 3773
rect 1689 3739 1723 3773
rect 1758 3739 1792 3773
rect 1827 3739 1861 3773
rect 1896 3739 1930 3773
rect 1965 3739 1999 3773
rect 2034 3739 2068 3773
rect 2103 3739 2137 3773
rect 2172 3739 2206 3773
rect 2241 3739 2275 3773
rect 654 3671 688 3705
rect 723 3671 757 3705
rect 792 3671 826 3705
rect 861 3671 895 3705
rect 930 3671 964 3705
rect 999 3671 1033 3705
rect 1068 3671 1102 3705
rect 1137 3671 1171 3705
rect 1206 3671 1240 3705
rect 1275 3671 1309 3705
rect 1344 3671 1378 3705
rect 1413 3671 1447 3705
rect 1482 3671 1516 3705
rect 1551 3671 1585 3705
rect 1620 3671 1654 3705
rect 1689 3671 1723 3705
rect 1758 3671 1792 3705
rect 1827 3671 1861 3705
rect 1896 3671 1930 3705
rect 1965 3671 1999 3705
rect 2034 3671 2068 3705
rect 2103 3671 2137 3705
rect 2172 3671 2206 3705
rect 2241 3671 2275 3705
<< poly >>
rect -172 5516 284 5532
rect -172 5482 -156 5516
rect -122 5482 -78 5516
rect -44 5482 0 5516
rect 34 5482 78 5516
rect 112 5482 156 5516
rect 190 5482 234 5516
rect 268 5482 284 5516
rect -172 5466 284 5482
rect 340 5516 796 5532
rect 340 5482 356 5516
rect 390 5482 434 5516
rect 468 5482 512 5516
rect 546 5482 590 5516
rect 624 5482 668 5516
rect 702 5482 746 5516
rect 780 5482 796 5516
rect 340 5466 796 5482
rect 852 5516 1308 5532
rect 852 5482 868 5516
rect 902 5482 946 5516
rect 980 5482 1024 5516
rect 1058 5482 1102 5516
rect 1136 5482 1180 5516
rect 1214 5482 1258 5516
rect 1292 5482 1308 5516
rect 852 5466 1308 5482
rect 1364 5516 1820 5532
rect 1364 5482 1380 5516
rect 1414 5482 1458 5516
rect 1492 5482 1536 5516
rect 1570 5482 1614 5516
rect 1648 5482 1692 5516
rect 1726 5482 1770 5516
rect 1804 5482 1820 5516
rect 1364 5466 1820 5482
rect 1162 4550 1458 4566
rect 1162 4516 1178 4550
rect 1212 4516 1255 4550
rect 1289 4516 1332 4550
rect 1366 4516 1408 4550
rect 1442 4516 1458 4550
rect 1162 4500 1458 4516
rect 1514 4550 1648 4566
rect 1514 4516 1530 4550
rect 1564 4516 1598 4550
rect 1632 4516 1648 4550
rect 1514 4500 1648 4516
rect 260 4361 394 4377
rect 260 4327 276 4361
rect 310 4327 344 4361
rect 378 4327 394 4361
rect 260 4311 394 4327
rect 450 4361 584 4377
rect 450 4327 466 4361
rect 500 4327 534 4361
rect 568 4327 584 4361
rect 450 4311 584 4327
rect 274 4186 570 4202
rect 274 4152 290 4186
rect 324 4152 367 4186
rect 401 4152 444 4186
rect 478 4152 520 4186
rect 554 4152 570 4186
rect 274 4136 570 4152
rect 2378 934 2444 950
rect 2378 900 2394 934
rect 2428 900 2444 934
rect 2378 866 2444 900
rect 2378 832 2394 866
rect 2428 832 2444 866
rect 2378 816 2444 832
rect 170 700 970 716
rect 170 666 186 700
rect 220 666 260 700
rect 294 666 334 700
rect 368 666 408 700
rect 442 666 482 700
rect 516 666 555 700
rect 589 666 628 700
rect 662 666 701 700
rect 735 666 774 700
rect 808 666 847 700
rect 881 666 920 700
rect 954 666 970 700
rect 170 650 970 666
rect 1026 700 2626 716
rect 1026 666 1042 700
rect 1076 666 1112 700
rect 1146 666 1182 700
rect 1216 666 1252 700
rect 1286 666 1322 700
rect 1356 666 1392 700
rect 1426 666 1462 700
rect 1496 666 1532 700
rect 1566 666 1602 700
rect 1636 666 1672 700
rect 1706 666 1742 700
rect 1776 666 1812 700
rect 1846 666 1882 700
rect 1916 666 1952 700
rect 1986 666 2022 700
rect 2056 666 2092 700
rect 2126 666 2162 700
rect 2196 666 2231 700
rect 2265 666 2300 700
rect 2334 666 2369 700
rect 2403 666 2438 700
rect 2472 666 2507 700
rect 2541 666 2576 700
rect 2610 666 2626 700
rect 1026 650 2626 666
rect 170 328 970 344
rect 170 294 186 328
rect 220 294 260 328
rect 294 294 334 328
rect 368 294 408 328
rect 442 294 482 328
rect 516 294 555 328
rect 589 294 628 328
rect 662 294 701 328
rect 735 294 774 328
rect 808 294 847 328
rect 881 294 920 328
rect 954 294 970 328
rect 170 278 970 294
rect 1026 328 2626 344
rect 1026 294 1042 328
rect 1076 294 1112 328
rect 1146 294 1182 328
rect 1216 294 1252 328
rect 1286 294 1322 328
rect 1356 294 1392 328
rect 1426 294 1462 328
rect 1496 294 1532 328
rect 1566 294 1602 328
rect 1636 294 1672 328
rect 1706 294 1742 328
rect 1776 294 1812 328
rect 1846 294 1882 328
rect 1916 294 1952 328
rect 1986 294 2022 328
rect 2056 294 2092 328
rect 2126 294 2162 328
rect 2196 294 2231 328
rect 2265 294 2300 328
rect 2334 294 2369 328
rect 2403 294 2438 328
rect 2472 294 2507 328
rect 2541 294 2576 328
rect 2610 294 2626 328
rect 1026 278 2626 294
rect 1956 -70 2356 -54
rect 1956 -104 1972 -70
rect 2006 -104 2056 -70
rect 2090 -104 2140 -70
rect 2174 -104 2223 -70
rect 2257 -104 2306 -70
rect 2340 -104 2356 -70
rect 1956 -120 2356 -104
rect 912 -242 978 -226
rect 912 -276 928 -242
rect 962 -276 978 -242
rect 912 -310 978 -276
rect 912 -344 928 -310
rect 962 -344 978 -310
rect 912 -360 978 -344
rect 912 -432 978 -416
rect 912 -466 928 -432
rect 962 -466 978 -432
rect 912 -500 978 -466
rect 1906 -442 2762 -426
rect 1906 -476 1922 -442
rect 1956 -476 1993 -442
rect 2027 -476 2064 -442
rect 2098 -476 2135 -442
rect 2169 -476 2206 -442
rect 2240 -476 2276 -442
rect 2310 -476 2346 -442
rect 2380 -476 2416 -442
rect 2450 -476 2486 -442
rect 2520 -476 2556 -442
rect 2590 -476 2626 -442
rect 2660 -476 2762 -442
rect 1906 -492 2762 -476
rect 912 -534 928 -500
rect 962 -534 978 -500
rect 912 -550 978 -534
<< polycont >>
rect -156 5482 -122 5516
rect -78 5482 -44 5516
rect 0 5482 34 5516
rect 78 5482 112 5516
rect 156 5482 190 5516
rect 234 5482 268 5516
rect 356 5482 390 5516
rect 434 5482 468 5516
rect 512 5482 546 5516
rect 590 5482 624 5516
rect 668 5482 702 5516
rect 746 5482 780 5516
rect 868 5482 902 5516
rect 946 5482 980 5516
rect 1024 5482 1058 5516
rect 1102 5482 1136 5516
rect 1180 5482 1214 5516
rect 1258 5482 1292 5516
rect 1380 5482 1414 5516
rect 1458 5482 1492 5516
rect 1536 5482 1570 5516
rect 1614 5482 1648 5516
rect 1692 5482 1726 5516
rect 1770 5482 1804 5516
rect 1178 4516 1212 4550
rect 1255 4516 1289 4550
rect 1332 4516 1366 4550
rect 1408 4516 1442 4550
rect 1530 4516 1564 4550
rect 1598 4516 1632 4550
rect 276 4327 310 4361
rect 344 4327 378 4361
rect 466 4327 500 4361
rect 534 4327 568 4361
rect 290 4152 324 4186
rect 367 4152 401 4186
rect 444 4152 478 4186
rect 520 4152 554 4186
rect 2394 900 2428 934
rect 2394 832 2428 866
rect 186 666 220 700
rect 260 666 294 700
rect 334 666 368 700
rect 408 666 442 700
rect 482 666 516 700
rect 555 666 589 700
rect 628 666 662 700
rect 701 666 735 700
rect 774 666 808 700
rect 847 666 881 700
rect 920 666 954 700
rect 1042 666 1076 700
rect 1112 666 1146 700
rect 1182 666 1216 700
rect 1252 666 1286 700
rect 1322 666 1356 700
rect 1392 666 1426 700
rect 1462 666 1496 700
rect 1532 666 1566 700
rect 1602 666 1636 700
rect 1672 666 1706 700
rect 1742 666 1776 700
rect 1812 666 1846 700
rect 1882 666 1916 700
rect 1952 666 1986 700
rect 2022 666 2056 700
rect 2092 666 2126 700
rect 2162 666 2196 700
rect 2231 666 2265 700
rect 2300 666 2334 700
rect 2369 666 2403 700
rect 2438 666 2472 700
rect 2507 666 2541 700
rect 2576 666 2610 700
rect 186 294 220 328
rect 260 294 294 328
rect 334 294 368 328
rect 408 294 442 328
rect 482 294 516 328
rect 555 294 589 328
rect 628 294 662 328
rect 701 294 735 328
rect 774 294 808 328
rect 847 294 881 328
rect 920 294 954 328
rect 1042 294 1076 328
rect 1112 294 1146 328
rect 1182 294 1216 328
rect 1252 294 1286 328
rect 1322 294 1356 328
rect 1392 294 1426 328
rect 1462 294 1496 328
rect 1532 294 1566 328
rect 1602 294 1636 328
rect 1672 294 1706 328
rect 1742 294 1776 328
rect 1812 294 1846 328
rect 1882 294 1916 328
rect 1952 294 1986 328
rect 2022 294 2056 328
rect 2092 294 2126 328
rect 2162 294 2196 328
rect 2231 294 2265 328
rect 2300 294 2334 328
rect 2369 294 2403 328
rect 2438 294 2472 328
rect 2507 294 2541 328
rect 2576 294 2610 328
rect 1972 -104 2006 -70
rect 2056 -104 2090 -70
rect 2140 -104 2174 -70
rect 2223 -104 2257 -70
rect 2306 -104 2340 -70
rect 928 -276 962 -242
rect 928 -344 962 -310
rect 928 -466 962 -432
rect 1922 -476 1956 -442
rect 1993 -476 2027 -442
rect 2064 -476 2098 -442
rect 2135 -476 2169 -442
rect 2206 -476 2240 -442
rect 2276 -476 2310 -442
rect 2346 -476 2380 -442
rect 2416 -476 2450 -442
rect 2486 -476 2520 -442
rect 2556 -476 2590 -442
rect 2626 -476 2660 -442
rect 928 -534 962 -500
<< locali >>
rect 210 5855 2303 5861
rect 210 5848 242 5855
rect -537 5821 242 5848
rect 276 5821 316 5855
rect 350 5821 390 5855
rect 424 5821 464 5855
rect 498 5821 538 5855
rect 572 5821 612 5855
rect 646 5821 686 5855
rect 720 5821 760 5855
rect 794 5821 834 5855
rect 868 5821 908 5855
rect 942 5821 982 5855
rect 1016 5821 1056 5855
rect 1090 5821 1130 5855
rect 1164 5821 1204 5855
rect 1238 5821 1278 5855
rect 1312 5821 1352 5855
rect 1386 5821 1426 5855
rect 1460 5821 1500 5855
rect 1534 5821 1574 5855
rect 1608 5821 1648 5855
rect 1682 5821 1722 5855
rect 1756 5821 1796 5855
rect 1830 5821 1870 5855
rect 1904 5821 1944 5855
rect 1978 5821 2018 5855
rect 2052 5821 2091 5855
rect 2125 5821 2164 5855
rect 2198 5821 2237 5855
rect 2271 5836 2303 5855
rect 2271 5821 2309 5836
rect -537 5814 2309 5821
rect -537 5802 -503 5814
rect -537 5768 -531 5802
rect -469 5780 -435 5814
rect -401 5780 -367 5814
rect -333 5802 -263 5814
rect -305 5780 -263 5802
rect -229 5780 -194 5814
rect -160 5780 -125 5814
rect -91 5780 -56 5814
rect -22 5780 13 5814
rect 47 5780 82 5814
rect 116 5780 151 5814
rect 185 5780 220 5814
rect 254 5780 289 5814
rect 323 5780 358 5814
rect 392 5780 427 5814
rect 461 5780 496 5814
rect 530 5780 565 5814
rect 599 5780 634 5814
rect 668 5780 703 5814
rect 737 5780 772 5814
rect 806 5780 841 5814
rect 875 5780 910 5814
rect 944 5780 979 5814
rect 1013 5780 1048 5814
rect 1082 5780 1117 5814
rect 1151 5780 1186 5814
rect 1220 5780 1255 5814
rect 1289 5780 1324 5814
rect 1358 5780 1393 5814
rect 1427 5780 1462 5814
rect 1496 5780 1531 5814
rect 1565 5780 1600 5814
rect 1634 5780 1669 5814
rect 1703 5780 1738 5814
rect 1772 5780 1807 5814
rect -497 5768 -435 5780
rect -401 5768 -339 5780
rect -305 5772 1807 5780
rect 1977 5802 2309 5814
rect 1977 5772 2037 5802
rect 2071 5772 2105 5802
rect 2139 5772 2173 5802
rect 2207 5772 2241 5802
rect -305 5768 242 5772
rect -537 5746 242 5768
rect 276 5746 316 5772
rect 350 5746 390 5772
rect 424 5746 464 5772
rect 498 5746 538 5772
rect 572 5746 612 5772
rect 646 5746 686 5772
rect 720 5746 760 5772
rect 794 5746 834 5772
rect 868 5746 908 5772
rect 942 5746 982 5772
rect 1016 5746 1056 5772
rect 1090 5746 1130 5772
rect 1164 5746 1204 5772
rect 1238 5746 1278 5772
rect 1312 5746 1352 5772
rect 1386 5746 1426 5772
rect 1460 5746 1500 5772
rect 1534 5746 1574 5772
rect 1608 5746 1648 5772
rect 1682 5746 1722 5772
rect 1756 5746 1796 5772
rect -537 5744 -263 5746
rect -537 5728 -503 5744
rect -537 5694 -531 5728
rect -469 5710 -435 5744
rect -401 5710 -367 5744
rect -333 5728 -263 5744
rect -305 5712 -263 5728
rect -229 5712 -194 5746
rect -160 5712 -125 5746
rect -91 5712 -56 5746
rect -22 5712 13 5746
rect 47 5712 82 5746
rect 116 5712 151 5746
rect 185 5712 220 5746
rect 276 5738 289 5746
rect 350 5738 358 5746
rect 424 5738 427 5746
rect 254 5712 289 5738
rect 323 5712 358 5738
rect 392 5712 427 5738
rect 461 5738 464 5746
rect 530 5738 538 5746
rect 599 5738 612 5746
rect 668 5738 686 5746
rect 737 5738 760 5746
rect 806 5738 834 5746
rect 875 5738 908 5746
rect 461 5712 496 5738
rect 530 5712 565 5738
rect 599 5712 634 5738
rect 668 5712 703 5738
rect 737 5712 772 5738
rect 806 5712 841 5738
rect 875 5712 910 5738
rect 944 5712 979 5746
rect 1016 5738 1048 5746
rect 1090 5738 1117 5746
rect 1164 5738 1186 5746
rect 1238 5738 1255 5746
rect 1312 5738 1324 5746
rect 1386 5738 1393 5746
rect 1460 5738 1462 5746
rect 1013 5712 1048 5738
rect 1082 5712 1117 5738
rect 1151 5712 1186 5738
rect 1220 5712 1255 5738
rect 1289 5712 1324 5738
rect 1358 5712 1393 5738
rect 1427 5712 1462 5738
rect 1496 5738 1500 5746
rect 1565 5738 1574 5746
rect 1634 5738 1648 5746
rect 1703 5738 1722 5746
rect 1772 5738 1796 5746
rect 1978 5738 2018 5772
rect 2071 5768 2091 5772
rect 2139 5768 2164 5772
rect 2207 5768 2237 5772
rect 2275 5768 2309 5802
rect 2052 5738 2091 5768
rect 2125 5738 2164 5768
rect 2198 5738 2237 5768
rect 2271 5738 2309 5768
rect 1496 5712 1531 5738
rect 1565 5712 1600 5738
rect 1634 5712 1669 5738
rect 1703 5712 1738 5738
rect 1772 5712 1807 5738
rect -497 5694 -435 5710
rect -401 5694 -339 5710
rect -305 5694 1807 5712
rect -537 5689 1807 5694
rect 1977 5731 2309 5738
rect 1977 5697 2037 5731
rect 2071 5697 2105 5731
rect 2139 5697 2173 5731
rect 2207 5697 2241 5731
rect 2275 5697 2309 5731
rect 1977 5689 2309 5697
rect -537 5678 242 5689
rect 276 5678 316 5689
rect 350 5678 390 5689
rect 424 5678 464 5689
rect 498 5678 538 5689
rect 572 5678 612 5689
rect 646 5678 686 5689
rect 720 5678 760 5689
rect 794 5678 834 5689
rect 868 5678 908 5689
rect 942 5678 982 5689
rect 1016 5678 1056 5689
rect 1090 5678 1130 5689
rect 1164 5678 1204 5689
rect 1238 5678 1278 5689
rect 1312 5678 1352 5689
rect 1386 5678 1426 5689
rect 1460 5678 1500 5689
rect 1534 5678 1574 5689
rect 1608 5678 1648 5689
rect 1682 5678 1722 5689
rect 1756 5678 1796 5689
rect -537 5674 -263 5678
rect -537 5654 -503 5674
rect -537 5620 -531 5654
rect -469 5640 -435 5674
rect -401 5640 -367 5674
rect -333 5654 -263 5674
rect -305 5644 -263 5654
rect -229 5644 -194 5678
rect -160 5644 -125 5678
rect -91 5644 -56 5678
rect -22 5644 13 5678
rect 47 5644 82 5678
rect 116 5644 151 5678
rect 185 5644 220 5678
rect 276 5655 289 5678
rect 350 5655 358 5678
rect 424 5655 427 5678
rect 254 5644 289 5655
rect 323 5644 358 5655
rect 392 5644 427 5655
rect 461 5655 464 5678
rect 530 5655 538 5678
rect 599 5655 612 5678
rect 668 5655 686 5678
rect 737 5655 760 5678
rect 806 5655 834 5678
rect 875 5655 908 5678
rect 461 5644 496 5655
rect 530 5644 565 5655
rect 599 5644 634 5655
rect 668 5644 703 5655
rect 737 5644 772 5655
rect 806 5644 841 5655
rect 875 5644 910 5655
rect 944 5644 979 5678
rect 1016 5655 1048 5678
rect 1090 5655 1117 5678
rect 1164 5655 1186 5678
rect 1238 5655 1255 5678
rect 1312 5655 1324 5678
rect 1386 5655 1393 5678
rect 1460 5655 1462 5678
rect 1013 5644 1048 5655
rect 1082 5644 1117 5655
rect 1151 5644 1186 5655
rect 1220 5644 1255 5655
rect 1289 5644 1324 5655
rect 1358 5644 1393 5655
rect 1427 5644 1462 5655
rect 1496 5655 1500 5678
rect 1565 5655 1574 5678
rect 1634 5655 1648 5678
rect 1703 5655 1722 5678
rect 1772 5655 1796 5678
rect 1978 5655 2018 5689
rect 2052 5660 2091 5689
rect 2125 5660 2164 5689
rect 2198 5660 2237 5689
rect 2271 5660 2309 5689
rect 2071 5655 2091 5660
rect 2139 5655 2164 5660
rect 2207 5655 2237 5660
rect 1496 5644 1531 5655
rect 1565 5644 1600 5655
rect 1634 5644 1669 5655
rect 1703 5644 1738 5655
rect 1772 5644 1807 5655
rect 1977 5644 2037 5655
rect -497 5620 -435 5640
rect -401 5620 -339 5640
rect -305 5626 2037 5644
rect 2071 5626 2105 5655
rect 2139 5626 2173 5655
rect 2207 5626 2241 5655
rect 2275 5626 2309 5660
rect -305 5620 2309 5626
rect -537 5610 2309 5620
rect -537 5609 -261 5610
rect -537 5604 -299 5609
rect -537 5580 -503 5604
rect -537 5546 -531 5580
rect -469 5570 -435 5604
rect -401 5570 -367 5604
rect -333 5580 -299 5604
rect -497 5546 -435 5570
rect -401 5546 -339 5570
rect -305 5546 -299 5580
rect -537 5534 -299 5546
rect -537 5506 -503 5534
rect -537 5472 -531 5506
rect -469 5500 -435 5534
rect -401 5500 -367 5534
rect -333 5506 -299 5534
rect 1970 5589 2309 5610
rect 1970 5577 2037 5589
rect 2071 5577 2105 5589
rect 2139 5577 2173 5589
rect 2207 5577 2241 5589
rect 2275 5577 2309 5589
rect 2004 5555 2037 5577
rect 2076 5555 2105 5577
rect 2148 5555 2173 5577
rect 2220 5555 2241 5577
rect 2004 5543 2042 5555
rect 2076 5543 2114 5555
rect 2148 5543 2186 5555
rect 2220 5543 2258 5555
rect 2292 5543 2309 5577
rect 1970 5518 2309 5543
rect 107 5516 156 5517
rect 190 5516 238 5517
rect 442 5516 527 5517
rect 898 5516 947 5517
rect 981 5516 1029 5517
rect 1479 5516 1528 5517
rect 1562 5516 1610 5517
rect -497 5472 -435 5500
rect -401 5472 -339 5500
rect -305 5472 -299 5506
rect -172 5482 -156 5516
rect -122 5482 -78 5516
rect -44 5482 0 5516
rect 34 5483 73 5516
rect 34 5482 78 5483
rect 112 5482 156 5516
rect 190 5482 234 5516
rect 272 5483 284 5516
rect 268 5482 284 5483
rect 340 5482 356 5516
rect 390 5483 408 5516
rect 390 5482 434 5483
rect 468 5482 512 5516
rect 561 5483 590 5516
rect 546 5482 590 5483
rect 624 5482 668 5516
rect 702 5482 746 5516
rect 780 5482 796 5516
rect 852 5483 864 5516
rect 852 5482 868 5483
rect 902 5482 946 5516
rect 981 5483 1024 5516
rect 1063 5483 1102 5516
rect 980 5482 1024 5483
rect 1058 5482 1102 5483
rect 1136 5482 1180 5516
rect 1214 5482 1258 5516
rect 1292 5482 1308 5516
rect 1364 5482 1380 5516
rect 1414 5483 1445 5516
rect 1492 5483 1528 5516
rect 1570 5483 1610 5516
rect 1414 5482 1458 5483
rect 1492 5482 1536 5483
rect 1570 5482 1614 5483
rect 1648 5482 1692 5516
rect 1726 5482 1770 5516
rect 1804 5482 1820 5516
rect 1970 5503 2037 5518
rect 2071 5503 2105 5518
rect 2139 5503 2173 5518
rect 2207 5503 2241 5518
rect 2275 5503 2309 5518
rect -537 5464 -299 5472
rect -537 5432 -503 5464
rect -537 5398 -531 5432
rect -469 5430 -435 5464
rect -401 5430 -367 5464
rect -333 5432 -299 5464
rect -497 5398 -435 5430
rect -401 5398 -339 5430
rect -305 5398 -299 5432
rect 2004 5484 2037 5503
rect 2076 5484 2105 5503
rect 2148 5484 2173 5503
rect 2220 5484 2241 5503
rect 2004 5469 2042 5484
rect 2076 5469 2114 5484
rect 2148 5469 2186 5484
rect 2220 5469 2258 5484
rect 2292 5469 2309 5503
rect 1970 5446 2309 5469
rect 1970 5428 2037 5446
rect 2071 5428 2105 5446
rect 2139 5428 2173 5446
rect 2207 5428 2241 5446
rect 2275 5428 2309 5446
rect -537 5394 -299 5398
rect -537 5360 -503 5394
rect -469 5360 -435 5394
rect -401 5360 -367 5394
rect -333 5360 -299 5394
rect -537 5358 -299 5360
rect -537 5324 -531 5358
rect -497 5324 -435 5358
rect -401 5324 -339 5358
rect -305 5324 -299 5358
rect -537 5290 -503 5324
rect -469 5290 -435 5324
rect -401 5290 -367 5324
rect -333 5290 -299 5324
rect 39 5334 73 5392
rect -537 5284 -299 5290
rect -537 5250 -531 5284
rect -497 5254 -435 5284
rect -401 5254 -339 5284
rect -537 5220 -503 5250
rect -469 5220 -435 5254
rect -401 5220 -367 5254
rect -305 5250 -299 5284
rect -333 5220 -299 5250
rect -537 5210 -299 5220
rect -537 5176 -531 5210
rect -497 5184 -435 5210
rect -401 5184 -339 5210
rect -537 5150 -503 5176
rect -469 5150 -435 5184
rect -401 5150 -367 5184
rect -305 5176 -299 5210
rect -333 5150 -299 5176
rect -537 5136 -299 5150
rect -537 5102 -531 5136
rect -497 5114 -435 5136
rect -401 5114 -339 5136
rect -537 5080 -503 5102
rect -469 5080 -435 5114
rect -401 5080 -367 5114
rect -305 5102 -299 5136
rect -333 5080 -299 5102
rect -537 5062 -299 5080
rect -537 5028 -531 5062
rect -497 5044 -435 5062
rect -401 5044 -339 5062
rect -537 5010 -503 5028
rect -469 5010 -435 5044
rect -401 5010 -367 5044
rect -305 5028 -299 5062
rect -333 5010 -299 5028
rect -537 4988 -299 5010
rect -537 4954 -531 4988
rect -497 4974 -435 4988
rect -401 4974 -339 4988
rect -537 4940 -503 4954
rect -469 4940 -435 4974
rect -401 4940 -367 4974
rect -305 4954 -299 4988
rect -333 4940 -299 4954
rect -537 4914 -299 4940
rect -537 4880 -531 4914
rect -497 4904 -435 4914
rect -401 4904 -339 4914
rect -537 4870 -503 4880
rect -469 4870 -435 4904
rect -401 4870 -367 4904
rect -305 4880 -299 4914
rect -333 4870 -299 4880
rect -537 4840 -299 4870
rect -217 5221 -183 5272
rect -217 5136 -183 5187
rect 551 5349 585 5392
rect 39 5241 73 5300
rect 39 5148 73 5207
rect 295 5221 329 5272
rect 295 5136 329 5187
rect -217 5051 -183 5102
rect -217 4966 -183 5017
rect -217 4880 -183 4932
rect 295 5051 329 5102
rect 295 4966 329 5017
rect 551 5271 585 5315
rect 1063 5349 1097 5392
rect 1063 5271 1097 5315
rect 1575 5349 1609 5392
rect 551 5193 585 5237
rect 551 5115 585 5159
rect 551 5037 585 5081
rect 807 5150 841 5205
rect 807 5060 841 5116
rect 295 4880 329 4932
rect 807 4970 841 5026
rect 1063 5193 1097 5237
rect 1063 5115 1097 5159
rect 1063 5037 1097 5081
rect 1319 5221 1353 5272
rect 1319 5136 1353 5187
rect 1319 5051 1353 5102
rect 807 4880 841 4936
rect 1319 4966 1353 5017
rect 1575 5271 1609 5315
rect 2004 5412 2037 5428
rect 2076 5412 2105 5428
rect 2148 5412 2173 5428
rect 2220 5412 2241 5428
rect 2004 5394 2042 5412
rect 2076 5394 2114 5412
rect 2148 5394 2186 5412
rect 2220 5394 2258 5412
rect 2292 5394 2309 5428
rect 1970 5374 2309 5394
rect 1970 5353 2037 5374
rect 2071 5353 2105 5374
rect 2139 5353 2173 5374
rect 2207 5353 2241 5374
rect 2275 5353 2309 5374
rect 2004 5340 2037 5353
rect 2076 5340 2105 5353
rect 2148 5340 2173 5353
rect 2220 5340 2241 5353
rect 2004 5319 2042 5340
rect 2076 5319 2114 5340
rect 2148 5319 2186 5340
rect 2220 5319 2258 5340
rect 2292 5319 2309 5353
rect 1970 5302 2309 5319
rect 1970 5278 2037 5302
rect 2071 5278 2105 5302
rect 2139 5278 2173 5302
rect 2207 5278 2241 5302
rect 2275 5278 2309 5302
rect 1575 5193 1609 5237
rect 1575 5115 1609 5159
rect 1575 5037 1609 5081
rect 1831 5176 1865 5215
rect 1831 5102 1865 5142
rect 1831 5028 1865 5068
rect 1319 4880 1353 4932
rect 1831 4954 1865 4994
rect 1831 4880 1865 4920
rect 2004 5268 2037 5278
rect 2076 5268 2105 5278
rect 2148 5268 2173 5278
rect 2220 5268 2241 5278
rect 2004 5244 2042 5268
rect 2076 5244 2114 5268
rect 2148 5244 2186 5268
rect 2220 5244 2258 5268
rect 2292 5244 2309 5278
rect 1970 5230 2309 5244
rect 1970 5203 2037 5230
rect 2071 5203 2105 5230
rect 2139 5203 2173 5230
rect 2207 5203 2241 5230
rect 2275 5203 2309 5230
rect 2004 5196 2037 5203
rect 2076 5196 2105 5203
rect 2148 5196 2173 5203
rect 2220 5196 2241 5203
rect 2004 5169 2042 5196
rect 2076 5169 2114 5196
rect 2148 5169 2186 5196
rect 2220 5169 2258 5196
rect 2292 5169 2309 5203
rect 1970 5158 2309 5169
rect 1970 5128 2037 5158
rect 2071 5128 2105 5158
rect 2139 5128 2173 5158
rect 2207 5128 2241 5158
rect 2275 5128 2309 5158
rect 2004 5124 2037 5128
rect 2076 5124 2105 5128
rect 2148 5124 2173 5128
rect 2220 5124 2241 5128
rect 2004 5094 2042 5124
rect 2076 5094 2114 5124
rect 2148 5094 2186 5124
rect 2220 5094 2258 5124
rect 2292 5094 2309 5128
rect 1970 5086 2309 5094
rect 1970 5053 2037 5086
rect 2071 5053 2105 5086
rect 2139 5053 2173 5086
rect 2207 5053 2241 5086
rect 2275 5053 2309 5086
rect 2004 5052 2037 5053
rect 2076 5052 2105 5053
rect 2148 5052 2173 5053
rect 2220 5052 2241 5053
rect 2004 5019 2042 5052
rect 2076 5019 2114 5052
rect 2148 5019 2186 5052
rect 2220 5019 2258 5052
rect 2292 5019 2309 5053
rect 1970 5014 2309 5019
rect 1970 4980 2037 5014
rect 2071 4980 2105 5014
rect 2139 4980 2173 5014
rect 2207 4980 2241 5014
rect 2275 4980 2309 5014
rect 1970 4978 2309 4980
rect 2004 4944 2042 4978
rect 2076 4944 2114 4978
rect 2148 4944 2186 4978
rect 2220 4944 2258 4978
rect 2292 4944 2309 4978
rect 1970 4942 2309 4944
rect 1970 4908 2037 4942
rect 2071 4908 2105 4942
rect 2139 4908 2173 4942
rect 2207 4908 2241 4942
rect 2275 4908 2309 4942
rect 1970 4903 2309 4908
rect 2004 4870 2042 4903
rect 2076 4870 2114 4903
rect 2148 4870 2186 4903
rect 2220 4870 2258 4903
rect 2004 4869 2037 4870
rect 2076 4869 2105 4870
rect 2148 4869 2173 4870
rect 2220 4869 2241 4870
rect 2292 4869 2309 4903
rect -537 4806 -531 4840
rect -497 4834 -435 4840
rect -401 4834 -339 4840
rect -537 4800 -503 4806
rect -469 4800 -435 4834
rect -401 4800 -367 4834
rect -305 4806 -299 4840
rect -333 4800 -299 4806
rect -537 4766 -299 4800
rect -537 4732 -531 4766
rect -497 4764 -435 4766
rect -401 4764 -339 4766
rect -537 4730 -503 4732
rect -469 4730 -435 4764
rect -401 4730 -367 4764
rect -305 4760 -299 4766
rect 1970 4836 2037 4869
rect 2071 4836 2105 4869
rect 2139 4836 2173 4869
rect 2207 4836 2241 4869
rect 2275 4836 2309 4869
rect 1970 4828 2309 4836
rect 2004 4798 2042 4828
rect 2076 4798 2114 4828
rect 2148 4798 2186 4828
rect 2220 4798 2258 4828
rect 2004 4794 2037 4798
rect 2076 4794 2105 4798
rect 2148 4794 2173 4798
rect 2220 4794 2241 4798
rect 2292 4794 2309 4828
rect 1970 4764 2037 4794
rect 2071 4764 2105 4794
rect 2139 4764 2173 4794
rect 2207 4764 2241 4794
rect 2275 4764 2309 4794
rect 1970 4760 2309 4764
rect -305 4732 2309 4760
rect -333 4730 2309 4732
rect -537 4729 2309 4730
rect -537 4726 -198 4729
rect -164 4726 -125 4729
rect -91 4726 -52 4729
rect -18 4726 21 4729
rect 55 4726 94 4729
rect 128 4726 167 4729
rect 201 4726 240 4729
rect 274 4726 312 4729
rect 346 4726 384 4729
rect 418 4726 456 4729
rect 490 4726 528 4729
rect -537 4694 -265 4726
rect -537 4692 -503 4694
rect -537 4658 -531 4692
rect -469 4660 -435 4694
rect -401 4660 -367 4694
rect -333 4692 -265 4694
rect -231 4695 -198 4726
rect -231 4692 -196 4695
rect -162 4692 -127 4726
rect -91 4695 -58 4726
rect -18 4695 11 4726
rect 55 4695 80 4726
rect 128 4695 149 4726
rect 201 4695 218 4726
rect 274 4695 287 4726
rect 346 4695 356 4726
rect 418 4695 425 4726
rect 490 4695 494 4726
rect -93 4692 -58 4695
rect -24 4692 11 4695
rect 45 4692 80 4695
rect 114 4692 149 4695
rect 183 4692 218 4695
rect 252 4692 287 4695
rect 321 4692 356 4695
rect 390 4692 425 4695
rect 459 4692 494 4695
rect 562 4726 600 4729
rect 634 4726 672 4729
rect 706 4726 744 4729
rect 778 4726 816 4729
rect 850 4726 888 4729
rect 922 4726 960 4729
rect 994 4726 1032 4729
rect 1066 4726 1104 4729
rect 1138 4726 1176 4729
rect 1210 4726 1248 4729
rect 1282 4726 1320 4729
rect 1354 4726 1392 4729
rect 1426 4726 1464 4729
rect 1498 4726 1536 4729
rect 1570 4726 1608 4729
rect 1642 4726 1680 4729
rect 1714 4726 1752 4729
rect 1786 4726 1824 4729
rect 1858 4726 1896 4729
rect 1930 4726 1968 4729
rect 2002 4726 2040 4729
rect 2074 4726 2309 4729
rect 562 4695 563 4726
rect 528 4692 563 4695
rect 597 4695 600 4726
rect 666 4695 672 4726
rect 735 4695 744 4726
rect 804 4695 816 4726
rect 873 4695 888 4726
rect 942 4695 960 4726
rect 1011 4695 1032 4726
rect 1080 4695 1104 4726
rect 1149 4695 1176 4726
rect 1218 4695 1248 4726
rect 1288 4695 1320 4726
rect 1358 4695 1392 4726
rect 597 4692 632 4695
rect 666 4692 701 4695
rect 735 4692 770 4695
rect 804 4692 839 4695
rect 873 4692 908 4695
rect 942 4692 977 4695
rect 1011 4692 1046 4695
rect 1080 4692 1115 4695
rect 1149 4692 1184 4695
rect 1218 4692 1254 4695
rect 1288 4692 1324 4695
rect 1358 4692 1394 4695
rect 1428 4692 1464 4726
rect 1498 4692 1534 4726
rect 1570 4695 1604 4726
rect 1642 4695 1674 4726
rect 1714 4695 1744 4726
rect 1786 4695 1814 4726
rect 1858 4695 1884 4726
rect 1930 4695 1954 4726
rect 2002 4695 2037 4726
rect 2074 4695 2105 4726
rect 1568 4692 1604 4695
rect 1638 4692 1674 4695
rect 1708 4692 1744 4695
rect 1778 4692 1814 4695
rect 1848 4692 1884 4695
rect 1918 4692 1954 4695
rect 1988 4692 2037 4695
rect 2071 4692 2105 4695
rect 2139 4692 2173 4726
rect 2207 4692 2241 4726
rect 2275 4692 2309 4726
rect -497 4658 -435 4660
rect -401 4658 -339 4660
rect -305 4658 2309 4692
rect -537 4624 -299 4658
rect -537 4618 -503 4624
rect -537 4584 -531 4618
rect -469 4590 -435 4624
rect -401 4590 -367 4624
rect -333 4618 -299 4624
rect -497 4584 -435 4590
rect -401 4584 -339 4590
rect -305 4584 -299 4618
rect 740 4640 842 4658
rect 740 4606 774 4640
rect 808 4606 842 4640
rect -537 4554 -299 4584
rect -537 4544 -503 4554
rect -537 4510 -531 4544
rect -469 4520 -435 4554
rect -401 4520 -367 4554
rect -333 4544 -299 4554
rect -497 4510 -435 4520
rect -401 4510 -339 4520
rect -305 4510 -299 4544
rect 405 4521 439 4559
rect -537 4484 -299 4510
rect -537 4470 -503 4484
rect -537 4436 -531 4470
rect -469 4450 -435 4484
rect -401 4450 -367 4484
rect -333 4470 -299 4484
rect -497 4436 -435 4450
rect -401 4436 -339 4450
rect -305 4436 -299 4470
rect -537 4413 -299 4436
rect -537 4396 -503 4413
rect -537 4362 -531 4396
rect -469 4379 -435 4413
rect -401 4379 -367 4413
rect -333 4396 -299 4413
rect 581 4521 615 4559
rect 740 4568 842 4606
rect 740 4534 774 4568
rect 808 4534 842 4568
rect 1799 4624 2309 4658
rect 1799 4590 1833 4624
rect 1867 4590 1901 4624
rect 1935 4590 1969 4624
rect 2003 4590 2037 4624
rect 2071 4590 2105 4624
rect 2139 4590 2173 4624
rect 2207 4590 2241 4624
rect 2275 4590 2309 4624
rect 1799 4563 2309 4590
rect 740 4496 842 4534
rect 1162 4516 1174 4550
rect 1212 4516 1248 4550
rect 1289 4516 1322 4550
rect 1366 4516 1408 4550
rect 1442 4516 1458 4550
rect 1514 4516 1526 4550
rect 1564 4516 1598 4550
rect 1632 4516 1648 4550
rect 1799 4529 1827 4563
rect 1861 4554 1899 4563
rect 1933 4554 1971 4563
rect 2005 4554 2043 4563
rect 2077 4554 2115 4563
rect 2149 4554 2187 4563
rect 2221 4554 2259 4563
rect 1867 4529 1899 4554
rect 1799 4520 1833 4529
rect 1867 4520 1901 4529
rect 1935 4520 1969 4554
rect 2005 4529 2037 4554
rect 2077 4529 2105 4554
rect 2149 4529 2173 4554
rect 2221 4529 2241 4554
rect 2293 4529 2309 4563
rect 2003 4520 2037 4529
rect 2071 4520 2105 4529
rect 2139 4520 2173 4529
rect 2207 4520 2241 4529
rect 2275 4520 2309 4529
rect 229 4441 263 4479
rect 740 4462 774 4496
rect 808 4462 842 4496
rect 740 4424 842 4462
rect -497 4362 -435 4379
rect -401 4362 -339 4379
rect -305 4362 -299 4396
rect -537 4342 -299 4362
rect 740 4390 774 4424
rect 808 4390 842 4424
rect -537 4322 -503 4342
rect -537 4288 -531 4322
rect -469 4308 -435 4342
rect -401 4308 -367 4342
rect -333 4322 -299 4342
rect 260 4327 272 4361
rect 310 4327 344 4361
rect 378 4327 394 4361
rect 450 4327 462 4361
rect 500 4327 534 4361
rect 568 4327 584 4361
rect 740 4352 842 4390
rect -497 4288 -435 4308
rect -401 4288 -339 4308
rect -305 4288 -299 4322
rect -537 4271 -299 4288
rect -537 4248 -503 4271
rect -537 4214 -531 4248
rect -469 4237 -435 4271
rect -401 4237 -367 4271
rect -333 4248 -299 4271
rect -497 4214 -435 4237
rect -401 4214 -339 4237
rect -305 4214 -299 4248
rect -537 4200 -299 4214
rect -537 4174 -503 4200
rect -537 4140 -531 4174
rect -469 4166 -435 4200
rect -401 4166 -367 4200
rect -333 4174 -299 4200
rect 740 4318 774 4352
rect 808 4318 842 4352
rect 1799 4487 2309 4520
rect 1799 4453 1827 4487
rect 1861 4484 1899 4487
rect 1933 4484 1971 4487
rect 2005 4484 2043 4487
rect 2077 4484 2115 4487
rect 2149 4484 2187 4487
rect 2221 4484 2259 4487
rect 1867 4453 1899 4484
rect 1799 4450 1833 4453
rect 1867 4450 1901 4453
rect 1935 4450 1969 4484
rect 2005 4453 2037 4484
rect 2077 4453 2105 4484
rect 2149 4453 2173 4484
rect 2221 4453 2241 4484
rect 2293 4453 2309 4487
rect 2003 4450 2037 4453
rect 2071 4450 2105 4453
rect 2139 4450 2173 4453
rect 2207 4450 2241 4453
rect 2275 4450 2309 4453
rect 1799 4413 2309 4450
rect 1799 4411 1833 4413
rect 1867 4411 1901 4413
rect 1799 4377 1827 4411
rect 1867 4379 1899 4411
rect 1935 4379 1969 4413
rect 2003 4411 2037 4413
rect 2071 4411 2105 4413
rect 2139 4411 2173 4413
rect 2207 4411 2241 4413
rect 2275 4411 2309 4413
rect 2005 4379 2037 4411
rect 2077 4379 2105 4411
rect 2149 4379 2173 4411
rect 2221 4379 2241 4411
rect 1861 4377 1899 4379
rect 1933 4377 1971 4379
rect 2005 4377 2043 4379
rect 2077 4377 2115 4379
rect 2149 4377 2187 4379
rect 2221 4377 2259 4379
rect 2293 4377 2309 4411
rect 740 4280 842 4318
rect 740 4246 774 4280
rect 808 4246 842 4280
rect 740 4208 842 4246
rect -497 4140 -435 4166
rect -401 4140 -339 4166
rect -305 4140 -299 4174
rect 274 4152 290 4186
rect 324 4152 367 4186
rect 401 4152 410 4186
rect 478 4152 482 4186
rect 516 4152 520 4186
rect 554 4152 570 4186
rect 740 4174 774 4208
rect 808 4174 842 4208
rect 1293 4206 1327 4271
rect -537 4129 -299 4140
rect -537 4100 -503 4129
rect -537 4066 -531 4100
rect -469 4095 -435 4129
rect -401 4095 -367 4129
rect -333 4100 -299 4129
rect -497 4066 -435 4095
rect -401 4066 -339 4095
rect -305 4066 -299 4100
rect 740 4136 842 4174
rect 740 4102 774 4136
rect 808 4102 842 4136
rect -537 4058 -299 4066
rect -537 4026 -503 4058
rect -537 3992 -531 4026
rect -469 4024 -435 4058
rect -401 4024 -367 4058
rect -333 4026 -299 4058
rect -497 3992 -435 4024
rect -401 3992 -339 4024
rect -305 3992 -299 4026
rect 405 4024 439 4062
rect 740 4064 842 4102
rect 740 4030 774 4064
rect 808 4030 842 4064
rect -537 3987 -299 3992
rect -537 3953 -503 3987
rect -469 3953 -435 3987
rect -401 3953 -367 3987
rect -333 3953 -299 3987
rect -537 3952 -299 3953
rect -537 3918 -531 3952
rect -497 3918 -435 3952
rect -401 3918 -339 3952
rect -305 3918 -299 3952
rect 229 3952 263 3990
rect 581 3952 615 3990
rect 740 3991 842 4030
rect 740 3957 774 3991
rect 808 3957 842 3991
rect 740 3918 842 3957
rect 1117 4080 1151 4149
rect 1645 4270 1679 4317
rect 1645 4188 1679 4236
rect 1293 4106 1327 4172
rect 1469 4080 1503 4149
rect 1117 3976 1151 4046
rect 1645 4106 1679 4154
rect 1799 4342 2309 4377
rect 1799 4335 1833 4342
rect 1867 4335 1901 4342
rect 1799 4301 1827 4335
rect 1867 4308 1899 4335
rect 1935 4308 1969 4342
rect 2003 4335 2037 4342
rect 2071 4335 2105 4342
rect 2139 4335 2173 4342
rect 2207 4335 2241 4342
rect 2275 4335 2309 4342
rect 2005 4308 2037 4335
rect 2077 4308 2105 4335
rect 2149 4308 2173 4335
rect 2221 4308 2241 4335
rect 1861 4301 1899 4308
rect 1933 4301 1971 4308
rect 2005 4301 2043 4308
rect 2077 4301 2115 4308
rect 2149 4301 2187 4308
rect 2221 4301 2259 4308
rect 2293 4301 2309 4335
rect 1799 4271 2309 4301
rect 1799 4259 1833 4271
rect 1867 4259 1901 4271
rect 1799 4225 1827 4259
rect 1867 4237 1899 4259
rect 1935 4237 1969 4271
rect 2003 4259 2037 4271
rect 2071 4259 2105 4271
rect 2139 4259 2173 4271
rect 2207 4259 2241 4271
rect 2275 4259 2309 4271
rect 2005 4237 2037 4259
rect 2077 4237 2105 4259
rect 2149 4237 2173 4259
rect 2221 4237 2241 4259
rect 1861 4225 1899 4237
rect 1933 4225 1971 4237
rect 2005 4225 2043 4237
rect 2077 4225 2115 4237
rect 2149 4225 2187 4237
rect 2221 4225 2259 4237
rect 2293 4225 2309 4259
rect 1799 4200 2309 4225
rect 1799 4183 1833 4200
rect 1867 4183 1901 4200
rect 1799 4149 1827 4183
rect 1867 4166 1899 4183
rect 1935 4166 1969 4200
rect 2003 4183 2037 4200
rect 2071 4183 2105 4200
rect 2139 4183 2173 4200
rect 2207 4183 2241 4200
rect 2275 4183 2309 4200
rect 2005 4166 2037 4183
rect 2077 4166 2105 4183
rect 2149 4166 2173 4183
rect 2221 4166 2241 4183
rect 1861 4149 1899 4166
rect 1933 4149 1971 4166
rect 2005 4149 2043 4166
rect 2077 4149 2115 4166
rect 2149 4149 2187 4166
rect 2221 4149 2259 4166
rect 2293 4149 2309 4183
rect 1799 4129 2309 4149
rect 1799 4107 1833 4129
rect 1867 4107 1901 4129
rect 1799 4073 1827 4107
rect 1867 4095 1899 4107
rect 1935 4095 1969 4129
rect 2003 4107 2037 4129
rect 2071 4107 2105 4129
rect 2139 4107 2173 4129
rect 2207 4107 2241 4129
rect 2275 4107 2309 4129
rect 2005 4095 2037 4107
rect 2077 4095 2105 4107
rect 2149 4095 2173 4107
rect 2221 4095 2241 4107
rect 1861 4073 1899 4095
rect 1933 4073 1971 4095
rect 2005 4073 2043 4095
rect 2077 4073 2115 4095
rect 2149 4073 2187 4095
rect 2221 4073 2259 4095
rect 2293 4073 2309 4107
rect 1469 3976 1503 4046
rect 1799 4058 2309 4073
rect 1799 4031 1833 4058
rect 1867 4031 1901 4058
rect 1799 3997 1827 4031
rect 1867 4024 1899 4031
rect 1935 4024 1969 4058
rect 2003 4031 2037 4058
rect 2071 4031 2105 4058
rect 2139 4031 2173 4058
rect 2207 4031 2241 4058
rect 2275 4031 2309 4058
rect 2005 4024 2037 4031
rect 2077 4024 2105 4031
rect 2149 4024 2173 4031
rect 2221 4024 2241 4031
rect 1861 3997 1899 4024
rect 1933 3997 1971 4024
rect 2005 3997 2043 4024
rect 2077 3997 2115 4024
rect 2149 3997 2187 4024
rect 2221 3997 2259 4024
rect 2293 3997 2309 4031
rect 1799 3987 2309 3997
rect 1799 3955 1833 3987
rect 1867 3955 1901 3987
rect -537 3916 -299 3918
rect -537 3882 -503 3916
rect -469 3882 -435 3916
rect -401 3882 -367 3916
rect -333 3882 -299 3916
rect -537 3878 -299 3882
rect -537 3844 -531 3878
rect -497 3845 -435 3878
rect -401 3845 -339 3878
rect -537 3811 -503 3844
rect -469 3811 -435 3845
rect -401 3811 -367 3845
rect -305 3844 -299 3878
rect -333 3811 -299 3844
rect -537 3807 -299 3811
rect 740 3884 774 3918
rect 808 3884 842 3918
rect 740 3845 842 3884
rect 740 3811 774 3845
rect 808 3811 842 3845
rect 740 3807 842 3811
rect 1799 3921 1827 3955
rect 1867 3953 1899 3955
rect 1935 3953 1969 3987
rect 2003 3955 2037 3987
rect 2071 3955 2105 3987
rect 2139 3955 2173 3987
rect 2207 3955 2241 3987
rect 2275 3955 2309 3987
rect 2005 3953 2037 3955
rect 2077 3953 2105 3955
rect 2149 3953 2173 3955
rect 2221 3953 2241 3955
rect 1861 3921 1899 3953
rect 1933 3921 1971 3953
rect 2005 3921 2043 3953
rect 2077 3921 2115 3953
rect 2149 3921 2187 3953
rect 2221 3921 2259 3953
rect 2293 3921 2309 3955
rect 1799 3916 2309 3921
rect 1799 3882 1833 3916
rect 1867 3882 1901 3916
rect 1935 3882 1969 3916
rect 2003 3882 2037 3916
rect 2071 3882 2105 3916
rect 2139 3882 2173 3916
rect 2207 3882 2241 3916
rect 2275 3882 2309 3916
rect 1799 3879 2309 3882
rect 1799 3845 1827 3879
rect 1861 3845 1899 3879
rect 1933 3845 1971 3879
rect 2005 3845 2043 3879
rect 2077 3845 2115 3879
rect 2149 3845 2187 3879
rect 2221 3845 2259 3879
rect 2293 3845 2309 3879
rect 1799 3811 1833 3845
rect 1867 3811 1901 3845
rect 1935 3811 1969 3845
rect 2003 3811 2037 3845
rect 2071 3811 2105 3845
rect 2139 3811 2173 3845
rect 2207 3811 2241 3845
rect 2275 3811 2309 3845
rect 1799 3807 2309 3811
rect -537 3803 2309 3807
rect -537 3769 -531 3803
rect -497 3773 -435 3803
rect -401 3773 -339 3803
rect -305 3802 2309 3803
rect -305 3773 1827 3802
rect 1861 3773 1899 3802
rect 1933 3773 1971 3802
rect 2005 3773 2043 3802
rect 2077 3773 2115 3802
rect 2149 3773 2187 3802
rect 2221 3773 2259 3802
rect -537 3728 -503 3769
rect 619 3739 654 3773
rect 688 3739 723 3773
rect 757 3739 792 3773
rect 826 3739 861 3773
rect 895 3739 930 3773
rect 964 3739 999 3773
rect 1033 3739 1068 3773
rect 1102 3739 1137 3773
rect 1171 3739 1206 3773
rect 1240 3739 1275 3773
rect 1309 3739 1344 3773
rect 1378 3739 1413 3773
rect 1447 3739 1482 3773
rect 1516 3739 1551 3773
rect 1585 3739 1620 3773
rect 1654 3739 1689 3773
rect 1723 3739 1758 3773
rect 1792 3739 1827 3773
rect 1861 3739 1896 3773
rect 1933 3768 1965 3773
rect 2005 3768 2034 3773
rect 2077 3768 2103 3773
rect 2149 3768 2172 3773
rect 2221 3768 2241 3773
rect 2293 3768 2309 3802
rect 1930 3739 1965 3768
rect 1999 3739 2034 3768
rect 2068 3739 2103 3768
rect 2137 3739 2172 3768
rect 2206 3739 2241 3768
rect 2275 3739 2309 3768
rect -537 3694 -531 3728
rect 619 3720 2309 3739
rect -537 3671 -503 3694
rect 619 3686 638 3720
rect 672 3705 711 3720
rect 745 3705 784 3720
rect 818 3705 857 3720
rect 891 3705 930 3720
rect 964 3705 1003 3720
rect 1037 3705 1076 3720
rect 1110 3705 1149 3720
rect 1183 3705 1222 3720
rect 1256 3705 1295 3720
rect 1329 3705 1368 3720
rect 1402 3705 1441 3720
rect 1475 3705 1514 3720
rect 1548 3705 1587 3720
rect 1621 3705 1660 3720
rect 1694 3705 1733 3720
rect 2271 3705 2309 3720
rect 688 3686 711 3705
rect 757 3686 784 3705
rect 826 3686 857 3705
rect 619 3671 654 3686
rect 688 3671 723 3686
rect 757 3671 792 3686
rect 826 3671 861 3686
rect 895 3671 930 3705
rect 964 3671 999 3705
rect 1037 3686 1068 3705
rect 1110 3686 1137 3705
rect 1183 3686 1206 3705
rect 1256 3686 1275 3705
rect 1329 3686 1344 3705
rect 1402 3686 1413 3705
rect 1475 3686 1482 3705
rect 1548 3686 1551 3705
rect 1033 3671 1068 3686
rect 1102 3671 1137 3686
rect 1171 3671 1206 3686
rect 1240 3671 1275 3686
rect 1309 3671 1344 3686
rect 1378 3671 1413 3686
rect 1447 3671 1482 3686
rect 1516 3671 1551 3686
rect 1585 3686 1587 3705
rect 1654 3686 1660 3705
rect 1585 3671 1620 3686
rect 1654 3671 1689 3686
rect 1723 3671 1733 3705
rect 2275 3671 2309 3705
rect -537 3653 1733 3671
rect -537 3619 -531 3653
rect -497 3619 -435 3653
rect -401 3619 -339 3653
rect -305 3648 1733 3653
rect -305 3619 -238 3648
rect -537 3614 -238 3619
rect -204 3614 -165 3648
rect -131 3614 -92 3648
rect -58 3614 -19 3648
rect 15 3614 54 3648
rect 88 3614 127 3648
rect 161 3614 200 3648
rect 234 3614 273 3648
rect 307 3614 346 3648
rect 380 3614 419 3648
rect 453 3614 492 3648
rect 526 3614 565 3648
rect 599 3614 638 3648
rect 672 3614 711 3648
rect 745 3614 784 3648
rect 818 3614 857 3648
rect 891 3614 930 3648
rect 964 3614 1003 3648
rect 1037 3614 1076 3648
rect 1110 3614 1149 3648
rect 1183 3614 1222 3648
rect 1256 3614 1295 3648
rect 1329 3614 1368 3648
rect 1402 3614 1441 3648
rect 1475 3614 1514 3648
rect 1548 3614 1587 3648
rect 1621 3614 1660 3648
rect 1694 3614 1733 3648
rect -537 3576 1733 3614
rect -537 3542 -238 3576
rect -204 3542 -165 3576
rect -131 3542 -92 3576
rect -58 3542 -19 3576
rect 15 3542 54 3576
rect 88 3542 127 3576
rect 161 3542 200 3576
rect 234 3542 273 3576
rect 307 3542 346 3576
rect 380 3542 419 3576
rect 453 3542 492 3576
rect 526 3542 565 3576
rect 599 3542 638 3576
rect 672 3542 711 3576
rect 745 3542 784 3576
rect 818 3542 857 3576
rect 891 3542 930 3576
rect 964 3542 1003 3576
rect 1037 3542 1076 3576
rect 1110 3542 1149 3576
rect 1183 3542 1222 3576
rect 1256 3542 1295 3576
rect 1329 3542 1368 3576
rect 1402 3542 1441 3576
rect 1475 3542 1514 3576
rect 1548 3542 1587 3576
rect 1621 3542 1660 3576
rect 1694 3542 1733 3576
rect 2271 3637 2309 3671
rect 2753 1071 2787 1095
rect 2753 999 2787 1037
rect 2394 934 2428 950
rect 2547 947 2585 981
rect 2394 866 2428 900
rect 2394 816 2428 828
rect 2753 927 2787 965
rect 2753 855 2787 893
rect 2528 772 2629 806
rect 2753 783 2787 821
rect 2753 711 2787 749
rect 170 666 186 700
rect 220 666 260 700
rect 294 666 334 700
rect 368 666 408 700
rect 442 666 482 700
rect 516 666 555 700
rect 589 666 628 700
rect 662 666 701 700
rect 735 666 742 700
rect 808 666 833 700
rect 881 666 920 700
rect 958 666 970 700
rect 1026 666 1038 700
rect 1076 666 1111 700
rect 1146 666 1182 700
rect 1218 666 1252 700
rect 1291 666 1322 700
rect 1364 666 1392 700
rect 1437 666 1462 700
rect 1510 666 1532 700
rect 1583 666 1602 700
rect 1656 666 1672 700
rect 1729 666 1742 700
rect 1802 666 1812 700
rect 1875 666 1882 700
rect 1948 666 1952 700
rect 1986 666 1987 700
rect 2021 666 2022 700
rect 2056 666 2060 700
rect 2126 666 2132 700
rect 2196 666 2204 700
rect 2265 666 2276 700
rect 2334 666 2369 700
rect 2403 666 2438 700
rect 2472 666 2507 700
rect 2541 666 2576 700
rect 2610 666 2626 700
rect 2753 638 2787 677
rect 2748 604 2753 616
rect 125 509 159 547
rect 2637 532 2671 570
rect 2637 460 2671 498
rect 2748 582 2756 604
rect 2790 582 2798 616
rect 2748 565 2798 582
rect 2748 531 2753 565
rect 2787 543 2798 565
rect 2748 509 2756 531
rect 2790 509 2798 543
rect 2748 492 2798 509
rect 2748 458 2753 492
rect 2787 470 2798 492
rect 2748 436 2756 458
rect 2790 436 2798 470
rect 2748 419 2798 436
rect 2748 385 2753 419
rect 2787 397 2798 419
rect 2748 363 2756 385
rect 2790 363 2798 397
rect 2748 346 2798 363
rect 170 294 186 328
rect 220 294 260 328
rect 328 294 334 328
rect 368 294 385 328
rect 442 294 476 328
rect 516 294 555 328
rect 589 294 628 328
rect 662 294 701 328
rect 735 294 774 328
rect 808 294 847 328
rect 881 294 920 328
rect 954 294 970 328
rect 1026 294 1038 328
rect 1076 294 1112 328
rect 1146 294 1182 328
rect 1220 294 1252 328
rect 1294 294 1322 328
rect 1368 294 1392 328
rect 1441 294 1462 328
rect 1514 294 1532 328
rect 1587 294 1602 328
rect 1660 294 1672 328
rect 1706 294 1742 328
rect 1776 294 1812 328
rect 1846 294 1882 328
rect 1916 294 1952 328
rect 1986 294 2022 328
rect 2056 294 2092 328
rect 2126 294 2162 328
rect 2196 294 2231 328
rect 2265 294 2300 328
rect 2334 294 2369 328
rect 2403 294 2438 328
rect 2472 294 2507 328
rect 2541 294 2576 328
rect 2610 294 2626 328
rect 2748 312 2753 346
rect 2787 324 2798 346
rect 2748 290 2756 312
rect 2790 290 2798 324
rect 2748 273 2798 290
rect 2748 239 2753 273
rect 2787 251 2798 273
rect 76 158 114 192
rect 2637 162 2671 200
rect 2637 90 2671 128
rect 2748 217 2756 239
rect 2790 217 2798 251
rect 2748 200 2798 217
rect 2748 166 2753 200
rect 2787 177 2798 200
rect 2748 143 2756 166
rect 2790 143 2798 177
rect 2748 127 2798 143
rect 2748 93 2753 127
rect 2787 103 2798 127
rect 2748 69 2756 93
rect 2790 69 2798 103
rect 2002 -70 2053 -68
rect 2087 -70 2138 -68
rect 2172 -70 2223 -68
rect 2257 -70 2308 -68
rect 1956 -102 1968 -70
rect 2006 -102 2053 -70
rect 2090 -102 2138 -70
rect 1956 -104 1972 -102
rect 2006 -104 2056 -102
rect 2090 -104 2140 -102
rect 2174 -104 2223 -70
rect 2257 -104 2306 -70
rect 2342 -102 2356 -70
rect 2340 -104 2356 -102
rect 928 -238 962 -226
rect 1052 -229 1098 -195
rect 1132 -229 1178 -195
rect 1212 -229 1259 -195
rect 1293 -229 1340 -195
rect 1374 -229 1421 -195
rect 1455 -229 1502 -195
rect 2368 -198 2406 -164
rect 928 -310 962 -276
rect 1911 -305 1945 -211
rect 928 -360 962 -344
rect 1052 -405 1096 -371
rect 1130 -405 1174 -371
rect 1208 -405 1252 -371
rect 1286 -405 1330 -371
rect 1364 -405 1408 -371
rect 1442 -405 1486 -371
rect 1520 -405 1564 -371
rect 928 -428 962 -416
rect 928 -500 962 -466
rect 1956 -476 1967 -442
rect 2027 -476 2040 -442
rect 2098 -476 2113 -442
rect 2169 -476 2186 -442
rect 2240 -476 2258 -442
rect 2310 -476 2330 -442
rect 2380 -476 2402 -442
rect 2450 -476 2474 -442
rect 2520 -476 2546 -442
rect 2590 -476 2618 -442
rect 2660 -476 2690 -442
rect 928 -550 962 -534
rect 1052 -581 1095 -547
rect 1129 -581 1172 -547
rect 1206 -581 1249 -547
rect 1283 -581 1326 -547
rect 1360 -581 1403 -547
rect 1437 -581 1480 -547
rect 1514 -581 1557 -547
rect 1895 -565 1941 -531
rect 2306 -606 2362 -519
rect 2559 -531 2781 -520
rect 2559 -565 2576 -531
rect 2610 -565 2648 -531
rect 2682 -565 2781 -531
rect 2559 -586 2781 -565
rect 2292 -640 2330 -606
<< viali >>
rect 242 5821 276 5855
rect 316 5821 350 5855
rect 390 5821 424 5855
rect 464 5821 498 5855
rect 538 5821 572 5855
rect 612 5821 646 5855
rect 686 5821 720 5855
rect 760 5821 794 5855
rect 834 5821 868 5855
rect 908 5821 942 5855
rect 982 5821 1016 5855
rect 1056 5821 1090 5855
rect 1130 5821 1164 5855
rect 1204 5821 1238 5855
rect 1278 5821 1312 5855
rect 1352 5821 1386 5855
rect 1426 5821 1460 5855
rect 1500 5821 1534 5855
rect 1574 5821 1608 5855
rect 1648 5821 1682 5855
rect 1722 5821 1756 5855
rect 1796 5821 1830 5855
rect 1870 5821 1904 5855
rect 1944 5821 1978 5855
rect 2018 5821 2052 5855
rect 2091 5821 2125 5855
rect 2164 5821 2198 5855
rect 2237 5821 2271 5855
rect -531 5780 -503 5802
rect -503 5780 -497 5802
rect -435 5780 -401 5802
rect -339 5780 -333 5802
rect -333 5780 -305 5802
rect -531 5768 -497 5780
rect -435 5768 -401 5780
rect -339 5768 -305 5780
rect 242 5746 276 5772
rect 316 5746 350 5772
rect 390 5746 424 5772
rect 464 5746 498 5772
rect 538 5746 572 5772
rect 612 5746 646 5772
rect 686 5746 720 5772
rect 760 5746 794 5772
rect 834 5746 868 5772
rect 908 5746 942 5772
rect 982 5746 1016 5772
rect 1056 5746 1090 5772
rect 1130 5746 1164 5772
rect 1204 5746 1238 5772
rect 1278 5746 1312 5772
rect 1352 5746 1386 5772
rect 1426 5746 1460 5772
rect 1500 5746 1534 5772
rect 1574 5746 1608 5772
rect 1648 5746 1682 5772
rect 1722 5746 1756 5772
rect -531 5710 -503 5728
rect -503 5710 -497 5728
rect -435 5710 -401 5728
rect -339 5710 -333 5728
rect -333 5710 -305 5728
rect 242 5738 254 5746
rect 254 5738 276 5746
rect 316 5738 323 5746
rect 323 5738 350 5746
rect 390 5738 392 5746
rect 392 5738 424 5746
rect 464 5738 496 5746
rect 496 5738 498 5746
rect 538 5738 565 5746
rect 565 5738 572 5746
rect 612 5738 634 5746
rect 634 5738 646 5746
rect 686 5738 703 5746
rect 703 5738 720 5746
rect 760 5738 772 5746
rect 772 5738 794 5746
rect 834 5738 841 5746
rect 841 5738 868 5746
rect 908 5738 910 5746
rect 910 5738 942 5746
rect 982 5738 1013 5746
rect 1013 5738 1016 5746
rect 1056 5738 1082 5746
rect 1082 5738 1090 5746
rect 1130 5738 1151 5746
rect 1151 5738 1164 5746
rect 1204 5738 1220 5746
rect 1220 5738 1238 5746
rect 1278 5738 1289 5746
rect 1289 5738 1312 5746
rect 1352 5738 1358 5746
rect 1358 5738 1386 5746
rect 1426 5738 1427 5746
rect 1427 5738 1460 5746
rect 1500 5738 1531 5746
rect 1531 5738 1534 5746
rect 1574 5738 1600 5746
rect 1600 5738 1608 5746
rect 1648 5738 1669 5746
rect 1669 5738 1682 5746
rect 1722 5738 1738 5746
rect 1738 5738 1756 5746
rect 1796 5738 1807 5772
rect 1807 5738 1830 5772
rect 1870 5738 1904 5772
rect 1944 5738 1977 5772
rect 1977 5738 1978 5772
rect 2018 5768 2037 5772
rect 2037 5768 2052 5772
rect 2091 5768 2105 5772
rect 2105 5768 2125 5772
rect 2164 5768 2173 5772
rect 2173 5768 2198 5772
rect 2237 5768 2241 5772
rect 2241 5768 2271 5772
rect 2018 5738 2052 5768
rect 2091 5738 2125 5768
rect 2164 5738 2198 5768
rect 2237 5738 2271 5768
rect -531 5694 -497 5710
rect -435 5694 -401 5710
rect -339 5694 -305 5710
rect 242 5678 276 5689
rect 316 5678 350 5689
rect 390 5678 424 5689
rect 464 5678 498 5689
rect 538 5678 572 5689
rect 612 5678 646 5689
rect 686 5678 720 5689
rect 760 5678 794 5689
rect 834 5678 868 5689
rect 908 5678 942 5689
rect 982 5678 1016 5689
rect 1056 5678 1090 5689
rect 1130 5678 1164 5689
rect 1204 5678 1238 5689
rect 1278 5678 1312 5689
rect 1352 5678 1386 5689
rect 1426 5678 1460 5689
rect 1500 5678 1534 5689
rect 1574 5678 1608 5689
rect 1648 5678 1682 5689
rect 1722 5678 1756 5689
rect -531 5640 -503 5654
rect -503 5640 -497 5654
rect -435 5640 -401 5654
rect -339 5640 -333 5654
rect -333 5640 -305 5654
rect 242 5655 254 5678
rect 254 5655 276 5678
rect 316 5655 323 5678
rect 323 5655 350 5678
rect 390 5655 392 5678
rect 392 5655 424 5678
rect 464 5655 496 5678
rect 496 5655 498 5678
rect 538 5655 565 5678
rect 565 5655 572 5678
rect 612 5655 634 5678
rect 634 5655 646 5678
rect 686 5655 703 5678
rect 703 5655 720 5678
rect 760 5655 772 5678
rect 772 5655 794 5678
rect 834 5655 841 5678
rect 841 5655 868 5678
rect 908 5655 910 5678
rect 910 5655 942 5678
rect 982 5655 1013 5678
rect 1013 5655 1016 5678
rect 1056 5655 1082 5678
rect 1082 5655 1090 5678
rect 1130 5655 1151 5678
rect 1151 5655 1164 5678
rect 1204 5655 1220 5678
rect 1220 5655 1238 5678
rect 1278 5655 1289 5678
rect 1289 5655 1312 5678
rect 1352 5655 1358 5678
rect 1358 5655 1386 5678
rect 1426 5655 1427 5678
rect 1427 5655 1460 5678
rect 1500 5655 1531 5678
rect 1531 5655 1534 5678
rect 1574 5655 1600 5678
rect 1600 5655 1608 5678
rect 1648 5655 1669 5678
rect 1669 5655 1682 5678
rect 1722 5655 1738 5678
rect 1738 5655 1756 5678
rect 1796 5655 1807 5689
rect 1807 5655 1830 5689
rect 1870 5655 1904 5689
rect 1944 5655 1977 5689
rect 1977 5655 1978 5689
rect 2018 5660 2052 5689
rect 2091 5660 2125 5689
rect 2164 5660 2198 5689
rect 2237 5660 2271 5689
rect 2018 5655 2037 5660
rect 2037 5655 2052 5660
rect 2091 5655 2105 5660
rect 2105 5655 2125 5660
rect 2164 5655 2173 5660
rect 2173 5655 2198 5660
rect 2237 5655 2241 5660
rect 2241 5655 2271 5660
rect -531 5620 -497 5640
rect -435 5620 -401 5640
rect -339 5620 -305 5640
rect -531 5570 -503 5580
rect -503 5570 -497 5580
rect -435 5570 -401 5580
rect -339 5570 -333 5580
rect -333 5570 -305 5580
rect -531 5546 -497 5570
rect -435 5546 -401 5570
rect -339 5546 -305 5570
rect -531 5500 -503 5506
rect -503 5500 -497 5506
rect -435 5500 -401 5506
rect 1970 5543 2004 5577
rect 2042 5555 2071 5577
rect 2071 5555 2076 5577
rect 2114 5555 2139 5577
rect 2139 5555 2148 5577
rect 2186 5555 2207 5577
rect 2207 5555 2220 5577
rect 2258 5555 2275 5577
rect 2275 5555 2292 5577
rect 2042 5543 2076 5555
rect 2114 5543 2148 5555
rect 2186 5543 2220 5555
rect 2258 5543 2292 5555
rect 73 5516 107 5517
rect 156 5516 190 5517
rect 238 5516 272 5517
rect 408 5516 442 5517
rect 527 5516 561 5517
rect 864 5516 898 5517
rect 947 5516 981 5517
rect 1029 5516 1063 5517
rect 1445 5516 1479 5517
rect 1528 5516 1562 5517
rect 1610 5516 1644 5517
rect -339 5500 -333 5506
rect -333 5500 -305 5506
rect -531 5472 -497 5500
rect -435 5472 -401 5500
rect -339 5472 -305 5500
rect 73 5483 78 5516
rect 78 5483 107 5516
rect 156 5483 190 5516
rect 238 5483 268 5516
rect 268 5483 272 5516
rect 408 5483 434 5516
rect 434 5483 442 5516
rect 527 5483 546 5516
rect 546 5483 561 5516
rect 864 5483 868 5516
rect 868 5483 898 5516
rect 947 5483 980 5516
rect 980 5483 981 5516
rect 1029 5483 1058 5516
rect 1058 5483 1063 5516
rect 1445 5483 1458 5516
rect 1458 5483 1479 5516
rect 1528 5483 1536 5516
rect 1536 5483 1562 5516
rect 1610 5483 1614 5516
rect 1614 5483 1644 5516
rect -531 5430 -503 5432
rect -503 5430 -497 5432
rect -435 5430 -401 5432
rect -339 5430 -333 5432
rect -333 5430 -305 5432
rect -531 5398 -497 5430
rect -435 5398 -401 5430
rect -339 5398 -305 5430
rect 1970 5469 2004 5503
rect 2042 5484 2071 5503
rect 2071 5484 2076 5503
rect 2114 5484 2139 5503
rect 2139 5484 2148 5503
rect 2186 5484 2207 5503
rect 2207 5484 2220 5503
rect 2258 5484 2275 5503
rect 2275 5484 2292 5503
rect 2042 5469 2076 5484
rect 2114 5469 2148 5484
rect 2186 5469 2220 5484
rect 2258 5469 2292 5484
rect -531 5324 -497 5358
rect -435 5324 -401 5358
rect -339 5324 -305 5358
rect 39 5392 73 5426
rect -531 5254 -497 5284
rect -435 5254 -401 5284
rect -339 5254 -305 5284
rect -531 5250 -503 5254
rect -503 5250 -497 5254
rect -435 5250 -401 5254
rect -339 5250 -333 5254
rect -333 5250 -305 5254
rect -531 5184 -497 5210
rect -435 5184 -401 5210
rect -339 5184 -305 5210
rect -531 5176 -503 5184
rect -503 5176 -497 5184
rect -435 5176 -401 5184
rect -339 5176 -333 5184
rect -333 5176 -305 5184
rect -531 5114 -497 5136
rect -435 5114 -401 5136
rect -339 5114 -305 5136
rect -531 5102 -503 5114
rect -503 5102 -497 5114
rect -435 5102 -401 5114
rect -339 5102 -333 5114
rect -333 5102 -305 5114
rect -531 5044 -497 5062
rect -435 5044 -401 5062
rect -339 5044 -305 5062
rect -531 5028 -503 5044
rect -503 5028 -497 5044
rect -435 5028 -401 5044
rect -339 5028 -333 5044
rect -333 5028 -305 5044
rect -531 4974 -497 4988
rect -435 4974 -401 4988
rect -339 4974 -305 4988
rect -531 4954 -503 4974
rect -503 4954 -497 4974
rect -435 4954 -401 4974
rect -339 4954 -333 4974
rect -333 4954 -305 4974
rect -531 4904 -497 4914
rect -435 4904 -401 4914
rect -339 4904 -305 4914
rect -531 4880 -503 4904
rect -503 4880 -497 4904
rect -435 4880 -401 4904
rect -339 4880 -333 4904
rect -333 4880 -305 4904
rect -217 5272 -183 5306
rect -217 5187 -183 5221
rect -217 5102 -183 5136
rect 39 5300 73 5334
rect 551 5392 585 5426
rect 551 5315 585 5349
rect 39 5207 73 5241
rect 39 5114 73 5148
rect 295 5272 329 5306
rect 295 5187 329 5221
rect -217 5017 -183 5051
rect -217 4932 -183 4966
rect -217 4846 -183 4880
rect 295 5102 329 5136
rect 295 5017 329 5051
rect 551 5237 585 5271
rect 1063 5392 1097 5426
rect 1063 5315 1097 5349
rect 1575 5392 1609 5426
rect 1575 5315 1609 5349
rect 551 5159 585 5193
rect 551 5081 585 5115
rect 551 5003 585 5037
rect 807 5205 841 5239
rect 807 5116 841 5150
rect 807 5026 841 5060
rect 295 4932 329 4966
rect 295 4846 329 4880
rect 1063 5237 1097 5271
rect 1063 5159 1097 5193
rect 1063 5081 1097 5115
rect 1063 5003 1097 5037
rect 1319 5272 1353 5306
rect 1319 5187 1353 5221
rect 1319 5102 1353 5136
rect 1319 5017 1353 5051
rect 807 4936 841 4970
rect 807 4846 841 4880
rect 1575 5237 1609 5271
rect 1970 5394 2004 5428
rect 2042 5412 2071 5428
rect 2071 5412 2076 5428
rect 2114 5412 2139 5428
rect 2139 5412 2148 5428
rect 2186 5412 2207 5428
rect 2207 5412 2220 5428
rect 2258 5412 2275 5428
rect 2275 5412 2292 5428
rect 2042 5394 2076 5412
rect 2114 5394 2148 5412
rect 2186 5394 2220 5412
rect 2258 5394 2292 5412
rect 1970 5319 2004 5353
rect 2042 5340 2071 5353
rect 2071 5340 2076 5353
rect 2114 5340 2139 5353
rect 2139 5340 2148 5353
rect 2186 5340 2207 5353
rect 2207 5340 2220 5353
rect 2258 5340 2275 5353
rect 2275 5340 2292 5353
rect 2042 5319 2076 5340
rect 2114 5319 2148 5340
rect 2186 5319 2220 5340
rect 2258 5319 2292 5340
rect 1575 5159 1609 5193
rect 1575 5081 1609 5115
rect 1575 5003 1609 5037
rect 1831 5215 1865 5249
rect 1831 5142 1865 5176
rect 1831 5068 1865 5102
rect 1319 4932 1353 4966
rect 1319 4846 1353 4880
rect 1831 4994 1865 5028
rect 1831 4920 1865 4954
rect 1831 4846 1865 4880
rect 1970 5244 2004 5278
rect 2042 5268 2071 5278
rect 2071 5268 2076 5278
rect 2114 5268 2139 5278
rect 2139 5268 2148 5278
rect 2186 5268 2207 5278
rect 2207 5268 2220 5278
rect 2258 5268 2275 5278
rect 2275 5268 2292 5278
rect 2042 5244 2076 5268
rect 2114 5244 2148 5268
rect 2186 5244 2220 5268
rect 2258 5244 2292 5268
rect 1970 5169 2004 5203
rect 2042 5196 2071 5203
rect 2071 5196 2076 5203
rect 2114 5196 2139 5203
rect 2139 5196 2148 5203
rect 2186 5196 2207 5203
rect 2207 5196 2220 5203
rect 2258 5196 2275 5203
rect 2275 5196 2292 5203
rect 2042 5169 2076 5196
rect 2114 5169 2148 5196
rect 2186 5169 2220 5196
rect 2258 5169 2292 5196
rect 1970 5094 2004 5128
rect 2042 5124 2071 5128
rect 2071 5124 2076 5128
rect 2114 5124 2139 5128
rect 2139 5124 2148 5128
rect 2186 5124 2207 5128
rect 2207 5124 2220 5128
rect 2258 5124 2275 5128
rect 2275 5124 2292 5128
rect 2042 5094 2076 5124
rect 2114 5094 2148 5124
rect 2186 5094 2220 5124
rect 2258 5094 2292 5124
rect 1970 5019 2004 5053
rect 2042 5052 2071 5053
rect 2071 5052 2076 5053
rect 2114 5052 2139 5053
rect 2139 5052 2148 5053
rect 2186 5052 2207 5053
rect 2207 5052 2220 5053
rect 2258 5052 2275 5053
rect 2275 5052 2292 5053
rect 2042 5019 2076 5052
rect 2114 5019 2148 5052
rect 2186 5019 2220 5052
rect 2258 5019 2292 5052
rect 1970 4944 2004 4978
rect 2042 4944 2076 4978
rect 2114 4944 2148 4978
rect 2186 4944 2220 4978
rect 2258 4944 2292 4978
rect 1970 4869 2004 4903
rect 2042 4870 2076 4903
rect 2114 4870 2148 4903
rect 2186 4870 2220 4903
rect 2258 4870 2292 4903
rect 2042 4869 2071 4870
rect 2071 4869 2076 4870
rect 2114 4869 2139 4870
rect 2139 4869 2148 4870
rect 2186 4869 2207 4870
rect 2207 4869 2220 4870
rect 2258 4869 2275 4870
rect 2275 4869 2292 4870
rect -531 4834 -497 4840
rect -435 4834 -401 4840
rect -339 4834 -305 4840
rect -531 4806 -503 4834
rect -503 4806 -497 4834
rect -435 4806 -401 4834
rect -339 4806 -333 4834
rect -333 4806 -305 4834
rect -531 4764 -497 4766
rect -435 4764 -401 4766
rect -339 4764 -305 4766
rect -531 4732 -503 4764
rect -503 4732 -497 4764
rect -435 4732 -401 4764
rect -339 4732 -333 4764
rect -333 4732 -305 4764
rect 1970 4794 2004 4828
rect 2042 4798 2076 4828
rect 2114 4798 2148 4828
rect 2186 4798 2220 4828
rect 2258 4798 2292 4828
rect 2042 4794 2071 4798
rect 2071 4794 2076 4798
rect 2114 4794 2139 4798
rect 2139 4794 2148 4798
rect 2186 4794 2207 4798
rect 2207 4794 2220 4798
rect 2258 4794 2275 4798
rect 2275 4794 2292 4798
rect -198 4726 -164 4729
rect -125 4726 -91 4729
rect -52 4726 -18 4729
rect 21 4726 55 4729
rect 94 4726 128 4729
rect 167 4726 201 4729
rect 240 4726 274 4729
rect 312 4726 346 4729
rect 384 4726 418 4729
rect 456 4726 490 4729
rect -531 4660 -503 4692
rect -503 4660 -497 4692
rect -435 4660 -401 4692
rect -198 4695 -196 4726
rect -196 4695 -164 4726
rect -125 4695 -93 4726
rect -93 4695 -91 4726
rect -52 4695 -24 4726
rect -24 4695 -18 4726
rect 21 4695 45 4726
rect 45 4695 55 4726
rect 94 4695 114 4726
rect 114 4695 128 4726
rect 167 4695 183 4726
rect 183 4695 201 4726
rect 240 4695 252 4726
rect 252 4695 274 4726
rect 312 4695 321 4726
rect 321 4695 346 4726
rect 384 4695 390 4726
rect 390 4695 418 4726
rect 456 4695 459 4726
rect 459 4695 490 4726
rect 528 4695 562 4729
rect 600 4726 634 4729
rect 672 4726 706 4729
rect 744 4726 778 4729
rect 816 4726 850 4729
rect 888 4726 922 4729
rect 960 4726 994 4729
rect 1032 4726 1066 4729
rect 1104 4726 1138 4729
rect 1176 4726 1210 4729
rect 1248 4726 1282 4729
rect 1320 4726 1354 4729
rect 1392 4726 1426 4729
rect 1464 4726 1498 4729
rect 1536 4726 1570 4729
rect 1608 4726 1642 4729
rect 1680 4726 1714 4729
rect 1752 4726 1786 4729
rect 1824 4726 1858 4729
rect 1896 4726 1930 4729
rect 1968 4726 2002 4729
rect 2040 4726 2074 4729
rect 600 4695 632 4726
rect 632 4695 634 4726
rect 672 4695 701 4726
rect 701 4695 706 4726
rect 744 4695 770 4726
rect 770 4695 778 4726
rect 816 4695 839 4726
rect 839 4695 850 4726
rect 888 4695 908 4726
rect 908 4695 922 4726
rect 960 4695 977 4726
rect 977 4695 994 4726
rect 1032 4695 1046 4726
rect 1046 4695 1066 4726
rect 1104 4695 1115 4726
rect 1115 4695 1138 4726
rect 1176 4695 1184 4726
rect 1184 4695 1210 4726
rect 1248 4695 1254 4726
rect 1254 4695 1282 4726
rect 1320 4695 1324 4726
rect 1324 4695 1354 4726
rect 1392 4695 1394 4726
rect 1394 4695 1426 4726
rect 1464 4695 1498 4726
rect 1536 4695 1568 4726
rect 1568 4695 1570 4726
rect 1608 4695 1638 4726
rect 1638 4695 1642 4726
rect 1680 4695 1708 4726
rect 1708 4695 1714 4726
rect 1752 4695 1778 4726
rect 1778 4695 1786 4726
rect 1824 4695 1848 4726
rect 1848 4695 1858 4726
rect 1896 4695 1918 4726
rect 1918 4695 1930 4726
rect 1968 4695 1988 4726
rect 1988 4695 2002 4726
rect 2040 4695 2071 4726
rect 2071 4695 2074 4726
rect -339 4660 -333 4692
rect -333 4660 -305 4692
rect -531 4658 -497 4660
rect -435 4658 -401 4660
rect -339 4658 -305 4660
rect -531 4590 -503 4618
rect -503 4590 -497 4618
rect -435 4590 -401 4618
rect -339 4590 -333 4618
rect -333 4590 -305 4618
rect -531 4584 -497 4590
rect -435 4584 -401 4590
rect -339 4584 -305 4590
rect -531 4520 -503 4544
rect -503 4520 -497 4544
rect -435 4520 -401 4544
rect -339 4520 -333 4544
rect -333 4520 -305 4544
rect -531 4510 -497 4520
rect -435 4510 -401 4520
rect -339 4510 -305 4520
rect 405 4559 439 4593
rect -531 4450 -503 4470
rect -503 4450 -497 4470
rect -435 4450 -401 4470
rect -339 4450 -333 4470
rect -333 4450 -305 4470
rect -531 4436 -497 4450
rect -435 4436 -401 4450
rect -339 4436 -305 4450
rect -531 4379 -503 4396
rect -503 4379 -497 4396
rect -435 4379 -401 4396
rect 229 4479 263 4513
rect 405 4487 439 4521
rect 581 4559 615 4593
rect 581 4487 615 4521
rect 1174 4516 1178 4550
rect 1178 4516 1208 4550
rect 1248 4516 1255 4550
rect 1255 4516 1282 4550
rect 1322 4516 1332 4550
rect 1332 4516 1356 4550
rect 1526 4516 1530 4550
rect 1530 4516 1560 4550
rect 1598 4516 1632 4550
rect 1827 4554 1861 4563
rect 1899 4554 1933 4563
rect 1971 4554 2005 4563
rect 2043 4554 2077 4563
rect 2115 4554 2149 4563
rect 2187 4554 2221 4563
rect 2259 4554 2293 4563
rect 1827 4529 1833 4554
rect 1833 4529 1861 4554
rect 1899 4529 1901 4554
rect 1901 4529 1933 4554
rect 1971 4529 2003 4554
rect 2003 4529 2005 4554
rect 2043 4529 2071 4554
rect 2071 4529 2077 4554
rect 2115 4529 2139 4554
rect 2139 4529 2149 4554
rect 2187 4529 2207 4554
rect 2207 4529 2221 4554
rect 2259 4529 2275 4554
rect 2275 4529 2293 4554
rect 229 4407 263 4441
rect -339 4379 -333 4396
rect -333 4379 -305 4396
rect -531 4362 -497 4379
rect -435 4362 -401 4379
rect -339 4362 -305 4379
rect -531 4308 -503 4322
rect -503 4308 -497 4322
rect -435 4308 -401 4322
rect 272 4327 276 4361
rect 276 4327 306 4361
rect 344 4327 378 4361
rect 462 4327 466 4361
rect 466 4327 496 4361
rect 534 4327 568 4361
rect -339 4308 -333 4322
rect -333 4308 -305 4322
rect -531 4288 -497 4308
rect -435 4288 -401 4308
rect -339 4288 -305 4308
rect -531 4237 -503 4248
rect -503 4237 -497 4248
rect -435 4237 -401 4248
rect -339 4237 -333 4248
rect -333 4237 -305 4248
rect -531 4214 -497 4237
rect -435 4214 -401 4237
rect -339 4214 -305 4237
rect -531 4166 -503 4174
rect -503 4166 -497 4174
rect -435 4166 -401 4174
rect 1827 4484 1861 4487
rect 1899 4484 1933 4487
rect 1971 4484 2005 4487
rect 2043 4484 2077 4487
rect 2115 4484 2149 4487
rect 2187 4484 2221 4487
rect 2259 4484 2293 4487
rect 1827 4453 1833 4484
rect 1833 4453 1861 4484
rect 1899 4453 1901 4484
rect 1901 4453 1933 4484
rect 1971 4453 2003 4484
rect 2003 4453 2005 4484
rect 2043 4453 2071 4484
rect 2071 4453 2077 4484
rect 2115 4453 2139 4484
rect 2139 4453 2149 4484
rect 2187 4453 2207 4484
rect 2207 4453 2221 4484
rect 2259 4453 2275 4484
rect 2275 4453 2293 4484
rect 1827 4379 1833 4411
rect 1833 4379 1861 4411
rect 1899 4379 1901 4411
rect 1901 4379 1933 4411
rect 1971 4379 2003 4411
rect 2003 4379 2005 4411
rect 2043 4379 2071 4411
rect 2071 4379 2077 4411
rect 2115 4379 2139 4411
rect 2139 4379 2149 4411
rect 2187 4379 2207 4411
rect 2207 4379 2221 4411
rect 2259 4379 2275 4411
rect 2275 4379 2293 4411
rect 1827 4377 1861 4379
rect 1899 4377 1933 4379
rect 1971 4377 2005 4379
rect 2043 4377 2077 4379
rect 2115 4377 2149 4379
rect 2187 4377 2221 4379
rect 2259 4377 2293 4379
rect 1645 4317 1679 4351
rect -339 4166 -333 4174
rect -333 4166 -305 4174
rect -531 4140 -497 4166
rect -435 4140 -401 4166
rect -339 4140 -305 4166
rect 410 4152 444 4186
rect 482 4152 516 4186
rect 1293 4271 1327 4305
rect -531 4095 -503 4100
rect -503 4095 -497 4100
rect -435 4095 -401 4100
rect -339 4095 -333 4100
rect -333 4095 -305 4100
rect -531 4066 -497 4095
rect -435 4066 -401 4095
rect -339 4066 -305 4095
rect -531 4024 -503 4026
rect -503 4024 -497 4026
rect -435 4024 -401 4026
rect -339 4024 -333 4026
rect -333 4024 -305 4026
rect -531 3992 -497 4024
rect -435 3992 -401 4024
rect -339 3992 -305 4024
rect 405 4062 439 4096
rect -531 3918 -497 3952
rect -435 3918 -401 3952
rect -339 3918 -305 3952
rect 229 3990 263 4024
rect 405 3990 439 4024
rect 581 3990 615 4024
rect 229 3918 263 3952
rect 581 3918 615 3952
rect 1117 4149 1151 4183
rect 1117 4046 1151 4080
rect 1293 4172 1327 4206
rect 1645 4236 1679 4270
rect 1293 4072 1327 4106
rect 1469 4149 1503 4183
rect 1117 3942 1151 3976
rect 1469 4046 1503 4080
rect 1645 4154 1679 4188
rect 1645 4072 1679 4106
rect 1827 4308 1833 4335
rect 1833 4308 1861 4335
rect 1899 4308 1901 4335
rect 1901 4308 1933 4335
rect 1971 4308 2003 4335
rect 2003 4308 2005 4335
rect 2043 4308 2071 4335
rect 2071 4308 2077 4335
rect 2115 4308 2139 4335
rect 2139 4308 2149 4335
rect 2187 4308 2207 4335
rect 2207 4308 2221 4335
rect 2259 4308 2275 4335
rect 2275 4308 2293 4335
rect 1827 4301 1861 4308
rect 1899 4301 1933 4308
rect 1971 4301 2005 4308
rect 2043 4301 2077 4308
rect 2115 4301 2149 4308
rect 2187 4301 2221 4308
rect 2259 4301 2293 4308
rect 1827 4237 1833 4259
rect 1833 4237 1861 4259
rect 1899 4237 1901 4259
rect 1901 4237 1933 4259
rect 1971 4237 2003 4259
rect 2003 4237 2005 4259
rect 2043 4237 2071 4259
rect 2071 4237 2077 4259
rect 2115 4237 2139 4259
rect 2139 4237 2149 4259
rect 2187 4237 2207 4259
rect 2207 4237 2221 4259
rect 2259 4237 2275 4259
rect 2275 4237 2293 4259
rect 1827 4225 1861 4237
rect 1899 4225 1933 4237
rect 1971 4225 2005 4237
rect 2043 4225 2077 4237
rect 2115 4225 2149 4237
rect 2187 4225 2221 4237
rect 2259 4225 2293 4237
rect 1827 4166 1833 4183
rect 1833 4166 1861 4183
rect 1899 4166 1901 4183
rect 1901 4166 1933 4183
rect 1971 4166 2003 4183
rect 2003 4166 2005 4183
rect 2043 4166 2071 4183
rect 2071 4166 2077 4183
rect 2115 4166 2139 4183
rect 2139 4166 2149 4183
rect 2187 4166 2207 4183
rect 2207 4166 2221 4183
rect 2259 4166 2275 4183
rect 2275 4166 2293 4183
rect 1827 4149 1861 4166
rect 1899 4149 1933 4166
rect 1971 4149 2005 4166
rect 2043 4149 2077 4166
rect 2115 4149 2149 4166
rect 2187 4149 2221 4166
rect 2259 4149 2293 4166
rect 1827 4095 1833 4107
rect 1833 4095 1861 4107
rect 1899 4095 1901 4107
rect 1901 4095 1933 4107
rect 1971 4095 2003 4107
rect 2003 4095 2005 4107
rect 2043 4095 2071 4107
rect 2071 4095 2077 4107
rect 2115 4095 2139 4107
rect 2139 4095 2149 4107
rect 2187 4095 2207 4107
rect 2207 4095 2221 4107
rect 2259 4095 2275 4107
rect 2275 4095 2293 4107
rect 1827 4073 1861 4095
rect 1899 4073 1933 4095
rect 1971 4073 2005 4095
rect 2043 4073 2077 4095
rect 2115 4073 2149 4095
rect 2187 4073 2221 4095
rect 2259 4073 2293 4095
rect 1469 3942 1503 3976
rect 1827 4024 1833 4031
rect 1833 4024 1861 4031
rect 1899 4024 1901 4031
rect 1901 4024 1933 4031
rect 1971 4024 2003 4031
rect 2003 4024 2005 4031
rect 2043 4024 2071 4031
rect 2071 4024 2077 4031
rect 2115 4024 2139 4031
rect 2139 4024 2149 4031
rect 2187 4024 2207 4031
rect 2207 4024 2221 4031
rect 2259 4024 2275 4031
rect 2275 4024 2293 4031
rect 1827 3997 1861 4024
rect 1899 3997 1933 4024
rect 1971 3997 2005 4024
rect 2043 3997 2077 4024
rect 2115 3997 2149 4024
rect 2187 3997 2221 4024
rect 2259 3997 2293 4024
rect -531 3845 -497 3878
rect -435 3845 -401 3878
rect -339 3845 -305 3878
rect -531 3844 -503 3845
rect -503 3844 -497 3845
rect -435 3844 -401 3845
rect -339 3844 -333 3845
rect -333 3844 -305 3845
rect 1827 3953 1833 3955
rect 1833 3953 1861 3955
rect 1899 3953 1901 3955
rect 1901 3953 1933 3955
rect 1971 3953 2003 3955
rect 2003 3953 2005 3955
rect 2043 3953 2071 3955
rect 2071 3953 2077 3955
rect 2115 3953 2139 3955
rect 2139 3953 2149 3955
rect 2187 3953 2207 3955
rect 2207 3953 2221 3955
rect 2259 3953 2275 3955
rect 2275 3953 2293 3955
rect 1827 3921 1861 3953
rect 1899 3921 1933 3953
rect 1971 3921 2005 3953
rect 2043 3921 2077 3953
rect 2115 3921 2149 3953
rect 2187 3921 2221 3953
rect 2259 3921 2293 3953
rect 1827 3845 1861 3879
rect 1899 3845 1933 3879
rect 1971 3845 2005 3879
rect 2043 3845 2077 3879
rect 2115 3845 2149 3879
rect 2187 3845 2221 3879
rect 2259 3845 2293 3879
rect -531 3773 -497 3803
rect -435 3773 -401 3803
rect -339 3773 -305 3803
rect 1827 3773 1861 3802
rect 1899 3773 1933 3802
rect 1971 3773 2005 3802
rect 2043 3773 2077 3802
rect 2115 3773 2149 3802
rect 2187 3773 2221 3802
rect 2259 3773 2293 3802
rect -531 3769 -503 3773
rect -503 3769 -497 3773
rect -435 3769 -401 3773
rect -339 3769 -305 3773
rect 1827 3768 1861 3773
rect 1899 3768 1930 3773
rect 1930 3768 1933 3773
rect 1971 3768 1999 3773
rect 1999 3768 2005 3773
rect 2043 3768 2068 3773
rect 2068 3768 2077 3773
rect 2115 3768 2137 3773
rect 2137 3768 2149 3773
rect 2187 3768 2206 3773
rect 2206 3768 2221 3773
rect 2259 3768 2275 3773
rect 2275 3768 2293 3773
rect -531 3694 -503 3728
rect -503 3694 -497 3728
rect -435 3694 -401 3728
rect -339 3694 -305 3728
rect -238 3686 -204 3720
rect -165 3686 -131 3720
rect -92 3686 -58 3720
rect -19 3686 15 3720
rect 54 3686 88 3720
rect 127 3686 161 3720
rect 200 3686 234 3720
rect 273 3686 307 3720
rect 346 3686 380 3720
rect 419 3686 453 3720
rect 492 3686 526 3720
rect 565 3686 599 3720
rect 638 3705 672 3720
rect 711 3705 745 3720
rect 784 3705 818 3720
rect 857 3705 891 3720
rect 930 3705 964 3720
rect 1003 3705 1037 3720
rect 1076 3705 1110 3720
rect 1149 3705 1183 3720
rect 1222 3705 1256 3720
rect 1295 3705 1329 3720
rect 1368 3705 1402 3720
rect 1441 3705 1475 3720
rect 1514 3705 1548 3720
rect 1587 3705 1621 3720
rect 1660 3705 1694 3720
rect 1733 3705 2271 3720
rect 638 3686 654 3705
rect 654 3686 672 3705
rect 711 3686 723 3705
rect 723 3686 745 3705
rect 784 3686 792 3705
rect 792 3686 818 3705
rect 857 3686 861 3705
rect 861 3686 891 3705
rect 930 3686 964 3705
rect 1003 3686 1033 3705
rect 1033 3686 1037 3705
rect 1076 3686 1102 3705
rect 1102 3686 1110 3705
rect 1149 3686 1171 3705
rect 1171 3686 1183 3705
rect 1222 3686 1240 3705
rect 1240 3686 1256 3705
rect 1295 3686 1309 3705
rect 1309 3686 1329 3705
rect 1368 3686 1378 3705
rect 1378 3686 1402 3705
rect 1441 3686 1447 3705
rect 1447 3686 1475 3705
rect 1514 3686 1516 3705
rect 1516 3686 1548 3705
rect 1587 3686 1620 3705
rect 1620 3686 1621 3705
rect 1660 3686 1689 3705
rect 1689 3686 1694 3705
rect 1733 3671 1758 3705
rect 1758 3671 1792 3705
rect 1792 3671 1827 3705
rect 1827 3671 1861 3705
rect 1861 3671 1896 3705
rect 1896 3671 1930 3705
rect 1930 3671 1965 3705
rect 1965 3671 1999 3705
rect 1999 3671 2034 3705
rect 2034 3671 2068 3705
rect 2068 3671 2103 3705
rect 2103 3671 2137 3705
rect 2137 3671 2172 3705
rect 2172 3671 2206 3705
rect 2206 3671 2241 3705
rect 2241 3671 2271 3705
rect -531 3619 -497 3653
rect -435 3619 -401 3653
rect -339 3619 -305 3653
rect -238 3614 -204 3648
rect -165 3614 -131 3648
rect -92 3614 -58 3648
rect -19 3614 15 3648
rect 54 3614 88 3648
rect 127 3614 161 3648
rect 200 3614 234 3648
rect 273 3614 307 3648
rect 346 3614 380 3648
rect 419 3614 453 3648
rect 492 3614 526 3648
rect 565 3614 599 3648
rect 638 3614 672 3648
rect 711 3614 745 3648
rect 784 3614 818 3648
rect 857 3614 891 3648
rect 930 3614 964 3648
rect 1003 3614 1037 3648
rect 1076 3614 1110 3648
rect 1149 3614 1183 3648
rect 1222 3614 1256 3648
rect 1295 3614 1329 3648
rect 1368 3614 1402 3648
rect 1441 3614 1475 3648
rect 1514 3614 1548 3648
rect 1587 3614 1621 3648
rect 1660 3614 1694 3648
rect -238 3542 -204 3576
rect -165 3542 -131 3576
rect -92 3542 -58 3576
rect -19 3542 15 3576
rect 54 3542 88 3576
rect 127 3542 161 3576
rect 200 3542 234 3576
rect 273 3542 307 3576
rect 346 3542 380 3576
rect 419 3542 453 3576
rect 492 3542 526 3576
rect 565 3542 599 3576
rect 638 3542 672 3576
rect 711 3542 745 3576
rect 784 3542 818 3576
rect 857 3542 891 3576
rect 930 3542 964 3576
rect 1003 3542 1037 3576
rect 1076 3542 1110 3576
rect 1149 3542 1183 3576
rect 1222 3542 1256 3576
rect 1295 3542 1329 3576
rect 1368 3542 1402 3576
rect 1441 3542 1475 3576
rect 1514 3542 1548 3576
rect 1587 3542 1621 3576
rect 1660 3542 1694 3576
rect 1733 3542 2271 3671
rect 2513 947 2547 981
rect 2585 947 2619 981
rect 2394 900 2428 934
rect 2394 832 2428 862
rect 2394 828 2428 832
rect 2494 772 2528 806
rect 2629 772 2663 806
rect 742 666 774 700
rect 774 666 776 700
rect 833 666 847 700
rect 847 666 867 700
rect 924 666 954 700
rect 954 666 958 700
rect 1038 666 1042 700
rect 1042 666 1072 700
rect 1111 666 1112 700
rect 1112 666 1145 700
rect 1184 666 1216 700
rect 1216 666 1218 700
rect 1257 666 1286 700
rect 1286 666 1291 700
rect 1330 666 1356 700
rect 1356 666 1364 700
rect 1403 666 1426 700
rect 1426 666 1437 700
rect 1476 666 1496 700
rect 1496 666 1510 700
rect 1549 666 1566 700
rect 1566 666 1583 700
rect 1622 666 1636 700
rect 1636 666 1656 700
rect 1695 666 1706 700
rect 1706 666 1729 700
rect 1768 666 1776 700
rect 1776 666 1802 700
rect 1841 666 1846 700
rect 1846 666 1875 700
rect 1914 666 1916 700
rect 1916 666 1948 700
rect 1987 666 2021 700
rect 2060 666 2092 700
rect 2092 666 2094 700
rect 2132 666 2162 700
rect 2162 666 2166 700
rect 2204 666 2231 700
rect 2231 666 2238 700
rect 2276 666 2300 700
rect 2300 666 2310 700
rect 2756 604 2787 616
rect 2787 604 2790 616
rect 125 547 159 581
rect 125 475 159 509
rect 2637 570 2671 604
rect 2637 498 2671 532
rect 2637 426 2671 460
rect 2756 582 2790 604
rect 2756 531 2787 543
rect 2787 531 2790 543
rect 2756 509 2790 531
rect 2756 458 2787 470
rect 2787 458 2790 470
rect 2756 436 2790 458
rect 2756 385 2787 397
rect 2787 385 2790 397
rect 2756 363 2790 385
rect 294 294 328 328
rect 385 294 408 328
rect 408 294 419 328
rect 476 294 482 328
rect 482 294 510 328
rect 1038 294 1042 328
rect 1042 294 1072 328
rect 1112 294 1146 328
rect 1186 294 1216 328
rect 1216 294 1220 328
rect 1260 294 1286 328
rect 1286 294 1294 328
rect 1334 294 1356 328
rect 1356 294 1368 328
rect 1407 294 1426 328
rect 1426 294 1441 328
rect 1480 294 1496 328
rect 1496 294 1514 328
rect 1553 294 1566 328
rect 1566 294 1587 328
rect 1626 294 1636 328
rect 1636 294 1660 328
rect 2756 312 2787 324
rect 2787 312 2790 324
rect 2756 290 2790 312
rect 2756 239 2787 251
rect 2787 239 2790 251
rect 2637 200 2671 234
rect 42 158 76 192
rect 114 158 148 192
rect 2637 128 2671 162
rect 2637 56 2671 90
rect 2756 217 2790 239
rect 2756 166 2787 177
rect 2787 166 2790 177
rect 2756 143 2790 166
rect 2756 93 2787 103
rect 2787 93 2790 103
rect 2756 69 2790 93
rect 1968 -70 2002 -68
rect 2053 -70 2087 -68
rect 2138 -70 2172 -68
rect 2223 -70 2257 -68
rect 2308 -70 2342 -68
rect 1968 -102 1972 -70
rect 1972 -102 2002 -70
rect 2053 -102 2056 -70
rect 2056 -102 2087 -70
rect 2138 -102 2140 -70
rect 2140 -102 2172 -70
rect 2223 -102 2257 -70
rect 2308 -102 2340 -70
rect 2340 -102 2342 -70
rect 1018 -229 1052 -195
rect 1098 -229 1132 -195
rect 1178 -229 1212 -195
rect 1259 -229 1293 -195
rect 1340 -229 1374 -195
rect 1421 -229 1455 -195
rect 1502 -229 1536 -195
rect 1911 -211 1945 -177
rect 2334 -198 2368 -164
rect 2406 -198 2440 -164
rect 928 -242 962 -238
rect 928 -272 962 -242
rect 928 -344 962 -310
rect 1911 -339 1945 -305
rect 1018 -405 1052 -371
rect 1096 -405 1130 -371
rect 1174 -405 1208 -371
rect 1252 -405 1286 -371
rect 1330 -405 1364 -371
rect 1408 -405 1442 -371
rect 1486 -405 1520 -371
rect 1564 -405 1598 -371
rect 928 -432 962 -428
rect 928 -462 962 -432
rect 1894 -476 1922 -442
rect 1922 -476 1928 -442
rect 1967 -476 1993 -442
rect 1993 -476 2001 -442
rect 2040 -476 2064 -442
rect 2064 -476 2074 -442
rect 2113 -476 2135 -442
rect 2135 -476 2147 -442
rect 2186 -476 2206 -442
rect 2206 -476 2220 -442
rect 2258 -476 2276 -442
rect 2276 -476 2292 -442
rect 2330 -476 2346 -442
rect 2346 -476 2364 -442
rect 2402 -476 2416 -442
rect 2416 -476 2436 -442
rect 2474 -476 2486 -442
rect 2486 -476 2508 -442
rect 2546 -476 2556 -442
rect 2556 -476 2580 -442
rect 2618 -476 2626 -442
rect 2626 -476 2652 -442
rect 2690 -476 2724 -442
rect 928 -534 962 -500
rect 1018 -581 1052 -547
rect 1095 -581 1129 -547
rect 1172 -581 1206 -547
rect 1249 -581 1283 -547
rect 1326 -581 1360 -547
rect 1403 -581 1437 -547
rect 1480 -581 1514 -547
rect 1557 -581 1591 -547
rect 1861 -565 1895 -531
rect 1941 -565 1975 -531
rect 2576 -565 2610 -531
rect 2648 -565 2682 -531
rect 2258 -640 2292 -606
rect 2330 -640 2364 -606
<< metal1 >>
rect -443 6004 -391 6010
rect -443 5927 -391 5952
tri -391 5921 -360 5952 sw
rect -391 5875 -181 5921
rect -443 5869 -181 5875
rect -129 5869 -104 5921
rect -52 5869 -46 5921
rect 24 5869 30 5921
rect 82 5869 107 5921
rect 159 5869 165 5921
tri 598 5869 623 5894 sw
rect 598 5861 623 5869
tri 623 5861 631 5869 sw
rect 210 5855 2303 5861
rect 210 5821 242 5855
rect 276 5821 316 5855
rect 350 5821 390 5855
rect 424 5821 464 5855
rect 498 5821 538 5855
rect 572 5821 612 5855
rect 646 5821 686 5855
rect 720 5821 760 5855
rect 794 5821 834 5855
rect 868 5821 908 5855
rect 942 5821 982 5855
rect 1016 5821 1056 5855
rect 1090 5821 1130 5855
rect 1164 5821 1204 5855
rect 1238 5821 1278 5855
rect 1312 5821 1352 5855
rect 1386 5821 1426 5855
rect 1460 5821 1500 5855
rect 1534 5821 1574 5855
rect 1608 5821 1648 5855
rect 1682 5821 1722 5855
rect 1756 5821 1796 5855
rect 1830 5821 1870 5855
rect 1904 5821 1944 5855
rect 1978 5821 2018 5855
rect 2052 5821 2091 5855
rect 2125 5821 2164 5855
rect 2198 5821 2237 5855
rect 2271 5821 2303 5855
rect -537 5802 -299 5814
rect -537 5768 -531 5802
rect -497 5768 -435 5802
rect -401 5768 -339 5802
rect -305 5768 -299 5802
rect -537 5728 -299 5768
rect -110 5763 -104 5815
rect -52 5763 -33 5815
rect 19 5763 38 5815
rect 90 5763 96 5815
rect 210 5772 2303 5821
rect -537 5694 -531 5728
rect -497 5694 -435 5728
rect -401 5694 -339 5728
rect -305 5694 -299 5728
rect -537 5654 -299 5694
rect 210 5738 242 5772
rect 276 5738 316 5772
rect 350 5738 390 5772
rect 424 5738 464 5772
rect 498 5738 538 5772
rect 572 5738 612 5772
rect 646 5738 686 5772
rect 720 5738 760 5772
rect 794 5738 834 5772
rect 868 5738 908 5772
rect 942 5738 982 5772
rect 1016 5738 1056 5772
rect 1090 5738 1130 5772
rect 1164 5738 1204 5772
rect 1238 5738 1278 5772
rect 1312 5738 1352 5772
rect 1386 5738 1426 5772
rect 1460 5738 1500 5772
rect 1534 5738 1574 5772
rect 1608 5738 1648 5772
rect 1682 5738 1722 5772
rect 1756 5738 1796 5772
rect 1830 5738 1870 5772
rect 1904 5738 1944 5772
rect 1978 5738 2018 5772
rect 2052 5738 2091 5772
rect 2125 5738 2164 5772
rect 2198 5738 2237 5772
rect 2271 5738 2303 5772
rect 210 5689 2303 5738
rect -537 5620 -531 5654
rect -497 5620 -435 5654
rect -401 5620 -339 5654
rect -305 5620 -299 5654
rect -537 5580 -299 5620
rect -110 5608 -104 5660
rect -52 5608 -33 5660
rect 19 5608 38 5660
rect 90 5608 96 5660
rect 210 5655 242 5689
rect 276 5655 316 5689
rect 350 5655 390 5689
rect 424 5655 464 5689
rect 498 5655 538 5689
rect 572 5655 612 5689
rect 646 5655 686 5689
rect 720 5655 760 5689
rect 794 5655 834 5689
rect 868 5655 908 5689
rect 942 5655 982 5689
rect 1016 5655 1056 5689
rect 1090 5655 1130 5689
rect 1164 5655 1204 5689
rect 1238 5655 1278 5689
rect 1312 5655 1352 5689
rect 1386 5655 1426 5689
rect 1460 5655 1500 5689
rect 1534 5655 1574 5689
rect 1608 5655 1648 5689
rect 1682 5655 1722 5689
rect 1756 5655 1796 5689
rect 1830 5655 1870 5689
rect 1904 5655 1944 5689
rect 1978 5655 2018 5689
rect 2052 5655 2091 5689
rect 2125 5655 2164 5689
rect 2198 5655 2237 5689
rect 2271 5655 2303 5689
rect 210 5649 2303 5655
tri 1722 5610 1761 5649 ne
rect 1761 5610 2302 5649
tri 2302 5648 2303 5649 nw
tri 787 5608 789 5610 se
rect 789 5608 1656 5610
tri 785 5606 787 5608 se
rect 787 5606 1656 5608
rect -537 5546 -531 5580
rect -497 5546 -435 5580
rect -401 5546 -339 5580
rect -305 5546 -299 5580
tri 265 5577 294 5606 se
rect 294 5577 470 5606
tri 255 5567 265 5577 se
rect 265 5567 470 5577
rect -537 5506 -299 5546
rect -537 5472 -531 5506
rect -497 5472 -435 5506
rect -401 5472 -339 5506
rect -305 5472 -299 5506
rect 61 5554 470 5567
rect 522 5554 559 5606
rect 611 5554 617 5606
tri 756 5577 785 5606 se
rect 785 5577 1656 5606
tri 1761 5577 1794 5610 ne
rect 1794 5577 2302 5610
tri 733 5554 756 5577 se
rect 756 5558 1656 5577
rect 756 5554 796 5558
rect 61 5543 305 5554
tri 305 5543 316 5554 nw
tri 722 5543 733 5554 se
rect 733 5543 796 5554
tri 796 5543 811 5558 nw
tri 1330 5543 1345 5558 ne
rect 1345 5543 1656 5558
tri 1794 5543 1828 5577 ne
rect 1828 5543 1970 5577
rect 2004 5543 2042 5577
rect 2076 5543 2114 5577
rect 2148 5543 2186 5577
rect 2220 5543 2258 5577
rect 2292 5543 2302 5577
rect 61 5523 285 5543
tri 285 5523 305 5543 nw
tri 715 5536 722 5543 se
rect 722 5536 789 5543
tri 789 5536 796 5543 nw
tri 1345 5536 1352 5543 ne
rect 1352 5536 1656 5543
tri 705 5526 715 5536 se
rect 715 5526 770 5536
rect 61 5517 284 5523
tri 284 5522 285 5523 nw
rect 61 5483 73 5517
rect 107 5483 156 5517
rect 190 5483 238 5517
rect 272 5483 284 5517
rect 61 5477 284 5483
rect 396 5474 402 5526
rect 454 5474 466 5526
rect 518 5517 573 5526
tri 696 5517 705 5526 se
rect 705 5517 770 5526
tri 770 5517 789 5536 nw
tri 1352 5526 1362 5536 ne
rect 1362 5526 1656 5536
rect 518 5483 527 5517
rect 561 5483 573 5517
tri 662 5483 696 5517 se
rect 696 5483 736 5517
tri 736 5483 770 5517 nw
rect 518 5474 573 5483
tri 653 5474 662 5483 se
rect 662 5474 722 5483
rect -537 5432 -299 5472
tri 648 5469 653 5474 se
rect 653 5469 722 5474
tri 722 5469 736 5483 nw
rect 852 5474 858 5526
rect 910 5474 922 5526
rect 974 5517 1075 5526
tri 1362 5524 1364 5526 ne
rect 981 5483 1029 5517
rect 1063 5483 1075 5517
rect 974 5474 1075 5483
rect 1364 5517 1656 5526
rect 1364 5483 1445 5517
rect 1479 5483 1528 5517
rect 1562 5483 1610 5517
rect 1644 5483 1656 5517
tri 1828 5504 1867 5543 ne
rect 1364 5477 1656 5483
rect 1867 5503 2302 5543
rect 1867 5469 1970 5503
rect 2004 5469 2042 5503
rect 2076 5469 2114 5503
rect 2148 5469 2186 5503
rect 2220 5469 2258 5503
rect 2292 5469 2302 5503
tri 641 5462 648 5469 se
rect 648 5462 715 5469
tri 715 5462 722 5469 nw
tri 619 5440 641 5462 se
rect 641 5440 691 5462
rect -537 5398 -531 5432
rect -497 5398 -435 5432
rect -401 5398 -339 5432
rect -305 5428 -299 5432
tri -299 5428 -287 5440 sw
tri 617 5438 619 5440 se
rect 619 5438 691 5440
tri 691 5438 715 5462 nw
rect 27 5428 681 5438
tri 681 5428 691 5438 nw
rect 771 5432 1615 5438
rect -305 5426 -287 5428
tri -287 5426 -285 5428 sw
rect 27 5426 679 5428
tri 679 5426 681 5428 nw
rect -305 5398 -285 5426
rect -537 5392 -285 5398
tri -285 5392 -251 5426 sw
rect 27 5392 39 5426
rect 73 5392 551 5426
rect 585 5392 645 5426
tri 645 5392 679 5426 nw
rect -537 5358 -251 5392
rect -537 5324 -531 5358
rect -497 5324 -435 5358
rect -401 5324 -339 5358
rect -305 5353 -251 5358
tri -251 5353 -212 5392 sw
rect 27 5386 639 5392
tri 639 5386 645 5392 nw
rect 27 5353 592 5386
tri 592 5353 625 5386 nw
rect 823 5426 1615 5432
rect 823 5392 1063 5426
rect 1097 5392 1575 5426
rect 1609 5392 1615 5426
rect 823 5380 1615 5392
rect 771 5368 1615 5380
rect -305 5349 -212 5353
tri -212 5349 -208 5353 sw
rect 27 5350 591 5353
tri 591 5352 592 5353 nw
rect 27 5349 112 5350
tri 112 5349 113 5350 nw
tri 511 5349 512 5350 ne
rect 512 5349 591 5350
rect -305 5334 -208 5349
tri -208 5334 -193 5349 sw
rect 27 5334 79 5349
rect -305 5324 -193 5334
rect -537 5318 -193 5324
tri -193 5318 -177 5334 sw
rect -537 5306 -177 5318
rect -537 5284 -217 5306
rect -537 5250 -531 5284
rect -497 5250 -435 5284
rect -401 5250 -339 5284
rect -305 5272 -217 5284
rect -183 5272 -177 5306
rect -305 5250 -177 5272
rect -537 5221 -177 5250
rect -537 5210 -217 5221
rect -537 5176 -531 5210
rect -497 5176 -435 5210
rect -401 5176 -339 5210
rect -305 5187 -217 5210
rect -183 5187 -177 5221
rect -305 5176 -177 5187
rect 27 5300 39 5334
rect 73 5300 79 5334
tri 79 5316 112 5349 nw
tri 512 5318 543 5349 ne
rect 543 5318 551 5349
rect 27 5241 79 5300
rect 27 5224 39 5241
rect 73 5224 79 5241
rect -537 5159 -177 5176
tri -177 5159 -157 5179 sw
rect 27 5160 79 5172
rect -537 5150 -157 5159
tri -157 5150 -148 5159 sw
rect -537 5148 -148 5150
tri -148 5148 -146 5150 sw
rect -537 5136 -146 5148
rect -537 5102 -531 5136
rect -497 5102 -435 5136
rect -401 5102 -339 5136
rect -305 5102 -217 5136
rect -183 5114 -146 5136
tri -146 5114 -112 5148 sw
rect -183 5102 -112 5114
tri -112 5102 -100 5114 sw
rect 27 5102 79 5108
rect 289 5306 335 5318
tri 543 5316 545 5318 ne
rect 289 5272 295 5306
rect 329 5272 335 5306
rect 289 5221 335 5272
rect 289 5187 295 5221
rect 329 5187 335 5221
rect 289 5136 335 5187
rect 289 5102 295 5136
rect 329 5102 335 5136
rect -537 5081 -100 5102
tri -100 5081 -79 5102 sw
rect -537 5068 -79 5081
tri -79 5068 -66 5081 sw
rect -537 5062 -66 5068
rect -537 5028 -531 5062
rect -497 5028 -435 5062
rect -401 5028 -339 5062
rect -305 5060 -66 5062
tri -66 5060 -58 5068 sw
rect -305 5051 -58 5060
tri -58 5051 -49 5060 sw
rect 289 5051 335 5102
rect -305 5028 -217 5051
rect -537 5017 -217 5028
rect -183 5017 -49 5051
tri -49 5017 -15 5051 sw
rect 289 5017 295 5051
rect 329 5017 335 5051
rect -537 5003 -15 5017
tri -15 5003 -1 5017 sw
rect -537 4994 -1 5003
tri -1 4994 8 5003 sw
rect -537 4988 8 4994
rect -537 4954 -531 4988
rect -497 4954 -435 4988
rect -401 4954 -339 4988
rect -305 4978 8 4988
tri 8 4978 24 4994 sw
tri 274 4978 289 4993 se
rect 289 4978 335 5017
rect 545 5315 551 5318
rect 585 5315 591 5349
rect 545 5271 591 5315
rect 823 5350 1615 5368
rect 823 5349 856 5350
tri 856 5349 857 5350 nw
tri 1023 5349 1024 5350 ne
rect 1024 5349 1136 5350
tri 1136 5349 1137 5350 nw
tri 1535 5349 1536 5350 ne
rect 1536 5349 1615 5350
tri 823 5316 856 5349 nw
tri 1024 5316 1057 5349 ne
rect 771 5310 823 5316
rect 1057 5315 1063 5349
rect 1097 5315 1103 5349
tri 1103 5316 1136 5349 nw
tri 1536 5318 1567 5349 ne
rect 1567 5318 1575 5349
rect 545 5237 551 5271
rect 585 5237 591 5271
rect 1057 5271 1103 5315
rect 545 5193 591 5237
rect 545 5159 551 5193
rect 585 5159 591 5193
rect 545 5115 591 5159
rect 545 5081 551 5115
rect 585 5081 591 5115
rect 545 5037 591 5081
rect 545 5003 551 5037
rect 585 5003 591 5037
tri 335 4978 350 4993 sw
rect 545 4991 591 5003
rect 801 5239 847 5251
rect 801 5205 807 5239
rect 841 5205 847 5239
rect 801 5150 847 5205
rect 801 5116 807 5150
rect 841 5116 847 5150
rect 801 5060 847 5116
rect 801 5026 807 5060
rect 841 5026 847 5060
tri 799 4991 801 4993 se
rect 801 4991 847 5026
rect 1057 5237 1063 5271
rect 1097 5237 1103 5271
rect 1057 5193 1103 5237
rect 1057 5159 1063 5193
rect 1097 5159 1103 5193
rect 1057 5115 1103 5159
rect 1057 5081 1063 5115
rect 1097 5081 1103 5115
rect 1057 5037 1103 5081
rect 1057 5003 1063 5037
rect 1097 5003 1103 5037
tri 786 4978 799 4991 se
rect 799 4978 847 4991
tri 847 4978 862 4993 sw
rect 1057 4991 1103 5003
rect 1313 5306 1359 5318
tri 1567 5316 1569 5318 ne
rect 1313 5272 1319 5306
rect 1353 5272 1359 5306
rect 1313 5221 1359 5272
rect 1313 5187 1319 5221
rect 1353 5187 1359 5221
rect 1313 5136 1359 5187
rect 1313 5102 1319 5136
rect 1353 5102 1359 5136
rect 1313 5051 1359 5102
rect 1313 5017 1319 5051
rect 1353 5017 1359 5051
tri 1311 4991 1313 4993 se
rect 1313 4991 1359 5017
rect 1569 5315 1575 5318
rect 1609 5315 1615 5349
rect 1569 5271 1615 5315
rect 1867 5428 2302 5469
rect 1867 5394 1970 5428
rect 2004 5394 2042 5428
rect 2076 5394 2114 5428
rect 2148 5394 2186 5428
rect 2220 5394 2258 5428
rect 2292 5394 2302 5428
rect 1867 5353 2302 5394
rect 1867 5319 1970 5353
rect 2004 5319 2042 5353
rect 2076 5319 2114 5353
rect 2148 5319 2186 5353
rect 2220 5319 2258 5353
rect 2292 5319 2302 5353
tri 1842 5278 1867 5303 se
rect 1867 5278 2302 5319
rect 1569 5237 1575 5271
rect 1609 5237 1615 5271
rect 1569 5193 1615 5237
rect 1569 5159 1575 5193
rect 1609 5159 1615 5193
rect 1569 5115 1615 5159
tri 1825 5261 1842 5278 se
rect 1842 5261 1970 5278
rect 1825 5249 1970 5261
rect 1825 5215 1831 5249
rect 1865 5244 1970 5249
rect 2004 5244 2042 5278
rect 2076 5244 2114 5278
rect 2148 5244 2186 5278
rect 2220 5244 2258 5278
rect 2292 5244 2302 5278
rect 1865 5215 2302 5244
rect 1825 5203 2302 5215
rect 1825 5176 1970 5203
rect 1825 5142 1831 5176
rect 1865 5169 1970 5176
rect 2004 5169 2042 5203
rect 2076 5169 2114 5203
rect 2148 5169 2186 5203
rect 2220 5169 2258 5203
rect 2292 5169 2302 5203
rect 1865 5142 2302 5169
rect 1825 5128 2302 5142
rect 1569 5081 1575 5115
rect 1609 5081 1615 5115
tri 1810 5102 1825 5117 se
rect 1825 5102 1970 5128
rect 1569 5037 1615 5081
tri 1776 5068 1810 5102 se
rect 1810 5068 1831 5102
rect 1865 5094 1970 5102
rect 2004 5094 2042 5128
rect 2076 5094 2114 5128
rect 2148 5094 2186 5128
rect 2220 5094 2258 5128
rect 2292 5094 2302 5128
rect 1865 5068 2302 5094
tri 1761 5053 1776 5068 se
rect 1776 5053 2302 5068
rect 1569 5003 1575 5037
rect 1609 5003 1615 5037
tri 1736 5028 1761 5053 se
rect 1761 5028 1970 5053
tri 1298 4978 1311 4991 se
rect 1311 4978 1359 4991
tri 1359 4978 1374 4993 sw
rect 1569 4991 1615 5003
tri 1702 4994 1736 5028 se
rect 1736 4994 1831 5028
rect 1865 5019 1970 5028
rect 2004 5019 2042 5053
rect 2076 5019 2114 5053
rect 2148 5019 2186 5053
rect 2220 5019 2258 5053
rect 2292 5019 2302 5053
rect 1865 4994 2302 5019
tri 1699 4991 1702 4994 se
rect 1702 4991 2302 4994
tri 1686 4978 1699 4991 se
rect 1699 4978 2302 4991
rect -305 4970 24 4978
tri 24 4970 32 4978 sw
tri 266 4970 274 4978 se
rect 274 4970 350 4978
tri 350 4970 358 4978 sw
tri 778 4970 786 4978 se
rect 786 4970 862 4978
rect -305 4966 32 4970
tri 32 4966 36 4970 sw
tri 262 4966 266 4970 se
rect 266 4966 358 4970
rect -305 4954 -217 4966
rect -537 4932 -217 4954
rect -183 4959 36 4966
tri 36 4959 43 4966 sw
tri 255 4959 262 4966 se
rect 262 4959 295 4966
rect -183 4932 295 4959
rect 329 4959 358 4966
tri 358 4959 369 4970 sw
tri 767 4959 778 4970 se
rect 778 4959 807 4970
rect 329 4936 807 4959
rect 841 4966 862 4970
tri 862 4966 874 4978 sw
tri 1286 4966 1298 4978 se
rect 1298 4966 1374 4978
rect 841 4959 874 4966
tri 874 4959 881 4966 sw
tri 1279 4959 1286 4966 se
rect 1286 4959 1319 4966
rect 841 4936 1319 4959
rect 329 4932 1319 4936
rect 1353 4959 1374 4966
tri 1374 4959 1393 4978 sw
tri 1667 4959 1686 4978 se
rect 1686 4959 1970 4978
rect 1353 4954 1970 4959
rect 1353 4932 1831 4954
rect -537 4920 1831 4932
rect 1865 4944 1970 4954
rect 2004 4944 2042 4978
rect 2076 4944 2114 4978
rect 2148 4944 2186 4978
rect 2220 4944 2258 4978
rect 2292 4944 2302 4978
rect 1865 4920 2302 4944
rect -537 4914 2302 4920
rect -537 4880 -531 4914
rect -497 4880 -435 4914
rect -401 4880 -339 4914
rect -305 4903 2302 4914
rect -305 4880 1970 4903
rect -537 4846 -217 4880
rect -183 4846 295 4880
rect 329 4846 807 4880
rect 841 4846 1319 4880
rect 1353 4846 1831 4880
rect 1865 4869 1970 4880
rect 2004 4869 2042 4903
rect 2076 4869 2114 4903
rect 2148 4869 2186 4903
rect 2220 4869 2258 4903
rect 2292 4869 2302 4903
rect 1865 4846 2302 4869
rect -537 4840 2302 4846
rect -537 4806 -531 4840
rect -497 4806 -435 4840
rect -401 4806 -339 4840
rect -305 4828 2302 4840
rect -305 4806 1970 4828
rect -537 4794 1970 4806
rect 2004 4794 2042 4828
rect 2076 4794 2114 4828
rect 2148 4794 2186 4828
rect 2220 4794 2258 4828
rect 2292 4794 2302 4828
rect -537 4766 2302 4794
rect -537 4732 -531 4766
rect -497 4732 -435 4766
rect -401 4732 -339 4766
rect -305 4732 2302 4766
rect -537 4729 2302 4732
rect -537 4695 -198 4729
rect -164 4695 -125 4729
rect -91 4695 -52 4729
rect -18 4695 21 4729
rect 55 4695 94 4729
rect 128 4695 167 4729
rect 201 4695 240 4729
rect 274 4695 312 4729
rect 346 4695 384 4729
rect 418 4695 456 4729
rect 490 4695 528 4729
rect 562 4695 600 4729
rect 634 4695 672 4729
rect 706 4695 744 4729
rect 778 4695 816 4729
rect 850 4695 888 4729
rect 922 4695 960 4729
rect 994 4695 1032 4729
rect 1066 4695 1104 4729
rect 1138 4695 1176 4729
rect 1210 4695 1248 4729
rect 1282 4695 1320 4729
rect 1354 4695 1392 4729
rect 1426 4695 1464 4729
rect 1498 4695 1536 4729
rect 1570 4695 1608 4729
rect 1642 4695 1680 4729
rect 1714 4695 1752 4729
rect 1786 4695 1824 4729
rect 1858 4695 1896 4729
rect 1930 4695 1968 4729
rect 2002 4695 2040 4729
rect 2074 4695 2302 4729
rect -537 4692 2302 4695
rect -537 4658 -531 4692
rect -497 4658 -435 4692
rect -401 4658 -339 4692
rect -305 4665 2302 4692
rect -305 4658 -137 4665
rect -537 4618 -137 4658
rect -537 4584 -531 4618
rect -497 4584 -435 4618
rect -401 4584 -339 4618
rect -305 4593 -137 4618
tri -137 4593 -65 4665 nw
tri 365 4631 399 4665 ne
rect 399 4593 445 4665
tri 445 4631 479 4665 nw
tri 1675 4631 1709 4665 ne
rect 1709 4631 2302 4665
tri 1709 4605 1735 4631 ne
rect 1735 4605 2302 4631
rect -305 4584 -171 4593
rect -537 4559 -171 4584
tri -171 4559 -137 4593 nw
rect 399 4559 405 4593
rect 439 4559 445 4593
rect -537 4550 -180 4559
tri -180 4550 -171 4559 nw
rect -537 4544 -209 4550
rect -537 4510 -531 4544
rect -497 4510 -435 4544
rect -401 4510 -339 4544
rect -305 4521 -209 4544
tri -209 4521 -180 4550 nw
rect -305 4513 -217 4521
tri -217 4513 -209 4521 nw
rect 223 4513 269 4525
rect -305 4510 -251 4513
rect -537 4479 -251 4510
tri -251 4479 -217 4513 nw
rect 223 4479 229 4513
rect 263 4479 269 4513
rect 399 4521 445 4559
rect 399 4487 405 4521
rect 439 4487 445 4521
rect -537 4470 -277 4479
rect -537 4436 -531 4470
rect -497 4436 -435 4470
rect -401 4436 -339 4470
rect -305 4453 -277 4470
tri -277 4453 -251 4479 nw
rect 223 4453 269 4479
tri 269 4453 297 4481 sw
rect 399 4475 445 4487
rect 575 4593 621 4605
tri 1735 4596 1744 4605 ne
rect 1744 4596 2302 4605
rect 575 4559 581 4593
rect 615 4563 621 4593
tri 621 4563 654 4596 sw
tri 1744 4563 1777 4596 ne
rect 1777 4563 2302 4596
rect 615 4562 654 4563
tri 654 4562 655 4563 sw
tri 1777 4562 1778 4563 ne
rect 1778 4562 1827 4563
rect 615 4559 1054 4562
rect 575 4521 1054 4559
rect 575 4487 581 4521
rect 615 4510 1054 4521
rect 1106 4510 1118 4562
rect 1170 4550 1368 4562
tri 1778 4556 1784 4562 ne
rect 1784 4556 1827 4562
tri 1485 4550 1491 4556 se
rect 1491 4550 1644 4556
rect 1170 4516 1174 4550
rect 1208 4516 1248 4550
rect 1282 4516 1322 4550
rect 1356 4516 1368 4550
tri 1451 4516 1485 4550 se
rect 1485 4516 1526 4550
rect 1560 4516 1598 4550
rect 1632 4516 1644 4550
tri 1784 4529 1811 4556 ne
rect 1811 4529 1827 4556
rect 1861 4529 1899 4563
rect 1933 4529 1971 4563
rect 2005 4529 2043 4563
rect 2077 4529 2115 4563
rect 2149 4529 2187 4563
rect 2221 4529 2259 4563
rect 2293 4529 2302 4563
tri 1811 4519 1821 4529 ne
rect 1170 4510 1368 4516
tri 1445 4510 1451 4516 se
rect 1451 4510 1644 4516
rect 615 4487 632 4510
tri 632 4487 655 4510 nw
tri 1424 4489 1445 4510 se
rect 1445 4489 1644 4510
tri 1422 4487 1424 4489 se
rect 1424 4487 1496 4489
tri 1496 4487 1498 4489 nw
rect 1821 4487 2302 4529
rect 575 4475 621 4487
tri 621 4476 632 4487 nw
tri 1411 4476 1422 4487 se
rect 1422 4476 1478 4487
tri 1410 4475 1411 4476 se
rect 1411 4475 1478 4476
tri 1404 4469 1410 4475 se
rect 1410 4469 1478 4475
tri 1478 4469 1496 4487 nw
tri 1388 4453 1404 4469 se
rect 1404 4453 1462 4469
tri 1462 4453 1478 4469 nw
rect 1821 4453 1827 4487
rect 1861 4453 1899 4487
rect 1933 4453 1971 4487
rect 2005 4453 2043 4487
rect 2077 4453 2115 4487
rect 2149 4453 2187 4487
rect 2221 4453 2259 4487
rect 2293 4453 2302 4487
rect -305 4441 -289 4453
tri -289 4441 -277 4453 nw
rect 27 4443 79 4449
rect -305 4436 -299 4441
rect -537 4396 -299 4436
tri -299 4431 -289 4441 nw
rect -537 4362 -531 4396
rect -497 4362 -435 4396
rect -401 4362 -339 4396
rect -305 4362 -299 4396
rect -537 4322 -299 4362
rect -537 4288 -531 4322
rect -497 4288 -435 4322
rect -401 4288 -339 4322
rect -305 4288 -299 4322
rect 223 4447 297 4453
tri 297 4447 303 4453 sw
tri 1382 4447 1388 4453 se
rect 1388 4447 1420 4453
rect 223 4441 1420 4447
rect 223 4407 229 4441
rect 263 4407 1204 4441
rect 27 4379 79 4391
tri 79 4377 103 4401 sw
rect 223 4395 1204 4407
tri 1170 4377 1188 4395 ne
rect 1188 4389 1204 4395
rect 1256 4411 1420 4441
tri 1420 4411 1462 4453 nw
rect 1821 4411 2302 4453
rect 1256 4395 1404 4411
tri 1404 4395 1420 4411 nw
rect 1256 4389 1272 4395
rect 1188 4377 1272 4389
tri 1272 4377 1290 4395 nw
rect 1821 4377 1827 4411
rect 1861 4377 1899 4411
rect 1933 4377 1971 4411
rect 2005 4377 2043 4411
rect 2077 4377 2115 4411
rect 2149 4377 2187 4411
rect 2221 4377 2259 4411
rect 2293 4377 2302 4411
rect 79 4367 103 4377
tri 103 4367 113 4377 sw
tri 1188 4367 1198 4377 ne
rect 1198 4367 1204 4377
rect 79 4361 390 4367
rect 79 4327 272 4361
rect 306 4327 344 4361
rect 378 4327 390 4361
rect 27 4321 390 4327
rect 450 4361 823 4367
tri 1198 4361 1204 4367 ne
rect 450 4327 462 4361
rect 496 4327 534 4361
rect 568 4327 771 4361
rect 450 4321 771 4327
tri 737 4317 741 4321 ne
rect 741 4317 771 4321
tri 741 4305 753 4317 ne
rect 753 4309 771 4317
tri 1256 4361 1272 4377 nw
rect 1204 4319 1256 4325
rect 1636 4351 1688 4363
rect 1636 4317 1645 4351
rect 1679 4317 1688 4351
rect 753 4305 823 4309
rect -537 4248 -299 4288
tri 753 4287 771 4305 ne
rect 771 4297 823 4305
rect -537 4214 -531 4248
rect -497 4214 -435 4248
rect -401 4214 -339 4248
rect -305 4214 -299 4248
rect 1287 4305 1339 4317
rect 771 4239 823 4245
rect 852 4268 904 4274
tri 851 4225 852 4226 se
rect -537 4174 -299 4214
tri 832 4206 851 4225 se
rect 851 4216 852 4225
rect 851 4206 904 4216
tri 818 4192 832 4206 se
rect 832 4204 904 4206
rect 832 4192 852 4204
rect -537 4140 -531 4174
rect -497 4140 -435 4174
rect -401 4140 -339 4174
rect -305 4140 -299 4174
rect 398 4186 852 4192
rect 398 4152 410 4186
rect 444 4152 482 4186
rect 516 4152 852 4186
rect 1287 4271 1293 4305
rect 1327 4271 1339 4305
rect 1287 4206 1339 4271
rect 398 4146 904 4152
rect 1111 4183 1157 4195
rect 1111 4149 1117 4183
rect 1151 4149 1157 4183
rect -537 4100 -299 4140
rect -537 4066 -531 4100
rect -497 4066 -435 4100
rect -401 4066 -339 4100
rect -305 4066 -299 4100
rect -537 4026 -299 4066
rect 396 4096 448 4108
rect 396 4087 405 4096
rect 439 4087 448 4096
rect -537 3992 -531 4026
rect -497 3992 -435 4026
rect -401 3992 -339 4026
rect -305 3992 -299 4026
rect -537 3952 -299 3992
rect -537 3918 -531 3952
rect -497 3918 -435 3952
rect -401 3918 -339 3952
rect -305 3918 -299 3952
rect 223 4024 269 4036
rect 223 3990 229 4024
rect 263 3990 269 4024
rect 223 3952 269 3990
rect 1111 4080 1157 4149
rect 1111 4046 1117 4080
rect 1151 4046 1157 4080
rect 1287 4182 1293 4206
rect 1327 4182 1339 4206
rect 1636 4270 1688 4317
rect 1636 4236 1645 4270
rect 1679 4236 1688 4270
rect 1287 4118 1339 4130
tri 1157 4046 1173 4062 sw
rect 1287 4060 1339 4066
rect 1463 4183 1509 4195
rect 1463 4149 1469 4183
rect 1503 4149 1509 4183
rect 1463 4080 1509 4149
tri 1461 4060 1463 4062 se
rect 1463 4060 1469 4080
tri 1447 4046 1461 4060 se
rect 1461 4046 1469 4060
rect 1503 4046 1509 4080
rect 1636 4188 1688 4236
rect 1636 4182 1645 4188
rect 1679 4182 1688 4188
rect 1636 4118 1688 4130
rect 396 4024 448 4035
rect 396 4023 405 4024
rect 439 4023 448 4024
rect 396 3965 448 3971
rect 575 4024 621 4036
rect 575 3990 581 4024
rect 615 3990 621 4024
tri -299 3918 -296 3921 sw
rect 223 3918 229 3952
rect 263 3918 269 3952
rect -537 3879 -296 3918
tri -296 3879 -257 3918 sw
rect -537 3878 -257 3879
rect -537 3844 -531 3878
rect -497 3844 -435 3878
rect -401 3844 -339 3878
rect -305 3845 -257 3878
tri -257 3845 -223 3879 sw
rect -305 3844 -223 3845
rect -537 3803 -223 3844
rect -537 3769 -531 3803
rect -497 3769 -435 3803
rect -401 3769 -339 3803
rect -305 3802 -223 3803
tri -223 3802 -180 3845 sw
rect -305 3769 -180 3802
rect -537 3768 -180 3769
tri -180 3768 -146 3802 sw
rect -537 3728 -146 3768
rect -537 3694 -531 3728
rect -497 3694 -435 3728
rect -401 3694 -339 3728
rect -305 3726 -146 3728
tri -146 3726 -104 3768 sw
tri 195 3726 223 3754 se
rect 223 3726 269 3918
rect 575 3952 621 3990
rect 575 3918 581 3952
rect 615 3918 621 3952
tri 269 3726 297 3754 sw
tri 547 3726 575 3754 se
rect 575 3726 621 3918
rect 1111 4031 1173 4046
tri 1173 4031 1188 4046 sw
tri 1432 4031 1447 4046 se
rect 1447 4031 1509 4046
tri 1509 4031 1540 4062 sw
rect 1636 4060 1688 4066
rect 1821 4335 2302 4377
rect 1821 4301 1827 4335
rect 1861 4301 1899 4335
rect 1933 4301 1971 4335
rect 2005 4301 2043 4335
rect 2077 4301 2115 4335
rect 2149 4301 2187 4335
rect 2221 4301 2259 4335
rect 2293 4301 2302 4335
rect 1821 4259 2302 4301
rect 1821 4225 1827 4259
rect 1861 4225 1899 4259
rect 1933 4225 1971 4259
rect 2005 4225 2043 4259
rect 2077 4225 2115 4259
rect 2149 4225 2187 4259
rect 2221 4225 2259 4259
rect 2293 4225 2302 4259
rect 1821 4183 2302 4225
rect 1821 4149 1827 4183
rect 1861 4149 1899 4183
rect 1933 4149 1971 4183
rect 2005 4149 2043 4183
rect 2077 4149 2115 4183
rect 2149 4149 2187 4183
rect 2221 4149 2259 4183
rect 2293 4149 2302 4183
rect 1821 4107 2302 4149
rect 1821 4073 1827 4107
rect 1861 4073 1899 4107
rect 1933 4073 1971 4107
rect 2005 4073 2043 4107
rect 2077 4073 2115 4107
rect 2149 4073 2187 4107
rect 2221 4073 2259 4107
rect 2293 4073 2302 4107
rect 1821 4031 2302 4073
rect 1111 4028 1188 4031
tri 1188 4028 1191 4031 sw
tri 1429 4028 1432 4031 se
rect 1432 4028 1540 4031
tri 1540 4028 1543 4031 sw
rect 1111 3976 1545 4028
rect 1111 3942 1117 3976
rect 1151 3942 1469 3976
rect 1503 3942 1545 3976
rect 1111 3802 1545 3942
rect 1821 3997 1827 4031
rect 1861 3997 1899 4031
rect 1933 3997 1971 4031
rect 2005 3997 2043 4031
rect 2077 3997 2115 4031
rect 2149 3997 2187 4031
rect 2221 3997 2259 4031
rect 2293 3997 2302 4031
rect 1821 3955 2302 3997
rect 1821 3921 1827 3955
rect 1861 3921 1899 3955
rect 1933 3921 1971 3955
rect 2005 3921 2043 3955
rect 2077 3921 2115 3955
rect 2149 3921 2187 3955
rect 2221 3921 2259 3955
rect 2293 3921 2302 3955
rect 1821 3879 2302 3921
rect 1821 3845 1827 3879
rect 1861 3845 1899 3879
rect 1933 3845 1971 3879
rect 2005 3845 2043 3879
rect 2077 3845 2115 3879
rect 2149 3845 2187 3879
rect 2221 3845 2259 3879
rect 2293 3845 2302 3879
tri 1810 3805 1821 3816 se
rect 1821 3805 2302 3845
tri 1545 3802 1548 3805 sw
tri 1807 3802 1810 3805 se
rect 1810 3802 2302 3805
tri 1085 3768 1111 3794 se
rect 1111 3768 1548 3802
tri 1548 3768 1582 3802 sw
tri 1773 3768 1807 3802 se
rect 1807 3768 1827 3802
rect 1861 3768 1899 3802
rect 1933 3768 1971 3802
rect 2005 3768 2043 3802
rect 2077 3768 2115 3802
rect 2149 3768 2187 3802
rect 2221 3768 2259 3802
rect 2293 3768 2302 3802
tri 1071 3754 1085 3768 se
rect 1085 3754 1582 3768
tri 621 3726 649 3754 sw
tri 1043 3726 1071 3754 se
rect 1071 3726 1582 3754
tri 1582 3726 1624 3768 sw
tri 1731 3726 1773 3768 se
rect 1773 3726 2302 3768
rect -305 3720 2302 3726
rect -305 3694 -238 3720
rect -537 3686 -238 3694
rect -204 3686 -165 3720
rect -131 3686 -92 3720
rect -58 3686 -19 3720
rect 15 3686 54 3720
rect 88 3686 127 3720
rect 161 3686 200 3720
rect 234 3686 273 3720
rect 307 3686 346 3720
rect 380 3686 419 3720
rect 453 3686 492 3720
rect 526 3686 565 3720
rect 599 3686 638 3720
rect 672 3686 711 3720
rect 745 3686 784 3720
rect 818 3686 857 3720
rect 891 3686 930 3720
rect 964 3686 1003 3720
rect 1037 3686 1076 3720
rect 1110 3686 1149 3720
rect 1183 3686 1222 3720
rect 1256 3686 1295 3720
rect 1329 3686 1368 3720
rect 1402 3686 1441 3720
rect 1475 3686 1514 3720
rect 1548 3686 1587 3720
rect 1621 3686 1660 3720
rect 1694 3686 1733 3720
rect -537 3653 1733 3686
rect -537 3619 -531 3653
rect -497 3619 -435 3653
rect -401 3619 -339 3653
rect -305 3648 1733 3653
rect -305 3619 -238 3648
rect -537 3614 -238 3619
rect -204 3614 -165 3648
rect -131 3614 -92 3648
rect -58 3614 -19 3648
rect 15 3614 54 3648
rect 88 3614 127 3648
rect 161 3614 200 3648
rect 234 3614 273 3648
rect 307 3614 346 3648
rect 380 3614 419 3648
rect 453 3614 492 3648
rect 526 3614 565 3648
rect 599 3614 638 3648
rect 672 3614 711 3648
rect 745 3614 784 3648
rect 818 3614 857 3648
rect 891 3614 930 3648
rect 964 3614 1003 3648
rect 1037 3614 1076 3648
rect 1110 3614 1149 3648
rect 1183 3614 1222 3648
rect 1256 3614 1295 3648
rect 1329 3614 1368 3648
rect 1402 3614 1441 3648
rect 1475 3614 1514 3648
rect 1548 3614 1587 3648
rect 1621 3614 1660 3648
rect 1694 3614 1733 3648
rect -537 3576 1733 3614
rect -537 3542 -238 3576
rect -204 3542 -165 3576
rect -131 3542 -92 3576
rect -58 3542 -19 3576
rect 15 3542 54 3576
rect 88 3542 127 3576
rect 161 3542 200 3576
rect 234 3542 273 3576
rect 307 3542 346 3576
rect 380 3542 419 3576
rect 453 3542 492 3576
rect 526 3542 565 3576
rect 599 3542 638 3576
rect 672 3542 711 3576
rect 745 3542 784 3576
rect 818 3542 857 3576
rect 891 3542 930 3576
rect 964 3542 1003 3576
rect 1037 3542 1076 3576
rect 1110 3542 1149 3576
rect 1183 3542 1222 3576
rect 1256 3542 1295 3576
rect 1329 3542 1368 3576
rect 1402 3542 1441 3576
rect 1475 3542 1514 3576
rect 1548 3542 1587 3576
rect 1621 3542 1660 3576
rect 1694 3542 1733 3576
rect 2271 3542 2302 3720
rect -537 3536 2302 3542
tri 894 3534 896 3536 ne
rect 896 3534 2302 3536
rect -2 1075 428 1367
tri 428 1075 720 1367 nw
tri 769 1123 817 1171 se
rect 817 1140 2456 1171
tri 2456 1140 2487 1171 sw
rect 817 1137 2487 1140
tri 817 1123 831 1137 nw
tri 2442 1123 2456 1137 ne
rect 2456 1123 2487 1137
tri 721 1075 769 1123 se
tri 769 1075 817 1123 nw
tri 2456 1092 2487 1123 ne
tri 2487 1092 2535 1140 sw
tri 2487 1078 2501 1092 ne
rect -2 981 334 1075
tri 334 981 428 1075 nw
tri 717 1071 721 1075 se
rect 721 1071 751 1075
rect -2 947 300 981
tri 300 947 334 981 nw
rect -2 934 287 947
tri 287 934 300 947 nw
rect -2 900 253 934
tri 253 900 287 934 nw
tri 715 900 717 902 se
rect 717 900 751 1071
tri 751 1057 769 1075 nw
rect 852 942 858 994
rect 910 942 922 994
rect 974 942 2437 994
tri 2342 934 2350 942 ne
rect 2350 940 2437 942
rect 2501 987 2535 1092
tri 2535 987 2578 1030 sw
rect 2501 981 2631 987
rect 2501 947 2513 981
rect 2547 947 2585 981
rect 2619 947 2631 981
rect 2501 941 2631 947
rect 2350 934 2385 940
tri 2350 900 2384 934 ne
rect 2384 900 2385 934
rect -2 862 215 900
tri 215 862 253 900 nw
tri 677 862 715 900 se
rect 715 888 751 900
tri 2384 899 2385 900 ne
rect 715 862 725 888
tri 725 862 751 888 nw
rect 2385 876 2437 888
rect -2 828 181 862
tri 181 828 215 862 nw
tri 669 854 677 862 se
rect 677 854 717 862
tri 717 854 725 862 nw
tri 643 828 669 854 se
rect 669 828 691 854
tri 691 828 717 854 nw
rect -2 824 177 828
tri 177 824 181 828 nw
tri 639 824 643 828 se
rect 643 824 678 828
rect -2 806 159 824
tri 159 806 177 824 nw
rect -2 772 125 806
tri 125 772 159 806 nw
rect 400 772 406 824
rect 458 772 470 824
rect 522 815 528 824
tri 528 815 537 824 sw
tri 630 815 639 824 se
rect 639 815 678 824
tri 678 815 691 828 nw
rect 2385 818 2437 824
tri 2791 818 2811 838 se
rect 2811 818 2863 859
tri 2386 816 2388 818 ne
rect 2388 816 2434 818
tri 2434 816 2436 818 nw
tri 2789 816 2791 818 se
rect 2791 816 2863 818
tri 2788 815 2789 816 se
rect 2789 815 2863 816
rect 522 806 669 815
tri 669 806 678 815 nw
tri 2785 812 2788 815 se
rect 2788 812 2863 815
rect 2482 806 2863 812
rect 522 781 644 806
tri 644 781 669 806 nw
rect 522 772 528 781
tri 528 772 537 781 nw
rect 2482 772 2494 806
rect 2528 772 2629 806
rect 2663 772 2863 806
rect -2 700 53 772
tri 53 700 125 772 nw
rect 2482 766 2863 772
tri 2776 731 2811 766 ne
rect 730 700 858 709
rect -2 666 19 700
tri 19 666 53 700 nw
rect 730 666 742 700
rect 776 666 833 700
tri -2 645 19 666 nw
rect 730 657 858 666
rect 910 657 922 709
rect 974 657 980 709
rect 1026 700 1865 706
rect 1917 700 1929 706
rect 1981 700 2322 706
rect 1026 666 1038 700
rect 1072 666 1111 700
rect 1145 666 1184 700
rect 1218 666 1257 700
rect 1291 666 1330 700
rect 1364 666 1403 700
rect 1437 666 1476 700
rect 1510 666 1549 700
rect 1583 666 1622 700
rect 1656 666 1695 700
rect 1729 666 1768 700
rect 1802 666 1841 700
rect 1981 666 1987 700
rect 2021 666 2060 700
rect 2094 666 2132 700
rect 2166 666 2204 700
rect 2238 666 2276 700
rect 2310 666 2322 700
rect 1026 654 1865 666
rect 1917 654 1929 666
rect 1981 660 2322 666
tri 2802 660 2811 669 se
rect 2811 660 2863 766
rect 1981 654 1987 660
tri 1901 645 1910 654 ne
rect 1910 645 1987 654
tri 1910 620 1935 645 ne
rect 119 581 165 593
rect 119 547 125 581
rect 159 547 165 581
rect 119 532 165 547
rect 771 569 823 575
tri 165 532 166 533 sw
tri 770 532 771 533 se
rect 119 509 166 532
rect 119 475 125 509
rect 159 499 166 509
tri 166 499 199 532 sw
tri 737 499 770 532 se
rect 770 517 771 532
tri 823 532 824 533 sw
rect 823 517 824 532
rect 770 505 824 517
rect 770 499 771 505
rect 159 475 771 499
rect 119 453 771 475
rect 823 499 824 505
tri 824 499 857 532 sw
rect 823 498 1018 499
tri 1018 498 1019 499 sw
rect 823 470 1019 498
tri 1019 470 1047 498 sw
rect 823 460 1047 470
tri 1047 460 1057 470 sw
rect 823 453 1057 460
rect 119 447 1057 453
tri 996 426 1017 447 ne
rect 1017 439 1057 447
tri 1057 439 1078 460 sw
rect 1017 426 1078 439
tri 1017 425 1018 426 ne
rect 1018 425 1078 426
tri 1018 417 1026 425 ne
rect 1026 363 1078 425
tri 1078 363 1083 368 sw
rect 282 328 402 337
rect 282 294 294 328
rect 328 294 385 328
rect 282 285 402 294
rect 454 285 466 337
rect 518 285 524 337
rect 1026 334 1083 363
tri 1083 334 1112 363 sw
rect 1026 328 1672 334
rect 1026 294 1038 328
rect 1072 294 1112 328
rect 1146 294 1186 328
rect 1220 294 1260 328
rect 1294 294 1334 328
rect 1368 294 1407 328
rect 1441 294 1480 328
rect 1514 294 1553 328
rect 1587 294 1626 328
rect 1660 294 1672 328
rect 1026 288 1672 294
tri 1908 251 1935 278 se
rect 1935 256 1987 645
tri 1987 626 2021 660 nw
tri 2770 628 2802 660 se
rect 2802 629 2863 660
tri 2863 629 2953 719 sw
rect 2802 628 2953 629
tri 2413 626 2415 628 se
rect 2415 626 2953 628
tri 2403 616 2413 626 se
rect 2413 616 2953 626
tri 2391 604 2403 616 se
rect 2403 604 2756 616
tri 2357 570 2391 604 se
rect 2391 570 2637 604
rect 2671 582 2756 604
rect 2790 582 2953 616
rect 2671 570 2953 582
tri 2330 543 2357 570 se
rect 2357 543 2953 570
tri 2319 532 2330 543 se
rect 2330 532 2756 543
rect 1935 251 1982 256
tri 1982 251 1987 256 nw
tri 2304 517 2319 532 se
rect 2319 517 2637 532
rect 2304 498 2637 517
rect 2671 509 2756 532
rect 2790 509 2953 543
rect 2671 498 2953 509
rect 2304 470 2953 498
rect 2304 460 2756 470
rect 2304 426 2637 460
rect 2671 436 2756 460
rect 2790 436 2953 470
rect 2671 426 2953 436
rect 2304 397 2953 426
rect 2304 363 2756 397
rect 2790 363 2953 397
rect 2304 324 2953 363
rect 2304 290 2756 324
rect 2790 290 2953 324
rect 2304 251 2953 290
tri 1891 234 1908 251 se
rect 1908 234 1965 251
tri 1965 234 1982 251 nw
rect 2304 234 2756 251
tri 1879 222 1891 234 se
rect 1891 222 1953 234
tri 1953 222 1965 234 nw
tri 1857 200 1879 222 se
rect 1879 200 1931 222
tri 1931 200 1953 222 nw
rect 2304 200 2637 234
rect 2671 217 2756 234
rect 2790 217 2953 251
rect 2671 200 2953 217
rect 27 148 33 200
rect 85 148 97 200
rect 149 148 886 200
rect 938 148 950 200
rect 1002 177 1908 200
tri 1908 177 1931 200 nw
rect 2304 177 2953 200
rect 1002 162 1893 177
tri 1893 162 1908 177 nw
rect 2304 162 2756 177
rect 1002 148 1879 162
tri 1879 148 1893 162 nw
rect 2304 128 2637 162
rect 2671 143 2756 162
rect 2790 143 2953 177
rect 2671 128 2953 143
rect 2304 103 2953 128
rect 2304 90 2756 103
rect 2304 56 2637 90
rect 2671 69 2756 90
rect 2790 69 2953 103
rect 2671 56 2953 69
rect 2304 13 2953 56
tri 2651 -42 2706 13 ne
rect 2706 -42 2953 13
rect 1048 -94 1054 -42
rect 1106 -94 1118 -42
rect 1170 -62 1985 -42
tri 1985 -62 2005 -42 sw
tri 2706 -62 2726 -42 ne
rect 2726 -62 2953 -42
rect 1170 -68 2354 -62
rect 1170 -94 1968 -68
tri 1942 -102 1950 -94 ne
rect 1950 -102 1968 -94
rect 2002 -102 2053 -68
rect 2087 -102 2138 -68
rect 2172 -102 2223 -68
rect 2257 -102 2308 -68
rect 2342 -102 2354 -68
tri 1950 -108 1956 -102 ne
rect 1956 -108 2354 -102
tri 2726 -108 2772 -62 ne
rect 2772 -108 2953 -62
tri 2772 -155 2819 -108 ne
rect 2819 -155 2953 -108
rect 1905 -177 1951 -165
tri 1197 -189 1204 -182 se
rect 1204 -189 1210 -182
rect 1006 -195 1210 -189
rect 1262 -195 1274 -182
rect 1326 -189 1332 -182
tri 1332 -189 1339 -182 sw
rect 1326 -195 1548 -189
rect 916 -232 968 -226
rect 1006 -229 1018 -195
rect 1052 -229 1098 -195
rect 1132 -229 1178 -195
rect 1326 -229 1340 -195
rect 1374 -229 1421 -195
rect 1455 -229 1502 -195
rect 1536 -229 1548 -195
rect 1905 -211 1911 -177
rect 1945 -211 1951 -177
rect 2321 -207 2327 -155
rect 2379 -207 2391 -155
rect 2443 -158 2449 -155
tri 2449 -158 2452 -155 sw
tri 2819 -156 2820 -155 ne
rect 2443 -204 2452 -158
rect 2443 -207 2449 -204
tri 2449 -207 2452 -204 nw
rect 1006 -234 1210 -229
rect 1262 -234 1274 -229
rect 1326 -234 1548 -229
rect 1006 -235 1548 -234
tri 1882 -235 1905 -212 se
rect 1905 -235 1951 -211
tri 1845 -272 1882 -235 se
rect 1882 -272 1951 -235
rect 916 -296 968 -284
rect 1404 -324 1410 -272
rect 1462 -324 1474 -272
rect 1526 -305 1951 -272
rect 1526 -324 1911 -305
tri 1879 -339 1894 -324 ne
rect 1894 -339 1911 -324
rect 1945 -339 1951 -305
rect 916 -354 968 -348
tri 1894 -350 1905 -339 ne
rect 1905 -351 1951 -339
tri 920 -356 922 -354 ne
rect 922 -356 968 -354
tri 1398 -365 1404 -359 se
rect 1404 -365 1410 -359
rect 1006 -371 1410 -365
rect 1006 -405 1018 -371
rect 1052 -405 1096 -371
rect 1130 -405 1174 -371
rect 1208 -405 1252 -371
rect 1286 -405 1330 -371
rect 1364 -405 1408 -371
rect 1006 -411 1410 -405
rect 1462 -411 1474 -359
rect 1526 -365 1532 -359
tri 1532 -365 1538 -359 sw
rect 1526 -371 1610 -365
rect 1526 -405 1564 -371
rect 1598 -405 1610 -371
rect 1526 -411 1610 -405
rect 771 -422 968 -416
rect 823 -428 968 -422
rect 823 -462 928 -428
rect 962 -462 968 -428
tri 1641 -442 1647 -436 se
rect 1647 -442 2736 -436
tri 1630 -453 1641 -442 se
rect 1641 -453 1894 -442
rect 823 -474 968 -462
rect 771 -486 968 -474
rect 823 -500 968 -486
rect 823 -534 928 -500
rect 962 -534 968 -500
rect 1204 -505 1210 -453
rect 1262 -505 1274 -453
rect 1326 -476 1894 -453
rect 1928 -476 1967 -442
rect 2001 -476 2040 -442
rect 2074 -476 2113 -442
rect 2147 -476 2186 -442
rect 2220 -476 2258 -442
rect 2292 -476 2330 -442
rect 2364 -476 2402 -442
rect 2436 -476 2474 -442
rect 2508 -476 2546 -442
rect 2580 -476 2618 -442
rect 2652 -476 2690 -442
rect 2724 -476 2736 -442
rect 1326 -482 2736 -476
rect 1326 -505 1644 -482
tri 1644 -505 1667 -482 nw
rect 823 -538 968 -534
rect 1849 -523 1901 -517
tri 1901 -525 1909 -517 sw
rect 1901 -531 2694 -525
rect 771 -546 968 -538
tri 1043 -541 1048 -536 se
rect 1048 -541 1054 -536
rect 1006 -547 1054 -541
rect 1106 -547 1118 -536
rect 1170 -541 1176 -536
tri 1176 -541 1181 -536 sw
rect 1170 -547 1603 -541
rect 1006 -581 1018 -547
rect 1052 -581 1054 -547
rect 1170 -581 1172 -547
rect 1206 -581 1249 -547
rect 1283 -581 1326 -547
rect 1360 -581 1403 -547
rect 1437 -581 1480 -547
rect 1514 -581 1557 -547
rect 1591 -581 1603 -547
rect 1006 -587 1054 -581
tri 1047 -588 1048 -587 ne
rect 1048 -588 1054 -587
rect 1106 -588 1118 -581
rect 1170 -587 1603 -581
rect 1901 -565 1941 -531
rect 1975 -565 2576 -531
rect 2610 -565 2648 -531
rect 2682 -565 2694 -531
rect 1901 -568 2694 -565
tri 2781 -568 2820 -529 se
rect 2820 -568 2953 -155
rect 1901 -571 1987 -568
tri 1987 -571 1990 -568 nw
tri 2561 -571 2564 -568 ne
rect 2564 -571 2694 -568
tri 2778 -571 2781 -568 se
rect 2781 -571 2953 -568
rect 1849 -587 1901 -575
rect 1170 -588 1176 -587
tri 1176 -588 1177 -587 nw
tri 1901 -599 1929 -571 nw
tri 2750 -599 2778 -571 se
rect 2778 -599 2953 -571
tri 2749 -600 2750 -599 se
rect 2750 -600 2953 -599
rect 1849 -645 1901 -639
tri 2223 -640 2246 -617 se
rect 2246 -640 2252 -600
tri 2218 -645 2223 -640 se
rect 2223 -645 2252 -640
tri 2186 -677 2218 -645 se
rect 2218 -652 2252 -645
rect 2304 -652 2318 -600
rect 2370 -652 2376 -600
tri 2723 -626 2749 -600 se
rect 2749 -626 2953 -600
rect 2218 -676 2376 -652
tri 2376 -676 2426 -626 sw
tri 2673 -676 2723 -626 se
rect 2723 -676 2953 -626
rect 2218 -677 2953 -676
tri 1356 -725 1404 -677 se
rect 1404 -701 2953 -677
rect 1404 -753 1410 -701
rect 1462 -753 1474 -701
rect 1526 -753 2953 -701
rect 1404 -778 2953 -753
<< via1 >>
rect -443 5952 -391 6004
rect -443 5875 -391 5927
rect -181 5869 -129 5921
rect -104 5869 -52 5921
rect 30 5869 82 5921
rect 107 5869 159 5921
rect -104 5763 -52 5815
rect -33 5763 19 5815
rect 38 5763 90 5815
rect -104 5608 -52 5660
rect -33 5608 19 5660
rect 38 5608 90 5660
rect 470 5554 522 5606
rect 559 5554 611 5606
rect 402 5517 454 5526
rect 402 5483 408 5517
rect 408 5483 442 5517
rect 442 5483 454 5517
rect 402 5474 454 5483
rect 466 5474 518 5526
rect 858 5517 910 5526
rect 858 5483 864 5517
rect 864 5483 898 5517
rect 898 5483 910 5517
rect 858 5474 910 5483
rect 922 5517 974 5526
rect 922 5483 947 5517
rect 947 5483 974 5517
rect 922 5474 974 5483
rect 771 5380 823 5432
rect 27 5207 39 5224
rect 39 5207 73 5224
rect 73 5207 79 5224
rect 27 5172 79 5207
rect 27 5148 79 5160
rect 27 5114 39 5148
rect 39 5114 73 5148
rect 73 5114 79 5148
rect 27 5108 79 5114
rect 771 5316 823 5368
rect 1054 4510 1106 4562
rect 1118 4510 1170 4562
rect 27 4391 79 4443
rect 27 4327 79 4379
rect 1204 4389 1256 4441
rect 771 4309 823 4361
rect 1204 4325 1256 4377
rect 771 4245 823 4297
rect 852 4216 904 4268
rect 852 4152 904 4204
rect 396 4062 405 4087
rect 405 4062 439 4087
rect 439 4062 448 4087
rect 396 4035 448 4062
rect 1287 4172 1293 4182
rect 1293 4172 1327 4182
rect 1327 4172 1339 4182
rect 1287 4130 1339 4172
rect 1287 4106 1339 4118
rect 1287 4072 1293 4106
rect 1293 4072 1327 4106
rect 1327 4072 1339 4106
rect 1287 4066 1339 4072
rect 1636 4154 1645 4182
rect 1645 4154 1679 4182
rect 1679 4154 1688 4182
rect 1636 4130 1688 4154
rect 1636 4106 1688 4118
rect 1636 4072 1645 4106
rect 1645 4072 1679 4106
rect 1679 4072 1688 4106
rect 1636 4066 1688 4072
rect 396 3990 405 4023
rect 405 3990 439 4023
rect 439 3990 448 4023
rect 396 3971 448 3990
rect 858 942 910 994
rect 922 942 974 994
rect 2385 934 2437 940
rect 2385 900 2394 934
rect 2394 900 2428 934
rect 2428 900 2437 934
rect 2385 888 2437 900
rect 2385 862 2437 876
rect 2385 828 2394 862
rect 2394 828 2428 862
rect 2428 828 2437 862
rect 406 772 458 824
rect 470 772 522 824
rect 2385 824 2437 828
rect 858 700 910 709
rect 858 666 867 700
rect 867 666 910 700
rect 858 657 910 666
rect 922 700 974 709
rect 922 666 924 700
rect 924 666 958 700
rect 958 666 974 700
rect 922 657 974 666
rect 1865 700 1917 706
rect 1929 700 1981 706
rect 1865 666 1875 700
rect 1875 666 1914 700
rect 1914 666 1917 700
rect 1929 666 1948 700
rect 1948 666 1981 700
rect 1865 654 1917 666
rect 1929 654 1981 666
rect 771 517 823 569
rect 771 453 823 505
rect 402 328 454 337
rect 402 294 419 328
rect 419 294 454 328
rect 402 285 454 294
rect 466 328 518 337
rect 466 294 476 328
rect 476 294 510 328
rect 510 294 518 328
rect 466 285 518 294
rect 33 192 85 200
rect 33 158 42 192
rect 42 158 76 192
rect 76 158 85 192
rect 33 148 85 158
rect 97 192 149 200
rect 97 158 114 192
rect 114 158 148 192
rect 148 158 149 192
rect 97 148 149 158
rect 886 148 938 200
rect 950 148 1002 200
rect 1054 -94 1106 -42
rect 1118 -94 1170 -42
rect 1210 -195 1262 -182
rect 1274 -195 1326 -182
rect 916 -238 968 -232
rect 1210 -229 1212 -195
rect 1212 -229 1259 -195
rect 1259 -229 1262 -195
rect 1274 -229 1293 -195
rect 1293 -229 1326 -195
rect 2327 -164 2379 -155
rect 2327 -198 2334 -164
rect 2334 -198 2368 -164
rect 2368 -198 2379 -164
rect 2327 -207 2379 -198
rect 2391 -164 2443 -155
rect 2391 -198 2406 -164
rect 2406 -198 2440 -164
rect 2440 -198 2443 -164
rect 2391 -207 2443 -198
rect 1210 -234 1262 -229
rect 1274 -234 1326 -229
rect 916 -272 928 -238
rect 928 -272 962 -238
rect 962 -272 968 -238
rect 916 -284 968 -272
rect 916 -310 968 -296
rect 916 -344 928 -310
rect 928 -344 962 -310
rect 962 -344 968 -310
rect 1410 -324 1462 -272
rect 1474 -324 1526 -272
rect 916 -348 968 -344
rect 1410 -371 1462 -359
rect 1410 -405 1442 -371
rect 1442 -405 1462 -371
rect 1410 -411 1462 -405
rect 1474 -371 1526 -359
rect 1474 -405 1486 -371
rect 1486 -405 1520 -371
rect 1520 -405 1526 -371
rect 1474 -411 1526 -405
rect 771 -474 823 -422
rect 771 -538 823 -486
rect 1210 -505 1262 -453
rect 1274 -505 1326 -453
rect 1849 -531 1901 -523
rect 1054 -547 1106 -536
rect 1118 -547 1170 -536
rect 1054 -581 1095 -547
rect 1095 -581 1106 -547
rect 1118 -581 1129 -547
rect 1129 -581 1170 -547
rect 1054 -588 1106 -581
rect 1118 -588 1170 -581
rect 1849 -565 1861 -531
rect 1861 -565 1895 -531
rect 1895 -565 1901 -531
rect 1849 -575 1901 -565
rect 1849 -639 1901 -587
rect 2252 -606 2304 -600
rect 2252 -640 2258 -606
rect 2258 -640 2292 -606
rect 2292 -640 2304 -606
rect 2252 -652 2304 -640
rect 2318 -606 2370 -600
rect 2318 -640 2330 -606
rect 2330 -640 2364 -606
rect 2364 -640 2370 -606
rect 2318 -652 2370 -640
rect 1410 -753 1462 -701
rect 1474 -753 1526 -701
<< metal2 >>
rect -443 6004 -391 6010
rect -443 5927 -391 5952
rect -443 5869 -391 5875
rect -187 5869 -181 5921
rect -129 5869 -104 5921
rect -52 5869 -46 5921
rect 24 5869 30 5921
rect 82 5869 107 5921
rect 159 5869 165 5921
tri -144 5835 -110 5869 ne
rect -110 5815 -46 5869
tri -46 5815 -12 5849 sw
rect -110 5763 -104 5815
rect -52 5763 -33 5815
rect 19 5763 38 5815
rect 90 5763 96 5815
tri -78 5729 -44 5763 ne
tri -78 5660 -44 5694 se
rect -44 5660 16 5763
tri 16 5729 50 5763 nw
tri 16 5660 50 5694 sw
tri 96 5660 125 5689 se
rect 125 5660 796 5689
rect -110 5608 -104 5660
rect -52 5608 -33 5660
rect 19 5608 38 5660
rect 90 5655 796 5660
tri 796 5655 830 5689 sw
rect 90 5637 830 5655
rect 90 5608 162 5637
tri 162 5608 191 5637 nw
tri 774 5608 803 5637 ne
rect 803 5608 830 5637
tri 803 5606 805 5608 ne
rect 805 5606 830 5608
rect 464 5554 470 5606
rect 522 5554 559 5606
rect 611 5572 715 5606
tri 715 5572 749 5606 sw
tri 805 5581 830 5606 ne
tri 830 5581 904 5655 sw
tri 830 5572 839 5581 ne
rect 839 5572 904 5581
rect 611 5554 749 5572
tri 693 5526 721 5554 ne
rect 721 5526 749 5554
tri 749 5526 795 5572 sw
tri 839 5559 852 5572 ne
rect 852 5526 904 5572
tri 904 5526 938 5560 sw
rect 396 5474 402 5526
rect 454 5474 466 5526
rect 518 5474 524 5526
tri 721 5498 749 5526 ne
rect 749 5498 795 5526
tri 795 5498 823 5526 sw
tri 749 5476 771 5498 ne
rect 27 5224 79 5230
rect 27 5160 79 5172
rect 27 4443 79 5108
rect 27 4379 79 4391
rect 27 200 79 4327
rect 396 4087 448 5474
tri 448 5440 482 5474 nw
rect 396 4023 448 4035
rect 396 824 448 3971
rect 771 5432 823 5498
rect 771 5368 823 5380
rect 771 4361 823 5316
rect 771 4297 823 4309
tri 448 824 482 858 sw
rect 396 772 406 824
rect 458 772 470 824
rect 522 772 528 824
rect 396 337 448 772
tri 448 738 482 772 nw
rect 771 569 823 4245
rect 852 5474 858 5526
rect 910 5474 922 5526
rect 974 5474 980 5526
rect 852 4268 904 5474
tri 904 5440 938 5474 nw
rect 1048 4510 1054 4562
rect 1106 4510 1118 4562
rect 1170 4510 1176 4562
tri 1090 4476 1124 4510 ne
rect 852 4204 904 4216
rect 852 994 904 4152
tri 904 994 938 1028 sw
rect 852 942 858 994
rect 910 942 922 994
rect 974 942 980 994
rect 852 940 936 942
tri 936 940 938 942 nw
rect 852 709 904 940
tri 904 908 936 940 nw
tri 904 709 938 743 sw
rect 852 657 858 709
rect 910 657 922 709
rect 974 657 980 709
rect 771 505 823 517
tri 448 337 482 371 sw
rect 396 285 402 337
rect 454 285 466 337
rect 518 285 524 337
tri 79 200 113 234 sw
rect 27 148 33 200
rect 85 148 97 200
rect 149 148 155 200
rect 771 -422 823 453
rect 880 148 886 200
rect 938 148 950 200
rect 1002 148 1008 200
tri 880 112 916 148 ne
rect 916 -232 968 148
tri 968 108 1008 148 nw
tri 1080 -42 1124 2 se
rect 1124 -42 1176 4510
rect 1048 -94 1054 -42
rect 1106 -94 1118 -42
rect 1170 -94 1176 -42
tri 1080 -138 1124 -94 ne
rect 916 -296 968 -284
rect 916 -356 968 -348
rect 771 -486 823 -474
tri 1121 -505 1124 -502 se
rect 1124 -505 1176 -94
rect 1204 4441 1256 4447
rect 1204 4377 1256 4389
rect 1204 -155 1256 4325
rect 1284 4182 1339 5975
rect 1284 4130 1287 4182
rect 1284 4118 1339 4130
rect 1284 4066 1287 4118
rect 1284 965 1339 4066
rect 1636 4182 1688 5974
rect 1636 4118 1688 4130
tri 1284 940 1309 965 ne
rect 1309 940 1339 965
tri 1339 940 1383 984 sw
tri 1309 910 1339 940 ne
rect 1339 939 1383 940
tri 1383 939 1384 940 sw
rect 1339 910 1384 939
tri 1339 888 1361 910 ne
rect 1361 888 1384 910
tri 1384 888 1435 939 sw
tri 1361 876 1373 888 ne
rect 1373 876 1435 888
tri 1435 876 1447 888 sw
tri 1373 865 1384 876 ne
rect 1384 865 1447 876
tri 1447 865 1458 876 sw
tri 1384 845 1404 865 ne
tri 1256 -155 1262 -149 sw
rect 1204 -182 1262 -155
tri 1262 -182 1289 -155 sw
rect 1204 -234 1210 -182
rect 1262 -234 1274 -182
rect 1326 -234 1332 -182
rect 1404 -207 1459 865
tri 1459 -207 1467 -199 sw
rect 1204 -411 1256 -234
tri 1256 -267 1289 -234 nw
rect 1404 -272 1467 -207
tri 1467 -272 1532 -207 sw
rect 1404 -324 1410 -272
rect 1462 -324 1474 -272
rect 1526 -324 1532 -272
tri 1256 -411 1290 -377 sw
rect 1404 -411 1410 -359
rect 1462 -411 1474 -359
rect 1526 -411 1532 -359
rect 1204 -453 1290 -411
tri 1290 -453 1332 -411 sw
rect 1204 -505 1210 -453
rect 1262 -505 1274 -453
rect 1326 -505 1332 -453
tri 1103 -523 1121 -505 se
rect 1121 -523 1176 -505
tri 1090 -536 1103 -523 se
rect 1103 -536 1176 -523
rect 771 -544 823 -538
rect 1048 -588 1054 -536
rect 1106 -588 1118 -536
rect 1170 -588 1176 -536
rect 1404 -701 1532 -411
rect 1636 -517 1688 4066
rect 2385 940 2437 946
rect 2385 876 2437 888
rect 2385 818 2437 824
rect 1859 654 1865 706
rect 1917 654 1929 706
rect 1981 654 1987 706
rect 2246 -207 2327 -155
rect 2379 -207 2391 -155
rect 2443 -207 2449 -155
tri 1688 -517 1714 -491 sw
rect 1636 -523 1901 -517
rect 1636 -575 1849 -523
rect 1636 -587 1901 -575
rect 1636 -639 1849 -587
rect 1636 -645 1901 -639
rect 2246 -600 2376 -207
tri 2376 -257 2426 -207 nw
rect 2246 -652 2252 -600
rect 2304 -652 2318 -600
rect 2370 -652 2376 -600
rect 2246 -662 2376 -652
rect 1404 -753 1410 -701
rect 1462 -753 1474 -701
rect 1526 -753 1532 -701
rect 1404 -778 1532 -753
<< comment >>
tri -86 6068 -81 6069 se
tri -81 6068 -76 6069 sw
tri 46 6068 51 6069 se
tri 51 6068 56 6069 sw
tri -90 6065 -86 6068 se
rect -86 6065 -76 6068
tri -76 6065 -71 6068 sw
tri 41 6065 46 6068 se
rect 46 6065 56 6068
tri 56 6065 61 6068 sw
tri -95 6060 -90 6065 se
rect -90 6060 -71 6065
tri -71 6060 -67 6065 sw
tri 37 6060 41 6065 se
rect 41 6060 61 6065
tri 61 6060 65 6065 sw
tri -100 6052 -95 6060 se
rect -95 6052 -67 6060
tri -67 6052 -62 6060 sw
tri 32 6052 37 6060 se
rect 37 6052 65 6060
tri 65 6052 70 6060 sw
tri -104 6043 -100 6052 se
rect -100 6043 -62 6052
tri -62 6043 -58 6052 sw
tri 28 6043 32 6052 se
rect 32 6043 70 6052
tri 70 6043 74 6052 sw
tri -108 6032 -104 6043 se
rect -104 6032 -58 6043
tri -58 6032 -54 6043 sw
tri 24 6032 28 6043 se
rect 28 6032 74 6043
tri 74 6032 78 6043 sw
tri -112 6019 -108 6032 se
rect -108 6019 -54 6032
tri -54 6019 -50 6032 sw
tri 20 6019 24 6032 se
rect 24 6019 78 6032
tri 78 6019 82 6032 sw
tri -115 6005 -112 6019 se
rect -112 6005 -50 6019
tri -50 6005 -46 6019 sw
tri 16 6005 20 6019 se
rect 20 6005 82 6019
tri 82 6005 86 6019 sw
tri -119 5989 -115 6005 se
rect -115 5989 -46 6005
tri -46 5989 -43 6005 sw
tri 13 5989 16 6005 se
rect 16 5989 86 6005
tri 86 5989 89 6005 sw
tri -122 5972 -119 5989 se
rect -119 5972 -43 5989
tri -43 5972 -40 5989 sw
tri 10 5972 13 5989 se
rect 13 5972 89 5989
tri 89 5972 92 5989 sw
tri -124 5953 -122 5972 se
rect -122 5953 -40 5972
tri -40 5953 -38 5972 sw
tri 8 5953 10 5972 se
rect 10 5953 92 5972
tri 92 5953 94 5972 sw
tri -126 5934 -124 5953 se
rect -124 5934 -38 5953
tri -38 5934 -36 5953 sw
tri 6 5934 8 5953 se
rect 8 5934 94 5953
tri 94 5934 96 5953 sw
tri -128 5914 -126 5934 se
rect -126 5914 -36 5934
tri -36 5914 -34 5934 sw
tri 4 5914 6 5934 se
rect 6 5914 96 5934
tri 96 5914 98 5934 sw
tri -129 5893 -128 5914 se
rect -128 5893 -34 5914
tri -34 5893 -33 5914 sw
tri 3 5893 4 5914 se
rect 4 5893 98 5914
tri 98 5893 99 5914 sw
tri -130 5872 -129 5893 se
rect -129 5872 -33 5893
tri -33 5872 -32 5893 sw
rect -130 5829 -32 5872
tri -130 5808 -129 5829 ne
rect -129 5808 -33 5829
tri -33 5808 -32 5829 nw
tri 2 5872 3 5893 se
rect 3 5872 99 5893
tri 99 5872 100 5893 sw
rect 2 5829 100 5872
tri 2 5808 3 5829 ne
rect 3 5808 99 5829
tri 99 5808 100 5829 nw
tri -129 5787 -128 5808 ne
rect -128 5787 -34 5808
tri -34 5787 -33 5808 nw
tri 3 5787 4 5808 ne
rect 4 5787 98 5808
tri 98 5787 99 5808 nw
tri -128 5767 -126 5787 ne
rect -126 5767 -36 5787
tri -36 5767 -34 5787 nw
tri 4 5767 6 5787 ne
rect 6 5767 96 5787
tri 96 5767 98 5787 nw
tri -126 5747 -124 5767 ne
rect -124 5747 -38 5767
tri -38 5747 -36 5767 nw
tri 6 5747 8 5767 ne
rect 8 5747 94 5767
tri 94 5747 96 5767 nw
tri -124 5729 -122 5747 ne
rect -122 5729 -40 5747
tri -40 5729 -38 5747 nw
tri 8 5729 10 5747 ne
rect 10 5729 92 5747
tri 92 5729 94 5747 nw
tri -122 5712 -119 5729 ne
rect -119 5712 -43 5729
tri -43 5712 -40 5729 nw
tri 10 5712 13 5729 ne
rect 13 5712 89 5729
tri 89 5712 92 5729 nw
tri -119 5696 -115 5712 ne
rect -115 5696 -46 5712
tri -46 5696 -43 5712 nw
tri 13 5696 16 5712 ne
rect 16 5696 86 5712
tri 86 5696 89 5712 nw
tri -115 5681 -112 5696 ne
rect -112 5681 -50 5696
tri -50 5681 -46 5696 nw
tri 16 5681 20 5696 ne
rect 20 5681 82 5696
tri 82 5681 86 5696 nw
tri -112 5669 -108 5681 ne
rect -108 5669 -54 5681
tri -54 5669 -50 5681 nw
tri 20 5669 24 5681 ne
rect 24 5669 78 5681
tri 78 5669 82 5681 nw
tri -108 5658 -104 5669 ne
rect -104 5658 -58 5669
tri -58 5658 -54 5669 nw
tri 24 5658 28 5669 ne
rect 28 5658 74 5669
tri 74 5658 78 5669 nw
tri -104 5648 -100 5658 ne
rect -100 5648 -62 5658
tri -62 5648 -58 5658 nw
tri 28 5648 32 5658 ne
rect 32 5648 70 5658
tri 70 5648 74 5658 nw
tri -100 5641 -95 5648 ne
rect -95 5641 -67 5648
tri -67 5641 -62 5648 nw
tri 32 5641 37 5648 ne
rect 37 5641 65 5648
tri 65 5641 70 5648 nw
tri -95 5636 -90 5641 ne
rect -90 5636 -71 5641
tri -71 5636 -67 5641 nw
tri 37 5636 41 5641 ne
rect 41 5636 61 5641
tri 61 5636 65 5641 nw
tri -90 5633 -86 5636 ne
rect -86 5633 -76 5636
tri -76 5633 -71 5636 nw
tri 41 5633 46 5636 ne
rect 46 5633 56 5636
tri 56 5633 61 5636 nw
tri -86 5632 -81 5633 ne
tri -81 5632 -76 5633 nw
tri 46 5632 51 5633 ne
tri 51 5632 56 5633 nw
use nfet_CDNS_5246887918540  nfet_CDNS_5246887918540_0
timestamp 1704896540
transform 0 1 2476 1 0 816
box -79 -32 199 232
use nfet_CDNS_5246887918541  nfet_CDNS_5246887918541_0
timestamp 1704896540
transform 0 1 1010 -1 0 -416
box -79 -32 199 632
use nfet_CDNS_5246887918541  nfet_CDNS_5246887918541_1
timestamp 1704896540
transform 0 1 1010 -1 0 -240
box -79 -32 199 632
use nfet_CDNS_52468879185481  nfet_CDNS_52468879185481_0
timestamp 1704896540
transform 1 0 1026 0 1 418
box -79 -32 1679 232
use nfet_CDNS_52468879185481  nfet_CDNS_52468879185481_1
timestamp 1704896540
transform 1 0 1026 0 1 46
box -79 -32 1679 232
use nfet_CDNS_52468879185482  nfet_CDNS_52468879185482_0
timestamp 1704896540
transform 1 0 170 0 1 418
box -79 -32 879 232
use nfet_CDNS_52468879185482  nfet_CDNS_52468879185482_1
timestamp 1704896540
transform 1 0 170 0 1 46
box -79 -32 879 232
use nfet_CDNS_52468879185483  nfet_CDNS_52468879185483_0
timestamp 1704896540
transform -1 0 2762 0 -1 -524
box -79 -32 935 116
use nfet_CDNS_52468879185484  nfet_CDNS_52468879185484_0
timestamp 1704896540
transform -1 0 2356 0 -1 -152
box -79 -32 479 116
use pfet_CDNS_5246887918533  pfet_CDNS_5246887918533_0
timestamp 1704896540
transform -1 0 1458 0 -1 4468
box -119 -66 415 666
use pfet_CDNS_5246887918536  pfet_CDNS_5246887918536_0
timestamp 1704896540
transform -1 0 1634 0 -1 4468
box -119 -66 239 666
use pfet_CDNS_52468879185664  pfet_CDNS_52468879185664_0
timestamp 1704896540
transform -1 0 570 0 -1 4104
box -119 -66 415 266
use pfet_CDNS_52468879185692  pfet_CDNS_52468879185692_0
timestamp 1704896540
transform -1 0 570 0 -1 4549
box -119 -66 415 206
use pfet_CDNS_524688791851448  pfet_CDNS_524688791851448_0
timestamp 1704896540
transform -1 0 1820 0 -1 5434
box -119 -66 2111 666
<< labels >>
flabel comment s 52 5542 52 5542 0 FreeSans 400 0 0 0 padlo
flabel comment s 52 5850 52 5850 0 FreeSans 400 90 0 0 ModA7B
flabel comment s -81 5850 -81 5850 0 FreeSans 400 90 0 0 ModA7
flabel comment s 590 153 590 153 0 FreeSans 1000 0 0 0 I51
flabel comment s 1766 153 1766 153 0 FreeSans 1000 0 0 0 I52
flabel comment s 590 531 590 531 0 FreeSans 1000 0 0 0 I69
flabel comment s 1754 531 1754 531 0 FreeSans 1000 0 0 0 I67
flabel comment s 1065 5245 1065 5245 0 FreeSans 600 0 0 0 I64
flabel comment s 562 5245 562 5245 0 FreeSans 600 0 0 0 I49
flabel comment s 1696 5245 1696 5245 0 FreeSans 600 0 0 0 I65
flabel comment s 56 5245 56 5245 0 FreeSans 600 0 0 0 I50
flabel comment s 562 4492 562 4492 0 FreeSans 600 0 0 0 I72
flabel comment s 1330 4492 1330 4492 0 FreeSans 600 0 0 0 I76
flabel comment s 1571 4492 1571 4492 0 FreeSans 600 0 0 0 I77
flabel comment s 329 4492 329 4492 0 FreeSans 600 0 0 0 I70
flabel comment s 434 4044 434 4044 0 FreeSans 600 0 0 0 I53
flabel metal1 s 2560 82 2950 546 0 FreeSans 600 0 0 0 vgnd
port 3 nsew
flabel metal1 s 1824 3889 2240 4002 0 FreeSans 600 0 0 0 vpwr
port 2 nsew
flabel metal2 s 1284 5915 1336 5974 0 FreeSans 200 0 0 0 p1g
port 4 nsew
flabel metal2 s 1636 5915 1688 5974 0 FreeSans 200 0 0 0 p2g
port 5 nsew
flabel metal2 s 108 5608 157 5660 0 FreeSans 200 0 0 0 padlo
port 6 nsew
<< properties >>
string GDS_END 89370560
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89254692
string path 30.750 107.975 30.750 111.175 
<< end >>
