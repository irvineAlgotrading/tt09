magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 217 607 711 1249
<< pwell >>
rect 286 -11 811 143
<< psubdiff >>
rect 312 83 785 117
rect 312 49 346 83
rect 380 49 421 83
rect 455 49 495 83
rect 529 49 569 83
rect 603 49 643 83
rect 677 49 717 83
rect 751 49 785 83
rect 312 15 785 49
<< psubdiffcont >>
rect 346 49 380 83
rect 421 49 455 83
rect 495 49 529 83
rect 569 49 603 83
rect 643 49 677 83
rect 717 49 751 83
<< poly >>
rect 336 595 612 611
rect 92 461 128 581
rect 336 561 352 595
rect 386 561 422 595
rect 456 561 492 595
rect 526 561 562 595
rect 596 561 612 595
rect 336 545 612 561
rect 37 445 428 461
rect 37 411 53 445
rect 87 411 121 445
rect 155 425 428 445
rect 155 411 171 425
rect 392 411 428 425
rect 484 411 520 545
rect 576 411 612 545
rect 800 533 836 581
rect 702 517 836 533
rect 702 503 718 517
rect 668 483 718 503
rect 752 483 786 517
rect 820 483 836 517
rect 668 467 836 483
rect 668 411 704 467
rect 37 395 171 411
<< polycont >>
rect 352 561 386 595
rect 422 561 456 595
rect 492 561 526 595
rect 562 561 596 595
rect 53 411 87 445
rect 121 411 155 445
rect 718 483 752 517
rect 786 483 820 517
<< locali >>
rect 24 517 102 1217
rect 139 787 325 1247
rect 447 947 481 985
rect 173 753 215 787
rect 249 753 291 787
rect 139 709 325 753
rect 173 675 215 709
rect 249 675 291 709
rect 603 787 789 1247
rect 637 753 679 787
rect 713 753 755 787
rect 603 709 789 753
rect 637 675 679 709
rect 713 675 755 709
rect 336 561 352 595
rect 412 561 422 595
rect 484 561 492 595
rect 526 561 562 595
rect 596 561 612 595
rect 58 483 96 517
rect 438 483 476 517
rect 702 483 716 517
rect 752 483 786 517
rect 822 483 836 517
rect 37 411 53 445
rect 87 411 121 445
rect 155 411 171 445
rect 339 199 392 377
rect 339 165 347 199
rect 381 165 392 199
rect 428 175 484 483
rect 521 199 574 377
rect 623 289 657 327
rect 339 117 392 165
rect 521 165 531 199
rect 565 165 574 199
rect 521 117 574 165
rect 704 199 757 377
rect 872 361 923 1217
rect 872 327 878 361
rect 912 327 923 361
rect 872 289 923 327
rect 872 255 878 289
rect 912 255 923 289
rect 872 243 923 255
rect 704 165 713 199
rect 747 165 757 199
rect 704 117 757 165
rect 312 83 785 117
rect 312 49 346 83
rect 380 73 421 83
rect 381 49 421 73
rect 455 49 495 83
rect 529 73 569 83
rect 529 49 531 73
rect 312 39 347 49
rect 381 39 531 49
rect 565 49 569 73
rect 603 49 643 83
rect 677 73 717 83
rect 677 49 713 73
rect 751 49 785 83
rect 565 39 713 49
rect 747 39 785 49
rect 312 15 785 39
<< viali >>
rect 447 985 481 1019
rect 447 913 481 947
rect 139 753 173 787
rect 215 753 249 787
rect 291 753 325 787
rect 139 675 173 709
rect 215 675 249 709
rect 291 675 325 709
rect 603 753 637 787
rect 679 753 713 787
rect 755 753 789 787
rect 603 675 637 709
rect 679 675 713 709
rect 755 675 789 709
rect 378 561 386 595
rect 386 561 412 595
rect 450 561 456 595
rect 456 561 484 595
rect 24 483 58 517
rect 96 483 130 517
rect 404 483 438 517
rect 476 483 510 517
rect 716 483 718 517
rect 718 483 750 517
rect 788 483 820 517
rect 820 483 822 517
rect 347 165 381 199
rect 623 327 657 361
rect 623 255 657 289
rect 531 165 565 199
rect 878 327 912 361
rect 878 255 912 289
rect 713 165 747 199
rect 347 49 380 73
rect 380 49 381 73
rect 347 39 381 49
rect 531 39 565 73
rect 713 49 717 73
rect 717 49 747 73
rect 713 39 747 49
<< metal1 >>
tri 435 1025 441 1031 se
rect 441 1025 487 1031
tri 487 1025 493 1031 sw
rect 0 1019 940 1025
rect 0 985 447 1019
rect 481 985 940 1019
rect 0 947 940 985
rect 0 913 447 947
rect 481 913 940 947
rect 0 901 940 913
rect 127 787 801 793
rect 127 753 139 787
rect 173 753 215 787
rect 249 753 291 787
rect 325 753 603 787
rect 637 753 679 787
rect 713 753 755 787
rect 789 753 801 787
rect 127 709 801 753
rect 127 675 139 709
rect 173 675 215 709
rect 249 675 291 709
rect 325 675 603 709
rect 637 675 679 709
rect 713 675 755 709
rect 789 675 801 709
rect 127 669 801 675
rect 0 595 940 601
rect 0 561 378 595
rect 412 561 450 595
rect 484 561 940 595
rect 0 555 940 561
rect 12 517 834 523
rect 12 483 24 517
rect 58 483 96 517
rect 130 483 404 517
rect 438 483 476 517
rect 510 483 716 517
rect 750 483 788 517
rect 822 483 834 517
rect 12 477 834 483
rect 617 361 663 373
tri 663 361 675 373 sw
tri 860 361 872 373 se
rect 872 361 918 373
rect 617 327 623 361
rect 657 331 675 361
tri 675 331 705 361 sw
tri 830 331 860 361 se
rect 860 331 878 361
rect 657 327 878 331
rect 912 327 918 361
rect 617 289 918 327
rect 617 255 623 289
rect 657 285 878 289
rect 657 255 675 285
tri 675 255 705 285 nw
tri 830 255 860 285 ne
rect 860 255 878 285
rect 912 255 918 289
rect 617 243 663 255
tri 663 243 675 255 nw
tri 860 243 872 255 ne
rect 872 243 918 255
rect 0 199 935 211
rect 0 165 347 199
rect 381 165 531 199
rect 565 165 713 199
rect 747 165 935 199
rect 0 73 935 165
rect 0 39 347 73
rect 381 39 531 73
rect 565 39 713 73
rect 747 39 935 73
rect 0 27 935 39
use nfet_CDNS_52468879185930  nfet_CDNS_52468879185930_0
timestamp 1704896540
transform -1 0 704 0 1 179
box -79 -32 115 232
use nfet_CDNS_52468879185930  nfet_CDNS_52468879185930_1
timestamp 1704896540
transform -1 0 520 0 1 179
box -79 -32 115 232
use nfet_CDNS_52468879185930  nfet_CDNS_52468879185930_2
timestamp 1704896540
transform 1 0 576 0 1 179
box -79 -32 115 232
use nfet_CDNS_52468879185930  nfet_CDNS_52468879185930_3
timestamp 1704896540
transform 1 0 392 0 1 179
box -79 -32 115 232
use pfet_CDNS_52468879185931  pfet_CDNS_52468879185931_0
timestamp 1704896540
transform -1 0 436 0 -1 1243
box -89 -36 189 636
use pfet_CDNS_52468879185931  pfet_CDNS_52468879185931_1
timestamp 1704896540
transform 1 0 492 0 -1 1243
box -89 -36 189 636
use pfet_CDNS_52468879185932  pfet_CDNS_52468879185932_0
timestamp 1704896540
transform -1 0 128 0 -1 1213
box -89 -36 125 636
use pfet_CDNS_52468879185932  pfet_CDNS_52468879185932_1
timestamp 1704896540
transform 1 0 800 0 -1 1213
box -89 -36 125 636
<< labels >>
flabel metal1 s 632 477 701 523 0 FreeSans 500 0 0 0 out_n
port 1 nsew
flabel metal1 s 741 285 795 331 0 FreeSans 500 0 0 0 out
port 2 nsew
flabel metal1 s 801 922 902 1004 0 FreeSans 500 0 0 0 vpwr
port 3 nsew
flabel metal1 s 608 69 686 173 0 FreeSans 500 0 0 0 vgnd
port 4 nsew
flabel metal1 s 825 555 934 601 0 FreeSans 500 0 0 0 in_dis
port 5 nsew
flabel locali s 85 411 129 445 0 FreeSans 500 0 0 0 in
port 6 nsew
<< properties >>
string GDS_END 80651646
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80643548
string path 7.800 1.650 19.625 1.650 
<< end >>
