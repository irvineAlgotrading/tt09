magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 37 3488 661 4329
<< pwell >>
rect -28 1922 1454 2008
rect -28 100 58 1922
rect 1368 100 1454 1922
rect -28 14 1454 100
<< mvpsubdiff >>
rect -2 1948 102 1982
rect 136 1948 170 1982
rect 204 1948 238 1982
rect 272 1948 306 1982
rect 340 1948 374 1982
rect 408 1948 442 1982
rect 476 1948 510 1982
rect 544 1948 578 1982
rect 612 1948 646 1982
rect 680 1948 714 1982
rect 748 1948 782 1982
rect 816 1948 850 1982
rect 884 1948 918 1982
rect 952 1948 986 1982
rect 1020 1948 1054 1982
rect 1088 1948 1122 1982
rect 1156 1948 1190 1982
rect 1224 1948 1258 1982
rect 1292 1948 1326 1982
rect 1360 1948 1428 1982
rect -2 1914 32 1948
rect 1394 1910 1428 1948
rect -2 1846 32 1880
rect 1394 1842 1428 1876
rect -2 1778 32 1812
rect -2 1710 32 1744
rect -2 1642 32 1676
rect -2 1574 32 1608
rect -2 1506 32 1540
rect -2 1438 32 1472
rect -2 1370 32 1404
rect -2 1302 32 1336
rect -2 1234 32 1268
rect -2 1166 32 1200
rect -2 1098 32 1132
rect -2 1030 32 1064
rect -2 962 32 996
rect -2 894 32 928
rect -2 826 32 860
rect 1394 1774 1428 1808
rect 1394 1706 1428 1740
rect 1394 1638 1428 1672
rect 1394 1570 1428 1604
rect 1394 1502 1428 1536
rect 1394 1434 1428 1468
rect 1394 1366 1428 1400
rect 1394 1298 1428 1332
rect 1394 1230 1428 1264
rect 1394 1162 1428 1196
rect 1394 1094 1428 1128
rect 1394 1026 1428 1060
rect 1394 958 1428 992
rect 1394 890 1428 924
rect -2 758 32 792
rect 1394 822 1428 856
rect -2 690 32 724
rect -2 622 32 656
rect -2 554 32 588
rect -2 486 32 520
rect 1394 754 1428 788
rect 1394 686 1428 720
rect 1394 618 1428 652
rect 1394 550 1428 584
rect 1394 482 1428 516
rect -2 418 32 452
rect 1394 414 1428 448
rect -2 350 32 384
rect -2 282 32 316
rect -2 214 32 248
rect -2 74 32 180
rect 1394 346 1428 380
rect 1394 278 1428 312
rect 1394 210 1428 244
rect 1394 142 1428 176
rect 1394 74 1428 108
rect -2 40 66 74
rect 100 40 134 74
rect 168 40 202 74
rect 236 40 270 74
rect 304 40 338 74
rect 372 40 406 74
rect 440 40 474 74
rect 508 40 542 74
rect 576 40 610 74
rect 644 40 678 74
rect 712 40 746 74
rect 780 40 814 74
rect 848 40 882 74
rect 916 40 950 74
rect 984 40 1018 74
rect 1052 40 1086 74
rect 1120 40 1154 74
rect 1188 40 1222 74
rect 1256 40 1290 74
rect 1324 40 1428 74
<< mvnsubdiff >>
rect 104 4228 138 4262
rect 172 4228 206 4262
rect 240 4228 274 4262
rect 308 4228 342 4262
rect 376 4228 410 4262
rect 444 4228 478 4262
rect 512 4228 594 4262
<< mvpsubdiffcont >>
rect 102 1948 136 1982
rect 170 1948 204 1982
rect 238 1948 272 1982
rect 306 1948 340 1982
rect 374 1948 408 1982
rect 442 1948 476 1982
rect 510 1948 544 1982
rect 578 1948 612 1982
rect 646 1948 680 1982
rect 714 1948 748 1982
rect 782 1948 816 1982
rect 850 1948 884 1982
rect 918 1948 952 1982
rect 986 1948 1020 1982
rect 1054 1948 1088 1982
rect 1122 1948 1156 1982
rect 1190 1948 1224 1982
rect 1258 1948 1292 1982
rect 1326 1948 1360 1982
rect -2 1880 32 1914
rect -2 1812 32 1846
rect 1394 1876 1428 1910
rect -2 1744 32 1778
rect -2 1676 32 1710
rect -2 1608 32 1642
rect -2 1540 32 1574
rect -2 1472 32 1506
rect -2 1404 32 1438
rect -2 1336 32 1370
rect -2 1268 32 1302
rect -2 1200 32 1234
rect -2 1132 32 1166
rect -2 1064 32 1098
rect -2 996 32 1030
rect -2 928 32 962
rect -2 860 32 894
rect 1394 1808 1428 1842
rect 1394 1740 1428 1774
rect 1394 1672 1428 1706
rect 1394 1604 1428 1638
rect 1394 1536 1428 1570
rect 1394 1468 1428 1502
rect 1394 1400 1428 1434
rect 1394 1332 1428 1366
rect 1394 1264 1428 1298
rect 1394 1196 1428 1230
rect 1394 1128 1428 1162
rect 1394 1060 1428 1094
rect 1394 992 1428 1026
rect 1394 924 1428 958
rect 1394 856 1428 890
rect -2 792 32 826
rect 1394 788 1428 822
rect -2 724 32 758
rect -2 656 32 690
rect -2 588 32 622
rect -2 520 32 554
rect -2 452 32 486
rect 1394 720 1428 754
rect 1394 652 1428 686
rect 1394 584 1428 618
rect 1394 516 1428 550
rect -2 384 32 418
rect 1394 448 1428 482
rect -2 316 32 350
rect -2 248 32 282
rect -2 180 32 214
rect 1394 380 1428 414
rect 1394 312 1428 346
rect 1394 244 1428 278
rect 1394 176 1428 210
rect 1394 108 1428 142
rect 66 40 100 74
rect 134 40 168 74
rect 202 40 236 74
rect 270 40 304 74
rect 338 40 372 74
rect 406 40 440 74
rect 474 40 508 74
rect 542 40 576 74
rect 610 40 644 74
rect 678 40 712 74
rect 746 40 780 74
rect 814 40 848 74
rect 882 40 916 74
rect 950 40 984 74
rect 1018 40 1052 74
rect 1086 40 1120 74
rect 1154 40 1188 74
rect 1222 40 1256 74
rect 1290 40 1324 74
<< mvnsubdiffcont >>
rect 138 4228 172 4262
rect 206 4228 240 4262
rect 274 4228 308 4262
rect 342 4228 376 4262
rect 410 4228 444 4262
rect 478 4228 512 4262
<< poly >>
rect 122 3956 256 3972
rect 122 3922 138 3956
rect 172 3922 206 3956
rect 240 3922 256 3956
rect 122 3906 256 3922
rect 156 3786 290 3802
rect 156 3752 172 3786
rect 206 3752 240 3786
rect 274 3752 290 3786
rect 156 3736 290 3752
rect 203 1872 609 1888
rect 203 1838 219 1872
rect 253 1838 287 1872
rect 321 1838 355 1872
rect 389 1838 423 1872
rect 457 1838 491 1872
rect 525 1838 559 1872
rect 593 1838 609 1872
rect 203 1822 609 1838
rect 651 1872 785 1888
rect 651 1838 667 1872
rect 701 1838 735 1872
rect 769 1838 785 1872
rect 651 1822 785 1838
rect 203 836 1091 852
rect 203 802 219 836
rect 253 802 287 836
rect 321 802 355 836
rect 389 802 423 836
rect 457 802 491 836
rect 525 802 559 836
rect 593 802 627 836
rect 661 802 696 836
rect 730 802 765 836
rect 799 802 834 836
rect 868 802 903 836
rect 937 802 972 836
rect 1006 802 1041 836
rect 1075 802 1091 836
rect 203 786 1091 802
rect 203 442 491 458
rect 203 408 219 442
rect 253 408 293 442
rect 327 408 367 442
rect 401 408 441 442
rect 475 408 491 442
rect 203 392 491 408
rect 547 442 835 458
rect 547 408 563 442
rect 597 408 637 442
rect 671 408 711 442
rect 745 408 785 442
rect 819 408 835 442
rect 547 392 835 408
<< polycont >>
rect 138 3922 172 3956
rect 206 3922 240 3956
rect 172 3752 206 3786
rect 240 3752 274 3786
rect 219 1838 253 1872
rect 287 1838 321 1872
rect 355 1838 389 1872
rect 423 1838 457 1872
rect 491 1838 525 1872
rect 559 1838 593 1872
rect 667 1838 701 1872
rect 735 1838 769 1872
rect 219 802 253 836
rect 287 802 321 836
rect 355 802 389 836
rect 423 802 457 836
rect 491 802 525 836
rect 559 802 593 836
rect 627 802 661 836
rect 696 802 730 836
rect 765 802 799 836
rect 834 802 868 836
rect 903 802 937 836
rect 972 802 1006 836
rect 1041 802 1075 836
rect 219 408 253 442
rect 293 408 327 442
rect 367 408 401 442
rect 441 408 475 442
rect 563 408 597 442
rect 637 408 671 442
rect 711 408 745 442
rect 785 408 819 442
<< locali >>
rect 172 4228 178 4262
rect 240 4228 252 4262
rect 308 4228 326 4262
rect 376 4228 400 4262
rect 444 4228 474 4262
rect 512 4228 548 4262
rect 582 4228 594 4262
rect 111 4050 145 4088
rect 267 4050 301 4088
rect 149 3956 187 3957
rect 172 3923 187 3956
rect 122 3922 138 3923
rect 172 3922 206 3923
rect 240 3922 256 3956
rect 156 3752 172 3786
rect 227 3752 240 3786
rect 111 3620 145 3658
rect 267 3600 301 3638
rect -8 1982 1434 1988
rect -8 1948 70 1982
rect 136 1948 143 1982
rect 204 1948 216 1982
rect 272 1948 289 1982
rect 340 1948 362 1982
rect 408 1948 442 1982
rect 505 1948 510 1982
rect 544 1948 548 1982
rect 612 1948 625 1982
rect 680 1948 702 1982
rect 748 1948 779 1982
rect 816 1948 850 1982
rect 890 1948 918 1982
rect 967 1948 986 1982
rect 1044 1948 1054 1982
rect 1156 1948 1166 1982
rect 1224 1948 1244 1982
rect 1292 1948 1322 1982
rect 1360 1948 1434 1982
rect -8 1942 1434 1948
rect -8 1914 38 1942
rect -8 1876 -2 1914
rect 32 1876 38 1914
rect -8 1846 38 1876
rect 1388 1910 1434 1942
rect 1388 1876 1394 1910
rect 1428 1876 1434 1910
rect -8 1802 -2 1846
rect 32 1802 38 1846
rect 203 1838 219 1872
rect 272 1838 287 1872
rect 351 1838 355 1872
rect 389 1838 397 1872
rect 457 1838 477 1872
rect 525 1838 557 1872
rect 593 1838 609 1872
rect 651 1838 667 1872
rect 701 1838 735 1872
rect 773 1838 785 1872
rect 1388 1842 1434 1876
rect -8 1778 38 1802
rect -8 1728 -2 1778
rect 32 1728 38 1778
rect -8 1710 38 1728
rect 1388 1804 1394 1842
rect 1428 1804 1434 1842
rect 1388 1774 1434 1804
rect 1388 1732 1394 1774
rect 1428 1732 1434 1774
rect -8 1654 -2 1710
rect 32 1654 38 1710
rect -8 1642 38 1654
rect -8 1580 -2 1642
rect 32 1580 38 1642
rect -8 1574 38 1580
rect -8 1472 -2 1574
rect 32 1472 38 1574
rect -8 1466 38 1472
rect -8 1404 -2 1466
rect 32 1404 38 1466
rect -8 1392 38 1404
rect -8 1336 -2 1392
rect 32 1336 38 1392
rect -8 1318 38 1336
rect -8 1268 -2 1318
rect 32 1268 38 1318
rect -8 1244 38 1268
rect -8 1200 -2 1244
rect 32 1200 38 1244
rect -8 1170 38 1200
rect 158 1635 192 1682
rect 158 1554 192 1601
rect 158 1473 192 1520
rect 158 1392 192 1439
rect 158 1312 192 1358
rect 158 1232 192 1278
rect 334 1635 368 1682
rect 334 1554 368 1601
rect 334 1473 368 1520
rect 334 1392 368 1439
rect 334 1312 368 1358
rect 334 1232 368 1278
rect 444 1635 478 1682
rect 444 1554 478 1601
rect 444 1473 478 1520
rect 444 1392 478 1439
rect 444 1312 478 1358
rect 444 1232 478 1278
rect 620 1635 654 1682
rect 620 1554 654 1601
rect 620 1473 654 1520
rect 620 1392 654 1439
rect 620 1312 654 1358
rect 620 1232 654 1278
rect 796 1635 830 1682
rect 796 1554 830 1601
rect 796 1473 830 1520
rect 796 1392 830 1439
rect 796 1312 830 1358
rect 796 1232 830 1278
rect 1388 1706 1434 1732
rect 1388 1660 1394 1706
rect 1428 1660 1434 1706
rect 1388 1638 1434 1660
rect 1388 1588 1394 1638
rect 1428 1588 1434 1638
rect 1388 1570 1434 1588
rect 1388 1516 1394 1570
rect 1428 1516 1434 1570
rect 1388 1502 1434 1516
rect 1388 1444 1394 1502
rect 1428 1444 1434 1502
rect 1388 1434 1434 1444
rect 1388 1372 1394 1434
rect 1428 1372 1434 1434
rect 1388 1366 1434 1372
rect 1388 1300 1394 1366
rect 1428 1300 1434 1366
rect 1388 1298 1434 1300
rect 1388 1264 1394 1298
rect 1428 1264 1434 1298
rect 1388 1262 1434 1264
rect -8 1132 -2 1170
rect 32 1132 38 1170
rect -8 1098 38 1132
rect -8 1062 -2 1098
rect 32 1062 38 1098
rect 1388 1196 1394 1262
rect 1428 1196 1434 1262
rect 1388 1190 1434 1196
rect 1388 1128 1394 1190
rect 1428 1128 1434 1190
rect 1388 1118 1434 1128
rect -8 1030 38 1062
rect -8 989 -2 1030
rect 32 989 38 1030
rect -8 962 38 989
rect 158 1010 192 1048
rect 630 1010 664 1048
rect -8 916 -2 962
rect 32 916 38 962
rect -8 894 38 916
rect 1102 1010 1136 1048
rect 394 930 428 968
rect 1388 1060 1394 1118
rect 1428 1060 1434 1118
rect 1388 1045 1434 1060
rect 1388 992 1394 1045
rect 1428 992 1434 1045
rect 866 930 900 968
rect 1388 972 1434 992
rect 1388 924 1394 972
rect 1428 924 1434 972
rect 1388 899 1434 924
rect -8 843 -2 894
rect 32 843 38 894
rect -8 826 38 843
rect 1388 856 1394 899
rect 1428 856 1434 899
rect -8 770 -2 826
rect 32 770 38 826
rect 203 802 219 836
rect 253 802 276 836
rect 321 802 355 836
rect 389 802 423 836
rect 468 802 491 836
rect 547 802 559 836
rect 626 802 627 836
rect 661 802 671 836
rect 730 802 751 836
rect 799 802 831 836
rect 868 802 903 836
rect 945 802 972 836
rect 1025 802 1041 836
rect 1075 802 1091 836
rect 1388 826 1434 856
rect -8 758 38 770
rect -8 697 -2 758
rect 32 697 38 758
rect 1388 788 1394 826
rect 1428 788 1434 826
rect 1388 754 1434 788
rect -8 690 38 697
rect -8 624 -2 690
rect 32 624 38 690
rect 394 680 428 718
rect -8 622 38 624
rect -8 588 -2 622
rect 32 588 38 622
rect -8 585 38 588
rect -8 520 -2 585
rect 32 520 38 585
rect 866 680 900 718
rect 158 600 192 638
rect 1388 719 1394 754
rect 1428 719 1434 754
rect 1388 686 1434 719
rect 630 600 664 638
rect 1102 600 1136 638
rect 1388 646 1394 686
rect 1428 646 1434 686
rect 1388 618 1434 646
rect 1388 573 1394 618
rect 1428 573 1434 618
rect -8 512 38 520
rect -8 452 -2 512
rect 32 452 38 512
rect -8 439 38 452
rect 1388 550 1434 573
rect 1388 500 1394 550
rect 1428 500 1434 550
rect 1388 482 1434 500
rect -8 384 -2 439
rect 32 384 38 439
rect 203 408 219 442
rect 286 408 293 442
rect 327 408 328 442
rect 362 408 367 442
rect 401 408 404 442
rect 438 408 441 442
rect 475 408 491 442
rect 547 408 563 442
rect 616 408 637 442
rect 692 408 711 442
rect 768 408 785 442
rect 819 408 835 442
rect 1388 427 1394 482
rect 1428 427 1434 482
rect 1388 414 1434 427
rect -8 366 38 384
rect -8 316 -2 366
rect 32 316 38 366
rect 1388 380 1394 414
rect 1428 380 1434 414
rect -8 293 38 316
rect -8 248 -2 293
rect 32 248 38 293
rect 244 282 278 320
rect -8 220 38 248
rect -8 180 -2 220
rect 32 180 38 220
rect -8 147 38 180
rect 416 282 450 320
rect 158 190 192 228
rect 588 282 622 320
rect 330 190 364 228
rect 760 282 794 320
rect 502 190 536 228
rect 1388 351 1434 380
rect 1388 312 1394 351
rect 1428 312 1434 351
rect 1388 278 1434 312
rect 674 190 708 228
rect 846 190 880 228
rect 1388 215 1394 278
rect 1428 215 1434 278
rect 1388 210 1434 215
rect 1388 176 1394 210
rect 1428 176 1434 210
rect -8 113 -2 147
rect 32 113 38 147
rect -8 80 38 113
rect 1388 146 1434 176
rect 1388 108 1394 146
rect 1428 108 1434 146
rect 1388 80 1434 108
rect -8 74 1434 80
rect -8 40 66 74
rect 104 40 134 74
rect 178 40 202 74
rect 252 40 270 74
rect 326 40 338 74
rect 400 40 406 74
rect 508 40 514 74
rect 576 40 588 74
rect 644 40 662 74
rect 712 40 736 74
rect 780 40 810 74
rect 848 40 882 74
rect 917 40 950 74
rect 990 40 1018 74
rect 1063 40 1086 74
rect 1136 40 1154 74
rect 1209 40 1222 74
rect 1282 40 1290 74
rect 1355 40 1434 74
rect -8 34 1434 40
<< viali >>
rect 104 4228 138 4262
rect 178 4228 206 4262
rect 206 4228 212 4262
rect 252 4228 274 4262
rect 274 4228 286 4262
rect 326 4228 342 4262
rect 342 4228 360 4262
rect 400 4228 410 4262
rect 410 4228 434 4262
rect 474 4228 478 4262
rect 478 4228 508 4262
rect 548 4228 582 4262
rect 111 4088 145 4122
rect 111 4016 145 4050
rect 267 4088 301 4122
rect 267 4016 301 4050
rect 115 3956 149 3957
rect 187 3956 221 3957
rect 115 3923 138 3956
rect 138 3923 149 3956
rect 187 3923 206 3956
rect 206 3923 221 3956
rect 193 3752 206 3786
rect 206 3752 227 3786
rect 265 3752 274 3786
rect 274 3752 299 3786
rect 111 3658 145 3692
rect 111 3586 145 3620
rect 267 3638 301 3672
rect 267 3566 301 3600
rect 70 1948 102 1982
rect 102 1948 104 1982
rect 143 1948 170 1982
rect 170 1948 177 1982
rect 216 1948 238 1982
rect 238 1948 250 1982
rect 289 1948 306 1982
rect 306 1948 323 1982
rect 362 1948 374 1982
rect 374 1948 396 1982
rect 471 1948 476 1982
rect 476 1948 505 1982
rect 548 1948 578 1982
rect 578 1948 582 1982
rect 625 1948 646 1982
rect 646 1948 659 1982
rect 702 1948 714 1982
rect 714 1948 736 1982
rect 779 1948 782 1982
rect 782 1948 813 1982
rect 856 1948 884 1982
rect 884 1948 890 1982
rect 933 1948 952 1982
rect 952 1948 967 1982
rect 1010 1948 1020 1982
rect 1020 1948 1044 1982
rect 1088 1948 1122 1982
rect 1166 1948 1190 1982
rect 1190 1948 1200 1982
rect 1244 1948 1258 1982
rect 1258 1948 1278 1982
rect 1322 1948 1326 1982
rect 1326 1948 1356 1982
rect -2 1880 32 1910
rect -2 1876 32 1880
rect 1394 1876 1428 1910
rect -2 1812 32 1836
rect -2 1802 32 1812
rect 238 1838 253 1872
rect 253 1838 272 1872
rect 317 1838 321 1872
rect 321 1838 351 1872
rect 397 1838 423 1872
rect 423 1838 431 1872
rect 477 1838 491 1872
rect 491 1838 511 1872
rect 557 1838 559 1872
rect 559 1838 591 1872
rect 667 1838 701 1872
rect 739 1838 769 1872
rect 769 1838 773 1872
rect -2 1744 32 1762
rect -2 1728 32 1744
rect 1394 1808 1428 1838
rect 1394 1804 1428 1808
rect 1394 1740 1428 1766
rect 1394 1732 1428 1740
rect -2 1676 32 1688
rect -2 1654 32 1676
rect -2 1608 32 1614
rect -2 1580 32 1608
rect -2 1506 32 1540
rect -2 1438 32 1466
rect -2 1432 32 1438
rect -2 1370 32 1392
rect -2 1358 32 1370
rect -2 1302 32 1318
rect -2 1284 32 1302
rect -2 1234 32 1244
rect -2 1210 32 1234
rect 158 1682 192 1716
rect 158 1601 192 1635
rect 158 1520 192 1554
rect 158 1439 192 1473
rect 158 1358 192 1392
rect 158 1278 192 1312
rect 158 1198 192 1232
rect 334 1682 368 1716
rect 334 1601 368 1635
rect 334 1520 368 1554
rect 334 1439 368 1473
rect 334 1358 368 1392
rect 334 1278 368 1312
rect 334 1198 368 1232
rect 444 1682 478 1716
rect 444 1601 478 1635
rect 444 1520 478 1554
rect 444 1439 478 1473
rect 444 1358 478 1392
rect 444 1278 478 1312
rect 444 1198 478 1232
rect 620 1682 654 1716
rect 620 1601 654 1635
rect 620 1520 654 1554
rect 620 1439 654 1473
rect 620 1358 654 1392
rect 620 1278 654 1312
rect 620 1198 654 1232
rect 796 1682 830 1716
rect 796 1601 830 1635
rect 796 1520 830 1554
rect 796 1439 830 1473
rect 796 1358 830 1392
rect 796 1278 830 1312
rect 796 1198 830 1232
rect 1394 1672 1428 1694
rect 1394 1660 1428 1672
rect 1394 1604 1428 1622
rect 1394 1588 1428 1604
rect 1394 1536 1428 1550
rect 1394 1516 1428 1536
rect 1394 1468 1428 1478
rect 1394 1444 1428 1468
rect 1394 1400 1428 1406
rect 1394 1372 1428 1400
rect 1394 1332 1428 1334
rect 1394 1300 1428 1332
rect -2 1166 32 1170
rect -2 1136 32 1166
rect -2 1064 32 1096
rect -2 1062 32 1064
rect 1394 1230 1428 1262
rect 1394 1228 1428 1230
rect 1394 1162 1428 1190
rect 1394 1156 1428 1162
rect -2 996 32 1023
rect -2 989 32 996
rect 158 1048 192 1082
rect 158 976 192 1010
rect 630 1048 664 1082
rect -2 928 32 950
rect -2 916 32 928
rect 394 968 428 1002
rect 630 976 664 1010
rect 1102 1048 1136 1082
rect 394 896 428 930
rect 866 968 900 1002
rect 1102 976 1136 1010
rect 1394 1094 1428 1118
rect 1394 1084 1428 1094
rect 1394 1026 1428 1045
rect 1394 1011 1428 1026
rect 866 896 900 930
rect 1394 958 1428 972
rect 1394 938 1428 958
rect -2 860 32 877
rect -2 843 32 860
rect 1394 890 1428 899
rect 1394 865 1428 890
rect -2 792 32 804
rect -2 770 32 792
rect 276 802 287 836
rect 287 802 310 836
rect 355 802 389 836
rect 434 802 457 836
rect 457 802 468 836
rect 513 802 525 836
rect 525 802 547 836
rect 592 802 593 836
rect 593 802 626 836
rect 671 802 696 836
rect 696 802 705 836
rect 751 802 765 836
rect 765 802 785 836
rect 831 802 834 836
rect 834 802 865 836
rect 911 802 937 836
rect 937 802 945 836
rect 991 802 1006 836
rect 1006 802 1025 836
rect -2 724 32 731
rect -2 697 32 724
rect 1394 822 1428 826
rect 1394 792 1428 822
rect -2 656 32 658
rect -2 624 32 656
rect 394 718 428 752
rect -2 554 32 585
rect -2 551 32 554
rect 158 638 192 672
rect 394 646 428 680
rect 866 718 900 752
rect 158 566 192 600
rect 630 638 664 672
rect 866 646 900 680
rect 1394 720 1428 753
rect 1394 719 1428 720
rect 630 566 664 600
rect 1102 638 1136 672
rect 1102 566 1136 600
rect 1394 652 1428 680
rect 1394 646 1428 652
rect 1394 584 1428 607
rect 1394 573 1428 584
rect -2 486 32 512
rect -2 478 32 486
rect 1394 516 1428 534
rect 1394 500 1428 516
rect -2 418 32 439
rect -2 405 32 418
rect 252 408 253 442
rect 253 408 286 442
rect 328 408 362 442
rect 404 408 438 442
rect 582 408 597 442
rect 597 408 616 442
rect 658 408 671 442
rect 671 408 692 442
rect 734 408 745 442
rect 745 408 768 442
rect 1394 448 1428 461
rect 1394 427 1428 448
rect -2 350 32 366
rect -2 332 32 350
rect -2 282 32 293
rect -2 259 32 282
rect 244 320 278 354
rect -2 214 32 220
rect -2 186 32 214
rect 158 228 192 262
rect 244 248 278 282
rect 416 320 450 354
rect 158 156 192 190
rect 330 228 364 262
rect 416 248 450 282
rect 588 320 622 354
rect 330 156 364 190
rect 502 228 536 262
rect 588 248 622 282
rect 760 320 794 354
rect 502 156 536 190
rect 674 228 708 262
rect 760 248 794 282
rect 1394 346 1428 351
rect 1394 317 1428 346
rect 674 156 708 190
rect 846 228 880 262
rect 846 156 880 190
rect 1394 244 1428 249
rect 1394 215 1428 244
rect -2 113 32 147
rect 1394 142 1428 146
rect 1394 112 1428 142
rect 70 40 100 74
rect 100 40 104 74
rect 144 40 168 74
rect 168 40 178 74
rect 218 40 236 74
rect 236 40 252 74
rect 292 40 304 74
rect 304 40 326 74
rect 366 40 372 74
rect 372 40 400 74
rect 440 40 474 74
rect 514 40 542 74
rect 542 40 548 74
rect 588 40 610 74
rect 610 40 622 74
rect 662 40 678 74
rect 678 40 696 74
rect 736 40 746 74
rect 746 40 770 74
rect 810 40 814 74
rect 814 40 844 74
rect 883 40 916 74
rect 916 40 917 74
rect 956 40 984 74
rect 984 40 990 74
rect 1029 40 1052 74
rect 1052 40 1063 74
rect 1102 40 1120 74
rect 1120 40 1136 74
rect 1175 40 1188 74
rect 1188 40 1209 74
rect 1248 40 1256 74
rect 1256 40 1282 74
rect 1321 40 1324 74
rect 1324 40 1355 74
<< metal1 >>
rect 91 4262 594 4268
rect 91 4228 104 4262
rect 138 4228 178 4262
rect 212 4228 252 4262
rect 286 4228 326 4262
rect 360 4228 400 4262
rect 434 4228 474 4262
rect 508 4228 548 4262
rect 582 4228 594 4262
rect 91 4222 594 4228
rect 91 4122 151 4222
tri 151 4188 185 4222 nw
rect 91 4088 111 4122
rect 145 4088 151 4122
rect 91 4050 151 4088
rect 91 4016 111 4050
rect 145 4016 151 4050
rect 91 4004 151 4016
rect 261 4122 313 4134
rect 261 4088 267 4122
rect 301 4088 313 4122
rect 261 4050 313 4088
rect 261 4016 267 4050
rect 301 4016 313 4050
rect 101 3957 233 3963
rect 101 3923 115 3957
rect 149 3923 187 3957
rect 221 3923 233 3957
rect 101 3917 233 3923
rect 101 3695 153 3917
tri 153 3883 187 3917 nw
rect 261 3868 313 4016
tri 227 3792 261 3826 se
rect 261 3804 313 3816
rect 181 3786 261 3792
rect 181 3752 193 3786
rect 227 3752 261 3786
rect 181 3746 313 3752
rect 101 3631 153 3643
rect 101 3573 153 3579
rect 261 3672 307 3684
rect 261 3638 267 3672
rect 301 3638 307 3672
rect 261 3600 307 3638
rect 261 3566 267 3600
rect 301 3566 307 3600
tri 227 3369 261 3403 se
rect 261 3369 307 3566
tri 307 3369 341 3403 sw
rect 137 3169 817 3369
rect 116 2938 267 2990
rect 319 2938 360 2990
rect 412 2938 1037 2990
rect 101 2858 107 2910
rect 159 2858 171 2910
rect 223 2858 1037 2910
rect 116 2772 1037 2830
rect 116 2720 824 2772
rect 876 2720 1037 2772
rect 116 2688 1037 2720
rect 116 2636 824 2688
rect 876 2636 1037 2688
rect 116 2630 1037 2636
rect 116 2538 674 2590
rect 726 2538 738 2590
rect 790 2538 1037 2590
rect 116 2458 211 2510
rect 263 2458 275 2510
rect 327 2458 1037 2510
rect -8 1982 1434 1988
rect -8 1948 70 1982
rect 104 1948 143 1982
rect 177 1948 216 1982
rect 250 1948 289 1982
rect 323 1948 362 1982
rect 396 1948 471 1982
rect 505 1948 548 1982
rect 582 1948 625 1982
rect 659 1948 702 1982
rect 736 1948 779 1982
rect 813 1948 856 1982
rect 890 1948 933 1982
rect 967 1948 1010 1982
rect 1044 1948 1088 1982
rect 1122 1948 1166 1982
rect 1200 1948 1244 1982
rect 1278 1948 1322 1982
rect 1356 1948 1434 1982
rect -8 1942 1434 1948
rect -8 1910 40 1942
tri 40 1910 72 1942 nw
tri 1354 1910 1386 1942 ne
rect 1386 1910 1434 1942
rect -8 1876 -2 1910
rect 32 1876 38 1910
tri 38 1908 40 1910 nw
tri 1386 1908 1388 1910 ne
rect -8 1836 38 1876
rect -8 1802 -2 1836
rect 32 1802 38 1836
rect 205 1829 211 1881
rect 263 1872 275 1881
rect 327 1872 603 1881
rect 272 1838 275 1872
rect 351 1838 397 1872
rect 431 1838 477 1872
rect 511 1838 557 1872
rect 591 1838 603 1872
rect 263 1829 275 1838
rect 327 1829 603 1838
rect 655 1829 663 1881
rect 715 1829 727 1881
rect 779 1829 785 1881
rect 1388 1876 1394 1910
rect 1428 1876 1434 1910
rect 1388 1838 1434 1876
rect -8 1762 38 1802
rect -8 1728 -2 1762
rect 32 1728 38 1762
rect 1388 1804 1394 1838
rect 1428 1804 1434 1838
rect 1388 1766 1434 1804
rect 1388 1732 1394 1766
rect 1428 1732 1434 1766
rect -8 1688 38 1728
rect -8 1654 -2 1688
rect 32 1654 38 1688
rect -8 1614 38 1654
rect -8 1580 -2 1614
rect 32 1580 38 1614
rect -8 1540 38 1580
rect -8 1506 -2 1540
rect 32 1506 38 1540
rect -8 1466 38 1506
rect -8 1432 -2 1466
rect 32 1432 38 1466
rect -8 1392 38 1432
rect -8 1358 -2 1392
rect 32 1358 38 1392
rect -8 1318 38 1358
rect -8 1284 -2 1318
rect 32 1284 38 1318
rect -8 1244 38 1284
rect -8 1210 -2 1244
rect 32 1210 38 1244
rect -8 1170 38 1210
rect 149 1716 201 1728
rect 149 1682 158 1716
rect 192 1682 201 1716
rect 149 1635 201 1682
rect 149 1601 158 1635
rect 192 1601 201 1635
rect 149 1554 201 1601
rect 149 1520 158 1554
rect 192 1520 201 1554
rect 149 1473 201 1520
rect 149 1439 158 1473
rect 192 1439 201 1473
rect 149 1392 201 1439
rect 149 1358 158 1392
rect 192 1358 201 1392
rect 149 1312 201 1358
rect 149 1308 158 1312
rect 192 1308 201 1312
rect 149 1244 201 1256
rect 149 1186 201 1192
rect 321 1716 374 1728
rect 321 1682 334 1716
rect 368 1682 374 1716
rect 321 1635 374 1682
rect 321 1601 334 1635
rect 368 1601 374 1635
rect 321 1557 374 1601
rect 373 1505 374 1557
rect 321 1493 374 1505
rect 373 1441 374 1493
rect 321 1439 334 1441
rect 368 1439 374 1441
rect 321 1392 374 1439
rect 321 1358 334 1392
rect 368 1358 374 1392
rect 321 1312 374 1358
rect 321 1278 334 1312
rect 368 1278 374 1312
rect 321 1232 374 1278
rect 321 1198 334 1232
rect 368 1198 374 1232
rect 321 1186 374 1198
rect 435 1716 487 1728
rect 435 1682 444 1716
rect 478 1682 487 1716
rect 435 1635 487 1682
rect 435 1601 444 1635
rect 478 1601 487 1635
rect 435 1554 487 1601
rect 435 1520 444 1554
rect 478 1520 487 1554
rect 435 1473 487 1520
rect 435 1439 444 1473
rect 478 1439 487 1473
rect 435 1392 487 1439
rect 435 1358 444 1392
rect 478 1358 487 1392
rect 435 1312 487 1358
rect 435 1308 444 1312
rect 478 1308 487 1312
rect 435 1244 487 1256
rect 435 1186 487 1192
rect 611 1716 663 1728
rect 611 1682 620 1716
rect 654 1682 663 1716
rect 611 1635 663 1682
rect 611 1601 620 1635
rect 654 1601 663 1635
rect 611 1600 663 1601
rect 611 1536 620 1548
rect 654 1536 663 1548
rect 611 1473 663 1484
rect 611 1439 620 1473
rect 654 1439 663 1473
rect 611 1392 663 1439
rect 611 1358 620 1392
rect 654 1358 663 1392
rect 611 1312 663 1358
rect 611 1278 620 1312
rect 654 1278 663 1312
rect 611 1232 663 1278
rect 611 1198 620 1232
rect 654 1198 663 1232
rect 611 1186 663 1198
rect 790 1716 836 1728
rect 790 1682 796 1716
rect 830 1682 836 1716
rect 790 1635 836 1682
rect 790 1601 796 1635
rect 830 1601 836 1635
rect 790 1554 836 1601
rect 790 1520 796 1554
rect 830 1520 836 1554
rect 790 1473 836 1520
rect 790 1439 796 1473
rect 830 1444 836 1473
rect 1388 1694 1434 1732
rect 1388 1660 1394 1694
rect 1428 1660 1434 1694
rect 1388 1622 1434 1660
rect 1388 1588 1394 1622
rect 1428 1588 1434 1622
rect 1388 1550 1434 1588
rect 1388 1516 1394 1550
rect 1428 1516 1434 1550
rect 1388 1478 1434 1516
tri 836 1444 859 1467 sw
tri 1365 1444 1388 1467 se
rect 1388 1444 1394 1478
rect 1428 1444 1434 1478
rect 830 1439 859 1444
rect 790 1433 859 1439
tri 859 1433 870 1444 sw
tri 1354 1433 1365 1444 se
rect 1365 1433 1434 1444
rect 790 1406 1434 1433
rect 790 1392 1394 1406
rect 790 1358 796 1392
rect 830 1372 1394 1392
rect 1428 1372 1434 1406
rect 830 1358 1434 1372
rect 790 1334 1434 1358
rect 790 1312 1394 1334
rect 790 1278 796 1312
rect 830 1300 1394 1312
rect 1428 1300 1434 1334
rect 830 1278 1434 1300
rect 790 1262 1434 1278
rect 790 1232 1394 1262
rect 790 1198 796 1232
rect 830 1228 1394 1232
rect 1428 1228 1434 1262
rect 830 1198 1434 1228
rect 790 1190 1434 1198
rect 790 1186 1394 1190
rect -8 1136 -2 1170
rect 32 1136 38 1170
tri 1354 1156 1384 1186 ne
rect 1384 1156 1394 1186
rect 1428 1156 1434 1190
tri 1384 1152 1388 1156 ne
rect -8 1096 38 1136
rect -8 1062 -2 1096
rect 32 1062 38 1096
rect 1388 1118 1434 1156
rect -8 1023 38 1062
rect -8 989 -2 1023
rect 32 989 38 1023
rect -8 950 38 989
rect 152 1082 441 1094
rect 152 1048 158 1082
rect 192 1048 441 1082
rect 152 1042 441 1048
rect 493 1042 505 1094
rect 557 1082 1142 1094
rect 557 1048 630 1082
rect 664 1048 1102 1082
rect 1136 1048 1142 1082
rect 557 1042 1142 1048
rect 152 1011 201 1042
tri 201 1011 232 1042 nw
tri 590 1014 618 1042 ne
rect 618 1014 673 1042
rect 152 1010 200 1011
tri 200 1010 201 1011 nw
rect 152 976 158 1010
rect 192 976 198 1010
tri 198 1008 200 1010 nw
rect 152 964 198 976
rect 388 1002 434 1014
tri 618 1011 621 1014 ne
rect 621 1011 673 1014
tri 673 1011 704 1042 nw
tri 1062 1014 1090 1042 ne
rect 1090 1014 1142 1042
tri 621 1010 622 1011 ne
rect 622 1010 672 1011
tri 672 1010 673 1011 nw
tri 622 1008 624 1010 ne
rect 388 968 394 1002
rect 428 968 434 1002
rect 624 976 630 1010
rect 664 976 670 1010
tri 670 1008 672 1010 nw
tri 434 968 436 970 sw
rect -8 916 -2 950
rect 32 916 38 950
rect -8 877 38 916
rect 388 938 436 968
tri 436 938 466 968 sw
rect 624 964 670 976
rect 860 1002 906 1014
tri 1090 1011 1093 1014 ne
rect 1093 1011 1142 1014
tri 1093 1010 1094 1011 ne
rect 1094 1010 1142 1011
tri 1094 1008 1096 1010 ne
tri 858 968 860 970 se
rect 860 968 866 1002
rect 900 968 906 1002
tri 854 964 858 968 se
rect 858 964 906 968
rect 1096 976 1102 1010
rect 1136 976 1142 1010
rect 1096 964 1142 976
rect 1388 1084 1394 1118
rect 1428 1084 1434 1118
rect 1388 1045 1434 1084
rect 1388 1011 1394 1045
rect 1428 1011 1434 1045
rect 1388 972 1434 1011
tri 828 938 854 964 se
rect 854 938 906 964
rect 388 936 466 938
tri 466 936 468 938 sw
tri 826 936 828 938 se
rect 828 936 906 938
rect 388 930 512 936
rect 388 896 394 930
rect 428 896 512 930
rect 388 884 512 896
rect 564 884 576 936
rect 628 930 906 936
rect 628 896 866 930
rect 900 896 906 930
rect 628 884 906 896
rect 1388 938 1394 972
rect 1428 938 1434 972
rect 1388 899 1434 938
rect -8 843 -2 877
rect 32 843 38 877
rect 1388 865 1394 899
rect 1428 865 1434 899
rect -8 804 38 843
rect -8 770 -2 804
rect 32 770 38 804
rect 264 836 672 847
rect 264 802 276 836
rect 310 802 355 836
rect 389 802 434 836
rect 468 802 513 836
rect 547 802 592 836
rect 626 802 671 836
rect 264 795 672 802
rect 724 795 736 847
rect 788 836 1037 847
rect 788 802 831 836
rect 865 802 911 836
rect 945 802 991 836
rect 1025 802 1037 836
rect 788 795 1037 802
rect 1388 826 1434 865
rect -8 731 38 770
rect 1388 792 1394 826
rect 1428 792 1434 826
rect -8 697 -2 731
rect 32 697 38 731
rect 314 712 320 764
rect 372 712 384 764
rect 436 752 906 764
rect 436 718 866 752
rect 900 718 906 752
rect 436 712 906 718
rect -8 658 38 697
tri 354 684 382 712 ne
rect 382 684 436 712
rect -8 624 -2 658
rect 32 624 38 658
rect -8 585 38 624
rect -8 551 -2 585
rect 32 551 38 585
rect 152 672 198 684
tri 382 680 386 684 ne
rect 386 680 436 684
tri 436 680 468 712 nw
tri 826 684 854 712 ne
rect 854 684 906 712
rect 1388 753 1434 792
rect 1388 719 1394 753
rect 1428 719 1434 753
tri 386 678 388 680 ne
rect 152 638 158 672
rect 192 638 198 672
rect 388 646 394 680
rect 428 646 434 680
tri 434 678 436 680 nw
tri 198 638 200 640 sw
rect 152 607 200 638
tri 200 607 231 638 sw
rect 388 634 434 646
rect 624 672 670 684
tri 854 680 858 684 ne
rect 858 680 906 684
tri 858 678 860 680 ne
tri 622 638 624 640 se
rect 624 638 630 672
rect 664 638 670 672
rect 860 646 866 680
rect 900 646 906 680
tri 670 638 672 640 sw
tri 618 634 622 638 se
rect 622 634 672 638
tri 591 607 618 634 se
rect 618 607 672 634
tri 672 607 703 638 sw
rect 860 634 906 646
rect 1096 672 1142 684
tri 1094 638 1096 640 se
rect 1096 638 1102 672
rect 1136 638 1142 672
tri 1090 634 1094 638 se
rect 1094 634 1142 638
tri 1063 607 1090 634 se
rect 1090 607 1142 634
rect 152 606 231 607
tri 231 606 232 607 sw
tri 590 606 591 607 se
rect 591 606 703 607
tri 703 606 704 607 sw
tri 1062 606 1063 607 se
rect 1063 606 1142 607
rect 152 554 158 606
rect 210 554 222 606
rect 274 600 1142 606
rect 274 566 630 600
rect 664 566 1102 600
rect 1136 566 1142 600
rect 274 554 1142 566
rect 1388 680 1434 719
rect 1388 646 1394 680
rect 1428 646 1434 680
rect 1388 607 1434 646
rect 1388 573 1394 607
rect 1428 573 1434 607
rect -8 512 38 551
rect 1388 534 1434 573
rect -8 478 -2 512
rect 32 478 38 512
tri 504 500 520 516 se
rect 520 500 906 516
rect -8 439 38 478
tri 465 461 504 500 se
rect 504 484 906 500
rect 1388 500 1394 534
rect 1428 500 1434 534
rect 504 461 523 484
tri 523 461 546 484 nw
rect 1388 461 1434 500
tri 462 458 465 461 se
rect 465 458 520 461
tri 520 458 523 461 nw
tri 452 448 462 458 se
rect 462 448 504 458
rect -8 405 -2 439
rect 32 405 38 439
rect -8 366 38 405
rect 240 442 504 448
tri 504 442 520 458 nw
rect 570 442 780 448
rect 240 408 252 442
rect 286 408 328 442
rect 362 408 404 442
rect 438 408 470 442
tri 470 408 504 442 nw
rect 570 408 582 442
rect 616 408 658 442
rect 692 408 734 442
rect 768 408 780 442
rect 240 402 464 408
tri 464 402 470 408 nw
rect 570 402 780 408
rect 1388 427 1394 461
rect 1428 427 1434 461
rect -8 332 -2 366
rect 32 332 38 366
rect -8 293 38 332
rect -8 259 -2 293
rect 32 259 38 293
rect 238 314 244 366
rect 296 314 308 366
rect 360 354 456 366
rect 360 320 416 354
rect 450 320 456 354
rect 360 314 456 320
rect 238 282 286 314
tri 286 282 318 314 nw
tri 376 282 408 314 ne
rect 408 282 456 314
rect -8 228 38 259
rect 152 262 198 274
tri 38 228 46 236 sw
tri 144 228 152 236 se
rect 152 228 158 262
rect 192 228 198 262
rect 238 248 244 282
rect 278 248 284 282
tri 284 280 286 282 nw
tri 408 280 410 282 ne
rect 238 236 284 248
rect 324 262 370 274
tri 198 228 206 236 sw
tri 316 228 324 236 se
rect 324 228 330 262
rect 364 228 370 262
rect 410 248 416 282
rect 450 248 456 282
rect 582 314 588 366
rect 640 314 652 366
rect 704 354 800 366
rect 704 320 760 354
rect 794 320 800 354
rect 704 314 800 320
rect 582 282 630 314
tri 630 282 662 314 nw
tri 720 282 752 314 ne
rect 752 282 800 314
rect 410 236 456 248
rect 496 262 542 274
tri 370 228 378 236 sw
tri 488 228 496 236 se
rect 496 228 502 262
rect 536 228 542 262
rect 582 248 588 282
rect 622 248 628 282
tri 628 280 630 282 nw
tri 752 280 754 282 ne
rect 582 236 628 248
rect 668 262 714 274
tri 542 228 550 236 sw
tri 660 228 668 236 se
rect 668 228 674 262
rect 708 228 714 262
rect 754 248 760 282
rect 794 248 800 282
rect 1388 351 1434 427
rect 1388 317 1394 351
rect 1428 317 1434 351
rect 754 236 800 248
rect 840 262 886 274
tri 714 228 722 236 sw
tri 832 228 840 236 se
rect 840 228 846 262
rect 880 228 886 262
rect 1388 249 1434 317
rect -8 220 46 228
rect -8 186 -2 220
rect 32 215 46 220
tri 46 215 59 228 sw
tri 131 215 144 228 se
rect 144 215 206 228
tri 206 215 219 228 sw
tri 303 215 316 228 se
rect 316 215 378 228
tri 378 215 391 228 sw
tri 475 215 488 228 se
rect 488 215 550 228
tri 550 215 563 228 sw
tri 647 215 660 228 se
rect 660 215 722 228
tri 722 215 735 228 sw
tri 819 215 832 228 se
rect 832 215 886 228
tri 886 215 907 236 sw
tri 1367 215 1388 236 se
rect 1388 215 1394 249
rect 1428 215 1434 249
rect 32 202 59 215
tri 59 202 72 215 sw
tri 118 202 131 215 se
rect 131 202 219 215
tri 219 202 232 215 sw
tri 290 202 303 215 se
rect 303 202 391 215
tri 391 202 404 215 sw
tri 462 202 475 215 se
rect 475 202 563 215
tri 563 202 576 215 sw
tri 634 202 647 215 se
rect 647 202 735 215
tri 735 202 748 215 sw
tri 806 202 819 215 se
rect 819 202 907 215
tri 907 202 920 215 sw
tri 1354 202 1367 215 se
rect 1367 202 1434 215
rect 32 190 1434 202
rect 32 186 158 190
rect -8 156 158 186
rect 192 156 330 190
rect 364 156 502 190
rect 536 156 674 190
rect 708 156 846 190
rect 880 156 1434 190
rect -8 147 1434 156
rect -8 113 -2 147
rect 32 146 1434 147
rect 32 113 1394 146
rect -8 112 1394 113
rect 1428 112 1434 146
rect -8 74 1434 112
rect -8 40 70 74
rect 104 40 144 74
rect 178 40 218 74
rect 252 40 292 74
rect 326 40 366 74
rect 400 40 440 74
rect 474 40 514 74
rect 548 40 588 74
rect 622 40 662 74
rect 696 40 736 74
rect 770 40 810 74
rect 844 40 883 74
rect 917 40 956 74
rect 990 40 1029 74
rect 1063 40 1102 74
rect 1136 40 1175 74
rect 1209 40 1248 74
rect 1282 40 1321 74
rect 1355 40 1434 74
rect -8 34 1434 40
<< via1 >>
rect 261 3816 313 3868
rect 261 3786 313 3804
rect 261 3752 265 3786
rect 265 3752 299 3786
rect 299 3752 313 3786
rect 101 3692 153 3695
rect 101 3658 111 3692
rect 111 3658 145 3692
rect 145 3658 153 3692
rect 101 3643 153 3658
rect 101 3620 153 3631
rect 101 3586 111 3620
rect 111 3586 145 3620
rect 145 3586 153 3620
rect 101 3579 153 3586
rect 267 2938 319 2990
rect 360 2938 412 2990
rect 107 2858 159 2910
rect 171 2858 223 2910
rect 824 2720 876 2772
rect 824 2636 876 2688
rect 674 2538 726 2590
rect 738 2538 790 2590
rect 211 2458 263 2510
rect 275 2458 327 2510
rect 211 1872 263 1881
rect 275 1872 327 1881
rect 211 1838 238 1872
rect 238 1838 263 1872
rect 275 1838 317 1872
rect 317 1838 327 1872
rect 211 1829 263 1838
rect 275 1829 327 1838
rect 663 1872 715 1881
rect 663 1838 667 1872
rect 667 1838 701 1872
rect 701 1838 715 1872
rect 663 1829 715 1838
rect 727 1872 779 1881
rect 727 1838 739 1872
rect 739 1838 773 1872
rect 773 1838 779 1872
rect 727 1829 779 1838
rect 149 1278 158 1308
rect 158 1278 192 1308
rect 192 1278 201 1308
rect 149 1256 201 1278
rect 149 1232 201 1244
rect 149 1198 158 1232
rect 158 1198 192 1232
rect 192 1198 201 1232
rect 149 1192 201 1198
rect 321 1554 373 1557
rect 321 1520 334 1554
rect 334 1520 368 1554
rect 368 1520 373 1554
rect 321 1505 373 1520
rect 321 1473 373 1493
rect 321 1441 334 1473
rect 334 1441 368 1473
rect 368 1441 373 1473
rect 435 1278 444 1308
rect 444 1278 478 1308
rect 478 1278 487 1308
rect 435 1256 487 1278
rect 435 1232 487 1244
rect 435 1198 444 1232
rect 444 1198 478 1232
rect 478 1198 487 1232
rect 435 1192 487 1198
rect 611 1554 663 1600
rect 611 1548 620 1554
rect 620 1548 654 1554
rect 654 1548 663 1554
rect 611 1520 620 1536
rect 620 1520 654 1536
rect 654 1520 663 1536
rect 611 1484 663 1520
rect 441 1042 493 1094
rect 505 1042 557 1094
rect 512 884 564 936
rect 576 884 628 936
rect 672 836 724 847
rect 672 802 705 836
rect 705 802 724 836
rect 672 795 724 802
rect 736 836 788 847
rect 736 802 751 836
rect 751 802 785 836
rect 785 802 788 836
rect 736 795 788 802
rect 320 712 372 764
rect 384 752 436 764
rect 384 718 394 752
rect 394 718 428 752
rect 428 718 436 752
rect 384 712 436 718
rect 158 600 210 606
rect 158 566 192 600
rect 192 566 210 600
rect 158 554 210 566
rect 222 554 274 606
rect 244 354 296 366
rect 244 320 278 354
rect 278 320 296 354
rect 244 314 296 320
rect 308 314 360 366
rect 588 354 640 366
rect 588 320 622 354
rect 622 320 640 354
rect 588 314 640 320
rect 652 314 704 366
<< metal2 >>
rect 261 3868 313 3874
rect 261 3804 313 3816
rect 101 3695 153 3701
rect 101 3631 153 3643
rect 101 2938 153 3579
rect 261 2990 313 3752
tri 313 2990 347 3024 sw
tri 153 2938 159 2944 sw
rect 261 2938 267 2990
rect 319 2938 360 2990
rect 412 2938 418 2990
rect 101 2910 159 2938
tri 159 2910 187 2938 sw
tri 332 2910 360 2938 ne
rect 360 2910 418 2938
rect 101 2858 107 2910
rect 159 2858 171 2910
rect 223 2858 229 2910
tri 360 2904 366 2910 ne
rect 101 1769 153 2858
tri 153 2824 187 2858 nw
rect 205 2458 211 2510
rect 263 2458 275 2510
rect 327 2458 333 2510
rect 205 1881 257 2458
tri 257 2424 291 2458 nw
rect 366 1929 418 2910
rect 824 2772 876 2778
rect 824 2688 876 2720
rect 668 2538 674 2590
rect 726 2538 738 2590
rect 790 2538 796 2590
tri 418 1929 420 1931 sw
tri 257 1881 291 1915 sw
rect 366 1902 420 1929
tri 366 1881 387 1902 ne
rect 387 1881 420 1902
tri 420 1881 468 1929 sw
tri 657 1881 668 1892 se
rect 668 1881 720 2538
tri 720 2504 754 2538 nw
tri 720 1881 754 1915 sw
rect 205 1829 211 1881
rect 263 1829 275 1881
rect 327 1829 333 1881
tri 387 1848 420 1881 ne
rect 420 1848 468 1881
tri 468 1848 501 1881 sw
tri 420 1829 439 1848 ne
rect 439 1829 501 1848
tri 501 1829 520 1848 sw
rect 657 1829 663 1881
rect 715 1829 727 1881
rect 779 1829 785 1881
tri 439 1791 477 1829 ne
rect 477 1791 520 1829
tri 101 1717 153 1769 ne
tri 153 1719 225 1791 sw
tri 477 1767 501 1791 ne
rect 501 1767 520 1791
tri 520 1767 582 1829 sw
tri 794 1773 824 1803 se
rect 824 1781 876 2636
rect 824 1773 868 1781
tri 868 1773 876 1781 nw
tri 788 1767 794 1773 se
tri 501 1719 549 1767 ne
rect 549 1719 582 1767
rect 153 1717 225 1719
tri 153 1645 225 1717 ne
tri 225 1645 299 1719 sw
tri 549 1686 582 1719 ne
tri 582 1686 663 1767 sw
tri 582 1657 611 1686 ne
tri 225 1600 270 1645 ne
rect 270 1600 299 1645
tri 299 1600 344 1645 sw
rect 611 1600 663 1686
tri 270 1571 299 1600 ne
rect 299 1571 344 1600
tri 344 1571 373 1600 sw
tri 299 1557 313 1571 ne
rect 313 1557 373 1571
tri 313 1549 321 1557 ne
rect 321 1493 373 1505
rect 611 1536 663 1548
rect 611 1478 663 1484
tri 742 1721 788 1767 se
rect 788 1721 794 1767
rect 321 1435 373 1441
rect 149 1308 201 1314
rect 149 1244 201 1256
rect 149 606 201 1192
rect 435 1308 487 1314
rect 435 1244 487 1256
rect 435 1094 487 1192
tri 487 1094 521 1128 sw
rect 435 1042 441 1094
rect 493 1042 505 1094
rect 557 1042 563 1094
rect 506 884 512 936
rect 564 884 576 936
rect 628 884 634 936
tri 548 850 582 884 ne
rect 314 712 320 764
rect 372 712 384 764
rect 436 712 442 764
tri 201 606 235 640 sw
rect 149 554 158 606
rect 210 554 222 606
rect 274 554 280 606
tri 286 366 314 394 se
rect 314 366 366 712
tri 366 678 400 712 nw
rect 238 314 244 366
rect 296 314 308 366
rect 360 314 366 366
rect 582 366 634 884
tri 708 847 742 881 se
rect 742 847 794 1721
tri 794 1699 868 1773 nw
rect 666 795 672 847
rect 724 795 736 847
rect 788 795 794 847
tri 634 366 662 394 sw
rect 582 314 588 366
rect 640 314 652 366
rect 704 314 710 366
use nfet_CDNS_5595914180818  nfet_CDNS_5595914180818_0
timestamp 1704896540
transform 1 0 665 0 1 1190
box -79 -32 199 632
use nfet_CDNS_5595914180818  nfet_CDNS_5595914180818_1
timestamp 1704896540
transform 1 0 489 0 1 1190
box -79 -32 199 632
use nfet_CDNS_5595914180818  nfet_CDNS_5595914180818_2
timestamp 1704896540
transform 1 0 203 0 1 1190
box -79 -32 199 632
use nfet_CDNS_5595914180820  nfet_CDNS_5595914180820_0
timestamp 1704896540
transform -1 0 1091 0 1 884
box -79 -32 967 232
use nfet_CDNS_5595914180820  nfet_CDNS_5595914180820_1
timestamp 1704896540
transform -1 0 1091 0 1 554
box -79 -32 967 232
use nfet_CDNS_5595914180821  nfet_CDNS_5595914180821_0
timestamp 1704896540
transform -1 0 491 0 1 160
box -79 -32 367 232
use nfet_CDNS_5595914180821  nfet_CDNS_5595914180821_1
timestamp 1704896540
transform -1 0 835 0 1 160
box -79 -32 367 232
use pfet_CDNS_5595914180822  pfet_CDNS_5595914180822_0
timestamp 1704896540
transform 1 0 156 0 1 4004
box -119 -66 219 216
use pfet_CDNS_5595914180822  pfet_CDNS_5595914180822_1
timestamp 1704896540
transform 1 0 156 0 1 3554
box -119 -66 219 216
<< labels >>
flabel metal1 s 146 2644 301 2738 3 FreeSans 200 0 0 0 vpwr_lv
port 2 nsew
flabel metal1 s 135 4234 228 4259 3 FreeSans 200 0 0 0 vpwr_hv
port 3 nsew
flabel metal1 s 144 2870 225 2900 3 FreeSans 200 0 0 0 fbk_n
port 4 nsew
flabel metal1 s 144 2947 244 2980 3 FreeSans 200 0 0 0 fbk
port 5 nsew
flabel metal1 s 146 2547 237 2581 3 FreeSans 200 0 0 0 reset
port 6 nsew
flabel metal1 s 143 2464 207 2501 3 FreeSans 200 0 0 0 hold
port 7 nsew
flabel metal1 s 637 412 732 437 3 FreeSans 200 0 0 0 switch_lv_n
port 8 nsew
flabel metal1 s 278 413 393 440 3 FreeSans 200 0 0 0 switch_lv
port 9 nsew
flabel metal1 s 133 67 301 127 3 FreeSans 200 0 0 0 vgnd
port 1 nsew
<< properties >>
string GDS_END 770478
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 729424
<< end >>
