magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< obsm2 >>
rect -6231 21500 -1085 23500
tri -1915 21330 -1745 21500 ne
rect -1745 21330 -1085 21500
tri -1085 21330 1085 23500 sw
tri -1745 18500 1085 21330 ne
tri 1085 20500 1915 21330 sw
rect 1085 18500 6008 20500
rect -6231 15500 -1085 17500
tri -1915 15330 -1745 15500 ne
rect -1745 15330 -1085 15500
tri -1085 15330 1085 17500 sw
tri -1745 12500 1085 15330 ne
tri 1085 14500 1915 15330 sw
rect 1085 12500 6008 14500
rect 9908 -1000 27500 1000
tri -1745 -18330 1085 -15500 se
rect 1085 -17500 6008 -15500
tri 1085 -18330 1915 -17500 nw
tri -1915 -18500 -1745 -18330 se
rect -1745 -18500 -1085 -18330
rect -6231 -20500 -1085 -18500
tri -1085 -20500 1085 -18330 nw
tri -1745 -24330 1085 -21500 se
rect 1085 -23500 6008 -21500
tri 1085 -24330 1915 -23500 nw
tri -1915 -24500 -1745 -24330 se
rect -1745 -24500 -1085 -24330
rect -6231 -26500 -1085 -24500
tri -1085 -26500 1085 -24330 nw
<< obsm3 >>
tri -13806 23672 -10978 26500 se
rect -10978 24500 10978 26500
tri 10978 24500 12978 26500 sw
tri -10978 23672 -10150 24500 nw
tri -15374 22104 -13806 23672 se
rect -13806 22290 -12360 23672
tri -12360 22290 -10978 23672 nw
tri 10150 23500 11150 24500 ne
rect 11150 23500 12978 24500
tri -10946 22290 -9736 23500 se
rect -9736 23253 -2202 23500
tri -2202 23253 -1955 23500 sw
rect -9736 22290 -1955 23253
rect -13806 22104 -13602 22290
tri -16634 20844 -15374 22104 se
rect -15374 21048 -13602 22104
tri -13602 21048 -12360 22290 nw
tri -12188 21048 -10946 22290 se
rect -10946 21747 -1955 22290
rect -10946 21500 -2202 21747
tri -2202 21500 -1955 21747 nw
rect -10946 21048 -10257 21500
rect -15374 20844 -14755 21048
tri -18107 19371 -16634 20844 se
rect -16634 19895 -14755 20844
tri -14755 19895 -13602 21048 nw
tri -13341 19895 -12188 21048 se
rect -12188 20151 -10257 21048
tri -10257 20151 -8908 21500 nw
tri -1745 20670 1085 23500 se
rect 1085 22290 9736 23500
tri 9736 22290 10946 23500 sw
tri 11150 22290 12360 23500 ne
rect 12360 22290 12978 23500
tri 12978 22290 15188 24500 sw
rect 1085 21500 10946 22290
tri 1085 20670 1915 21500 nw
tri -1915 20500 -1745 20670 se
rect -1745 20500 -1085 20670
tri -8842 20151 -8493 20500 se
rect -8493 20151 -1085 20500
rect -12188 19895 -11561 20151
rect -16634 19371 -15803 19895
tri -19462 18016 -18107 19371 se
rect -18107 18847 -15803 19371
tri -15803 18847 -14755 19895 nw
tri -14389 18847 -13341 19895 se
rect -13341 18847 -11561 19895
tri -11561 18847 -10257 20151 nw
tri -10146 18847 -8842 20151 se
rect -8842 18847 -1085 20151
rect -18107 18016 -16806 18847
tri -20849 16629 -19462 18016 se
rect -19462 17844 -16806 18016
tri -16806 17844 -15803 18847 nw
tri -15392 17844 -14389 18847 se
rect -14389 17844 -12736 18847
rect -19462 16629 -18220 17844
tri -22290 15188 -20849 16629 se
rect -20849 16430 -18220 16629
tri -18220 16430 -16806 17844 nw
tri -16806 16430 -15392 17844 se
rect -15392 17672 -12736 17844
tri -12736 17672 -11561 18847 nw
tri -11321 17672 -10146 18847 se
rect -10146 18500 -1085 18847
tri -1085 18500 1085 20670 nw
tri 8908 20500 9908 21500 ne
rect 9908 21048 10946 21500
tri 10946 21048 12188 22290 sw
tri 12360 21048 13602 22290 ne
rect 13602 21048 15188 22290
rect 9908 20500 12188 21048
tri 1732 20253 1979 20500 se
rect 1979 20253 8493 20500
rect 1732 19462 8493 20253
tri 8493 19462 9531 20500 sw
tri 9908 19462 10946 20500 ne
rect 10946 19634 12188 20500
tri 12188 19634 13602 21048 sw
tri 13602 19634 15016 21048 ne
rect 15016 19634 15188 21048
rect 10946 19462 13602 19634
rect 1732 18747 9531 19462
tri 1732 18500 1979 18747 ne
rect 1979 18500 9531 18747
rect -10146 17672 -9012 18500
rect -15392 16430 -14149 17672
rect -20849 15188 -19634 16430
tri -23849 13629 -22290 15188 se
rect -22290 15016 -19634 15188
tri -19634 15016 -18220 16430 nw
tri -18220 15016 -16806 16430 se
rect -16806 16259 -14149 16430
tri -14149 16259 -12736 17672 nw
tri -12734 16259 -11321 17672 se
rect -11321 17153 -9012 17672
tri -9012 17153 -7665 18500 nw
tri -7598 17153 -7251 17500 se
rect -7251 17253 -2202 17500
tri -2202 17253 -1955 17500 sw
rect -7251 17153 -1955 17253
rect -11321 16259 -10316 17153
rect -16806 15016 -15564 16259
rect -22290 13629 -21048 15016
tri -26500 10978 -23849 13629 se
rect -23849 13602 -21048 13629
tri -21048 13602 -19634 15016 nw
tri -19634 13602 -18220 15016 se
rect -18220 14844 -15564 15016
tri -15564 14844 -14149 16259 nw
tri -14149 14844 -12734 16259 se
rect -12734 15849 -10316 16259
tri -10316 15849 -9012 17153 nw
tri -8902 15849 -7598 17153 se
rect -7598 15849 -1955 17153
rect -12734 14844 -11493 15849
rect -18220 13602 -16977 14844
rect -23849 12188 -22462 13602
tri -22462 12188 -21048 13602 nw
tri -21048 12188 -19634 13602 se
rect -19634 13431 -16977 13602
tri -16977 13431 -15564 14844 nw
tri -15562 13431 -14149 14844 se
rect -14149 14672 -11493 14844
tri -11493 14672 -10316 15849 nw
tri -10079 14672 -8902 15849 se
rect -8902 15747 -1955 15849
rect -8902 15500 -2202 15747
tri -2202 15500 -1955 15747 nw
rect -8902 14672 -7774 15500
rect -14149 13431 -12907 14672
rect -19634 12188 -18392 13431
rect -23849 10978 -23672 12188
tri -23672 10978 -22462 12188 nw
tri -22258 10978 -21048 12188 se
rect -21048 12016 -18392 12188
tri -18392 12016 -16977 13431 nw
tri -16977 12016 -15562 13431 se
rect -15562 13258 -12907 13431
tri -12907 13258 -11493 14672 nw
tri -11493 13258 -10079 14672 se
rect -10079 14149 -7774 14672
tri -7774 14149 -6423 15500 nw
tri -1745 14670 1085 17500 se
rect 1085 17149 7251 17500
tri 7251 17149 7602 17500 sw
tri 7665 17149 9016 18500 ne
rect 9016 18220 9531 18500
tri 9531 18220 10773 19462 sw
tri 10946 18220 12188 19462 ne
rect 12188 18220 13602 19462
tri 13602 18220 15016 19634 sw
tri 15016 19462 15188 19634 ne
tri 15188 19462 18016 22290 sw
tri 15188 18220 16430 19462 ne
rect 16430 18220 18016 19462
rect 9016 17149 10773 18220
rect 1085 15735 7602 17149
tri 7602 15735 9016 17149 sw
tri 9016 15735 10430 17149 ne
rect 10430 16977 10773 17149
tri 10773 16977 12016 18220 sw
tri 12188 16977 13431 18220 ne
rect 13431 16977 15016 18220
rect 10430 15735 12016 16977
rect 1085 15500 9016 15735
tri 1085 14670 1915 15500 nw
tri -1915 14500 -1745 14670 se
rect -1745 14500 -1085 14670
tri -6359 14149 -6008 14500 se
rect -6008 14149 -1085 14500
rect -10079 13258 -9074 14149
rect -15562 12016 -14321 13258
rect -21048 10978 -19805 12016
rect -26500 -10978 -24500 10978
tri -24500 10150 -23672 10978 nw
tri -23500 9736 -22258 10978 se
rect -22258 10603 -19805 10978
tri -19805 10603 -18392 12016 nw
tri -18390 10603 -16977 12016 se
rect -16977 11844 -14321 12016
tri -14321 11844 -12907 13258 nw
tri -12907 11844 -11493 13258 se
rect -11493 12849 -9074 13258
tri -9074 12849 -7774 14149 nw
tri -7659 12849 -6359 14149 se
rect -6359 12849 -1085 14149
rect -11493 11844 -10259 12849
rect -16977 10603 -15735 11844
rect -22258 9736 -21220 10603
rect -23500 9188 -21220 9736
tri -21220 9188 -19805 10603 nw
tri -19805 9188 -18390 10603 se
rect -18390 10430 -15735 10603
tri -15735 10430 -14321 11844 nw
tri -14321 10430 -12907 11844 se
rect -12907 11664 -10259 11844
tri -10259 11664 -9074 12849 nw
tri -8844 11664 -7659 12849 se
rect -7659 12500 -1085 12849
tri -1085 12500 1085 14670 nw
tri 1732 14253 1979 14500 se
rect 1979 14253 6008 14500
rect 1732 14149 6008 14253
tri 6008 14149 6359 14500 sw
tri 6423 14149 7774 15500 ne
rect 7774 14321 9016 15500
tri 9016 14321 10430 15735 sw
tri 10430 14321 11844 15735 ne
rect 11844 15564 12016 15735
tri 12016 15564 13429 16977 sw
tri 13431 15564 14844 16977 ne
rect 14844 16806 15016 16977
tri 15016 16806 16430 18220 sw
tri 16430 16806 17844 18220 ne
rect 17844 16806 18016 18220
rect 14844 15564 16430 16806
rect 11844 14321 13429 15564
rect 7774 14149 10430 14321
rect 1732 12907 6359 14149
tri 6359 12907 7601 14149 sw
tri 7774 12907 9016 14149 ne
rect 9016 12907 10430 14149
tri 10430 12907 11844 14321 sw
tri 11844 12907 13258 14321 ne
rect 13258 14149 13429 14321
tri 13429 14149 14844 15564 sw
tri 14844 14149 16259 15564 ne
rect 16259 15392 16430 15564
tri 16430 15392 17844 16806 sw
tri 17844 16634 18016 16806 ne
tri 18016 16634 20844 19462 sw
tri 18016 15392 19258 16634 ne
rect 19258 15392 20844 16634
rect 16259 14149 17844 15392
rect 13258 12907 14844 14149
rect 1732 12747 7601 12907
tri 1732 12500 1979 12747 ne
rect 1979 12500 7601 12747
rect -7659 11664 -7601 12500
rect -12907 10430 -11664 11664
rect -18390 9188 -17149 10430
rect -23500 -9736 -21500 9188
tri -21500 8908 -21220 9188 nw
tri -20500 8493 -19805 9188 se
rect -19805 9016 -17149 9188
tri -17149 9016 -15735 10430 nw
tri -15735 9016 -14321 10430 se
rect -14321 10259 -11664 10430
tri -11664 10259 -10259 11664 nw
tri -10249 10259 -8844 11664 se
rect -8844 10259 -7601 11664
rect -14321 9016 -13079 10259
rect -19805 8493 -18500 9016
rect -20500 -8493 -18500 8493
tri -18500 7665 -17149 9016 nw
tri -17086 7665 -15735 9016 se
rect -15735 8844 -13079 9016
tri -13079 8844 -11664 10259 nw
tri -11664 8844 -10249 10259 se
rect -10249 10079 -7601 10259
tri -7601 10079 -5180 12500 nw
tri 5180 10079 7601 12500 ne
tri 7601 11664 8844 12907 sw
tri 9016 11664 10259 12907 ne
rect 10259 11664 11844 12907
rect 7601 10251 8844 11664
tri 8844 10251 10257 11664 sw
tri 10259 10251 11672 11664 ne
rect 11672 11493 11844 11664
tri 11844 11493 13258 12907 sw
tri 13258 11493 14672 12907 ne
rect 14672 12736 14844 12907
tri 14844 12736 16257 14149 sw
tri 16259 12736 17672 14149 ne
rect 17672 13978 17844 14149
tri 17844 13978 19258 15392 sw
tri 19258 13978 20672 15392 ne
rect 20672 13978 20844 15392
rect 17672 12736 19258 13978
rect 14672 11493 16257 12736
rect 11672 10251 13258 11493
rect 7601 10079 10257 10251
rect -10249 8844 -10015 10079
rect -15735 7665 -14492 8844
tri -17500 7251 -17086 7665 se
rect -17086 7431 -14492 7665
tri -14492 7431 -13079 8844 nw
tri -13077 7431 -11664 8844 se
rect -11664 7665 -10015 8844
tri -10015 7665 -7601 10079 nw
tri 7601 7665 10015 10079 ne
rect 10015 8836 10257 10079
tri 10257 8836 11672 10251 sw
tri 11672 8836 13087 10251 ne
rect 13087 10079 13258 10251
tri 13258 10079 14672 11493 sw
tri 14672 10079 16086 11493 ne
rect 16086 11321 16257 11493
tri 16257 11321 17672 12736 sw
tri 17672 11321 19087 12736 ne
rect 19087 12564 19258 12736
tri 19258 12564 20672 13978 sw
tri 20672 13806 20844 13978 ne
tri 20844 13806 23672 16634 sw
tri 20844 12564 22086 13806 ne
rect 22086 12564 23672 13806
rect 19087 11321 20672 12564
rect 16086 10079 17672 11321
rect 13087 8836 14672 10079
rect 10015 7665 11672 8836
rect -17086 7251 -15500 7431
rect -17500 -7251 -15500 7251
tri -15500 6423 -14492 7431 nw
tri -14085 6423 -13077 7431 se
rect -13077 6423 -11664 7431
tri -14500 6008 -14085 6423 se
rect -14085 6016 -11664 6423
tri -11664 6016 -10015 7665 nw
rect -14085 6008 -12500 6016
rect -14500 1000 -12500 6008
tri -12500 5180 -11664 6016 nw
tri 10015 6008 11672 7665 ne
tri 11672 7423 13085 8836 sw
tri 13087 7423 14500 8836 ne
rect 14500 8665 14672 8836
tri 14672 8665 16086 10079 sw
tri 16086 8665 17500 10079 ne
rect 17500 9908 17672 10079
tri 17672 9908 19085 11321 sw
tri 19087 9908 20500 11321 ne
rect 20500 11150 20672 11321
tri 20672 11150 22086 12564 sw
tri 22086 11150 23500 12564 ne
rect 23500 11150 23672 12564
rect 20500 9908 22086 11150
rect 17500 8665 19085 9908
rect 14500 7423 16086 8665
rect 11672 6008 13085 7423
tri 13085 6008 14500 7423 sw
tri 14500 6423 15500 7423 ne
rect 15500 7251 16086 7423
tri 16086 7251 17500 8665 sw
tri 17500 7665 18500 8665 ne
rect 18500 8493 19085 8665
tri 19085 8493 20500 9908 sw
tri 20500 8908 21500 9908 ne
rect 21500 9736 22086 9908
tri 22086 9736 23500 11150 sw
tri 23500 10978 23672 11150 ne
tri 23672 10978 26500 13806 sw
tri 23672 10150 24500 10978 ne
tri 11672 5180 12500 6008 ne
rect -14500 -1000 11500 1000
rect -14500 -6008 -12500 -1000
tri -26500 -12360 -25118 -10978 ne
rect -25118 -11150 -24500 -10978
tri -24500 -11150 -23500 -10150 sw
tri -23500 -11150 -22086 -9736 ne
rect -22086 -9908 -21500 -9736
tri -21500 -9908 -20500 -8908 sw
tri -20500 -9908 -19085 -8493 ne
rect -19085 -8665 -18500 -8493
tri -18500 -8665 -17500 -7665 sw
tri -17500 -8665 -16086 -7251 ne
rect -16086 -7423 -15500 -7251
tri -15500 -7423 -14500 -6423 sw
tri -14500 -7423 -13085 -6008 ne
rect -13085 -7423 -12500 -6008
rect -16086 -8665 -14500 -7423
rect -19085 -9908 -17500 -8665
rect -22086 -11150 -20500 -9908
rect -25118 -12360 -23500 -11150
tri -25118 -13806 -23672 -12360 ne
rect -23672 -12564 -23500 -12360
tri -23500 -12564 -22086 -11150 sw
tri -22086 -12564 -20672 -11150 ne
rect -20672 -11321 -20500 -11150
tri -20500 -11321 -19087 -9908 sw
tri -19085 -11321 -17672 -9908 ne
rect -17672 -10079 -17500 -9908
tri -17500 -10079 -16086 -8665 sw
tri -16086 -10079 -14672 -8665 ne
rect -14672 -8836 -14500 -8665
tri -14500 -8836 -13087 -7423 sw
tri -13085 -7665 -12843 -7423 ne
rect -12843 -7665 -12500 -7423
tri -12500 -7665 -10015 -5180 sw
tri 10429 -7251 12500 -5180 se
rect 12500 -6008 14500 6008
rect 12500 -7251 13257 -6008
tri 13257 -7251 14500 -6008 nw
tri 14672 -7251 15500 -6423 se
rect 15500 -7251 17500 7251
rect -14672 -9016 -13087 -8836
tri -13087 -9016 -12907 -8836 sw
tri -12843 -9016 -11492 -7665 ne
rect -11492 -9016 -10015 -7665
rect -14672 -10079 -12907 -9016
rect -17672 -11321 -16086 -10079
rect -20672 -12564 -19087 -11321
rect -23672 -13806 -22086 -12564
tri -23672 -15188 -22290 -13806 ne
rect -22290 -13978 -22086 -13806
tri -22086 -13978 -20672 -12564 sw
tri -20672 -13978 -19258 -12564 ne
rect -19258 -12736 -19087 -12564
tri -19087 -12736 -17672 -11321 sw
tri -17672 -12736 -16257 -11321 ne
rect -16257 -11493 -16086 -11321
tri -16086 -11493 -14672 -10079 sw
tri -14672 -11493 -13258 -10079 ne
rect -13258 -10251 -12907 -10079
tri -12907 -10251 -11672 -9016 sw
tri -11492 -10251 -10257 -9016 ne
rect -10257 -10150 -10015 -9016
tri -10015 -10150 -7530 -7665 sw
tri 7601 -10079 10429 -7251 se
rect 10429 -8493 12015 -7251
tri 12015 -8493 13257 -7251 nw
tri 13430 -8493 14672 -7251 se
rect 14672 -8493 16086 -7251
rect 10429 -9736 10772 -8493
tri 10772 -9736 12015 -8493 nw
tri 12187 -9736 13430 -8493 se
rect 13430 -8665 16086 -8493
tri 16086 -8665 17500 -7251 nw
tri 17500 -8665 18500 -7665 se
rect 18500 -8493 20500 8493
rect 18500 -8665 19257 -8493
rect 13430 -9736 15015 -8665
tri 15015 -9736 16086 -8665 nw
tri 16429 -9736 17500 -8665 se
rect 17500 -9736 19257 -8665
tri 19257 -9736 20500 -8493 nw
tri 20672 -9736 21500 -8908 se
rect 21500 -9736 23500 9736
rect 24500 5000 26500 10978
rect 24500 3000 27500 5000
tri 10429 -10079 10772 -9736 nw
tri 11844 -10079 12187 -9736 se
rect 12187 -10079 13773 -9736
rect -10257 -10251 -7530 -10150
rect -13258 -11493 -11672 -10251
rect -16257 -12736 -14672 -11493
rect -19258 -13978 -17672 -12736
rect -22290 -15188 -20672 -13978
tri -22290 -16634 -20844 -15188 ne
rect -20844 -15392 -20672 -15188
tri -20672 -15392 -19258 -13978 sw
tri -19258 -15392 -17844 -13978 ne
rect -17844 -14149 -17672 -13978
tri -17672 -14149 -16259 -12736 sw
tri -16257 -14149 -14844 -12736 ne
rect -14844 -12907 -14672 -12736
tri -14672 -12907 -13258 -11493 sw
tri -13258 -12907 -11844 -11493 ne
rect -11844 -11664 -11672 -11493
tri -11672 -11664 -10259 -10251 sw
tri -10257 -11664 -8844 -10251 ne
rect -8844 -11664 -7530 -10251
rect -11844 -12907 -10259 -11664
rect -14844 -14149 -13258 -12907
rect -17844 -15392 -16259 -14149
rect -20844 -16634 -19258 -15392
tri -20844 -18016 -19462 -16634 ne
rect -19462 -16806 -19258 -16634
tri -19258 -16806 -17844 -15392 sw
tri -17844 -16806 -16430 -15392 ne
rect -16430 -15564 -16259 -15392
tri -16259 -15564 -14844 -14149 sw
tri -14844 -15564 -13429 -14149 ne
rect -13429 -14321 -13258 -14149
tri -13258 -14321 -11844 -12907 sw
tri -11844 -14321 -10430 -12907 ne
rect -10430 -13079 -10259 -12907
tri -10259 -13079 -8844 -11664 sw
tri -8844 -12907 -7601 -11664 ne
rect -7601 -12500 -7530 -11664
tri -7530 -12500 -5180 -10150 sw
tri 5180 -12500 7601 -10079 se
rect 7601 -11321 9187 -10079
tri 9187 -11321 10429 -10079 nw
tri 10602 -11321 11844 -10079 se
rect 11844 -10978 13773 -10079
tri 13773 -10978 15015 -9736 nw
tri 15187 -10978 16429 -9736 se
rect 16429 -10978 18015 -9736
tri 18015 -10978 19257 -9736 nw
tri 19430 -10978 20672 -9736 se
rect 20672 -10978 22086 -9736
rect 11844 -11321 12391 -10978
rect 7601 -12500 7944 -11321
rect -7601 -12564 7944 -12500
tri 7944 -12564 9187 -11321 nw
tri 9359 -12564 10602 -11321 se
rect 10602 -12360 12391 -11321
tri 12391 -12360 13773 -10978 nw
tri 13805 -12360 15187 -10978 se
rect 15187 -12360 16633 -10978
tri 16633 -12360 18015 -10978 nw
tri 18048 -12360 19430 -10978 se
rect 19430 -11150 22086 -10978
tri 22086 -11150 23500 -9736 nw
rect 24500 -5000 27500 -3000
tri 23500 -11150 24500 -10150 se
rect 24500 -10978 26500 -5000
rect 24500 -11150 25118 -10978
rect 19430 -12360 20876 -11150
tri 20876 -12360 22086 -11150 nw
tri 22290 -12360 23500 -11150 se
rect 23500 -12360 25118 -11150
tri 25118 -12360 26500 -10978 nw
rect 10602 -12564 11493 -12360
rect -7601 -12907 6702 -12564
rect -10430 -14149 -8844 -13079
tri -8844 -14149 -7774 -13079 sw
tri -7601 -14149 -6359 -12907 ne
rect -6359 -13806 6702 -12907
tri 6702 -13806 7944 -12564 nw
tri 8117 -13806 9359 -12564 se
rect 9359 -13258 11493 -12564
tri 11493 -13258 12391 -12360 nw
tri 12907 -13258 13805 -12360 se
rect 13805 -13258 15562 -12360
rect 9359 -13806 10079 -13258
rect -6359 -14149 6008 -13806
rect -10430 -14321 -7774 -14149
rect -13429 -15564 -11844 -14321
rect -16430 -16806 -14844 -15564
rect -19462 -18016 -17844 -16806
tri -19462 -19628 -17850 -18016 ne
rect -17850 -18220 -17844 -18016
tri -17844 -18220 -16430 -16806 sw
tri -16430 -18220 -15016 -16806 ne
rect -15016 -16977 -14844 -16806
tri -14844 -16977 -13431 -15564 sw
tri -13429 -16977 -12016 -15564 ne
rect -12016 -15735 -11844 -15564
tri -11844 -15735 -10430 -14321 sw
tri -10430 -15735 -9016 -14321 ne
rect -9016 -15500 -7774 -14321
tri -7774 -15500 -6423 -14149 sw
tri -6359 -14500 -6008 -14149 ne
rect -6008 -14500 6008 -14149
tri 6008 -14500 6702 -13806 nw
tri 7423 -14500 8117 -13806 se
rect 8117 -14500 10079 -13806
tri 6423 -15500 7423 -14500 se
rect 7423 -14672 10079 -14500
tri 10079 -14672 11493 -13258 nw
tri 11493 -14672 12907 -13258 se
rect 12907 -13431 15562 -13258
tri 15562 -13431 16633 -12360 nw
tri 16977 -13431 18048 -12360 se
rect 18048 -13431 19634 -12360
rect 12907 -14672 14149 -13431
rect 7423 -15500 8665 -14672
rect -9016 -15735 -1085 -15500
rect -12016 -16977 -10430 -15735
rect -15016 -18220 -13431 -16977
rect -17850 -19628 -16430 -18220
tri -17850 -20844 -16634 -19628 ne
rect -16634 -19634 -16430 -19628
tri -16430 -19634 -15016 -18220 sw
tri -15016 -19634 -13602 -18220 ne
rect -13602 -18392 -13431 -18220
tri -13431 -18392 -12016 -16977 sw
tri -12016 -18392 -10601 -16977 ne
rect -10601 -17149 -10430 -16977
tri -10430 -17149 -9016 -15735 sw
tri -9016 -17149 -7602 -15735 ne
rect -7602 -17149 -1085 -15735
rect -10601 -18392 -9016 -17149
rect -13602 -19634 -12016 -18392
rect -16634 -20844 -15016 -19634
tri -16634 -22372 -15106 -20844 ne
rect -15106 -21048 -15016 -20844
tri -15016 -21048 -13602 -19634 sw
tri -13602 -21048 -12188 -19634 ne
rect -12188 -19805 -12016 -19634
tri -12016 -19805 -10603 -18392 sw
tri -10601 -19805 -9188 -18392 ne
rect -9188 -18500 -9016 -18392
tri -9016 -18500 -7665 -17149 sw
tri -7602 -17500 -7251 -17149 ne
rect -7251 -17500 -1085 -17149
tri -1915 -18220 -1195 -17500 ne
rect -1195 -18016 -1085 -17500
tri -1085 -18016 1431 -15500 sw
tri 1732 -15747 1979 -15500 se
rect 1979 -15747 8665 -15500
rect 1732 -16086 8665 -15747
tri 8665 -16086 10079 -14672 nw
tri 10079 -16086 11493 -14672 se
rect 11493 -14844 14149 -14672
tri 14149 -14844 15562 -13431 nw
tri 15564 -14844 16977 -13431 se
rect 16977 -13602 19634 -13431
tri 19634 -13602 20876 -12360 nw
tri 21048 -13602 22290 -12360 se
rect 16977 -14844 18220 -13602
rect 11493 -16086 12734 -14844
rect 1732 -17253 7251 -16086
tri 1732 -17500 1979 -17253 ne
rect 1979 -17500 7251 -17253
tri 7251 -17500 8665 -16086 nw
tri 8665 -17500 10079 -16086 se
rect 10079 -16259 12734 -16086
tri 12734 -16259 14149 -14844 nw
tri 14149 -16259 15564 -14844 se
rect 15564 -15016 18220 -14844
tri 18220 -15016 19634 -13602 nw
tri 19634 -15016 21048 -13602 se
rect 21048 -15016 22290 -13602
rect 15564 -16259 16806 -15016
rect 10079 -17500 11321 -16259
rect -1195 -18220 1431 -18016
rect -9188 -18747 -2202 -18500
tri -2202 -18747 -1955 -18500 sw
rect -9188 -19805 -1955 -18747
rect -12188 -21048 -10603 -19805
tri -10603 -21048 -9360 -19805 sw
tri -9188 -20500 -8493 -19805 ne
rect -8493 -20253 -1955 -19805
rect -8493 -20500 -2202 -20253
tri -2202 -20500 -1955 -20253 nw
tri -1195 -20500 1085 -18220 ne
rect 1085 -18500 1431 -18220
tri 1431 -18500 1915 -18016 sw
tri 7665 -18500 8665 -17500 se
rect 8665 -17672 11321 -17500
tri 11321 -17672 12734 -16259 nw
tri 12736 -17672 14149 -16259 se
rect 14149 -16430 16806 -16259
tri 16806 -16430 18220 -15016 nw
tri 19462 -15188 19634 -15016 se
rect 19634 -15188 22290 -15016
tri 22290 -15188 25118 -12360 nw
tri 18220 -16430 19462 -15188 se
rect 14149 -17672 15392 -16430
rect 8665 -18500 9906 -17672
rect 1085 -19087 9906 -18500
tri 9906 -19087 11321 -17672 nw
tri 11321 -19087 12736 -17672 se
rect 12736 -17844 15392 -17672
tri 15392 -17844 16806 -16430 nw
tri 16806 -17844 18220 -16430 se
rect 18220 -17844 19462 -16430
rect 12736 -19087 13978 -17844
rect 1085 -20500 8493 -19087
tri 8493 -20500 9906 -19087 nw
tri 9908 -20500 11321 -19087 se
rect 11321 -19258 13978 -19087
tri 13978 -19258 15392 -17844 nw
tri 16634 -18016 16806 -17844 se
rect 16806 -18016 19462 -17844
tri 19462 -18016 22290 -15188 nw
tri 15392 -19258 16634 -18016 se
rect 11321 -20500 12564 -19258
rect -15106 -22372 -13602 -21048
tri -15106 -23672 -13806 -22372 ne
rect -13806 -22462 -13602 -22372
tri -13602 -22462 -12188 -21048 sw
tri -12188 -22462 -10774 -21048 ne
rect -10774 -21500 -9360 -21048
tri -9360 -21500 -8908 -21048 sw
tri 8908 -21500 9908 -20500 se
rect 9908 -20672 12564 -20500
tri 12564 -20672 13978 -19258 nw
tri 13978 -20672 15392 -19258 se
rect 15392 -20672 16634 -19258
rect 9908 -21500 11150 -20672
rect -10774 -22462 -1085 -21500
rect -13806 -23672 -12188 -22462
tri -12188 -23672 -10978 -22462 sw
tri -10774 -23500 -9736 -22462 ne
rect -9736 -23500 -1085 -22462
tri -1915 -23672 -1743 -23500 ne
rect -1743 -23672 -1085 -23500
tri -1085 -23672 1087 -21500 sw
tri 1732 -21747 1979 -21500 se
rect 1979 -21747 11150 -21500
rect 1732 -22086 11150 -21747
tri 11150 -22086 12564 -20672 nw
tri 13806 -20844 13978 -20672 se
rect 13978 -20844 16634 -20672
tri 16634 -20844 19462 -18016 nw
tri 12564 -22086 13806 -20844 se
rect 1732 -23253 9736 -22086
tri 1732 -23500 1979 -23253 ne
rect 1979 -23500 9736 -23253
tri 9736 -23500 11150 -22086 nw
tri 11150 -23500 12564 -22086 se
rect 12564 -23500 13806 -22086
tri 10978 -23672 11150 -23500 se
rect 11150 -23672 13806 -23500
tri 13806 -23672 16634 -20844 nw
tri -13806 -26500 -10978 -23672 ne
tri -10978 -24500 -10150 -23672 sw
rect -10978 -24747 -2202 -24500
tri -2202 -24747 -1955 -24500 sw
rect -10978 -26253 -1955 -24747
rect -10978 -26500 -2202 -26253
tri -2202 -26500 -1955 -26253 nw
tri -1743 -26500 1085 -23672 ne
rect 1085 -24500 1087 -23672
tri 1087 -24500 1915 -23672 sw
tri 10150 -24500 10978 -23672 se
rect 1085 -26500 10978 -24500
tri 10978 -26500 13806 -23672 nw
<< properties >>
string FIXED_BBOX -26500 -26500 27500 26500
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__rf_test_coil2
string library sky130
string parameter m=1
string GDS_END 10379688
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10361220
<< end >>
