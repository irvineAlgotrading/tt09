magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< locali >>
rect 0 1397 1278 1431
rect 430 708 464 1167
rect 430 674 559 708
rect 875 674 909 708
rect 345 485 379 551
rect 212 361 246 427
rect 79 237 113 303
rect 0 -17 1278 17
use sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_5  sky130_sram_1kbyte_1rw1r_8x1024_8_pdriver_5_0
timestamp 1704896540
transform 1 0 478 0 1 0
box -36 -17 836 1471
use sky130_sram_1kbyte_1rw1r_8x1024_8_pnand3  sky130_sram_1kbyte_1rw1r_8x1024_8_pnand3_0
timestamp 1704896540
transform 1 0 0 0 1 0
box -36 -17 514 1471
<< labels >>
rlabel locali s 892 691 892 691 4 Z
rlabel locali s 96 270 96 270 4 A
rlabel locali s 229 394 229 394 4 B
rlabel locali s 362 518 362 518 4 C
rlabel locali s 639 0 639 0 4 gnd
rlabel locali s 639 1414 639 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1278 1414
string GDS_END 6089524
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 6088276
<< end >>
