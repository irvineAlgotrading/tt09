magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 519 366
<< mvpmos >>
rect 0 0 400 300
<< mvpdiff >>
rect -50 0 0 300
rect 400 0 450 300
<< poly >>
rect 0 300 400 326
rect 0 -26 400 0
<< metal1 >>
rect -51 -16 -5 258
rect 405 -16 451 258
use hvDFM1sd_CDNS_52468879185274  hvDFM1sd_CDNS_52468879185274_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 336
use hvDFM1sd_CDNS_52468879185274  hvDFM1sd_CDNS_52468879185274_1
timestamp 1704896540
transform 1 0 400 0 1 0
box -36 -36 89 336
<< labels >>
flabel comment s -28 121 -28 121 0 FreeSans 300 0 0 0 S
flabel comment s 428 121 428 121 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86838552
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86837534
<< end >>
