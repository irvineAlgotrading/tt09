magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 154
rect 125 0 128 154
<< via1 >>
rect 3 0 125 154
<< metal2 >>
rect 0 0 3 154
rect 125 0 128 154
<< properties >>
string GDS_END 85243784
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85242372
<< end >>
