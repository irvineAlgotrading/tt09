magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -1442 120 -694 483
rect 458 120 478 482
rect -2594 14 1034 120
rect 74 -348 94 14
rect -2088 -877 613 -869
rect -2263 -1578 613 -877
rect 1234 -988 3386 -548
rect 2622 -1119 3386 -988
rect 2622 -2005 3502 -1119
rect 1467 -3217 1831 -2749
<< pwell >>
rect -2556 852 1092 938
rect -1404 765 -732 852
rect -1388 551 -743 765
rect -2556 -804 996 -718
rect -2188 -1910 573 -1683
rect -2263 -1996 582 -1910
rect 4350 -2117 4684 -2013
rect 1505 -2379 1793 -2293
<< scnmos >>
rect -1309 577 -1279 745
rect -1223 577 -1193 745
rect -1137 577 -1107 745
rect -1059 577 -1029 745
rect -913 577 -883 745
<< scpmoshvt >>
rect -1309 195 -1279 447
rect -1231 195 -1201 447
rect -1141 195 -1111 447
rect -1055 195 -1025 447
rect -842 195 -812 447
<< mvnmos >>
rect -2109 -1849 -1989 -1709
rect -1933 -1849 -1813 -1709
rect -1757 -1849 -1637 -1709
rect -1581 -1849 -1461 -1709
rect -1206 -1849 -1086 -1709
rect -1030 -1849 -910 -1709
rect -741 -1849 -621 -1709
rect -565 -1849 -445 -1709
rect -273 -1849 -153 -1709
rect -97 -1849 23 -1709
rect 198 -1849 318 -1709
rect 374 -1849 494 -1709
<< mvpmos >>
rect -2109 -1243 -1989 -1043
rect -1933 -1243 -1813 -1043
rect -1757 -1243 -1637 -1043
rect -1581 -1243 -1461 -1043
rect -1206 -1243 -1086 -1043
rect -1030 -1243 -910 -1043
rect -741 -1243 -621 -1043
rect -565 -1243 -445 -1043
rect -273 -1243 -153 -1043
rect -97 -1243 23 -1043
rect 198 -1243 318 -1043
rect 374 -1243 494 -1043
rect -2109 -1511 -1989 -1311
rect -1933 -1511 -1813 -1311
rect -1757 -1511 -1637 -1311
rect -1581 -1511 -1461 -1311
rect -1206 -1511 -1086 -1311
rect -1030 -1511 -910 -1311
rect -741 -1511 -621 -1311
rect -565 -1511 -445 -1311
rect -273 -1511 -153 -1311
rect -97 -1511 23 -1311
rect 198 -1511 318 -1311
rect 374 -1511 494 -1311
<< ndiff >>
rect -1362 733 -1309 745
rect -1362 699 -1354 733
rect -1320 699 -1309 733
rect -1362 656 -1309 699
rect -1362 622 -1354 656
rect -1320 622 -1309 656
rect -1362 577 -1309 622
rect -1279 731 -1223 745
rect -1279 697 -1268 731
rect -1234 697 -1223 731
rect -1279 640 -1223 697
rect -1279 606 -1268 640
rect -1234 606 -1223 640
rect -1279 577 -1223 606
rect -1193 716 -1137 745
rect -1193 682 -1182 716
rect -1148 682 -1137 716
rect -1193 577 -1137 682
rect -1107 577 -1059 745
rect -1029 695 -913 745
rect -1029 661 -980 695
rect -946 661 -913 695
rect -1029 619 -913 661
rect -1029 585 -980 619
rect -946 585 -913 619
rect -1029 577 -913 585
rect -883 733 -769 745
rect -883 699 -811 733
rect -777 699 -769 733
rect -883 652 -769 699
rect -883 618 -811 652
rect -777 618 -769 652
rect -883 577 -769 618
<< pdiff >>
rect -1362 401 -1309 447
rect -1362 367 -1354 401
rect -1320 367 -1309 401
rect -1362 323 -1309 367
rect -1362 289 -1354 323
rect -1320 289 -1309 323
rect -1362 249 -1309 289
rect -1362 215 -1354 249
rect -1320 215 -1309 249
rect -1362 195 -1309 215
rect -1279 195 -1231 447
rect -1201 317 -1141 447
rect -1201 283 -1190 317
rect -1156 283 -1141 317
rect -1201 241 -1141 283
rect -1201 207 -1190 241
rect -1156 207 -1141 241
rect -1201 195 -1141 207
rect -1111 333 -1055 447
rect -1111 299 -1100 333
rect -1066 299 -1055 333
rect -1111 241 -1055 299
rect -1111 207 -1100 241
rect -1066 207 -1055 241
rect -1111 195 -1055 207
rect -1025 227 -953 447
rect -1025 195 -995 227
rect -1003 193 -995 195
rect -961 193 -953 227
rect -899 439 -842 447
rect -899 405 -887 439
rect -853 405 -842 439
rect -899 195 -842 405
rect -812 279 -759 447
rect -812 245 -801 279
rect -767 245 -759 279
rect -812 195 -759 245
rect -1003 175 -953 193
<< mvndiff >>
rect -2162 -1721 -2109 -1709
rect -2162 -1755 -2154 -1721
rect -2120 -1755 -2109 -1721
rect -2162 -1789 -2109 -1755
rect -2162 -1823 -2154 -1789
rect -2120 -1823 -2109 -1789
rect -2162 -1849 -2109 -1823
rect -1989 -1849 -1933 -1709
rect -1813 -1721 -1757 -1709
rect -1813 -1755 -1802 -1721
rect -1768 -1755 -1757 -1721
rect -1813 -1789 -1757 -1755
rect -1813 -1823 -1802 -1789
rect -1768 -1823 -1757 -1789
rect -1813 -1849 -1757 -1823
rect -1637 -1849 -1581 -1709
rect -1461 -1721 -1408 -1709
rect -1461 -1755 -1450 -1721
rect -1416 -1755 -1408 -1721
rect -1461 -1789 -1408 -1755
rect -1461 -1823 -1450 -1789
rect -1416 -1823 -1408 -1789
rect -1461 -1849 -1408 -1823
rect -1259 -1721 -1206 -1709
rect -1259 -1755 -1251 -1721
rect -1217 -1755 -1206 -1721
rect -1259 -1789 -1206 -1755
rect -1259 -1823 -1251 -1789
rect -1217 -1823 -1206 -1789
rect -1259 -1849 -1206 -1823
rect -1086 -1849 -1030 -1709
rect -910 -1721 -857 -1709
rect -910 -1755 -899 -1721
rect -865 -1755 -857 -1721
rect -910 -1789 -857 -1755
rect -910 -1823 -899 -1789
rect -865 -1823 -857 -1789
rect -910 -1849 -857 -1823
rect -794 -1721 -741 -1709
rect -794 -1755 -786 -1721
rect -752 -1755 -741 -1721
rect -794 -1789 -741 -1755
rect -794 -1823 -786 -1789
rect -752 -1823 -741 -1789
rect -794 -1849 -741 -1823
rect -621 -1849 -565 -1709
rect -445 -1721 -392 -1709
rect -445 -1755 -434 -1721
rect -400 -1755 -392 -1721
rect -445 -1789 -392 -1755
rect -445 -1823 -434 -1789
rect -400 -1823 -392 -1789
rect -445 -1849 -392 -1823
rect -326 -1721 -273 -1709
rect -326 -1755 -318 -1721
rect -284 -1755 -273 -1721
rect -326 -1789 -273 -1755
rect -326 -1823 -318 -1789
rect -284 -1823 -273 -1789
rect -326 -1849 -273 -1823
rect -153 -1721 -97 -1709
rect -153 -1755 -142 -1721
rect -108 -1755 -97 -1721
rect -153 -1789 -97 -1755
rect -153 -1823 -142 -1789
rect -108 -1823 -97 -1789
rect -153 -1849 -97 -1823
rect 23 -1721 79 -1709
rect 23 -1755 34 -1721
rect 68 -1755 79 -1721
rect 23 -1789 79 -1755
rect 23 -1823 34 -1789
rect 68 -1823 79 -1789
rect 23 -1849 79 -1823
rect 142 -1721 198 -1709
rect 142 -1755 153 -1721
rect 187 -1755 198 -1721
rect 142 -1789 198 -1755
rect 142 -1823 153 -1789
rect 187 -1823 198 -1789
rect 142 -1849 198 -1823
rect 318 -1721 374 -1709
rect 318 -1755 329 -1721
rect 363 -1755 374 -1721
rect 318 -1789 374 -1755
rect 318 -1823 329 -1789
rect 363 -1823 374 -1789
rect 318 -1849 374 -1823
rect 494 -1721 547 -1709
rect 494 -1755 505 -1721
rect 539 -1755 547 -1721
rect 494 -1789 547 -1755
rect 494 -1823 505 -1789
rect 539 -1823 547 -1789
rect 494 -1849 547 -1823
<< mvpdiff >>
rect -2162 -1061 -2109 -1043
rect -2162 -1095 -2154 -1061
rect -2120 -1095 -2109 -1061
rect -2162 -1129 -2109 -1095
rect -2162 -1163 -2154 -1129
rect -2120 -1163 -2109 -1129
rect -2162 -1197 -2109 -1163
rect -2162 -1231 -2154 -1197
rect -2120 -1231 -2109 -1197
rect -2162 -1243 -2109 -1231
rect -1989 -1061 -1933 -1043
rect -1989 -1095 -1978 -1061
rect -1944 -1095 -1933 -1061
rect -1989 -1129 -1933 -1095
rect -1989 -1163 -1978 -1129
rect -1944 -1163 -1933 -1129
rect -1989 -1197 -1933 -1163
rect -1989 -1231 -1978 -1197
rect -1944 -1231 -1933 -1197
rect -1989 -1243 -1933 -1231
rect -1813 -1061 -1757 -1043
rect -1813 -1095 -1802 -1061
rect -1768 -1095 -1757 -1061
rect -1813 -1129 -1757 -1095
rect -1813 -1163 -1802 -1129
rect -1768 -1163 -1757 -1129
rect -1813 -1197 -1757 -1163
rect -1813 -1231 -1802 -1197
rect -1768 -1231 -1757 -1197
rect -1813 -1243 -1757 -1231
rect -1637 -1061 -1581 -1043
rect -1637 -1095 -1626 -1061
rect -1592 -1095 -1581 -1061
rect -1637 -1129 -1581 -1095
rect -1637 -1163 -1626 -1129
rect -1592 -1163 -1581 -1129
rect -1637 -1197 -1581 -1163
rect -1637 -1231 -1626 -1197
rect -1592 -1231 -1581 -1197
rect -1637 -1243 -1581 -1231
rect -1461 -1061 -1408 -1043
rect -1461 -1095 -1450 -1061
rect -1416 -1095 -1408 -1061
rect -1461 -1129 -1408 -1095
rect -1461 -1163 -1450 -1129
rect -1416 -1163 -1408 -1129
rect -1461 -1197 -1408 -1163
rect -1461 -1231 -1450 -1197
rect -1416 -1231 -1408 -1197
rect -1461 -1243 -1408 -1231
rect -1259 -1061 -1206 -1043
rect -1259 -1095 -1251 -1061
rect -1217 -1095 -1206 -1061
rect -1259 -1129 -1206 -1095
rect -1259 -1163 -1251 -1129
rect -1217 -1163 -1206 -1129
rect -1259 -1197 -1206 -1163
rect -1259 -1231 -1251 -1197
rect -1217 -1231 -1206 -1197
rect -1259 -1243 -1206 -1231
rect -1086 -1061 -1030 -1043
rect -1086 -1095 -1075 -1061
rect -1041 -1095 -1030 -1061
rect -1086 -1129 -1030 -1095
rect -1086 -1163 -1075 -1129
rect -1041 -1163 -1030 -1129
rect -1086 -1197 -1030 -1163
rect -1086 -1231 -1075 -1197
rect -1041 -1231 -1030 -1197
rect -1086 -1243 -1030 -1231
rect -910 -1061 -857 -1043
rect -910 -1095 -899 -1061
rect -865 -1095 -857 -1061
rect -910 -1129 -857 -1095
rect -910 -1163 -899 -1129
rect -865 -1163 -857 -1129
rect -910 -1197 -857 -1163
rect -910 -1231 -899 -1197
rect -865 -1231 -857 -1197
rect -910 -1243 -857 -1231
rect -794 -1061 -741 -1043
rect -794 -1095 -786 -1061
rect -752 -1095 -741 -1061
rect -794 -1129 -741 -1095
rect -794 -1163 -786 -1129
rect -752 -1163 -741 -1129
rect -794 -1197 -741 -1163
rect -794 -1231 -786 -1197
rect -752 -1231 -741 -1197
rect -794 -1243 -741 -1231
rect -621 -1061 -565 -1043
rect -621 -1095 -610 -1061
rect -576 -1095 -565 -1061
rect -621 -1129 -565 -1095
rect -621 -1163 -610 -1129
rect -576 -1163 -565 -1129
rect -621 -1197 -565 -1163
rect -621 -1231 -610 -1197
rect -576 -1231 -565 -1197
rect -621 -1243 -565 -1231
rect -445 -1061 -392 -1043
rect -445 -1095 -434 -1061
rect -400 -1095 -392 -1061
rect -445 -1129 -392 -1095
rect -445 -1163 -434 -1129
rect -400 -1163 -392 -1129
rect -445 -1197 -392 -1163
rect -445 -1231 -434 -1197
rect -400 -1231 -392 -1197
rect -445 -1243 -392 -1231
rect -326 -1061 -273 -1043
rect -326 -1095 -318 -1061
rect -284 -1095 -273 -1061
rect -326 -1129 -273 -1095
rect -326 -1163 -318 -1129
rect -284 -1163 -273 -1129
rect -326 -1197 -273 -1163
rect -326 -1231 -318 -1197
rect -284 -1231 -273 -1197
rect -326 -1243 -273 -1231
rect -153 -1061 -97 -1043
rect -153 -1095 -142 -1061
rect -108 -1095 -97 -1061
rect -153 -1129 -97 -1095
rect -153 -1163 -142 -1129
rect -108 -1163 -97 -1129
rect -153 -1197 -97 -1163
rect -153 -1231 -142 -1197
rect -108 -1231 -97 -1197
rect -153 -1243 -97 -1231
rect 23 -1061 76 -1043
rect 23 -1095 34 -1061
rect 68 -1095 76 -1061
rect 23 -1129 76 -1095
rect 23 -1163 34 -1129
rect 68 -1163 76 -1129
rect 23 -1197 76 -1163
rect 23 -1231 34 -1197
rect 68 -1231 76 -1197
rect 23 -1243 76 -1231
rect 145 -1061 198 -1043
rect 145 -1095 153 -1061
rect 187 -1095 198 -1061
rect 145 -1129 198 -1095
rect 145 -1163 153 -1129
rect 187 -1163 198 -1129
rect 145 -1197 198 -1163
rect 145 -1231 153 -1197
rect 187 -1231 198 -1197
rect 145 -1243 198 -1231
rect 318 -1061 374 -1043
rect 318 -1095 329 -1061
rect 363 -1095 374 -1061
rect 318 -1129 374 -1095
rect 318 -1163 329 -1129
rect 363 -1163 374 -1129
rect 318 -1197 374 -1163
rect 318 -1231 329 -1197
rect 363 -1231 374 -1197
rect 318 -1243 374 -1231
rect 494 -1061 547 -1043
rect 494 -1095 505 -1061
rect 539 -1095 547 -1061
rect 494 -1129 547 -1095
rect 494 -1163 505 -1129
rect 539 -1163 547 -1129
rect 494 -1197 547 -1163
rect 494 -1231 505 -1197
rect 539 -1231 547 -1197
rect 494 -1243 547 -1231
rect -2162 -1323 -2109 -1311
rect -2162 -1357 -2154 -1323
rect -2120 -1357 -2109 -1323
rect -2162 -1391 -2109 -1357
rect -2162 -1425 -2154 -1391
rect -2120 -1425 -2109 -1391
rect -2162 -1459 -2109 -1425
rect -2162 -1493 -2154 -1459
rect -2120 -1493 -2109 -1459
rect -2162 -1511 -2109 -1493
rect -1989 -1323 -1933 -1311
rect -1989 -1357 -1978 -1323
rect -1944 -1357 -1933 -1323
rect -1989 -1391 -1933 -1357
rect -1989 -1425 -1978 -1391
rect -1944 -1425 -1933 -1391
rect -1989 -1459 -1933 -1425
rect -1989 -1493 -1978 -1459
rect -1944 -1493 -1933 -1459
rect -1989 -1511 -1933 -1493
rect -1813 -1323 -1757 -1311
rect -1813 -1357 -1802 -1323
rect -1768 -1357 -1757 -1323
rect -1813 -1391 -1757 -1357
rect -1813 -1425 -1802 -1391
rect -1768 -1425 -1757 -1391
rect -1813 -1459 -1757 -1425
rect -1813 -1493 -1802 -1459
rect -1768 -1493 -1757 -1459
rect -1813 -1511 -1757 -1493
rect -1637 -1323 -1581 -1311
rect -1637 -1357 -1626 -1323
rect -1592 -1357 -1581 -1323
rect -1637 -1391 -1581 -1357
rect -1637 -1425 -1626 -1391
rect -1592 -1425 -1581 -1391
rect -1637 -1459 -1581 -1425
rect -1637 -1493 -1626 -1459
rect -1592 -1493 -1581 -1459
rect -1637 -1511 -1581 -1493
rect -1461 -1323 -1408 -1311
rect -1461 -1357 -1450 -1323
rect -1416 -1357 -1408 -1323
rect -1461 -1391 -1408 -1357
rect -1461 -1425 -1450 -1391
rect -1416 -1425 -1408 -1391
rect -1461 -1459 -1408 -1425
rect -1461 -1493 -1450 -1459
rect -1416 -1493 -1408 -1459
rect -1461 -1511 -1408 -1493
rect -1259 -1323 -1206 -1311
rect -1259 -1357 -1251 -1323
rect -1217 -1357 -1206 -1323
rect -1259 -1391 -1206 -1357
rect -1259 -1425 -1251 -1391
rect -1217 -1425 -1206 -1391
rect -1259 -1459 -1206 -1425
rect -1259 -1493 -1251 -1459
rect -1217 -1493 -1206 -1459
rect -1259 -1511 -1206 -1493
rect -1086 -1323 -1030 -1311
rect -1086 -1357 -1075 -1323
rect -1041 -1357 -1030 -1323
rect -1086 -1391 -1030 -1357
rect -1086 -1425 -1075 -1391
rect -1041 -1425 -1030 -1391
rect -1086 -1459 -1030 -1425
rect -1086 -1493 -1075 -1459
rect -1041 -1493 -1030 -1459
rect -1086 -1511 -1030 -1493
rect -910 -1323 -857 -1311
rect -910 -1357 -899 -1323
rect -865 -1357 -857 -1323
rect -910 -1391 -857 -1357
rect -910 -1425 -899 -1391
rect -865 -1425 -857 -1391
rect -910 -1459 -857 -1425
rect -910 -1493 -899 -1459
rect -865 -1493 -857 -1459
rect -910 -1511 -857 -1493
rect -794 -1323 -741 -1311
rect -794 -1357 -786 -1323
rect -752 -1357 -741 -1323
rect -794 -1391 -741 -1357
rect -794 -1425 -786 -1391
rect -752 -1425 -741 -1391
rect -794 -1459 -741 -1425
rect -794 -1493 -786 -1459
rect -752 -1493 -741 -1459
rect -794 -1511 -741 -1493
rect -621 -1323 -565 -1311
rect -621 -1357 -610 -1323
rect -576 -1357 -565 -1323
rect -621 -1391 -565 -1357
rect -621 -1425 -610 -1391
rect -576 -1425 -565 -1391
rect -621 -1459 -565 -1425
rect -621 -1493 -610 -1459
rect -576 -1493 -565 -1459
rect -621 -1511 -565 -1493
rect -445 -1323 -392 -1311
rect -445 -1357 -434 -1323
rect -400 -1357 -392 -1323
rect -445 -1391 -392 -1357
rect -445 -1425 -434 -1391
rect -400 -1425 -392 -1391
rect -445 -1459 -392 -1425
rect -445 -1493 -434 -1459
rect -400 -1493 -392 -1459
rect -445 -1511 -392 -1493
rect -326 -1323 -273 -1311
rect -326 -1357 -318 -1323
rect -284 -1357 -273 -1323
rect -326 -1391 -273 -1357
rect -326 -1425 -318 -1391
rect -284 -1425 -273 -1391
rect -326 -1459 -273 -1425
rect -326 -1493 -318 -1459
rect -284 -1493 -273 -1459
rect -326 -1511 -273 -1493
rect -153 -1323 -97 -1311
rect -153 -1357 -142 -1323
rect -108 -1357 -97 -1323
rect -153 -1391 -97 -1357
rect -153 -1425 -142 -1391
rect -108 -1425 -97 -1391
rect -153 -1511 -97 -1425
rect 23 -1323 76 -1311
rect 23 -1357 34 -1323
rect 68 -1357 76 -1323
rect 23 -1391 76 -1357
rect 23 -1425 34 -1391
rect 68 -1425 76 -1391
rect 23 -1459 76 -1425
rect 23 -1493 34 -1459
rect 68 -1493 76 -1459
rect 23 -1511 76 -1493
rect 145 -1323 198 -1311
rect 145 -1357 153 -1323
rect 187 -1357 198 -1323
rect 145 -1391 198 -1357
rect 145 -1425 153 -1391
rect 187 -1425 198 -1391
rect 145 -1459 198 -1425
rect 145 -1493 153 -1459
rect 187 -1493 198 -1459
rect 145 -1511 198 -1493
rect 318 -1323 374 -1311
rect 318 -1357 329 -1323
rect 363 -1357 374 -1323
rect 318 -1391 374 -1357
rect 318 -1425 329 -1391
rect 363 -1425 374 -1391
rect 318 -1511 374 -1425
rect 494 -1323 547 -1311
rect 494 -1357 505 -1323
rect 539 -1357 547 -1323
rect 494 -1391 547 -1357
rect 494 -1425 505 -1391
rect 539 -1425 547 -1391
rect 494 -1459 547 -1425
rect 494 -1493 505 -1459
rect 539 -1493 547 -1459
rect 494 -1511 547 -1493
<< ndiffc >>
rect -1354 699 -1320 733
rect -1354 622 -1320 656
rect -1268 697 -1234 731
rect -1268 606 -1234 640
rect -1182 682 -1148 716
rect -980 661 -946 695
rect -980 585 -946 619
rect -811 699 -777 733
rect -811 618 -777 652
<< pdiffc >>
rect -1354 367 -1320 401
rect -1354 289 -1320 323
rect -1354 215 -1320 249
rect -1190 283 -1156 317
rect -1190 207 -1156 241
rect -1100 299 -1066 333
rect -1100 207 -1066 241
rect -995 193 -961 227
rect -887 405 -853 439
rect -801 245 -767 279
<< mvndiffc >>
rect -2154 -1755 -2120 -1721
rect -2154 -1823 -2120 -1789
rect -1802 -1755 -1768 -1721
rect -1802 -1823 -1768 -1789
rect -1450 -1755 -1416 -1721
rect -1450 -1823 -1416 -1789
rect -1251 -1755 -1217 -1721
rect -1251 -1823 -1217 -1789
rect -899 -1755 -865 -1721
rect -899 -1823 -865 -1789
rect -786 -1755 -752 -1721
rect -786 -1823 -752 -1789
rect -434 -1755 -400 -1721
rect -434 -1823 -400 -1789
rect -318 -1755 -284 -1721
rect -318 -1823 -284 -1789
rect -142 -1755 -108 -1721
rect -142 -1823 -108 -1789
rect 34 -1755 68 -1721
rect 34 -1823 68 -1789
rect 153 -1755 187 -1721
rect 153 -1823 187 -1789
rect 329 -1755 363 -1721
rect 329 -1823 363 -1789
rect 505 -1755 539 -1721
rect 505 -1823 539 -1789
<< mvpdiffc >>
rect -2154 -1095 -2120 -1061
rect -2154 -1163 -2120 -1129
rect -2154 -1231 -2120 -1197
rect -1978 -1095 -1944 -1061
rect -1978 -1163 -1944 -1129
rect -1978 -1231 -1944 -1197
rect -1802 -1095 -1768 -1061
rect -1802 -1163 -1768 -1129
rect -1802 -1231 -1768 -1197
rect -1626 -1095 -1592 -1061
rect -1626 -1163 -1592 -1129
rect -1626 -1231 -1592 -1197
rect -1450 -1095 -1416 -1061
rect -1450 -1163 -1416 -1129
rect -1450 -1231 -1416 -1197
rect -1251 -1095 -1217 -1061
rect -1251 -1163 -1217 -1129
rect -1251 -1231 -1217 -1197
rect -1075 -1095 -1041 -1061
rect -1075 -1163 -1041 -1129
rect -1075 -1231 -1041 -1197
rect -899 -1095 -865 -1061
rect -899 -1163 -865 -1129
rect -899 -1231 -865 -1197
rect -786 -1095 -752 -1061
rect -786 -1163 -752 -1129
rect -786 -1231 -752 -1197
rect -610 -1095 -576 -1061
rect -610 -1163 -576 -1129
rect -610 -1231 -576 -1197
rect -434 -1095 -400 -1061
rect -434 -1163 -400 -1129
rect -434 -1231 -400 -1197
rect -318 -1095 -284 -1061
rect -318 -1163 -284 -1129
rect -318 -1231 -284 -1197
rect -142 -1095 -108 -1061
rect -142 -1163 -108 -1129
rect -142 -1231 -108 -1197
rect 34 -1095 68 -1061
rect 34 -1163 68 -1129
rect 34 -1231 68 -1197
rect 153 -1095 187 -1061
rect 153 -1163 187 -1129
rect 153 -1231 187 -1197
rect 329 -1095 363 -1061
rect 329 -1163 363 -1129
rect 329 -1231 363 -1197
rect 505 -1095 539 -1061
rect 505 -1163 539 -1129
rect 505 -1231 539 -1197
rect -2154 -1357 -2120 -1323
rect -2154 -1425 -2120 -1391
rect -2154 -1493 -2120 -1459
rect -1978 -1357 -1944 -1323
rect -1978 -1425 -1944 -1391
rect -1978 -1493 -1944 -1459
rect -1802 -1357 -1768 -1323
rect -1802 -1425 -1768 -1391
rect -1802 -1493 -1768 -1459
rect -1626 -1357 -1592 -1323
rect -1626 -1425 -1592 -1391
rect -1626 -1493 -1592 -1459
rect -1450 -1357 -1416 -1323
rect -1450 -1425 -1416 -1391
rect -1450 -1493 -1416 -1459
rect -1251 -1357 -1217 -1323
rect -1251 -1425 -1217 -1391
rect -1251 -1493 -1217 -1459
rect -1075 -1357 -1041 -1323
rect -1075 -1425 -1041 -1391
rect -1075 -1493 -1041 -1459
rect -899 -1357 -865 -1323
rect -899 -1425 -865 -1391
rect -899 -1493 -865 -1459
rect -786 -1357 -752 -1323
rect -786 -1425 -752 -1391
rect -786 -1493 -752 -1459
rect -610 -1357 -576 -1323
rect -610 -1425 -576 -1391
rect -610 -1493 -576 -1459
rect -434 -1357 -400 -1323
rect -434 -1425 -400 -1391
rect -434 -1493 -400 -1459
rect -318 -1357 -284 -1323
rect -318 -1425 -284 -1391
rect -318 -1493 -284 -1459
rect -142 -1357 -108 -1323
rect -142 -1425 -108 -1391
rect 34 -1357 68 -1323
rect 34 -1425 68 -1391
rect 34 -1493 68 -1459
rect 153 -1357 187 -1323
rect 153 -1425 187 -1391
rect 153 -1493 187 -1459
rect 329 -1357 363 -1323
rect 329 -1425 363 -1391
rect 505 -1357 539 -1323
rect 505 -1425 539 -1391
rect 505 -1493 539 -1459
<< psubdiff >>
rect -2530 878 -2506 912
rect -2472 878 -2365 912
rect -2331 878 -2224 912
rect -2190 878 -2083 912
rect -2049 878 -1942 912
rect -1908 878 -1801 912
rect -1767 878 -1660 912
rect -1626 878 -1519 912
rect -1485 878 -1378 912
rect -1344 878 -1237 912
rect -1203 878 -1096 912
rect -1062 878 -955 912
rect -921 878 -814 912
rect -780 878 -673 912
rect -639 878 -532 912
rect -498 878 -392 912
rect -358 878 -252 912
rect -218 878 -112 912
rect -78 878 28 912
rect 62 878 168 912
rect 202 878 308 912
rect 342 878 448 912
rect 482 878 588 912
rect 622 878 728 912
rect 762 878 868 912
rect 902 878 1008 912
rect 1042 878 1066 912
rect -2530 -778 -2506 -744
rect -2472 -778 -2369 -744
rect -2335 -778 -2232 -744
rect -2198 -778 -2095 -744
rect -2061 -778 -1958 -744
rect -1924 -778 -1821 -744
rect -1787 -778 -1684 -744
rect -1650 -778 -1547 -744
rect -1513 -778 -1410 -744
rect -1376 -778 -1273 -744
rect -1239 -778 -1136 -744
rect -1102 -778 -999 -744
rect -965 -778 -862 -744
rect -828 -778 -725 -744
rect -691 -778 -588 -744
rect -554 -778 -451 -744
rect -417 -778 -314 -744
rect -280 -778 -177 -744
rect -143 -778 -40 -744
rect -6 -778 96 -744
rect 130 -778 232 -744
rect 266 -778 368 -744
rect 402 -778 504 -744
rect 538 -778 640 -744
rect 674 -778 776 -744
rect 810 -778 912 -744
rect 946 -778 970 -744
rect 1531 -2353 1555 -2319
rect 1589 -2353 1709 -2319
rect 1743 -2353 1767 -2319
<< nsubdiff >>
rect -2558 50 -2534 84
rect -2500 50 -2465 84
rect -2431 50 -2396 84
rect -2362 50 -2327 84
rect -2293 50 -2258 84
rect -2224 50 -2189 84
rect -2155 50 -2120 84
rect -2086 50 -2052 84
rect -2018 50 -1984 84
rect -1950 50 -1916 84
rect -1882 50 -1848 84
rect -1814 50 -1780 84
rect -1746 50 -1712 84
rect -1678 50 -1644 84
rect -1610 50 -1576 84
rect -1542 50 -1508 84
rect -1474 50 -1440 84
rect -1406 50 -1372 84
rect -1338 50 -1304 84
rect -1270 50 -1236 84
rect -1202 50 -1168 84
rect -1134 50 -1100 84
rect -1066 50 -1032 84
rect -998 50 -964 84
rect -930 50 -896 84
rect -862 50 -828 84
rect -794 50 -760 84
rect -726 50 -692 84
rect -658 50 -624 84
rect -590 50 -556 84
rect -522 50 -488 84
rect -454 50 -420 84
rect -386 50 -352 84
rect -318 50 -284 84
rect -250 50 -216 84
rect -182 50 -148 84
rect -114 50 -80 84
rect -46 50 -12 84
rect 22 50 56 84
rect 90 50 124 84
rect 158 50 192 84
rect 226 50 260 84
rect 294 50 328 84
rect 362 50 396 84
rect 430 50 464 84
rect 498 50 532 84
rect 566 50 600 84
rect 634 50 668 84
rect 702 50 736 84
rect 770 50 804 84
rect 838 50 872 84
rect 906 50 940 84
rect 974 50 998 84
rect 1531 -3181 1555 -3147
rect 1589 -3181 1632 -3147
rect 1666 -3181 1709 -3147
rect 1743 -3181 1767 -3147
<< mvpsubdiff >>
rect -2237 -1970 -2213 -1936
rect -2179 -1970 -2070 -1936
rect -2036 -1970 -1927 -1936
rect -1893 -1970 -1784 -1936
rect -1750 -1970 -1641 -1936
rect -1607 -1970 -1498 -1936
rect -1464 -1970 -1355 -1936
rect -1321 -1970 -1212 -1936
rect -1178 -1970 -1069 -1936
rect -1035 -1970 -926 -1936
rect -892 -1970 -783 -1936
rect -749 -1970 -640 -1936
rect -606 -1970 -497 -1936
rect -463 -1970 -354 -1936
rect -320 -1970 -212 -1936
rect -178 -1970 -70 -1936
rect -36 -1970 72 -1936
rect 106 -1970 214 -1936
rect 248 -1970 356 -1936
rect 390 -1970 498 -1936
rect 532 -1970 556 -1936
<< mvnsubdiff >>
rect -2022 -969 -1998 -935
rect -1964 -969 -1928 -935
rect -1894 -969 -1858 -935
rect -1824 -969 -1788 -935
rect -1754 -969 -1719 -935
rect -1685 -969 -1650 -935
rect -1616 -969 -1581 -935
rect -1547 -969 -1512 -935
rect -1478 -969 -1443 -935
rect -1409 -969 -1374 -935
rect -1340 -969 -1305 -935
rect -1271 -969 -1236 -935
rect -1202 -969 -1167 -935
rect -1133 -969 -1098 -935
rect -1064 -969 -1029 -935
rect -995 -969 -960 -935
rect -926 -969 -891 -935
rect -857 -969 -822 -935
rect -788 -969 -753 -935
rect -719 -969 -684 -935
rect -650 -969 -615 -935
rect -581 -969 -546 -935
rect -512 -969 -477 -935
rect -443 -969 -408 -935
rect -374 -969 -339 -935
rect -305 -969 -270 -935
rect -236 -969 -201 -935
rect -167 -969 -132 -935
rect -98 -969 -63 -935
rect -29 -969 6 -935
rect 40 -969 75 -935
rect 109 -969 144 -935
rect 178 -969 213 -935
rect 247 -969 282 -935
rect 316 -969 351 -935
rect 385 -969 420 -935
rect 454 -969 489 -935
rect 523 -969 547 -935
<< psubdiffcont >>
rect -2506 878 -2472 912
rect -2365 878 -2331 912
rect -2224 878 -2190 912
rect -2083 878 -2049 912
rect -1942 878 -1908 912
rect -1801 878 -1767 912
rect -1660 878 -1626 912
rect -1519 878 -1485 912
rect -1378 878 -1344 912
rect -1237 878 -1203 912
rect -1096 878 -1062 912
rect -955 878 -921 912
rect -814 878 -780 912
rect -673 878 -639 912
rect -532 878 -498 912
rect -392 878 -358 912
rect -252 878 -218 912
rect -112 878 -78 912
rect 28 878 62 912
rect 168 878 202 912
rect 308 878 342 912
rect 448 878 482 912
rect 588 878 622 912
rect 728 878 762 912
rect 868 878 902 912
rect 1008 878 1042 912
rect -2506 -778 -2472 -744
rect -2369 -778 -2335 -744
rect -2232 -778 -2198 -744
rect -2095 -778 -2061 -744
rect -1958 -778 -1924 -744
rect -1821 -778 -1787 -744
rect -1684 -778 -1650 -744
rect -1547 -778 -1513 -744
rect -1410 -778 -1376 -744
rect -1273 -778 -1239 -744
rect -1136 -778 -1102 -744
rect -999 -778 -965 -744
rect -862 -778 -828 -744
rect -725 -778 -691 -744
rect -588 -778 -554 -744
rect -451 -778 -417 -744
rect -314 -778 -280 -744
rect -177 -778 -143 -744
rect -40 -778 -6 -744
rect 96 -778 130 -744
rect 232 -778 266 -744
rect 368 -778 402 -744
rect 504 -778 538 -744
rect 640 -778 674 -744
rect 776 -778 810 -744
rect 912 -778 946 -744
rect 1555 -2353 1589 -2319
rect 1709 -2353 1743 -2319
<< nsubdiffcont >>
rect -2534 50 -2500 84
rect -2465 50 -2431 84
rect -2396 50 -2362 84
rect -2327 50 -2293 84
rect -2258 50 -2224 84
rect -2189 50 -2155 84
rect -2120 50 -2086 84
rect -2052 50 -2018 84
rect -1984 50 -1950 84
rect -1916 50 -1882 84
rect -1848 50 -1814 84
rect -1780 50 -1746 84
rect -1712 50 -1678 84
rect -1644 50 -1610 84
rect -1576 50 -1542 84
rect -1508 50 -1474 84
rect -1440 50 -1406 84
rect -1372 50 -1338 84
rect -1304 50 -1270 84
rect -1236 50 -1202 84
rect -1168 50 -1134 84
rect -1100 50 -1066 84
rect -1032 50 -998 84
rect -964 50 -930 84
rect -896 50 -862 84
rect -828 50 -794 84
rect -760 50 -726 84
rect -692 50 -658 84
rect -624 50 -590 84
rect -556 50 -522 84
rect -488 50 -454 84
rect -420 50 -386 84
rect -352 50 -318 84
rect -284 50 -250 84
rect -216 50 -182 84
rect -148 50 -114 84
rect -80 50 -46 84
rect -12 50 22 84
rect 56 50 90 84
rect 124 50 158 84
rect 192 50 226 84
rect 260 50 294 84
rect 328 50 362 84
rect 396 50 430 84
rect 464 50 498 84
rect 532 50 566 84
rect 600 50 634 84
rect 668 50 702 84
rect 736 50 770 84
rect 804 50 838 84
rect 872 50 906 84
rect 940 50 974 84
rect 1555 -3181 1589 -3147
rect 1632 -3181 1666 -3147
rect 1709 -3181 1743 -3147
<< mvpsubdiffcont >>
rect -2213 -1970 -2179 -1936
rect -2070 -1970 -2036 -1936
rect -1927 -1970 -1893 -1936
rect -1784 -1970 -1750 -1936
rect -1641 -1970 -1607 -1936
rect -1498 -1970 -1464 -1936
rect -1355 -1970 -1321 -1936
rect -1212 -1970 -1178 -1936
rect -1069 -1970 -1035 -1936
rect -926 -1970 -892 -1936
rect -783 -1970 -749 -1936
rect -640 -1970 -606 -1936
rect -497 -1970 -463 -1936
rect -354 -1970 -320 -1936
rect -212 -1970 -178 -1936
rect -70 -1970 -36 -1936
rect 72 -1970 106 -1936
rect 214 -1970 248 -1936
rect 356 -1970 390 -1936
rect 498 -1970 532 -1936
<< mvnsubdiffcont >>
rect -1998 -969 -1964 -935
rect -1928 -969 -1894 -935
rect -1858 -969 -1824 -935
rect -1788 -969 -1754 -935
rect -1719 -969 -1685 -935
rect -1650 -969 -1616 -935
rect -1581 -969 -1547 -935
rect -1512 -969 -1478 -935
rect -1443 -969 -1409 -935
rect -1374 -969 -1340 -935
rect -1305 -969 -1271 -935
rect -1236 -969 -1202 -935
rect -1167 -969 -1133 -935
rect -1098 -969 -1064 -935
rect -1029 -969 -995 -935
rect -960 -969 -926 -935
rect -891 -969 -857 -935
rect -822 -969 -788 -935
rect -753 -969 -719 -935
rect -684 -969 -650 -935
rect -615 -969 -581 -935
rect -546 -969 -512 -935
rect -477 -969 -443 -935
rect -408 -969 -374 -935
rect -339 -969 -305 -935
rect -270 -969 -236 -935
rect -201 -969 -167 -935
rect -132 -969 -98 -935
rect -63 -969 -29 -935
rect 6 -969 40 -935
rect 75 -969 109 -935
rect 144 -969 178 -935
rect 213 -969 247 -935
rect 282 -969 316 -935
rect 351 -969 385 -935
rect 420 -969 454 -935
rect 489 -969 523 -935
<< poly >>
rect -1309 745 -1279 771
rect -1223 745 -1193 771
rect -1137 745 -1107 771
rect -1059 745 -1029 771
rect -913 745 -883 771
rect -1309 555 -1279 577
rect -1223 555 -1193 577
rect -1137 555 -1107 577
rect -1379 539 -1279 555
rect -1379 505 -1363 539
rect -1329 505 -1279 539
rect -1379 489 -1279 505
rect -1237 539 -1103 555
rect -1237 505 -1221 539
rect -1187 505 -1153 539
rect -1119 505 -1103 539
rect -1237 489 -1103 505
rect -1059 545 -1029 577
rect -913 555 -883 577
rect -1059 529 -965 545
rect -1059 495 -1015 529
rect -981 495 -965 529
rect -913 539 -757 555
rect -913 525 -807 539
rect -1309 447 -1279 489
rect -1231 447 -1201 489
rect -1141 447 -1111 489
rect -1059 479 -965 495
rect -842 505 -807 525
rect -773 505 -757 539
rect -842 489 -757 505
rect -1055 447 -1025 479
rect -842 447 -812 489
rect -1309 169 -1279 195
rect -1231 169 -1201 195
rect -1141 169 -1111 195
rect -1055 169 -1025 195
rect -842 169 -812 195
rect -2109 -1043 -1989 -1017
rect -1933 -1043 -1813 -1017
rect -1757 -1043 -1637 -1017
rect -1581 -1043 -1461 -1017
rect -1206 -1043 -1086 -1017
rect -1030 -1043 -910 -1017
rect -741 -1043 -621 -1017
rect -565 -1043 -445 -1017
rect -273 -1043 -153 -1017
rect -97 -1043 23 -1017
rect 198 -1043 318 -1017
rect 374 -1043 494 -1017
rect -2109 -1311 -1989 -1243
rect -1933 -1311 -1813 -1243
rect -1757 -1311 -1637 -1243
rect -1581 -1311 -1461 -1243
rect -1206 -1311 -1086 -1243
rect -1030 -1311 -910 -1243
rect -741 -1311 -621 -1243
rect -565 -1311 -445 -1243
rect -273 -1311 -153 -1243
rect -97 -1311 23 -1243
rect 198 -1311 318 -1243
rect 374 -1311 494 -1243
rect -2109 -1559 -1989 -1511
rect -2109 -1593 -2064 -1559
rect -2030 -1593 -1989 -1559
rect -2109 -1627 -1989 -1593
rect -2109 -1661 -2064 -1627
rect -2030 -1661 -1989 -1627
rect -2109 -1709 -1989 -1661
rect -1933 -1559 -1813 -1511
rect -1933 -1593 -1893 -1559
rect -1859 -1593 -1813 -1559
rect -1933 -1627 -1813 -1593
rect -1933 -1661 -1893 -1627
rect -1859 -1661 -1813 -1627
rect -1933 -1709 -1813 -1661
rect -1757 -1559 -1637 -1511
rect -1757 -1593 -1711 -1559
rect -1677 -1593 -1637 -1559
rect -1757 -1627 -1637 -1593
rect -1757 -1661 -1711 -1627
rect -1677 -1661 -1637 -1627
rect -1757 -1709 -1637 -1661
rect -1581 -1559 -1461 -1511
rect -1581 -1593 -1540 -1559
rect -1506 -1593 -1461 -1559
rect -1581 -1627 -1461 -1593
rect -1581 -1661 -1540 -1627
rect -1506 -1661 -1461 -1627
rect -1581 -1709 -1461 -1661
rect -1206 -1559 -1086 -1511
rect -1206 -1593 -1161 -1559
rect -1127 -1593 -1086 -1559
rect -1206 -1627 -1086 -1593
rect -1206 -1661 -1161 -1627
rect -1127 -1661 -1086 -1627
rect -1206 -1709 -1086 -1661
rect -1030 -1559 -910 -1511
rect -1030 -1593 -990 -1559
rect -956 -1593 -910 -1559
rect -1030 -1627 -910 -1593
rect -1030 -1661 -990 -1627
rect -956 -1661 -910 -1627
rect -1030 -1709 -910 -1661
rect -741 -1559 -621 -1511
rect -741 -1593 -696 -1559
rect -662 -1593 -621 -1559
rect -741 -1627 -621 -1593
rect -741 -1661 -696 -1627
rect -662 -1661 -621 -1627
rect -741 -1709 -621 -1661
rect -565 -1559 -445 -1511
rect -565 -1593 -525 -1559
rect -491 -1593 -445 -1559
rect -565 -1627 -445 -1593
rect -565 -1661 -525 -1627
rect -491 -1661 -445 -1627
rect -565 -1709 -445 -1661
rect -273 -1559 -153 -1511
rect -273 -1593 -230 -1559
rect -196 -1593 -153 -1559
rect -273 -1627 -153 -1593
rect -273 -1661 -230 -1627
rect -196 -1661 -153 -1627
rect -273 -1709 -153 -1661
rect -97 -1559 23 -1511
rect -97 -1593 -52 -1559
rect -18 -1593 23 -1559
rect -97 -1627 23 -1593
rect -97 -1661 -52 -1627
rect -18 -1661 23 -1627
rect -97 -1709 23 -1661
rect 198 -1559 318 -1511
rect 198 -1593 239 -1559
rect 273 -1593 318 -1559
rect 198 -1627 318 -1593
rect 198 -1661 239 -1627
rect 273 -1661 318 -1627
rect 198 -1709 318 -1661
rect 374 -1559 494 -1511
rect 374 -1593 417 -1559
rect 451 -1593 494 -1559
rect 374 -1627 494 -1593
rect 374 -1661 417 -1627
rect 451 -1661 494 -1627
rect 374 -1709 494 -1661
rect -2109 -1875 -1989 -1849
rect -1933 -1875 -1813 -1849
rect -1757 -1875 -1637 -1849
rect -1581 -1875 -1461 -1849
rect -1206 -1875 -1086 -1849
rect -1030 -1875 -910 -1849
rect -741 -1875 -621 -1849
rect -565 -1875 -445 -1849
rect -273 -1875 -153 -1849
rect -97 -1875 23 -1849
rect 198 -1875 318 -1849
rect 374 -1875 494 -1849
<< polycont >>
rect -1363 505 -1329 539
rect -1221 505 -1187 539
rect -1153 505 -1119 539
rect -1015 495 -981 529
rect -807 505 -773 539
rect -2064 -1593 -2030 -1559
rect -2064 -1661 -2030 -1627
rect -1893 -1593 -1859 -1559
rect -1893 -1661 -1859 -1627
rect -1711 -1593 -1677 -1559
rect -1711 -1661 -1677 -1627
rect -1540 -1593 -1506 -1559
rect -1540 -1661 -1506 -1627
rect -1161 -1593 -1127 -1559
rect -1161 -1661 -1127 -1627
rect -990 -1593 -956 -1559
rect -990 -1661 -956 -1627
rect -696 -1593 -662 -1559
rect -696 -1661 -662 -1627
rect -525 -1593 -491 -1559
rect -525 -1661 -491 -1627
rect -230 -1593 -196 -1559
rect -230 -1661 -196 -1627
rect -52 -1593 -18 -1559
rect -52 -1661 -18 -1627
rect 239 -1593 273 -1559
rect 239 -1661 273 -1627
rect 417 -1593 451 -1559
rect 417 -1661 451 -1627
<< locali >>
rect -2530 879 -2506 912
rect -2556 878 -2506 879
rect -2472 878 -2365 912
rect -2331 878 -2224 912
rect -2190 878 -2083 912
rect -2049 878 -1942 912
rect -1908 878 -1801 912
rect -1767 878 -1660 912
rect -1626 878 -1519 912
rect -1485 878 -1378 912
rect -1344 878 -1237 912
rect -1203 878 -1096 912
rect -1062 878 -955 912
rect -921 878 -814 912
rect -780 878 -673 912
rect -639 878 -532 912
rect -498 878 -392 912
rect -358 878 -252 912
rect -218 878 -112 912
rect -78 878 28 912
rect 62 878 168 912
rect 202 878 308 912
rect 342 878 448 912
rect 482 878 588 912
rect 622 878 728 912
rect 762 878 868 912
rect 902 878 1008 912
rect 1042 879 1066 912
rect 1042 878 1092 879
rect -2556 831 1092 878
rect -1404 797 -1373 831
rect -1339 797 -1277 831
rect -1243 797 -1181 831
rect -1147 797 -1085 831
rect -1051 797 -989 831
rect -955 797 -893 831
rect -859 797 -797 831
rect -763 797 -732 831
rect 420 797 516 831
rect -2062 651 -2028 689
rect -1724 612 -1629 744
rect -1667 595 -1629 612
rect -1370 733 -1318 797
rect -1370 699 -1354 733
rect -1320 699 -1318 733
rect -1370 656 -1318 699
rect -1370 622 -1354 656
rect -1320 622 -1318 656
rect -1370 606 -1318 622
rect -1284 731 -1232 747
rect -1284 697 -1268 731
rect -1234 697 -1232 731
rect -1284 640 -1232 697
rect -1198 716 -1132 797
rect -1198 682 -1182 716
rect -1148 682 -1132 716
rect -1198 674 -1132 682
rect -1064 729 -845 763
rect -1064 640 -1030 729
rect -1284 606 -1268 640
rect -1234 606 -1030 640
rect -996 661 -980 695
rect -946 661 -913 695
rect -996 619 -913 661
rect -996 585 -980 619
rect -946 585 -913 619
rect -996 581 -913 585
rect -2487 466 -2449 500
rect -2293 458 -2243 554
rect -2196 511 -2153 545
rect -1728 538 -1722 572
rect -1959 484 -1942 504
rect -1908 504 -1902 518
rect -1621 515 -1583 549
rect -1387 539 -1313 572
rect -1387 505 -1363 539
rect -1329 505 -1313 539
rect -1908 484 -1893 504
rect -1489 410 -1455 448
rect -1387 469 -1313 505
rect -1279 539 -1051 572
rect -947 558 -913 581
rect -1279 537 -1221 539
rect -1187 537 -1153 539
rect -1279 503 -1226 537
rect -1187 505 -1154 537
rect -1119 505 -1051 539
rect -1192 503 -1154 505
rect -1120 503 -1051 505
rect -1017 529 -981 545
rect -1017 495 -1015 529
rect -1017 469 -981 495
rect -1353 435 -1313 469
rect -1279 435 -981 469
rect -879 568 -845 729
rect -811 733 -761 797
rect -777 699 -761 733
rect -811 652 -761 699
rect -495 694 -457 728
rect 1430 723 1464 761
rect -777 618 -761 652
rect -811 602 -761 618
rect 1584 723 1618 761
rect 1736 723 1770 761
rect 2678 723 2712 761
rect 2824 723 2858 761
rect 2978 700 3012 738
rect -230 642 -196 685
rect -113 576 -79 614
rect -879 539 -757 568
rect -879 534 -807 539
rect -947 500 -913 524
rect -823 505 -807 534
rect -773 505 -757 539
rect -662 523 -657 557
rect -475 523 -466 557
rect -363 514 -320 548
rect -947 483 -857 500
rect -823 489 -757 505
rect -913 455 -857 483
rect -913 439 -837 455
rect -913 405 -887 439
rect -853 405 -837 439
rect -913 401 -837 405
rect -1853 332 -1819 370
rect -1370 367 -1354 401
rect -1320 367 -982 401
rect -791 367 -757 489
rect 60 489 94 528
rect 175 550 209 562
rect 259 489 293 528
rect 352 542 386 552
rect 560 480 594 518
rect 779 458 836 554
rect 985 481 1023 515
rect -1370 323 -1304 367
rect -1016 333 -757 367
rect -1370 289 -1354 323
rect -1320 289 -1304 323
rect -1370 249 -1304 289
rect -1370 215 -1354 249
rect -1320 215 -1304 249
rect -1370 199 -1304 215
rect -1206 317 -1150 333
rect -1206 283 -1190 317
rect -1156 283 -1150 317
rect -1206 241 -1150 283
rect -1206 207 -1190 241
rect -1156 207 -1150 241
rect -1206 165 -1150 207
rect -1116 299 -1100 333
rect -1066 299 -1050 333
rect -1116 279 -751 299
rect -1116 265 -801 279
rect -1116 241 -1050 265
rect -1116 207 -1100 241
rect -1066 207 -1050 241
rect -817 245 -801 265
rect -767 245 -751 279
rect -1116 199 -1050 207
rect -1011 227 -945 231
rect -817 229 -751 245
rect 811 233 849 267
rect -1011 193 -995 227
rect -961 193 -945 227
rect -1011 165 -945 193
rect -1404 131 -1373 165
rect -1339 131 -1277 165
rect -1243 131 -1181 165
rect -1147 131 -1085 165
rect -1051 131 -989 165
rect -955 131 -893 165
rect -859 131 -797 165
rect -763 131 -732 165
rect 420 131 516 165
rect -2510 84 -2471 90
rect -2437 84 -2398 90
rect -2364 84 -2325 90
rect -2291 84 -2252 90
rect -2218 84 -2179 90
rect -2145 84 -2106 90
rect -2072 84 -2033 90
rect -1999 84 -1960 90
rect -1926 84 -1887 90
rect -1853 84 -1814 90
rect -2558 56 -2544 84
rect -2500 56 -2471 84
rect -2431 56 -2398 84
rect -2558 50 -2534 56
rect -2500 50 -2465 56
rect -2431 50 -2396 56
rect -2362 50 -2327 84
rect -2291 56 -2258 84
rect -2218 56 -2189 84
rect -2145 56 -2120 84
rect -2072 56 -2052 84
rect -1999 56 -1984 84
rect -1926 56 -1916 84
rect -1853 56 -1848 84
rect -2293 50 -2258 56
rect -2224 50 -2189 56
rect -2155 50 -2120 56
rect -2086 50 -2052 56
rect -2018 50 -1984 56
rect -1950 50 -1916 56
rect -1882 50 -1848 56
rect -1780 84 -1741 90
rect -1707 84 -1668 90
rect -1634 84 -1595 90
rect -1561 84 -1522 90
rect -1488 84 -1449 90
rect -1415 84 -1376 90
rect -1342 84 -1303 90
rect -1269 84 -1230 90
rect -1196 84 -1157 90
rect -1123 84 -1084 90
rect -1050 84 -1011 90
rect -977 84 -938 90
rect -904 84 -865 90
rect -831 84 -792 90
rect -758 84 -719 90
rect -685 84 -646 90
rect -612 84 -573 90
rect -539 84 -500 90
rect -466 84 -427 90
rect -393 84 -354 90
rect -320 84 -281 90
rect -247 84 -208 90
rect -174 84 -135 90
rect -101 84 -62 90
rect -28 84 11 90
rect 45 84 84 90
rect 118 84 157 90
rect 191 84 230 90
rect 264 84 303 90
rect 337 84 376 90
rect 410 84 448 90
rect 482 84 520 90
rect 554 84 592 90
rect 626 84 664 90
rect 698 84 736 90
rect 770 84 808 90
rect 842 84 880 90
rect 914 84 952 90
rect -1814 50 -1780 56
rect -1746 56 -1741 84
rect -1678 56 -1668 84
rect -1610 56 -1595 84
rect -1542 56 -1522 84
rect -1474 56 -1449 84
rect -1406 56 -1376 84
rect -1746 50 -1712 56
rect -1678 50 -1644 56
rect -1610 50 -1576 56
rect -1542 50 -1508 56
rect -1474 50 -1440 56
rect -1406 50 -1372 56
rect -1338 50 -1304 84
rect -1269 56 -1236 84
rect -1196 56 -1168 84
rect -1123 56 -1100 84
rect -1050 56 -1032 84
rect -977 56 -964 84
rect -904 56 -896 84
rect -831 56 -828 84
rect -1270 50 -1236 56
rect -1202 50 -1168 56
rect -1134 50 -1100 56
rect -1066 50 -1032 56
rect -998 50 -964 56
rect -930 50 -896 56
rect -862 50 -828 56
rect -794 56 -792 84
rect -726 56 -719 84
rect -658 56 -646 84
rect -590 56 -573 84
rect -522 56 -500 84
rect -454 56 -427 84
rect -386 56 -354 84
rect -794 50 -760 56
rect -726 50 -692 56
rect -658 50 -624 56
rect -590 50 -556 56
rect -522 50 -488 56
rect -454 50 -420 56
rect -386 50 -352 56
rect -318 50 -284 84
rect -247 56 -216 84
rect -174 56 -148 84
rect -101 56 -80 84
rect -28 56 -12 84
rect 45 56 56 84
rect 118 56 124 84
rect 191 56 192 84
rect -250 50 -216 56
rect -182 50 -148 56
rect -114 50 -80 56
rect -46 50 -12 56
rect 22 50 56 56
rect 90 50 124 56
rect 158 50 192 56
rect 226 56 230 84
rect 294 56 303 84
rect 362 56 376 84
rect 430 56 448 84
rect 498 56 520 84
rect 566 56 592 84
rect 634 56 664 84
rect 226 50 260 56
rect 294 50 328 56
rect 362 50 396 56
rect 430 50 464 56
rect 498 50 532 56
rect 566 50 600 56
rect 634 50 668 56
rect 702 50 736 84
rect 770 50 804 84
rect 842 56 872 84
rect 914 56 940 84
rect 986 56 998 84
rect 838 50 872 56
rect 906 50 940 56
rect 974 50 998 56
rect 36 -31 132 3
rect -2293 -290 -2205 -84
rect -2048 -239 -2014 -201
rect -853 -256 -765 -84
rect -2338 -346 -2304 -333
rect -2525 -374 -2491 -361
rect -2258 -335 -2205 -290
rect -2258 -369 -2232 -335
rect -2198 -369 -2160 -335
rect -1851 -346 -1817 -306
rect -850 -290 -811 -256
rect -777 -290 -765 -256
rect -277 -290 -189 -84
rect 169 -175 203 -137
rect -2258 -420 -2205 -369
rect -1767 -346 -1733 -333
rect -1617 -369 -1579 -335
rect -1469 -346 -1435 -308
rect -1331 -369 -1293 -335
rect -1141 -380 -1091 -324
rect -1913 -414 -1900 -380
rect -1129 -414 -1091 -380
rect -912 -381 -891 -347
rect -753 -369 -715 -335
rect -618 -348 -592 -314
rect -321 -357 -287 -326
rect -472 -414 -459 -380
rect -242 -360 -189 -290
rect 452 -175 486 -137
rect -33 -280 1 -242
rect -242 -394 -223 -360
rect -189 -394 -151 -360
rect -1141 -420 -1091 -414
rect -242 -420 -189 -394
rect 389 -420 451 -324
rect 834 -344 868 -306
rect 597 -385 635 -351
rect 729 -384 744 -350
rect 778 -384 795 -350
rect 1033 -344 1067 -306
rect 909 -378 1033 -350
rect 729 -444 795 -384
rect 909 -444 1067 -378
rect 36 -697 132 -663
rect -2484 -744 -2445 -735
rect -2530 -769 -2518 -744
rect -2472 -769 -2445 -744
rect -2411 -769 -2372 -735
rect -2338 -744 -2299 -735
rect -2335 -769 -2299 -744
rect -2265 -744 -2226 -735
rect -2265 -769 -2232 -744
rect -2192 -769 -2153 -735
rect -2119 -744 -2080 -735
rect -2119 -769 -2095 -744
rect -2046 -769 -2007 -735
rect -1973 -744 -1934 -735
rect -1973 -769 -1958 -744
rect -1900 -769 -1861 -735
rect -1827 -744 -1788 -735
rect -1827 -769 -1821 -744
rect -1754 -769 -1715 -735
rect -1681 -744 -1642 -735
rect -1650 -769 -1642 -744
rect -1608 -769 -1570 -735
rect -1536 -744 -1498 -735
rect -1513 -769 -1498 -744
rect -1464 -769 -1426 -735
rect -1392 -744 -1354 -735
rect -1376 -769 -1354 -744
rect -1320 -769 -1282 -735
rect -1248 -744 -1210 -735
rect -1239 -769 -1210 -744
rect -1176 -769 -1138 -735
rect -1104 -744 -1066 -735
rect -1102 -769 -1066 -744
rect -1032 -744 -994 -735
rect -1032 -769 -999 -744
rect -960 -769 -922 -735
rect -888 -744 -850 -735
rect -888 -769 -862 -744
rect -816 -769 -778 -735
rect -744 -744 -706 -735
rect -744 -769 -725 -744
rect -672 -769 -634 -735
rect -600 -744 -562 -735
rect -600 -769 -588 -744
rect -528 -769 -490 -735
rect -456 -744 -418 -735
rect -456 -769 -451 -744
rect -384 -769 -346 -735
rect -312 -744 -274 -735
rect -280 -769 -274 -744
rect -240 -769 -202 -735
rect -168 -744 -130 -735
rect -143 -769 -130 -744
rect -96 -769 -58 -735
rect -24 -744 14 -735
rect -6 -769 14 -744
rect 48 -769 86 -735
rect 120 -744 158 -735
rect 130 -769 158 -744
rect 192 -769 230 -735
rect 264 -744 302 -735
rect 266 -769 302 -744
rect 336 -744 374 -735
rect 336 -769 368 -744
rect 408 -769 446 -735
rect 480 -744 518 -735
rect 480 -769 504 -744
rect 552 -769 590 -735
rect 624 -744 662 -735
rect 624 -769 640 -744
rect 696 -769 734 -735
rect 768 -744 806 -735
rect 768 -769 776 -744
rect 840 -769 878 -735
rect 912 -744 950 -735
rect -2530 -778 -2506 -769
rect -2472 -778 -2369 -769
rect -2335 -778 -2232 -769
rect -2198 -778 -2095 -769
rect -2061 -778 -1958 -769
rect -1924 -778 -1821 -769
rect -1787 -778 -1684 -769
rect -1650 -778 -1547 -769
rect -1513 -778 -1410 -769
rect -1376 -778 -1273 -769
rect -1239 -778 -1136 -769
rect -1102 -778 -999 -769
rect -965 -778 -862 -769
rect -828 -778 -725 -769
rect -691 -778 -588 -769
rect -554 -778 -451 -769
rect -417 -778 -314 -769
rect -280 -778 -177 -769
rect -143 -778 -40 -769
rect -6 -778 96 -769
rect 130 -778 232 -769
rect 266 -778 368 -769
rect 402 -778 504 -769
rect 538 -778 640 -769
rect 674 -778 776 -769
rect 810 -778 912 -769
rect 946 -769 950 -744
rect 946 -778 970 -769
rect -2205 -969 -2165 -935
rect -2131 -969 -2091 -935
rect -2057 -969 -2017 -935
rect -1964 -969 -1943 -935
rect -1894 -969 -1869 -935
rect -1824 -969 -1795 -935
rect -1754 -969 -1721 -935
rect -1685 -969 -1650 -935
rect -1613 -969 -1581 -935
rect -1540 -969 -1512 -935
rect -1467 -969 -1443 -935
rect -1394 -969 -1374 -935
rect -1321 -969 -1305 -935
rect -1248 -969 -1236 -935
rect -1175 -969 -1167 -935
rect -1102 -969 -1098 -935
rect -1064 -969 -1063 -935
rect -995 -969 -990 -935
rect -926 -969 -917 -935
rect -857 -969 -844 -935
rect -788 -969 -771 -935
rect -719 -969 -698 -935
rect -650 -969 -625 -935
rect -581 -969 -552 -935
rect -512 -969 -479 -935
rect -443 -969 -408 -935
rect -372 -969 -339 -935
rect -299 -969 -270 -935
rect -226 -969 -201 -935
rect -153 -969 -132 -935
rect -80 -969 -63 -935
rect -7 -969 6 -935
rect 66 -969 75 -935
rect 139 -969 144 -935
rect 212 -969 213 -935
rect 247 -969 282 -935
rect 316 -969 351 -935
rect 385 -969 420 -935
rect 454 -969 489 -935
rect 523 -969 547 -935
rect -2154 -1061 -2120 -1049
rect -2154 -1129 -2120 -1121
rect -2154 -1197 -2120 -1163
rect -2154 -1323 -2120 -1231
rect -1978 -1061 -1944 -1043
rect -1978 -1129 -1944 -1095
rect -1978 -1197 -1944 -1163
rect -1978 -1323 -1944 -1231
rect -1802 -1061 -1768 -1049
rect -1802 -1129 -1768 -1121
rect -1802 -1197 -1768 -1163
rect -1802 -1323 -1768 -1231
rect -2154 -1391 -2120 -1357
rect -1944 -1357 -1936 -1337
rect -1974 -1371 -1936 -1357
rect -2154 -1459 -2120 -1425
rect -2154 -1509 -2120 -1493
rect -1978 -1391 -1944 -1371
rect -1978 -1459 -1944 -1425
rect -2080 -1577 -2070 -1559
rect -2080 -1593 -2064 -1577
rect -2030 -1593 -2014 -1559
rect -2080 -1615 -2014 -1593
rect -2080 -1649 -2070 -1615
rect -2036 -1627 -2014 -1615
rect -2080 -1661 -2064 -1649
rect -2030 -1661 -2014 -1627
rect -2154 -1721 -2120 -1705
rect -1978 -1732 -1944 -1493
rect -1802 -1391 -1768 -1357
rect -1802 -1459 -1768 -1425
rect -1802 -1509 -1768 -1493
rect -1626 -1061 -1592 -1043
rect -1626 -1129 -1592 -1095
rect -1626 -1197 -1592 -1163
rect -1450 -1061 -1416 -1049
rect -1450 -1129 -1416 -1121
rect -1626 -1323 -1592 -1231
rect -1626 -1391 -1592 -1357
rect -1626 -1459 -1592 -1425
rect -1909 -1593 -1893 -1559
rect -1859 -1573 -1855 -1559
rect -1626 -1543 -1592 -1493
rect -1859 -1593 -1821 -1573
rect -1909 -1611 -1821 -1593
rect -1909 -1627 -1855 -1611
rect -1909 -1661 -1893 -1627
rect -1859 -1645 -1855 -1627
rect -1727 -1577 -1725 -1559
rect -1727 -1593 -1711 -1577
rect -1677 -1593 -1661 -1559
rect -1727 -1615 -1661 -1593
rect -1859 -1661 -1843 -1645
rect -1727 -1649 -1725 -1615
rect -1691 -1627 -1661 -1615
rect -1727 -1661 -1711 -1649
rect -1677 -1661 -1661 -1627
rect -1626 -1615 -1592 -1577
rect -2120 -1755 -1944 -1732
rect -2154 -1766 -1944 -1755
rect -1802 -1721 -1768 -1705
rect -1802 -1766 -1768 -1755
rect -1626 -1732 -1592 -1649
rect -1556 -1182 -1490 -1169
rect -1556 -1216 -1539 -1182
rect -1505 -1216 -1490 -1182
rect -1556 -1254 -1490 -1216
rect -1556 -1288 -1539 -1254
rect -1505 -1288 -1490 -1254
rect -1556 -1559 -1490 -1288
rect -1450 -1197 -1416 -1163
rect -1450 -1323 -1416 -1231
rect -1450 -1391 -1416 -1357
rect -1450 -1459 -1416 -1425
rect -1450 -1509 -1416 -1493
rect -1251 -1061 -1217 -1049
rect -1251 -1129 -1217 -1121
rect -1251 -1197 -1217 -1163
rect -1251 -1323 -1217 -1231
rect -1075 -1061 -1041 -1043
rect -1075 -1129 -1041 -1095
rect -1075 -1197 -1041 -1163
rect -1251 -1391 -1217 -1357
rect -1251 -1459 -1217 -1425
rect -1251 -1509 -1217 -1493
rect -1178 -1319 -1111 -1312
rect -1178 -1353 -1159 -1319
rect -1125 -1353 -1111 -1319
rect -1178 -1391 -1111 -1353
rect -1178 -1425 -1159 -1391
rect -1125 -1425 -1111 -1391
rect -1556 -1593 -1540 -1559
rect -1506 -1593 -1490 -1559
rect -1556 -1627 -1490 -1593
rect -1556 -1661 -1540 -1627
rect -1506 -1661 -1490 -1627
rect -1178 -1559 -1111 -1425
rect -1178 -1593 -1161 -1559
rect -1127 -1593 -1111 -1559
rect -1178 -1627 -1111 -1593
rect -1178 -1661 -1161 -1627
rect -1127 -1661 -1111 -1627
rect -1075 -1323 -1041 -1231
rect -899 -1061 -865 -1049
rect -899 -1129 -865 -1121
rect -899 -1197 -865 -1163
rect -1075 -1391 -1041 -1357
rect -1075 -1459 -1041 -1425
rect -1450 -1721 -1416 -1705
rect -1289 -1720 -1251 -1686
rect -1626 -1755 -1450 -1732
rect -1626 -1766 -1416 -1755
rect -2154 -1789 -2115 -1766
rect -2120 -1823 -2115 -1789
rect -2154 -1839 -2115 -1823
rect -1802 -1838 -1768 -1823
rect -1455 -1789 -1416 -1766
rect -1455 -1823 -1450 -1789
rect -1455 -1839 -1416 -1823
rect -1251 -1721 -1217 -1720
rect -1075 -1732 -1041 -1493
rect -1006 -1260 -940 -1247
rect -1006 -1294 -993 -1260
rect -959 -1294 -940 -1260
rect -1006 -1332 -940 -1294
rect -1006 -1366 -993 -1332
rect -959 -1366 -940 -1332
rect -1006 -1559 -940 -1366
rect -899 -1323 -865 -1231
rect -899 -1391 -865 -1357
rect -899 -1459 -865 -1425
rect -899 -1509 -865 -1493
rect -786 -1061 -752 -1049
rect -786 -1129 -752 -1121
rect -786 -1197 -752 -1163
rect -786 -1323 -752 -1231
rect -610 -1061 -576 -1043
rect -610 -1129 -576 -1095
rect -610 -1197 -576 -1163
rect -610 -1323 -576 -1231
rect -786 -1391 -752 -1357
rect -786 -1459 -752 -1425
rect -786 -1509 -752 -1493
rect -712 -1368 -695 -1334
rect -661 -1368 -646 -1334
rect -712 -1406 -646 -1368
rect -712 -1440 -695 -1406
rect -661 -1440 -646 -1406
rect -1006 -1593 -990 -1559
rect -956 -1593 -940 -1559
rect -1006 -1627 -940 -1593
rect -1006 -1661 -990 -1627
rect -956 -1661 -940 -1627
rect -847 -1577 -809 -1543
rect -775 -1577 -752 -1543
rect -881 -1631 -752 -1577
rect -1217 -1755 -1041 -1732
rect -1251 -1766 -1041 -1755
rect -899 -1721 -865 -1705
rect -899 -1766 -865 -1755
rect -1251 -1789 -1212 -1766
rect -1217 -1823 -1212 -1789
rect -1251 -1839 -1212 -1823
rect -899 -1838 -865 -1823
rect -786 -1721 -752 -1631
rect -712 -1559 -646 -1440
rect -712 -1593 -696 -1559
rect -662 -1593 -646 -1559
rect -712 -1627 -646 -1593
rect -712 -1661 -696 -1627
rect -662 -1661 -646 -1627
rect -434 -1061 -400 -1049
rect -434 -1129 -400 -1121
rect -434 -1197 -400 -1163
rect -434 -1323 -400 -1231
rect -610 -1391 -576 -1357
rect -610 -1459 -576 -1425
rect -610 -1732 -576 -1493
rect -541 -1368 -519 -1334
rect -485 -1368 -475 -1334
rect -541 -1406 -475 -1368
rect -541 -1440 -519 -1406
rect -485 -1440 -475 -1406
rect -541 -1559 -475 -1440
rect -434 -1391 -400 -1357
rect -434 -1459 -400 -1425
rect -434 -1509 -400 -1493
rect -318 -1061 -284 -1049
rect -318 -1129 -284 -1121
rect -318 -1197 -284 -1163
rect -318 -1323 -284 -1231
rect -318 -1391 -284 -1357
rect -318 -1459 -284 -1425
rect -142 -1061 -108 -1045
rect -142 -1129 -108 -1095
rect -142 -1197 -108 -1163
rect -142 -1323 -108 -1231
rect -142 -1391 -108 -1357
rect -142 -1441 -108 -1425
rect 34 -1061 68 -1015
rect 34 -1129 68 -1095
rect 34 -1197 68 -1163
rect 153 -1061 187 -1015
rect 153 -1129 187 -1095
rect 153 -1176 187 -1163
rect 329 -1061 363 -1045
rect 329 -1129 363 -1095
rect 155 -1197 193 -1176
rect 187 -1210 193 -1197
rect 329 -1197 363 -1163
rect 505 -1061 539 -1049
rect 505 -1129 539 -1121
rect 34 -1323 68 -1231
rect 34 -1391 68 -1357
rect 34 -1459 68 -1425
rect -142 -1476 34 -1475
rect -318 -1509 -284 -1493
rect -176 -1510 -138 -1476
rect -104 -1493 34 -1476
rect -104 -1509 68 -1493
rect 153 -1323 187 -1231
rect 153 -1391 187 -1357
rect 153 -1459 187 -1425
rect 329 -1323 363 -1231
rect 329 -1391 363 -1357
rect 329 -1441 363 -1425
rect 401 -1210 415 -1176
rect 449 -1210 467 -1176
rect 401 -1248 467 -1210
rect 401 -1282 415 -1248
rect 449 -1282 467 -1248
rect 187 -1493 363 -1475
rect 153 -1509 363 -1493
rect -541 -1593 -525 -1559
rect -491 -1593 -475 -1559
rect -541 -1627 -475 -1593
rect -541 -1661 -525 -1627
rect -491 -1661 -475 -1627
rect -286 -1593 -230 -1559
rect -196 -1593 -180 -1559
rect -286 -1610 -180 -1593
rect -252 -1627 -214 -1610
rect -252 -1644 -230 -1627
rect -286 -1661 -230 -1644
rect -196 -1661 -180 -1644
rect -752 -1755 -576 -1732
rect -786 -1766 -576 -1755
rect -434 -1721 -400 -1705
rect -434 -1766 -400 -1755
rect -786 -1789 -747 -1766
rect -752 -1823 -747 -1789
rect -786 -1839 -747 -1823
rect -434 -1838 -400 -1823
rect -318 -1721 -284 -1705
rect -318 -1766 -284 -1755
rect -318 -1838 -284 -1823
rect -142 -1721 -108 -1510
rect -68 -1593 -52 -1559
rect -18 -1593 -2 -1559
rect -68 -1610 -2 -1593
rect 223 -1593 239 -1559
rect 273 -1593 289 -1559
rect -68 -1644 -67 -1610
rect -33 -1627 5 -1610
rect -18 -1644 5 -1627
rect 223 -1613 289 -1593
rect -68 -1661 -52 -1644
rect -18 -1661 -2 -1644
rect 217 -1627 255 -1613
rect 217 -1647 239 -1627
rect 223 -1661 239 -1647
rect 273 -1661 289 -1647
rect -142 -1789 -108 -1755
rect -142 -1839 -108 -1823
rect 34 -1721 68 -1705
rect 34 -1766 68 -1755
rect 34 -1838 68 -1823
rect 153 -1721 187 -1705
rect 153 -1766 187 -1755
rect 153 -1838 187 -1823
rect 329 -1721 363 -1509
rect 401 -1559 467 -1282
rect 505 -1197 539 -1163
rect 4702 -1164 4846 -1151
rect 1324 -1200 1362 -1166
rect 4736 -1198 4774 -1164
rect 4808 -1198 4846 -1164
rect 4702 -1205 4846 -1198
rect 505 -1323 539 -1231
rect 4639 -1320 4846 -1307
rect 1324 -1355 1362 -1321
rect 4673 -1354 4711 -1320
rect 4745 -1354 4846 -1320
rect 505 -1391 539 -1357
rect 4639 -1361 4846 -1354
rect 505 -1459 539 -1425
rect 505 -1509 539 -1493
rect 1324 -1505 1362 -1471
rect 4556 -1473 4846 -1463
rect 4590 -1507 4628 -1473
rect 4662 -1507 4846 -1473
rect 4556 -1517 4846 -1507
rect 401 -1593 417 -1559
rect 451 -1593 467 -1559
rect 401 -1627 467 -1593
rect 401 -1661 417 -1627
rect 451 -1661 467 -1627
rect 1324 -1661 1362 -1627
rect 4561 -1630 4846 -1619
rect 4561 -1664 4562 -1630
rect 4596 -1664 4634 -1630
rect 4668 -1664 4846 -1630
rect 4561 -1673 4846 -1664
rect 329 -1789 363 -1755
rect 329 -1839 363 -1823
rect 505 -1721 539 -1705
rect 505 -1766 539 -1755
rect 505 -1838 539 -1823
rect -2237 -1970 -2213 -1936
rect -2151 -1970 -2111 -1936
rect -2077 -1970 -2070 -1936
rect -2003 -1970 -1963 -1936
rect -1929 -1970 -1927 -1936
rect -1893 -1970 -1889 -1936
rect -1855 -1970 -1815 -1936
rect -1750 -1970 -1741 -1936
rect -1707 -1970 -1667 -1936
rect -1607 -1970 -1593 -1936
rect -1559 -1970 -1519 -1936
rect -1464 -1970 -1445 -1936
rect -1411 -1970 -1372 -1936
rect -1321 -1970 -1299 -1936
rect -1265 -1970 -1226 -1936
rect -1178 -1970 -1153 -1936
rect -1119 -1970 -1080 -1936
rect -1035 -1970 -1007 -1936
rect -973 -1970 -934 -1936
rect -892 -1970 -861 -1936
rect -827 -1970 -788 -1936
rect -749 -1970 -715 -1936
rect -681 -1970 -642 -1936
rect -606 -1970 -569 -1936
rect -535 -1970 -497 -1936
rect -462 -1970 -423 -1936
rect -389 -1970 -354 -1936
rect -316 -1970 -277 -1936
rect -243 -1970 -212 -1936
rect -170 -1970 -131 -1936
rect -97 -1970 -70 -1936
rect -24 -1970 15 -1936
rect 49 -1970 72 -1936
rect 122 -1970 161 -1936
rect 195 -1970 214 -1936
rect 268 -1970 307 -1936
rect 341 -1970 356 -1936
rect 414 -1970 453 -1936
rect 487 -1970 498 -1936
rect 1505 -2353 1555 -2319
rect 1589 -2353 1709 -2319
rect 1743 -2353 1793 -2319
rect 1505 -2400 1793 -2353
rect 1715 -2619 1749 -2581
rect 1583 -2738 1621 -2704
rect 1505 -3147 1793 -3066
rect 1505 -3181 1555 -3147
rect 1589 -3181 1632 -3147
rect 1666 -3181 1709 -3147
rect 1743 -3181 1793 -3147
<< viali >>
rect -1373 797 -1339 831
rect -1277 797 -1243 831
rect -1181 797 -1147 831
rect -1085 797 -1051 831
rect -989 797 -955 831
rect -893 797 -859 831
rect -797 797 -763 831
rect -2062 689 -2028 723
rect -2062 617 -2028 651
rect -2521 466 -2487 500
rect -2449 466 -2415 500
rect -2230 511 -2196 545
rect -2153 511 -2119 545
rect -1762 538 -1728 572
rect -1942 484 -1908 518
rect -1655 515 -1621 549
rect -1583 515 -1549 549
rect -1489 448 -1455 482
rect -1226 505 -1221 537
rect -1221 505 -1192 537
rect -1154 505 -1153 537
rect -1153 505 -1120 537
rect -1226 503 -1192 505
rect -1154 503 -1120 505
rect -1387 435 -1353 469
rect -1313 435 -1279 469
rect -947 524 -913 558
rect 1430 761 1464 795
rect -529 694 -495 728
rect -457 694 -423 728
rect -230 685 -196 719
rect 1430 689 1464 723
rect 1584 761 1618 795
rect 1584 689 1618 723
rect 1736 761 1770 795
rect 1736 689 1770 723
rect 2678 761 2712 795
rect 2678 689 2712 723
rect 2824 761 2858 795
rect 2824 689 2858 723
rect 2978 738 3012 772
rect 2978 666 3012 700
rect -230 608 -196 642
rect -113 614 -79 648
rect -696 523 -662 557
rect -509 523 -475 557
rect -397 514 -363 548
rect -320 514 -286 548
rect -113 542 -79 576
rect 60 528 94 562
rect -947 449 -913 483
rect -1853 370 -1819 404
rect -1489 376 -1455 410
rect -1853 298 -1819 332
rect 175 516 209 550
rect 259 528 293 562
rect 60 455 94 489
rect 352 508 386 542
rect 560 518 594 552
rect 259 455 293 489
rect 560 446 594 480
rect 951 481 985 515
rect 1023 481 1057 515
rect 777 233 811 267
rect 849 233 883 267
rect -1373 131 -1339 165
rect -1277 131 -1243 165
rect -1181 131 -1147 165
rect -1085 131 -1051 165
rect -989 131 -955 165
rect -893 131 -859 165
rect -797 131 -763 165
rect -2544 84 -2510 90
rect -2471 84 -2437 90
rect -2398 84 -2364 90
rect -2325 84 -2291 90
rect -2252 84 -2218 90
rect -2179 84 -2145 90
rect -2106 84 -2072 90
rect -2033 84 -1999 90
rect -1960 84 -1926 90
rect -1887 84 -1853 90
rect -2544 56 -2534 84
rect -2534 56 -2510 84
rect -2471 56 -2465 84
rect -2465 56 -2437 84
rect -2398 56 -2396 84
rect -2396 56 -2364 84
rect -2325 56 -2293 84
rect -2293 56 -2291 84
rect -2252 56 -2224 84
rect -2224 56 -2218 84
rect -2179 56 -2155 84
rect -2155 56 -2145 84
rect -2106 56 -2086 84
rect -2086 56 -2072 84
rect -2033 56 -2018 84
rect -2018 56 -1999 84
rect -1960 56 -1950 84
rect -1950 56 -1926 84
rect -1887 56 -1882 84
rect -1882 56 -1853 84
rect -1814 56 -1780 90
rect -1741 84 -1707 90
rect -1668 84 -1634 90
rect -1595 84 -1561 90
rect -1522 84 -1488 90
rect -1449 84 -1415 90
rect -1376 84 -1342 90
rect -1303 84 -1269 90
rect -1230 84 -1196 90
rect -1157 84 -1123 90
rect -1084 84 -1050 90
rect -1011 84 -977 90
rect -938 84 -904 90
rect -865 84 -831 90
rect -792 84 -758 90
rect -719 84 -685 90
rect -646 84 -612 90
rect -573 84 -539 90
rect -500 84 -466 90
rect -427 84 -393 90
rect -354 84 -320 90
rect -281 84 -247 90
rect -208 84 -174 90
rect -135 84 -101 90
rect -62 84 -28 90
rect 11 84 45 90
rect 84 84 118 90
rect 157 84 191 90
rect 230 84 264 90
rect 303 84 337 90
rect 376 84 410 90
rect 448 84 482 90
rect 520 84 554 90
rect 592 84 626 90
rect 664 84 698 90
rect 736 84 770 90
rect 808 84 842 90
rect 880 84 914 90
rect 952 84 986 90
rect -1741 56 -1712 84
rect -1712 56 -1707 84
rect -1668 56 -1644 84
rect -1644 56 -1634 84
rect -1595 56 -1576 84
rect -1576 56 -1561 84
rect -1522 56 -1508 84
rect -1508 56 -1488 84
rect -1449 56 -1440 84
rect -1440 56 -1415 84
rect -1376 56 -1372 84
rect -1372 56 -1342 84
rect -1303 56 -1270 84
rect -1270 56 -1269 84
rect -1230 56 -1202 84
rect -1202 56 -1196 84
rect -1157 56 -1134 84
rect -1134 56 -1123 84
rect -1084 56 -1066 84
rect -1066 56 -1050 84
rect -1011 56 -998 84
rect -998 56 -977 84
rect -938 56 -930 84
rect -930 56 -904 84
rect -865 56 -862 84
rect -862 56 -831 84
rect -792 56 -760 84
rect -760 56 -758 84
rect -719 56 -692 84
rect -692 56 -685 84
rect -646 56 -624 84
rect -624 56 -612 84
rect -573 56 -556 84
rect -556 56 -539 84
rect -500 56 -488 84
rect -488 56 -466 84
rect -427 56 -420 84
rect -420 56 -393 84
rect -354 56 -352 84
rect -352 56 -320 84
rect -281 56 -250 84
rect -250 56 -247 84
rect -208 56 -182 84
rect -182 56 -174 84
rect -135 56 -114 84
rect -114 56 -101 84
rect -62 56 -46 84
rect -46 56 -28 84
rect 11 56 22 84
rect 22 56 45 84
rect 84 56 90 84
rect 90 56 118 84
rect 157 56 158 84
rect 158 56 191 84
rect 230 56 260 84
rect 260 56 264 84
rect 303 56 328 84
rect 328 56 337 84
rect 376 56 396 84
rect 396 56 410 84
rect 448 56 464 84
rect 464 56 482 84
rect 520 56 532 84
rect 532 56 554 84
rect 592 56 600 84
rect 600 56 626 84
rect 664 56 668 84
rect 668 56 698 84
rect 736 56 770 84
rect 808 56 838 84
rect 838 56 842 84
rect 880 56 906 84
rect 906 56 914 84
rect 952 56 974 84
rect 974 56 986 84
rect -2048 -201 -2014 -167
rect -2048 -273 -2014 -239
rect -2525 -408 -2491 -374
rect -2338 -380 -2304 -346
rect -1851 -306 -1817 -272
rect -2232 -369 -2198 -335
rect -2160 -369 -2126 -335
rect -1469 -308 -1435 -274
rect -884 -290 -850 -256
rect -811 -290 -777 -256
rect 169 -137 203 -103
rect -1851 -380 -1817 -346
rect -1767 -380 -1733 -346
rect -1651 -369 -1617 -335
rect -1579 -369 -1545 -335
rect -1469 -380 -1435 -346
rect -1365 -369 -1331 -335
rect -1293 -369 -1259 -335
rect -1947 -414 -1913 -380
rect -1163 -414 -1129 -380
rect -1091 -414 -1057 -380
rect -891 -381 -857 -347
rect -787 -369 -753 -335
rect -715 -369 -681 -335
rect -592 -348 -558 -314
rect -506 -414 -472 -380
rect -321 -391 -287 -357
rect -33 -242 1 -208
rect 169 -209 203 -175
rect 452 -137 486 -103
rect 452 -209 486 -175
rect -33 -314 1 -280
rect 834 -306 868 -272
rect -223 -394 -189 -360
rect -151 -394 -117 -360
rect 563 -385 597 -351
rect 635 -385 669 -351
rect 744 -384 778 -350
rect 834 -378 868 -344
rect 1033 -306 1067 -272
rect 1033 -378 1067 -344
rect -2518 -744 -2484 -735
rect -2518 -769 -2506 -744
rect -2506 -769 -2484 -744
rect -2445 -769 -2411 -735
rect -2372 -744 -2338 -735
rect -2372 -769 -2369 -744
rect -2369 -769 -2338 -744
rect -2299 -769 -2265 -735
rect -2226 -744 -2192 -735
rect -2226 -769 -2198 -744
rect -2198 -769 -2192 -744
rect -2153 -769 -2119 -735
rect -2080 -744 -2046 -735
rect -2080 -769 -2061 -744
rect -2061 -769 -2046 -744
rect -2007 -769 -1973 -735
rect -1934 -744 -1900 -735
rect -1934 -769 -1924 -744
rect -1924 -769 -1900 -744
rect -1861 -769 -1827 -735
rect -1788 -744 -1754 -735
rect -1788 -769 -1787 -744
rect -1787 -769 -1754 -744
rect -1715 -744 -1681 -735
rect -1715 -769 -1684 -744
rect -1684 -769 -1681 -744
rect -1642 -769 -1608 -735
rect -1570 -744 -1536 -735
rect -1570 -769 -1547 -744
rect -1547 -769 -1536 -744
rect -1498 -769 -1464 -735
rect -1426 -744 -1392 -735
rect -1426 -769 -1410 -744
rect -1410 -769 -1392 -744
rect -1354 -769 -1320 -735
rect -1282 -744 -1248 -735
rect -1282 -769 -1273 -744
rect -1273 -769 -1248 -744
rect -1210 -769 -1176 -735
rect -1138 -744 -1104 -735
rect -1138 -769 -1136 -744
rect -1136 -769 -1104 -744
rect -1066 -769 -1032 -735
rect -994 -744 -960 -735
rect -994 -769 -965 -744
rect -965 -769 -960 -744
rect -922 -769 -888 -735
rect -850 -744 -816 -735
rect -850 -769 -828 -744
rect -828 -769 -816 -744
rect -778 -769 -744 -735
rect -706 -744 -672 -735
rect -706 -769 -691 -744
rect -691 -769 -672 -744
rect -634 -769 -600 -735
rect -562 -744 -528 -735
rect -562 -769 -554 -744
rect -554 -769 -528 -744
rect -490 -769 -456 -735
rect -418 -744 -384 -735
rect -418 -769 -417 -744
rect -417 -769 -384 -744
rect -346 -744 -312 -735
rect -346 -769 -314 -744
rect -314 -769 -312 -744
rect -274 -769 -240 -735
rect -202 -744 -168 -735
rect -202 -769 -177 -744
rect -177 -769 -168 -744
rect -130 -769 -96 -735
rect -58 -744 -24 -735
rect -58 -769 -40 -744
rect -40 -769 -24 -744
rect 14 -769 48 -735
rect 86 -744 120 -735
rect 86 -769 96 -744
rect 96 -769 120 -744
rect 158 -769 192 -735
rect 230 -744 264 -735
rect 230 -769 232 -744
rect 232 -769 264 -744
rect 302 -769 336 -735
rect 374 -744 408 -735
rect 374 -769 402 -744
rect 402 -769 408 -744
rect 446 -769 480 -735
rect 518 -744 552 -735
rect 518 -769 538 -744
rect 538 -769 552 -744
rect 590 -769 624 -735
rect 662 -744 696 -735
rect 662 -769 674 -744
rect 674 -769 696 -744
rect 734 -769 768 -735
rect 806 -744 840 -735
rect 806 -769 810 -744
rect 810 -769 840 -744
rect 878 -769 912 -735
rect 950 -769 984 -735
rect -2239 -969 -2205 -935
rect -2165 -969 -2131 -935
rect -2091 -969 -2057 -935
rect -2017 -969 -1998 -935
rect -1998 -969 -1983 -935
rect -1943 -969 -1928 -935
rect -1928 -969 -1909 -935
rect -1869 -969 -1858 -935
rect -1858 -969 -1835 -935
rect -1795 -969 -1788 -935
rect -1788 -969 -1761 -935
rect -1721 -969 -1719 -935
rect -1719 -969 -1687 -935
rect -1647 -969 -1616 -935
rect -1616 -969 -1613 -935
rect -1574 -969 -1547 -935
rect -1547 -969 -1540 -935
rect -1501 -969 -1478 -935
rect -1478 -969 -1467 -935
rect -1428 -969 -1409 -935
rect -1409 -969 -1394 -935
rect -1355 -969 -1340 -935
rect -1340 -969 -1321 -935
rect -1282 -969 -1271 -935
rect -1271 -969 -1248 -935
rect -1209 -969 -1202 -935
rect -1202 -969 -1175 -935
rect -1136 -969 -1133 -935
rect -1133 -969 -1102 -935
rect -1063 -969 -1029 -935
rect -990 -969 -960 -935
rect -960 -969 -956 -935
rect -917 -969 -891 -935
rect -891 -969 -883 -935
rect -844 -969 -822 -935
rect -822 -969 -810 -935
rect -771 -969 -753 -935
rect -753 -969 -737 -935
rect -698 -969 -684 -935
rect -684 -969 -664 -935
rect -625 -969 -615 -935
rect -615 -969 -591 -935
rect -552 -969 -546 -935
rect -546 -969 -518 -935
rect -479 -969 -477 -935
rect -477 -969 -445 -935
rect -406 -969 -374 -935
rect -374 -969 -372 -935
rect -333 -969 -305 -935
rect -305 -969 -299 -935
rect -260 -969 -236 -935
rect -236 -969 -226 -935
rect -187 -969 -167 -935
rect -167 -969 -153 -935
rect -114 -969 -98 -935
rect -98 -969 -80 -935
rect -41 -969 -29 -935
rect -29 -969 -7 -935
rect 32 -969 40 -935
rect 40 -969 66 -935
rect 105 -969 109 -935
rect 109 -969 139 -935
rect 178 -969 212 -935
rect -2154 -1049 -2120 -1015
rect -2154 -1095 -2120 -1087
rect -2154 -1121 -2120 -1095
rect -1802 -1049 -1768 -1015
rect -1802 -1095 -1768 -1087
rect -1802 -1121 -1768 -1095
rect -2008 -1357 -1978 -1337
rect -1978 -1357 -1974 -1337
rect -2008 -1371 -1974 -1357
rect -1936 -1371 -1902 -1337
rect -2070 -1559 -2036 -1543
rect -2070 -1577 -2064 -1559
rect -2064 -1577 -2036 -1559
rect -2070 -1627 -2036 -1615
rect -2070 -1649 -2064 -1627
rect -2064 -1649 -2036 -1627
rect -1450 -1049 -1416 -1015
rect -1450 -1095 -1416 -1087
rect -1450 -1121 -1416 -1095
rect -1855 -1573 -1821 -1539
rect -1725 -1559 -1691 -1543
rect -1855 -1645 -1821 -1611
rect -1725 -1577 -1711 -1559
rect -1711 -1577 -1691 -1559
rect -1725 -1627 -1691 -1615
rect -1725 -1649 -1711 -1627
rect -1711 -1649 -1691 -1627
rect -1626 -1577 -1592 -1543
rect -1626 -1649 -1592 -1615
rect -1539 -1216 -1505 -1182
rect -1539 -1288 -1505 -1254
rect -1251 -1049 -1217 -1015
rect -1251 -1095 -1217 -1087
rect -1251 -1121 -1217 -1095
rect -1159 -1353 -1125 -1319
rect -1159 -1425 -1125 -1391
rect -899 -1049 -865 -1015
rect -899 -1095 -865 -1087
rect -899 -1121 -865 -1095
rect -1323 -1720 -1289 -1686
rect -1251 -1720 -1217 -1686
rect -1802 -1789 -1768 -1766
rect -1802 -1800 -1768 -1789
rect -1802 -1872 -1768 -1838
rect -993 -1294 -959 -1260
rect -993 -1366 -959 -1332
rect -786 -1049 -752 -1015
rect -786 -1095 -752 -1087
rect -786 -1121 -752 -1095
rect -695 -1368 -661 -1334
rect -695 -1440 -661 -1406
rect -881 -1577 -847 -1543
rect -809 -1577 -775 -1543
rect -899 -1789 -865 -1766
rect -899 -1800 -865 -1789
rect -899 -1872 -865 -1838
rect -434 -1049 -400 -1015
rect -434 -1095 -400 -1087
rect -434 -1121 -400 -1095
rect -519 -1368 -485 -1334
rect -519 -1440 -485 -1406
rect -318 -1049 -284 -1015
rect -318 -1095 -284 -1087
rect -318 -1121 -284 -1095
rect 121 -1197 155 -1176
rect 121 -1210 153 -1197
rect 153 -1210 155 -1197
rect 193 -1210 227 -1176
rect 505 -1049 539 -1015
rect 505 -1095 539 -1087
rect 505 -1121 539 -1095
rect -210 -1510 -176 -1476
rect -138 -1510 -104 -1476
rect 415 -1210 449 -1176
rect 415 -1282 449 -1248
rect -286 -1644 -252 -1610
rect -214 -1627 -180 -1610
rect -214 -1644 -196 -1627
rect -196 -1644 -180 -1627
rect -434 -1789 -400 -1766
rect -434 -1800 -400 -1789
rect -434 -1872 -400 -1838
rect -318 -1789 -284 -1766
rect -318 -1800 -284 -1789
rect -318 -1872 -284 -1838
rect -67 -1627 -33 -1610
rect -67 -1644 -52 -1627
rect -52 -1644 -33 -1627
rect 5 -1644 39 -1610
rect 183 -1647 217 -1613
rect 255 -1627 289 -1613
rect 255 -1647 273 -1627
rect 273 -1647 289 -1627
rect 34 -1789 68 -1766
rect 34 -1800 68 -1789
rect 34 -1872 68 -1838
rect 153 -1789 187 -1766
rect 153 -1800 187 -1789
rect 153 -1872 187 -1838
rect 1290 -1200 1324 -1166
rect 1362 -1200 1396 -1166
rect 4702 -1198 4736 -1164
rect 4774 -1198 4808 -1164
rect 1290 -1355 1324 -1321
rect 1362 -1355 1396 -1321
rect 4639 -1354 4673 -1320
rect 4711 -1354 4745 -1320
rect 1290 -1505 1324 -1471
rect 1362 -1505 1396 -1471
rect 4556 -1507 4590 -1473
rect 4628 -1507 4662 -1473
rect 1290 -1661 1324 -1627
rect 1362 -1661 1396 -1627
rect 4562 -1664 4596 -1630
rect 4634 -1664 4668 -1630
rect 505 -1789 539 -1766
rect 505 -1800 539 -1789
rect 505 -1872 539 -1838
rect -2185 -1970 -2179 -1936
rect -2179 -1970 -2151 -1936
rect -2111 -1970 -2077 -1936
rect -2037 -1970 -2036 -1936
rect -2036 -1970 -2003 -1936
rect -1963 -1970 -1929 -1936
rect -1889 -1970 -1855 -1936
rect -1815 -1970 -1784 -1936
rect -1784 -1970 -1781 -1936
rect -1741 -1970 -1707 -1936
rect -1667 -1970 -1641 -1936
rect -1641 -1970 -1633 -1936
rect -1593 -1970 -1559 -1936
rect -1519 -1970 -1498 -1936
rect -1498 -1970 -1485 -1936
rect -1445 -1970 -1411 -1936
rect -1372 -1970 -1355 -1936
rect -1355 -1970 -1338 -1936
rect -1299 -1970 -1265 -1936
rect -1226 -1970 -1212 -1936
rect -1212 -1970 -1192 -1936
rect -1153 -1970 -1119 -1936
rect -1080 -1970 -1069 -1936
rect -1069 -1970 -1046 -1936
rect -1007 -1970 -973 -1936
rect -934 -1970 -926 -1936
rect -926 -1970 -900 -1936
rect -861 -1970 -827 -1936
rect -788 -1970 -783 -1936
rect -783 -1970 -754 -1936
rect -715 -1970 -681 -1936
rect -642 -1970 -640 -1936
rect -640 -1970 -608 -1936
rect -569 -1970 -535 -1936
rect -496 -1970 -463 -1936
rect -463 -1970 -462 -1936
rect -423 -1970 -389 -1936
rect -350 -1970 -320 -1936
rect -320 -1970 -316 -1936
rect -277 -1970 -243 -1936
rect -204 -1970 -178 -1936
rect -178 -1970 -170 -1936
rect -131 -1970 -97 -1936
rect -58 -1970 -36 -1936
rect -36 -1970 -24 -1936
rect 15 -1970 49 -1936
rect 88 -1970 106 -1936
rect 106 -1970 122 -1936
rect 161 -1970 195 -1936
rect 234 -1970 248 -1936
rect 248 -1970 268 -1936
rect 307 -1970 341 -1936
rect 380 -1970 390 -1936
rect 390 -1970 414 -1936
rect 453 -1970 487 -1936
rect 526 -1970 532 -1936
rect 532 -1970 560 -1936
rect 1715 -2581 1749 -2547
rect 1715 -2653 1749 -2619
rect 1549 -2738 1583 -2704
rect 1621 -2738 1655 -2704
<< metal1 >>
rect -2660 1070 -492 1104
rect -2660 728 -2626 1070
rect -526 990 -492 1070
rect -526 956 -398 990
rect -404 938 -398 956
rect -346 938 -334 990
rect -282 973 308 990
rect -282 956 186 973
rect -282 938 -276 956
rect 180 921 186 956
rect 238 921 250 973
rect 302 921 308 973
rect -1404 831 -732 863
rect -1404 797 -1373 831
rect -1339 797 -1277 831
rect -1243 797 -1181 831
rect -1147 797 -1085 831
rect -1051 797 -989 831
rect -955 797 -893 831
rect -859 797 -797 831
rect -763 797 -732 831
rect -1404 765 -732 797
rect 420 765 516 863
rect 646 773 674 801
rect 1333 796 1385 802
rect -2659 676 -2653 728
rect -2601 676 -2589 728
rect -2537 676 -2531 728
rect -2068 723 -2022 735
rect -2068 689 -2062 723
rect -2028 689 -2022 723
rect -2068 657 -2022 689
rect -1813 685 -1807 737
rect -1755 685 -1743 737
rect -1691 735 -1685 737
rect -1691 728 -411 735
rect 1333 732 1385 744
rect -1691 694 -529 728
rect -495 694 -457 728
rect -423 694 -411 728
rect -1691 685 -411 694
rect -236 730 -190 731
rect -236 719 1333 730
rect -236 685 -230 719
rect -196 690 1333 719
rect -196 685 -190 690
rect -2068 651 -690 657
rect -2068 617 -2062 651
rect -2028 648 -690 651
tri -690 648 -681 657 sw
rect -2028 642 -681 648
tri -681 642 -675 648 sw
rect -236 642 -190 685
rect 1333 674 1385 680
rect 1421 801 1473 807
rect 1421 735 1473 749
rect 1421 677 1473 683
rect 1575 801 1627 807
rect 1575 735 1627 749
rect 1575 677 1627 683
rect 1727 801 1779 807
rect 1727 735 1779 749
rect 1727 677 1779 683
rect 2669 801 2721 807
rect 2818 795 2864 807
rect 2818 791 2824 795
rect 2669 735 2721 749
rect 2669 677 2721 683
rect 2815 785 2824 791
rect 2858 791 2864 795
rect 2858 785 2867 791
rect 2972 772 3018 784
rect 2972 740 2978 772
rect 3012 740 3018 772
rect 2815 723 2867 733
rect 2815 719 2824 723
rect 2858 719 2867 723
rect 2936 688 2942 740
rect 2994 700 3008 738
rect 3060 688 3066 740
rect 2815 661 2867 667
rect 2972 666 2978 688
rect 3012 666 3018 688
rect -2028 627 -675 642
rect -2028 617 -2022 627
rect -2068 605 -2022 617
tri -724 611 -708 627 ne
rect -708 610 -675 627
tri -675 610 -643 642 sw
tri -2010 576 -2006 580 se
rect -2006 576 -1710 580
tri -2014 572 -2010 576 se
rect -2010 572 -1710 576
tri -2035 551 -2014 572 se
rect -2014 552 -1762 572
rect -2014 551 -1995 552
tri -1995 551 -1994 552 nw
tri -1780 551 -1779 552 ne
rect -1779 551 -1762 552
rect -2242 545 -2008 551
rect -2242 511 -2230 545
rect -2196 511 -2153 545
rect -2119 538 -2008 545
tri -2008 538 -1995 551 nw
tri -1779 546 -1774 551 ne
rect -1774 538 -1762 551
rect -1728 538 -1710 572
rect -1660 555 -1654 561
rect -2119 518 -2028 538
tri -2028 518 -2008 538 nw
rect -1774 532 -1710 538
rect -1667 549 -1654 555
rect -1954 518 -1807 524
rect -2119 511 -2041 518
rect -2533 500 -2403 506
rect -2242 505 -2041 511
tri -2041 505 -2028 518 nw
rect -2533 466 -2521 500
rect -2487 466 -2449 500
rect -2415 466 -2403 500
rect -1954 484 -1942 518
rect -1908 515 -1807 518
tri -1807 515 -1798 524 sw
rect -1667 515 -1655 549
rect -1908 503 -1798 515
tri -1798 503 -1786 515 sw
rect -1667 509 -1654 515
rect -1602 509 -1590 561
rect -1538 509 -1532 561
rect -953 558 -907 570
rect -1238 537 -1108 543
rect -1382 523 -1330 529
rect -1908 500 -1786 503
tri -1786 500 -1783 503 sw
rect -1908 489 -1783 500
tri -1783 489 -1772 500 sw
rect -1908 484 -1772 489
rect -1954 483 -1772 484
tri -1772 483 -1766 489 sw
rect -1954 482 -1766 483
tri -1766 482 -1765 483 sw
rect -1495 482 -1449 494
rect -1954 478 -1765 482
rect -2533 460 -2403 466
tri -1832 460 -1814 478 ne
rect -1814 460 -1765 478
tri -1814 448 -1802 460 ne
rect -1802 448 -1765 460
tri -1765 448 -1731 482 sw
rect -1495 448 -1489 482
rect -1455 448 -1449 482
tri -1802 435 -1789 448 ne
rect -1789 435 -1731 448
tri -1731 435 -1718 448 sw
tri -1789 429 -1783 435 ne
rect -1783 429 -1718 435
tri -1718 429 -1712 435 sw
tri -1783 416 -1770 429 ne
rect -1770 416 -1712 429
rect -1495 425 -1449 448
rect -1399 471 -1382 475
rect -1238 503 -1226 537
rect -1192 503 -1154 537
rect -1120 503 -1108 537
rect -1238 497 -1108 503
rect -1330 471 -1267 475
rect -1399 469 -1267 471
rect -1399 435 -1387 469
rect -1353 459 -1313 469
rect -1330 435 -1313 459
rect -1279 435 -1267 469
rect -1399 429 -1382 435
rect -1878 404 -1813 416
tri -1770 412 -1766 416 ne
rect -1878 370 -1853 404
rect -1819 370 -1813 404
rect -1878 332 -1813 370
rect -1878 298 -1853 332
rect -1819 298 -1813 332
rect -1766 334 -1712 416
rect -1660 421 -1449 425
rect -1660 369 -1654 421
rect -1602 369 -1590 421
rect -1538 410 -1449 421
rect -1538 376 -1489 410
rect -1455 376 -1449 410
rect -1330 429 -1267 435
rect -1382 401 -1330 407
rect -1160 401 -1108 497
rect -953 524 -947 558
rect -913 524 -907 558
rect -953 483 -907 524
rect -796 559 -744 565
rect -708 563 -643 610
rect -236 608 -230 642
rect -196 608 -190 642
rect -236 596 -190 608
rect -119 654 -67 660
rect -119 590 -67 602
rect -708 557 -645 563
rect -708 523 -696 557
rect -662 523 -645 557
rect -708 517 -645 523
rect -521 557 -454 563
rect -521 523 -509 557
rect -475 523 -454 557
tri -522 508 -521 509 se
rect -521 508 -454 523
rect -796 495 -744 507
rect -953 449 -947 483
rect -913 449 -796 483
rect -953 443 -796 449
tri -541 489 -522 508 se
rect -522 489 -454 508
rect -409 507 -403 559
rect -351 507 -339 559
rect -287 554 -281 559
rect -287 548 -274 554
rect -286 514 -274 548
rect 166 629 218 635
rect 263 606 269 658
rect 321 606 333 658
rect 385 650 391 658
rect 2972 654 3018 666
rect 385 640 1211 650
rect 385 618 1388 640
rect 385 606 391 618
rect 1179 608 1388 618
rect -119 532 -67 538
rect 48 568 100 574
rect -119 530 -73 532
rect -287 508 -274 514
rect -287 507 -281 508
tri -547 483 -541 489 se
rect -541 486 -454 489
rect -541 483 -485 486
rect -744 455 -485 483
tri -485 455 -454 486 nw
rect 48 504 100 516
rect 166 565 218 577
rect 4426 597 4432 649
rect 4484 597 4498 649
rect 4550 597 4556 649
rect 166 507 218 513
rect 253 568 318 574
rect 253 562 266 568
rect 253 528 259 562
rect 253 516 266 528
rect 169 504 215 507
rect 253 504 318 516
rect -744 446 -494 455
tri -494 446 -485 455 nw
rect 48 446 100 452
rect -744 443 -503 446
rect -953 437 -503 443
tri -503 437 -494 446 nw
rect 54 443 100 446
rect 253 489 266 504
rect 253 455 259 489
rect 253 452 266 455
rect 253 446 318 452
rect 346 542 392 564
rect 346 508 352 542
rect 386 508 392 542
rect 253 443 299 446
rect -1538 369 -1449 376
rect -1160 377 185 401
tri 185 377 209 401 sw
tri 327 377 346 396 se
rect 346 377 392 508
rect 554 552 600 564
rect 554 518 560 552
rect 594 518 600 552
rect 1234 522 1286 528
rect 554 480 600 518
rect 554 446 560 480
rect 594 446 600 480
rect 939 515 1069 521
rect 939 481 951 515
rect 985 481 1023 515
rect 1057 481 1069 515
rect 939 475 1069 481
tri 553 397 554 398 se
rect 554 397 600 446
rect 1234 458 1286 470
tri 392 377 412 397 sw
tri 533 377 553 397 se
rect 553 377 600 397
rect -1160 373 600 377
rect -1660 364 -1449 369
tri 160 364 169 373 ne
rect 169 364 576 373
tri 169 349 184 364 ne
rect 184 349 576 364
tri 576 349 600 373 nw
tri 636 406 664 434 se
rect 664 406 1234 434
rect 2143 457 2171 485
rect 2973 474 3025 480
rect 636 404 1286 406
rect -796 334 -790 345
rect -1766 306 -790 334
rect -1878 265 -1813 298
rect -796 293 -790 306
rect -738 293 -726 345
rect -674 293 -668 345
rect -572 293 -566 345
rect -514 293 -502 345
rect -450 309 -148 345
tri -148 309 -112 345 sw
tri 634 343 636 345 se
rect 636 343 666 404
tri 666 393 677 404 nw
rect 1234 400 1286 404
rect 2973 408 3025 422
rect 1076 368 1128 374
rect -450 308 -112 309
rect -450 293 -444 308
tri -159 293 -144 308 ne
rect -144 293 -112 308
tri -144 278 -129 293 ne
rect -129 278 -112 293
rect -330 265 -324 278
rect -1878 235 -324 265
rect -330 226 -324 235
rect -272 226 -260 278
rect -208 265 -202 278
tri -129 267 -118 278 ne
rect -118 267 -112 278
tri -112 267 -70 309 sw
rect -34 291 -28 343
rect 24 291 36 343
rect 88 321 94 343
tri 612 321 634 343 se
rect 634 327 666 343
rect 634 321 660 327
tri 660 321 666 327 nw
tri 705 321 732 348 se
rect 732 321 1076 348
rect 88 291 630 321
tri 630 291 660 321 nw
tri 692 308 705 321 se
rect 705 320 1076 321
rect 705 308 732 320
tri 732 308 744 320 nw
rect 4426 459 4556 597
rect 4426 407 4432 459
rect 4484 407 4498 459
rect 4550 407 4556 459
tri 675 291 692 308 se
tri 662 278 675 291 se
rect 675 278 692 291
tri 652 268 662 278 se
rect 662 268 692 278
tri 692 268 732 308 nw
rect 1076 304 1128 316
rect 833 273 839 279
tri 651 267 652 268 se
rect 652 267 691 268
tri 691 267 692 268 nw
rect 765 267 839 273
tri -118 265 -116 267 ne
rect -116 265 -70 267
rect -208 235 -201 265
tri -116 261 -112 265 ne
rect -112 261 -70 265
tri -70 261 -64 267 sw
tri 645 261 651 267 se
rect 651 261 657 267
tri -112 235 -86 261 ne
rect -86 235 657 261
rect -208 226 -202 235
tri -86 233 -84 235 ne
rect -84 233 657 235
tri 657 233 691 267 nw
rect 765 233 777 267
rect 811 233 839 267
rect 765 227 839 233
rect 891 227 903 279
rect 955 227 961 279
rect 1076 246 1128 252
rect 2505 316 2557 322
rect 2505 252 2557 264
rect -1404 195 -732 197
rect -2556 187 1092 195
rect 2505 194 2557 200
rect -2556 165 -790 187
rect -2556 131 -1373 165
rect -1339 131 -1277 165
rect -1243 131 -1181 165
rect -1147 131 -1085 165
rect -1051 131 -989 165
rect -955 131 -893 165
rect -859 131 -797 165
rect -738 135 -725 187
rect -673 135 -660 187
rect -608 135 -595 187
rect -543 135 -530 187
rect -478 135 -465 187
rect -413 135 -400 187
rect -348 135 -335 187
rect -283 135 -270 187
rect -218 135 1092 187
rect -763 131 1092 135
rect -2556 123 1092 131
rect -2556 90 -790 123
rect -2556 56 -2544 90
rect -2510 56 -2471 90
rect -2437 56 -2398 90
rect -2364 56 -2325 90
rect -2291 56 -2252 90
rect -2218 56 -2179 90
rect -2145 56 -2106 90
rect -2072 56 -2033 90
rect -1999 56 -1960 90
rect -1926 56 -1887 90
rect -1853 56 -1814 90
rect -1780 56 -1741 90
rect -1707 56 -1668 90
rect -1634 56 -1595 90
rect -1561 56 -1522 90
rect -1488 56 -1449 90
rect -1415 56 -1376 90
rect -1342 56 -1303 90
rect -1269 56 -1230 90
rect -1196 56 -1157 90
rect -1123 56 -1084 90
rect -1050 56 -1011 90
rect -977 56 -938 90
rect -904 56 -865 90
rect -831 56 -792 90
rect -738 71 -725 123
rect -673 71 -660 123
rect -608 71 -595 123
rect -543 90 -530 123
rect -478 90 -465 123
rect -413 90 -400 123
rect -348 90 -335 123
rect -283 90 -270 123
rect -218 90 1092 123
rect -539 71 -530 90
rect -466 71 -465 90
rect -283 71 -281 90
rect -218 71 -208 90
rect -758 59 -719 71
rect -685 59 -646 71
rect -612 59 -573 71
rect -539 59 -500 71
rect -466 59 -427 71
rect -393 59 -354 71
rect -320 59 -281 71
rect -247 59 -208 71
rect -2556 7 -790 56
rect -738 7 -725 59
rect -673 7 -660 59
rect -608 7 -595 59
rect -539 56 -530 59
rect -466 56 -465 59
rect -283 56 -281 59
rect -218 56 -208 59
rect -174 56 -135 90
rect -101 56 -62 90
rect -28 56 11 90
rect 45 56 84 90
rect 118 56 157 90
rect 191 56 230 90
rect 264 56 303 90
rect 337 56 376 90
rect 410 56 448 90
rect 482 56 520 90
rect 554 56 592 90
rect 626 56 664 90
rect 698 56 736 90
rect 770 56 808 90
rect 842 56 880 90
rect 914 56 952 90
rect 986 56 1092 90
rect -543 7 -530 56
rect -478 7 -465 56
rect -413 7 -400 56
rect -348 7 -335 56
rect -283 7 -270 56
rect -218 7 1092 56
rect -2556 -5 1092 7
rect -2556 -57 -790 -5
rect -738 -57 -725 -5
rect -673 -57 -660 -5
rect -608 -57 -595 -5
rect -543 -57 -530 -5
rect -478 -57 -465 -5
rect -413 -57 -400 -5
rect -348 -57 -335 -5
rect -283 -57 -270 -5
rect -218 -57 1092 -5
rect -2556 -63 1092 -57
rect -1254 -143 -1246 -91
rect -1194 -143 -1182 -91
rect -1130 -97 238 -91
rect -1130 -103 186 -97
rect -1130 -137 169 -103
rect -1130 -143 186 -137
rect 163 -149 186 -143
rect -2057 -161 -2005 -155
rect 163 -161 238 -149
rect 163 -175 186 -161
rect 39 -182 91 -176
rect -2057 -225 -2005 -213
rect -2057 -283 -2005 -277
rect -1953 -190 -1901 -184
rect -1255 -234 -1249 -182
rect -1197 -234 -1185 -182
rect -1133 -214 -391 -182
rect -1133 -234 -1127 -214
rect -397 -234 -391 -214
rect -339 -234 -327 -182
rect -275 -234 -269 -182
rect -191 -202 7 -196
rect -1953 -254 -1901 -242
rect -2054 -285 -2008 -283
rect -1901 -272 -1811 -260
rect -1901 -306 -1851 -272
rect -1817 -306 -1811 -272
rect -1953 -312 -1811 -306
rect -2344 -333 -2298 -321
rect -2531 -374 -2485 -349
rect -2531 -408 -2525 -374
rect -2491 -408 -2485 -374
rect -2425 -385 -2419 -333
rect -2367 -385 -2355 -333
rect -2303 -385 -2297 -333
rect -2244 -381 -2238 -329
rect -2186 -381 -2174 -329
rect -2122 -375 -2114 -329
rect -1857 -346 -1811 -312
rect -2122 -381 -2116 -375
rect -1959 -380 -1888 -374
rect -2344 -392 -2298 -385
rect -2531 -420 -2485 -408
rect -1959 -414 -1947 -380
rect -1913 -414 -1888 -380
rect -1857 -380 -1851 -346
rect -1817 -380 -1811 -346
rect -1857 -392 -1811 -380
rect -1776 -270 -1724 -264
rect -1776 -334 -1724 -322
rect -1776 -392 -1724 -386
rect -1663 -270 -1611 -264
rect -1663 -329 -1611 -322
rect -1478 -268 -1426 -262
rect -896 -298 -890 -246
rect -838 -298 -823 -246
rect -771 -298 -765 -246
rect -721 -251 -669 -245
rect -1663 -334 -1533 -329
rect -1611 -335 -1533 -334
rect -1611 -369 -1579 -335
rect -1545 -369 -1533 -335
rect -1611 -375 -1533 -369
rect -1478 -334 -1426 -320
rect -139 -208 7 -202
rect -139 -242 -33 -208
rect 1 -242 7 -208
rect -139 -254 7 -242
rect -191 -266 7 -254
rect -333 -281 -281 -275
rect -721 -317 -669 -303
rect -1663 -392 -1611 -386
rect -1377 -335 -1247 -329
rect -1377 -369 -1365 -335
rect -1331 -369 -1293 -335
rect -1259 -369 -1247 -335
rect -799 -335 -721 -329
rect -1377 -375 -1247 -369
rect -1478 -392 -1426 -386
rect -1175 -380 -1045 -374
rect -1959 -420 -1888 -414
rect -1175 -414 -1163 -380
rect -1129 -414 -1091 -380
rect -1057 -414 -1045 -380
rect -959 -391 -953 -339
rect -901 -347 -889 -339
rect -901 -381 -891 -347
rect -901 -391 -889 -381
rect -837 -391 -831 -339
rect -799 -369 -787 -335
rect -753 -369 -721 -335
rect -630 -345 -624 -293
rect -572 -314 -560 -293
rect -508 -345 -502 -293
rect -139 -280 7 -266
rect -139 -314 -33 -280
rect 1 -314 7 -280
rect -139 -318 7 -314
rect -191 -324 7 -318
rect -39 -326 7 -324
rect 163 -209 169 -175
rect 163 -213 186 -209
rect 163 -219 238 -213
rect 446 -103 659 -91
rect 446 -137 452 -103
rect 486 -137 659 -103
rect 446 -143 659 -137
rect 711 -143 723 -91
rect 775 -143 781 -91
rect 446 -175 492 -143
rect 446 -209 452 -175
rect 486 -209 492 -175
rect 163 -221 209 -219
rect 446 -221 492 -209
rect 2973 -196 3025 356
rect 3132 -76 3138 -24
rect 3190 -76 3202 -24
rect 3254 -76 3733 -24
rect 3146 -156 3152 -104
rect 3204 -156 3217 -104
rect 3269 -156 3733 -104
rect 3845 -119 3897 -113
rect 3845 -184 3897 -171
rect 39 -246 91 -234
rect 3146 -242 3152 -190
rect 3204 -242 3217 -190
rect 3269 -236 3845 -190
rect 3269 -242 3897 -236
rect 6433 -241 6485 -235
rect 39 -304 91 -298
rect -333 -345 -281 -333
rect -630 -348 -592 -345
rect -558 -348 -546 -345
rect -630 -354 -546 -348
rect -799 -375 -669 -369
rect 39 -354 77 -304
rect 125 -312 131 -260
rect 183 -312 195 -260
rect 247 -312 483 -260
rect 535 -312 547 -260
rect 599 -312 605 -260
rect 729 -262 781 -256
rect 1885 -259 1937 -253
rect 828 -262 874 -260
rect 961 -262 1073 -260
rect 729 -326 781 -314
rect -518 -380 -447 -374
rect -1175 -420 -1045 -414
rect -518 -414 -506 -380
rect -472 -414 -447 -380
rect -333 -403 -281 -397
rect -235 -360 77 -354
rect -235 -394 -223 -360
rect -189 -394 -151 -360
rect -117 -388 77 -360
rect 551 -351 681 -345
rect 551 -385 563 -351
rect 597 -385 635 -351
rect 669 -385 681 -351
rect -117 -394 -105 -388
rect 551 -391 681 -385
rect 719 -378 729 -344
rect 825 -268 877 -262
rect 825 -332 877 -320
rect 781 -378 790 -344
rect 719 -384 744 -378
rect 778 -384 790 -378
rect 719 -390 790 -384
rect 825 -390 877 -384
rect 909 -268 1073 -262
rect 961 -272 1073 -268
rect 961 -306 1033 -272
rect 1067 -306 1073 -272
rect 961 -320 1073 -306
rect 909 -332 1073 -320
rect 961 -344 1073 -332
rect 1885 -323 1937 -311
rect 2973 -262 3025 -248
rect 2973 -320 3025 -314
rect 3268 -280 3661 -274
rect 961 -378 1033 -344
rect 1067 -378 1073 -344
rect 961 -384 1073 -378
rect 909 -390 1073 -384
rect 1139 -340 1191 -334
rect -235 -400 -105 -394
rect 1885 -381 1937 -375
rect 3320 -332 3609 -280
rect 3268 -334 3661 -332
rect 3268 -344 3320 -334
rect -518 -420 -447 -414
rect -2531 -448 -447 -420
rect 1139 -404 1191 -392
rect 3268 -402 3320 -396
rect 3609 -344 3661 -334
rect 3609 -402 3661 -396
rect 6433 -305 6485 -293
tri -365 -448 -348 -431 se
rect -348 -448 1139 -431
tri -395 -478 -365 -448 se
rect -365 -456 1139 -448
rect -365 -463 1191 -456
rect 3183 -440 3235 -434
rect -365 -478 -337 -463
tri -337 -478 -322 -463 nw
rect -2244 -530 -2238 -478
rect -2186 -530 -2174 -478
rect -2122 -510 -369 -478
tri -369 -510 -337 -478 nw
rect -227 -493 1188 -491
rect -2122 -530 -2116 -510
rect -1663 -597 -1657 -545
rect -1605 -597 -1593 -545
rect -1541 -597 -1241 -545
rect -1189 -597 -1177 -545
rect -1125 -597 -1119 -545
rect -916 -591 -910 -539
rect -858 -591 -846 -539
rect -794 -575 -769 -539
tri -769 -575 -733 -539 sw
rect -227 -545 -221 -493
rect -169 -545 -157 -493
rect -105 -497 1188 -493
rect -105 -522 1136 -497
rect -105 -545 -99 -522
tri 723 -575 747 -551 se
rect 747 -575 755 -551
rect -794 -591 755 -575
tri -788 -597 -782 -591 ne
rect -782 -597 755 -591
tri -782 -603 -776 -597 ne
rect -776 -603 755 -597
rect 807 -603 819 -551
rect 871 -603 878 -551
rect 1136 -561 1188 -549
rect 3235 -448 3661 -442
rect 3235 -492 3609 -448
rect 3183 -500 3609 -492
rect 3183 -502 3661 -500
rect 3183 -504 3235 -502
rect 3183 -562 3235 -556
rect 3609 -512 3661 -502
rect 3609 -570 3661 -564
rect 3693 -528 3745 -522
rect 3693 -592 3745 -580
rect 1136 -619 1188 -613
rect -2556 -735 996 -631
rect 3140 -644 3693 -598
rect 3140 -650 3745 -644
rect 6433 -609 6485 -357
rect 6433 -661 6639 -609
rect 6431 -716 6483 -710
rect -2556 -769 -2518 -735
rect -2484 -769 -2445 -735
rect -2411 -769 -2372 -735
rect -2338 -769 -2299 -735
rect -2265 -769 -2226 -735
rect -2192 -769 -2153 -735
rect -2119 -769 -2080 -735
rect -2046 -769 -2007 -735
rect -1973 -769 -1934 -735
rect -1900 -769 -1861 -735
rect -1827 -769 -1788 -735
rect -1754 -769 -1715 -735
rect -1681 -769 -1642 -735
rect -1608 -769 -1570 -735
rect -1536 -769 -1498 -735
rect -1464 -769 -1426 -735
rect -1392 -769 -1354 -735
rect -1320 -769 -1282 -735
rect -1248 -769 -1210 -735
rect -1176 -769 -1138 -735
rect -1104 -769 -1066 -735
rect -1032 -769 -994 -735
rect -960 -769 -922 -735
rect -888 -769 -850 -735
rect -816 -769 -778 -735
rect -744 -769 -706 -735
rect -672 -769 -634 -735
rect -600 -769 -562 -735
rect -528 -769 -490 -735
rect -456 -769 -418 -735
rect -384 -769 -346 -735
rect -312 -769 -274 -735
rect -240 -769 -202 -735
rect -168 -769 -130 -735
rect -96 -769 -58 -735
rect -24 -769 14 -735
rect 48 -769 86 -735
rect 120 -769 158 -735
rect 192 -769 230 -735
rect 264 -769 302 -735
rect 336 -769 374 -735
rect 408 -769 446 -735
rect 480 -769 518 -735
rect 552 -769 590 -735
rect 624 -769 662 -735
rect 696 -769 734 -735
rect 768 -769 806 -735
rect 840 -769 878 -735
rect 912 -769 950 -735
rect 984 -769 996 -735
rect -2556 -775 996 -769
tri 3289 -775 3331 -733 se
rect 3331 -773 5020 -733
tri 5020 -773 5060 -733 sw
rect 3331 -775 5060 -773
tri 3248 -816 3289 -775 se
rect 3289 -816 5060 -775
rect 6113 -798 6119 -746
rect 6171 -798 6183 -746
rect 6235 -768 6431 -746
rect 6235 -780 6483 -768
rect 6235 -798 6431 -780
rect -2571 -868 -2565 -816
rect -2513 -868 -2501 -816
rect -2449 -868 -2443 -816
tri 3236 -828 3248 -816 se
rect 3248 -823 5060 -816
rect 3248 -828 3337 -823
rect 327 -834 333 -828
rect -2657 -1036 -2651 -984
rect -2599 -1036 -2587 -984
rect -2535 -1036 -2529 -984
rect -2574 -1599 -2529 -1036
rect -2487 -1510 -2443 -868
rect -2395 -874 333 -834
rect -2395 -900 -2355 -874
rect 327 -880 333 -874
rect 385 -880 397 -828
rect 449 -880 455 -828
tri 3188 -876 3236 -828 se
rect 3236 -876 3337 -828
tri 639 -880 643 -876 se
rect 643 -880 1072 -876
tri 1072 -880 1076 -876 sw
tri 3184 -880 3188 -876 se
rect 3188 -880 3337 -876
tri 3337 -880 3394 -823 nw
tri 4879 -852 4908 -823 ne
rect 4908 -852 5060 -823
rect 6431 -838 6483 -832
rect -2407 -906 -2355 -900
tri 590 -929 639 -880 se
rect 639 -929 3250 -880
rect -2251 -931 224 -929
tri 588 -931 590 -929 se
rect 590 -931 3250 -929
rect -2251 -932 3250 -931
rect -2407 -970 -2355 -958
rect -2407 -1028 -2355 -1022
rect -2255 -935 3250 -932
rect -2255 -969 -2239 -935
rect -2205 -969 -2165 -935
rect -2131 -969 -2091 -935
rect -2057 -969 -2017 -935
rect -1983 -969 -1943 -935
rect -1909 -969 -1869 -935
rect -1835 -969 -1795 -935
rect -1761 -969 -1721 -935
rect -1687 -969 -1647 -935
rect -1613 -969 -1574 -935
rect -1540 -969 -1501 -935
rect -1467 -969 -1428 -935
rect -1394 -969 -1355 -935
rect -1321 -969 -1282 -935
rect -1248 -969 -1209 -935
rect -1175 -969 -1136 -935
rect -1102 -969 -1063 -935
rect -1029 -969 -990 -935
rect -956 -969 -917 -935
rect -883 -969 -844 -935
rect -810 -942 -771 -935
rect -737 -942 -698 -935
rect -664 -942 -625 -935
rect -591 -942 -552 -935
rect -518 -942 -479 -935
rect -445 -942 -406 -935
rect -372 -942 -333 -935
rect -299 -942 -260 -935
rect -226 -942 -187 -935
rect -810 -969 -790 -942
rect -737 -969 -725 -942
rect -664 -969 -660 -942
rect -413 -969 -406 -942
rect -2255 -994 -790 -969
rect -738 -994 -725 -969
rect -673 -994 -660 -969
rect -608 -994 -595 -969
rect -543 -994 -530 -969
rect -478 -994 -465 -969
rect -413 -994 -400 -969
rect -348 -994 -335 -942
rect -283 -994 -270 -942
rect -218 -969 -187 -942
rect -153 -969 -114 -935
rect -80 -969 -41 -935
rect -7 -969 32 -935
rect 66 -969 105 -935
rect 139 -969 178 -935
rect 212 -967 3250 -935
tri 3250 -967 3337 -880 nw
rect 4403 -904 4409 -852
rect 4461 -904 4473 -852
rect 4525 -886 4531 -852
tri 4531 -886 4565 -852 sw
tri 4908 -881 4937 -852 ne
rect 4525 -904 4565 -886
tri 4467 -950 4513 -904 ne
rect 212 -969 3164 -967
rect -218 -974 3164 -969
rect -218 -994 662 -974
rect -2255 -1010 662 -994
rect -2255 -1015 -790 -1010
rect -2255 -1049 -2154 -1015
rect -2120 -1049 -1802 -1015
rect -1768 -1049 -1450 -1015
rect -1416 -1049 -1251 -1015
rect -1217 -1049 -899 -1015
rect -865 -1049 -790 -1015
rect -2255 -1062 -790 -1049
rect -738 -1062 -725 -1010
rect -673 -1062 -660 -1010
rect -608 -1062 -595 -1010
rect -543 -1062 -530 -1010
rect -478 -1062 -465 -1010
rect -413 -1015 -400 -1010
rect -413 -1062 -400 -1049
rect -348 -1062 -335 -1010
rect -283 -1062 -270 -1010
rect -218 -1015 662 -1010
rect -218 -1049 505 -1015
rect 539 -1049 662 -1015
tri 662 -1025 713 -974 nw
tri 2914 -1002 2942 -974 ne
rect 2942 -1000 3164 -974
tri 3164 -1000 3197 -967 nw
rect 2942 -1002 2957 -1000
rect -218 -1062 662 -1049
rect -2255 -1078 662 -1062
rect -2255 -1087 -790 -1078
rect -2255 -1121 -2154 -1087
rect -2120 -1121 -1802 -1087
rect -1768 -1121 -1450 -1087
rect -1416 -1121 -1251 -1087
rect -1217 -1121 -899 -1087
rect -865 -1121 -790 -1087
rect -2255 -1130 -790 -1121
rect -738 -1130 -725 -1078
rect -673 -1130 -660 -1078
rect -608 -1130 -595 -1078
rect -543 -1130 -530 -1078
rect -478 -1130 -465 -1078
rect -413 -1087 -400 -1078
rect -413 -1130 -400 -1121
rect -348 -1130 -335 -1078
rect -283 -1130 -270 -1078
rect -218 -1087 662 -1078
rect -218 -1121 505 -1087
rect 539 -1121 662 -1087
rect -218 -1130 662 -1121
rect -2255 -1134 662 -1130
rect 1148 -1030 1902 -1002
tri 2942 -1016 2956 -1002 ne
rect 2956 -1008 2957 -1002
rect 1148 -1036 1704 -1030
rect 1200 -1045 1704 -1036
rect 1148 -1112 1200 -1088
rect 1450 -1125 1456 -1073
rect 1508 -1125 1520 -1073
rect 1572 -1125 1578 -1073
rect 1698 -1082 1704 -1045
rect 1756 -1082 1774 -1030
rect 1826 -1082 1844 -1030
rect 1896 -1082 1902 -1030
rect 1529 -1155 1578 -1125
rect 2956 -1126 3168 -1008
rect 3211 -1059 3217 -1007
rect 3269 -1059 3281 -1007
rect 3333 -1013 3349 -1007
tri 3349 -1013 3355 -1007 sw
rect 3333 -1059 3355 -1013
tri 4497 -1153 4513 -1137 se
rect 4513 -1153 4565 -904
rect 4937 -911 5060 -852
rect 6588 -944 6639 -661
rect 6587 -950 6639 -944
rect 6587 -1014 6639 -1002
rect -1545 -1176 239 -1170
rect -1545 -1182 121 -1176
rect -1545 -1216 -1539 -1182
rect -1505 -1210 121 -1182
rect 155 -1210 193 -1176
rect 227 -1210 239 -1176
rect -1505 -1216 239 -1210
rect 327 -1216 333 -1164
rect 385 -1216 397 -1164
rect 449 -1216 455 -1164
rect 1148 -1170 1200 -1164
rect 1278 -1208 1284 -1156
rect 1336 -1208 1357 -1156
rect 1409 -1208 1415 -1156
rect 1529 -1191 2354 -1155
rect -2040 -1237 -1886 -1235
rect -2040 -1289 -2034 -1237
rect -1982 -1289 -1944 -1237
rect -1892 -1255 -1886 -1237
rect -1545 -1254 -1499 -1216
rect 409 -1248 455 -1216
tri 1256 -1236 1278 -1214 se
rect 1278 -1236 1408 -1208
rect -1892 -1289 -1732 -1255
rect -2040 -1291 -1732 -1289
rect -2040 -1328 -1886 -1326
rect -2040 -1380 -2034 -1328
rect -1982 -1337 -1944 -1328
rect -1974 -1371 -1944 -1337
rect -1982 -1380 -1944 -1371
rect -1892 -1380 -1886 -1328
rect -2040 -1382 -1886 -1380
rect -1768 -1394 -1732 -1291
rect -1545 -1288 -1539 -1254
rect -1505 -1288 -1499 -1254
rect -1545 -1300 -1499 -1288
rect -999 -1260 286 -1248
rect -999 -1294 -993 -1260
rect -959 -1264 286 -1260
tri 286 -1264 302 -1248 sw
rect -959 -1282 302 -1264
tri 302 -1282 320 -1264 sw
rect 409 -1282 415 -1248
rect 449 -1282 455 -1248
rect -959 -1294 320 -1282
rect -1165 -1319 -1119 -1307
rect -1165 -1353 -1159 -1319
rect -1125 -1353 -1119 -1319
rect -1165 -1391 -1119 -1353
rect -999 -1332 -953 -1294
tri 268 -1320 294 -1294 ne
rect 294 -1320 320 -1294
tri 320 -1320 358 -1282 sw
rect 409 -1294 455 -1282
tri 508 -1294 566 -1236 se
rect 566 -1282 1408 -1236
rect 566 -1294 571 -1282
tri 482 -1320 508 -1294 se
rect 508 -1320 571 -1294
tri 571 -1320 609 -1282 nw
tri 636 -1320 644 -1312 se
rect 644 -1320 1284 -1312
tri 294 -1321 295 -1320 ne
rect 295 -1321 358 -1320
tri 358 -1321 359 -1320 sw
tri 481 -1321 482 -1320 se
rect 482 -1321 570 -1320
tri 570 -1321 571 -1320 nw
tri 635 -1321 636 -1320 se
rect 636 -1321 1284 -1320
tri 295 -1322 296 -1321 ne
rect 296 -1322 359 -1321
rect -999 -1366 -993 -1332
rect -959 -1366 -953 -1332
rect -999 -1378 -953 -1366
rect -701 -1334 -655 -1322
rect -701 -1368 -695 -1334
rect -661 -1368 -655 -1334
rect -1768 -1401 -1277 -1394
rect -1165 -1401 -1159 -1391
rect -1768 -1425 -1159 -1401
rect -1125 -1425 -1119 -1391
rect -1768 -1430 -1119 -1425
rect -1313 -1437 -1119 -1430
rect -701 -1406 -655 -1368
rect -701 -1440 -695 -1406
rect -661 -1440 -655 -1406
rect -701 -1452 -655 -1440
rect -525 -1334 235 -1322
rect -525 -1368 -519 -1334
rect -485 -1346 235 -1334
tri 235 -1346 259 -1322 sw
tri 296 -1328 302 -1322 ne
rect 302 -1328 359 -1322
tri 359 -1328 366 -1321 sw
tri 477 -1325 481 -1321 se
rect 481 -1325 566 -1321
tri 566 -1325 570 -1321 nw
tri 631 -1325 635 -1321 se
rect 635 -1325 1284 -1321
tri 474 -1328 477 -1325 se
rect 477 -1328 536 -1325
tri 302 -1346 320 -1328 ne
rect 320 -1346 536 -1328
rect -485 -1355 259 -1346
tri 259 -1355 268 -1346 sw
tri 320 -1355 329 -1346 ne
rect 329 -1355 536 -1346
tri 536 -1355 566 -1325 nw
tri 601 -1355 631 -1325 se
rect 631 -1355 1284 -1325
rect -485 -1368 268 -1355
rect -525 -1406 -479 -1368
rect -525 -1440 -519 -1406
rect -485 -1440 -479 -1406
tri 217 -1410 259 -1368 ne
rect 259 -1375 268 -1368
tri 268 -1375 288 -1355 sw
tri 329 -1375 349 -1355 ne
rect 349 -1375 516 -1355
tri 516 -1375 536 -1355 nw
tri 581 -1375 601 -1355 se
rect 601 -1358 1284 -1355
rect 601 -1375 644 -1358
rect 259 -1410 288 -1375
tri 288 -1410 323 -1375 sw
tri 546 -1410 581 -1375 se
rect 581 -1401 644 -1375
tri 644 -1401 687 -1358 nw
rect 1278 -1364 1284 -1358
rect 1336 -1364 1350 -1312
rect 1402 -1364 1408 -1312
rect 581 -1410 588 -1401
rect -525 -1452 -479 -1440
tri 259 -1452 301 -1410 ne
rect 301 -1452 588 -1410
tri 301 -1457 306 -1452 ne
rect 306 -1457 588 -1452
tri 588 -1457 644 -1401 nw
rect -2076 -1470 -1408 -1459
tri -1408 -1470 -1397 -1459 sw
rect -2076 -1471 -725 -1470
tri -725 -1471 -724 -1470 sw
tri -428 -1471 -427 -1470 se
rect -427 -1471 -92 -1470
rect -2076 -1476 -724 -1471
tri -724 -1476 -719 -1471 sw
tri -433 -1476 -428 -1471 se
rect -428 -1476 -92 -1471
rect -2076 -1480 -719 -1476
tri -719 -1480 -715 -1476 sw
tri -437 -1480 -433 -1476 se
rect -433 -1480 -210 -1476
tri -2443 -1510 -2413 -1480 sw
rect -2076 -1490 -210 -1480
rect -2076 -1510 -2023 -1490
tri -2023 -1510 -2003 -1490 nw
tri -1442 -1508 -1424 -1490 ne
rect -1424 -1508 -210 -1490
tri -752 -1510 -750 -1508 ne
rect -750 -1510 -210 -1508
rect -176 -1510 -138 -1476
rect -104 -1510 -92 -1476
rect -2487 -1512 -2413 -1510
tri -2413 -1512 -2411 -1510 sw
rect -2487 -1564 -2481 -1512
rect -2429 -1564 -2417 -1512
rect -2365 -1564 -2359 -1512
rect -2076 -1543 -2030 -1510
tri -2030 -1517 -2023 -1510 nw
tri -750 -1516 -744 -1510 ne
rect -744 -1516 -92 -1510
rect 1278 -1514 1284 -1462
rect 1336 -1514 1350 -1462
rect 1402 -1514 1408 -1462
rect -1861 -1529 -1815 -1527
rect -2076 -1577 -2070 -1543
rect -2036 -1577 -2030 -1543
rect -2574 -1640 -2112 -1599
rect -2157 -1692 -2112 -1640
rect -2076 -1615 -2030 -1577
rect -2076 -1649 -2070 -1615
rect -2036 -1649 -2030 -1615
rect -2076 -1661 -2030 -1649
rect -1864 -1535 -1812 -1529
rect -1864 -1599 -1812 -1587
rect -1864 -1657 -1812 -1651
rect -1739 -1531 -1687 -1529
rect -1739 -1535 -1685 -1531
rect -1687 -1587 -1685 -1535
rect -1739 -1599 -1685 -1587
rect -1687 -1651 -1685 -1599
rect -1739 -1657 -1685 -1651
rect -1731 -1661 -1685 -1657
rect -1632 -1537 -1580 -1531
rect -893 -1543 -763 -1537
rect -893 -1577 -881 -1543
rect -847 -1577 -809 -1543
rect -775 -1545 -763 -1543
rect -775 -1575 301 -1545
rect -775 -1577 -763 -1575
rect -893 -1583 -763 -1577
tri 138 -1583 146 -1575 ne
rect 146 -1583 301 -1575
rect -1632 -1603 -1580 -1589
tri 146 -1604 167 -1583 ne
rect 167 -1604 301 -1583
rect -298 -1610 -168 -1604
rect -298 -1620 -286 -1610
tri -1483 -1644 -1459 -1620 se
rect -1459 -1644 -286 -1620
rect -252 -1644 -214 -1610
rect -180 -1644 -168 -1610
tri -1486 -1647 -1483 -1644 se
rect -1483 -1647 -168 -1644
rect -1632 -1661 -1580 -1655
tri -1500 -1661 -1486 -1647 se
rect -1486 -1650 -168 -1647
rect -79 -1610 51 -1604
tri 167 -1608 171 -1604 ne
rect -79 -1644 -67 -1610
rect -33 -1644 5 -1610
rect 39 -1644 51 -1610
rect -79 -1650 51 -1644
rect 171 -1613 301 -1604
rect 171 -1647 183 -1613
rect 217 -1647 255 -1613
rect 289 -1647 301 -1613
rect -1486 -1661 -1444 -1650
tri -1444 -1661 -1433 -1650 nw
tri -1503 -1664 -1500 -1661 se
rect -1500 -1664 -1447 -1661
tri -1447 -1664 -1444 -1661 nw
tri -1515 -1676 -1503 -1664 se
rect -1503 -1676 -1459 -1664
tri -1459 -1676 -1447 -1664 nw
tri -1525 -1686 -1515 -1676 se
rect -1515 -1686 -1469 -1676
tri -1469 -1686 -1459 -1676 nw
rect -79 -1680 -32 -1650
rect 171 -1653 301 -1647
rect 1278 -1669 1284 -1617
rect 1336 -1669 1350 -1617
rect 1402 -1669 1408 -1617
rect -1335 -1686 -32 -1680
tri -1531 -1692 -1525 -1686 se
rect -1525 -1692 -1503 -1686
rect -2157 -1720 -1503 -1692
tri -1503 -1720 -1469 -1686 nw
rect -1335 -1720 -1323 -1686
rect -1289 -1720 -1251 -1686
rect -1217 -1720 -32 -1686
rect -2157 -1722 -1505 -1720
tri -1505 -1722 -1503 -1720 nw
rect -1335 -1726 -32 -1720
rect -2197 -1766 572 -1754
rect -2197 -1800 -1802 -1766
rect -1768 -1800 -899 -1766
rect -865 -1800 -434 -1766
rect -400 -1800 -318 -1766
rect -284 -1800 34 -1766
rect 68 -1800 153 -1766
rect 187 -1800 505 -1766
rect 539 -1800 572 -1766
rect 2316 -1775 2354 -1191
rect 3760 -1202 4565 -1153
rect 4851 -1066 4903 -1060
rect 6587 -1072 6639 -1066
rect 4851 -1130 4903 -1118
rect 3760 -1777 3812 -1202
tri 3812 -1238 3848 -1202 nw
rect 4690 -1208 4696 -1156
rect 4748 -1208 4762 -1156
rect 4814 -1208 4820 -1156
rect 4627 -1360 4633 -1308
rect 4685 -1360 4699 -1308
rect 4751 -1360 4757 -1308
rect 4544 -1516 4550 -1464
rect 4602 -1516 4621 -1464
rect 4673 -1516 4679 -1464
rect 4550 -1672 4556 -1620
rect 4608 -1672 4626 -1620
rect 4678 -1672 4684 -1620
rect -2197 -1838 572 -1800
rect -2197 -1872 -1802 -1838
rect -1768 -1872 -899 -1838
rect -865 -1872 -434 -1838
rect -400 -1872 -318 -1838
rect -284 -1872 34 -1838
rect 68 -1872 153 -1838
rect 187 -1872 505 -1838
rect 539 -1872 572 -1838
rect -2197 -1936 572 -1872
rect -2197 -1970 -2185 -1936
rect -2151 -1970 -2111 -1936
rect -2077 -1970 -2037 -1936
rect -2003 -1970 -1963 -1936
rect -1929 -1970 -1889 -1936
rect -1855 -1970 -1815 -1936
rect -1781 -1970 -1741 -1936
rect -1707 -1970 -1667 -1936
rect -1633 -1970 -1593 -1936
rect -1559 -1970 -1519 -1936
rect -1485 -1970 -1445 -1936
rect -1411 -1970 -1372 -1936
rect -1338 -1970 -1299 -1936
rect -1265 -1970 -1226 -1936
rect -1192 -1970 -1153 -1936
rect -1119 -1970 -1080 -1936
rect -1046 -1970 -1007 -1936
rect -973 -1970 -934 -1936
rect -900 -1970 -861 -1936
rect -827 -1970 -788 -1936
rect -754 -1970 -715 -1936
rect -681 -1970 -642 -1936
rect -608 -1970 -569 -1936
rect -535 -1970 -496 -1936
rect -462 -1970 -423 -1936
rect -389 -1970 -350 -1936
rect -316 -1970 -277 -1936
rect -243 -1970 -204 -1936
rect -170 -1970 -131 -1936
rect -97 -1970 -58 -1936
rect -24 -1970 15 -1936
rect 49 -1970 88 -1936
rect 122 -1970 161 -1936
rect 195 -1970 234 -1936
rect 268 -1970 307 -1936
rect 341 -1970 380 -1936
rect 414 -1970 453 -1936
rect 487 -1970 526 -1936
rect 560 -1970 572 -1936
rect -2197 -1976 572 -1970
rect 4723 -2054 4757 -1360
rect 4786 -1981 4820 -1208
rect 4851 -1621 4903 -1182
rect 4851 -1685 4903 -1673
rect 4851 -1743 4903 -1737
rect 4786 -2015 4968 -1981
rect 4723 -2088 4967 -2054
rect 1148 -2306 1403 -2300
rect 1200 -2358 1403 -2306
rect 1148 -2382 1403 -2358
rect 1200 -2434 1403 -2382
rect 1148 -2440 1403 -2434
rect 1357 -2698 1403 -2440
rect 1706 -2541 1758 -2535
rect 1706 -2607 1758 -2593
rect 1706 -2665 1758 -2659
rect 1357 -2704 1667 -2698
rect 1357 -2738 1549 -2704
rect 1583 -2738 1621 -2704
rect 1655 -2738 1667 -2704
rect 1357 -2744 1667 -2738
rect 1505 -3987 1633 -3132
tri 1633 -3189 1690 -3132 nw
rect 1505 -4039 1511 -3987
rect 1563 -4039 1575 -3987
rect 1627 -4039 1633 -3987
rect 1505 -4041 1633 -4039
<< via1 >>
rect -398 938 -346 990
rect -334 938 -282 990
rect 186 921 238 973
rect 250 921 302 973
rect 1333 744 1385 796
rect -2653 676 -2601 728
rect -2589 676 -2537 728
rect -1807 685 -1755 737
rect -1743 685 -1691 737
rect 1333 680 1385 732
rect 1421 795 1473 801
rect 1421 761 1430 795
rect 1430 761 1464 795
rect 1464 761 1473 795
rect 1421 749 1473 761
rect 1421 723 1473 735
rect 1421 689 1430 723
rect 1430 689 1464 723
rect 1464 689 1473 723
rect 1421 683 1473 689
rect 1575 795 1627 801
rect 1575 761 1584 795
rect 1584 761 1618 795
rect 1618 761 1627 795
rect 1575 749 1627 761
rect 1575 723 1627 735
rect 1575 689 1584 723
rect 1584 689 1618 723
rect 1618 689 1627 723
rect 1575 683 1627 689
rect 1727 795 1779 801
rect 1727 761 1736 795
rect 1736 761 1770 795
rect 1770 761 1779 795
rect 1727 749 1779 761
rect 1727 723 1779 735
rect 1727 689 1736 723
rect 1736 689 1770 723
rect 1770 689 1779 723
rect 1727 683 1779 689
rect 2669 795 2721 801
rect 2669 761 2678 795
rect 2678 761 2712 795
rect 2712 761 2721 795
rect 2669 749 2721 761
rect 2669 723 2721 735
rect 2669 689 2678 723
rect 2678 689 2712 723
rect 2712 689 2721 723
rect 2669 683 2721 689
rect 2815 761 2824 785
rect 2824 761 2858 785
rect 2858 761 2867 785
rect 2815 733 2867 761
rect 2815 689 2824 719
rect 2824 689 2858 719
rect 2858 689 2867 719
rect 2815 667 2867 689
rect 2942 738 2978 740
rect 2978 738 2994 740
rect 3008 738 3012 740
rect 3012 738 3060 740
rect 2942 700 2994 738
rect 3008 700 3060 738
rect 2942 688 2978 700
rect 2978 688 2994 700
rect 3008 688 3012 700
rect 3012 688 3060 700
rect -1654 549 -1602 561
rect -1654 515 -1621 549
rect -1621 515 -1602 549
rect -1654 509 -1602 515
rect -1590 549 -1538 561
rect -1590 515 -1583 549
rect -1583 515 -1549 549
rect -1549 515 -1538 549
rect -1590 509 -1538 515
rect -1382 471 -1330 523
rect -1382 435 -1353 459
rect -1353 435 -1330 459
rect -1654 369 -1602 421
rect -1590 369 -1538 421
rect -1382 407 -1330 435
rect -796 507 -744 559
rect -119 648 -67 654
rect -119 614 -113 648
rect -113 614 -79 648
rect -79 614 -67 648
rect -119 602 -67 614
rect -119 576 -67 590
rect -796 443 -744 495
rect -403 548 -351 559
rect -403 514 -397 548
rect -397 514 -363 548
rect -363 514 -351 548
rect -403 507 -351 514
rect -339 548 -287 559
rect -339 514 -320 548
rect -320 514 -287 548
rect -119 542 -113 576
rect -113 542 -79 576
rect -79 542 -67 576
rect 166 577 218 629
rect 269 606 321 658
rect 333 606 385 658
rect -119 538 -67 542
rect 48 562 100 568
rect -339 507 -287 514
rect 48 528 60 562
rect 60 528 94 562
rect 94 528 100 562
rect 48 516 100 528
rect 4432 597 4484 649
rect 4498 597 4550 649
rect 166 550 218 565
rect 166 516 175 550
rect 175 516 209 550
rect 209 516 218 550
rect 166 513 218 516
rect 266 562 318 568
rect 266 528 293 562
rect 293 528 318 562
rect 266 516 318 528
rect 48 489 100 504
rect 48 455 60 489
rect 60 455 94 489
rect 94 455 100 489
rect 48 452 100 455
rect 266 489 318 504
rect 266 455 293 489
rect 293 455 318 489
rect 266 452 318 455
rect 1234 470 1286 522
rect 1234 406 1286 458
rect -790 293 -738 345
rect -726 293 -674 345
rect -566 293 -514 345
rect -502 293 -450 345
rect 2973 422 3025 474
rect -324 226 -272 278
rect -260 226 -208 278
rect -28 291 24 343
rect 36 291 88 343
rect 1076 316 1128 368
rect 2973 356 3025 408
rect 4432 407 4484 459
rect 4498 407 4550 459
rect 839 267 891 279
rect 839 233 849 267
rect 849 233 883 267
rect 883 233 891 267
rect 839 227 891 233
rect 903 227 955 279
rect 1076 252 1128 304
rect 2505 264 2557 316
rect 2505 200 2557 252
rect -790 165 -738 187
rect -790 135 -763 165
rect -763 135 -738 165
rect -725 135 -673 187
rect -660 135 -608 187
rect -595 135 -543 187
rect -530 135 -478 187
rect -465 135 -413 187
rect -400 135 -348 187
rect -335 135 -283 187
rect -270 135 -218 187
rect -790 90 -738 123
rect -790 71 -758 90
rect -758 71 -738 90
rect -725 90 -673 123
rect -725 71 -719 90
rect -719 71 -685 90
rect -685 71 -673 90
rect -660 90 -608 123
rect -660 71 -646 90
rect -646 71 -612 90
rect -612 71 -608 90
rect -595 90 -543 123
rect -530 90 -478 123
rect -465 90 -413 123
rect -400 90 -348 123
rect -335 90 -283 123
rect -270 90 -218 123
rect -595 71 -573 90
rect -573 71 -543 90
rect -530 71 -500 90
rect -500 71 -478 90
rect -465 71 -427 90
rect -427 71 -413 90
rect -400 71 -393 90
rect -393 71 -354 90
rect -354 71 -348 90
rect -335 71 -320 90
rect -320 71 -283 90
rect -270 71 -247 90
rect -247 71 -218 90
rect -790 56 -758 59
rect -758 56 -738 59
rect -790 7 -738 56
rect -725 56 -719 59
rect -719 56 -685 59
rect -685 56 -673 59
rect -725 7 -673 56
rect -660 56 -646 59
rect -646 56 -612 59
rect -612 56 -608 59
rect -660 7 -608 56
rect -595 56 -573 59
rect -573 56 -543 59
rect -530 56 -500 59
rect -500 56 -478 59
rect -465 56 -427 59
rect -427 56 -413 59
rect -400 56 -393 59
rect -393 56 -354 59
rect -354 56 -348 59
rect -335 56 -320 59
rect -320 56 -283 59
rect -270 56 -247 59
rect -247 56 -218 59
rect -595 7 -543 56
rect -530 7 -478 56
rect -465 7 -413 56
rect -400 7 -348 56
rect -335 7 -283 56
rect -270 7 -218 56
rect -790 -57 -738 -5
rect -725 -57 -673 -5
rect -660 -57 -608 -5
rect -595 -57 -543 -5
rect -530 -57 -478 -5
rect -465 -57 -413 -5
rect -400 -57 -348 -5
rect -335 -57 -283 -5
rect -270 -57 -218 -5
rect -1246 -143 -1194 -91
rect -1182 -143 -1130 -91
rect 186 -103 238 -97
rect 186 -137 203 -103
rect 203 -137 238 -103
rect 186 -149 238 -137
rect -2057 -167 -2005 -161
rect -2057 -201 -2048 -167
rect -2048 -201 -2014 -167
rect -2014 -201 -2005 -167
rect 186 -175 238 -161
rect -2057 -213 -2005 -201
rect -2057 -239 -2005 -225
rect -2057 -273 -2048 -239
rect -2048 -273 -2014 -239
rect -2014 -273 -2005 -239
rect -2057 -277 -2005 -273
rect -1953 -242 -1901 -190
rect -1249 -234 -1197 -182
rect -1185 -234 -1133 -182
rect -391 -234 -339 -182
rect -327 -234 -275 -182
rect -1953 -306 -1901 -254
rect -2419 -385 -2367 -333
rect -2355 -346 -2303 -333
rect -2355 -380 -2338 -346
rect -2338 -380 -2304 -346
rect -2304 -380 -2303 -346
rect -2355 -385 -2303 -380
rect -2238 -335 -2186 -329
rect -2238 -369 -2232 -335
rect -2232 -369 -2198 -335
rect -2198 -369 -2186 -335
rect -2238 -381 -2186 -369
rect -2174 -335 -2122 -329
rect -2174 -369 -2160 -335
rect -2160 -369 -2126 -335
rect -2126 -369 -2122 -335
rect -2174 -381 -2122 -369
rect -1776 -322 -1724 -270
rect -1776 -346 -1724 -334
rect -1776 -380 -1767 -346
rect -1767 -380 -1733 -346
rect -1733 -380 -1724 -346
rect -1776 -386 -1724 -380
rect -1663 -322 -1611 -270
rect -1478 -274 -1426 -268
rect -1478 -308 -1469 -274
rect -1469 -308 -1435 -274
rect -1435 -308 -1426 -274
rect -890 -256 -838 -246
rect -890 -290 -884 -256
rect -884 -290 -850 -256
rect -850 -290 -838 -256
rect -890 -298 -838 -290
rect -823 -256 -771 -246
rect -823 -290 -811 -256
rect -811 -290 -777 -256
rect -777 -290 -771 -256
rect -823 -298 -771 -290
rect -1478 -320 -1426 -308
rect -1663 -335 -1611 -334
rect -1663 -369 -1651 -335
rect -1651 -369 -1617 -335
rect -1617 -369 -1611 -335
rect -1663 -386 -1611 -369
rect -721 -303 -669 -251
rect -191 -254 -139 -202
rect -1478 -346 -1426 -334
rect -1478 -380 -1469 -346
rect -1469 -380 -1435 -346
rect -1435 -380 -1426 -346
rect -721 -335 -669 -317
rect -1478 -386 -1426 -380
rect -953 -391 -901 -339
rect -889 -347 -837 -339
rect -889 -381 -857 -347
rect -857 -381 -837 -347
rect -889 -391 -837 -381
rect -721 -369 -715 -335
rect -715 -369 -681 -335
rect -681 -369 -669 -335
rect -624 -314 -572 -293
rect -560 -314 -508 -293
rect -624 -345 -592 -314
rect -592 -345 -572 -314
rect -560 -345 -558 -314
rect -558 -345 -508 -314
rect -333 -333 -281 -281
rect -191 -318 -139 -266
rect 39 -234 91 -182
rect 186 -209 203 -175
rect 203 -209 238 -175
rect 186 -213 238 -209
rect 659 -143 711 -91
rect 723 -143 775 -91
rect 3138 -76 3190 -24
rect 3202 -76 3254 -24
rect 3152 -156 3204 -104
rect 3217 -156 3269 -104
rect 3845 -171 3897 -119
rect 39 -298 91 -246
rect 2973 -248 3025 -196
rect 3152 -242 3204 -190
rect 3217 -242 3269 -190
rect 3845 -236 3897 -184
rect -333 -357 -281 -345
rect 131 -312 183 -260
rect 195 -312 247 -260
rect 483 -312 535 -260
rect 547 -312 599 -260
rect 729 -314 781 -262
rect -333 -391 -321 -357
rect -321 -391 -287 -357
rect -287 -391 -281 -357
rect -333 -397 -281 -391
rect 729 -350 781 -326
rect 825 -272 877 -268
rect 825 -306 834 -272
rect 834 -306 868 -272
rect 868 -306 877 -272
rect 825 -320 877 -306
rect 825 -344 877 -332
rect 729 -378 744 -350
rect 744 -378 778 -350
rect 778 -378 781 -350
rect 825 -378 834 -344
rect 834 -378 868 -344
rect 868 -378 877 -344
rect 825 -384 877 -378
rect 909 -320 961 -268
rect 909 -384 961 -332
rect 1885 -311 1937 -259
rect 2973 -314 3025 -262
rect 1139 -392 1191 -340
rect 1885 -375 1937 -323
rect 3268 -332 3320 -280
rect 3609 -332 3661 -280
rect 3268 -396 3320 -344
rect 3609 -396 3661 -344
rect 6433 -293 6485 -241
rect 6433 -357 6485 -305
rect 1139 -456 1191 -404
rect -2238 -530 -2186 -478
rect -2174 -530 -2122 -478
rect -1657 -597 -1605 -545
rect -1593 -597 -1541 -545
rect -1241 -597 -1189 -545
rect -1177 -597 -1125 -545
rect -910 -591 -858 -539
rect -846 -591 -794 -539
rect -221 -545 -169 -493
rect -157 -545 -105 -493
rect 1136 -549 1188 -497
rect 755 -603 807 -551
rect 819 -603 871 -551
rect 1136 -613 1188 -561
rect 3183 -492 3235 -440
rect 3609 -500 3661 -448
rect 3183 -556 3235 -504
rect 3609 -564 3661 -512
rect 3693 -580 3745 -528
rect 3693 -644 3745 -592
rect 6119 -798 6171 -746
rect 6183 -798 6235 -746
rect 6431 -768 6483 -716
rect -2565 -868 -2513 -816
rect -2501 -868 -2449 -816
rect -2651 -1036 -2599 -984
rect -2587 -1036 -2535 -984
rect 333 -880 385 -828
rect 397 -880 449 -828
rect 6431 -832 6483 -780
rect -2407 -958 -2355 -906
rect -2407 -1022 -2355 -970
rect -790 -969 -771 -942
rect -771 -969 -738 -942
rect -725 -969 -698 -942
rect -698 -969 -673 -942
rect -660 -969 -625 -942
rect -625 -969 -608 -942
rect -595 -969 -591 -942
rect -591 -969 -552 -942
rect -552 -969 -543 -942
rect -530 -969 -518 -942
rect -518 -969 -479 -942
rect -479 -969 -478 -942
rect -465 -969 -445 -942
rect -445 -969 -413 -942
rect -400 -969 -372 -942
rect -372 -969 -348 -942
rect -790 -994 -738 -969
rect -725 -994 -673 -969
rect -660 -994 -608 -969
rect -595 -994 -543 -969
rect -530 -994 -478 -969
rect -465 -994 -413 -969
rect -400 -994 -348 -969
rect -335 -969 -333 -942
rect -333 -969 -299 -942
rect -299 -969 -283 -942
rect -335 -994 -283 -969
rect -270 -969 -260 -942
rect -260 -969 -226 -942
rect -226 -969 -218 -942
rect 4409 -904 4461 -852
rect 4473 -904 4525 -852
rect -270 -994 -218 -969
rect -790 -1015 -738 -1010
rect -790 -1049 -786 -1015
rect -786 -1049 -752 -1015
rect -752 -1049 -738 -1015
rect -790 -1062 -738 -1049
rect -725 -1062 -673 -1010
rect -660 -1062 -608 -1010
rect -595 -1062 -543 -1010
rect -530 -1062 -478 -1010
rect -465 -1015 -413 -1010
rect -465 -1049 -434 -1015
rect -434 -1049 -413 -1015
rect -465 -1062 -413 -1049
rect -400 -1062 -348 -1010
rect -335 -1015 -283 -1010
rect -335 -1049 -318 -1015
rect -318 -1049 -284 -1015
rect -284 -1049 -283 -1015
rect -335 -1062 -283 -1049
rect -270 -1062 -218 -1010
rect -790 -1087 -738 -1078
rect -790 -1121 -786 -1087
rect -786 -1121 -752 -1087
rect -752 -1121 -738 -1087
rect -790 -1130 -738 -1121
rect -725 -1130 -673 -1078
rect -660 -1130 -608 -1078
rect -595 -1130 -543 -1078
rect -530 -1130 -478 -1078
rect -465 -1087 -413 -1078
rect -465 -1121 -434 -1087
rect -434 -1121 -413 -1087
rect -465 -1130 -413 -1121
rect -400 -1130 -348 -1078
rect -335 -1087 -283 -1078
rect -335 -1121 -318 -1087
rect -318 -1121 -284 -1087
rect -284 -1121 -283 -1087
rect -335 -1130 -283 -1121
rect -270 -1130 -218 -1078
rect 1148 -1088 1200 -1036
rect 1148 -1164 1200 -1112
rect 1456 -1125 1508 -1073
rect 1520 -1125 1572 -1073
rect 1704 -1082 1756 -1030
rect 1774 -1082 1826 -1030
rect 1844 -1082 1896 -1030
rect 3217 -1059 3269 -1007
rect 3281 -1059 3333 -1007
rect 6587 -1002 6639 -950
rect 333 -1216 385 -1164
rect 397 -1176 449 -1164
rect 397 -1210 415 -1176
rect 415 -1210 449 -1176
rect 397 -1216 449 -1210
rect 1284 -1166 1336 -1156
rect 1284 -1200 1290 -1166
rect 1290 -1200 1324 -1166
rect 1324 -1200 1336 -1166
rect 1284 -1208 1336 -1200
rect 1357 -1166 1409 -1156
rect 1357 -1200 1362 -1166
rect 1362 -1200 1396 -1166
rect 1396 -1200 1409 -1166
rect 1357 -1208 1409 -1200
rect -2034 -1289 -1982 -1237
rect -1944 -1289 -1892 -1237
rect -2034 -1337 -1982 -1328
rect -1944 -1337 -1892 -1328
rect -2034 -1371 -2008 -1337
rect -2008 -1371 -1982 -1337
rect -1944 -1371 -1936 -1337
rect -1936 -1371 -1902 -1337
rect -1902 -1371 -1892 -1337
rect -2034 -1380 -1982 -1371
rect -1944 -1380 -1892 -1371
rect 1284 -1321 1336 -1312
rect 1284 -1355 1290 -1321
rect 1290 -1355 1324 -1321
rect 1324 -1355 1336 -1321
rect 1284 -1364 1336 -1355
rect 1350 -1321 1402 -1312
rect 1350 -1355 1362 -1321
rect 1362 -1355 1396 -1321
rect 1396 -1355 1402 -1321
rect 1350 -1364 1402 -1355
rect -2481 -1564 -2429 -1512
rect -2417 -1564 -2365 -1512
rect 1284 -1471 1336 -1462
rect 1284 -1505 1290 -1471
rect 1290 -1505 1324 -1471
rect 1324 -1505 1336 -1471
rect 1284 -1514 1336 -1505
rect 1350 -1471 1402 -1462
rect 1350 -1505 1362 -1471
rect 1362 -1505 1396 -1471
rect 1396 -1505 1402 -1471
rect 1350 -1514 1402 -1505
rect -1864 -1539 -1812 -1535
rect -1864 -1573 -1855 -1539
rect -1855 -1573 -1821 -1539
rect -1821 -1573 -1812 -1539
rect -1864 -1587 -1812 -1573
rect -1864 -1611 -1812 -1599
rect -1864 -1645 -1855 -1611
rect -1855 -1645 -1821 -1611
rect -1821 -1645 -1812 -1611
rect -1864 -1651 -1812 -1645
rect -1739 -1543 -1687 -1535
rect -1739 -1577 -1725 -1543
rect -1725 -1577 -1691 -1543
rect -1691 -1577 -1687 -1543
rect -1739 -1587 -1687 -1577
rect -1739 -1615 -1687 -1599
rect -1739 -1649 -1725 -1615
rect -1725 -1649 -1691 -1615
rect -1691 -1649 -1687 -1615
rect -1739 -1651 -1687 -1649
rect -1632 -1543 -1580 -1537
rect -1632 -1577 -1626 -1543
rect -1626 -1577 -1592 -1543
rect -1592 -1577 -1580 -1543
rect -1632 -1589 -1580 -1577
rect -1632 -1615 -1580 -1603
rect -1632 -1649 -1626 -1615
rect -1626 -1649 -1592 -1615
rect -1592 -1649 -1580 -1615
rect -1632 -1655 -1580 -1649
rect 1284 -1627 1336 -1617
rect 1284 -1661 1290 -1627
rect 1290 -1661 1324 -1627
rect 1324 -1661 1336 -1627
rect 1284 -1669 1336 -1661
rect 1350 -1627 1402 -1617
rect 1350 -1661 1362 -1627
rect 1362 -1661 1396 -1627
rect 1396 -1661 1402 -1627
rect 1350 -1669 1402 -1661
rect 4851 -1118 4903 -1066
rect 6587 -1066 6639 -1014
rect 4696 -1164 4748 -1156
rect 4696 -1198 4702 -1164
rect 4702 -1198 4736 -1164
rect 4736 -1198 4748 -1164
rect 4696 -1208 4748 -1198
rect 4762 -1164 4814 -1156
rect 4762 -1198 4774 -1164
rect 4774 -1198 4808 -1164
rect 4808 -1198 4814 -1164
rect 4762 -1208 4814 -1198
rect 4633 -1320 4685 -1308
rect 4633 -1354 4639 -1320
rect 4639 -1354 4673 -1320
rect 4673 -1354 4685 -1320
rect 4633 -1360 4685 -1354
rect 4699 -1320 4751 -1308
rect 4699 -1354 4711 -1320
rect 4711 -1354 4745 -1320
rect 4745 -1354 4751 -1320
rect 4699 -1360 4751 -1354
rect 4550 -1473 4602 -1464
rect 4550 -1507 4556 -1473
rect 4556 -1507 4590 -1473
rect 4590 -1507 4602 -1473
rect 4550 -1516 4602 -1507
rect 4621 -1473 4673 -1464
rect 4621 -1507 4628 -1473
rect 4628 -1507 4662 -1473
rect 4662 -1507 4673 -1473
rect 4621 -1516 4673 -1507
rect 4556 -1630 4608 -1620
rect 4556 -1664 4562 -1630
rect 4562 -1664 4596 -1630
rect 4596 -1664 4608 -1630
rect 4556 -1672 4608 -1664
rect 4626 -1630 4678 -1620
rect 4626 -1664 4634 -1630
rect 4634 -1664 4668 -1630
rect 4668 -1664 4678 -1630
rect 4626 -1672 4678 -1664
rect 4851 -1182 4903 -1130
rect 4851 -1673 4903 -1621
rect 4851 -1737 4903 -1685
rect 1148 -2358 1200 -2306
rect 1148 -2434 1200 -2382
rect 1706 -2547 1758 -2541
rect 1706 -2581 1715 -2547
rect 1715 -2581 1749 -2547
rect 1749 -2581 1758 -2547
rect 1706 -2593 1758 -2581
rect 1706 -2619 1758 -2607
rect 1706 -2653 1715 -2619
rect 1715 -2653 1749 -2619
rect 1749 -2653 1758 -2619
rect 1706 -2659 1758 -2653
rect 1511 -4039 1563 -3987
rect 1575 -4039 1627 -3987
<< metal2 >>
rect -2619 759 -2294 811
rect -2238 768 -1600 809
rect -2659 676 -2653 728
rect -2601 676 -2589 728
rect -2537 676 -2531 728
rect -1813 685 -1807 737
rect -1755 685 -1743 737
rect -1691 728 -1685 737
rect -1741 648 -1685 672
rect -2168 604 -2112 613
rect -1741 583 -1685 592
rect -1640 561 -1600 768
rect -2168 517 -2112 548
rect -1660 509 -1654 561
rect -1602 509 -1590 561
rect -1538 509 -1532 561
rect -1382 523 -1330 529
rect -2168 421 -2112 461
rect -1382 459 -1330 471
rect -2168 369 -1654 421
rect -1602 369 -1590 421
rect -1538 369 -1532 421
rect -1330 407 -1200 458
rect -1382 401 -1200 407
rect -2353 88 -1821 144
rect -1765 88 -1741 144
rect -1685 88 -1676 144
rect -2353 -333 -2297 88
rect -2057 -103 -1750 -47
rect -1694 -103 -1670 -47
rect -1614 -103 -1605 -47
rect -1252 -91 -1200 401
rect -2057 -161 -2005 -103
rect -1867 -143 -1298 -137
tri -1298 -143 -1292 -137 sw
rect -1252 -143 -1246 -91
rect -1194 -143 -1182 -91
rect -1130 -143 -1124 -91
rect -1867 -146 -1292 -143
rect -2057 -225 -2005 -213
rect -2057 -283 -2005 -277
rect -1953 -190 -1901 -184
rect -1953 -254 -1901 -242
rect -1811 -149 -1292 -146
tri -1292 -149 -1286 -143 sw
rect -1811 -156 -1286 -149
tri -1286 -156 -1279 -149 sw
rect -1811 -161 -1279 -156
tri -1279 -161 -1274 -156 sw
rect -1811 -169 -1274 -161
tri -1340 -182 -1327 -169 ne
rect -1327 -182 -1274 -169
tri -1274 -182 -1253 -161 sw
rect -949 -169 -917 934
rect -872 261 -840 1059
rect 48 1043 1434 1059
tri 1434 1043 1450 1059 sw
rect 48 1018 3309 1043
rect -404 938 -398 990
rect -346 938 -334 990
rect -282 938 -276 990
rect -796 559 -744 565
rect -404 559 -370 938
rect -119 654 -67 660
rect -119 590 -67 602
rect -409 507 -403 559
rect -351 507 -339 559
rect -287 507 -281 559
rect 48 568 100 1018
tri 100 986 132 1018 nw
tri 1396 1002 1412 1018 ne
rect 1412 1002 3309 1018
tri 3276 986 3292 1002 ne
rect 3292 993 3309 1002
tri 3309 993 3359 1043 sw
rect 3292 986 3359 993
tri 3292 973 3305 986 ne
rect 3305 973 3359 986
rect 180 921 186 973
rect 238 921 250 973
rect 302 921 308 973
tri 3305 969 3309 973 ne
rect 3309 969 3359 973
tri 3309 964 3314 969 ne
rect 3314 964 3359 969
rect 263 658 308 921
tri 1726 911 1779 964 se
rect 1779 928 3257 964
rect 1726 807 1779 911
tri 1779 872 1835 928 nw
tri 3224 895 3257 928 ne
tri 3257 923 3298 964 sw
tri 3314 923 3355 964 ne
rect 3355 923 3359 964
rect 3257 919 3298 923
tri 3298 919 3302 923 sw
tri 3355 919 3359 923 ne
tri 3359 919 3433 993 sw
rect 3257 895 3302 919
tri 3257 880 3272 895 ne
rect 3272 880 3302 895
tri 2707 872 2715 880 se
rect 2715 872 3213 880
rect 1333 796 1385 802
rect 1333 732 1385 744
rect -67 538 12 564
rect -119 532 12 538
rect -796 495 -744 507
rect -796 345 -744 443
rect -20 416 12 532
rect 48 504 100 516
rect 48 446 100 452
rect 166 629 218 635
rect 263 606 269 658
rect 321 606 333 658
rect 385 606 391 658
rect 166 565 218 577
rect 166 452 218 513
rect 266 568 331 574
rect 318 516 331 568
rect 1333 538 1385 680
rect 1421 801 1473 807
rect 1421 735 1473 749
rect 1421 602 1473 683
rect 1575 801 1627 807
rect 1575 735 1627 749
rect 1575 642 1627 683
rect 1727 801 1779 807
rect 1727 735 1779 749
rect 1727 677 1779 683
tri 2669 834 2707 872 se
rect 2707 854 3213 872
tri 3213 854 3239 880 sw
tri 3272 854 3298 880 ne
rect 3298 862 3302 880
tri 3302 862 3359 919 sw
tri 3359 862 3416 919 ne
rect 3416 862 3433 919
rect 3298 854 3359 862
rect 2707 844 3239 854
rect 2707 834 2721 844
rect 2669 801 2721 834
tri 2721 794 2771 844 nw
tri 3180 815 3209 844 ne
rect 3209 817 3239 844
tri 3239 817 3276 854 sw
tri 3298 817 3335 854 ne
rect 3335 845 3359 854
tri 3359 845 3376 862 sw
tri 3416 845 3433 862 ne
tri 3433 845 3507 919 sw
rect 3335 817 3376 845
rect 3209 815 3276 817
tri 2818 794 2839 815 se
rect 2839 811 3150 815
tri 3150 811 3154 815 sw
tri 3209 811 3213 815 ne
rect 3213 811 3276 815
rect 2839 794 3154 811
rect 2669 735 2721 749
rect 2669 677 2721 683
tri 2815 791 2818 794 se
rect 2818 791 3154 794
rect 2815 785 3154 791
rect 2867 779 3154 785
tri 2867 758 2888 779 nw
tri 3112 758 3133 779 ne
rect 3133 777 3154 779
tri 3154 777 3188 811 sw
tri 3213 777 3247 811 ne
rect 3247 795 3276 811
tri 3276 795 3298 817 sw
tri 3335 795 3357 817 ne
rect 3357 795 3376 817
rect 3247 777 3298 795
rect 3133 758 3188 777
tri 3133 741 3150 758 ne
rect 3150 752 3188 758
tri 3188 752 3213 777 sw
tri 3247 752 3272 777 ne
rect 3272 752 3298 777
rect 3150 741 3213 752
tri 3150 740 3151 741 ne
rect 3151 740 3213 741
rect 2815 719 2867 733
rect 2936 688 2942 740
rect 2994 688 3008 740
rect 3060 688 3066 740
tri 3151 703 3188 740 ne
rect 3188 703 3213 740
tri 3213 703 3262 752 sw
tri 3272 748 3276 752 ne
rect 3276 748 3298 752
tri 3298 748 3345 795 sw
tri 3357 785 3367 795 ne
rect 3367 788 3376 795
tri 3376 788 3433 845 sw
tri 3433 788 3490 845 ne
rect 3490 788 3507 845
rect 3367 785 3433 788
tri 3367 748 3404 785 ne
rect 3404 771 3433 785
tri 3433 771 3450 788 sw
tri 3490 771 3507 788 ne
tri 3507 771 3581 845 sw
rect 3404 748 3450 771
tri 3276 703 3321 748 ne
rect 3321 726 3345 748
tri 3345 726 3367 748 sw
tri 3404 726 3426 748 ne
rect 3426 726 3450 748
rect 3321 703 3367 726
tri 3188 688 3203 703 ne
rect 3203 689 3262 703
tri 3262 689 3276 703 sw
tri 3321 689 3335 703 ne
rect 3335 689 3367 703
rect 3203 688 3276 689
tri 2814 649 2815 650 se
rect 2815 649 2867 667
tri 1627 642 1634 649 sw
tri 2807 642 2814 649 se
rect 2814 642 2867 649
rect 1575 628 2867 642
rect 1575 627 2841 628
tri 1575 624 1578 627 ne
rect 1578 624 2841 627
tri 1473 602 1495 624 sw
tri 1578 602 1600 624 ne
rect 1600 602 2841 624
tri 2841 602 2867 628 nw
tri 2945 602 2969 626 se
rect 2969 604 3021 688
tri 3203 649 3242 688 ne
rect 3242 679 3276 688
tri 3276 679 3286 689 sw
tri 3335 679 3345 689 ne
rect 3345 679 3367 689
tri 3367 679 3414 726 sw
tri 3426 716 3436 726 ne
rect 3436 716 3450 726
tri 3450 716 3505 771 sw
tri 3507 716 3562 771 ne
rect 3562 716 3581 771
tri 3436 679 3473 716 ne
rect 3473 714 3505 716
tri 3505 714 3507 716 sw
tri 3562 714 3564 716 ne
rect 3564 714 3581 716
rect 3473 697 3507 714
tri 3507 697 3524 714 sw
tri 3564 697 3581 714 ne
tri 3581 697 3655 771 sw
rect 3473 679 3524 697
rect 3242 649 3286 679
tri 3286 649 3316 679 sw
tri 3345 649 3375 679 ne
rect 3375 657 3414 679
tri 3414 657 3436 679 sw
tri 3473 657 3495 679 ne
rect 3495 657 3524 679
rect 3375 649 3436 657
tri 3436 649 3444 657 sw
tri 3495 649 3503 657 ne
rect 3503 649 3524 657
tri 3524 649 3572 697 sw
tri 3581 669 3609 697 ne
tri 3242 629 3262 649 ne
rect 3262 629 3316 649
tri 3316 629 3336 649 sw
tri 3375 629 3395 649 ne
rect 3395 629 3444 649
rect 2969 602 3014 604
tri 1421 597 1426 602 ne
rect 1426 597 1495 602
tri 1495 597 1500 602 sw
tri 2940 597 2945 602 se
rect 2945 597 3014 602
tri 3014 597 3021 604 nw
tri 3262 597 3294 629 ne
rect 3294 620 3336 629
tri 3336 620 3345 629 sw
tri 3395 620 3404 629 ne
rect 3404 620 3444 629
rect 3294 610 3345 620
tri 3345 610 3355 620 sw
tri 3404 610 3414 620 ne
rect 3414 610 3444 620
tri 3444 610 3483 649 sw
tri 3503 647 3505 649 ne
rect 3505 647 3572 649
tri 3572 647 3574 649 sw
tri 3505 618 3534 647 ne
rect 3294 597 3355 610
tri 3355 597 3368 610 sw
tri 3414 597 3427 610 ne
rect 3427 597 3483 610
tri 1426 574 1449 597 ne
rect 1449 574 1500 597
tri 1385 538 1421 574 sw
tri 1449 538 1485 574 ne
rect 1485 564 1500 574
tri 1500 564 1533 597 sw
tri 2929 586 2940 597 se
rect 2940 586 3003 597
tri 3003 586 3014 597 nw
tri 3294 586 3305 597 ne
rect 3305 586 3368 597
tri 2907 564 2929 586 se
rect 1485 538 2929 564
rect 1333 532 1421 538
tri 1333 528 1337 532 ne
rect 1337 528 1421 532
rect 266 504 331 516
tri 218 452 238 472 sw
rect 166 448 238 452
tri 166 446 168 448 ne
rect 168 446 238 448
rect 318 452 331 504
rect 266 446 331 452
tri 168 428 186 446 ne
rect -20 384 157 416
rect -796 293 -790 345
rect -738 293 -726 345
rect -674 293 -668 345
tri -578 293 -572 299 se
rect -572 293 -566 345
rect -514 293 -502 345
rect -450 293 -444 345
tri -580 291 -578 293 se
rect -578 291 -526 293
tri -526 291 -524 293 nw
rect -34 291 -28 343
rect 24 291 36 343
rect 88 291 94 343
tri -592 279 -580 291 se
rect -580 279 -538 291
tri -538 279 -526 291 nw
tri -593 278 -592 279 se
rect -592 278 -539 279
tri -539 278 -538 279 nw
tri -610 261 -593 278 se
rect -593 261 -556 278
tri -556 261 -539 278 nw
rect -872 227 -590 261
tri -590 227 -556 261 nw
rect -872 -92 -840 227
rect -330 226 -324 278
rect -272 226 -260 278
rect -208 226 -134 278
rect -796 135 -790 187
rect -738 173 -725 187
rect -673 173 -660 187
rect -608 173 -595 187
rect -543 173 -530 187
rect -478 173 -465 187
rect -413 173 -400 187
rect -348 173 -335 187
rect -283 173 -270 187
rect -729 135 -725 173
rect -543 135 -532 173
rect -476 135 -465 173
rect -283 135 -280 173
rect -218 135 -212 187
rect -796 123 -785 135
rect -729 123 -700 135
rect -644 123 -616 135
rect -560 123 -532 135
rect -476 123 -448 135
rect -392 123 -364 135
rect -308 123 -280 135
rect -224 123 -212 135
rect -796 71 -790 123
rect -729 117 -725 123
rect -543 117 -532 123
rect -476 117 -465 123
rect -283 117 -280 123
rect -738 93 -725 117
rect -673 93 -660 117
rect -608 93 -595 117
rect -543 93 -530 117
rect -478 93 -465 117
rect -413 93 -400 117
rect -348 93 -335 117
rect -283 93 -270 117
rect -729 71 -725 93
rect -543 71 -532 93
rect -476 71 -465 93
rect -283 71 -280 93
rect -218 71 -212 123
rect -796 59 -785 71
rect -729 59 -700 71
rect -644 59 -616 71
rect -560 59 -532 71
rect -476 59 -448 71
rect -392 59 -364 71
rect -308 59 -280 71
rect -224 59 -212 71
rect -796 7 -790 59
rect -729 37 -725 59
rect -543 37 -532 59
rect -476 37 -465 59
rect -283 37 -280 59
rect -738 13 -725 37
rect -673 13 -660 37
rect -608 13 -595 37
rect -543 13 -530 37
rect -478 13 -465 37
rect -413 13 -400 37
rect -348 13 -335 37
rect -283 13 -270 37
rect -729 7 -725 13
rect -543 7 -532 13
rect -476 7 -465 13
rect -283 7 -280 13
rect -218 7 -212 59
rect -796 -5 -785 7
rect -729 -5 -700 7
rect -644 -5 -616 7
rect -560 -5 -532 7
rect -476 -5 -448 7
rect -392 -5 -364 7
rect -308 -5 -280 7
rect -224 -5 -212 7
rect -796 -57 -790 -5
rect -729 -43 -725 -5
rect -543 -43 -532 -5
rect -476 -43 -465 -5
rect -283 -43 -280 -5
rect -738 -57 -725 -43
rect -673 -57 -660 -43
rect -608 -57 -595 -43
rect -543 -57 -530 -43
rect -478 -57 -465 -43
rect -413 -57 -400 -43
rect -348 -57 -335 -43
rect -283 -57 -270 -43
rect -218 -57 -212 -5
rect -166 -71 -134 226
rect -872 -124 -428 -92
rect -166 -103 -72 -71
tri -1327 -201 -1308 -182 ne
rect -1308 -201 -1249 -182
rect -1867 -226 -1811 -202
rect -1867 -291 -1811 -282
rect -1776 -233 -1365 -201
tri -1308 -211 -1298 -201 ne
rect -1298 -211 -1249 -201
rect -1776 -270 -1724 -233
rect -2425 -385 -2419 -333
rect -2367 -385 -2355 -333
rect -2303 -385 -2297 -333
rect -2244 -381 -2238 -329
rect -2186 -381 -2174 -329
rect -2122 -381 -2116 -329
rect -2347 -476 -2295 -385
rect -2244 -478 -2116 -381
rect -2244 -530 -2238 -478
rect -2186 -530 -2174 -478
rect -2122 -530 -2116 -478
rect -2589 -868 -2565 -816
rect -2513 -868 -2501 -816
rect -2449 -868 -2443 -816
rect -2407 -906 -2355 -900
rect -2407 -970 -2355 -958
rect -2657 -1036 -2651 -984
rect -2599 -1036 -2587 -984
rect -2535 -1036 -2529 -984
rect -1953 -931 -1901 -306
rect -1776 -334 -1724 -322
rect -1776 -392 -1724 -386
rect -1663 -270 -1611 -264
rect -1663 -334 -1611 -322
rect -1663 -545 -1611 -386
rect -1478 -268 -1426 -262
rect -1478 -334 -1426 -320
rect -1663 -597 -1657 -545
rect -1605 -597 -1593 -545
rect -1541 -597 -1535 -545
tri -1901 -931 -1891 -921 sw
rect -1953 -942 -1891 -931
tri -1891 -942 -1880 -931 sw
rect -1953 -943 -1880 -942
tri -1953 -994 -1902 -943 ne
rect -1902 -994 -1880 -943
tri -1880 -994 -1828 -942 sw
tri -1902 -1002 -1894 -994 ne
rect -1894 -1002 -1828 -994
tri -1828 -1002 -1820 -994 sw
tri -1894 -1005 -1891 -1002 ne
rect -1891 -1005 -1820 -1002
tri -1820 -1005 -1817 -1002 sw
tri -1891 -1007 -1889 -1005 ne
rect -1889 -1007 -1589 -1005
tri -1589 -1007 -1587 -1005 sw
tri -1889 -1010 -1886 -1007 ne
rect -1886 -1010 -1587 -1007
tri -1587 -1010 -1584 -1007 sw
rect -2407 -1028 -2355 -1022
tri -1886 -1028 -1868 -1010 ne
rect -1868 -1028 -1584 -1010
tri -1868 -1036 -1860 -1028 ne
rect -1860 -1034 -1584 -1028
tri -1584 -1034 -1560 -1010 sw
rect -1860 -1036 -1560 -1034
tri -1860 -1057 -1839 -1036 ne
rect -1839 -1057 -1560 -1036
tri -1611 -1062 -1606 -1057 ne
rect -1606 -1062 -1560 -1057
tri -1560 -1062 -1532 -1034 sw
rect -1478 -1044 -1426 -386
rect -1397 -455 -1365 -233
tri -1298 -234 -1275 -211 ne
rect -1275 -234 -1249 -211
rect -1197 -234 -1185 -182
rect -1133 -234 -1127 -182
rect -949 -201 -573 -169
rect -896 -298 -890 -246
rect -838 -298 -823 -246
rect -771 -298 -765 -246
rect -959 -391 -953 -339
rect -901 -391 -889 -339
rect -837 -391 -831 -339
rect -1397 -487 -1058 -455
rect -1247 -597 -1241 -545
rect -1189 -597 -1177 -545
rect -1125 -597 -1119 -545
rect -1156 -770 -1128 -597
rect -1090 -705 -1058 -487
rect -916 -539 -864 -391
rect -793 -437 -765 -298
rect -721 -251 -669 -245
rect -605 -293 -573 -201
rect -721 -317 -669 -303
rect -630 -345 -624 -293
rect -572 -345 -560 -293
rect -508 -345 -502 -293
rect -721 -388 -669 -369
rect -460 -388 -428 -124
rect -397 -234 -391 -182
rect -339 -234 -327 -182
rect -275 -202 -269 -182
rect -191 -202 -139 -196
rect -275 -234 -191 -202
rect -191 -266 -139 -254
rect -721 -420 -428 -388
rect -333 -281 -281 -275
rect -191 -324 -139 -318
rect -333 -345 -281 -333
tri -137 -371 -104 -338 se
rect -104 -352 -72 -103
rect 44 -176 76 291
rect 39 -182 91 -176
rect 39 -246 91 -234
rect 39 -304 91 -298
rect 125 -260 157 384
rect 186 -97 238 446
rect 186 -161 238 -149
rect 186 -219 238 -213
rect 125 -312 131 -260
rect 183 -312 195 -260
rect 247 -312 253 -260
rect -104 -371 -91 -352
tri -91 -371 -72 -352 nw
rect -281 -378 -98 -371
tri -98 -378 -91 -371 nw
rect -281 -384 -104 -378
tri -104 -384 -98 -378 nw
rect -281 -392 -112 -384
tri -112 -392 -104 -384 nw
rect 299 -386 331 446
rect 1234 522 1286 528
tri 1337 480 1385 528 ne
rect 1385 480 1421 528
tri 1421 480 1479 538 sw
tri 1485 528 1495 538 ne
rect 1495 528 2929 538
tri 1495 512 1511 528 ne
rect 1511 512 2929 528
tri 2929 512 3003 586 nw
tri 3305 555 3336 586 ne
rect 3336 555 3368 586
tri 3368 555 3410 597 sw
tri 3427 581 3443 597 ne
tri 3336 531 3360 555 ne
tri 1385 474 1391 480 ne
rect 1391 474 3025 480
rect 1234 458 1286 470
tri 1391 431 1434 474 ne
rect 1434 431 2973 474
tri 628 368 658 398 se
rect 658 370 950 398
rect 658 368 678 370
tri 678 368 680 370 nw
tri 928 368 930 370 ne
rect 930 368 950 370
tri 950 368 980 398 sw
rect 1076 369 1132 378
tri 608 348 628 368 se
rect 628 348 658 368
tri 658 348 678 368 nw
tri 930 348 950 368 ne
rect 950 352 980 368
tri 980 352 996 368 sw
rect 950 348 996 352
tri 577 317 608 348 se
rect 608 317 627 348
tri 627 317 658 348 nw
tri 950 317 981 348 ne
rect 981 317 996 348
rect 577 316 626 317
tri 626 316 627 317 nw
tri 981 316 982 317 ne
rect 982 316 996 317
tri 996 316 1032 352 sw
rect 1234 356 1286 406
rect 2973 408 3025 422
tri 1286 356 1294 364 sw
rect 1234 327 1294 356
tri 1234 316 1245 327 ne
rect 1245 322 1294 327
tri 1294 322 1328 356 sw
rect 2973 350 3025 356
rect 1245 316 2557 322
rect 577 304 614 316
tri 614 304 626 316 nw
tri 982 304 994 316 ne
rect 994 304 1032 316
tri 1032 304 1044 316 sw
rect 1076 304 1132 313
rect 577 -260 605 304
tri 605 295 614 304 nw
tri 994 302 996 304 ne
rect 996 302 1044 304
tri 1044 302 1046 304 sw
tri 996 295 1003 302 ne
rect 1003 295 1046 302
tri 1003 280 1018 295 ne
rect 833 227 839 279
rect 891 227 903 279
rect 955 227 961 279
rect 653 -143 659 -91
rect 711 -143 723 -91
rect 775 -143 781 -91
rect 477 -312 483 -260
rect 535 -312 547 -260
rect 599 -312 605 -260
rect -281 -396 -116 -392
tri -116 -396 -112 -392 nw
rect -281 -397 -123 -396
rect -333 -403 -123 -397
tri -123 -403 -116 -396 nw
rect 103 -418 331 -386
tri -765 -437 -762 -434 sw
rect -793 -446 -762 -437
tri -793 -456 -783 -446 ne
rect -783 -456 -762 -446
tri -762 -456 -743 -437 sw
tri -783 -477 -762 -456 ne
rect -762 -477 -743 -456
tri -743 -477 -722 -456 sw
tri -762 -492 -747 -477 ne
rect -747 -492 -722 -477
tri -722 -492 -707 -477 sw
tri -747 -493 -746 -492 ne
rect -746 -493 -707 -492
tri -707 -493 -706 -492 sw
tri -746 -517 -722 -493 ne
rect -722 -517 -706 -493
tri -706 -517 -682 -493 sw
rect -227 -517 -221 -493
tri -722 -539 -700 -517 ne
rect -700 -539 -221 -517
rect -916 -591 -910 -539
rect -858 -591 -846 -539
rect -794 -591 -788 -539
tri -700 -545 -694 -539 ne
rect -694 -545 -221 -539
rect -169 -545 -157 -493
rect -105 -545 -99 -493
rect 103 -705 135 -418
rect 577 -655 605 -312
rect 729 -262 781 -143
rect 729 -326 781 -314
rect 729 -384 781 -378
rect 825 -268 877 -262
rect 825 -332 877 -320
rect 825 -390 877 -384
rect 909 -268 961 227
rect 1018 44 1046 295
rect 1128 289 1132 304
tri 1245 277 1284 316 ne
rect 1284 277 2505 316
tri 2471 264 2484 277 ne
rect 2484 264 2505 277
tri 2484 252 2496 264 ne
rect 2496 252 2557 264
tri 2496 243 2505 252 ne
rect 1076 224 1132 233
rect 2505 194 2557 200
tri 1046 44 1068 66 sw
tri 1018 12 1050 44 ne
rect 1050 12 3281 44
tri 3267 -2 3281 12 ne
tri 3281 3 3322 44 sw
rect 3281 -2 3322 3
tri 3281 -11 3290 -2 ne
tri 3112 -44 3132 -24 se
rect 3132 -44 3138 -24
rect 909 -332 961 -320
rect 909 -390 961 -384
tri 1015 -62 1033 -44 se
rect 1033 -62 3138 -44
rect 1015 -76 3138 -62
rect 3190 -76 3202 -24
rect 3254 -76 3260 -24
rect 826 -551 877 -390
rect 749 -603 755 -551
rect 807 -603 819 -551
rect 871 -603 877 -551
rect -1090 -737 135 -705
rect 181 -683 605 -655
rect 181 -770 209 -683
rect -1156 -798 209 -770
rect 327 -880 333 -828
rect 385 -880 397 -828
rect 449 -880 455 -828
rect -796 -994 -790 -942
rect -738 -944 -725 -942
rect -673 -944 -660 -942
rect -608 -944 -595 -942
rect -543 -944 -530 -942
rect -478 -944 -465 -942
rect -413 -944 -400 -942
rect -348 -944 -335 -942
rect -283 -944 -270 -942
rect -729 -994 -725 -944
rect -543 -994 -532 -944
rect -476 -994 -465 -944
rect -283 -994 -280 -944
rect -218 -994 -212 -942
rect -796 -1000 -785 -994
rect -729 -1000 -700 -994
rect -644 -1000 -616 -994
rect -560 -1000 -532 -994
rect -476 -1000 -448 -994
rect -392 -1000 -364 -994
rect -308 -1000 -280 -994
rect -224 -1000 -212 -994
rect -796 -1010 -212 -1000
tri -1426 -1044 -1425 -1043 sw
rect -1478 -1047 -1425 -1044
tri -1478 -1062 -1463 -1047 ne
rect -1463 -1062 -1425 -1047
tri -1425 -1062 -1407 -1044 sw
rect -796 -1062 -790 -1010
rect -738 -1062 -725 -1010
rect -673 -1062 -660 -1010
rect -608 -1062 -595 -1010
rect -543 -1062 -530 -1010
rect -478 -1062 -465 -1010
rect -413 -1062 -400 -1010
rect -348 -1062 -335 -1010
rect -283 -1062 -270 -1010
rect -218 -1062 -212 -1010
tri -1606 -1078 -1590 -1062 ne
rect -1590 -1078 -1532 -1062
tri -1532 -1078 -1516 -1062 sw
tri -1463 -1078 -1447 -1062 ne
rect -1447 -1078 -1407 -1062
tri -1407 -1078 -1391 -1062 sw
rect -796 -1072 -212 -1062
rect -796 -1078 -785 -1072
rect -729 -1078 -700 -1072
rect -644 -1078 -616 -1072
rect -560 -1078 -532 -1072
rect -476 -1078 -448 -1072
rect -392 -1078 -364 -1072
rect -308 -1078 -280 -1072
rect -224 -1078 -212 -1072
tri -1590 -1108 -1560 -1078 ne
rect -1560 -1108 -1516 -1078
tri -1516 -1108 -1486 -1078 sw
tri -1447 -1100 -1425 -1078 ne
rect -1425 -1100 -1391 -1078
tri -1391 -1100 -1369 -1078 sw
tri -1425 -1108 -1417 -1100 ne
rect -1417 -1108 -1369 -1100
tri -1560 -1130 -1538 -1108 ne
rect -1538 -1130 -1486 -1108
tri -1486 -1130 -1464 -1108 sw
tri -1417 -1130 -1395 -1108 ne
rect -1395 -1130 -1369 -1108
tri -1369 -1130 -1339 -1100 sw
rect -796 -1130 -790 -1078
rect -729 -1128 -725 -1078
rect -543 -1128 -532 -1078
rect -476 -1128 -465 -1078
rect -283 -1128 -280 -1078
rect -738 -1130 -725 -1128
rect -673 -1130 -660 -1128
rect -608 -1130 -595 -1128
rect -543 -1130 -530 -1128
rect -478 -1130 -465 -1128
rect -413 -1130 -400 -1128
rect -348 -1130 -335 -1128
rect -283 -1130 -270 -1128
rect -218 -1130 -212 -1078
tri -1538 -1164 -1504 -1130 ne
rect -1504 -1156 -1464 -1130
tri -1464 -1156 -1438 -1130 sw
tri -1395 -1156 -1369 -1130 ne
rect -1369 -1156 -1339 -1130
tri -1339 -1156 -1313 -1130 sw
rect -1504 -1164 -1438 -1156
tri -1438 -1164 -1430 -1156 sw
tri -1369 -1164 -1361 -1156 ne
rect -1361 -1164 -1313 -1156
tri -1313 -1164 -1305 -1156 sw
rect 327 -1164 455 -880
tri -1504 -1182 -1486 -1164 ne
rect -1486 -1182 -1430 -1164
tri -1430 -1182 -1412 -1164 sw
tri -1361 -1182 -1343 -1164 ne
rect -1343 -1182 -1305 -1164
tri -1486 -1216 -1452 -1182 ne
rect -1452 -1212 -1412 -1182
tri -1412 -1212 -1382 -1182 sw
tri -1343 -1212 -1313 -1182 ne
rect -1313 -1212 -1305 -1182
tri -1305 -1212 -1257 -1164 sw
rect -1452 -1216 -1382 -1212
tri -1382 -1216 -1378 -1212 sw
tri -1313 -1216 -1309 -1212 ne
rect -1309 -1216 -1257 -1212
tri -1257 -1216 -1253 -1212 sw
rect 327 -1216 333 -1164
rect 385 -1216 397 -1164
rect 449 -1216 455 -1164
tri -1452 -1235 -1433 -1216 ne
rect -1433 -1235 -1378 -1216
rect -2534 -1237 -1886 -1235
rect -2534 -1289 -2034 -1237
rect -1982 -1289 -1944 -1237
rect -1892 -1289 -1886 -1237
tri -1433 -1256 -1412 -1235 ne
rect -1412 -1256 -1378 -1235
tri -1378 -1256 -1338 -1216 sw
tri -1309 -1256 -1269 -1216 ne
rect -1269 -1256 -1253 -1216
rect -2534 -1291 -1886 -1289
tri -1412 -1291 -1377 -1256 ne
rect -1377 -1268 -1338 -1256
tri -1338 -1268 -1326 -1256 sw
tri -1269 -1268 -1257 -1256 ne
rect -1257 -1268 -1253 -1256
tri -1253 -1268 -1201 -1216 sw
tri 988 -1268 1015 -1241 se
rect 1015 -1268 1047 -76
tri 1047 -103 1074 -76 nw
tri 3273 -103 3290 -86 se
rect 3290 -103 3322 -2
tri 3272 -104 3273 -103 se
rect 3273 -104 3322 -103
rect -1377 -1291 -1326 -1268
tri -1377 -1308 -1360 -1291 ne
rect -1360 -1308 -1326 -1291
tri -1326 -1308 -1286 -1268 sw
tri -1257 -1300 -1225 -1268 ne
rect -1225 -1282 1047 -1268
rect -1225 -1300 1029 -1282
tri 1029 -1300 1047 -1282 nw
tri 1075 -122 1093 -104 se
rect 1093 -115 2868 -104
tri 2868 -115 2879 -104 sw
rect 1093 -122 2879 -115
rect 1075 -136 2879 -122
rect 1075 -156 1114 -136
tri 1114 -156 1134 -136 nw
tri 2850 -156 2870 -136 ne
rect 2870 -156 2879 -136
tri 2879 -156 2920 -115 sw
rect 3146 -156 3152 -104
rect 3204 -156 3217 -104
rect 3269 -130 3322 -104
rect 3269 -156 3296 -130
tri 3296 -156 3322 -130 nw
tri 1070 -1308 1075 -1303 se
rect 1075 -1308 1107 -156
tri 1107 -163 1114 -156 nw
tri 2870 -163 2877 -156 ne
rect 2877 -163 2920 -156
tri 2877 -165 2879 -163 ne
rect 2879 -165 2920 -163
tri 2920 -165 2929 -156 sw
tri 2879 -171 2885 -165 ne
rect 2885 -171 2929 -165
tri 2885 -177 2891 -171 ne
rect 1885 -255 1937 -253
rect 1139 -259 1937 -255
rect 1139 -307 1885 -259
rect 1139 -340 1191 -307
rect 1885 -323 1937 -311
rect 1885 -381 1937 -375
rect 1139 -404 1191 -392
rect 2891 -385 2929 -171
rect 2973 -196 3152 -190
rect 3025 -242 3152 -196
rect 3204 -242 3217 -190
rect 3269 -242 3275 -190
rect 2973 -262 3025 -248
rect 2973 -320 3025 -314
rect 3268 -280 3320 -274
rect 3268 -344 3320 -332
tri 2929 -385 2934 -380 sw
rect 2891 -391 2934 -385
tri 2891 -396 2896 -391 ne
rect 2896 -396 2934 -391
tri 2934 -396 2945 -385 sw
tri 2896 -434 2934 -396 ne
rect 2934 -434 2945 -396
tri 2945 -434 2983 -396 sw
tri 2934 -440 2940 -434 ne
rect 2940 -440 3235 -434
rect 1139 -462 1191 -456
tri 2940 -462 2962 -440 ne
rect 2962 -462 3183 -440
tri 2962 -469 2969 -462 ne
rect 2969 -469 3183 -462
rect 1136 -497 1188 -491
rect 1136 -561 1188 -549
rect 3183 -504 3235 -492
rect 3183 -562 3235 -556
rect 1136 -619 1188 -613
rect 1136 -898 1185 -619
tri 1185 -622 1188 -619 nw
tri 1185 -898 1204 -879 sw
rect 1136 -904 1307 -898
tri 1307 -904 1313 -898 sw
rect 1136 -908 1313 -904
tri 1313 -908 1317 -904 sw
rect 1136 -920 1317 -908
tri 1136 -943 1159 -920 ne
rect 1159 -943 1317 -920
tri 1252 -950 1259 -943 ne
rect 1259 -950 1317 -943
tri 1259 -956 1265 -950 ne
rect 1146 -1027 1202 -1018
rect 1146 -1088 1148 -1083
rect 1200 -1088 1202 -1083
rect 1146 -1107 1202 -1088
rect 1265 -1073 1317 -950
rect 3268 -1007 3320 -396
rect 3360 -878 3410 555
rect 3443 -832 3483 597
rect 3534 -746 3574 647
rect 3609 -274 3655 697
rect 4426 597 4432 649
rect 4484 597 4498 649
rect 4550 597 6485 649
rect 3845 407 4432 459
rect 4484 407 4498 459
rect 4550 407 4556 459
rect 3845 -119 3897 407
rect 3845 -184 3897 -171
rect 3845 -242 3897 -236
rect 6433 -241 6485 597
tri 3655 -274 3661 -268 sw
rect 3609 -280 3661 -274
rect 3609 -344 3661 -332
rect 6433 -305 6485 -293
rect 6433 -363 6485 -357
rect 3609 -403 3661 -396
rect 3609 -448 3661 -442
rect 3609 -512 3661 -500
rect 3609 -689 3661 -564
rect 3693 -528 3745 -522
rect 3693 -592 3745 -580
rect 3693 -650 3745 -644
tri 3745 -650 3767 -628 sw
tri 3693 -667 3710 -650 ne
rect 3710 -667 3767 -650
tri 3609 -716 3636 -689 ne
rect 3636 -699 3661 -689
tri 3661 -699 3693 -667 sw
tri 3710 -699 3742 -667 ne
rect 3742 -699 3767 -667
rect 3636 -716 3693 -699
tri 3693 -716 3710 -699 sw
tri 3742 -716 3759 -699 ne
rect 3759 -716 3767 -699
tri 3767 -716 3833 -650 sw
rect 6431 -716 6483 -710
tri 3636 -741 3661 -716 ne
rect 3661 -724 3710 -716
tri 3710 -724 3718 -716 sw
tri 3759 -724 3767 -716 ne
rect 3767 -724 3833 -716
tri 3833 -724 3841 -716 sw
rect 3661 -741 3718 -724
tri 3661 -743 3663 -741 ne
rect 3663 -743 3718 -741
tri 3574 -746 3577 -743 sw
tri 3663 -746 3666 -743 ne
rect 3666 -746 3718 -743
tri 3718 -746 3740 -724 sw
tri 3767 -746 3789 -724 ne
rect 3789 -746 3841 -724
tri 3841 -746 3863 -724 sw
rect 3534 -777 3577 -746
tri 3534 -798 3555 -777 ne
rect 3555 -785 3577 -777
tri 3577 -785 3616 -746 sw
tri 3666 -778 3698 -746 ne
rect 3698 -773 3740 -746
tri 3740 -773 3767 -746 sw
tri 3789 -773 3816 -746 ne
rect 3816 -773 6119 -746
rect 3698 -778 3767 -773
tri 3698 -785 3705 -778 ne
rect 3705 -785 3767 -778
rect 3555 -798 3616 -785
tri 3616 -798 3629 -785 sw
tri 3705 -798 3718 -785 ne
rect 3718 -798 3767 -785
tri 3767 -798 3792 -773 sw
tri 3816 -798 3841 -773 ne
rect 3841 -798 6119 -773
rect 6171 -798 6183 -746
rect 6235 -798 6241 -746
rect 6431 -780 6483 -768
tri 3555 -804 3561 -798 ne
rect 3561 -804 3629 -798
tri 3483 -832 3511 -804 sw
tri 3561 -817 3574 -804 ne
rect 3574 -817 3629 -804
tri 3574 -832 3589 -817 ne
rect 3589 -832 3629 -817
tri 3629 -832 3663 -798 sw
tri 3718 -832 3752 -798 ne
rect 3752 -832 3792 -798
tri 3792 -832 3826 -798 sw
rect 3443 -838 3511 -832
tri 3443 -852 3457 -838 ne
rect 3457 -849 3511 -838
tri 3511 -849 3528 -832 sw
tri 3589 -849 3606 -832 ne
rect 3606 -849 3663 -832
rect 3457 -852 3528 -849
tri 3528 -852 3531 -849 sw
tri 3606 -852 3609 -849 ne
rect 3609 -852 3663 -849
tri 3663 -852 3683 -832 sw
tri 3752 -852 3772 -832 ne
rect 3772 -852 3826 -832
tri 3826 -852 3846 -832 sw
rect 6431 -838 6483 -832
tri 3457 -855 3460 -852 ne
rect 3460 -855 3531 -852
tri 3410 -878 3433 -855 sw
tri 3460 -878 3483 -855 ne
rect 3483 -859 3531 -855
tri 3531 -859 3538 -852 sw
tri 3609 -859 3616 -852 ne
rect 3616 -859 3683 -852
tri 3683 -859 3690 -852 sw
tri 3772 -859 3779 -852 ne
rect 3779 -859 4409 -852
rect 3483 -878 3538 -859
rect 3360 -879 3433 -878
tri 3360 -904 3385 -879 ne
rect 3385 -904 3433 -879
tri 3433 -904 3459 -878 sw
tri 3483 -904 3509 -878 ne
rect 3509 -904 3538 -878
tri 3538 -904 3583 -859 sw
tri 3616 -904 3661 -859 ne
rect 3661 -904 3690 -859
tri 3690 -904 3735 -859 sw
tri 3779 -904 3824 -859 ne
rect 3824 -904 4409 -859
rect 4461 -904 4473 -852
rect 4525 -904 4531 -852
tri 3385 -929 3410 -904 ne
rect 3410 -923 3459 -904
tri 3459 -923 3478 -904 sw
tri 3509 -923 3528 -904 ne
rect 3528 -923 3583 -904
tri 3583 -923 3602 -904 sw
tri 3661 -923 3680 -904 ne
rect 3680 -923 3735 -904
rect 3410 -929 3478 -923
tri 3410 -950 3431 -929 ne
rect 3431 -950 3478 -929
tri 3478 -950 3505 -923 sw
tri 3528 -950 3555 -923 ne
rect 3555 -933 3602 -923
tri 3602 -933 3612 -923 sw
tri 3680 -933 3690 -923 ne
rect 3690 -933 3735 -923
tri 3735 -933 3764 -904 sw
rect 3555 -950 3612 -933
tri 3612 -950 3629 -933 sw
tri 3690 -950 3707 -933 ne
rect 3707 -950 4918 -933
tri 3431 -986 3467 -950 ne
rect 3467 -973 3505 -950
tri 3505 -973 3528 -950 sw
tri 3555 -973 3578 -950 ne
rect 3578 -973 3629 -950
rect 3467 -986 3528 -973
tri 3467 -997 3478 -986 ne
rect 3478 -997 3528 -986
tri 3528 -997 3552 -973 sw
tri 3578 -997 3602 -973 ne
rect 3602 -997 3629 -973
tri 3629 -997 3676 -950 sw
tri 3707 -967 3724 -950 ne
rect 3724 -967 4918 -950
rect 6587 -950 6639 -944
tri 3478 -1002 3483 -997 ne
rect 3483 -1002 3552 -997
tri 3552 -1002 3557 -997 sw
tri 3602 -1002 3607 -997 ne
rect 3607 -1002 4916 -997
tri 3483 -1007 3488 -1002 ne
rect 3488 -1007 3557 -1002
tri 1317 -1073 1330 -1060 sw
rect 1265 -1103 1456 -1073
tri 1265 -1125 1287 -1103 ne
rect 1287 -1125 1456 -1103
rect 1508 -1125 1520 -1073
rect 1572 -1125 1578 -1073
rect 1698 -1082 1704 -1030
rect 1756 -1082 1774 -1030
rect 1826 -1082 1844 -1030
rect 1896 -1082 1902 -1030
rect 3211 -1059 3217 -1007
rect 3269 -1059 3281 -1007
rect 3333 -1059 3339 -1007
tri 3488 -1014 3495 -1007 ne
rect 3495 -1014 3557 -1007
tri 3557 -1014 3569 -1002 sw
tri 3607 -1014 3619 -1002 ne
rect 3619 -1014 4916 -1002
tri 3495 -1059 3540 -1014 ne
rect 3540 -1031 3569 -1014
tri 3569 -1031 3586 -1014 sw
tri 3619 -1031 3636 -1014 ne
rect 3636 -1031 4916 -1014
rect 6587 -1014 6639 -1002
rect 3540 -1059 3586 -1031
tri 3540 -1060 3541 -1059 ne
rect 3541 -1060 3586 -1059
tri 3586 -1060 3615 -1031 sw
tri 3541 -1066 3547 -1060 ne
rect 3547 -1066 4903 -1060
tri 3547 -1082 3563 -1066 ne
rect 3563 -1082 4851 -1066
tri 3563 -1112 3593 -1082 ne
rect 3593 -1112 4851 -1082
tri 4833 -1118 4839 -1112 ne
rect 4839 -1118 4851 -1112
rect 6587 -1072 6639 -1066
tri 4839 -1125 4846 -1118 ne
rect 4846 -1125 4903 -1118
tri 4846 -1130 4851 -1125 ne
rect 4851 -1130 4903 -1125
tri 2121 -1156 2131 -1146 se
rect 2131 -1156 3874 -1146
tri 3874 -1156 3884 -1146 sw
rect 1146 -1164 1148 -1163
rect 1200 -1164 1202 -1163
rect 1146 -1172 1202 -1164
rect 1278 -1208 1284 -1156
rect 1336 -1208 1357 -1156
rect 1409 -1198 4696 -1156
rect 1409 -1208 2183 -1198
tri 2183 -1208 2193 -1198 nw
tri 3812 -1208 3822 -1198 ne
rect 3822 -1208 4696 -1198
rect 4748 -1208 4762 -1156
rect 4814 -1208 4820 -1156
rect 4851 -1188 4903 -1182
tri -1360 -1312 -1356 -1308 ne
rect -1356 -1312 -1286 -1308
tri -1286 -1312 -1282 -1308 sw
tri 1066 -1312 1070 -1308 se
rect 1070 -1312 1107 -1308
rect 4627 -1312 4633 -1308
tri -1356 -1326 -1342 -1312 ne
rect -1342 -1326 -1282 -1312
rect -2040 -1328 -1886 -1326
rect -2040 -1380 -2034 -1328
rect -1982 -1380 -1944 -1328
rect -1892 -1336 -1886 -1328
tri -1342 -1330 -1338 -1326 ne
rect -1338 -1330 -1282 -1326
tri -1282 -1330 -1264 -1312 sw
tri 1048 -1330 1066 -1312 se
rect 1066 -1330 1107 -1312
tri -1338 -1336 -1332 -1330 ne
rect -1332 -1336 1107 -1330
rect -1892 -1338 -1403 -1336
tri -1403 -1338 -1401 -1336 sw
tri -1332 -1338 -1330 -1336 ne
rect -1330 -1338 1107 -1336
rect -1892 -1364 -1401 -1338
tri -1401 -1364 -1375 -1338 sw
tri -1330 -1362 -1306 -1338 ne
rect -1306 -1344 1107 -1338
rect -1306 -1362 1089 -1344
tri 1089 -1362 1107 -1344 nw
rect 1278 -1364 1284 -1312
rect 1336 -1364 1350 -1312
rect 1402 -1360 4633 -1312
rect 4685 -1360 4699 -1308
rect 4751 -1360 4757 -1308
rect 1402 -1364 4757 -1360
rect -1892 -1372 -1375 -1364
rect -1892 -1380 -1886 -1372
rect -2040 -1382 -1886 -1380
tri -1423 -1382 -1413 -1372 ne
rect -1413 -1382 -1375 -1372
tri -1413 -1394 -1401 -1382 ne
rect -1401 -1394 -1375 -1382
tri -1375 -1394 -1345 -1364 sw
tri -1401 -1417 -1378 -1394 ne
rect -1378 -1417 4924 -1394
tri -2586 -1462 -2541 -1417 se
rect -2541 -1462 -1464 -1417
tri -1464 -1462 -1419 -1417 sw
tri -1378 -1430 -1365 -1417 ne
rect -1365 -1430 4924 -1417
tri -2631 -1507 -2586 -1462 se
rect -2586 -1469 1284 -1462
rect -2586 -1507 -2539 -1469
tri -2539 -1507 -2501 -1469 nw
tri -1514 -1507 -1476 -1469 ne
rect -1476 -1507 1284 -1469
rect -2609 -1512 -2544 -1507
tri -2544 -1512 -2539 -1507 nw
rect -2609 -1559 -2591 -1512
tri -2591 -1559 -2544 -1512 nw
rect -2487 -1564 -2481 -1512
rect -2429 -1564 -2417 -1512
rect -2365 -1514 -1936 -1512
tri -1936 -1514 -1934 -1512 sw
rect -2365 -1516 -1934 -1514
tri -1934 -1516 -1932 -1514 sw
rect -1867 -1516 -1811 -1507
rect -2365 -1535 -1932 -1516
tri -1932 -1535 -1913 -1516 sw
rect -2365 -1538 -1913 -1535
tri -1913 -1538 -1910 -1535 sw
rect -2365 -1564 -1910 -1538
tri -1973 -1582 -1955 -1564 ne
rect -2604 -1638 -1998 -1602
rect -2034 -1781 -1998 -1638
rect -1955 -1669 -1910 -1564
rect -1867 -1587 -1864 -1572
rect -1812 -1587 -1811 -1572
rect -1867 -1596 -1811 -1587
rect -1867 -1661 -1811 -1652
rect -1741 -1516 -1685 -1507
tri -1476 -1514 -1469 -1507 ne
rect -1469 -1514 1284 -1507
rect 1336 -1514 1350 -1462
rect 1402 -1464 4679 -1462
rect 1402 -1514 4550 -1464
rect 4544 -1516 4550 -1514
rect 4602 -1516 4621 -1464
rect 4673 -1516 4679 -1464
rect -1741 -1587 -1739 -1572
rect -1687 -1587 -1685 -1572
rect -1741 -1596 -1685 -1587
rect -1741 -1661 -1685 -1652
rect -1632 -1537 -1580 -1531
rect -1580 -1581 4926 -1545
rect -1632 -1603 -1580 -1589
rect -1632 -1661 -1580 -1655
tri -1315 -1661 -1271 -1617 se
rect -1271 -1661 1284 -1617
tri -1321 -1667 -1315 -1661 se
rect -1315 -1667 1284 -1661
tri -1910 -1669 -1908 -1667 sw
tri -1323 -1669 -1321 -1667 se
rect -1321 -1669 1284 -1667
rect 1336 -1669 1350 -1617
rect 1402 -1620 4684 -1617
rect 1402 -1669 4556 -1620
rect -1955 -1672 -1908 -1669
tri -1908 -1672 -1905 -1669 sw
tri -1326 -1672 -1323 -1669 se
rect -1323 -1672 -1250 -1669
tri -1250 -1672 -1247 -1669 nw
rect 4550 -1672 4556 -1669
rect 4608 -1672 4626 -1620
rect 4678 -1672 4684 -1620
rect 4851 -1621 4903 -1615
rect -1955 -1673 -1905 -1672
tri -1905 -1673 -1904 -1672 sw
tri -1327 -1673 -1326 -1672 se
rect -1326 -1673 -1251 -1672
tri -1251 -1673 -1250 -1672 nw
rect -1955 -1685 -1904 -1673
tri -1904 -1685 -1892 -1673 sw
tri -1339 -1685 -1327 -1673 se
rect -1327 -1685 -1263 -1673
tri -1263 -1685 -1251 -1673 nw
rect 4851 -1685 4903 -1673
rect -1955 -1691 -1892 -1685
tri -1892 -1691 -1886 -1685 sw
tri -1345 -1691 -1339 -1685 se
rect -1339 -1691 -1269 -1685
tri -1269 -1691 -1263 -1685 nw
rect -1955 -1719 -1315 -1691
tri -1955 -1737 -1937 -1719 ne
rect -1937 -1737 -1315 -1719
tri -1315 -1737 -1269 -1691 nw
tri -1262 -1737 -1232 -1707 se
rect -1232 -1737 4851 -1707
tri -1937 -1739 -1935 -1737 ne
rect -1935 -1739 -1317 -1737
tri -1317 -1739 -1315 -1737 nw
tri -1264 -1739 -1262 -1737 se
rect -1262 -1739 4903 -1737
tri -1268 -1743 -1264 -1739 se
rect -1264 -1743 4903 -1739
tri -1300 -1775 -1268 -1743 se
rect -1268 -1775 -1232 -1743
tri -1232 -1775 -1200 -1743 nw
tri -1306 -1781 -1300 -1775 se
rect -1300 -1781 -1274 -1775
rect -2034 -1817 -1274 -1781
tri -1274 -1817 -1232 -1775 nw
rect 1146 -2306 1202 -2299
rect 1146 -2308 1148 -2306
rect 1200 -2308 1202 -2306
rect 1146 -2382 1202 -2364
rect 1146 -2388 1148 -2382
rect 1200 -2388 1202 -2382
rect 1146 -2453 1202 -2444
rect 1011 -2507 1067 -2498
rect 1067 -2541 1758 -2535
rect 1067 -2563 1706 -2541
rect 1011 -2575 1706 -2563
rect 1011 -2587 1067 -2575
rect 1011 -2652 1067 -2643
rect 1706 -2607 1758 -2593
rect 1706 -2665 1758 -2659
rect -801 -4041 -792 -3985
rect -736 -4041 -705 -3985
rect -649 -4041 -618 -3985
rect -562 -4041 -532 -3985
rect -476 -4041 -446 -3985
rect -390 -4041 -360 -3985
rect -304 -4041 -274 -3985
rect -218 -3987 1633 -3985
rect -218 -4039 1511 -3987
rect 1563 -4039 1575 -3987
rect 1627 -4039 1633 -3987
rect -218 -4041 1633 -4039
<< via2 >>
rect -1741 685 -1691 728
rect -1691 685 -1685 728
rect -1741 672 -1685 685
rect -2168 548 -2112 604
rect -1741 592 -1685 648
rect -2168 461 -2112 517
rect -1821 88 -1765 144
rect -1741 88 -1685 144
rect -1750 -103 -1694 -47
rect -1670 -103 -1614 -47
rect -1867 -202 -1811 -146
rect -785 135 -738 173
rect -738 135 -729 173
rect -700 135 -673 173
rect -673 135 -660 173
rect -660 135 -644 173
rect -616 135 -608 173
rect -608 135 -595 173
rect -595 135 -560 173
rect -532 135 -530 173
rect -530 135 -478 173
rect -478 135 -476 173
rect -448 135 -413 173
rect -413 135 -400 173
rect -400 135 -392 173
rect -364 135 -348 173
rect -348 135 -335 173
rect -335 135 -308 173
rect -280 135 -270 173
rect -270 135 -224 173
rect -785 123 -729 135
rect -700 123 -644 135
rect -616 123 -560 135
rect -532 123 -476 135
rect -448 123 -392 135
rect -364 123 -308 135
rect -280 123 -224 135
rect -785 117 -738 123
rect -738 117 -729 123
rect -700 117 -673 123
rect -673 117 -660 123
rect -660 117 -644 123
rect -616 117 -608 123
rect -608 117 -595 123
rect -595 117 -560 123
rect -532 117 -530 123
rect -530 117 -478 123
rect -478 117 -476 123
rect -448 117 -413 123
rect -413 117 -400 123
rect -400 117 -392 123
rect -364 117 -348 123
rect -348 117 -335 123
rect -335 117 -308 123
rect -280 117 -270 123
rect -270 117 -224 123
rect -785 71 -738 93
rect -738 71 -729 93
rect -700 71 -673 93
rect -673 71 -660 93
rect -660 71 -644 93
rect -616 71 -608 93
rect -608 71 -595 93
rect -595 71 -560 93
rect -532 71 -530 93
rect -530 71 -478 93
rect -478 71 -476 93
rect -448 71 -413 93
rect -413 71 -400 93
rect -400 71 -392 93
rect -364 71 -348 93
rect -348 71 -335 93
rect -335 71 -308 93
rect -280 71 -270 93
rect -270 71 -224 93
rect -785 59 -729 71
rect -700 59 -644 71
rect -616 59 -560 71
rect -532 59 -476 71
rect -448 59 -392 71
rect -364 59 -308 71
rect -280 59 -224 71
rect -785 37 -738 59
rect -738 37 -729 59
rect -700 37 -673 59
rect -673 37 -660 59
rect -660 37 -644 59
rect -616 37 -608 59
rect -608 37 -595 59
rect -595 37 -560 59
rect -532 37 -530 59
rect -530 37 -478 59
rect -478 37 -476 59
rect -448 37 -413 59
rect -413 37 -400 59
rect -400 37 -392 59
rect -364 37 -348 59
rect -348 37 -335 59
rect -335 37 -308 59
rect -280 37 -270 59
rect -270 37 -224 59
rect -785 7 -738 13
rect -738 7 -729 13
rect -700 7 -673 13
rect -673 7 -660 13
rect -660 7 -644 13
rect -616 7 -608 13
rect -608 7 -595 13
rect -595 7 -560 13
rect -532 7 -530 13
rect -530 7 -478 13
rect -478 7 -476 13
rect -448 7 -413 13
rect -413 7 -400 13
rect -400 7 -392 13
rect -364 7 -348 13
rect -348 7 -335 13
rect -335 7 -308 13
rect -280 7 -270 13
rect -270 7 -224 13
rect -785 -5 -729 7
rect -700 -5 -644 7
rect -616 -5 -560 7
rect -532 -5 -476 7
rect -448 -5 -392 7
rect -364 -5 -308 7
rect -280 -5 -224 7
rect -785 -43 -738 -5
rect -738 -43 -729 -5
rect -700 -43 -673 -5
rect -673 -43 -660 -5
rect -660 -43 -644 -5
rect -616 -43 -608 -5
rect -608 -43 -595 -5
rect -595 -43 -560 -5
rect -532 -43 -530 -5
rect -530 -43 -478 -5
rect -478 -43 -476 -5
rect -448 -43 -413 -5
rect -413 -43 -400 -5
rect -400 -43 -392 -5
rect -364 -43 -348 -5
rect -348 -43 -335 -5
rect -335 -43 -308 -5
rect -280 -43 -270 -5
rect -270 -43 -224 -5
rect -1867 -282 -1811 -226
rect 1076 368 1132 369
rect 1076 316 1128 368
rect 1128 316 1132 368
rect 1076 313 1132 316
rect 1076 252 1128 289
rect 1128 252 1132 289
rect 1076 233 1132 252
rect -785 -994 -738 -944
rect -738 -994 -729 -944
rect -700 -994 -673 -944
rect -673 -994 -660 -944
rect -660 -994 -644 -944
rect -616 -994 -608 -944
rect -608 -994 -595 -944
rect -595 -994 -560 -944
rect -532 -994 -530 -944
rect -530 -994 -478 -944
rect -478 -994 -476 -944
rect -448 -994 -413 -944
rect -413 -994 -400 -944
rect -400 -994 -392 -944
rect -364 -994 -348 -944
rect -348 -994 -335 -944
rect -335 -994 -308 -944
rect -280 -994 -270 -944
rect -270 -994 -224 -944
rect -785 -1000 -729 -994
rect -700 -1000 -644 -994
rect -616 -1000 -560 -994
rect -532 -1000 -476 -994
rect -448 -1000 -392 -994
rect -364 -1000 -308 -994
rect -280 -1000 -224 -994
rect -785 -1078 -729 -1072
rect -700 -1078 -644 -1072
rect -616 -1078 -560 -1072
rect -532 -1078 -476 -1072
rect -448 -1078 -392 -1072
rect -364 -1078 -308 -1072
rect -280 -1078 -224 -1072
rect -785 -1128 -738 -1078
rect -738 -1128 -729 -1078
rect -700 -1128 -673 -1078
rect -673 -1128 -660 -1078
rect -660 -1128 -644 -1078
rect -616 -1128 -608 -1078
rect -608 -1128 -595 -1078
rect -595 -1128 -560 -1078
rect -532 -1128 -530 -1078
rect -530 -1128 -478 -1078
rect -478 -1128 -476 -1078
rect -448 -1128 -413 -1078
rect -413 -1128 -400 -1078
rect -400 -1128 -392 -1078
rect -364 -1128 -348 -1078
rect -348 -1128 -335 -1078
rect -335 -1128 -308 -1078
rect -280 -1128 -270 -1078
rect -270 -1128 -224 -1078
rect 1146 -1036 1202 -1027
rect 1146 -1083 1148 -1036
rect 1148 -1083 1200 -1036
rect 1200 -1083 1202 -1036
rect 1146 -1112 1202 -1107
rect 1146 -1163 1148 -1112
rect 1148 -1163 1200 -1112
rect 1200 -1163 1202 -1112
rect -1867 -1535 -1811 -1516
rect -1867 -1572 -1864 -1535
rect -1864 -1572 -1812 -1535
rect -1812 -1572 -1811 -1535
rect -1867 -1599 -1811 -1596
rect -1867 -1651 -1864 -1599
rect -1864 -1651 -1812 -1599
rect -1812 -1651 -1811 -1599
rect -1867 -1652 -1811 -1651
rect -1741 -1535 -1685 -1516
rect -1741 -1572 -1739 -1535
rect -1739 -1572 -1687 -1535
rect -1687 -1572 -1685 -1535
rect -1741 -1599 -1685 -1596
rect -1741 -1651 -1739 -1599
rect -1739 -1651 -1687 -1599
rect -1687 -1651 -1685 -1599
rect -1741 -1652 -1685 -1651
rect 1146 -2358 1148 -2308
rect 1148 -2358 1200 -2308
rect 1200 -2358 1202 -2308
rect 1146 -2364 1202 -2358
rect 1146 -2434 1148 -2388
rect 1148 -2434 1200 -2388
rect 1200 -2434 1202 -2388
rect 1146 -2444 1202 -2434
rect 1011 -2563 1067 -2507
rect 1011 -2643 1067 -2587
rect -792 -4041 -736 -3985
rect -705 -4041 -649 -3985
rect -618 -4041 -562 -3985
rect -532 -4041 -476 -3985
rect -446 -4041 -390 -3985
rect -360 -4041 -304 -3985
rect -274 -4041 -218 -3985
<< metal3 >>
rect -1746 728 -1680 733
rect -1746 672 -1741 728
rect -1685 672 -1680 728
rect -1746 648 -1680 672
rect -2173 604 -2107 609
rect -2173 548 -2168 604
rect -2112 548 -2107 604
rect -2173 517 -2107 548
rect -2173 461 -2168 517
rect -2112 461 -2107 517
rect -2173 456 -2107 461
rect -1746 592 -1741 648
rect -1685 592 -1680 648
rect -1746 149 -1680 592
rect 1071 369 1137 374
rect 1071 313 1076 369
rect 1132 313 1137 369
rect 1071 294 1137 313
rect 1006 289 1137 294
rect 1006 233 1076 289
rect 1132 233 1137 289
rect 1006 228 1137 233
rect -1826 144 -1680 149
rect -1826 88 -1821 144
rect -1765 88 -1741 144
rect -1685 88 -1680 144
rect -1826 83 -1680 88
rect -801 173 -209 195
rect -801 117 -785 173
rect -729 117 -700 173
rect -644 117 -616 173
rect -560 117 -532 173
rect -476 117 -448 173
rect -392 117 -364 173
rect -308 117 -280 173
rect -224 117 -209 173
rect -801 93 -209 117
rect -801 37 -785 93
rect -729 37 -700 93
rect -644 37 -616 93
rect -560 37 -532 93
rect -476 37 -448 93
rect -392 37 -364 93
rect -308 37 -280 93
rect -224 37 -209 93
rect -801 13 -209 37
rect -1755 -47 -1609 -42
rect -1755 -103 -1750 -47
rect -1694 -103 -1670 -47
rect -1614 -103 -1609 -47
rect -1755 -108 -1609 -103
rect -801 -43 -785 13
rect -729 -43 -700 13
rect -644 -43 -616 13
rect -560 -43 -532 13
rect -476 -43 -448 13
rect -392 -43 -364 13
rect -308 -43 -280 13
rect -224 -43 -209 13
rect -1872 -146 -1806 -141
rect -1872 -202 -1867 -146
rect -1811 -202 -1806 -146
rect -1872 -226 -1806 -202
rect -1872 -282 -1867 -226
rect -1811 -282 -1806 -226
rect -1872 -1516 -1806 -282
rect -1872 -1572 -1867 -1516
rect -1811 -1572 -1806 -1516
rect -1872 -1596 -1806 -1572
rect -1872 -1652 -1867 -1596
rect -1811 -1652 -1806 -1596
rect -1872 -1657 -1806 -1652
rect -1746 -1516 -1680 -108
rect -801 -944 -209 -43
rect -801 -1000 -785 -944
rect -729 -1000 -700 -944
rect -644 -1000 -616 -944
rect -560 -1000 -532 -944
rect -476 -1000 -448 -944
rect -392 -1000 -364 -944
rect -308 -1000 -280 -944
rect -224 -1000 -209 -944
rect -801 -1072 -209 -1000
rect -801 -1128 -785 -1072
rect -729 -1128 -700 -1072
rect -644 -1128 -616 -1072
rect -560 -1128 -532 -1072
rect -476 -1128 -448 -1072
rect -392 -1128 -364 -1072
rect -308 -1128 -280 -1072
rect -224 -1128 -209 -1072
rect -801 -1133 -209 -1128
rect -1746 -1572 -1741 -1516
rect -1685 -1572 -1680 -1516
rect -1746 -1596 -1680 -1572
rect -1746 -1652 -1741 -1596
rect -1685 -1652 -1680 -1596
rect -1746 -1657 -1680 -1652
rect 1006 -2507 1072 228
rect 1141 -1027 1207 -1022
rect 1141 -1083 1146 -1027
rect 1202 -1083 1207 -1027
rect 1141 -1107 1207 -1083
rect 1141 -1163 1146 -1107
rect 1202 -1163 1207 -1107
rect 1141 -2308 1207 -1163
rect 1141 -2364 1146 -2308
rect 1202 -2364 1207 -2308
rect 1141 -2388 1207 -2364
rect 1141 -2444 1146 -2388
rect 1202 -2444 1207 -2388
rect 1141 -2449 1207 -2444
rect 1006 -2563 1011 -2507
rect 1067 -2563 1072 -2507
rect 1006 -2587 1072 -2563
rect 1006 -2643 1011 -2587
rect 1067 -2643 1072 -2587
rect 1006 -2673 1072 -2643
rect -797 -3985 -213 -3980
rect -797 -4041 -792 -3985
rect -736 -4041 -705 -3985
rect -649 -4041 -618 -3985
rect -562 -4041 -532 -3985
rect -476 -4041 -446 -3985
rect -390 -4041 -360 -3985
rect -304 -4041 -274 -3985
rect -218 -4041 -213 -3985
rect -797 -4046 -213 -4041
use sky130_fd_io__gpio_ovtv2_amux_nand4  sky130_fd_io__gpio_ovtv2_amux_nand4_0
timestamp 1704896540
transform -1 0 2247 0 -1 834
box -44 33 1013 1822
use sky130_fd_io__gpio_ovtv2_amux_nand4  sky130_fd_io__gpio_ovtv2_amux_nand4_1
timestamp 1704896540
transform 1 0 2195 0 -1 834
box -44 33 1013 1822
use sky130_fd_io__gpio_ovtv2_amux_nand5  sky130_fd_io__gpio_ovtv2_amux_nand5_0
timestamp 1704896540
transform 0 -1 4886 1 0 -2138
box 33 38 1194 1846
use sky130_fd_io__gpio_ovtv2_amux_nand5  sky130_fd_io__gpio_ovtv2_amux_nand5_1
timestamp 1704896540
transform 0 1 1238 1 0 -2138
box 33 38 1194 1846
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1704896540
transform -1 0 -791 0 1 -1993
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1704896540
transform -1 0 -326 0 1 -1993
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1704896540
transform 1 0 -1876 0 1 -1993
box 107 226 460 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1704896540
transform -1 0 -1694 0 1 -1993
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1704896540
transform -1 0 613 0 1 -1993
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1704896540
transform 1 0 -392 0 1 -1993
box 107 226 460 873
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_0
timestamp 1704896540
transform 1 0 1505 0 -1 -2417
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_1
timestamp 1704896540
transform 1 0 -252 0 1 -680
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_2
timestamp 1704896540
transform 1 0 -2556 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_3
timestamp 1704896540
transform 1 0 -2268 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_4
timestamp 1704896540
transform -1 0 804 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_5
timestamp 1704896540
transform -1 0 1092 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_6
timestamp 1704896540
transform 1 0 -444 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_7
timestamp 1704896540
transform 1 0 -1692 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_8
timestamp 1704896540
transform 1 0 -1404 0 1 -680
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_9
timestamp 1704896540
transform -1 0 132 0 -1 814
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_10
timestamp 1704896540
transform -1 0 708 0 1 -680
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_11
timestamp 1704896540
transform -1 0 420 0 1 -680
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_12
timestamp 1704896540
transform 1 0 -2268 0 1 -680
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_13
timestamp 1704896540
transform 1 0 -1692 0 1 -680
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_14
timestamp 1704896540
transform 1 0 -828 0 1 -680
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_0
timestamp 1704896540
transform 1 0 132 0 -1 814
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_1
timestamp 1704896540
transform 1 0 708 0 1 -680
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_2
timestamp 1704896540
transform 1 0 -1980 0 -1 814
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_3
timestamp 1704896540
transform 1 0 -732 0 -1 814
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_0
timestamp 1704896540
transform 1 0 -1116 0 1 -680
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_1
timestamp 1704896540
transform 1 0 -540 0 1 -680
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_2
timestamp 1704896540
transform 1 0 -1980 0 1 -680
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_3
timestamp 1704896540
transform 1 0 -2556 0 1 -680
box -38 -49 326 715
use sky130_fd_io__xor2_1  sky130_fd_io__xor2_1_0
timestamp 1704896540
transform 1 0 -1404 0 -1 814
box 0 0 1 1
<< labels >>
flabel metal3 s -528 -820 -500 -792 3 FreeSans 280 0 0 0 VCCD
port 1 nsew
flabel comment s 629 -114 629 -114 0 FreeSans 280 0 0 0 OUT_I_N
flabel comment s -2049 674 -2049 674 0 FreeSans 280 90 0 0 ANA_SEL_I
flabel comment s 1244 618 1244 618 0 FreeSans 280 0 0 0 INT_AMUXB_ON
flabel comment s -1463 532 -1463 532 0 FreeSans 280 90 0 0 INT_AMUXA_ON
flabel comment s 1070 422 1070 422 0 FreeSans 280 0 0 0 INT_AMUXA_ON
flabel comment s -433 369 -433 369 0 FreeSans 280 0 0 0 ANA_POL_I
flabel comment s 999 -1716 999 -1716 0 FreeSans 280 0 0 0 PD_CSD_VSWITCH_H_N
flabel comment s 4835 -1561 4835 -1561 0 FreeSans 280 0 0 0 NMIDB_ON_N
flabel comment s 4802 -1410 4802 -1410 0 FreeSans 280 0 0 0 NMIDA_ON_N
flabel comment s 478 -950 478 -950 0 FreeSans 280 0 0 0 LV_NET
flabel comment s -2343 -1703 -2343 -1703 0 FreeSans 280 0 0 0 NGA_PAD_VSWITCH_H
flabel metal1 s 262 -666 290 -638 3 FreeSans 280 0 0 0 VSSD
port 2 nsew
flabel metal1 s 646 773 674 801 3 FreeSans 280 0 0 0 VSSD
port 2 nsew
flabel metal1 s -26 -266 2 -238 3 FreeSans 280 0 0 0 AMUXBUSA_ON_N
port 3 nsew
flabel metal1 s -213 -391 -185 -363 3 FreeSans 280 0 0 0 AMUXBUSA_ON
port 4 nsew
flabel metal1 s 262 -3 290 25 3 FreeSans 280 0 0 0 VCCD
port 1 nsew
flabel metal1 s -2522 465 -2494 493 3 FreeSans 280 0 0 0 ANALOG_SEL
port 5 nsew
flabel metal1 s 1030 482 1058 510 3 FreeSans 280 0 0 0 ANALOG_POL
port 6 nsew
flabel metal1 s -1370 -361 -1342 -333 3 FreeSans 280 0 0 0 ANALOG_EN
port 7 nsew
flabel metal1 s 646 -382 674 -354 3 FreeSans 280 0 0 0 OUT
port 8 nsew
flabel metal1 s -2042 -210 -2014 -182 3 FreeSans 280 0 0 0 AMUXBUSB_ON_N
port 9 nsew
flabel metal1 s -2234 -361 -2206 -333 3 FreeSans 280 0 0 0 AMUXBUSB_ON
port 10 nsew
flabel metal1 s -1466 -295 -1438 -267 3 FreeSans 280 0 0 0 PU_ON_N
port 11 nsew
flabel metal1 s -1658 -361 -1630 -333 3 FreeSans 280 0 0 0 PU_ON
port 12 nsew
flabel metal1 s -602 -321 -574 -293 3 FreeSans 280 0 0 0 PD_ON_N
port 13 nsew
flabel metal1 s -794 -361 -766 -333 3 FreeSans 280 0 0 0 PD_ON
port 14 nsew
flabel metal1 s -217 -1646 -189 -1618 3 FreeSans 280 90 0 0 NGA_PAD_VSWITCH_H
port 15 nsew
flabel metal1 s -460 -1034 -432 -1006 3 FreeSans 280 0 0 0 VCCD
port 1 nsew
flabel metal1 s -429 -1857 -401 -1829 3 FreeSans 280 0 0 0 VSSD
port 2 nsew
flabel metal1 s -991 -1315 -963 -1287 3 FreeSans 280 90 0 0 PGA_PAD_VDDIOQ_H_N
port 16 nsew
flabel metal1 s -1156 -1414 -1128 -1386 3 FreeSans 280 90 0 0 PGA_AMX_VDDA_H_N
port 17 nsew
flabel metal1 s -513 -1420 -485 -1392 3 FreeSans 280 90 0 0 PGB_PAD_VDDIOQ_H_N
port 18 nsew
flabel metal1 s -698 -1366 -670 -1338 3 FreeSans 280 270 0 0 PGB_AMX_VDDA_H_N
port 19 nsew
flabel metal1 s -1621 -1612 -1593 -1584 3 FreeSans 280 0 0 0 D_B
port 20 nsew
flabel metal1 s -1971 -1361 -1943 -1333 3 FreeSans 280 0 0 0 NMIDA_ON_N
port 21 nsew
flabel metal1 s 410 -1228 438 -1200 3 FreeSans 280 180 0 0 NGB_PAD_VSWITCH_H
port 22 nsew
flabel metal1 s 1741 697 1769 725 3 FreeSans 280 0 0 0 D_B
port 20 nsew
flabel metal1 s 1429 697 1457 725 3 FreeSans 280 0 0 0 PU_VDDIOQ_H_N
port 23 nsew
flabel metal1 s 4561 -1662 4589 -1634 3 FreeSans 280 0 0 0 NGB_PAD_VSWITCH_H_N
port 24 nsew
flabel metal1 s 2143 457 2171 485 3 FreeSans 280 0 0 0 VSSD
port 2 nsew
flabel metal1 s 1770 -957 1798 -929 3 FreeSans 280 0 0 0 VCCD
port 1 nsew
flabel metal1 s 4571 -1506 4599 -1478 3 FreeSans 280 0 0 0 NGA_PAD_VSWITCH_H_N
port 25 nsew
flabel metal1 s 1585 697 1613 725 3 FreeSans 280 0 0 0 PD_VSWITCH_H_N
port 26 nsew
flabel metal1 s 2673 697 2701 725 3 FreeSans 280 0 0 0 NMIDA_VCCD_N
port 27 nsew
<< properties >>
string FIXED_BBOX -1404 148 -732 814
string GDS_END 64983414
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 64877712
<< end >>
