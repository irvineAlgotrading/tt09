magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 415 206
<< mvpmos >>
rect 0 0 120 140
rect 176 0 296 140
<< mvpdiff >>
rect -53 114 0 140
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 120 114 176 140
rect 120 80 131 114
rect 165 80 176 114
rect 120 46 176 80
rect 120 12 131 46
rect 165 12 176 46
rect 120 0 176 12
rect 296 114 349 140
rect 296 80 307 114
rect 341 80 349 114
rect 296 46 349 80
rect 296 12 307 46
rect 341 12 349 46
rect 296 0 349 12
<< mvpdiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 131 80 165 114
rect 131 12 165 46
rect 307 80 341 114
rect 307 12 341 46
<< poly >>
rect 0 140 120 172
rect 176 140 296 172
rect 0 -32 120 0
rect 176 -32 296 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 80
rect -45 -4 -11 12
rect 131 114 165 130
rect 131 46 165 80
rect 131 -4 165 12
rect 307 114 341 130
rect 307 46 341 80
rect 307 -4 341 12
use DFL1sd2_CDNS_52468879185693  DFL1sd2_CDNS_52468879185693_0
timestamp 1704896540
transform 1 0 120 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185486  DFL1sd_CDNS_52468879185486_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185486  DFL1sd_CDNS_52468879185486_1
timestamp 1704896540
transform 1 0 296 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
flabel comment s 148 63 148 63 0 FreeSans 300 0 0 0 D
flabel comment s 324 63 324 63 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 89239406
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89237894
<< end >>
