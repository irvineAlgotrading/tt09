magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_0
timestamp 1704896540
transform -1 0 -16 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_1
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 9656940
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 9655954
<< end >>
