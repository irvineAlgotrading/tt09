magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 450 897
<< pwell >>
rect 16 43 378 295
rect -26 -43 410 43
<< obsli1 >>
rect 0 797 384 831
rect 50 537 340 751
rect 95 250 161 406
rect 203 340 269 537
rect 95 169 356 250
rect 34 73 356 169
rect 0 -17 384 17
<< metal1 >>
rect 0 791 384 837
rect 0 689 384 763
rect 0 51 384 125
rect 0 -23 384 23
<< labels >>
rlabel metal1 s 0 51 384 125 6 VGND
port 1 nsew ground bidirectional
rlabel metal1 s 0 -23 384 23 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s -26 -43 410 43 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s 16 43 378 295 6 VNB
port 2 nsew ground bidirectional
rlabel metal1 s 0 791 384 837 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -66 377 450 897 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 689 384 763 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 384 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 959862
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 955112
<< end >>
