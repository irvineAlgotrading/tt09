magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< metal4 >>
tri 226 14000 766 14540 se
rect 766 14000 11234 14540
tri 11234 14000 11774 14540 sw
tri 0 13774 226 14000 se
tri -540 13234 0 13774 se
rect 0 13236 226 13774
tri 226 13236 990 14000 nw
tri 11010 13774 11236 14000 ne
rect 11236 13774 11774 14000
tri 11774 13774 12000 14000 sw
tri 11236 13236 11774 13774 ne
rect 11774 13236 12000 13774
rect -540 766 0 13234
tri 0 13010 226 13236 nw
tri 11774 13010 12000 13236 ne
tri 12000 13234 12540 13774 sw
tri -540 226 0 766 ne
tri 0 226 764 990 sw
tri 11774 764 12000 990 se
rect 12000 766 12540 13234
tri 11236 226 11774 764 se
rect 11774 226 12000 764
tri 12000 226 12540 766 nw
tri 0 0 226 226 ne
rect 226 0 764 226
tri 764 0 990 226 sw
tri 11010 0 11236 226 se
rect 11236 0 11774 226
tri 11774 0 12000 226 nw
tri 226 -540 766 0 ne
rect 766 -540 11234 0
tri 11234 -540 11774 0 nw
<< metal5 >>
tri -540 13234 766 14540 se
rect 766 13234 11234 14540
tri 11234 13234 12540 14540 sw
rect -540 766 12540 13234
tri -540 -540 766 766 ne
rect 766 -540 11234 766
tri 11234 -540 12540 766 nw
<< glass >>
tri 0 13010 990 14000 se
rect 990 13010 11010 14000
tri 11010 13010 12000 14000 sw
rect 0 990 12000 13010
tri 0 0 990 990 ne
rect 990 0 11010 990
tri 11010 0 12000 990 nw
use genDLring_CDNS_5246887918517  genDLring_CDNS_5246887918517_0
timestamp 1704896540
transform 1 0 0 0 1 0
box 0 0 1 1
use genRivetDLring_CDNS_5246887918518  genRivetDLring_CDNS_5246887918518_0
timestamp 1704896540
transform 1 0 -478 0 1 -478
box -38 -38 12994 14994
<< labels >>
flabel comment s 6000 7000 6000 7000 0 FreeSans 1600 0 0 0 plastic
flabel comment s 6000 7000 6000 7000 0 FreeSans 1600 0 0 0 plastic
flabel comment s 6000 6666 6000 6666 0 FreeSans 1600 0 0 0 HP
<< properties >>
string GDS_END 85509582
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85508748
<< end >>
