magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -54 284 204 454
rect -59 116 209 284
rect -54 -54 204 116
<< scpmos >>
rect 60 0 90 400
<< pdiff >>
rect 0 217 60 400
rect 0 183 8 217
rect 42 183 60 217
rect 0 0 60 183
rect 90 217 150 400
rect 90 183 108 217
rect 142 183 150 217
rect 90 0 150 183
<< pdiffc >>
rect 8 183 42 217
rect 108 183 142 217
<< poly >>
rect 60 400 90 426
rect 60 -26 90 0
<< locali >>
rect 8 217 42 233
rect 8 167 42 183
rect 108 217 142 233
rect 108 167 142 183
use contact_11  contact_11_0
timestamp 1704896540
transform 1 0 100 0 1 167
box 0 0 1 1
use contact_11  contact_11_1
timestamp 1704896540
transform 1 0 0 0 1 167
box 0 0 1 1
<< labels >>
rlabel locali s 125 200 125 200 4 D
port 1 nsew
rlabel locali s 25 200 25 200 4 S
port 2 nsew
rlabel poly s 75 200 75 200 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -54 204 116
string GDS_END 58898
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 58082
<< end >>
