magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 203
rect 29 -17 63 21
<< locali >>
rect 118 291 168 425
rect 17 212 84 257
rect 118 119 156 291
rect 207 289 247 422
rect 207 265 241 289
rect 191 231 241 265
rect 191 199 225 231
rect 652 152 719 324
<< obsli1 >>
rect 0 527 736 561
rect 24 459 315 493
rect 24 291 84 459
rect 17 93 69 177
rect 281 330 315 459
rect 349 367 395 527
rect 457 330 523 493
rect 281 296 523 330
rect 572 262 617 493
rect 659 367 718 527
rect 277 215 617 262
rect 259 165 524 177
rect 191 143 524 165
rect 191 131 304 143
rect 17 85 88 93
rect 193 85 361 93
rect 17 51 361 85
rect 395 17 429 109
rect 477 51 524 143
rect 560 97 617 215
rect 560 51 633 97
rect 667 17 711 109
rect 0 -17 736 17
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 17 212 84 257 6 A0
port 1 nsew signal input
rlabel locali s 191 199 225 231 6 A1
port 2 nsew signal input
rlabel locali s 191 231 241 265 6 A1
port 2 nsew signal input
rlabel locali s 207 265 241 289 6 A1
port 2 nsew signal input
rlabel locali s 207 289 247 422 6 A1
port 2 nsew signal input
rlabel locali s 652 152 719 324 6 S
port 3 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 735 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 118 119 156 291 6 Y
port 8 nsew signal output
rlabel locali s 118 291 168 425 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1705468
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1698572
<< end >>
