magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 131 0 160
rect -50 97 -34 131
rect -50 63 0 97
rect -50 29 -34 63
rect -50 0 0 29
rect 1200 131 1250 160
rect 1234 97 1250 131
rect 1200 63 1250 97
rect 1234 29 1250 63
rect 1200 0 1250 29
<< polycont >>
rect -34 97 0 131
rect -34 29 0 63
rect 1200 97 1234 131
rect 1200 29 1234 63
<< npolyres >>
rect 0 0 1200 160
<< locali >>
rect -34 131 0 147
rect -34 63 0 97
rect -34 13 0 29
rect 1200 131 1234 147
rect 1200 63 1234 97
rect 1200 13 1234 29
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 1 0 1184 0 1 13
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 1 0 -50 0 1 13
box 0 0 1 1
<< properties >>
string GDS_END 90828934
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90828450
<< end >>
