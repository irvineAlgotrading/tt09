magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 336 12495 18396 17444
<< nwell >>
rect 256 17220 18476 17524
rect 256 12719 560 17220
rect 18172 12719 18476 17220
rect 256 12415 18476 12719
rect 10069 3490 15897 3792
rect 10069 359 10371 3490
rect 15595 359 15897 3490
rect 10069 0 15897 359
<< pwell >>
rect -26 17631 18805 17853
rect -26 12275 196 17631
rect 620 16938 18112 17160
rect 620 13001 842 16938
rect 10405 16718 15676 16938
rect 15045 16106 15676 16718
rect 15045 15981 15608 16106
rect 15155 15139 15608 15981
rect 15056 13867 15608 15139
rect 15135 13241 15608 13867
rect 15252 13001 15608 13241
rect 17890 13001 18112 16938
rect 620 12779 18112 13001
rect 18583 12275 18805 17631
rect -26 12053 18805 12275
rect 11946 7717 12168 12053
rect 17894 7717 18116 12053
rect 11946 7495 18116 7717
rect 10465 3208 15535 3430
rect 10465 724 10687 3208
rect 15313 724 15535 3208
rect 10465 502 15535 724
<< psubdiff >>
rect 0 17793 102 17827
rect 15640 17793 15675 17827
rect 15709 17793 15744 17827
rect 15778 17793 15813 17827
rect 15847 17793 15882 17827
rect 15916 17793 15951 17827
rect 15985 17793 16020 17827
rect 16054 17793 16089 17827
rect 16123 17793 16158 17827
rect 16192 17793 16227 17827
rect 16261 17793 16296 17827
rect 16330 17793 16365 17827
rect 16399 17793 16434 17827
rect 16468 17793 16503 17827
rect 16537 17793 16572 17827
rect 16606 17793 16641 17827
rect 16675 17793 16710 17827
rect 16744 17793 16779 17827
rect 16813 17793 16848 17827
rect 16882 17793 16917 17827
rect 16951 17793 16986 17827
rect 17020 17793 17055 17827
rect 17089 17793 17124 17827
rect 17158 17793 17193 17827
rect 17227 17793 17262 17827
rect 17296 17793 17331 17827
rect 17365 17793 17400 17827
rect 17434 17793 17469 17827
rect 17503 17793 17538 17827
rect 17572 17793 17607 17827
rect 17641 17793 17676 17827
rect 17710 17793 17745 17827
rect 17779 17793 17814 17827
rect 17848 17793 17883 17827
rect 17917 17793 17952 17827
rect 17986 17793 18021 17827
rect 18055 17793 18090 17827
rect 18124 17793 18159 17827
rect 18193 17793 18228 17827
rect 18262 17793 18297 17827
rect 18331 17793 18366 17827
rect 18400 17793 18435 17827
rect 18469 17793 18504 17827
rect 18538 17793 18573 17827
rect 18607 17793 18642 17827
rect 18676 17793 18711 17827
rect 18745 17793 18779 17827
rect 34 17759 102 17793
rect 15606 17759 18779 17793
rect 0 17725 68 17759
rect 15606 17725 15641 17759
rect 15675 17725 15710 17759
rect 15744 17725 15779 17759
rect 15813 17725 15848 17759
rect 15882 17725 15917 17759
rect 15951 17725 15986 17759
rect 16020 17725 16055 17759
rect 16089 17725 16124 17759
rect 16158 17725 16193 17759
rect 16227 17725 16262 17759
rect 16296 17725 16331 17759
rect 16365 17725 16400 17759
rect 16434 17725 16469 17759
rect 16503 17725 16538 17759
rect 16572 17725 16607 17759
rect 16641 17725 16676 17759
rect 16710 17725 16745 17759
rect 16779 17725 16814 17759
rect 16848 17725 16883 17759
rect 16917 17725 16952 17759
rect 16986 17725 17021 17759
rect 17055 17725 17090 17759
rect 17124 17725 17159 17759
rect 17193 17725 17228 17759
rect 17262 17725 17297 17759
rect 17331 17725 17366 17759
rect 17400 17725 17435 17759
rect 17469 17725 17504 17759
rect 17538 17725 17573 17759
rect 17607 17725 17642 17759
rect 17676 17725 17711 17759
rect 17745 17725 17780 17759
rect 17814 17725 17849 17759
rect 17883 17725 17918 17759
rect 17952 17725 17987 17759
rect 18021 17725 18056 17759
rect 18090 17725 18125 17759
rect 18159 17725 18194 17759
rect 18228 17725 18263 17759
rect 18297 17725 18332 17759
rect 18366 17725 18401 17759
rect 18435 17725 18470 17759
rect 18504 17725 18539 17759
rect 18573 17725 18608 17759
rect 18642 17725 18677 17759
rect 18711 17725 18779 17759
rect 0 17723 136 17725
rect 34 17690 136 17723
rect 34 17689 68 17690
rect 0 17656 68 17689
rect 102 17657 136 17690
rect 15538 17691 18677 17725
rect 15538 17657 15573 17691
rect 15607 17657 15642 17691
rect 15676 17657 15711 17691
rect 15745 17657 15780 17691
rect 15814 17657 15849 17691
rect 15883 17657 15918 17691
rect 15952 17657 15987 17691
rect 16021 17657 16056 17691
rect 16090 17657 16125 17691
rect 16159 17657 16194 17691
rect 16228 17657 16263 17691
rect 16297 17657 16332 17691
rect 16366 17657 16401 17691
rect 16435 17657 16470 17691
rect 16504 17657 16539 17691
rect 16573 17657 16608 17691
rect 16642 17657 16677 17691
rect 16711 17657 16746 17691
rect 16780 17657 16815 17691
rect 16849 17657 16884 17691
rect 16918 17657 16953 17691
rect 16987 17657 17022 17691
rect 17056 17657 17091 17691
rect 17125 17657 17160 17691
rect 17194 17657 17229 17691
rect 17263 17657 17298 17691
rect 17332 17657 17367 17691
rect 17401 17657 17436 17691
rect 17470 17657 17505 17691
rect 17539 17657 17574 17691
rect 17608 17657 17643 17691
rect 17677 17657 17712 17691
rect 17746 17657 17781 17691
rect 17815 17657 17850 17691
rect 17884 17657 17919 17691
rect 17953 17657 17988 17691
rect 18022 17657 18057 17691
rect 18091 17657 18126 17691
rect 18160 17657 18195 17691
rect 18229 17657 18264 17691
rect 18298 17657 18333 17691
rect 18367 17657 18402 17691
rect 18436 17657 18471 17691
rect 18505 17657 18540 17691
rect 18574 17657 18609 17691
rect 102 17656 170 17657
rect 0 17653 170 17656
rect 34 17622 170 17653
rect 34 17621 136 17622
rect 34 17619 68 17621
rect 0 17587 68 17619
rect 102 17588 136 17621
rect 102 17587 170 17588
rect 0 17583 170 17587
rect 34 17553 170 17583
rect 34 17552 136 17553
rect 34 17549 68 17552
rect 0 17518 68 17549
rect 102 17519 136 17552
rect 102 17518 170 17519
rect 0 17513 170 17518
rect 34 17484 170 17513
rect 34 17483 136 17484
rect 34 17479 68 17483
rect 0 17449 68 17479
rect 102 17450 136 17483
rect 102 17449 170 17450
rect 0 17443 170 17449
rect 34 17415 170 17443
rect 34 17414 136 17415
rect 34 17409 68 17414
rect 0 17380 68 17409
rect 102 17381 136 17414
rect 102 17380 170 17381
rect 0 17373 170 17380
rect 34 17346 170 17373
rect 34 17345 136 17346
rect 34 17339 68 17345
rect 0 17311 68 17339
rect 102 17312 136 17345
rect 102 17311 170 17312
rect 0 17303 170 17311
rect 34 17277 170 17303
rect 34 17276 136 17277
rect 34 17269 68 17276
rect 0 17242 68 17269
rect 102 17243 136 17276
rect 102 17242 170 17243
rect 0 17233 170 17242
rect 34 17208 170 17233
rect 34 17207 136 17208
rect 34 17199 68 17207
rect 0 17173 68 17199
rect 102 17174 136 17207
rect 102 17173 170 17174
rect 0 17164 170 17173
rect 34 17139 170 17164
rect 34 17138 136 17139
rect 34 17130 68 17138
rect 0 17104 68 17130
rect 102 17105 136 17138
rect 102 17104 170 17105
rect 0 17095 170 17104
rect 34 17070 170 17095
rect 34 17069 136 17070
rect 34 17061 68 17069
rect 0 17035 68 17061
rect 102 17036 136 17069
rect 102 17035 170 17036
rect 0 17026 170 17035
rect 34 17001 170 17026
rect 34 17000 136 17001
rect 34 16992 68 17000
rect 0 16966 68 16992
rect 102 16967 136 17000
rect 102 16966 170 16967
rect 0 16957 170 16966
rect 34 16932 170 16957
rect 34 16931 136 16932
rect 34 16923 68 16931
rect 0 16897 68 16923
rect 102 16898 136 16931
rect 102 16897 170 16898
rect 0 16888 170 16897
rect 34 16863 170 16888
rect 34 16862 136 16863
rect 34 16854 68 16862
rect 0 16828 68 16854
rect 102 16829 136 16862
rect 102 16828 170 16829
rect 0 16819 170 16828
rect 34 16794 170 16819
rect 34 16793 136 16794
rect 34 16785 68 16793
rect 0 16759 68 16785
rect 102 16760 136 16793
rect 102 16759 170 16760
rect 0 16750 170 16759
rect 34 16725 170 16750
rect 34 16724 136 16725
rect 34 16716 68 16724
rect 0 16690 68 16716
rect 102 16691 136 16724
rect 102 16690 170 16691
rect 0 16681 170 16690
rect 34 16656 170 16681
rect 34 16655 136 16656
rect 34 16647 68 16655
rect 0 16621 68 16647
rect 102 16622 136 16655
rect 102 16621 170 16622
rect 0 16612 170 16621
rect 34 16587 170 16612
rect 34 16586 136 16587
rect 34 16578 68 16586
rect 0 16552 68 16578
rect 102 16553 136 16586
rect 102 16552 170 16553
rect 0 16543 170 16552
rect 34 16518 170 16543
rect 34 16517 136 16518
rect 34 16509 68 16517
rect 0 16483 68 16509
rect 102 16484 136 16517
rect 102 16483 170 16484
rect 0 16474 170 16483
rect 34 16449 170 16474
rect 34 16448 136 16449
rect 34 16440 68 16448
rect 0 16414 68 16440
rect 102 16415 136 16448
rect 102 16414 170 16415
rect 0 16405 170 16414
rect 34 16380 170 16405
rect 34 16379 136 16380
rect 34 16371 68 16379
rect 0 16345 68 16371
rect 102 16346 136 16379
rect 102 16345 170 16346
rect 0 16336 170 16345
rect 34 16311 170 16336
rect 34 16310 136 16311
rect 34 16302 68 16310
rect 0 16276 68 16302
rect 102 16277 136 16310
rect 102 16276 170 16277
rect 0 16267 170 16276
rect 34 16242 170 16267
rect 34 16241 136 16242
rect 34 16233 68 16241
rect 0 16207 68 16233
rect 102 16208 136 16241
rect 102 16207 170 16208
rect 0 16198 170 16207
rect 34 16173 170 16198
rect 34 16172 136 16173
rect 34 16164 68 16172
rect 0 16138 68 16164
rect 102 16139 136 16172
rect 102 16138 170 16139
rect 0 16129 170 16138
rect 34 16104 170 16129
rect 34 16103 136 16104
rect 34 16095 68 16103
rect 0 16069 68 16095
rect 102 16070 136 16103
rect 102 16069 170 16070
rect 0 16060 170 16069
rect 34 16035 170 16060
rect 34 16034 136 16035
rect 34 16026 68 16034
rect 0 16000 68 16026
rect 102 16001 136 16034
rect 102 16000 170 16001
rect 0 15991 170 16000
rect 34 15966 170 15991
rect 34 15965 136 15966
rect 34 15957 68 15965
rect 0 15931 68 15957
rect 102 15932 136 15965
rect 102 15931 170 15932
rect 0 15922 170 15931
rect 34 15897 170 15922
rect 34 15896 136 15897
rect 34 15888 68 15896
rect 0 15862 68 15888
rect 102 15863 136 15896
rect 102 15862 170 15863
rect 0 15853 170 15862
rect 34 15828 170 15853
rect 34 15827 136 15828
rect 34 15819 68 15827
rect 0 15793 68 15819
rect 102 15794 136 15827
rect 102 15793 170 15794
rect 0 15784 170 15793
rect 34 15759 170 15784
rect 34 15758 136 15759
rect 34 15750 68 15758
rect 0 15724 68 15750
rect 102 15725 136 15758
rect 102 15724 170 15725
rect 0 15715 170 15724
rect 34 15690 170 15715
rect 34 15681 68 15690
rect 0 15646 68 15681
rect 34 15612 68 15646
rect 0 15577 68 15612
rect 34 15543 68 15577
rect 0 15508 68 15543
rect 34 15474 68 15508
rect 0 15439 68 15474
rect 34 15405 68 15439
rect 0 15370 68 15405
rect 34 15336 68 15370
rect 0 15301 68 15336
rect 34 15267 68 15301
rect 0 15232 68 15267
rect 34 15198 68 15232
rect 0 15163 68 15198
rect 34 15129 68 15163
rect 0 15094 68 15129
rect 34 15060 68 15094
rect 0 15025 68 15060
rect 34 14991 68 15025
rect 0 14956 68 14991
rect 34 14922 68 14956
rect 0 14887 68 14922
rect 34 14853 68 14887
rect 0 14818 68 14853
rect 34 14784 68 14818
rect 0 14749 68 14784
rect 34 14715 68 14749
rect 0 14680 68 14715
rect 34 14646 68 14680
rect 0 14611 68 14646
rect 34 14577 68 14611
rect 0 14542 68 14577
rect 34 14508 68 14542
rect 0 14473 68 14508
rect 34 14439 68 14473
rect 0 14404 68 14439
rect 34 14370 68 14404
rect 0 14335 68 14370
rect 34 14301 68 14335
rect 0 14266 68 14301
rect 34 14232 68 14266
rect 0 14197 68 14232
rect 34 14163 68 14197
rect 0 14128 68 14163
rect 34 14094 68 14128
rect 0 14059 68 14094
rect 34 14025 68 14059
rect 0 13990 68 14025
rect 34 13956 68 13990
rect 0 13888 170 13956
rect 34 13854 68 13888
rect 102 13854 136 13888
rect 0 13819 170 13854
rect 34 13785 68 13819
rect 102 13785 136 13819
rect 0 13750 170 13785
rect 34 13716 68 13750
rect 102 13716 136 13750
rect 0 13681 170 13716
rect 34 13647 68 13681
rect 102 13647 136 13681
rect 0 13612 170 13647
rect 34 13578 68 13612
rect 102 13578 136 13612
rect 0 13543 170 13578
rect 646 17100 748 17134
rect 13498 17100 13533 17134
rect 13567 17100 13602 17134
rect 13636 17100 13671 17134
rect 13705 17100 13740 17134
rect 13774 17100 13809 17134
rect 13843 17100 13878 17134
rect 13912 17100 13947 17134
rect 13981 17100 14016 17134
rect 14050 17100 14085 17134
rect 14119 17100 14154 17134
rect 14188 17100 14223 17134
rect 14257 17100 14292 17134
rect 14326 17100 14361 17134
rect 14395 17100 14430 17134
rect 14464 17100 14499 17134
rect 14533 17100 14568 17134
rect 14602 17100 14637 17134
rect 14671 17100 14706 17134
rect 14740 17100 14775 17134
rect 14809 17100 14844 17134
rect 14878 17100 14913 17134
rect 14947 17100 14982 17134
rect 15016 17100 15051 17134
rect 15085 17100 15120 17134
rect 15154 17100 15189 17134
rect 15223 17100 15258 17134
rect 15292 17100 15327 17134
rect 15361 17100 15396 17134
rect 15430 17100 15465 17134
rect 15499 17100 15534 17134
rect 15568 17100 15603 17134
rect 15637 17100 15672 17134
rect 15706 17100 15741 17134
rect 15775 17100 15810 17134
rect 15844 17100 15879 17134
rect 15913 17100 15948 17134
rect 15982 17100 16017 17134
rect 16051 17100 16086 17134
rect 16120 17100 16155 17134
rect 16189 17100 16224 17134
rect 16258 17100 16293 17134
rect 16327 17100 16362 17134
rect 16396 17100 16431 17134
rect 16465 17100 16500 17134
rect 16534 17100 16569 17134
rect 16603 17100 16638 17134
rect 16672 17100 16707 17134
rect 16741 17100 16776 17134
rect 16810 17100 16845 17134
rect 16879 17100 16914 17134
rect 16948 17100 16983 17134
rect 17017 17100 17052 17134
rect 17086 17100 17121 17134
rect 17155 17100 17190 17134
rect 17224 17100 17259 17134
rect 17293 17100 17328 17134
rect 17362 17100 17397 17134
rect 17431 17100 17466 17134
rect 17500 17100 17535 17134
rect 17569 17100 17604 17134
rect 17638 17100 17673 17134
rect 17707 17100 17742 17134
rect 17776 17100 17811 17134
rect 17845 17100 17880 17134
rect 17914 17100 17949 17134
rect 17983 17100 18018 17134
rect 18052 17100 18086 17134
rect 680 17066 748 17100
rect 13464 17066 18086 17100
rect 646 17032 714 17066
rect 13464 17032 13499 17066
rect 13533 17032 13568 17066
rect 13602 17032 13637 17066
rect 13671 17032 13706 17066
rect 13740 17032 13775 17066
rect 13809 17032 13844 17066
rect 13878 17032 13913 17066
rect 13947 17032 13982 17066
rect 14016 17032 14051 17066
rect 14085 17032 14120 17066
rect 14154 17032 14189 17066
rect 14223 17032 14258 17066
rect 14292 17032 14327 17066
rect 14361 17032 14396 17066
rect 14430 17032 14465 17066
rect 14499 17032 14534 17066
rect 14568 17032 14603 17066
rect 14637 17032 14672 17066
rect 14706 17032 14741 17066
rect 14775 17032 14810 17066
rect 14844 17032 14879 17066
rect 14913 17032 14948 17066
rect 14982 17032 15017 17066
rect 15051 17032 15086 17066
rect 15120 17032 15155 17066
rect 15189 17032 15224 17066
rect 15258 17032 15293 17066
rect 15327 17032 15362 17066
rect 15396 17032 15431 17066
rect 15465 17032 15500 17066
rect 15534 17032 15569 17066
rect 15603 17032 15638 17066
rect 15672 17032 15707 17066
rect 15741 17032 15776 17066
rect 15810 17032 15845 17066
rect 15879 17032 15914 17066
rect 15948 17032 15983 17066
rect 16017 17032 16052 17066
rect 16086 17032 16121 17066
rect 16155 17032 16190 17066
rect 16224 17032 16259 17066
rect 16293 17032 16328 17066
rect 16362 17032 16397 17066
rect 16431 17032 16466 17066
rect 16500 17032 16535 17066
rect 16569 17032 16604 17066
rect 16638 17032 16673 17066
rect 16707 17032 16742 17066
rect 16776 17032 16811 17066
rect 16845 17032 16880 17066
rect 16914 17032 16949 17066
rect 16983 17032 17018 17066
rect 17052 17032 17087 17066
rect 17121 17032 17156 17066
rect 17190 17032 17225 17066
rect 17259 17032 17294 17066
rect 17328 17032 17363 17066
rect 17397 17032 17432 17066
rect 17466 17032 17501 17066
rect 17535 17032 17570 17066
rect 17604 17032 17639 17066
rect 17673 17032 17708 17066
rect 17742 17032 17777 17066
rect 17811 17032 17846 17066
rect 17880 17032 17915 17066
rect 17949 17032 17984 17066
rect 18018 17032 18086 17066
rect 646 17031 782 17032
rect 680 16997 782 17031
rect 646 16963 714 16997
rect 748 16964 782 16997
rect 13396 16998 17984 17032
rect 13396 16964 13431 16998
rect 13465 16964 13500 16998
rect 13534 16964 13569 16998
rect 13603 16964 13638 16998
rect 13672 16964 13707 16998
rect 13741 16964 13776 16998
rect 13810 16964 13845 16998
rect 13879 16964 13914 16998
rect 13948 16964 13983 16998
rect 14017 16964 14052 16998
rect 14086 16964 14121 16998
rect 14155 16964 14190 16998
rect 14224 16964 14259 16998
rect 14293 16964 14328 16998
rect 14362 16964 14397 16998
rect 14431 16964 14466 16998
rect 14500 16964 14535 16998
rect 14569 16964 14604 16998
rect 14638 16964 14673 16998
rect 14707 16964 14742 16998
rect 14776 16964 14811 16998
rect 14845 16964 14880 16998
rect 14914 16964 14949 16998
rect 14983 16964 15018 16998
rect 15052 16964 15087 16998
rect 15121 16964 15156 16998
rect 15190 16964 15225 16998
rect 15259 16964 15294 16998
rect 15328 16964 15363 16998
rect 15397 16964 15432 16998
rect 15466 16964 15501 16998
rect 15535 16964 15570 16998
rect 15604 16964 15639 16998
rect 15673 16964 15708 16998
rect 15742 16964 15777 16998
rect 15811 16964 15846 16998
rect 15880 16964 15915 16998
rect 15949 16964 15984 16998
rect 16018 16964 16053 16998
rect 16087 16964 16122 16998
rect 16156 16964 16191 16998
rect 16225 16964 16260 16998
rect 16294 16964 16329 16998
rect 16363 16964 16398 16998
rect 16432 16964 16467 16998
rect 16501 16964 16536 16998
rect 16570 16964 16605 16998
rect 16639 16964 16674 16998
rect 16708 16964 16743 16998
rect 16777 16964 16812 16998
rect 16846 16964 16881 16998
rect 16915 16964 16950 16998
rect 16984 16964 17019 16998
rect 17053 16964 17088 16998
rect 17122 16964 17157 16998
rect 17191 16964 17226 16998
rect 17260 16964 17295 16998
rect 17329 16964 17364 16998
rect 17398 16964 17433 16998
rect 17467 16964 17502 16998
rect 17536 16964 17571 16998
rect 17605 16964 17640 16998
rect 17674 16964 17709 16998
rect 17743 16964 17778 16998
rect 17812 16964 17847 16998
rect 17881 16964 17916 16998
rect 748 16963 816 16964
rect 646 16962 816 16963
rect 680 16929 816 16962
rect 680 16928 782 16929
rect 646 16894 714 16928
rect 748 16895 782 16928
rect 748 16894 816 16895
rect 646 16893 816 16894
rect 680 16860 816 16893
rect 680 16859 782 16860
rect 646 16825 714 16859
rect 748 16826 782 16859
rect 748 16825 816 16826
rect 646 16824 816 16825
rect 680 16791 816 16824
rect 680 16790 782 16791
rect 646 16756 714 16790
rect 748 16757 782 16790
rect 748 16756 816 16757
rect 646 16755 816 16756
rect 680 16722 816 16755
rect 10431 16930 15650 16964
rect 10431 16896 10494 16930
rect 10528 16896 10563 16930
rect 10597 16896 10632 16930
rect 10666 16896 10701 16930
rect 10735 16896 10770 16930
rect 10804 16896 10839 16930
rect 10873 16896 10908 16930
rect 10942 16896 10977 16930
rect 11011 16896 11046 16930
rect 11080 16896 11115 16930
rect 11149 16896 11184 16930
rect 11218 16896 11253 16930
rect 11287 16896 11322 16930
rect 11356 16896 11391 16930
rect 11425 16896 11460 16930
rect 11494 16896 11529 16930
rect 11563 16896 11598 16930
rect 11632 16896 11667 16930
rect 11701 16896 11736 16930
rect 11770 16896 11805 16930
rect 11839 16896 11874 16930
rect 11908 16896 11943 16930
rect 11977 16896 12012 16930
rect 12046 16896 12081 16930
rect 12115 16896 12150 16930
rect 12184 16896 12219 16930
rect 12253 16896 12288 16930
rect 12322 16896 12357 16930
rect 12391 16896 12426 16930
rect 12460 16896 12495 16930
rect 12529 16896 12564 16930
rect 12598 16896 12633 16930
rect 12667 16896 12702 16930
rect 12736 16896 12771 16930
rect 12805 16896 12840 16930
rect 12874 16896 12909 16930
rect 12943 16896 12978 16930
rect 13012 16896 13047 16930
rect 13081 16896 13116 16930
rect 13150 16896 13185 16930
rect 13219 16896 13254 16930
rect 13288 16896 13323 16930
rect 13357 16896 13392 16930
rect 13426 16896 13461 16930
rect 13495 16896 13530 16930
rect 13564 16896 13599 16930
rect 13633 16896 13668 16930
rect 13702 16896 13737 16930
rect 13771 16896 13806 16930
rect 13840 16896 13875 16930
rect 13909 16896 13944 16930
rect 13978 16896 14013 16930
rect 14047 16896 14082 16930
rect 14116 16896 14151 16930
rect 14185 16896 14220 16930
rect 14254 16896 14289 16930
rect 14323 16896 14358 16930
rect 14392 16896 14427 16930
rect 14461 16896 14496 16930
rect 10431 16862 14496 16896
rect 10431 16828 10494 16862
rect 10528 16828 10563 16862
rect 10597 16828 10632 16862
rect 10666 16828 10701 16862
rect 10735 16828 10770 16862
rect 10804 16828 10839 16862
rect 10873 16828 10908 16862
rect 10942 16828 10977 16862
rect 11011 16828 11046 16862
rect 11080 16828 11115 16862
rect 11149 16828 11184 16862
rect 11218 16828 11253 16862
rect 11287 16828 11322 16862
rect 11356 16828 11391 16862
rect 11425 16828 11460 16862
rect 11494 16828 11529 16862
rect 11563 16828 11598 16862
rect 11632 16828 11667 16862
rect 11701 16828 11736 16862
rect 11770 16828 11805 16862
rect 11839 16828 11874 16862
rect 11908 16828 11943 16862
rect 11977 16828 12012 16862
rect 12046 16828 12081 16862
rect 12115 16828 12150 16862
rect 12184 16828 12219 16862
rect 12253 16828 12288 16862
rect 12322 16828 12357 16862
rect 12391 16828 12426 16862
rect 12460 16828 12495 16862
rect 12529 16828 12564 16862
rect 12598 16828 12633 16862
rect 12667 16828 12702 16862
rect 12736 16828 12771 16862
rect 12805 16828 12840 16862
rect 12874 16828 12909 16862
rect 12943 16828 12978 16862
rect 13012 16828 13047 16862
rect 13081 16828 13116 16862
rect 13150 16828 13185 16862
rect 13219 16828 13254 16862
rect 13288 16828 13323 16862
rect 13357 16828 13392 16862
rect 13426 16828 13461 16862
rect 13495 16828 13530 16862
rect 13564 16828 13599 16862
rect 13633 16828 13668 16862
rect 13702 16828 13737 16862
rect 13771 16828 13806 16862
rect 13840 16828 13875 16862
rect 13909 16828 13944 16862
rect 13978 16828 14013 16862
rect 14047 16828 14082 16862
rect 14116 16828 14151 16862
rect 14185 16828 14220 16862
rect 14254 16828 14289 16862
rect 14323 16828 14358 16862
rect 14392 16828 14427 16862
rect 14461 16828 14496 16862
rect 10431 16794 14496 16828
rect 10431 16760 10494 16794
rect 10528 16760 10563 16794
rect 10597 16760 10632 16794
rect 10666 16760 10701 16794
rect 10735 16760 10770 16794
rect 10804 16760 10839 16794
rect 10873 16760 10908 16794
rect 10942 16760 10977 16794
rect 11011 16760 11046 16794
rect 11080 16760 11115 16794
rect 11149 16760 11184 16794
rect 11218 16760 11253 16794
rect 11287 16760 11322 16794
rect 11356 16760 11391 16794
rect 11425 16760 11460 16794
rect 11494 16760 11529 16794
rect 11563 16760 11598 16794
rect 11632 16760 11667 16794
rect 11701 16760 11736 16794
rect 11770 16760 11805 16794
rect 11839 16760 11874 16794
rect 11908 16760 11943 16794
rect 11977 16760 12012 16794
rect 12046 16760 12081 16794
rect 12115 16760 12150 16794
rect 12184 16760 12219 16794
rect 12253 16760 12288 16794
rect 12322 16760 12357 16794
rect 12391 16760 12426 16794
rect 12460 16760 12495 16794
rect 12529 16760 12564 16794
rect 12598 16760 12633 16794
rect 12667 16760 12702 16794
rect 12736 16760 12771 16794
rect 12805 16760 12840 16794
rect 12874 16760 12909 16794
rect 12943 16760 12978 16794
rect 13012 16760 13047 16794
rect 13081 16760 13116 16794
rect 13150 16760 13185 16794
rect 13219 16760 13254 16794
rect 13288 16760 13323 16794
rect 13357 16760 13392 16794
rect 13426 16760 13461 16794
rect 13495 16760 13530 16794
rect 13564 16760 13599 16794
rect 13633 16760 13668 16794
rect 13702 16760 13737 16794
rect 13771 16760 13806 16794
rect 13840 16760 13875 16794
rect 13909 16760 13944 16794
rect 13978 16760 14013 16794
rect 14047 16760 14082 16794
rect 14116 16760 14151 16794
rect 14185 16760 14220 16794
rect 14254 16760 14289 16794
rect 14323 16760 14358 16794
rect 14392 16760 14427 16794
rect 14461 16760 14496 16794
rect 15210 16760 15260 16930
rect 10431 16744 15260 16760
rect 680 16721 782 16722
rect 646 16687 714 16721
rect 748 16688 782 16721
rect 748 16687 816 16688
rect 646 16686 816 16687
rect 680 16653 816 16686
rect 680 16652 782 16653
rect 646 16618 714 16652
rect 748 16619 782 16652
rect 748 16618 816 16619
rect 646 16617 816 16618
rect 680 16584 816 16617
rect 680 16583 782 16584
rect 646 16549 714 16583
rect 748 16550 782 16583
rect 748 16549 816 16550
rect 646 16548 816 16549
rect 680 16515 816 16548
rect 680 16514 782 16515
rect 646 16480 714 16514
rect 748 16481 782 16514
rect 748 16480 816 16481
rect 646 16479 816 16480
rect 680 16446 816 16479
rect 680 16445 782 16446
rect 646 16411 714 16445
rect 748 16412 782 16445
rect 748 16411 816 16412
rect 646 16410 816 16411
rect 680 16377 816 16410
rect 680 16376 782 16377
rect 646 16342 714 16376
rect 748 16343 782 16376
rect 748 16342 816 16343
rect 646 16341 816 16342
rect 680 16308 816 16341
rect 680 16307 782 16308
rect 748 16274 782 16307
rect 748 16239 816 16274
rect 15071 16007 15260 16744
rect 15181 15113 15260 16007
rect 15082 14788 15260 15113
rect 15430 16904 15650 16930
rect 15430 16870 15464 16904
rect 15498 16870 15532 16904
rect 15566 16870 15600 16904
rect 15634 16870 15650 16904
rect 15430 16832 15650 16870
rect 15430 16798 15464 16832
rect 15498 16798 15532 16832
rect 15566 16798 15600 16832
rect 15634 16798 15650 16832
rect 15430 16760 15650 16798
rect 15430 16726 15464 16760
rect 15498 16726 15532 16760
rect 15566 16726 15600 16760
rect 15634 16726 15650 16760
rect 15430 16688 15650 16726
rect 15430 16654 15464 16688
rect 15498 16654 15532 16688
rect 15566 16654 15600 16688
rect 15634 16654 15650 16688
rect 15430 16616 15650 16654
rect 15430 16582 15464 16616
rect 15498 16582 15532 16616
rect 15566 16582 15600 16616
rect 15634 16582 15650 16616
rect 15430 16544 15650 16582
rect 15430 16510 15464 16544
rect 15498 16510 15532 16544
rect 15566 16510 15600 16544
rect 15634 16510 15650 16544
rect 15430 16472 15650 16510
rect 15430 16438 15464 16472
rect 15498 16438 15532 16472
rect 15566 16438 15600 16472
rect 15634 16438 15650 16472
rect 15430 16400 15650 16438
rect 15430 16366 15464 16400
rect 15498 16366 15532 16400
rect 15566 16366 15600 16400
rect 15634 16366 15650 16400
rect 15430 16328 15650 16366
rect 15430 16294 15464 16328
rect 15498 16294 15532 16328
rect 15566 16294 15600 16328
rect 15634 16294 15650 16328
rect 15430 16255 15650 16294
rect 15430 16221 15464 16255
rect 15498 16221 15532 16255
rect 15566 16221 15600 16255
rect 15634 16221 15650 16255
rect 15430 16132 15650 16221
rect 17916 16590 18052 16624
rect 17916 16589 18086 16590
rect 17950 16555 17984 16589
rect 18018 16556 18086 16589
rect 18018 16555 18052 16556
rect 17916 16522 18052 16555
rect 17916 16520 18086 16522
rect 17950 16486 17984 16520
rect 18018 16488 18086 16520
rect 18018 16486 18052 16488
rect 17916 16454 18052 16486
rect 17916 16451 18086 16454
rect 17950 16417 17984 16451
rect 18018 16420 18086 16451
rect 18018 16417 18052 16420
rect 17916 16386 18052 16417
rect 17916 16382 18086 16386
rect 17950 16348 17984 16382
rect 18018 16352 18086 16382
rect 18018 16348 18052 16352
rect 17916 16318 18052 16348
rect 17916 16313 18086 16318
rect 17950 16279 17984 16313
rect 18018 16284 18086 16313
rect 18018 16279 18052 16284
rect 17916 16250 18052 16279
rect 17916 16244 18086 16250
rect 17950 16210 17984 16244
rect 18018 16216 18086 16244
rect 18018 16210 18052 16216
rect 17916 16182 18052 16210
rect 17916 16175 18086 16182
rect 17950 16141 17984 16175
rect 18018 16148 18086 16175
rect 18018 16141 18052 16148
rect 15430 14788 15582 16132
rect 17916 16114 18052 16141
rect 17916 16106 18086 16114
rect 17950 16072 17984 16106
rect 18018 16080 18086 16106
rect 18018 16072 18052 16080
rect 17916 16046 18052 16072
rect 17916 16037 18086 16046
rect 17950 16003 17984 16037
rect 18018 16012 18086 16037
rect 18018 16003 18052 16012
rect 17916 15978 18052 16003
rect 17916 15968 18086 15978
rect 17950 15934 17984 15968
rect 18018 15944 18086 15968
rect 18018 15934 18052 15944
rect 17916 15910 18052 15934
rect 17916 15899 18086 15910
rect 17950 15865 17984 15899
rect 18018 15876 18086 15899
rect 18018 15865 18052 15876
rect 17916 15842 18052 15865
rect 17916 15830 18086 15842
rect 17950 15796 17984 15830
rect 18018 15808 18086 15830
rect 18018 15796 18052 15808
rect 17916 15774 18052 15796
rect 17916 15761 18086 15774
rect 17950 15727 17984 15761
rect 18018 15740 18086 15761
rect 18018 15727 18052 15740
rect 17916 15706 18052 15727
rect 17916 15692 18086 15706
rect 17950 15658 17984 15692
rect 18018 15672 18086 15692
rect 18018 15658 18052 15672
rect 17916 15638 18052 15658
rect 17916 15623 18086 15638
rect 17950 15589 17984 15623
rect 18018 15604 18086 15623
rect 18018 15589 18052 15604
rect 17916 15570 18052 15589
rect 17916 15554 18086 15570
rect 17950 15520 17984 15554
rect 18018 15536 18086 15554
rect 18018 15520 18052 15536
rect 17916 15502 18052 15520
rect 17916 15485 18086 15502
rect 17950 15451 17984 15485
rect 18018 15468 18086 15485
rect 18018 15451 18052 15468
rect 17916 15434 18052 15451
rect 17916 15416 18086 15434
rect 17950 15382 17984 15416
rect 18018 15400 18086 15416
rect 18018 15382 18052 15400
rect 17916 15366 18052 15382
rect 17916 15347 18086 15366
rect 17950 15313 17984 15347
rect 18018 15332 18086 15347
rect 18018 15313 18052 15332
rect 17916 15298 18052 15313
rect 17916 15278 18086 15298
rect 17950 15244 17984 15278
rect 18018 15264 18086 15278
rect 18018 15244 18052 15264
rect 17916 15230 18052 15244
rect 17916 15209 18086 15230
rect 17950 15175 17984 15209
rect 18018 15196 18086 15209
rect 18018 15175 18052 15196
rect 17916 15162 18052 15175
rect 17916 15140 18086 15162
rect 17950 15106 17984 15140
rect 18018 15128 18086 15140
rect 18018 15106 18052 15128
rect 17916 15094 18052 15106
rect 17916 15071 18086 15094
rect 17950 15037 17984 15071
rect 18018 15060 18086 15071
rect 18018 15037 18052 15060
rect 17916 15026 18052 15037
rect 17916 15002 18086 15026
rect 15082 14753 15582 14788
rect 15082 14719 15260 14753
rect 15294 14719 15328 14753
rect 15362 14719 15396 14753
rect 15430 14719 15582 14753
rect 17950 14968 17984 15002
rect 18018 14992 18086 15002
rect 18018 14968 18052 14992
rect 17916 14958 18052 14968
rect 17916 14933 18086 14958
rect 17950 14899 17984 14933
rect 18018 14924 18086 14933
rect 18018 14899 18052 14924
rect 17916 14890 18052 14899
rect 17916 14864 18086 14890
rect 17950 14830 17984 14864
rect 18018 14856 18086 14864
rect 18018 14830 18052 14856
rect 17916 14822 18052 14830
rect 17916 14795 18086 14822
rect 17950 14761 17984 14795
rect 18018 14788 18086 14795
rect 18018 14761 18052 14788
rect 17916 14754 18052 14761
rect 17916 14726 18086 14754
rect 15082 14684 15582 14719
rect 15082 14650 15260 14684
rect 15294 14650 15328 14684
rect 15362 14650 15396 14684
rect 15430 14650 15582 14684
rect 15082 14615 15582 14650
rect 15082 14581 15260 14615
rect 15294 14581 15328 14615
rect 15362 14581 15396 14615
rect 15430 14581 15582 14615
rect 15082 14546 15582 14581
rect 15082 14512 15260 14546
rect 15294 14512 15328 14546
rect 15362 14512 15396 14546
rect 15430 14512 15582 14546
rect 15082 14477 15582 14512
rect 15082 14443 15260 14477
rect 15294 14443 15328 14477
rect 15362 14443 15396 14477
rect 15430 14443 15582 14477
rect 15082 14408 15582 14443
rect 15082 14374 15260 14408
rect 15294 14374 15328 14408
rect 15362 14374 15396 14408
rect 15430 14374 15582 14408
rect 15082 14340 15582 14374
rect 15082 14306 15396 14340
rect 15430 14306 15582 14340
rect 15082 14269 15582 14306
rect 15082 14235 15396 14269
rect 15430 14235 15582 14269
rect 15082 14198 15582 14235
rect 15082 14164 15396 14198
rect 15430 14164 15582 14198
rect 15082 14127 15582 14164
rect 15082 14093 15396 14127
rect 15430 14093 15582 14127
rect 15082 14056 15582 14093
rect 15082 14022 15396 14056
rect 15430 14022 15582 14056
rect 15082 13985 15582 14022
rect 15082 13951 15396 13985
rect 15430 13951 15582 13985
rect 15082 13914 15582 13951
rect 15082 13893 15396 13914
rect 15161 13880 15396 13893
rect 15430 13880 15582 13914
rect 15161 13843 15582 13880
rect 15161 13809 15396 13843
rect 15430 13809 15582 13843
rect 15161 13772 15582 13809
rect 15161 13738 15396 13772
rect 15430 13738 15582 13772
rect 15161 13701 15582 13738
rect 15161 13667 15396 13701
rect 15430 13667 15582 13701
rect 15161 13630 15582 13667
rect 15161 13596 15396 13630
rect 15430 13596 15582 13630
rect 17950 14692 17984 14726
rect 18018 14720 18086 14726
rect 18018 14692 18052 14720
rect 17916 14686 18052 14692
rect 17916 14657 18086 14686
rect 17950 14623 17984 14657
rect 18018 14652 18086 14657
rect 18018 14623 18052 14652
rect 17916 14618 18052 14623
rect 17916 14588 18086 14618
rect 17950 14554 17984 14588
rect 18018 14584 18086 14588
rect 18018 14554 18052 14584
rect 17916 14550 18052 14554
rect 17916 14519 18086 14550
rect 17950 14485 17984 14519
rect 18018 14516 18086 14519
rect 18018 14485 18052 14516
rect 17916 14482 18052 14485
rect 17916 14450 18086 14482
rect 17950 14416 17984 14450
rect 18018 14448 18086 14450
rect 18018 14416 18052 14448
rect 17916 14414 18052 14416
rect 17916 14381 18086 14414
rect 17950 14347 17984 14381
rect 18018 14380 18086 14381
rect 18018 14347 18052 14380
rect 17916 14346 18052 14347
rect 17916 14312 18086 14346
rect 17950 14278 17984 14312
rect 18018 14278 18052 14312
rect 17916 14243 18086 14278
rect 17950 14209 17984 14243
rect 18018 14209 18052 14243
rect 17916 14174 18086 14209
rect 17950 14140 17984 14174
rect 18018 14140 18052 14174
rect 17916 14105 18086 14140
rect 17950 14071 17984 14105
rect 18018 14071 18052 14105
rect 17916 14036 18086 14071
rect 17950 14002 17984 14036
rect 18018 14002 18052 14036
rect 17916 13967 18086 14002
rect 17950 13933 17984 13967
rect 18018 13933 18052 13967
rect 17916 13898 18086 13933
rect 17950 13864 17984 13898
rect 18018 13864 18052 13898
rect 17916 13829 18086 13864
rect 17950 13795 17984 13829
rect 18018 13795 18052 13829
rect 17916 13760 18086 13795
rect 17950 13726 17984 13760
rect 18018 13726 18052 13760
rect 17916 13691 18086 13726
rect 17950 13657 17984 13691
rect 18018 13657 18052 13691
rect 15161 13559 15582 13596
rect 15161 13525 15396 13559
rect 15430 13525 15582 13559
rect 15161 13488 15582 13525
rect 15161 13454 15396 13488
rect 15430 13454 15582 13488
rect 15161 13417 15582 13454
rect 15161 13383 15396 13417
rect 15430 13383 15582 13417
rect 15161 13346 15582 13383
rect 17916 13622 18086 13657
rect 17950 13588 17984 13622
rect 18018 13588 18052 13622
rect 17916 13553 18086 13588
rect 17950 13519 17984 13553
rect 18018 13519 18052 13553
rect 17916 13484 18086 13519
rect 17950 13450 17984 13484
rect 18018 13450 18052 13484
rect 17916 13415 18086 13450
rect 17950 13381 17984 13415
rect 18018 13381 18052 13415
rect 15161 13312 15396 13346
rect 15430 13312 15582 13346
rect 15161 13275 15582 13312
rect 15161 13267 15396 13275
rect 15278 13241 15396 13267
rect 15430 13241 15582 13275
rect 15278 12975 15582 13241
rect 17916 13346 18086 13381
rect 17950 13312 17984 13346
rect 18018 13312 18052 13346
rect 17916 13277 18086 13312
rect 17950 13243 17984 13277
rect 18018 13243 18052 13277
rect 17916 13208 18086 13243
rect 17950 13174 17984 13208
rect 18018 13174 18052 13208
rect 17916 13139 18086 13174
rect 17950 13105 17984 13139
rect 18018 13105 18052 13139
rect 17916 13070 18086 13105
rect 17950 13036 17984 13070
rect 18018 13036 18052 13070
rect 17916 13001 18086 13036
rect 816 12941 851 12975
rect 885 12941 920 12975
rect 954 12941 989 12975
rect 1023 12941 1058 12975
rect 1092 12941 1127 12975
rect 1161 12941 1196 12975
rect 1230 12941 1265 12975
rect 1299 12941 1334 12975
rect 1368 12941 1403 12975
rect 1437 12941 1472 12975
rect 1506 12941 1541 12975
rect 1575 12941 1610 12975
rect 1644 12941 1679 12975
rect 1713 12941 1748 12975
rect 1782 12941 1817 12975
rect 1851 12941 1886 12975
rect 1920 12941 1955 12975
rect 1989 12941 2024 12975
rect 2058 12941 2093 12975
rect 2127 12941 2162 12975
rect 2196 12941 2231 12975
rect 2265 12941 2300 12975
rect 2334 12941 2369 12975
rect 2403 12941 2438 12975
rect 748 12907 2438 12941
rect 646 12873 714 12907
rect 748 12873 783 12907
rect 817 12873 852 12907
rect 886 12873 921 12907
rect 955 12873 990 12907
rect 1024 12873 1059 12907
rect 1093 12873 1128 12907
rect 1162 12873 1197 12907
rect 1231 12873 1266 12907
rect 1300 12873 1335 12907
rect 1369 12873 1404 12907
rect 1438 12873 1473 12907
rect 1507 12873 1542 12907
rect 1576 12873 1611 12907
rect 1645 12873 1680 12907
rect 1714 12873 1749 12907
rect 1783 12873 1818 12907
rect 1852 12873 1887 12907
rect 1921 12873 1956 12907
rect 1990 12873 2025 12907
rect 2059 12873 2094 12907
rect 2128 12873 2163 12907
rect 2197 12873 2232 12907
rect 2266 12873 2301 12907
rect 2335 12873 2370 12907
rect 2404 12873 2438 12907
rect 17840 12967 17916 12975
rect 17950 12967 17984 13001
rect 18018 12967 18052 13001
rect 17840 12932 18086 12967
rect 17840 12898 17916 12932
rect 17950 12898 17984 12932
rect 18018 12898 18052 12932
rect 646 12839 4682 12873
rect 646 12805 680 12839
rect 714 12805 749 12839
rect 783 12805 818 12839
rect 852 12805 887 12839
rect 921 12805 956 12839
rect 990 12805 1025 12839
rect 1059 12805 1094 12839
rect 1128 12805 1163 12839
rect 1197 12805 1232 12839
rect 1266 12805 1301 12839
rect 1335 12805 1370 12839
rect 1404 12805 1439 12839
rect 1473 12805 1508 12839
rect 1542 12805 1577 12839
rect 1611 12805 1646 12839
rect 1680 12805 1715 12839
rect 1749 12805 1784 12839
rect 1818 12805 1853 12839
rect 1887 12805 1922 12839
rect 1956 12805 1991 12839
rect 2025 12805 2060 12839
rect 2094 12805 2129 12839
rect 2163 12805 2198 12839
rect 2232 12805 2267 12839
rect 2301 12805 2336 12839
rect 2370 12805 2405 12839
rect 2439 12805 2474 12839
rect 2508 12805 2543 12839
rect 2577 12805 2612 12839
rect 2646 12805 2681 12839
rect 2715 12805 2750 12839
rect 2784 12805 2819 12839
rect 2853 12805 2888 12839
rect 2922 12805 2957 12839
rect 2991 12805 3026 12839
rect 3060 12805 3095 12839
rect 3129 12805 3164 12839
rect 3198 12805 3233 12839
rect 3267 12805 3302 12839
rect 3336 12805 3371 12839
rect 3405 12805 3440 12839
rect 3474 12805 3509 12839
rect 3543 12805 3578 12839
rect 3612 12805 3647 12839
rect 3681 12805 3716 12839
rect 3750 12805 3785 12839
rect 3819 12805 3854 12839
rect 3888 12805 3923 12839
rect 3957 12805 3992 12839
rect 4026 12805 4061 12839
rect 4095 12805 4130 12839
rect 4164 12805 4199 12839
rect 4233 12805 4268 12839
rect 4302 12805 4337 12839
rect 4371 12805 4406 12839
rect 4440 12805 4475 12839
rect 4509 12805 4544 12839
rect 4578 12805 4613 12839
rect 4647 12805 4682 12839
rect 17840 12863 18086 12898
rect 17840 12829 17916 12863
rect 17950 12829 17984 12863
rect 18018 12829 18052 12863
rect 17840 12805 18086 12829
rect 0 12249 170 12285
rect 18609 12318 18677 12353
rect 18643 12285 18677 12318
rect 18643 12284 18745 12285
rect 18609 12251 18745 12284
rect 18609 12250 18779 12251
rect 18609 12249 18677 12250
rect 0 12215 18124 12249
rect 18158 12215 18194 12249
rect 18228 12215 18264 12249
rect 18298 12215 18333 12249
rect 18367 12215 18402 12249
rect 18436 12215 18471 12249
rect 18505 12215 18540 12249
rect 18574 12215 18609 12249
rect 18643 12216 18677 12249
rect 18711 12216 18779 12250
rect 18643 12215 18745 12216
rect 0 12182 18745 12215
rect 0 12181 18779 12182
rect 0 12147 18124 12181
rect 18158 12147 18194 12181
rect 18228 12147 18263 12181
rect 18297 12147 18332 12181
rect 18366 12147 18401 12181
rect 18435 12147 18470 12181
rect 18504 12147 18539 12181
rect 18573 12147 18608 12181
rect 18642 12147 18677 12181
rect 18711 12147 18779 12181
rect 0 12113 18745 12147
rect 0 12079 18124 12113
rect 18158 12079 18197 12113
rect 18231 12079 18270 12113
rect 18304 12079 18343 12113
rect 18377 12079 18416 12113
rect 18450 12079 18489 12113
rect 18523 12079 18562 12113
rect 18596 12079 18635 12113
rect 18669 12079 18779 12113
rect 11972 7691 12142 12079
rect 17920 7691 18090 12079
rect 11972 7521 18090 7691
<< mvpsubdiff >>
rect 10491 3380 10737 3404
rect 10525 3346 10559 3380
rect 10593 3346 10627 3380
rect 10661 3346 10737 3380
rect 10491 3311 10737 3346
rect 10491 3310 10559 3311
rect 10525 3277 10559 3310
rect 10593 3277 10627 3311
rect 10661 3277 10737 3311
rect 12267 3370 12301 3404
rect 12335 3370 12369 3404
rect 12403 3370 12437 3404
rect 12471 3370 12505 3404
rect 12539 3370 12573 3404
rect 12607 3370 12641 3404
rect 12675 3370 12709 3404
rect 12743 3370 12777 3404
rect 12811 3370 12845 3404
rect 12879 3370 12913 3404
rect 12947 3370 12981 3404
rect 13015 3370 13049 3404
rect 13083 3370 13117 3404
rect 13151 3370 13185 3404
rect 13219 3370 13253 3404
rect 13287 3370 13321 3404
rect 13355 3370 13389 3404
rect 13423 3370 13457 3404
rect 13491 3370 13525 3404
rect 13559 3370 13593 3404
rect 13627 3370 13661 3404
rect 13695 3370 13729 3404
rect 13763 3370 13797 3404
rect 13831 3370 13865 3404
rect 13899 3370 13933 3404
rect 13967 3370 14001 3404
rect 14035 3370 14069 3404
rect 14103 3370 14137 3404
rect 14171 3370 14205 3404
rect 14239 3370 14273 3404
rect 14307 3370 14341 3404
rect 14375 3370 14409 3404
rect 14443 3370 14477 3404
rect 14511 3370 14545 3404
rect 14579 3370 14613 3404
rect 14647 3370 14682 3404
rect 14716 3370 14751 3404
rect 14785 3370 14820 3404
rect 14854 3370 14889 3404
rect 14923 3370 14958 3404
rect 14992 3370 15027 3404
rect 15061 3370 15096 3404
rect 15130 3370 15165 3404
rect 15199 3370 15234 3404
rect 15268 3370 15303 3404
rect 15337 3370 15372 3404
rect 15406 3370 15441 3404
rect 15475 3370 15509 3404
rect 12267 3336 15509 3370
rect 12267 3302 12302 3336
rect 12336 3302 12371 3336
rect 12405 3302 12440 3336
rect 12474 3302 12509 3336
rect 12543 3302 12578 3336
rect 12612 3302 12647 3336
rect 12681 3302 12716 3336
rect 12750 3302 12785 3336
rect 12819 3302 12854 3336
rect 12888 3302 12923 3336
rect 12957 3302 12992 3336
rect 13026 3302 13061 3336
rect 13095 3302 13130 3336
rect 13164 3302 13199 3336
rect 13233 3302 13268 3336
rect 13302 3302 13337 3336
rect 13371 3302 13406 3336
rect 13440 3302 13475 3336
rect 13509 3302 13544 3336
rect 13578 3302 13613 3336
rect 13647 3302 13682 3336
rect 13716 3302 13751 3336
rect 13785 3302 13820 3336
rect 13854 3302 13889 3336
rect 13923 3302 13958 3336
rect 13992 3302 14027 3336
rect 14061 3302 14096 3336
rect 14130 3302 14165 3336
rect 14199 3302 14234 3336
rect 14268 3302 14303 3336
rect 14337 3302 14372 3336
rect 14406 3302 14441 3336
rect 14475 3302 14510 3336
rect 14544 3302 14579 3336
rect 14613 3302 14648 3336
rect 14682 3302 14717 3336
rect 14751 3302 14786 3336
rect 14820 3302 14855 3336
rect 14889 3302 14924 3336
rect 14958 3302 14993 3336
rect 15027 3302 15062 3336
rect 15096 3302 15131 3336
rect 15165 3302 15200 3336
rect 15234 3302 15269 3336
rect 15303 3302 15338 3336
rect 15372 3302 15407 3336
rect 15441 3302 15509 3336
rect 10525 3276 10737 3277
rect 10491 3242 10737 3276
rect 10491 3240 10559 3242
rect 10525 3208 10559 3240
rect 10593 3208 10627 3242
rect 10661 3234 10737 3242
rect 12199 3300 15509 3302
rect 12199 3268 15475 3300
rect 12199 3234 12234 3268
rect 12268 3234 12303 3268
rect 12337 3234 12372 3268
rect 12406 3234 12441 3268
rect 12475 3234 12510 3268
rect 12544 3234 12579 3268
rect 12613 3234 12648 3268
rect 12682 3234 12717 3268
rect 12751 3234 12786 3268
rect 12820 3234 12855 3268
rect 12889 3234 12924 3268
rect 12958 3234 12993 3268
rect 13027 3234 13062 3268
rect 13096 3234 13131 3268
rect 13165 3234 13200 3268
rect 13234 3234 13269 3268
rect 13303 3234 13338 3268
rect 13372 3234 13407 3268
rect 13441 3234 13476 3268
rect 13510 3234 13545 3268
rect 13579 3234 13614 3268
rect 13648 3234 13683 3268
rect 13717 3234 13752 3268
rect 13786 3234 13821 3268
rect 13855 3234 13890 3268
rect 13924 3234 13959 3268
rect 13993 3234 14028 3268
rect 14062 3234 14097 3268
rect 14131 3234 14166 3268
rect 14200 3234 14235 3268
rect 14269 3234 14304 3268
rect 14338 3234 14373 3268
rect 14407 3234 14442 3268
rect 14476 3234 14511 3268
rect 14545 3234 14580 3268
rect 14614 3234 14649 3268
rect 14683 3234 14718 3268
rect 14752 3234 14787 3268
rect 14821 3234 14856 3268
rect 14890 3234 14925 3268
rect 14959 3234 14994 3268
rect 15028 3234 15063 3268
rect 15097 3234 15132 3268
rect 15166 3234 15201 3268
rect 15235 3234 15270 3268
rect 15304 3234 15339 3268
rect 15373 3267 15475 3268
rect 15373 3234 15407 3267
rect 10525 3206 10661 3208
rect 10491 3173 10661 3206
rect 10491 3170 10559 3173
rect 10525 3139 10559 3170
rect 10593 3139 10627 3173
rect 10525 3136 10661 3139
rect 10491 3104 10661 3136
rect 10491 3100 10559 3104
rect 10525 3070 10559 3100
rect 10593 3070 10627 3104
rect 10525 3066 10661 3070
rect 10491 3035 10661 3066
rect 10491 3030 10559 3035
rect 10525 3001 10559 3030
rect 10593 3001 10627 3035
rect 10525 2996 10661 3001
rect 10491 2966 10661 2996
rect 10491 2960 10559 2966
rect 10525 2932 10559 2960
rect 10593 2932 10627 2966
rect 10525 2926 10661 2932
rect 10491 2897 10661 2926
rect 10491 2890 10559 2897
rect 10525 2863 10559 2890
rect 10593 2863 10627 2897
rect 10525 2856 10661 2863
rect 10491 2828 10661 2856
rect 10491 2820 10559 2828
rect 10525 2794 10559 2820
rect 10593 2794 10627 2828
rect 10525 2786 10661 2794
rect 10491 2759 10661 2786
rect 10491 2750 10559 2759
rect 10525 2725 10559 2750
rect 10593 2725 10627 2759
rect 10525 2716 10661 2725
rect 10491 2690 10661 2716
rect 10491 2680 10559 2690
rect 10525 2656 10559 2680
rect 10593 2656 10627 2690
rect 10525 2646 10661 2656
rect 10491 2621 10661 2646
rect 10491 2610 10559 2621
rect 10525 2587 10559 2610
rect 10593 2587 10627 2621
rect 10525 2576 10661 2587
rect 10491 2552 10661 2576
rect 10491 2540 10559 2552
rect 10525 2518 10559 2540
rect 10593 2518 10627 2552
rect 10525 2506 10661 2518
rect 10491 2483 10661 2506
rect 10491 2470 10559 2483
rect 10525 2449 10559 2470
rect 10593 2449 10627 2483
rect 10525 2436 10661 2449
rect 10491 2414 10661 2436
rect 10491 2400 10559 2414
rect 10525 2380 10559 2400
rect 10593 2380 10627 2414
rect 10525 2366 10661 2380
rect 10491 2345 10661 2366
rect 10491 2330 10559 2345
rect 10525 2311 10559 2330
rect 10593 2311 10627 2345
rect 10525 2296 10661 2311
rect 10491 2276 10661 2296
rect 10491 2260 10559 2276
rect 10525 2242 10559 2260
rect 10593 2242 10627 2276
rect 10525 2226 10661 2242
rect 10491 2207 10661 2226
rect 10491 2190 10559 2207
rect 10525 2173 10559 2190
rect 10593 2173 10627 2207
rect 10525 2156 10661 2173
rect 10491 2138 10661 2156
rect 10491 2120 10559 2138
rect 10525 2104 10559 2120
rect 10593 2104 10627 2138
rect 10525 2086 10661 2104
rect 10491 2069 10661 2086
rect 10491 2050 10559 2069
rect 10525 2035 10559 2050
rect 10593 2035 10627 2069
rect 10525 2016 10661 2035
rect 10491 2000 10661 2016
rect 10491 1980 10559 2000
rect 10525 1966 10559 1980
rect 10593 1966 10627 2000
rect 10525 1946 10661 1966
rect 10491 1931 10661 1946
rect 10491 1910 10559 1931
rect 10525 1897 10559 1910
rect 10593 1897 10627 1931
rect 10525 1876 10661 1897
rect 10491 1862 10661 1876
rect 10491 1840 10559 1862
rect 10525 1828 10559 1840
rect 10593 1828 10627 1862
rect 10525 1806 10661 1828
rect 10491 1793 10661 1806
rect 10491 1770 10559 1793
rect 10525 1759 10559 1770
rect 10593 1759 10627 1793
rect 10525 1736 10661 1759
rect 10491 1724 10661 1736
rect 10491 1701 10559 1724
rect 10525 1690 10559 1701
rect 10593 1690 10627 1724
rect 10525 1667 10661 1690
rect 10491 1655 10661 1667
rect 10491 1632 10559 1655
rect 10525 1621 10559 1632
rect 10593 1621 10627 1655
rect 10525 1598 10661 1621
rect 10491 1586 10661 1598
rect 10491 1563 10559 1586
rect 10525 1552 10559 1563
rect 10593 1552 10627 1586
rect 10525 1529 10661 1552
rect 10491 1517 10661 1529
rect 10491 1494 10559 1517
rect 10525 1483 10559 1494
rect 10593 1483 10627 1517
rect 10525 1460 10661 1483
rect 10491 1448 10661 1460
rect 10491 1425 10559 1448
rect 10525 1414 10559 1425
rect 10593 1414 10627 1448
rect 10525 1391 10661 1414
rect 10491 1379 10661 1391
rect 10491 1356 10559 1379
rect 10525 1345 10559 1356
rect 10593 1345 10627 1379
rect 10525 1322 10661 1345
rect 10491 1310 10661 1322
rect 10491 1287 10559 1310
rect 10525 1253 10559 1287
rect 10491 1218 10559 1253
rect 10525 1184 10559 1218
rect 10491 1149 10559 1184
rect 10525 1115 10559 1149
rect 10491 1080 10559 1115
rect 10525 1046 10559 1080
rect 10491 1011 10559 1046
rect 10525 977 10559 1011
rect 10491 942 10559 977
rect 10525 908 10559 942
rect 10491 873 10559 908
rect 10525 839 10559 873
rect 10491 804 10559 839
rect 10525 770 10559 804
rect 10491 735 10559 770
rect 10525 701 10559 735
rect 10491 666 10559 701
rect 10525 664 10559 666
rect 15339 3233 15407 3234
rect 15441 3266 15475 3267
rect 15441 3233 15509 3266
rect 15339 3231 15509 3233
rect 15339 3199 15475 3231
rect 15373 3198 15475 3199
rect 15373 3165 15407 3198
rect 15339 3164 15407 3165
rect 15441 3197 15475 3198
rect 15441 3164 15509 3197
rect 15339 3162 15509 3164
rect 15339 3130 15475 3162
rect 15373 3129 15475 3130
rect 15373 3096 15407 3129
rect 15339 3095 15407 3096
rect 15441 3128 15475 3129
rect 15441 3095 15509 3128
rect 15339 3093 15509 3095
rect 15339 3061 15475 3093
rect 15373 3060 15475 3061
rect 15373 3027 15407 3060
rect 15339 3026 15407 3027
rect 15441 3059 15475 3060
rect 15441 3026 15509 3059
rect 15339 3024 15509 3026
rect 15339 2992 15475 3024
rect 15373 2991 15475 2992
rect 15373 2958 15407 2991
rect 15339 2957 15407 2958
rect 15441 2990 15475 2991
rect 15441 2957 15509 2990
rect 15339 2955 15509 2957
rect 15339 2923 15475 2955
rect 15373 2922 15475 2923
rect 15373 2889 15407 2922
rect 15339 2888 15407 2889
rect 15441 2921 15475 2922
rect 15441 2888 15509 2921
rect 15339 2886 15509 2888
rect 15339 2854 15475 2886
rect 15373 2853 15475 2854
rect 15373 2820 15407 2853
rect 15339 2819 15407 2820
rect 15441 2852 15475 2853
rect 15441 2819 15509 2852
rect 15339 2817 15509 2819
rect 15339 2785 15475 2817
rect 15373 2784 15475 2785
rect 15373 2751 15407 2784
rect 15339 2750 15407 2751
rect 15441 2783 15475 2784
rect 15441 2750 15509 2783
rect 15339 2748 15509 2750
rect 15339 2716 15475 2748
rect 15373 2715 15475 2716
rect 15373 2682 15407 2715
rect 15339 2681 15407 2682
rect 15441 2714 15475 2715
rect 15441 2681 15509 2714
rect 15339 2679 15509 2681
rect 15339 2647 15475 2679
rect 15373 2646 15475 2647
rect 15373 2613 15407 2646
rect 15339 2612 15407 2613
rect 15441 2645 15475 2646
rect 15441 2612 15509 2645
rect 15339 2610 15509 2612
rect 15339 2578 15475 2610
rect 15373 2577 15475 2578
rect 15373 2544 15407 2577
rect 15339 2543 15407 2544
rect 15441 2576 15475 2577
rect 15441 2543 15509 2576
rect 15339 2541 15509 2543
rect 15339 2509 15475 2541
rect 15373 2508 15475 2509
rect 15373 2475 15407 2508
rect 15339 2474 15407 2475
rect 15441 2507 15475 2508
rect 15441 2474 15509 2507
rect 15339 2472 15509 2474
rect 15339 2440 15475 2472
rect 15373 2439 15475 2440
rect 15373 2406 15407 2439
rect 15339 2405 15407 2406
rect 15441 2438 15475 2439
rect 15441 2405 15509 2438
rect 15339 2403 15509 2405
rect 15339 2371 15475 2403
rect 15373 2370 15475 2371
rect 15373 2337 15407 2370
rect 15339 2336 15407 2337
rect 15441 2369 15475 2370
rect 15441 2336 15509 2369
rect 15339 2334 15509 2336
rect 15339 2302 15475 2334
rect 15373 2301 15475 2302
rect 15373 2268 15407 2301
rect 15339 2267 15407 2268
rect 15441 2300 15475 2301
rect 15441 2267 15509 2300
rect 15339 2265 15509 2267
rect 15339 2233 15475 2265
rect 15373 2232 15475 2233
rect 15373 2199 15407 2232
rect 15339 2198 15407 2199
rect 15441 2231 15475 2232
rect 15441 2198 15509 2231
rect 15339 2196 15509 2198
rect 15339 2164 15475 2196
rect 15373 2163 15475 2164
rect 15373 2130 15407 2163
rect 15339 2129 15407 2130
rect 15441 2162 15475 2163
rect 15441 2129 15509 2162
rect 15339 2127 15509 2129
rect 15339 2095 15475 2127
rect 15373 2094 15475 2095
rect 15373 2061 15407 2094
rect 15339 2060 15407 2061
rect 15441 2093 15475 2094
rect 15441 2060 15509 2093
rect 15339 2058 15509 2060
rect 15339 2026 15475 2058
rect 15373 2025 15475 2026
rect 15373 1992 15407 2025
rect 15339 1991 15407 1992
rect 15441 2024 15475 2025
rect 15441 1991 15509 2024
rect 15339 1989 15509 1991
rect 15339 1957 15475 1989
rect 15373 1956 15475 1957
rect 15373 1923 15407 1956
rect 15339 1922 15407 1923
rect 15441 1955 15475 1956
rect 15441 1922 15509 1955
rect 15339 1920 15509 1922
rect 15339 1888 15475 1920
rect 15373 1887 15475 1888
rect 15373 1854 15407 1887
rect 15339 1853 15407 1854
rect 15441 1886 15475 1887
rect 15441 1853 15509 1886
rect 15339 1851 15509 1853
rect 15339 1818 15475 1851
rect 15373 1784 15407 1818
rect 15441 1817 15475 1818
rect 15441 1784 15509 1817
rect 15339 1782 15509 1784
rect 15339 1749 15475 1782
rect 15339 1748 15407 1749
rect 15373 1715 15407 1748
rect 15441 1748 15475 1749
rect 15441 1715 15509 1748
rect 15373 1714 15509 1715
rect 15339 1713 15509 1714
rect 15339 1680 15475 1713
rect 15339 1678 15407 1680
rect 15373 1646 15407 1678
rect 15441 1679 15475 1680
rect 15441 1646 15509 1679
rect 15373 1644 15509 1646
rect 15339 1610 15475 1644
rect 15339 1608 15407 1610
rect 15373 1576 15407 1608
rect 15441 1576 15509 1610
rect 15373 1575 15509 1576
rect 15373 1574 15475 1575
rect 15339 1541 15475 1574
rect 15339 1540 15509 1541
rect 15339 1538 15407 1540
rect 15373 1506 15407 1538
rect 15441 1506 15509 1540
rect 15373 1504 15475 1506
rect 15339 1472 15475 1504
rect 15339 1470 15509 1472
rect 15339 1468 15407 1470
rect 15373 1436 15407 1468
rect 15441 1436 15509 1470
rect 15373 1434 15475 1436
rect 15339 1402 15475 1434
rect 15339 1400 15509 1402
rect 15339 1398 15407 1400
rect 15373 1366 15407 1398
rect 15441 1366 15509 1400
rect 15373 1364 15475 1366
rect 15339 1332 15475 1364
rect 15339 1330 15509 1332
rect 15339 1328 15407 1330
rect 15373 1296 15407 1328
rect 15441 1296 15509 1330
rect 15373 1294 15475 1296
rect 15339 1262 15475 1294
rect 15339 1260 15509 1262
rect 15339 1258 15407 1260
rect 15373 1226 15407 1258
rect 15441 1226 15509 1260
rect 15373 1224 15475 1226
rect 15339 1192 15475 1224
rect 15339 1190 15509 1192
rect 15339 1188 15407 1190
rect 15373 1156 15407 1188
rect 15441 1156 15509 1190
rect 15373 1154 15475 1156
rect 15339 1122 15475 1154
rect 15339 1120 15509 1122
rect 15339 1118 15407 1120
rect 15373 1086 15407 1118
rect 15441 1086 15509 1120
rect 15373 1084 15475 1086
rect 15339 1052 15475 1084
rect 15339 1050 15509 1052
rect 15339 1048 15407 1050
rect 15373 1016 15407 1048
rect 15441 1016 15509 1050
rect 15373 1014 15475 1016
rect 15339 982 15475 1014
rect 15339 980 15509 982
rect 15339 978 15407 980
rect 15373 946 15407 978
rect 15441 946 15509 980
rect 15373 944 15475 946
rect 15339 912 15475 944
rect 15339 910 15509 912
rect 15339 908 15407 910
rect 15373 876 15407 908
rect 15441 876 15509 910
rect 15373 874 15475 876
rect 15339 842 15475 874
rect 15339 840 15509 842
rect 15339 838 15407 840
rect 15373 806 15407 838
rect 15441 806 15509 840
rect 15373 804 15475 806
rect 15339 772 15475 804
rect 15339 770 15509 772
rect 15339 768 15407 770
rect 15373 736 15407 768
rect 15441 736 15509 770
rect 15373 734 15475 736
rect 15339 702 15475 734
rect 15339 700 15509 702
rect 15339 698 15407 700
rect 10661 664 10696 698
rect 10730 664 10765 698
rect 10799 664 10834 698
rect 10868 664 10903 698
rect 10937 664 10972 698
rect 11006 664 11041 698
rect 11075 664 11110 698
rect 11144 664 11179 698
rect 11213 664 11248 698
rect 11282 664 11317 698
rect 11351 664 11386 698
rect 11420 664 11455 698
rect 11489 664 11524 698
rect 11558 664 11593 698
rect 11627 664 11662 698
rect 11696 664 11731 698
rect 11765 664 11800 698
rect 11834 664 11869 698
rect 11903 664 11938 698
rect 11972 664 12007 698
rect 10525 632 12007 664
rect 10491 630 12007 632
rect 15373 666 15407 698
rect 15441 666 15509 700
rect 15373 632 15475 666
rect 15373 630 15509 632
rect 10491 596 10559 630
rect 10593 596 10628 630
rect 10662 596 10697 630
rect 10731 596 10766 630
rect 10800 596 10835 630
rect 10869 596 10904 630
rect 10938 596 10973 630
rect 11007 596 11042 630
rect 11076 596 11111 630
rect 11145 596 11180 630
rect 11214 596 11249 630
rect 11283 596 11318 630
rect 11352 596 11387 630
rect 11421 596 11456 630
rect 11490 596 11525 630
rect 11559 596 11594 630
rect 11628 596 11663 630
rect 11697 596 11732 630
rect 11766 596 11801 630
rect 11835 596 11870 630
rect 11904 596 11939 630
rect 15441 596 15509 630
rect 10491 562 11939 596
rect 15407 562 15475 596
rect 10491 528 10525 562
rect 10559 528 10594 562
rect 10628 528 10663 562
rect 10697 528 10732 562
rect 10766 528 10801 562
rect 10835 528 10870 562
rect 10904 528 10939 562
rect 10973 528 11008 562
rect 11042 528 11077 562
rect 11111 528 11146 562
rect 11180 528 11215 562
rect 11249 528 11284 562
rect 11318 528 11353 562
rect 11387 528 11422 562
rect 11456 528 11491 562
rect 11525 528 11560 562
rect 11594 528 11629 562
rect 11663 528 11698 562
rect 11732 528 11767 562
rect 11801 528 11836 562
rect 11870 528 11905 562
rect 15407 528 15509 562
<< mvnsubdiff >>
rect 323 17423 425 17457
rect 16167 17423 16202 17457
rect 16236 17423 16271 17457
rect 16305 17423 16340 17457
rect 16374 17423 16409 17457
rect 16443 17423 16478 17457
rect 16512 17423 16547 17457
rect 16581 17423 16616 17457
rect 16650 17423 16685 17457
rect 16719 17423 16754 17457
rect 16788 17423 16823 17457
rect 16857 17423 16892 17457
rect 16926 17423 16961 17457
rect 16995 17423 17030 17457
rect 17064 17423 17099 17457
rect 17133 17423 17168 17457
rect 17202 17423 17237 17457
rect 17271 17423 17306 17457
rect 17340 17423 17375 17457
rect 17409 17423 17444 17457
rect 17478 17423 17513 17457
rect 17547 17423 17582 17457
rect 17616 17423 17651 17457
rect 17685 17423 17720 17457
rect 17754 17423 17789 17457
rect 17823 17423 17858 17457
rect 17892 17423 17927 17457
rect 17961 17423 17996 17457
rect 18030 17423 18065 17457
rect 18099 17423 18134 17457
rect 18168 17423 18203 17457
rect 18237 17423 18272 17457
rect 18306 17423 18341 17457
rect 18375 17423 18409 17457
rect 357 17389 425 17423
rect 16133 17389 18409 17423
rect 323 17355 391 17389
rect 16133 17355 16168 17389
rect 16202 17355 16237 17389
rect 16271 17355 16306 17389
rect 16340 17355 16375 17389
rect 16409 17355 16444 17389
rect 16478 17355 16513 17389
rect 16547 17355 16582 17389
rect 16616 17355 16651 17389
rect 16685 17355 16720 17389
rect 16754 17355 16789 17389
rect 16823 17355 16858 17389
rect 16892 17355 16927 17389
rect 16961 17355 16996 17389
rect 17030 17355 17065 17389
rect 17099 17355 17134 17389
rect 17168 17355 17203 17389
rect 17237 17355 17272 17389
rect 17306 17355 17341 17389
rect 17375 17355 17410 17389
rect 17444 17355 17479 17389
rect 17513 17355 17548 17389
rect 17582 17355 17617 17389
rect 17651 17355 17686 17389
rect 17720 17355 17755 17389
rect 17789 17355 17824 17389
rect 17858 17355 17893 17389
rect 17927 17355 17962 17389
rect 17996 17355 18031 17389
rect 18065 17355 18100 17389
rect 18134 17355 18169 17389
rect 18203 17355 18238 17389
rect 18272 17355 18307 17389
rect 18341 17355 18409 17389
rect 323 17354 459 17355
rect 357 17320 459 17354
rect 323 17286 391 17320
rect 425 17287 459 17320
rect 16065 17321 18307 17355
rect 16065 17287 16100 17321
rect 16134 17287 16169 17321
rect 16203 17287 16238 17321
rect 16272 17287 16307 17321
rect 16341 17287 16376 17321
rect 16410 17287 16445 17321
rect 16479 17287 16514 17321
rect 16548 17287 16583 17321
rect 16617 17287 16652 17321
rect 16686 17287 16721 17321
rect 16755 17287 16790 17321
rect 16824 17287 16859 17321
rect 16893 17287 16928 17321
rect 16962 17287 16997 17321
rect 17031 17287 17066 17321
rect 17100 17287 17135 17321
rect 17169 17287 17204 17321
rect 17238 17287 17273 17321
rect 17307 17287 17342 17321
rect 17376 17287 17411 17321
rect 17445 17287 17480 17321
rect 17514 17287 17549 17321
rect 17583 17287 17618 17321
rect 17652 17287 17687 17321
rect 17721 17287 17756 17321
rect 17790 17287 17825 17321
rect 17859 17287 17894 17321
rect 17928 17287 17963 17321
rect 17997 17287 18032 17321
rect 18066 17287 18101 17321
rect 18135 17287 18170 17321
rect 18204 17287 18239 17321
rect 425 17286 493 17287
rect 323 17285 493 17286
rect 357 17252 493 17285
rect 357 17251 459 17252
rect 323 17217 391 17251
rect 425 17218 459 17251
rect 425 17217 493 17218
rect 323 17216 493 17217
rect 357 17183 493 17216
rect 357 17182 459 17183
rect 323 17148 391 17182
rect 425 17149 459 17182
rect 425 17148 493 17149
rect 323 17147 493 17148
rect 357 17114 493 17147
rect 357 17113 459 17114
rect 323 17079 391 17113
rect 425 17080 459 17113
rect 425 17079 493 17080
rect 323 17078 493 17079
rect 357 17045 493 17078
rect 357 17044 459 17045
rect 323 17010 391 17044
rect 425 17011 459 17044
rect 425 17010 493 17011
rect 323 17009 493 17010
rect 357 16976 493 17009
rect 357 16975 459 16976
rect 323 16941 391 16975
rect 425 16942 459 16975
rect 425 16941 493 16942
rect 323 16940 493 16941
rect 357 16907 493 16940
rect 357 16906 459 16907
rect 323 16872 391 16906
rect 425 16873 459 16906
rect 425 16872 493 16873
rect 323 16871 493 16872
rect 357 16838 493 16871
rect 357 16837 459 16838
rect 323 16803 391 16837
rect 425 16804 459 16837
rect 425 16803 493 16804
rect 323 16802 493 16803
rect 357 16769 493 16802
rect 357 16768 391 16769
rect 323 16733 391 16768
rect 357 16699 391 16733
rect 323 16664 391 16699
rect 357 16630 391 16664
rect 323 16595 391 16630
rect 357 16561 391 16595
rect 323 16526 391 16561
rect 357 16492 391 16526
rect 323 16457 391 16492
rect 357 16423 391 16457
rect 323 16388 391 16423
rect 357 16354 391 16388
rect 323 16319 391 16354
rect 357 16285 391 16319
rect 323 16250 391 16285
rect 357 16216 391 16250
rect 323 16181 391 16216
rect 357 16147 391 16181
rect 323 16112 391 16147
rect 357 16078 391 16112
rect 323 16043 391 16078
rect 357 16009 391 16043
rect 323 15974 391 16009
rect 357 15940 391 15974
rect 323 15905 391 15940
rect 357 15871 391 15905
rect 323 15836 391 15871
rect 357 15802 391 15836
rect 323 15767 391 15802
rect 357 15733 391 15767
rect 323 15698 391 15733
rect 357 15664 391 15698
rect 323 15629 391 15664
rect 357 15595 391 15629
rect 323 15560 391 15595
rect 357 15526 391 15560
rect 323 15491 391 15526
rect 357 15457 391 15491
rect 323 15422 391 15457
rect 357 15388 391 15422
rect 323 15353 391 15388
rect 357 15319 391 15353
rect 323 15284 391 15319
rect 357 15250 391 15284
rect 323 15215 391 15250
rect 357 15181 391 15215
rect 323 15146 391 15181
rect 357 15112 391 15146
rect 323 15077 391 15112
rect 357 15043 391 15077
rect 323 15008 391 15043
rect 357 14974 391 15008
rect 323 14939 391 14974
rect 357 14905 391 14939
rect 323 14870 391 14905
rect 357 14836 391 14870
rect 323 14801 391 14836
rect 357 14767 391 14801
rect 323 14732 391 14767
rect 357 14698 391 14732
rect 323 14663 391 14698
rect 357 14629 391 14663
rect 323 14594 391 14629
rect 357 14560 391 14594
rect 323 14525 391 14560
rect 323 13879 493 13947
rect 357 13845 391 13879
rect 425 13845 459 13879
rect 323 13810 493 13845
rect 323 13809 391 13810
rect 357 13776 391 13809
rect 425 13776 459 13810
rect 357 13775 493 13776
rect 323 13741 493 13775
rect 323 13739 391 13741
rect 357 13707 391 13739
rect 425 13707 459 13741
rect 357 13705 493 13707
rect 323 13672 493 13705
rect 323 13669 391 13672
rect 357 13635 391 13669
rect 323 13599 391 13635
rect 357 13565 391 13599
rect 323 13529 391 13565
rect 357 13495 391 13529
rect 323 13459 391 13495
rect 357 13425 391 13459
rect 323 13389 391 13425
rect 357 13355 391 13389
rect 323 13319 391 13355
rect 357 13285 391 13319
rect 323 13249 391 13285
rect 357 13215 391 13249
rect 323 13179 391 13215
rect 357 13145 391 13179
rect 323 13109 391 13145
rect 357 13075 391 13109
rect 323 13039 391 13075
rect 357 13005 391 13039
rect 323 12969 391 13005
rect 357 12935 391 12969
rect 323 12899 391 12935
rect 357 12865 391 12899
rect 323 12829 391 12865
rect 357 12795 391 12829
rect 323 12759 391 12795
rect 357 12725 391 12759
rect 323 12689 391 12725
rect 357 12655 391 12689
rect 323 12620 391 12655
rect 357 12618 391 12620
rect 18239 15688 18307 15723
rect 18273 15655 18307 15688
rect 18273 15654 18375 15655
rect 18239 15621 18375 15654
rect 18239 15620 18409 15621
rect 18239 15619 18307 15620
rect 18273 15586 18307 15619
rect 18341 15586 18409 15620
rect 18273 15585 18375 15586
rect 18239 15552 18375 15585
rect 18239 15551 18409 15552
rect 18239 15550 18307 15551
rect 18273 15517 18307 15550
rect 18341 15517 18409 15551
rect 18273 15516 18375 15517
rect 18239 15483 18375 15516
rect 18239 15482 18409 15483
rect 18239 15481 18307 15482
rect 18273 15448 18307 15481
rect 18341 15448 18409 15482
rect 18273 15447 18375 15448
rect 18239 15414 18375 15447
rect 18239 15413 18409 15414
rect 18239 15412 18307 15413
rect 18273 15379 18307 15412
rect 18341 15379 18409 15413
rect 18273 15378 18375 15379
rect 18239 15345 18375 15378
rect 18239 15344 18409 15345
rect 18239 15343 18307 15344
rect 18273 15310 18307 15343
rect 18341 15310 18409 15344
rect 18273 15309 18375 15310
rect 18239 15276 18375 15309
rect 18239 15275 18409 15276
rect 18239 15274 18307 15275
rect 18273 15241 18307 15274
rect 18341 15241 18409 15275
rect 18273 15240 18375 15241
rect 18239 15207 18375 15240
rect 18239 15206 18409 15207
rect 18239 15205 18307 15206
rect 18273 15172 18307 15205
rect 18341 15172 18409 15206
rect 18273 15171 18375 15172
rect 18239 15138 18375 15171
rect 18239 15137 18409 15138
rect 18239 15136 18307 15137
rect 18273 15103 18307 15136
rect 18341 15103 18409 15137
rect 18273 15102 18375 15103
rect 18239 15069 18375 15102
rect 18239 15068 18409 15069
rect 18239 15067 18307 15068
rect 18273 15034 18307 15067
rect 18341 15034 18409 15068
rect 18273 15033 18375 15034
rect 18239 15000 18375 15033
rect 18239 14999 18409 15000
rect 18239 14998 18307 14999
rect 18273 14965 18307 14998
rect 18341 14965 18409 14999
rect 18273 14964 18375 14965
rect 18239 14931 18375 14964
rect 18239 14930 18409 14931
rect 18239 14929 18307 14930
rect 18273 14896 18307 14929
rect 18341 14896 18409 14930
rect 18273 14895 18375 14896
rect 18239 14862 18375 14895
rect 18239 14861 18409 14862
rect 18239 14860 18307 14861
rect 18273 14827 18307 14860
rect 18341 14827 18409 14861
rect 18273 14826 18375 14827
rect 18239 14793 18375 14826
rect 18239 14792 18409 14793
rect 18239 14791 18307 14792
rect 18273 14758 18307 14791
rect 18341 14758 18409 14792
rect 18273 14757 18375 14758
rect 18239 14724 18375 14757
rect 18239 14723 18409 14724
rect 18239 14722 18307 14723
rect 18273 14689 18307 14722
rect 18341 14689 18409 14723
rect 18273 14688 18375 14689
rect 18239 14655 18375 14688
rect 18239 14654 18409 14655
rect 18239 14653 18307 14654
rect 18273 14620 18307 14653
rect 18341 14620 18409 14654
rect 18273 14619 18375 14620
rect 18239 14586 18375 14619
rect 18239 14585 18409 14586
rect 18239 14584 18307 14585
rect 18273 14551 18307 14584
rect 18341 14551 18409 14585
rect 18273 14550 18375 14551
rect 18239 14517 18375 14550
rect 18239 14516 18409 14517
rect 18239 14515 18307 14516
rect 18273 14482 18307 14515
rect 18341 14482 18409 14516
rect 18273 14481 18375 14482
rect 18239 14448 18375 14481
rect 18239 14447 18409 14448
rect 18239 14446 18307 14447
rect 18273 14413 18307 14446
rect 18341 14413 18409 14447
rect 18273 14412 18375 14413
rect 18239 14379 18375 14412
rect 18239 14378 18409 14379
rect 18239 14377 18307 14378
rect 18273 14344 18307 14377
rect 18341 14344 18409 14378
rect 18273 14343 18375 14344
rect 18239 14310 18375 14343
rect 18239 14309 18409 14310
rect 18239 14308 18307 14309
rect 18273 14275 18307 14308
rect 18341 14275 18409 14309
rect 18273 14274 18375 14275
rect 18239 14241 18375 14274
rect 18239 14240 18409 14241
rect 18239 14239 18307 14240
rect 18273 14206 18307 14239
rect 18341 14206 18409 14240
rect 18273 14205 18375 14206
rect 18239 14172 18375 14205
rect 18239 14171 18409 14172
rect 18239 14170 18307 14171
rect 18273 14137 18307 14170
rect 18341 14137 18409 14171
rect 18273 14136 18375 14137
rect 18239 14103 18375 14136
rect 18239 14102 18409 14103
rect 18239 14101 18307 14102
rect 18273 14068 18307 14101
rect 18341 14068 18409 14102
rect 18273 14067 18375 14068
rect 18239 14034 18375 14067
rect 18239 14033 18409 14034
rect 18239 14032 18307 14033
rect 18273 13999 18307 14032
rect 18341 13999 18409 14033
rect 18273 13998 18375 13999
rect 18239 13965 18375 13998
rect 18239 13964 18409 13965
rect 18239 13963 18307 13964
rect 18273 13930 18307 13963
rect 18341 13930 18409 13964
rect 18273 13929 18375 13930
rect 18239 13896 18375 13929
rect 18239 13895 18409 13896
rect 18239 13894 18307 13895
rect 18273 13861 18307 13894
rect 18341 13861 18409 13895
rect 18273 13860 18375 13861
rect 18239 13827 18375 13860
rect 18239 13826 18409 13827
rect 18239 13825 18307 13826
rect 18273 13792 18307 13825
rect 18341 13792 18409 13826
rect 18273 13791 18375 13792
rect 18239 13758 18375 13791
rect 18239 13757 18409 13758
rect 18239 13756 18307 13757
rect 18273 13723 18307 13756
rect 18341 13723 18409 13757
rect 18273 13722 18375 13723
rect 18239 13689 18375 13722
rect 18239 13688 18409 13689
rect 18239 13687 18307 13688
rect 18273 13654 18307 13687
rect 18341 13654 18409 13688
rect 18273 13653 18375 13654
rect 18239 13620 18375 13653
rect 18239 13619 18409 13620
rect 18239 13618 18307 13619
rect 18273 13585 18307 13618
rect 18341 13585 18409 13619
rect 18273 13584 18375 13585
rect 18239 13551 18375 13584
rect 18239 13550 18409 13551
rect 18239 13549 18307 13550
rect 18273 13516 18307 13549
rect 18341 13516 18409 13550
rect 18273 13515 18375 13516
rect 18239 13482 18375 13515
rect 18239 13481 18409 13482
rect 18239 13480 18307 13481
rect 18273 13447 18307 13480
rect 18341 13447 18409 13481
rect 18273 13446 18375 13447
rect 18239 13413 18375 13446
rect 18239 13412 18409 13413
rect 18239 13411 18307 13412
rect 18273 13378 18307 13411
rect 18341 13378 18409 13412
rect 18273 13377 18375 13378
rect 18239 13344 18375 13377
rect 18239 13343 18409 13344
rect 18239 13342 18307 13343
rect 18273 13309 18307 13342
rect 18341 13309 18409 13343
rect 18273 13308 18375 13309
rect 18239 13275 18375 13308
rect 18239 13274 18409 13275
rect 18239 13273 18307 13274
rect 18273 13240 18307 13273
rect 18341 13240 18409 13274
rect 18273 13239 18375 13240
rect 18239 13206 18375 13239
rect 18239 13205 18409 13206
rect 18239 13204 18307 13205
rect 18273 13171 18307 13204
rect 18341 13171 18409 13205
rect 18273 13170 18375 13171
rect 18239 13137 18375 13170
rect 18239 13136 18409 13137
rect 18239 13135 18307 13136
rect 18273 13102 18307 13135
rect 18341 13102 18409 13136
rect 18273 13101 18375 13102
rect 18239 13068 18375 13101
rect 18239 13067 18409 13068
rect 18239 13066 18307 13067
rect 18273 13033 18307 13066
rect 18341 13033 18409 13067
rect 18273 13032 18375 13033
rect 18239 12999 18375 13032
rect 18239 12998 18409 12999
rect 18239 12997 18307 12998
rect 18273 12964 18307 12997
rect 18341 12964 18409 12998
rect 18273 12963 18375 12964
rect 18239 12930 18375 12963
rect 18239 12929 18409 12930
rect 18239 12928 18307 12929
rect 18273 12895 18307 12928
rect 18341 12895 18409 12929
rect 18273 12894 18375 12895
rect 18239 12861 18375 12894
rect 18239 12860 18409 12861
rect 18239 12859 18307 12860
rect 18273 12826 18307 12859
rect 18341 12826 18409 12860
rect 18273 12825 18375 12826
rect 18239 12792 18375 12825
rect 18239 12791 18409 12792
rect 18239 12790 18307 12791
rect 18273 12757 18307 12790
rect 18341 12757 18409 12791
rect 18273 12756 18375 12757
rect 18239 12723 18375 12756
rect 18239 12722 18409 12723
rect 18239 12721 18307 12722
rect 18273 12688 18307 12721
rect 18341 12688 18409 12722
rect 18273 12687 18375 12688
rect 18239 12654 18375 12687
rect 18239 12653 18409 12654
rect 18239 12652 18307 12653
rect 493 12618 528 12652
rect 562 12618 597 12652
rect 631 12618 666 12652
rect 700 12618 735 12652
rect 769 12618 804 12652
rect 838 12618 873 12652
rect 907 12618 942 12652
rect 976 12618 1011 12652
rect 1045 12618 1080 12652
rect 1114 12618 1149 12652
rect 1183 12618 1218 12652
rect 1252 12618 1287 12652
rect 1321 12618 1356 12652
rect 1390 12618 1425 12652
rect 1459 12618 1494 12652
rect 1528 12618 1563 12652
rect 1597 12618 1632 12652
rect 1666 12618 1701 12652
rect 1735 12618 1770 12652
rect 1804 12618 1839 12652
rect 1873 12618 1908 12652
rect 1942 12618 1977 12652
rect 2011 12618 2046 12652
rect 2080 12618 2115 12652
rect 2149 12618 2184 12652
rect 2218 12618 2253 12652
rect 2287 12618 2322 12652
rect 2356 12618 2391 12652
rect 2425 12618 2460 12652
rect 2494 12618 2529 12652
rect 2563 12618 2598 12652
rect 2632 12618 2667 12652
rect 357 12586 2667 12618
rect 323 12584 2667 12586
rect 18273 12619 18307 12652
rect 18341 12619 18409 12653
rect 18273 12585 18375 12619
rect 18273 12584 18409 12585
rect 323 12550 391 12584
rect 425 12550 460 12584
rect 494 12550 529 12584
rect 563 12550 598 12584
rect 632 12550 667 12584
rect 701 12550 736 12584
rect 770 12550 805 12584
rect 839 12550 874 12584
rect 908 12550 943 12584
rect 977 12550 1012 12584
rect 1046 12550 1081 12584
rect 1115 12550 1150 12584
rect 1184 12550 1219 12584
rect 1253 12550 1288 12584
rect 1322 12550 1357 12584
rect 1391 12550 1426 12584
rect 1460 12550 1495 12584
rect 1529 12550 1564 12584
rect 1598 12550 1633 12584
rect 1667 12550 1702 12584
rect 1736 12550 1771 12584
rect 1805 12550 1840 12584
rect 1874 12550 1909 12584
rect 1943 12550 1978 12584
rect 2012 12550 2047 12584
rect 2081 12550 2116 12584
rect 2150 12550 2185 12584
rect 2219 12550 2254 12584
rect 2288 12550 2323 12584
rect 2357 12550 2392 12584
rect 2426 12550 2461 12584
rect 2495 12550 2530 12584
rect 2564 12550 2599 12584
rect 18341 12550 18409 12584
rect 323 12516 2599 12550
rect 18307 12516 18375 12550
rect 323 12482 357 12516
rect 391 12482 426 12516
rect 460 12482 495 12516
rect 529 12482 564 12516
rect 598 12482 633 12516
rect 667 12482 702 12516
rect 736 12482 771 12516
rect 805 12482 840 12516
rect 874 12482 909 12516
rect 943 12482 978 12516
rect 1012 12482 1047 12516
rect 1081 12482 1116 12516
rect 1150 12482 1185 12516
rect 1219 12482 1254 12516
rect 1288 12482 1323 12516
rect 1357 12482 1392 12516
rect 1426 12482 1461 12516
rect 1495 12482 1530 12516
rect 1564 12482 1599 12516
rect 1633 12482 1668 12516
rect 1702 12482 1737 12516
rect 1771 12482 1806 12516
rect 1840 12482 1875 12516
rect 1909 12482 1944 12516
rect 1978 12482 2013 12516
rect 2047 12482 2082 12516
rect 2116 12482 2151 12516
rect 2185 12482 2220 12516
rect 2254 12482 2289 12516
rect 2323 12482 2358 12516
rect 2392 12482 2427 12516
rect 2461 12482 2496 12516
rect 2530 12482 2565 12516
rect 18307 12482 18409 12516
rect 10135 3692 10237 3726
rect 14555 3692 14590 3726
rect 14624 3692 14659 3726
rect 14693 3692 14728 3726
rect 14762 3692 14797 3726
rect 14831 3692 14866 3726
rect 14900 3692 14935 3726
rect 14969 3692 15004 3726
rect 15038 3692 15073 3726
rect 15107 3692 15142 3726
rect 15176 3692 15211 3726
rect 15245 3692 15280 3726
rect 15314 3692 15349 3726
rect 15383 3692 15418 3726
rect 15452 3692 15487 3726
rect 15521 3692 15556 3726
rect 15590 3692 15625 3726
rect 15659 3692 15694 3726
rect 15728 3692 15763 3726
rect 15797 3692 15831 3726
rect 10169 3658 10237 3692
rect 14521 3658 15831 3692
rect 10135 3624 10203 3658
rect 14521 3624 14556 3658
rect 14590 3624 14625 3658
rect 14659 3624 14694 3658
rect 14728 3624 14763 3658
rect 14797 3624 14832 3658
rect 14866 3624 14901 3658
rect 14935 3624 14970 3658
rect 15004 3624 15039 3658
rect 15073 3624 15108 3658
rect 15142 3624 15177 3658
rect 15211 3624 15246 3658
rect 15280 3624 15315 3658
rect 15349 3624 15384 3658
rect 15418 3624 15453 3658
rect 15487 3624 15522 3658
rect 15556 3624 15591 3658
rect 15625 3624 15660 3658
rect 15694 3624 15729 3658
rect 15763 3624 15831 3658
rect 10135 3617 10271 3624
rect 10169 3587 10271 3617
rect 10169 3583 10203 3587
rect 10135 3553 10203 3583
rect 10237 3556 10271 3587
rect 14453 3590 15797 3624
rect 14453 3556 14488 3590
rect 14522 3556 14557 3590
rect 14591 3556 14626 3590
rect 14660 3556 14695 3590
rect 14729 3556 14764 3590
rect 14798 3556 14833 3590
rect 14867 3556 14902 3590
rect 14936 3556 14971 3590
rect 15005 3556 15040 3590
rect 15074 3556 15109 3590
rect 15143 3556 15178 3590
rect 15212 3556 15247 3590
rect 15281 3556 15316 3590
rect 15350 3556 15385 3590
rect 15419 3556 15454 3590
rect 15488 3556 15523 3590
rect 15557 3556 15592 3590
rect 15626 3556 15661 3590
rect 15695 3589 15831 3590
rect 15695 3556 15729 3589
rect 10237 3553 10305 3556
rect 10135 3543 10305 3553
rect 10169 3519 10305 3543
rect 10169 3516 10271 3519
rect 10169 3509 10203 3516
rect 10135 3482 10203 3509
rect 10237 3485 10271 3516
rect 10237 3482 10305 3485
rect 10135 3469 10305 3482
rect 10169 3448 10305 3469
rect 10169 3445 10271 3448
rect 10169 3435 10203 3445
rect 10135 3411 10203 3435
rect 10237 3414 10271 3445
rect 10237 3411 10305 3414
rect 10135 3395 10305 3411
rect 15661 3555 15729 3556
rect 15763 3556 15831 3589
rect 15763 3555 15797 3556
rect 15661 3522 15797 3555
rect 15661 3521 15831 3522
rect 15695 3520 15831 3521
rect 15695 3487 15729 3520
rect 15661 3486 15729 3487
rect 15763 3488 15831 3520
rect 15763 3486 15797 3488
rect 15661 3454 15797 3486
rect 15661 3452 15831 3454
rect 15695 3451 15831 3452
rect 15695 3418 15729 3451
rect 15661 3417 15729 3418
rect 15763 3420 15831 3451
rect 15763 3417 15797 3420
rect 10169 3377 10305 3395
rect 10169 3374 10271 3377
rect 10169 3361 10203 3374
rect 10135 3340 10203 3361
rect 10237 3343 10271 3374
rect 10237 3340 10305 3343
rect 10135 3321 10305 3340
rect 10169 3306 10305 3321
rect 10169 3303 10271 3306
rect 10169 3287 10203 3303
rect 10135 3269 10203 3287
rect 10237 3272 10271 3303
rect 10237 3269 10305 3272
rect 10135 3247 10305 3269
rect 10169 3235 10305 3247
rect 10169 3232 10271 3235
rect 10169 3213 10203 3232
rect 10135 3198 10203 3213
rect 10237 3201 10271 3232
rect 10237 3198 10305 3201
rect 10135 3173 10305 3198
rect 10169 3164 10305 3173
rect 10169 3161 10271 3164
rect 10169 3139 10203 3161
rect 10135 3127 10203 3139
rect 10237 3130 10271 3161
rect 10237 3127 10305 3130
rect 10135 3099 10305 3127
rect 10169 3093 10305 3099
rect 10169 3091 10271 3093
rect 10169 3065 10203 3091
rect 10135 3057 10203 3065
rect 10237 3059 10271 3091
rect 10237 3057 10305 3059
rect 10135 3025 10305 3057
rect 10169 3022 10305 3025
rect 10169 3021 10271 3022
rect 10169 2991 10203 3021
rect 10135 2987 10203 2991
rect 10237 2988 10271 3021
rect 10237 2987 10305 2988
rect 10135 2951 10305 2987
rect 10169 2917 10203 2951
rect 10237 2917 10271 2951
rect 10135 236 10305 2917
rect 15661 3386 15797 3417
rect 15661 3383 15831 3386
rect 15695 3382 15831 3383
rect 15695 3349 15729 3382
rect 15661 3348 15729 3349
rect 15763 3352 15831 3382
rect 15763 3348 15797 3352
rect 15661 3318 15797 3348
rect 15661 3314 15831 3318
rect 15695 3313 15831 3314
rect 15695 3280 15729 3313
rect 15661 3279 15729 3280
rect 15763 3284 15831 3313
rect 15763 3279 15797 3284
rect 15661 3250 15797 3279
rect 15661 3245 15831 3250
rect 15695 3244 15831 3245
rect 15695 3211 15729 3244
rect 15661 3210 15729 3211
rect 15763 3216 15831 3244
rect 15763 3210 15797 3216
rect 15661 3182 15797 3210
rect 15661 3176 15831 3182
rect 15695 3175 15831 3176
rect 15695 3142 15729 3175
rect 15661 3141 15729 3142
rect 15763 3148 15831 3175
rect 15763 3141 15797 3148
rect 15661 3114 15797 3141
rect 15661 3107 15831 3114
rect 15695 3106 15831 3107
rect 15695 3073 15729 3106
rect 15661 3072 15729 3073
rect 15763 3080 15831 3106
rect 15763 3072 15797 3080
rect 15661 3046 15797 3072
rect 15661 3038 15831 3046
rect 15695 3037 15831 3038
rect 15695 3004 15729 3037
rect 15661 3003 15729 3004
rect 15763 3012 15831 3037
rect 15763 3003 15797 3012
rect 15661 2978 15797 3003
rect 15661 2969 15831 2978
rect 15695 2968 15831 2969
rect 15695 2935 15729 2968
rect 15661 2934 15729 2935
rect 15763 2944 15831 2968
rect 15763 2934 15797 2944
rect 15661 2910 15797 2934
rect 15661 2900 15831 2910
rect 15695 2899 15831 2900
rect 15695 2866 15729 2899
rect 15661 2865 15729 2866
rect 15763 2876 15831 2899
rect 15763 2865 15797 2876
rect 15661 2842 15797 2865
rect 15661 2831 15831 2842
rect 15695 2830 15831 2831
rect 15695 2797 15729 2830
rect 15661 2796 15729 2797
rect 15763 2808 15831 2830
rect 15763 2796 15797 2808
rect 15661 2774 15797 2796
rect 15661 2762 15831 2774
rect 15695 2761 15831 2762
rect 15695 2728 15729 2761
rect 15661 2727 15729 2728
rect 15763 2740 15831 2761
rect 15763 2727 15797 2740
rect 15661 2706 15797 2727
rect 15661 2693 15831 2706
rect 15695 2692 15831 2693
rect 15695 2659 15729 2692
rect 15661 2658 15729 2659
rect 15763 2672 15831 2692
rect 15763 2658 15797 2672
rect 15661 2638 15797 2658
rect 15661 2624 15831 2638
rect 15695 2623 15831 2624
rect 15695 2590 15729 2623
rect 15661 2589 15729 2590
rect 15763 2604 15831 2623
rect 15763 2589 15797 2604
rect 15661 2570 15797 2589
rect 15661 2555 15831 2570
rect 15695 2554 15831 2555
rect 15695 2521 15729 2554
rect 15661 2520 15729 2521
rect 15763 2536 15831 2554
rect 15763 2520 15797 2536
rect 15661 2502 15797 2520
rect 15661 2486 15831 2502
rect 15695 2485 15831 2486
rect 15695 2452 15729 2485
rect 15661 2451 15729 2452
rect 15763 2468 15831 2485
rect 15763 2451 15797 2468
rect 15661 2434 15797 2451
rect 15661 2417 15831 2434
rect 15695 2416 15831 2417
rect 15695 2383 15729 2416
rect 15661 2382 15729 2383
rect 15763 2400 15831 2416
rect 15763 2382 15797 2400
rect 15661 2366 15797 2382
rect 15661 2348 15831 2366
rect 15695 2347 15831 2348
rect 15695 2314 15729 2347
rect 15661 2313 15729 2314
rect 15763 2331 15831 2347
rect 15763 2313 15797 2331
rect 15661 2297 15797 2313
rect 15661 2279 15831 2297
rect 15695 2278 15831 2279
rect 15695 2245 15729 2278
rect 15661 2244 15729 2245
rect 15763 2262 15831 2278
rect 15763 2244 15797 2262
rect 15661 2228 15797 2244
rect 15661 2210 15831 2228
rect 15695 2209 15831 2210
rect 15695 2176 15729 2209
rect 15661 2175 15729 2176
rect 15763 2193 15831 2209
rect 15763 2175 15797 2193
rect 15661 2159 15797 2175
rect 15661 2141 15831 2159
rect 15695 2140 15831 2141
rect 15695 2107 15729 2140
rect 15661 2106 15729 2107
rect 15763 2124 15831 2140
rect 15763 2106 15797 2124
rect 15661 2090 15797 2106
rect 15661 2072 15831 2090
rect 15695 2071 15831 2072
rect 15695 2038 15729 2071
rect 15661 2037 15729 2038
rect 15763 2055 15831 2071
rect 15763 2037 15797 2055
rect 15661 2021 15797 2037
rect 15661 2003 15831 2021
rect 15695 2002 15831 2003
rect 15695 1969 15729 2002
rect 15661 1968 15729 1969
rect 15763 1986 15831 2002
rect 15763 1968 15797 1986
rect 15661 1952 15797 1968
rect 15661 1934 15831 1952
rect 15695 1933 15831 1934
rect 15695 1900 15729 1933
rect 15661 1899 15729 1900
rect 15763 1917 15831 1933
rect 15763 1899 15797 1917
rect 15661 1883 15797 1899
rect 15661 1865 15831 1883
rect 15695 1864 15831 1865
rect 15695 1831 15729 1864
rect 15661 1830 15729 1831
rect 15763 1848 15831 1864
rect 15763 1830 15797 1848
rect 15661 1814 15797 1830
rect 15661 1796 15831 1814
rect 15695 1795 15831 1796
rect 15695 1762 15729 1795
rect 15661 1761 15729 1762
rect 15763 1779 15831 1795
rect 15763 1761 15797 1779
rect 15661 1745 15797 1761
rect 15661 1727 15831 1745
rect 15695 1726 15831 1727
rect 15695 1693 15729 1726
rect 15661 1692 15729 1693
rect 15763 1710 15831 1726
rect 15763 1692 15797 1710
rect 15661 1676 15797 1692
rect 15661 1658 15831 1676
rect 15695 1657 15831 1658
rect 15695 1624 15729 1657
rect 15661 1623 15729 1624
rect 15763 1641 15831 1657
rect 15763 1623 15797 1641
rect 15661 1607 15797 1623
rect 15661 1589 15831 1607
rect 15695 1588 15831 1589
rect 15695 1555 15729 1588
rect 15661 1554 15729 1555
rect 15763 1572 15831 1588
rect 15763 1554 15797 1572
rect 15661 1538 15797 1554
rect 15661 1520 15831 1538
rect 15695 1519 15831 1520
rect 15695 1486 15729 1519
rect 15661 1485 15729 1486
rect 15763 1503 15831 1519
rect 15763 1485 15797 1503
rect 15661 1469 15797 1485
rect 15661 1450 15831 1469
rect 15695 1416 15729 1450
rect 15763 1434 15831 1450
rect 15763 1416 15797 1434
rect 15661 1400 15797 1416
rect 15661 1380 15831 1400
rect 15695 1346 15729 1380
rect 15763 1365 15831 1380
rect 15763 1346 15797 1365
rect 15661 1331 15797 1346
rect 15661 1310 15831 1331
rect 15695 1276 15729 1310
rect 15763 1296 15831 1310
rect 15763 1276 15797 1296
rect 15661 1262 15797 1276
rect 15661 1240 15831 1262
rect 15695 1206 15729 1240
rect 15763 1227 15831 1240
rect 15763 1206 15797 1227
rect 15661 1193 15797 1206
rect 15661 1170 15831 1193
rect 15695 1136 15729 1170
rect 15763 1158 15831 1170
rect 15763 1136 15797 1158
rect 15661 1124 15797 1136
rect 15661 1100 15831 1124
rect 15695 1066 15729 1100
rect 15763 1089 15831 1100
rect 15763 1066 15797 1089
rect 15661 1055 15797 1066
rect 15661 1030 15831 1055
rect 15695 996 15729 1030
rect 15763 1020 15831 1030
rect 15763 996 15797 1020
rect 15661 986 15797 996
rect 15661 960 15831 986
rect 15695 926 15729 960
rect 15763 951 15831 960
rect 15763 926 15797 951
rect 15661 917 15797 926
rect 15661 890 15831 917
rect 15695 856 15729 890
rect 15763 882 15831 890
rect 15763 856 15797 882
rect 15661 848 15797 856
rect 15661 820 15831 848
rect 15695 786 15729 820
rect 15763 813 15831 820
rect 15763 786 15797 813
rect 15661 779 15797 786
rect 15661 750 15831 779
rect 15695 716 15729 750
rect 15763 744 15831 750
rect 15763 716 15797 744
rect 15661 710 15797 716
rect 15661 680 15831 710
rect 15695 646 15729 680
rect 15763 675 15831 680
rect 15763 646 15797 675
rect 15661 641 15797 646
rect 15661 610 15831 641
rect 15695 576 15729 610
rect 15763 606 15831 610
rect 15763 576 15797 606
rect 15661 572 15797 576
rect 15661 540 15831 572
rect 15695 506 15729 540
rect 15763 537 15831 540
rect 15763 506 15797 537
rect 15661 503 15797 506
rect 15661 470 15831 503
rect 15695 436 15729 470
rect 15763 468 15831 470
rect 15763 436 15797 468
rect 15661 434 15797 436
rect 15661 400 15831 434
rect 15695 366 15729 400
rect 15763 399 15831 400
rect 15763 366 15797 399
rect 15661 365 15797 366
rect 15661 330 15831 365
rect 15695 296 15729 330
rect 15763 296 15797 330
rect 15661 236 15831 296
rect 10135 66 15831 236
<< psubdiffcont >>
rect 102 17793 15640 17827
rect 15675 17793 15709 17827
rect 15744 17793 15778 17827
rect 15813 17793 15847 17827
rect 15882 17793 15916 17827
rect 15951 17793 15985 17827
rect 16020 17793 16054 17827
rect 16089 17793 16123 17827
rect 16158 17793 16192 17827
rect 16227 17793 16261 17827
rect 16296 17793 16330 17827
rect 16365 17793 16399 17827
rect 16434 17793 16468 17827
rect 16503 17793 16537 17827
rect 16572 17793 16606 17827
rect 16641 17793 16675 17827
rect 16710 17793 16744 17827
rect 16779 17793 16813 17827
rect 16848 17793 16882 17827
rect 16917 17793 16951 17827
rect 16986 17793 17020 17827
rect 17055 17793 17089 17827
rect 17124 17793 17158 17827
rect 17193 17793 17227 17827
rect 17262 17793 17296 17827
rect 17331 17793 17365 17827
rect 17400 17793 17434 17827
rect 17469 17793 17503 17827
rect 17538 17793 17572 17827
rect 17607 17793 17641 17827
rect 17676 17793 17710 17827
rect 17745 17793 17779 17827
rect 17814 17793 17848 17827
rect 17883 17793 17917 17827
rect 17952 17793 17986 17827
rect 18021 17793 18055 17827
rect 18090 17793 18124 17827
rect 18159 17793 18193 17827
rect 18228 17793 18262 17827
rect 18297 17793 18331 17827
rect 18366 17793 18400 17827
rect 18435 17793 18469 17827
rect 18504 17793 18538 17827
rect 18573 17793 18607 17827
rect 18642 17793 18676 17827
rect 18711 17793 18745 17827
rect 0 17759 34 17793
rect 102 17759 15606 17793
rect 68 17725 15606 17759
rect 15641 17725 15675 17759
rect 15710 17725 15744 17759
rect 15779 17725 15813 17759
rect 15848 17725 15882 17759
rect 15917 17725 15951 17759
rect 15986 17725 16020 17759
rect 16055 17725 16089 17759
rect 16124 17725 16158 17759
rect 16193 17725 16227 17759
rect 16262 17725 16296 17759
rect 16331 17725 16365 17759
rect 16400 17725 16434 17759
rect 16469 17725 16503 17759
rect 16538 17725 16572 17759
rect 16607 17725 16641 17759
rect 16676 17725 16710 17759
rect 16745 17725 16779 17759
rect 16814 17725 16848 17759
rect 16883 17725 16917 17759
rect 16952 17725 16986 17759
rect 17021 17725 17055 17759
rect 17090 17725 17124 17759
rect 17159 17725 17193 17759
rect 17228 17725 17262 17759
rect 17297 17725 17331 17759
rect 17366 17725 17400 17759
rect 17435 17725 17469 17759
rect 17504 17725 17538 17759
rect 17573 17725 17607 17759
rect 17642 17725 17676 17759
rect 17711 17725 17745 17759
rect 17780 17725 17814 17759
rect 17849 17725 17883 17759
rect 17918 17725 17952 17759
rect 17987 17725 18021 17759
rect 18056 17725 18090 17759
rect 18125 17725 18159 17759
rect 18194 17725 18228 17759
rect 18263 17725 18297 17759
rect 18332 17725 18366 17759
rect 18401 17725 18435 17759
rect 18470 17725 18504 17759
rect 18539 17725 18573 17759
rect 18608 17725 18642 17759
rect 18677 17725 18711 17759
rect 0 17689 34 17723
rect 68 17656 102 17690
rect 136 17657 15538 17725
rect 18677 17691 18779 17725
rect 15573 17657 15607 17691
rect 15642 17657 15676 17691
rect 15711 17657 15745 17691
rect 15780 17657 15814 17691
rect 15849 17657 15883 17691
rect 15918 17657 15952 17691
rect 15987 17657 16021 17691
rect 16056 17657 16090 17691
rect 16125 17657 16159 17691
rect 16194 17657 16228 17691
rect 16263 17657 16297 17691
rect 16332 17657 16366 17691
rect 16401 17657 16435 17691
rect 16470 17657 16504 17691
rect 16539 17657 16573 17691
rect 16608 17657 16642 17691
rect 16677 17657 16711 17691
rect 16746 17657 16780 17691
rect 16815 17657 16849 17691
rect 16884 17657 16918 17691
rect 16953 17657 16987 17691
rect 17022 17657 17056 17691
rect 17091 17657 17125 17691
rect 17160 17657 17194 17691
rect 17229 17657 17263 17691
rect 17298 17657 17332 17691
rect 17367 17657 17401 17691
rect 17436 17657 17470 17691
rect 17505 17657 17539 17691
rect 17574 17657 17608 17691
rect 17643 17657 17677 17691
rect 17712 17657 17746 17691
rect 17781 17657 17815 17691
rect 17850 17657 17884 17691
rect 17919 17657 17953 17691
rect 17988 17657 18022 17691
rect 18057 17657 18091 17691
rect 18126 17657 18160 17691
rect 18195 17657 18229 17691
rect 18264 17657 18298 17691
rect 18333 17657 18367 17691
rect 18402 17657 18436 17691
rect 18471 17657 18505 17691
rect 18540 17657 18574 17691
rect 0 17619 34 17653
rect 68 17587 102 17621
rect 136 17588 170 17622
rect 0 17549 34 17583
rect 68 17518 102 17552
rect 136 17519 170 17553
rect 0 17479 34 17513
rect 68 17449 102 17483
rect 136 17450 170 17484
rect 0 17409 34 17443
rect 68 17380 102 17414
rect 136 17381 170 17415
rect 0 17339 34 17373
rect 68 17311 102 17345
rect 136 17312 170 17346
rect 0 17269 34 17303
rect 68 17242 102 17276
rect 136 17243 170 17277
rect 0 17199 34 17233
rect 68 17173 102 17207
rect 136 17174 170 17208
rect 0 17130 34 17164
rect 68 17104 102 17138
rect 136 17105 170 17139
rect 0 17061 34 17095
rect 68 17035 102 17069
rect 136 17036 170 17070
rect 0 16992 34 17026
rect 68 16966 102 17000
rect 136 16967 170 17001
rect 0 16923 34 16957
rect 68 16897 102 16931
rect 136 16898 170 16932
rect 0 16854 34 16888
rect 68 16828 102 16862
rect 136 16829 170 16863
rect 0 16785 34 16819
rect 68 16759 102 16793
rect 136 16760 170 16794
rect 0 16716 34 16750
rect 68 16690 102 16724
rect 136 16691 170 16725
rect 0 16647 34 16681
rect 68 16621 102 16655
rect 136 16622 170 16656
rect 0 16578 34 16612
rect 68 16552 102 16586
rect 136 16553 170 16587
rect 0 16509 34 16543
rect 68 16483 102 16517
rect 136 16484 170 16518
rect 0 16440 34 16474
rect 68 16414 102 16448
rect 136 16415 170 16449
rect 0 16371 34 16405
rect 68 16345 102 16379
rect 136 16346 170 16380
rect 0 16302 34 16336
rect 68 16276 102 16310
rect 136 16277 170 16311
rect 0 16233 34 16267
rect 68 16207 102 16241
rect 136 16208 170 16242
rect 0 16164 34 16198
rect 68 16138 102 16172
rect 136 16139 170 16173
rect 0 16095 34 16129
rect 68 16069 102 16103
rect 136 16070 170 16104
rect 0 16026 34 16060
rect 68 16000 102 16034
rect 136 16001 170 16035
rect 0 15957 34 15991
rect 68 15931 102 15965
rect 136 15932 170 15966
rect 0 15888 34 15922
rect 68 15862 102 15896
rect 136 15863 170 15897
rect 0 15819 34 15853
rect 68 15793 102 15827
rect 136 15794 170 15828
rect 0 15750 34 15784
rect 68 15724 102 15758
rect 136 15725 170 15759
rect 0 15681 34 15715
rect 0 15612 34 15646
rect 0 15543 34 15577
rect 0 15474 34 15508
rect 0 15405 34 15439
rect 0 15336 34 15370
rect 0 15267 34 15301
rect 0 15198 34 15232
rect 0 15129 34 15163
rect 0 15060 34 15094
rect 0 14991 34 15025
rect 0 14922 34 14956
rect 0 14853 34 14887
rect 0 14784 34 14818
rect 0 14715 34 14749
rect 0 14646 34 14680
rect 0 14577 34 14611
rect 0 14508 34 14542
rect 0 14439 34 14473
rect 0 14370 34 14404
rect 0 14301 34 14335
rect 0 14232 34 14266
rect 0 14163 34 14197
rect 0 14094 34 14128
rect 0 14025 34 14059
rect 0 13956 34 13990
rect 68 13956 170 15690
rect 0 13854 34 13888
rect 68 13854 102 13888
rect 136 13854 170 13888
rect 0 13785 34 13819
rect 68 13785 102 13819
rect 136 13785 170 13819
rect 0 13716 34 13750
rect 68 13716 102 13750
rect 136 13716 170 13750
rect 0 13647 34 13681
rect 68 13647 102 13681
rect 136 13647 170 13681
rect 0 13578 34 13612
rect 68 13578 102 13612
rect 136 13578 170 13612
rect 0 12285 170 13543
rect 748 17100 13498 17134
rect 13533 17100 13567 17134
rect 13602 17100 13636 17134
rect 13671 17100 13705 17134
rect 13740 17100 13774 17134
rect 13809 17100 13843 17134
rect 13878 17100 13912 17134
rect 13947 17100 13981 17134
rect 14016 17100 14050 17134
rect 14085 17100 14119 17134
rect 14154 17100 14188 17134
rect 14223 17100 14257 17134
rect 14292 17100 14326 17134
rect 14361 17100 14395 17134
rect 14430 17100 14464 17134
rect 14499 17100 14533 17134
rect 14568 17100 14602 17134
rect 14637 17100 14671 17134
rect 14706 17100 14740 17134
rect 14775 17100 14809 17134
rect 14844 17100 14878 17134
rect 14913 17100 14947 17134
rect 14982 17100 15016 17134
rect 15051 17100 15085 17134
rect 15120 17100 15154 17134
rect 15189 17100 15223 17134
rect 15258 17100 15292 17134
rect 15327 17100 15361 17134
rect 15396 17100 15430 17134
rect 15465 17100 15499 17134
rect 15534 17100 15568 17134
rect 15603 17100 15637 17134
rect 15672 17100 15706 17134
rect 15741 17100 15775 17134
rect 15810 17100 15844 17134
rect 15879 17100 15913 17134
rect 15948 17100 15982 17134
rect 16017 17100 16051 17134
rect 16086 17100 16120 17134
rect 16155 17100 16189 17134
rect 16224 17100 16258 17134
rect 16293 17100 16327 17134
rect 16362 17100 16396 17134
rect 16431 17100 16465 17134
rect 16500 17100 16534 17134
rect 16569 17100 16603 17134
rect 16638 17100 16672 17134
rect 16707 17100 16741 17134
rect 16776 17100 16810 17134
rect 16845 17100 16879 17134
rect 16914 17100 16948 17134
rect 16983 17100 17017 17134
rect 17052 17100 17086 17134
rect 17121 17100 17155 17134
rect 17190 17100 17224 17134
rect 17259 17100 17293 17134
rect 17328 17100 17362 17134
rect 17397 17100 17431 17134
rect 17466 17100 17500 17134
rect 17535 17100 17569 17134
rect 17604 17100 17638 17134
rect 17673 17100 17707 17134
rect 17742 17100 17776 17134
rect 17811 17100 17845 17134
rect 17880 17100 17914 17134
rect 17949 17100 17983 17134
rect 18018 17100 18052 17134
rect 646 17066 680 17100
rect 748 17066 13464 17100
rect 714 17032 13464 17066
rect 13499 17032 13533 17066
rect 13568 17032 13602 17066
rect 13637 17032 13671 17066
rect 13706 17032 13740 17066
rect 13775 17032 13809 17066
rect 13844 17032 13878 17066
rect 13913 17032 13947 17066
rect 13982 17032 14016 17066
rect 14051 17032 14085 17066
rect 14120 17032 14154 17066
rect 14189 17032 14223 17066
rect 14258 17032 14292 17066
rect 14327 17032 14361 17066
rect 14396 17032 14430 17066
rect 14465 17032 14499 17066
rect 14534 17032 14568 17066
rect 14603 17032 14637 17066
rect 14672 17032 14706 17066
rect 14741 17032 14775 17066
rect 14810 17032 14844 17066
rect 14879 17032 14913 17066
rect 14948 17032 14982 17066
rect 15017 17032 15051 17066
rect 15086 17032 15120 17066
rect 15155 17032 15189 17066
rect 15224 17032 15258 17066
rect 15293 17032 15327 17066
rect 15362 17032 15396 17066
rect 15431 17032 15465 17066
rect 15500 17032 15534 17066
rect 15569 17032 15603 17066
rect 15638 17032 15672 17066
rect 15707 17032 15741 17066
rect 15776 17032 15810 17066
rect 15845 17032 15879 17066
rect 15914 17032 15948 17066
rect 15983 17032 16017 17066
rect 16052 17032 16086 17066
rect 16121 17032 16155 17066
rect 16190 17032 16224 17066
rect 16259 17032 16293 17066
rect 16328 17032 16362 17066
rect 16397 17032 16431 17066
rect 16466 17032 16500 17066
rect 16535 17032 16569 17066
rect 16604 17032 16638 17066
rect 16673 17032 16707 17066
rect 16742 17032 16776 17066
rect 16811 17032 16845 17066
rect 16880 17032 16914 17066
rect 16949 17032 16983 17066
rect 17018 17032 17052 17066
rect 17087 17032 17121 17066
rect 17156 17032 17190 17066
rect 17225 17032 17259 17066
rect 17294 17032 17328 17066
rect 17363 17032 17397 17066
rect 17432 17032 17466 17066
rect 17501 17032 17535 17066
rect 17570 17032 17604 17066
rect 17639 17032 17673 17066
rect 17708 17032 17742 17066
rect 17777 17032 17811 17066
rect 17846 17032 17880 17066
rect 17915 17032 17949 17066
rect 17984 17032 18018 17066
rect 646 16997 680 17031
rect 714 16963 748 16997
rect 782 16964 13396 17032
rect 17984 16998 18086 17032
rect 13431 16964 13465 16998
rect 13500 16964 13534 16998
rect 13569 16964 13603 16998
rect 13638 16964 13672 16998
rect 13707 16964 13741 16998
rect 13776 16964 13810 16998
rect 13845 16964 13879 16998
rect 13914 16964 13948 16998
rect 13983 16964 14017 16998
rect 14052 16964 14086 16998
rect 14121 16964 14155 16998
rect 14190 16964 14224 16998
rect 14259 16964 14293 16998
rect 14328 16964 14362 16998
rect 14397 16964 14431 16998
rect 14466 16964 14500 16998
rect 14535 16964 14569 16998
rect 14604 16964 14638 16998
rect 14673 16964 14707 16998
rect 14742 16964 14776 16998
rect 14811 16964 14845 16998
rect 14880 16964 14914 16998
rect 14949 16964 14983 16998
rect 15018 16964 15052 16998
rect 15087 16964 15121 16998
rect 15156 16964 15190 16998
rect 15225 16964 15259 16998
rect 15294 16964 15328 16998
rect 15363 16964 15397 16998
rect 15432 16964 15466 16998
rect 15501 16964 15535 16998
rect 15570 16964 15604 16998
rect 15639 16964 15673 16998
rect 15708 16964 15742 16998
rect 15777 16964 15811 16998
rect 15846 16964 15880 16998
rect 15915 16964 15949 16998
rect 15984 16964 16018 16998
rect 16053 16964 16087 16998
rect 16122 16964 16156 16998
rect 16191 16964 16225 16998
rect 16260 16964 16294 16998
rect 16329 16964 16363 16998
rect 16398 16964 16432 16998
rect 16467 16964 16501 16998
rect 16536 16964 16570 16998
rect 16605 16964 16639 16998
rect 16674 16964 16708 16998
rect 16743 16964 16777 16998
rect 16812 16964 16846 16998
rect 16881 16964 16915 16998
rect 16950 16964 16984 16998
rect 17019 16964 17053 16998
rect 17088 16964 17122 16998
rect 17157 16964 17191 16998
rect 17226 16964 17260 16998
rect 17295 16964 17329 16998
rect 17364 16964 17398 16998
rect 17433 16964 17467 16998
rect 17502 16964 17536 16998
rect 17571 16964 17605 16998
rect 17640 16964 17674 16998
rect 17709 16964 17743 16998
rect 17778 16964 17812 16998
rect 17847 16964 17881 16998
rect 646 16928 680 16962
rect 714 16894 748 16928
rect 782 16895 816 16929
rect 646 16859 680 16893
rect 714 16825 748 16859
rect 782 16826 816 16860
rect 646 16790 680 16824
rect 714 16756 748 16790
rect 782 16757 816 16791
rect 646 16721 680 16755
rect 10494 16896 10528 16930
rect 10563 16896 10597 16930
rect 10632 16896 10666 16930
rect 10701 16896 10735 16930
rect 10770 16896 10804 16930
rect 10839 16896 10873 16930
rect 10908 16896 10942 16930
rect 10977 16896 11011 16930
rect 11046 16896 11080 16930
rect 11115 16896 11149 16930
rect 11184 16896 11218 16930
rect 11253 16896 11287 16930
rect 11322 16896 11356 16930
rect 11391 16896 11425 16930
rect 11460 16896 11494 16930
rect 11529 16896 11563 16930
rect 11598 16896 11632 16930
rect 11667 16896 11701 16930
rect 11736 16896 11770 16930
rect 11805 16896 11839 16930
rect 11874 16896 11908 16930
rect 11943 16896 11977 16930
rect 12012 16896 12046 16930
rect 12081 16896 12115 16930
rect 12150 16896 12184 16930
rect 12219 16896 12253 16930
rect 12288 16896 12322 16930
rect 12357 16896 12391 16930
rect 12426 16896 12460 16930
rect 12495 16896 12529 16930
rect 12564 16896 12598 16930
rect 12633 16896 12667 16930
rect 12702 16896 12736 16930
rect 12771 16896 12805 16930
rect 12840 16896 12874 16930
rect 12909 16896 12943 16930
rect 12978 16896 13012 16930
rect 13047 16896 13081 16930
rect 13116 16896 13150 16930
rect 13185 16896 13219 16930
rect 13254 16896 13288 16930
rect 13323 16896 13357 16930
rect 13392 16896 13426 16930
rect 13461 16896 13495 16930
rect 13530 16896 13564 16930
rect 13599 16896 13633 16930
rect 13668 16896 13702 16930
rect 13737 16896 13771 16930
rect 13806 16896 13840 16930
rect 13875 16896 13909 16930
rect 13944 16896 13978 16930
rect 14013 16896 14047 16930
rect 14082 16896 14116 16930
rect 14151 16896 14185 16930
rect 14220 16896 14254 16930
rect 14289 16896 14323 16930
rect 14358 16896 14392 16930
rect 14427 16896 14461 16930
rect 10494 16828 10528 16862
rect 10563 16828 10597 16862
rect 10632 16828 10666 16862
rect 10701 16828 10735 16862
rect 10770 16828 10804 16862
rect 10839 16828 10873 16862
rect 10908 16828 10942 16862
rect 10977 16828 11011 16862
rect 11046 16828 11080 16862
rect 11115 16828 11149 16862
rect 11184 16828 11218 16862
rect 11253 16828 11287 16862
rect 11322 16828 11356 16862
rect 11391 16828 11425 16862
rect 11460 16828 11494 16862
rect 11529 16828 11563 16862
rect 11598 16828 11632 16862
rect 11667 16828 11701 16862
rect 11736 16828 11770 16862
rect 11805 16828 11839 16862
rect 11874 16828 11908 16862
rect 11943 16828 11977 16862
rect 12012 16828 12046 16862
rect 12081 16828 12115 16862
rect 12150 16828 12184 16862
rect 12219 16828 12253 16862
rect 12288 16828 12322 16862
rect 12357 16828 12391 16862
rect 12426 16828 12460 16862
rect 12495 16828 12529 16862
rect 12564 16828 12598 16862
rect 12633 16828 12667 16862
rect 12702 16828 12736 16862
rect 12771 16828 12805 16862
rect 12840 16828 12874 16862
rect 12909 16828 12943 16862
rect 12978 16828 13012 16862
rect 13047 16828 13081 16862
rect 13116 16828 13150 16862
rect 13185 16828 13219 16862
rect 13254 16828 13288 16862
rect 13323 16828 13357 16862
rect 13392 16828 13426 16862
rect 13461 16828 13495 16862
rect 13530 16828 13564 16862
rect 13599 16828 13633 16862
rect 13668 16828 13702 16862
rect 13737 16828 13771 16862
rect 13806 16828 13840 16862
rect 13875 16828 13909 16862
rect 13944 16828 13978 16862
rect 14013 16828 14047 16862
rect 14082 16828 14116 16862
rect 14151 16828 14185 16862
rect 14220 16828 14254 16862
rect 14289 16828 14323 16862
rect 14358 16828 14392 16862
rect 14427 16828 14461 16862
rect 10494 16760 10528 16794
rect 10563 16760 10597 16794
rect 10632 16760 10666 16794
rect 10701 16760 10735 16794
rect 10770 16760 10804 16794
rect 10839 16760 10873 16794
rect 10908 16760 10942 16794
rect 10977 16760 11011 16794
rect 11046 16760 11080 16794
rect 11115 16760 11149 16794
rect 11184 16760 11218 16794
rect 11253 16760 11287 16794
rect 11322 16760 11356 16794
rect 11391 16760 11425 16794
rect 11460 16760 11494 16794
rect 11529 16760 11563 16794
rect 11598 16760 11632 16794
rect 11667 16760 11701 16794
rect 11736 16760 11770 16794
rect 11805 16760 11839 16794
rect 11874 16760 11908 16794
rect 11943 16760 11977 16794
rect 12012 16760 12046 16794
rect 12081 16760 12115 16794
rect 12150 16760 12184 16794
rect 12219 16760 12253 16794
rect 12288 16760 12322 16794
rect 12357 16760 12391 16794
rect 12426 16760 12460 16794
rect 12495 16760 12529 16794
rect 12564 16760 12598 16794
rect 12633 16760 12667 16794
rect 12702 16760 12736 16794
rect 12771 16760 12805 16794
rect 12840 16760 12874 16794
rect 12909 16760 12943 16794
rect 12978 16760 13012 16794
rect 13047 16760 13081 16794
rect 13116 16760 13150 16794
rect 13185 16760 13219 16794
rect 13254 16760 13288 16794
rect 13323 16760 13357 16794
rect 13392 16760 13426 16794
rect 13461 16760 13495 16794
rect 13530 16760 13564 16794
rect 13599 16760 13633 16794
rect 13668 16760 13702 16794
rect 13737 16760 13771 16794
rect 13806 16760 13840 16794
rect 13875 16760 13909 16794
rect 13944 16760 13978 16794
rect 14013 16760 14047 16794
rect 14082 16760 14116 16794
rect 14151 16760 14185 16794
rect 14220 16760 14254 16794
rect 14289 16760 14323 16794
rect 14358 16760 14392 16794
rect 14427 16760 14461 16794
rect 14496 16760 15210 16930
rect 714 16687 748 16721
rect 782 16688 816 16722
rect 646 16652 680 16686
rect 714 16618 748 16652
rect 782 16619 816 16653
rect 646 16583 680 16617
rect 714 16549 748 16583
rect 782 16550 816 16584
rect 646 16514 680 16548
rect 714 16480 748 16514
rect 782 16481 816 16515
rect 646 16445 680 16479
rect 714 16411 748 16445
rect 782 16412 816 16446
rect 646 16376 680 16410
rect 714 16342 748 16376
rect 782 16343 816 16377
rect 646 16307 680 16341
rect 646 16239 748 16307
rect 782 16274 816 16308
rect 646 12941 816 16239
rect 15260 14788 15430 16930
rect 15464 16870 15498 16904
rect 15532 16870 15566 16904
rect 15600 16870 15634 16904
rect 15464 16798 15498 16832
rect 15532 16798 15566 16832
rect 15600 16798 15634 16832
rect 15464 16726 15498 16760
rect 15532 16726 15566 16760
rect 15600 16726 15634 16760
rect 15464 16654 15498 16688
rect 15532 16654 15566 16688
rect 15600 16654 15634 16688
rect 15464 16582 15498 16616
rect 15532 16582 15566 16616
rect 15600 16582 15634 16616
rect 15464 16510 15498 16544
rect 15532 16510 15566 16544
rect 15600 16510 15634 16544
rect 15464 16438 15498 16472
rect 15532 16438 15566 16472
rect 15600 16438 15634 16472
rect 15464 16366 15498 16400
rect 15532 16366 15566 16400
rect 15600 16366 15634 16400
rect 15464 16294 15498 16328
rect 15532 16294 15566 16328
rect 15600 16294 15634 16328
rect 15464 16221 15498 16255
rect 15532 16221 15566 16255
rect 15600 16221 15634 16255
rect 17916 16624 18086 16998
rect 18052 16590 18086 16624
rect 17916 16555 17950 16589
rect 17984 16555 18018 16589
rect 18052 16522 18086 16556
rect 17916 16486 17950 16520
rect 17984 16486 18018 16520
rect 18052 16454 18086 16488
rect 17916 16417 17950 16451
rect 17984 16417 18018 16451
rect 18052 16386 18086 16420
rect 17916 16348 17950 16382
rect 17984 16348 18018 16382
rect 18052 16318 18086 16352
rect 17916 16279 17950 16313
rect 17984 16279 18018 16313
rect 18052 16250 18086 16284
rect 17916 16210 17950 16244
rect 17984 16210 18018 16244
rect 18052 16182 18086 16216
rect 17916 16141 17950 16175
rect 17984 16141 18018 16175
rect 18052 16114 18086 16148
rect 17916 16072 17950 16106
rect 17984 16072 18018 16106
rect 18052 16046 18086 16080
rect 17916 16003 17950 16037
rect 17984 16003 18018 16037
rect 18052 15978 18086 16012
rect 17916 15934 17950 15968
rect 17984 15934 18018 15968
rect 18052 15910 18086 15944
rect 17916 15865 17950 15899
rect 17984 15865 18018 15899
rect 18052 15842 18086 15876
rect 17916 15796 17950 15830
rect 17984 15796 18018 15830
rect 18052 15774 18086 15808
rect 17916 15727 17950 15761
rect 17984 15727 18018 15761
rect 18052 15706 18086 15740
rect 17916 15658 17950 15692
rect 17984 15658 18018 15692
rect 18052 15638 18086 15672
rect 17916 15589 17950 15623
rect 17984 15589 18018 15623
rect 18052 15570 18086 15604
rect 17916 15520 17950 15554
rect 17984 15520 18018 15554
rect 18052 15502 18086 15536
rect 17916 15451 17950 15485
rect 17984 15451 18018 15485
rect 18052 15434 18086 15468
rect 17916 15382 17950 15416
rect 17984 15382 18018 15416
rect 18052 15366 18086 15400
rect 17916 15313 17950 15347
rect 17984 15313 18018 15347
rect 18052 15298 18086 15332
rect 17916 15244 17950 15278
rect 17984 15244 18018 15278
rect 18052 15230 18086 15264
rect 17916 15175 17950 15209
rect 17984 15175 18018 15209
rect 18052 15162 18086 15196
rect 17916 15106 17950 15140
rect 17984 15106 18018 15140
rect 18052 15094 18086 15128
rect 17916 15037 17950 15071
rect 17984 15037 18018 15071
rect 18052 15026 18086 15060
rect 15260 14719 15294 14753
rect 15328 14719 15362 14753
rect 15396 14719 15430 14753
rect 17916 14968 17950 15002
rect 17984 14968 18018 15002
rect 18052 14958 18086 14992
rect 17916 14899 17950 14933
rect 17984 14899 18018 14933
rect 18052 14890 18086 14924
rect 17916 14830 17950 14864
rect 17984 14830 18018 14864
rect 18052 14822 18086 14856
rect 17916 14761 17950 14795
rect 17984 14761 18018 14795
rect 18052 14754 18086 14788
rect 15260 14650 15294 14684
rect 15328 14650 15362 14684
rect 15396 14650 15430 14684
rect 15260 14581 15294 14615
rect 15328 14581 15362 14615
rect 15396 14581 15430 14615
rect 15260 14512 15294 14546
rect 15328 14512 15362 14546
rect 15396 14512 15430 14546
rect 15260 14443 15294 14477
rect 15328 14443 15362 14477
rect 15396 14443 15430 14477
rect 15260 14374 15294 14408
rect 15328 14374 15362 14408
rect 15396 14374 15430 14408
rect 15396 14306 15430 14340
rect 15396 14235 15430 14269
rect 15396 14164 15430 14198
rect 15396 14093 15430 14127
rect 15396 14022 15430 14056
rect 15396 13951 15430 13985
rect 15396 13880 15430 13914
rect 15396 13809 15430 13843
rect 15396 13738 15430 13772
rect 15396 13667 15430 13701
rect 15396 13596 15430 13630
rect 17916 14692 17950 14726
rect 17984 14692 18018 14726
rect 18052 14686 18086 14720
rect 17916 14623 17950 14657
rect 17984 14623 18018 14657
rect 18052 14618 18086 14652
rect 17916 14554 17950 14588
rect 17984 14554 18018 14588
rect 18052 14550 18086 14584
rect 17916 14485 17950 14519
rect 17984 14485 18018 14519
rect 18052 14482 18086 14516
rect 17916 14416 17950 14450
rect 17984 14416 18018 14450
rect 18052 14414 18086 14448
rect 17916 14347 17950 14381
rect 17984 14347 18018 14381
rect 18052 14346 18086 14380
rect 17916 14278 17950 14312
rect 17984 14278 18018 14312
rect 18052 14278 18086 14312
rect 17916 14209 17950 14243
rect 17984 14209 18018 14243
rect 18052 14209 18086 14243
rect 17916 14140 17950 14174
rect 17984 14140 18018 14174
rect 18052 14140 18086 14174
rect 17916 14071 17950 14105
rect 17984 14071 18018 14105
rect 18052 14071 18086 14105
rect 17916 14002 17950 14036
rect 17984 14002 18018 14036
rect 18052 14002 18086 14036
rect 17916 13933 17950 13967
rect 17984 13933 18018 13967
rect 18052 13933 18086 13967
rect 17916 13864 17950 13898
rect 17984 13864 18018 13898
rect 18052 13864 18086 13898
rect 17916 13795 17950 13829
rect 17984 13795 18018 13829
rect 18052 13795 18086 13829
rect 17916 13726 17950 13760
rect 17984 13726 18018 13760
rect 18052 13726 18086 13760
rect 17916 13657 17950 13691
rect 17984 13657 18018 13691
rect 18052 13657 18086 13691
rect 15396 13525 15430 13559
rect 15396 13454 15430 13488
rect 15396 13383 15430 13417
rect 17916 13588 17950 13622
rect 17984 13588 18018 13622
rect 18052 13588 18086 13622
rect 17916 13519 17950 13553
rect 17984 13519 18018 13553
rect 18052 13519 18086 13553
rect 17916 13450 17950 13484
rect 17984 13450 18018 13484
rect 18052 13450 18086 13484
rect 17916 13381 17950 13415
rect 17984 13381 18018 13415
rect 18052 13381 18086 13415
rect 15396 13312 15430 13346
rect 15396 13241 15430 13275
rect 17916 13312 17950 13346
rect 17984 13312 18018 13346
rect 18052 13312 18086 13346
rect 17916 13243 17950 13277
rect 17984 13243 18018 13277
rect 18052 13243 18086 13277
rect 17916 13174 17950 13208
rect 17984 13174 18018 13208
rect 18052 13174 18086 13208
rect 17916 13105 17950 13139
rect 17984 13105 18018 13139
rect 18052 13105 18086 13139
rect 17916 13036 17950 13070
rect 17984 13036 18018 13070
rect 18052 13036 18086 13070
rect 851 12941 885 12975
rect 920 12941 954 12975
rect 989 12941 1023 12975
rect 1058 12941 1092 12975
rect 1127 12941 1161 12975
rect 1196 12941 1230 12975
rect 1265 12941 1299 12975
rect 1334 12941 1368 12975
rect 1403 12941 1437 12975
rect 1472 12941 1506 12975
rect 1541 12941 1575 12975
rect 1610 12941 1644 12975
rect 1679 12941 1713 12975
rect 1748 12941 1782 12975
rect 1817 12941 1851 12975
rect 1886 12941 1920 12975
rect 1955 12941 1989 12975
rect 2024 12941 2058 12975
rect 2093 12941 2127 12975
rect 2162 12941 2196 12975
rect 2231 12941 2265 12975
rect 2300 12941 2334 12975
rect 2369 12941 2403 12975
rect 646 12907 748 12941
rect 714 12873 748 12907
rect 783 12873 817 12907
rect 852 12873 886 12907
rect 921 12873 955 12907
rect 990 12873 1024 12907
rect 1059 12873 1093 12907
rect 1128 12873 1162 12907
rect 1197 12873 1231 12907
rect 1266 12873 1300 12907
rect 1335 12873 1369 12907
rect 1404 12873 1438 12907
rect 1473 12873 1507 12907
rect 1542 12873 1576 12907
rect 1611 12873 1645 12907
rect 1680 12873 1714 12907
rect 1749 12873 1783 12907
rect 1818 12873 1852 12907
rect 1887 12873 1921 12907
rect 1956 12873 1990 12907
rect 2025 12873 2059 12907
rect 2094 12873 2128 12907
rect 2163 12873 2197 12907
rect 2232 12873 2266 12907
rect 2301 12873 2335 12907
rect 2370 12873 2404 12907
rect 2438 12873 17840 12975
rect 17916 12967 17950 13001
rect 17984 12967 18018 13001
rect 18052 12967 18086 13001
rect 17916 12898 17950 12932
rect 17984 12898 18018 12932
rect 18052 12898 18086 12932
rect 680 12805 714 12839
rect 749 12805 783 12839
rect 818 12805 852 12839
rect 887 12805 921 12839
rect 956 12805 990 12839
rect 1025 12805 1059 12839
rect 1094 12805 1128 12839
rect 1163 12805 1197 12839
rect 1232 12805 1266 12839
rect 1301 12805 1335 12839
rect 1370 12805 1404 12839
rect 1439 12805 1473 12839
rect 1508 12805 1542 12839
rect 1577 12805 1611 12839
rect 1646 12805 1680 12839
rect 1715 12805 1749 12839
rect 1784 12805 1818 12839
rect 1853 12805 1887 12839
rect 1922 12805 1956 12839
rect 1991 12805 2025 12839
rect 2060 12805 2094 12839
rect 2129 12805 2163 12839
rect 2198 12805 2232 12839
rect 2267 12805 2301 12839
rect 2336 12805 2370 12839
rect 2405 12805 2439 12839
rect 2474 12805 2508 12839
rect 2543 12805 2577 12839
rect 2612 12805 2646 12839
rect 2681 12805 2715 12839
rect 2750 12805 2784 12839
rect 2819 12805 2853 12839
rect 2888 12805 2922 12839
rect 2957 12805 2991 12839
rect 3026 12805 3060 12839
rect 3095 12805 3129 12839
rect 3164 12805 3198 12839
rect 3233 12805 3267 12839
rect 3302 12805 3336 12839
rect 3371 12805 3405 12839
rect 3440 12805 3474 12839
rect 3509 12805 3543 12839
rect 3578 12805 3612 12839
rect 3647 12805 3681 12839
rect 3716 12805 3750 12839
rect 3785 12805 3819 12839
rect 3854 12805 3888 12839
rect 3923 12805 3957 12839
rect 3992 12805 4026 12839
rect 4061 12805 4095 12839
rect 4130 12805 4164 12839
rect 4199 12805 4233 12839
rect 4268 12805 4302 12839
rect 4337 12805 4371 12839
rect 4406 12805 4440 12839
rect 4475 12805 4509 12839
rect 4544 12805 4578 12839
rect 4613 12805 4647 12839
rect 4682 12805 17840 12873
rect 17916 12829 17950 12863
rect 17984 12829 18018 12863
rect 18052 12829 18086 12863
rect 18609 12353 18779 17691
rect 18609 12284 18643 12318
rect 18677 12285 18779 12353
rect 18745 12251 18779 12285
rect 18124 12215 18158 12249
rect 18194 12215 18228 12249
rect 18264 12215 18298 12249
rect 18333 12215 18367 12249
rect 18402 12215 18436 12249
rect 18471 12215 18505 12249
rect 18540 12215 18574 12249
rect 18609 12215 18643 12249
rect 18677 12216 18711 12250
rect 18745 12182 18779 12216
rect 18124 12147 18158 12181
rect 18194 12147 18228 12181
rect 18263 12147 18297 12181
rect 18332 12147 18366 12181
rect 18401 12147 18435 12181
rect 18470 12147 18504 12181
rect 18539 12147 18573 12181
rect 18608 12147 18642 12181
rect 18677 12147 18711 12181
rect 18745 12113 18779 12147
rect 18124 12079 18158 12113
rect 18197 12079 18231 12113
rect 18270 12079 18304 12113
rect 18343 12079 18377 12113
rect 18416 12079 18450 12113
rect 18489 12079 18523 12113
rect 18562 12079 18596 12113
rect 18635 12079 18669 12113
<< mvpsubdiffcont >>
rect 10491 3346 10525 3380
rect 10559 3346 10593 3380
rect 10627 3346 10661 3380
rect 10491 3276 10525 3310
rect 10559 3277 10593 3311
rect 10627 3277 10661 3311
rect 10737 3302 12267 3404
rect 12301 3370 12335 3404
rect 12369 3370 12403 3404
rect 12437 3370 12471 3404
rect 12505 3370 12539 3404
rect 12573 3370 12607 3404
rect 12641 3370 12675 3404
rect 12709 3370 12743 3404
rect 12777 3370 12811 3404
rect 12845 3370 12879 3404
rect 12913 3370 12947 3404
rect 12981 3370 13015 3404
rect 13049 3370 13083 3404
rect 13117 3370 13151 3404
rect 13185 3370 13219 3404
rect 13253 3370 13287 3404
rect 13321 3370 13355 3404
rect 13389 3370 13423 3404
rect 13457 3370 13491 3404
rect 13525 3370 13559 3404
rect 13593 3370 13627 3404
rect 13661 3370 13695 3404
rect 13729 3370 13763 3404
rect 13797 3370 13831 3404
rect 13865 3370 13899 3404
rect 13933 3370 13967 3404
rect 14001 3370 14035 3404
rect 14069 3370 14103 3404
rect 14137 3370 14171 3404
rect 14205 3370 14239 3404
rect 14273 3370 14307 3404
rect 14341 3370 14375 3404
rect 14409 3370 14443 3404
rect 14477 3370 14511 3404
rect 14545 3370 14579 3404
rect 14613 3370 14647 3404
rect 14682 3370 14716 3404
rect 14751 3370 14785 3404
rect 14820 3370 14854 3404
rect 14889 3370 14923 3404
rect 14958 3370 14992 3404
rect 15027 3370 15061 3404
rect 15096 3370 15130 3404
rect 15165 3370 15199 3404
rect 15234 3370 15268 3404
rect 15303 3370 15337 3404
rect 15372 3370 15406 3404
rect 15441 3370 15475 3404
rect 12302 3302 12336 3336
rect 12371 3302 12405 3336
rect 12440 3302 12474 3336
rect 12509 3302 12543 3336
rect 12578 3302 12612 3336
rect 12647 3302 12681 3336
rect 12716 3302 12750 3336
rect 12785 3302 12819 3336
rect 12854 3302 12888 3336
rect 12923 3302 12957 3336
rect 12992 3302 13026 3336
rect 13061 3302 13095 3336
rect 13130 3302 13164 3336
rect 13199 3302 13233 3336
rect 13268 3302 13302 3336
rect 13337 3302 13371 3336
rect 13406 3302 13440 3336
rect 13475 3302 13509 3336
rect 13544 3302 13578 3336
rect 13613 3302 13647 3336
rect 13682 3302 13716 3336
rect 13751 3302 13785 3336
rect 13820 3302 13854 3336
rect 13889 3302 13923 3336
rect 13958 3302 13992 3336
rect 14027 3302 14061 3336
rect 14096 3302 14130 3336
rect 14165 3302 14199 3336
rect 14234 3302 14268 3336
rect 14303 3302 14337 3336
rect 14372 3302 14406 3336
rect 14441 3302 14475 3336
rect 14510 3302 14544 3336
rect 14579 3302 14613 3336
rect 14648 3302 14682 3336
rect 14717 3302 14751 3336
rect 14786 3302 14820 3336
rect 14855 3302 14889 3336
rect 14924 3302 14958 3336
rect 14993 3302 15027 3336
rect 15062 3302 15096 3336
rect 15131 3302 15165 3336
rect 15200 3302 15234 3336
rect 15269 3302 15303 3336
rect 15338 3302 15372 3336
rect 15407 3302 15441 3336
rect 10491 3206 10525 3240
rect 10559 3208 10593 3242
rect 10627 3208 10661 3242
rect 10737 3234 12199 3302
rect 12234 3234 12268 3268
rect 12303 3234 12337 3268
rect 12372 3234 12406 3268
rect 12441 3234 12475 3268
rect 12510 3234 12544 3268
rect 12579 3234 12613 3268
rect 12648 3234 12682 3268
rect 12717 3234 12751 3268
rect 12786 3234 12820 3268
rect 12855 3234 12889 3268
rect 12924 3234 12958 3268
rect 12993 3234 13027 3268
rect 13062 3234 13096 3268
rect 13131 3234 13165 3268
rect 13200 3234 13234 3268
rect 13269 3234 13303 3268
rect 13338 3234 13372 3268
rect 13407 3234 13441 3268
rect 13476 3234 13510 3268
rect 13545 3234 13579 3268
rect 13614 3234 13648 3268
rect 13683 3234 13717 3268
rect 13752 3234 13786 3268
rect 13821 3234 13855 3268
rect 13890 3234 13924 3268
rect 13959 3234 13993 3268
rect 14028 3234 14062 3268
rect 14097 3234 14131 3268
rect 14166 3234 14200 3268
rect 14235 3234 14269 3268
rect 14304 3234 14338 3268
rect 14373 3234 14407 3268
rect 14442 3234 14476 3268
rect 14511 3234 14545 3268
rect 14580 3234 14614 3268
rect 14649 3234 14683 3268
rect 14718 3234 14752 3268
rect 14787 3234 14821 3268
rect 14856 3234 14890 3268
rect 14925 3234 14959 3268
rect 14994 3234 15028 3268
rect 15063 3234 15097 3268
rect 15132 3234 15166 3268
rect 15201 3234 15235 3268
rect 15270 3234 15304 3268
rect 15339 3234 15373 3268
rect 10491 3136 10525 3170
rect 10559 3139 10593 3173
rect 10627 3139 10661 3173
rect 10491 3066 10525 3100
rect 10559 3070 10593 3104
rect 10627 3070 10661 3104
rect 10491 2996 10525 3030
rect 10559 3001 10593 3035
rect 10627 3001 10661 3035
rect 10491 2926 10525 2960
rect 10559 2932 10593 2966
rect 10627 2932 10661 2966
rect 10491 2856 10525 2890
rect 10559 2863 10593 2897
rect 10627 2863 10661 2897
rect 10491 2786 10525 2820
rect 10559 2794 10593 2828
rect 10627 2794 10661 2828
rect 10491 2716 10525 2750
rect 10559 2725 10593 2759
rect 10627 2725 10661 2759
rect 10491 2646 10525 2680
rect 10559 2656 10593 2690
rect 10627 2656 10661 2690
rect 10491 2576 10525 2610
rect 10559 2587 10593 2621
rect 10627 2587 10661 2621
rect 10491 2506 10525 2540
rect 10559 2518 10593 2552
rect 10627 2518 10661 2552
rect 10491 2436 10525 2470
rect 10559 2449 10593 2483
rect 10627 2449 10661 2483
rect 10491 2366 10525 2400
rect 10559 2380 10593 2414
rect 10627 2380 10661 2414
rect 10491 2296 10525 2330
rect 10559 2311 10593 2345
rect 10627 2311 10661 2345
rect 10491 2226 10525 2260
rect 10559 2242 10593 2276
rect 10627 2242 10661 2276
rect 10491 2156 10525 2190
rect 10559 2173 10593 2207
rect 10627 2173 10661 2207
rect 10491 2086 10525 2120
rect 10559 2104 10593 2138
rect 10627 2104 10661 2138
rect 10491 2016 10525 2050
rect 10559 2035 10593 2069
rect 10627 2035 10661 2069
rect 10491 1946 10525 1980
rect 10559 1966 10593 2000
rect 10627 1966 10661 2000
rect 10491 1876 10525 1910
rect 10559 1897 10593 1931
rect 10627 1897 10661 1931
rect 10491 1806 10525 1840
rect 10559 1828 10593 1862
rect 10627 1828 10661 1862
rect 10491 1736 10525 1770
rect 10559 1759 10593 1793
rect 10627 1759 10661 1793
rect 10491 1667 10525 1701
rect 10559 1690 10593 1724
rect 10627 1690 10661 1724
rect 10491 1598 10525 1632
rect 10559 1621 10593 1655
rect 10627 1621 10661 1655
rect 10491 1529 10525 1563
rect 10559 1552 10593 1586
rect 10627 1552 10661 1586
rect 10491 1460 10525 1494
rect 10559 1483 10593 1517
rect 10627 1483 10661 1517
rect 10491 1391 10525 1425
rect 10559 1414 10593 1448
rect 10627 1414 10661 1448
rect 10491 1322 10525 1356
rect 10559 1345 10593 1379
rect 10627 1345 10661 1379
rect 10491 1253 10525 1287
rect 10491 1184 10525 1218
rect 10491 1115 10525 1149
rect 10491 1046 10525 1080
rect 10491 977 10525 1011
rect 10491 908 10525 942
rect 10491 839 10525 873
rect 10491 770 10525 804
rect 10491 701 10525 735
rect 10491 632 10525 666
rect 10559 664 10661 1310
rect 15407 3233 15441 3267
rect 15475 3266 15509 3300
rect 15339 3165 15373 3199
rect 15407 3164 15441 3198
rect 15475 3197 15509 3231
rect 15339 3096 15373 3130
rect 15407 3095 15441 3129
rect 15475 3128 15509 3162
rect 15339 3027 15373 3061
rect 15407 3026 15441 3060
rect 15475 3059 15509 3093
rect 15339 2958 15373 2992
rect 15407 2957 15441 2991
rect 15475 2990 15509 3024
rect 15339 2889 15373 2923
rect 15407 2888 15441 2922
rect 15475 2921 15509 2955
rect 15339 2820 15373 2854
rect 15407 2819 15441 2853
rect 15475 2852 15509 2886
rect 15339 2751 15373 2785
rect 15407 2750 15441 2784
rect 15475 2783 15509 2817
rect 15339 2682 15373 2716
rect 15407 2681 15441 2715
rect 15475 2714 15509 2748
rect 15339 2613 15373 2647
rect 15407 2612 15441 2646
rect 15475 2645 15509 2679
rect 15339 2544 15373 2578
rect 15407 2543 15441 2577
rect 15475 2576 15509 2610
rect 15339 2475 15373 2509
rect 15407 2474 15441 2508
rect 15475 2507 15509 2541
rect 15339 2406 15373 2440
rect 15407 2405 15441 2439
rect 15475 2438 15509 2472
rect 15339 2337 15373 2371
rect 15407 2336 15441 2370
rect 15475 2369 15509 2403
rect 15339 2268 15373 2302
rect 15407 2267 15441 2301
rect 15475 2300 15509 2334
rect 15339 2199 15373 2233
rect 15407 2198 15441 2232
rect 15475 2231 15509 2265
rect 15339 2130 15373 2164
rect 15407 2129 15441 2163
rect 15475 2162 15509 2196
rect 15339 2061 15373 2095
rect 15407 2060 15441 2094
rect 15475 2093 15509 2127
rect 15339 1992 15373 2026
rect 15407 1991 15441 2025
rect 15475 2024 15509 2058
rect 15339 1923 15373 1957
rect 15407 1922 15441 1956
rect 15475 1955 15509 1989
rect 15339 1854 15373 1888
rect 15407 1853 15441 1887
rect 15475 1886 15509 1920
rect 15339 1784 15373 1818
rect 15407 1784 15441 1818
rect 15475 1817 15509 1851
rect 15339 1714 15373 1748
rect 15407 1715 15441 1749
rect 15475 1748 15509 1782
rect 15339 1644 15373 1678
rect 15407 1646 15441 1680
rect 15475 1679 15509 1713
rect 15475 1610 15509 1644
rect 15339 1574 15373 1608
rect 15407 1576 15441 1610
rect 15475 1541 15509 1575
rect 15339 1504 15373 1538
rect 15407 1506 15441 1540
rect 15475 1472 15509 1506
rect 15339 1434 15373 1468
rect 15407 1436 15441 1470
rect 15475 1402 15509 1436
rect 15339 1364 15373 1398
rect 15407 1366 15441 1400
rect 15475 1332 15509 1366
rect 15339 1294 15373 1328
rect 15407 1296 15441 1330
rect 15475 1262 15509 1296
rect 15339 1224 15373 1258
rect 15407 1226 15441 1260
rect 15475 1192 15509 1226
rect 15339 1154 15373 1188
rect 15407 1156 15441 1190
rect 15475 1122 15509 1156
rect 15339 1084 15373 1118
rect 15407 1086 15441 1120
rect 15475 1052 15509 1086
rect 15339 1014 15373 1048
rect 15407 1016 15441 1050
rect 15475 982 15509 1016
rect 15339 944 15373 978
rect 15407 946 15441 980
rect 15475 912 15509 946
rect 15339 874 15373 908
rect 15407 876 15441 910
rect 15475 842 15509 876
rect 15339 804 15373 838
rect 15407 806 15441 840
rect 15475 772 15509 806
rect 15339 734 15373 768
rect 15407 736 15441 770
rect 15475 702 15509 736
rect 10696 664 10730 698
rect 10765 664 10799 698
rect 10834 664 10868 698
rect 10903 664 10937 698
rect 10972 664 11006 698
rect 11041 664 11075 698
rect 11110 664 11144 698
rect 11179 664 11213 698
rect 11248 664 11282 698
rect 11317 664 11351 698
rect 11386 664 11420 698
rect 11455 664 11489 698
rect 11524 664 11558 698
rect 11593 664 11627 698
rect 11662 664 11696 698
rect 11731 664 11765 698
rect 11800 664 11834 698
rect 11869 664 11903 698
rect 11938 664 11972 698
rect 12007 630 15373 698
rect 15407 666 15441 700
rect 15475 632 15509 666
rect 10559 596 10593 630
rect 10628 596 10662 630
rect 10697 596 10731 630
rect 10766 596 10800 630
rect 10835 596 10869 630
rect 10904 596 10938 630
rect 10973 596 11007 630
rect 11042 596 11076 630
rect 11111 596 11145 630
rect 11180 596 11214 630
rect 11249 596 11283 630
rect 11318 596 11352 630
rect 11387 596 11421 630
rect 11456 596 11490 630
rect 11525 596 11559 630
rect 11594 596 11628 630
rect 11663 596 11697 630
rect 11732 596 11766 630
rect 11801 596 11835 630
rect 11870 596 11904 630
rect 11939 596 15441 630
rect 11939 562 15407 596
rect 15475 562 15509 596
rect 10525 528 10559 562
rect 10594 528 10628 562
rect 10663 528 10697 562
rect 10732 528 10766 562
rect 10801 528 10835 562
rect 10870 528 10904 562
rect 10939 528 10973 562
rect 11008 528 11042 562
rect 11077 528 11111 562
rect 11146 528 11180 562
rect 11215 528 11249 562
rect 11284 528 11318 562
rect 11353 528 11387 562
rect 11422 528 11456 562
rect 11491 528 11525 562
rect 11560 528 11594 562
rect 11629 528 11663 562
rect 11698 528 11732 562
rect 11767 528 11801 562
rect 11836 528 11870 562
rect 11905 528 15407 562
<< mvnsubdiffcont >>
rect 425 17423 16167 17457
rect 16202 17423 16236 17457
rect 16271 17423 16305 17457
rect 16340 17423 16374 17457
rect 16409 17423 16443 17457
rect 16478 17423 16512 17457
rect 16547 17423 16581 17457
rect 16616 17423 16650 17457
rect 16685 17423 16719 17457
rect 16754 17423 16788 17457
rect 16823 17423 16857 17457
rect 16892 17423 16926 17457
rect 16961 17423 16995 17457
rect 17030 17423 17064 17457
rect 17099 17423 17133 17457
rect 17168 17423 17202 17457
rect 17237 17423 17271 17457
rect 17306 17423 17340 17457
rect 17375 17423 17409 17457
rect 17444 17423 17478 17457
rect 17513 17423 17547 17457
rect 17582 17423 17616 17457
rect 17651 17423 17685 17457
rect 17720 17423 17754 17457
rect 17789 17423 17823 17457
rect 17858 17423 17892 17457
rect 17927 17423 17961 17457
rect 17996 17423 18030 17457
rect 18065 17423 18099 17457
rect 18134 17423 18168 17457
rect 18203 17423 18237 17457
rect 18272 17423 18306 17457
rect 18341 17423 18375 17457
rect 323 17389 357 17423
rect 425 17389 16133 17423
rect 391 17355 16133 17389
rect 16168 17355 16202 17389
rect 16237 17355 16271 17389
rect 16306 17355 16340 17389
rect 16375 17355 16409 17389
rect 16444 17355 16478 17389
rect 16513 17355 16547 17389
rect 16582 17355 16616 17389
rect 16651 17355 16685 17389
rect 16720 17355 16754 17389
rect 16789 17355 16823 17389
rect 16858 17355 16892 17389
rect 16927 17355 16961 17389
rect 16996 17355 17030 17389
rect 17065 17355 17099 17389
rect 17134 17355 17168 17389
rect 17203 17355 17237 17389
rect 17272 17355 17306 17389
rect 17341 17355 17375 17389
rect 17410 17355 17444 17389
rect 17479 17355 17513 17389
rect 17548 17355 17582 17389
rect 17617 17355 17651 17389
rect 17686 17355 17720 17389
rect 17755 17355 17789 17389
rect 17824 17355 17858 17389
rect 17893 17355 17927 17389
rect 17962 17355 17996 17389
rect 18031 17355 18065 17389
rect 18100 17355 18134 17389
rect 18169 17355 18203 17389
rect 18238 17355 18272 17389
rect 18307 17355 18341 17389
rect 323 17320 357 17354
rect 391 17286 425 17320
rect 459 17287 16065 17355
rect 18307 17321 18409 17355
rect 16100 17287 16134 17321
rect 16169 17287 16203 17321
rect 16238 17287 16272 17321
rect 16307 17287 16341 17321
rect 16376 17287 16410 17321
rect 16445 17287 16479 17321
rect 16514 17287 16548 17321
rect 16583 17287 16617 17321
rect 16652 17287 16686 17321
rect 16721 17287 16755 17321
rect 16790 17287 16824 17321
rect 16859 17287 16893 17321
rect 16928 17287 16962 17321
rect 16997 17287 17031 17321
rect 17066 17287 17100 17321
rect 17135 17287 17169 17321
rect 17204 17287 17238 17321
rect 17273 17287 17307 17321
rect 17342 17287 17376 17321
rect 17411 17287 17445 17321
rect 17480 17287 17514 17321
rect 17549 17287 17583 17321
rect 17618 17287 17652 17321
rect 17687 17287 17721 17321
rect 17756 17287 17790 17321
rect 17825 17287 17859 17321
rect 17894 17287 17928 17321
rect 17963 17287 17997 17321
rect 18032 17287 18066 17321
rect 18101 17287 18135 17321
rect 18170 17287 18204 17321
rect 323 17251 357 17285
rect 391 17217 425 17251
rect 459 17218 493 17252
rect 323 17182 357 17216
rect 391 17148 425 17182
rect 459 17149 493 17183
rect 323 17113 357 17147
rect 391 17079 425 17113
rect 459 17080 493 17114
rect 323 17044 357 17078
rect 391 17010 425 17044
rect 459 17011 493 17045
rect 323 16975 357 17009
rect 391 16941 425 16975
rect 459 16942 493 16976
rect 323 16906 357 16940
rect 391 16872 425 16906
rect 459 16873 493 16907
rect 323 16837 357 16871
rect 391 16803 425 16837
rect 459 16804 493 16838
rect 323 16768 357 16802
rect 323 16699 357 16733
rect 323 16630 357 16664
rect 323 16561 357 16595
rect 323 16492 357 16526
rect 323 16423 357 16457
rect 323 16354 357 16388
rect 323 16285 357 16319
rect 323 16216 357 16250
rect 323 16147 357 16181
rect 323 16078 357 16112
rect 323 16009 357 16043
rect 323 15940 357 15974
rect 323 15871 357 15905
rect 323 15802 357 15836
rect 323 15733 357 15767
rect 323 15664 357 15698
rect 323 15595 357 15629
rect 323 15526 357 15560
rect 323 15457 357 15491
rect 323 15388 357 15422
rect 323 15319 357 15353
rect 323 15250 357 15284
rect 323 15181 357 15215
rect 323 15112 357 15146
rect 323 15043 357 15077
rect 323 14974 357 15008
rect 323 14905 357 14939
rect 323 14836 357 14870
rect 323 14767 357 14801
rect 323 14698 357 14732
rect 323 14629 357 14663
rect 323 14560 357 14594
rect 391 14525 493 16769
rect 323 13947 493 14525
rect 323 13845 357 13879
rect 391 13845 425 13879
rect 459 13845 493 13879
rect 323 13775 357 13809
rect 391 13776 425 13810
rect 459 13776 493 13810
rect 323 13705 357 13739
rect 391 13707 425 13741
rect 459 13707 493 13741
rect 323 13635 357 13669
rect 323 13565 357 13599
rect 323 13495 357 13529
rect 323 13425 357 13459
rect 323 13355 357 13389
rect 323 13285 357 13319
rect 323 13215 357 13249
rect 323 13145 357 13179
rect 323 13075 357 13109
rect 323 13005 357 13039
rect 323 12935 357 12969
rect 323 12865 357 12899
rect 323 12795 357 12829
rect 323 12725 357 12759
rect 323 12655 357 12689
rect 323 12586 357 12620
rect 391 12618 493 13672
rect 18239 15723 18409 17321
rect 18239 15654 18273 15688
rect 18307 15655 18409 15723
rect 18375 15621 18409 15655
rect 18239 15585 18273 15619
rect 18307 15586 18341 15620
rect 18375 15552 18409 15586
rect 18239 15516 18273 15550
rect 18307 15517 18341 15551
rect 18375 15483 18409 15517
rect 18239 15447 18273 15481
rect 18307 15448 18341 15482
rect 18375 15414 18409 15448
rect 18239 15378 18273 15412
rect 18307 15379 18341 15413
rect 18375 15345 18409 15379
rect 18239 15309 18273 15343
rect 18307 15310 18341 15344
rect 18375 15276 18409 15310
rect 18239 15240 18273 15274
rect 18307 15241 18341 15275
rect 18375 15207 18409 15241
rect 18239 15171 18273 15205
rect 18307 15172 18341 15206
rect 18375 15138 18409 15172
rect 18239 15102 18273 15136
rect 18307 15103 18341 15137
rect 18375 15069 18409 15103
rect 18239 15033 18273 15067
rect 18307 15034 18341 15068
rect 18375 15000 18409 15034
rect 18239 14964 18273 14998
rect 18307 14965 18341 14999
rect 18375 14931 18409 14965
rect 18239 14895 18273 14929
rect 18307 14896 18341 14930
rect 18375 14862 18409 14896
rect 18239 14826 18273 14860
rect 18307 14827 18341 14861
rect 18375 14793 18409 14827
rect 18239 14757 18273 14791
rect 18307 14758 18341 14792
rect 18375 14724 18409 14758
rect 18239 14688 18273 14722
rect 18307 14689 18341 14723
rect 18375 14655 18409 14689
rect 18239 14619 18273 14653
rect 18307 14620 18341 14654
rect 18375 14586 18409 14620
rect 18239 14550 18273 14584
rect 18307 14551 18341 14585
rect 18375 14517 18409 14551
rect 18239 14481 18273 14515
rect 18307 14482 18341 14516
rect 18375 14448 18409 14482
rect 18239 14412 18273 14446
rect 18307 14413 18341 14447
rect 18375 14379 18409 14413
rect 18239 14343 18273 14377
rect 18307 14344 18341 14378
rect 18375 14310 18409 14344
rect 18239 14274 18273 14308
rect 18307 14275 18341 14309
rect 18375 14241 18409 14275
rect 18239 14205 18273 14239
rect 18307 14206 18341 14240
rect 18375 14172 18409 14206
rect 18239 14136 18273 14170
rect 18307 14137 18341 14171
rect 18375 14103 18409 14137
rect 18239 14067 18273 14101
rect 18307 14068 18341 14102
rect 18375 14034 18409 14068
rect 18239 13998 18273 14032
rect 18307 13999 18341 14033
rect 18375 13965 18409 13999
rect 18239 13929 18273 13963
rect 18307 13930 18341 13964
rect 18375 13896 18409 13930
rect 18239 13860 18273 13894
rect 18307 13861 18341 13895
rect 18375 13827 18409 13861
rect 18239 13791 18273 13825
rect 18307 13792 18341 13826
rect 18375 13758 18409 13792
rect 18239 13722 18273 13756
rect 18307 13723 18341 13757
rect 18375 13689 18409 13723
rect 18239 13653 18273 13687
rect 18307 13654 18341 13688
rect 18375 13620 18409 13654
rect 18239 13584 18273 13618
rect 18307 13585 18341 13619
rect 18375 13551 18409 13585
rect 18239 13515 18273 13549
rect 18307 13516 18341 13550
rect 18375 13482 18409 13516
rect 18239 13446 18273 13480
rect 18307 13447 18341 13481
rect 18375 13413 18409 13447
rect 18239 13377 18273 13411
rect 18307 13378 18341 13412
rect 18375 13344 18409 13378
rect 18239 13308 18273 13342
rect 18307 13309 18341 13343
rect 18375 13275 18409 13309
rect 18239 13239 18273 13273
rect 18307 13240 18341 13274
rect 18375 13206 18409 13240
rect 18239 13170 18273 13204
rect 18307 13171 18341 13205
rect 18375 13137 18409 13171
rect 18239 13101 18273 13135
rect 18307 13102 18341 13136
rect 18375 13068 18409 13102
rect 18239 13032 18273 13066
rect 18307 13033 18341 13067
rect 18375 12999 18409 13033
rect 18239 12963 18273 12997
rect 18307 12964 18341 12998
rect 18375 12930 18409 12964
rect 18239 12894 18273 12928
rect 18307 12895 18341 12929
rect 18375 12861 18409 12895
rect 18239 12825 18273 12859
rect 18307 12826 18341 12860
rect 18375 12792 18409 12826
rect 18239 12756 18273 12790
rect 18307 12757 18341 12791
rect 18375 12723 18409 12757
rect 18239 12687 18273 12721
rect 18307 12688 18341 12722
rect 18375 12654 18409 12688
rect 528 12618 562 12652
rect 597 12618 631 12652
rect 666 12618 700 12652
rect 735 12618 769 12652
rect 804 12618 838 12652
rect 873 12618 907 12652
rect 942 12618 976 12652
rect 1011 12618 1045 12652
rect 1080 12618 1114 12652
rect 1149 12618 1183 12652
rect 1218 12618 1252 12652
rect 1287 12618 1321 12652
rect 1356 12618 1390 12652
rect 1425 12618 1459 12652
rect 1494 12618 1528 12652
rect 1563 12618 1597 12652
rect 1632 12618 1666 12652
rect 1701 12618 1735 12652
rect 1770 12618 1804 12652
rect 1839 12618 1873 12652
rect 1908 12618 1942 12652
rect 1977 12618 2011 12652
rect 2046 12618 2080 12652
rect 2115 12618 2149 12652
rect 2184 12618 2218 12652
rect 2253 12618 2287 12652
rect 2322 12618 2356 12652
rect 2391 12618 2425 12652
rect 2460 12618 2494 12652
rect 2529 12618 2563 12652
rect 2598 12618 2632 12652
rect 2667 12584 18273 12652
rect 18307 12619 18341 12653
rect 18375 12585 18409 12619
rect 391 12550 425 12584
rect 460 12550 494 12584
rect 529 12550 563 12584
rect 598 12550 632 12584
rect 667 12550 701 12584
rect 736 12550 770 12584
rect 805 12550 839 12584
rect 874 12550 908 12584
rect 943 12550 977 12584
rect 1012 12550 1046 12584
rect 1081 12550 1115 12584
rect 1150 12550 1184 12584
rect 1219 12550 1253 12584
rect 1288 12550 1322 12584
rect 1357 12550 1391 12584
rect 1426 12550 1460 12584
rect 1495 12550 1529 12584
rect 1564 12550 1598 12584
rect 1633 12550 1667 12584
rect 1702 12550 1736 12584
rect 1771 12550 1805 12584
rect 1840 12550 1874 12584
rect 1909 12550 1943 12584
rect 1978 12550 2012 12584
rect 2047 12550 2081 12584
rect 2116 12550 2150 12584
rect 2185 12550 2219 12584
rect 2254 12550 2288 12584
rect 2323 12550 2357 12584
rect 2392 12550 2426 12584
rect 2461 12550 2495 12584
rect 2530 12550 2564 12584
rect 2599 12550 18341 12584
rect 2599 12516 18307 12550
rect 18375 12516 18409 12550
rect 357 12482 391 12516
rect 426 12482 460 12516
rect 495 12482 529 12516
rect 564 12482 598 12516
rect 633 12482 667 12516
rect 702 12482 736 12516
rect 771 12482 805 12516
rect 840 12482 874 12516
rect 909 12482 943 12516
rect 978 12482 1012 12516
rect 1047 12482 1081 12516
rect 1116 12482 1150 12516
rect 1185 12482 1219 12516
rect 1254 12482 1288 12516
rect 1323 12482 1357 12516
rect 1392 12482 1426 12516
rect 1461 12482 1495 12516
rect 1530 12482 1564 12516
rect 1599 12482 1633 12516
rect 1668 12482 1702 12516
rect 1737 12482 1771 12516
rect 1806 12482 1840 12516
rect 1875 12482 1909 12516
rect 1944 12482 1978 12516
rect 2013 12482 2047 12516
rect 2082 12482 2116 12516
rect 2151 12482 2185 12516
rect 2220 12482 2254 12516
rect 2289 12482 2323 12516
rect 2358 12482 2392 12516
rect 2427 12482 2461 12516
rect 2496 12482 2530 12516
rect 2565 12482 18307 12516
rect 10237 3692 14555 3726
rect 14590 3692 14624 3726
rect 14659 3692 14693 3726
rect 14728 3692 14762 3726
rect 14797 3692 14831 3726
rect 14866 3692 14900 3726
rect 14935 3692 14969 3726
rect 15004 3692 15038 3726
rect 15073 3692 15107 3726
rect 15142 3692 15176 3726
rect 15211 3692 15245 3726
rect 15280 3692 15314 3726
rect 15349 3692 15383 3726
rect 15418 3692 15452 3726
rect 15487 3692 15521 3726
rect 15556 3692 15590 3726
rect 15625 3692 15659 3726
rect 15694 3692 15728 3726
rect 15763 3692 15797 3726
rect 10135 3658 10169 3692
rect 10237 3658 14521 3692
rect 10203 3624 14521 3658
rect 14556 3624 14590 3658
rect 14625 3624 14659 3658
rect 14694 3624 14728 3658
rect 14763 3624 14797 3658
rect 14832 3624 14866 3658
rect 14901 3624 14935 3658
rect 14970 3624 15004 3658
rect 15039 3624 15073 3658
rect 15108 3624 15142 3658
rect 15177 3624 15211 3658
rect 15246 3624 15280 3658
rect 15315 3624 15349 3658
rect 15384 3624 15418 3658
rect 15453 3624 15487 3658
rect 15522 3624 15556 3658
rect 15591 3624 15625 3658
rect 15660 3624 15694 3658
rect 15729 3624 15763 3658
rect 10135 3583 10169 3617
rect 10203 3553 10237 3587
rect 10271 3556 14453 3624
rect 15797 3590 15831 3624
rect 14488 3556 14522 3590
rect 14557 3556 14591 3590
rect 14626 3556 14660 3590
rect 14695 3556 14729 3590
rect 14764 3556 14798 3590
rect 14833 3556 14867 3590
rect 14902 3556 14936 3590
rect 14971 3556 15005 3590
rect 15040 3556 15074 3590
rect 15109 3556 15143 3590
rect 15178 3556 15212 3590
rect 15247 3556 15281 3590
rect 15316 3556 15350 3590
rect 15385 3556 15419 3590
rect 15454 3556 15488 3590
rect 15523 3556 15557 3590
rect 15592 3556 15626 3590
rect 15661 3556 15695 3590
rect 10135 3509 10169 3543
rect 10203 3482 10237 3516
rect 10271 3485 10305 3519
rect 10135 3435 10169 3469
rect 10203 3411 10237 3445
rect 10271 3414 10305 3448
rect 15729 3555 15763 3589
rect 15797 3522 15831 3556
rect 15661 3487 15695 3521
rect 15729 3486 15763 3520
rect 15797 3454 15831 3488
rect 15661 3418 15695 3452
rect 15729 3417 15763 3451
rect 10135 3361 10169 3395
rect 10203 3340 10237 3374
rect 10271 3343 10305 3377
rect 10135 3287 10169 3321
rect 10203 3269 10237 3303
rect 10271 3272 10305 3306
rect 10135 3213 10169 3247
rect 10203 3198 10237 3232
rect 10271 3201 10305 3235
rect 10135 3139 10169 3173
rect 10203 3127 10237 3161
rect 10271 3130 10305 3164
rect 10135 3065 10169 3099
rect 10203 3057 10237 3091
rect 10271 3059 10305 3093
rect 10135 2991 10169 3025
rect 10203 2987 10237 3021
rect 10271 2988 10305 3022
rect 10135 2917 10169 2951
rect 10203 2917 10237 2951
rect 10271 2917 10305 2951
rect 15797 3386 15831 3420
rect 15661 3349 15695 3383
rect 15729 3348 15763 3382
rect 15797 3318 15831 3352
rect 15661 3280 15695 3314
rect 15729 3279 15763 3313
rect 15797 3250 15831 3284
rect 15661 3211 15695 3245
rect 15729 3210 15763 3244
rect 15797 3182 15831 3216
rect 15661 3142 15695 3176
rect 15729 3141 15763 3175
rect 15797 3114 15831 3148
rect 15661 3073 15695 3107
rect 15729 3072 15763 3106
rect 15797 3046 15831 3080
rect 15661 3004 15695 3038
rect 15729 3003 15763 3037
rect 15797 2978 15831 3012
rect 15661 2935 15695 2969
rect 15729 2934 15763 2968
rect 15797 2910 15831 2944
rect 15661 2866 15695 2900
rect 15729 2865 15763 2899
rect 15797 2842 15831 2876
rect 15661 2797 15695 2831
rect 15729 2796 15763 2830
rect 15797 2774 15831 2808
rect 15661 2728 15695 2762
rect 15729 2727 15763 2761
rect 15797 2706 15831 2740
rect 15661 2659 15695 2693
rect 15729 2658 15763 2692
rect 15797 2638 15831 2672
rect 15661 2590 15695 2624
rect 15729 2589 15763 2623
rect 15797 2570 15831 2604
rect 15661 2521 15695 2555
rect 15729 2520 15763 2554
rect 15797 2502 15831 2536
rect 15661 2452 15695 2486
rect 15729 2451 15763 2485
rect 15797 2434 15831 2468
rect 15661 2383 15695 2417
rect 15729 2382 15763 2416
rect 15797 2366 15831 2400
rect 15661 2314 15695 2348
rect 15729 2313 15763 2347
rect 15797 2297 15831 2331
rect 15661 2245 15695 2279
rect 15729 2244 15763 2278
rect 15797 2228 15831 2262
rect 15661 2176 15695 2210
rect 15729 2175 15763 2209
rect 15797 2159 15831 2193
rect 15661 2107 15695 2141
rect 15729 2106 15763 2140
rect 15797 2090 15831 2124
rect 15661 2038 15695 2072
rect 15729 2037 15763 2071
rect 15797 2021 15831 2055
rect 15661 1969 15695 2003
rect 15729 1968 15763 2002
rect 15797 1952 15831 1986
rect 15661 1900 15695 1934
rect 15729 1899 15763 1933
rect 15797 1883 15831 1917
rect 15661 1831 15695 1865
rect 15729 1830 15763 1864
rect 15797 1814 15831 1848
rect 15661 1762 15695 1796
rect 15729 1761 15763 1795
rect 15797 1745 15831 1779
rect 15661 1693 15695 1727
rect 15729 1692 15763 1726
rect 15797 1676 15831 1710
rect 15661 1624 15695 1658
rect 15729 1623 15763 1657
rect 15797 1607 15831 1641
rect 15661 1555 15695 1589
rect 15729 1554 15763 1588
rect 15797 1538 15831 1572
rect 15661 1486 15695 1520
rect 15729 1485 15763 1519
rect 15797 1469 15831 1503
rect 15661 1416 15695 1450
rect 15729 1416 15763 1450
rect 15797 1400 15831 1434
rect 15661 1346 15695 1380
rect 15729 1346 15763 1380
rect 15797 1331 15831 1365
rect 15661 1276 15695 1310
rect 15729 1276 15763 1310
rect 15797 1262 15831 1296
rect 15661 1206 15695 1240
rect 15729 1206 15763 1240
rect 15797 1193 15831 1227
rect 15661 1136 15695 1170
rect 15729 1136 15763 1170
rect 15797 1124 15831 1158
rect 15661 1066 15695 1100
rect 15729 1066 15763 1100
rect 15797 1055 15831 1089
rect 15661 996 15695 1030
rect 15729 996 15763 1030
rect 15797 986 15831 1020
rect 15661 926 15695 960
rect 15729 926 15763 960
rect 15797 917 15831 951
rect 15661 856 15695 890
rect 15729 856 15763 890
rect 15797 848 15831 882
rect 15661 786 15695 820
rect 15729 786 15763 820
rect 15797 779 15831 813
rect 15661 716 15695 750
rect 15729 716 15763 750
rect 15797 710 15831 744
rect 15661 646 15695 680
rect 15729 646 15763 680
rect 15797 641 15831 675
rect 15661 576 15695 610
rect 15729 576 15763 610
rect 15797 572 15831 606
rect 15661 506 15695 540
rect 15729 506 15763 540
rect 15797 503 15831 537
rect 15661 436 15695 470
rect 15729 436 15763 470
rect 15797 434 15831 468
rect 15661 366 15695 400
rect 15729 366 15763 400
rect 15797 365 15831 399
rect 15661 296 15695 330
rect 15729 296 15763 330
rect 15797 296 15831 330
<< poly >>
rect 12702 15900 12768 15916
rect 12702 15866 12718 15900
rect 12752 15866 12768 15900
rect 12702 15803 12768 15866
rect 12702 15769 12718 15803
rect 12752 15769 12768 15803
rect 12702 15706 12768 15769
rect 12702 15672 12718 15706
rect 12752 15672 12768 15706
rect 12702 15656 12768 15672
rect 15058 15900 15124 15916
rect 15058 15866 15074 15900
rect 15108 15866 15124 15900
rect 15058 15803 15124 15866
rect 15058 15769 15074 15803
rect 15108 15769 15124 15803
rect 15058 15706 15124 15769
rect 15058 15672 15074 15706
rect 15108 15672 15124 15706
rect 15058 15656 15124 15672
rect 10346 14948 10393 15428
rect 15058 15412 15124 15428
rect 15058 15378 15074 15412
rect 15108 15378 15124 15412
rect 15058 15315 15124 15378
rect 15058 15281 15074 15315
rect 15108 15281 15124 15315
rect 15058 15218 15124 15281
rect 15058 15184 15074 15218
rect 15108 15184 15124 15218
rect 15058 15168 15124 15184
rect 15622 16065 15688 16081
rect 15622 16031 15638 16065
rect 15672 16031 15688 16065
rect 15622 15968 15688 16031
rect 15622 15934 15638 15968
rect 15672 15934 15688 15968
rect 15622 15871 15688 15934
rect 15622 15837 15638 15871
rect 15672 15837 15688 15871
rect 15622 15821 15688 15837
rect 15622 14969 15688 14985
rect 15622 14935 15638 14969
rect 15672 14935 15688 14969
rect 15622 14872 15688 14935
rect 15622 14838 15638 14872
rect 15672 14838 15688 14872
rect 15622 14775 15688 14838
rect 15622 14741 15638 14775
rect 15672 14741 15688 14775
rect 15622 14725 15688 14741
rect 10346 13366 10393 13846
rect 15058 13830 15124 13846
rect 15058 13796 15074 13830
rect 15108 13796 15124 13830
rect 15058 13733 15124 13796
rect 15058 13699 15074 13733
rect 15108 13699 15124 13733
rect 15058 13636 15124 13699
rect 15058 13602 15074 13636
rect 15108 13602 15124 13636
rect 15058 13586 15124 13602
rect 15622 13607 15688 13623
rect 15622 13573 15638 13607
rect 15672 13573 15688 13607
rect 15622 13510 15688 13573
rect 15622 13476 15638 13510
rect 15672 13476 15688 13510
rect 15622 13413 15688 13476
rect 15622 13379 15638 13413
rect 15672 13379 15688 13413
rect 15622 13363 15688 13379
rect 12969 13138 13037 13171
rect 12969 13104 12985 13138
rect 13019 13104 13037 13138
rect 12969 13071 13037 13104
rect 15177 13138 15245 13171
rect 15177 13104 15195 13138
rect 15229 13104 15245 13138
rect 15177 13071 15245 13104
rect 10795 399 10863 432
rect 10795 365 10811 399
rect 10845 365 10863 399
rect 10795 332 10863 365
rect 13003 399 13071 432
rect 13003 365 13021 399
rect 13055 365 13071 399
rect 13003 332 13071 365
<< polycont >>
rect 12718 15866 12752 15900
rect 12718 15769 12752 15803
rect 12718 15672 12752 15706
rect 15074 15866 15108 15900
rect 15074 15769 15108 15803
rect 15074 15672 15108 15706
rect 15074 15378 15108 15412
rect 15074 15281 15108 15315
rect 15074 15184 15108 15218
rect 15638 16031 15672 16065
rect 15638 15934 15672 15968
rect 15638 15837 15672 15871
rect 15638 14935 15672 14969
rect 15638 14838 15672 14872
rect 15638 14741 15672 14775
rect 15074 13796 15108 13830
rect 15074 13699 15108 13733
rect 15074 13602 15108 13636
rect 15638 13573 15672 13607
rect 15638 13476 15672 13510
rect 15638 13379 15672 13413
rect 12985 13104 13019 13138
rect 15195 13104 15229 13138
rect 10811 365 10845 399
rect 13021 365 13055 399
<< locali >>
rect 0 17793 102 17827
rect 15640 17793 15675 17827
rect 15709 17793 15744 17827
rect 15778 17793 15813 17827
rect 15847 17793 15882 17827
rect 15916 17793 15951 17827
rect 15985 17793 16020 17827
rect 16054 17793 16089 17827
rect 16123 17793 16158 17827
rect 16192 17793 16227 17827
rect 16261 17793 16296 17827
rect 16330 17793 16365 17827
rect 16399 17793 16434 17827
rect 16468 17793 16503 17827
rect 16537 17793 16572 17827
rect 16606 17793 16641 17827
rect 16675 17793 16710 17827
rect 16744 17793 16779 17827
rect 16813 17793 16848 17827
rect 16882 17793 16917 17827
rect 16951 17793 16986 17827
rect 17020 17793 17055 17827
rect 17089 17793 17124 17827
rect 17158 17793 17193 17827
rect 17227 17793 17262 17827
rect 17296 17793 17331 17827
rect 17365 17793 17400 17827
rect 17434 17793 17469 17827
rect 17503 17793 17538 17827
rect 17572 17793 17607 17827
rect 17641 17793 17676 17827
rect 17710 17793 17745 17827
rect 17779 17793 17814 17827
rect 17848 17793 17883 17827
rect 17917 17793 17952 17827
rect 17986 17793 18021 17827
rect 18055 17793 18090 17827
rect 18124 17793 18159 17827
rect 18193 17793 18228 17827
rect 18262 17793 18297 17827
rect 18331 17793 18366 17827
rect 18400 17793 18435 17827
rect 18469 17793 18504 17827
rect 18538 17793 18573 17827
rect 18607 17793 18642 17827
rect 18676 17793 18711 17827
rect 18745 17793 18779 17827
rect 34 17759 102 17793
rect 15606 17759 18779 17793
rect 0 17725 68 17759
rect 15606 17725 15641 17759
rect 15675 17725 15710 17759
rect 15744 17725 15779 17759
rect 15813 17725 15848 17759
rect 15882 17725 15917 17759
rect 15951 17725 15986 17759
rect 16020 17725 16055 17759
rect 16089 17725 16124 17759
rect 16158 17725 16193 17759
rect 16227 17725 16262 17759
rect 16296 17725 16331 17759
rect 16365 17725 16400 17759
rect 16434 17725 16469 17759
rect 16503 17725 16538 17759
rect 16572 17725 16607 17759
rect 16641 17725 16676 17759
rect 16710 17725 16745 17759
rect 16779 17725 16814 17759
rect 16848 17725 16883 17759
rect 16917 17725 16952 17759
rect 16986 17725 17021 17759
rect 17055 17725 17090 17759
rect 17124 17725 17159 17759
rect 17193 17725 17228 17759
rect 17262 17725 17297 17759
rect 17331 17725 17366 17759
rect 17400 17725 17435 17759
rect 17469 17725 17504 17759
rect 17538 17725 17573 17759
rect 17607 17725 17642 17759
rect 17676 17725 17711 17759
rect 17745 17725 17780 17759
rect 17814 17725 17849 17759
rect 17883 17725 17918 17759
rect 17952 17725 17987 17759
rect 18021 17725 18056 17759
rect 18090 17725 18125 17759
rect 18159 17725 18194 17759
rect 18228 17725 18263 17759
rect 18297 17725 18332 17759
rect 18366 17725 18401 17759
rect 18435 17725 18470 17759
rect 18504 17725 18539 17759
rect 18573 17725 18608 17759
rect 18642 17725 18677 17759
rect 18711 17725 18779 17759
rect 0 17723 136 17725
rect 34 17690 136 17723
rect 34 17689 68 17690
rect 0 17656 68 17689
rect 102 17657 136 17690
rect 15538 17691 18677 17725
rect 15538 17657 15573 17691
rect 15607 17657 15642 17691
rect 15676 17657 15711 17691
rect 15745 17657 15780 17691
rect 15814 17657 15849 17691
rect 15883 17657 15918 17691
rect 15952 17657 15987 17691
rect 16021 17657 16056 17691
rect 16090 17657 16125 17691
rect 16159 17657 16194 17691
rect 16228 17657 16263 17691
rect 16297 17657 16332 17691
rect 16366 17657 16401 17691
rect 16435 17657 16470 17691
rect 16504 17657 16539 17691
rect 16573 17657 16608 17691
rect 16642 17657 16677 17691
rect 16711 17657 16746 17691
rect 16780 17657 16815 17691
rect 16849 17657 16884 17691
rect 16918 17657 16953 17691
rect 16987 17657 17022 17691
rect 17056 17657 17091 17691
rect 17125 17657 17160 17691
rect 17194 17657 17229 17691
rect 17263 17657 17298 17691
rect 17332 17657 17367 17691
rect 17401 17657 17436 17691
rect 17470 17657 17505 17691
rect 17539 17657 17574 17691
rect 17608 17657 17643 17691
rect 17677 17657 17712 17691
rect 17746 17657 17781 17691
rect 17815 17657 17850 17691
rect 17884 17657 17919 17691
rect 17953 17657 17988 17691
rect 18022 17657 18057 17691
rect 18091 17657 18126 17691
rect 18160 17657 18195 17691
rect 18229 17657 18264 17691
rect 18298 17657 18333 17691
rect 18367 17657 18402 17691
rect 18436 17657 18471 17691
rect 18505 17657 18540 17691
rect 18574 17657 18609 17691
rect 102 17656 170 17657
rect 0 17653 170 17656
rect 34 17622 170 17653
rect 34 17621 136 17622
rect 34 17619 68 17621
rect 0 17587 68 17619
rect 102 17588 136 17621
rect 102 17587 170 17588
rect 0 17583 170 17587
rect 34 17553 170 17583
rect 34 17552 136 17553
rect 34 17549 68 17552
rect 0 17518 68 17549
rect 102 17519 136 17552
rect 102 17518 170 17519
rect 0 17513 170 17518
rect 34 17484 170 17513
rect 34 17483 136 17484
rect 34 17479 68 17483
rect 0 17449 68 17479
rect 102 17450 136 17483
rect 102 17449 170 17450
rect 0 17443 170 17449
rect 34 17415 170 17443
rect 34 17414 136 17415
rect 34 17409 68 17414
rect 0 17380 68 17409
rect 102 17381 136 17414
rect 102 17380 170 17381
rect 0 17373 170 17380
rect 34 17346 170 17373
rect 34 17345 136 17346
rect 34 17339 68 17345
rect 0 17311 68 17339
rect 102 17312 136 17345
rect 102 17311 170 17312
rect 0 17303 170 17311
rect 34 17277 170 17303
rect 34 17276 136 17277
rect 34 17269 68 17276
rect 0 17242 68 17269
rect 102 17243 136 17276
rect 102 17242 170 17243
rect 0 17233 170 17242
rect 34 17208 170 17233
rect 34 17207 136 17208
rect 34 17199 68 17207
rect 0 17173 68 17199
rect 102 17174 136 17207
rect 102 17173 170 17174
rect 0 17164 170 17173
rect 34 17139 170 17164
rect 34 17138 136 17139
rect 34 17130 68 17138
rect 0 17104 68 17130
rect 102 17105 136 17138
rect 102 17104 170 17105
rect 0 17095 170 17104
rect 34 17070 170 17095
rect 34 17069 136 17070
rect 34 17061 68 17069
rect 0 17035 68 17061
rect 102 17036 136 17069
rect 102 17035 170 17036
rect 0 17026 170 17035
rect 34 17001 170 17026
rect 34 17000 136 17001
rect 34 16992 68 17000
rect 0 16966 68 16992
rect 102 16967 136 17000
rect 102 16966 170 16967
rect 0 16957 170 16966
rect 34 16932 170 16957
rect 34 16931 136 16932
rect 34 16923 68 16931
rect 0 16897 68 16923
rect 102 16898 136 16931
rect 102 16897 170 16898
rect 0 16888 170 16897
rect 34 16863 170 16888
rect 34 16862 136 16863
rect 34 16854 68 16862
rect 0 16828 68 16854
rect 102 16829 136 16862
rect 102 16828 170 16829
rect 0 16819 170 16828
rect 34 16794 170 16819
rect 34 16793 136 16794
rect 34 16785 68 16793
rect 0 16759 68 16785
rect 102 16760 136 16793
rect 102 16759 170 16760
rect 0 16750 170 16759
rect 34 16725 170 16750
rect 34 16724 136 16725
rect 34 16716 68 16724
rect 0 16690 68 16716
rect 102 16691 136 16724
rect 102 16690 170 16691
rect 0 16681 170 16690
rect 34 16656 170 16681
rect 34 16655 136 16656
rect 34 16647 68 16655
rect 0 16621 68 16647
rect 102 16622 136 16655
rect 102 16621 170 16622
rect 0 16612 170 16621
rect 34 16587 170 16612
rect 34 16586 136 16587
rect 34 16578 68 16586
rect 0 16552 68 16578
rect 102 16553 136 16586
rect 102 16552 170 16553
rect 0 16543 170 16552
rect 34 16518 170 16543
rect 34 16517 136 16518
rect 34 16509 68 16517
rect 0 16483 68 16509
rect 102 16484 136 16517
rect 102 16483 170 16484
rect 0 16474 170 16483
rect 34 16449 170 16474
rect 34 16448 136 16449
rect 34 16440 68 16448
rect 0 16414 68 16440
rect 102 16415 136 16448
rect 102 16414 170 16415
rect 0 16405 170 16414
rect 34 16380 170 16405
rect 34 16379 136 16380
rect 34 16371 68 16379
rect 0 16345 68 16371
rect 102 16346 136 16379
rect 102 16345 170 16346
rect 0 16336 170 16345
rect 34 16311 170 16336
rect 34 16310 136 16311
rect 34 16302 68 16310
rect 0 16276 68 16302
rect 102 16277 136 16310
rect 102 16276 170 16277
rect 0 16267 170 16276
rect 34 16242 170 16267
rect 34 16241 136 16242
rect 34 16233 68 16241
rect 0 16207 68 16233
rect 102 16208 136 16241
rect 102 16207 170 16208
rect 0 16198 170 16207
rect 34 16173 170 16198
rect 34 16172 136 16173
rect 34 16164 68 16172
rect 0 16138 68 16164
rect 102 16139 136 16172
rect 102 16138 170 16139
rect 0 16129 170 16138
rect 34 16104 170 16129
rect 34 16103 136 16104
rect 34 16095 68 16103
rect 0 16069 68 16095
rect 102 16070 136 16103
rect 102 16069 170 16070
rect 0 16060 170 16069
rect 34 16035 170 16060
rect 34 16034 136 16035
rect 34 16026 68 16034
rect 0 16000 68 16026
rect 102 16001 136 16034
rect 102 16000 170 16001
rect 0 15991 170 16000
rect 34 15966 170 15991
rect 34 15965 136 15966
rect 34 15957 68 15965
rect 0 15931 68 15957
rect 102 15932 136 15965
rect 102 15931 170 15932
rect 0 15922 170 15931
rect 34 15897 170 15922
rect 34 15896 136 15897
rect 34 15888 68 15896
rect 0 15862 68 15888
rect 102 15863 136 15896
rect 102 15862 170 15863
rect 0 15853 170 15862
rect 34 15828 170 15853
rect 34 15827 136 15828
rect 34 15819 68 15827
rect 0 15793 68 15819
rect 102 15794 136 15827
rect 102 15793 170 15794
rect 0 15784 170 15793
rect 34 15759 170 15784
rect 34 15758 136 15759
rect 34 15750 68 15758
rect 0 15724 68 15750
rect 102 15725 136 15758
rect 102 15724 170 15725
rect 0 15715 170 15724
rect 34 15690 170 15715
rect 34 15681 68 15690
rect 0 15646 68 15681
rect 34 15612 68 15646
rect 0 15577 68 15612
rect 34 15543 68 15577
rect 0 15508 68 15543
rect 34 15474 68 15508
rect 0 15439 68 15474
rect 34 15405 68 15439
rect 0 15370 68 15405
rect 34 15336 68 15370
rect 0 15301 68 15336
rect 34 15267 68 15301
rect 0 15232 68 15267
rect 34 15198 68 15232
rect 0 15163 68 15198
rect 34 15129 68 15163
rect 0 15094 68 15129
rect 34 15060 68 15094
rect 0 15025 68 15060
rect 34 14991 68 15025
rect 0 14956 68 14991
rect 34 14922 68 14956
rect 0 14887 68 14922
rect 34 14853 68 14887
rect 0 14818 68 14853
rect 34 14784 68 14818
rect 0 14749 68 14784
rect 34 14715 68 14749
rect 0 14680 68 14715
rect 34 14646 68 14680
rect 0 14611 68 14646
rect 34 14577 68 14611
rect 0 14542 68 14577
rect 34 14508 68 14542
rect 0 14473 68 14508
rect 34 14439 68 14473
rect 0 14404 68 14439
rect 34 14370 68 14404
rect 0 14335 68 14370
rect 34 14301 68 14335
rect 0 14266 68 14301
rect 34 14232 68 14266
rect 0 14197 68 14232
rect 34 14163 68 14197
rect 0 14128 68 14163
rect 34 14094 68 14128
rect 0 14059 68 14094
rect 34 14025 68 14059
rect 0 13990 68 14025
rect 34 13956 68 13990
rect 0 13888 170 13956
rect 34 13854 68 13888
rect 102 13854 136 13888
rect 0 13819 170 13854
rect 34 13785 68 13819
rect 102 13785 136 13819
rect 0 13750 170 13785
rect 34 13716 68 13750
rect 102 13716 136 13750
rect 0 13681 170 13716
rect 34 13647 68 13681
rect 102 13647 136 13681
rect 0 13612 170 13647
rect 34 13578 68 13612
rect 102 13578 136 13612
rect 0 13543 170 13578
rect 323 17425 425 17457
rect 16167 17425 16202 17457
rect 16236 17425 16271 17457
rect 16305 17425 16340 17457
rect 16374 17425 16409 17457
rect 16443 17425 16478 17457
rect 16512 17425 16547 17457
rect 323 17423 393 17425
rect 357 17391 393 17423
rect 16543 17423 16547 17425
rect 16581 17423 16616 17457
rect 16650 17423 16685 17457
rect 16719 17423 16754 17457
rect 16788 17423 16823 17457
rect 16857 17423 16892 17457
rect 16926 17423 16961 17457
rect 16995 17425 17030 17457
rect 17064 17425 17099 17457
rect 17133 17425 17168 17457
rect 17202 17425 17237 17457
rect 17271 17425 17306 17457
rect 17340 17425 17375 17457
rect 17409 17425 17444 17457
rect 16997 17423 17030 17425
rect 17071 17423 17099 17425
rect 17145 17423 17168 17425
rect 17219 17423 17237 17425
rect 17293 17423 17306 17425
rect 17367 17423 17375 17425
rect 17441 17423 17444 17425
rect 17478 17425 17513 17457
rect 17547 17425 17582 17457
rect 17616 17425 17651 17457
rect 17685 17425 17720 17457
rect 17754 17425 17789 17457
rect 17823 17425 17858 17457
rect 17478 17423 17481 17425
rect 17547 17423 17555 17425
rect 17616 17423 17630 17425
rect 17685 17423 17705 17425
rect 17754 17423 17780 17425
rect 17823 17423 17855 17425
rect 17892 17423 17927 17457
rect 17961 17425 17996 17457
rect 18030 17425 18065 17457
rect 18099 17425 18134 17457
rect 18168 17425 18203 17457
rect 18237 17425 18272 17457
rect 18306 17425 18341 17457
rect 17964 17423 17996 17425
rect 18039 17423 18065 17425
rect 18114 17423 18134 17425
rect 18189 17423 18203 17425
rect 18264 17423 18272 17425
rect 18339 17423 18341 17425
rect 18375 17423 18409 17457
rect 357 17389 425 17391
rect 323 17355 391 17389
rect 16543 17391 16963 17423
rect 16997 17391 17037 17423
rect 17071 17391 17111 17423
rect 17145 17391 17185 17423
rect 17219 17391 17259 17423
rect 17293 17391 17333 17423
rect 17367 17391 17407 17423
rect 17441 17391 17481 17423
rect 17515 17391 17555 17423
rect 17589 17391 17630 17423
rect 17664 17391 17705 17423
rect 17739 17391 17780 17423
rect 17814 17391 17855 17423
rect 17889 17391 17930 17423
rect 17964 17391 18005 17423
rect 18039 17391 18080 17423
rect 18114 17391 18155 17423
rect 18189 17391 18230 17423
rect 18264 17391 18305 17423
rect 18339 17391 18409 17423
rect 16543 17389 18409 17391
rect 16547 17355 16582 17389
rect 16616 17355 16651 17389
rect 16685 17355 16720 17389
rect 16754 17355 16789 17389
rect 16823 17355 16858 17389
rect 16892 17355 16927 17389
rect 16961 17355 16996 17389
rect 17030 17355 17065 17389
rect 17099 17355 17134 17389
rect 17168 17355 17203 17389
rect 17237 17355 17272 17389
rect 17306 17355 17341 17389
rect 17375 17355 17410 17389
rect 17444 17355 17479 17389
rect 17513 17355 17548 17389
rect 17582 17355 17617 17389
rect 17651 17355 17686 17389
rect 17720 17355 17755 17389
rect 17789 17355 17824 17389
rect 17858 17355 17893 17389
rect 17927 17355 17962 17389
rect 17996 17355 18031 17389
rect 18065 17355 18100 17389
rect 18134 17355 18169 17389
rect 18203 17355 18238 17389
rect 18272 17355 18307 17389
rect 18341 17355 18409 17389
rect 323 17354 459 17355
rect 357 17353 459 17354
rect 357 17320 427 17353
rect 323 17309 391 17320
rect 323 17285 355 17309
rect 389 17286 391 17309
rect 425 17319 427 17320
rect 16543 17353 18307 17355
rect 16543 17321 16963 17353
rect 425 17287 459 17319
rect 16065 17287 16100 17319
rect 16134 17287 16169 17319
rect 16203 17287 16238 17319
rect 16272 17287 16307 17319
rect 16341 17287 16376 17319
rect 16410 17287 16445 17319
rect 16479 17287 16514 17319
rect 16548 17287 16583 17321
rect 16617 17287 16652 17321
rect 16686 17287 16721 17321
rect 16755 17287 16790 17321
rect 16824 17287 16859 17321
rect 16893 17287 16928 17321
rect 16962 17319 16963 17321
rect 16997 17321 17035 17353
rect 17069 17321 17107 17353
rect 17141 17321 17179 17353
rect 17213 17321 17251 17353
rect 17285 17321 17323 17353
rect 17357 17321 17395 17353
rect 17429 17321 17468 17353
rect 17502 17321 17541 17353
rect 17575 17321 17614 17353
rect 17648 17321 17687 17353
rect 17721 17321 17760 17353
rect 17794 17321 17833 17353
rect 17867 17321 17906 17353
rect 17940 17321 17979 17353
rect 18013 17321 18052 17353
rect 18086 17321 18125 17353
rect 18159 17321 18198 17353
rect 18232 17321 18271 17353
rect 18305 17321 18307 17353
rect 16962 17287 16997 17319
rect 17031 17319 17035 17321
rect 17100 17319 17107 17321
rect 17169 17319 17179 17321
rect 17238 17319 17251 17321
rect 17307 17319 17323 17321
rect 17376 17319 17395 17321
rect 17445 17319 17468 17321
rect 17514 17319 17541 17321
rect 17583 17319 17614 17321
rect 17031 17287 17066 17319
rect 17100 17287 17135 17319
rect 17169 17287 17204 17319
rect 17238 17287 17273 17319
rect 17307 17287 17342 17319
rect 17376 17287 17411 17319
rect 17445 17287 17480 17319
rect 17514 17287 17549 17319
rect 17583 17287 17618 17319
rect 17652 17287 17687 17321
rect 17721 17287 17756 17321
rect 17794 17319 17825 17321
rect 17867 17319 17894 17321
rect 17940 17319 17963 17321
rect 18013 17319 18032 17321
rect 18086 17319 18101 17321
rect 18159 17319 18170 17321
rect 18232 17319 18239 17321
rect 17790 17287 17825 17319
rect 17859 17287 17894 17319
rect 17928 17287 17963 17319
rect 17997 17287 18032 17319
rect 18066 17287 18101 17319
rect 18135 17287 18170 17319
rect 18204 17287 18239 17319
rect 425 17286 493 17287
rect 389 17280 493 17286
rect 389 17275 427 17280
rect 357 17251 427 17275
rect 461 17252 493 17280
rect 323 17234 391 17251
rect 323 17216 355 17234
rect 389 17217 391 17234
rect 425 17246 427 17251
rect 425 17218 459 17246
rect 425 17217 493 17218
rect 389 17207 493 17217
rect 389 17200 427 17207
rect 357 17182 427 17200
rect 461 17183 493 17207
rect 323 17158 391 17182
rect 323 17147 355 17158
rect 389 17148 391 17158
rect 425 17173 427 17182
rect 425 17149 459 17173
rect 425 17148 493 17149
rect 389 17134 493 17148
rect 678 17134 716 17140
rect 750 17134 789 17140
rect 823 17134 862 17140
rect 896 17134 935 17140
rect 969 17134 1008 17140
rect 1042 17134 1081 17140
rect 1115 17134 1154 17140
rect 1188 17134 1227 17140
rect 1261 17134 1300 17140
rect 1334 17134 1373 17140
rect 1407 17134 1446 17140
rect 1480 17134 1519 17140
rect 1553 17134 1592 17140
rect 1626 17134 1665 17140
rect 1699 17134 1738 17140
rect 1772 17134 1811 17140
rect 1845 17134 1884 17140
rect 1918 17134 1957 17140
rect 1991 17134 2030 17140
rect 2064 17134 2103 17140
rect 2137 17134 2176 17140
rect 2210 17134 2249 17140
rect 2283 17134 2322 17140
rect 2356 17134 2395 17140
rect 2429 17134 2468 17140
rect 2502 17134 2541 17140
rect 2575 17134 2614 17140
rect 2648 17134 2687 17140
rect 2721 17134 2760 17140
rect 2794 17134 2833 17140
rect 2867 17134 2906 17140
rect 2940 17134 2979 17140
rect 3013 17134 3052 17140
rect 3086 17134 3125 17140
rect 3159 17134 3197 17140
rect 3231 17134 3269 17140
rect 3303 17134 3341 17140
rect 3375 17134 3413 17140
rect 3447 17134 3485 17140
rect 3519 17134 3557 17140
rect 3591 17134 3629 17140
rect 3663 17134 3701 17140
rect 3735 17134 3773 17140
rect 3807 17134 3845 17140
rect 3879 17134 3917 17140
rect 3951 17134 3989 17140
rect 4023 17134 4061 17140
rect 4095 17134 4133 17140
rect 4167 17134 4205 17140
rect 4239 17134 4277 17140
rect 4311 17134 4349 17140
rect 4383 17134 4421 17140
rect 4455 17134 4493 17140
rect 4527 17134 4565 17140
rect 4599 17134 4637 17140
rect 4671 17134 4709 17140
rect 4743 17134 4781 17140
rect 4815 17134 4853 17140
rect 4887 17134 4925 17140
rect 4959 17134 4997 17140
rect 5031 17134 5069 17140
rect 5103 17134 5141 17140
rect 5175 17134 5213 17140
rect 5247 17134 5285 17140
rect 5319 17134 5357 17140
rect 5391 17134 5429 17140
rect 5463 17134 5501 17140
rect 5535 17134 5573 17140
rect 5607 17134 5645 17140
rect 5679 17134 5717 17140
rect 5751 17134 5789 17140
rect 5823 17134 5861 17140
rect 5895 17134 5933 17140
rect 389 17124 427 17134
rect 357 17113 427 17124
rect 461 17114 493 17134
rect 323 17082 391 17113
rect 323 17078 355 17082
rect 389 17079 391 17082
rect 425 17100 427 17113
rect 425 17080 459 17100
rect 425 17079 493 17080
rect 389 17061 493 17079
rect 389 17048 427 17061
rect 357 17044 427 17048
rect 461 17045 493 17061
rect 323 17010 391 17044
rect 425 17027 427 17044
rect 425 17011 459 17027
rect 425 17010 493 17011
rect 323 17009 493 17010
rect 357 17006 493 17009
rect 389 16988 493 17006
rect 389 16975 427 16988
rect 461 16976 493 16988
rect 323 16972 355 16975
rect 389 16972 391 16975
rect 323 16941 391 16972
rect 425 16954 427 16975
rect 425 16942 459 16954
rect 425 16941 493 16942
rect 323 16940 493 16941
rect 357 16930 493 16940
rect 389 16915 493 16930
rect 389 16906 427 16915
rect 461 16907 493 16915
rect 323 16896 355 16906
rect 389 16896 391 16906
rect 323 16872 391 16896
rect 425 16881 427 16906
rect 425 16873 459 16881
rect 425 16872 493 16873
rect 323 16871 493 16872
rect 357 16854 493 16871
rect 389 16842 493 16854
rect 389 16837 427 16842
rect 461 16838 493 16842
rect 323 16820 355 16837
rect 389 16820 391 16837
rect 323 16803 391 16820
rect 425 16808 427 16837
rect 425 16804 459 16808
rect 425 16803 493 16804
rect 323 16802 493 16803
rect 357 16778 493 16802
rect 389 16769 493 16778
rect 323 16744 355 16768
rect 389 16744 391 16769
rect 323 16733 391 16744
rect 357 16702 391 16733
rect 323 16668 355 16699
rect 389 16668 391 16702
rect 323 16664 391 16668
rect 357 16630 391 16664
rect 323 16626 391 16630
rect 323 16595 355 16626
rect 389 16592 391 16626
rect 357 16561 391 16592
rect 323 16550 391 16561
rect 323 16526 355 16550
rect 389 16516 391 16550
rect 357 16492 391 16516
rect 323 16474 391 16492
rect 323 16457 355 16474
rect 389 16440 391 16474
rect 357 16423 391 16440
rect 323 16388 391 16423
rect 357 16354 391 16388
rect 323 16319 391 16354
rect 357 16285 391 16319
rect 323 16250 391 16285
rect 357 16216 391 16250
rect 323 16181 391 16216
rect 357 16147 391 16181
rect 323 16112 391 16147
rect 357 16078 391 16112
rect 323 16043 391 16078
rect 357 16009 391 16043
rect 323 15974 391 16009
rect 357 15940 391 15974
rect 323 15905 391 15940
rect 357 15871 391 15905
rect 323 15847 391 15871
rect 323 15836 357 15847
rect 357 15802 391 15813
rect 323 15773 391 15802
rect 323 15767 357 15773
rect 357 15733 391 15739
rect 323 15699 391 15733
rect 323 15698 357 15699
rect 357 15664 391 15665
rect 323 15629 391 15664
rect 357 15625 391 15629
rect 323 15591 357 15595
rect 323 15560 391 15591
rect 357 15551 391 15560
rect 323 15517 357 15526
rect 323 15491 391 15517
rect 357 15477 391 15491
rect 323 15443 357 15457
rect 323 15422 391 15443
rect 357 15403 391 15422
rect 323 15369 357 15388
rect 323 15353 391 15369
rect 357 15329 391 15353
rect 323 15295 357 15319
rect 323 15284 391 15295
rect 357 15255 391 15284
rect 323 15221 357 15250
rect 323 15215 391 15221
rect 357 15181 391 15215
rect 323 15147 357 15181
rect 323 15146 391 15147
rect 357 15112 391 15146
rect 323 15107 391 15112
rect 323 15077 357 15107
rect 357 15043 391 15073
rect 323 15033 391 15043
rect 323 15008 357 15033
rect 357 14974 391 14999
rect 323 14959 391 14974
rect 323 14939 357 14959
rect 357 14905 391 14925
rect 323 14885 391 14905
rect 323 14870 357 14885
rect 357 14836 391 14851
rect 323 14811 391 14836
rect 323 14801 357 14811
rect 357 14767 391 14777
rect 323 14737 391 14767
rect 323 14732 357 14737
rect 357 14698 391 14703
rect 323 14663 391 14698
rect 323 14594 391 14629
rect 357 14589 391 14594
rect 323 14555 357 14560
rect 323 14525 391 14555
rect 323 13923 493 13947
rect 323 13889 357 13923
rect 391 13889 429 13923
rect 463 13889 493 13923
rect 323 13879 493 13889
rect 357 13850 391 13879
rect 323 13816 357 13845
rect 425 13850 459 13879
rect 425 13845 429 13850
rect 391 13816 429 13845
rect 463 13816 493 13845
rect 323 13810 493 13816
rect 323 13809 391 13810
rect 357 13777 391 13809
rect 323 13743 357 13775
rect 425 13777 459 13810
rect 425 13776 429 13777
rect 391 13743 429 13776
rect 463 13743 493 13776
rect 323 13741 493 13743
rect 323 13739 391 13741
rect 357 13707 391 13739
rect 425 13707 459 13741
rect 357 13705 493 13707
rect 323 13704 493 13705
rect 323 13670 357 13704
rect 391 13672 429 13704
rect 463 13672 493 13704
rect 323 13669 391 13670
rect 357 13635 391 13669
rect 323 13631 391 13635
rect 323 13599 357 13631
rect 357 13565 391 13597
rect 323 13558 391 13565
rect 323 13529 357 13558
rect 357 13495 391 13524
rect 323 13485 391 13495
rect 323 13459 357 13485
rect 357 13425 391 13451
rect 323 13412 391 13425
rect 323 13389 357 13412
rect 357 13355 391 13378
rect 323 13339 391 13355
rect 323 13319 357 13339
rect 357 13285 391 13305
rect 323 13266 391 13285
rect 323 13249 357 13266
rect 357 13215 391 13232
rect 323 13193 391 13215
rect 323 13179 357 13193
rect 357 13145 391 13159
rect 323 13120 391 13145
rect 323 13109 357 13120
rect 357 13075 391 13086
rect 323 13047 391 13075
rect 323 13039 357 13047
rect 357 13005 391 13013
rect 323 12974 391 13005
rect 323 12969 357 12974
rect 357 12935 391 12940
rect 323 12901 391 12935
rect 323 12899 357 12901
rect 357 12865 391 12867
rect 323 12829 391 12865
rect 357 12828 391 12829
rect 323 12794 357 12795
rect 646 17106 716 17134
rect 646 17100 748 17106
rect 680 17066 748 17100
rect 16407 17100 16431 17134
rect 16465 17100 16500 17134
rect 16534 17100 16569 17134
rect 16603 17100 16638 17134
rect 16672 17100 16707 17134
rect 16741 17100 16776 17134
rect 16810 17100 16845 17134
rect 16879 17100 16914 17134
rect 16948 17100 16983 17134
rect 17017 17100 17052 17134
rect 17086 17100 17121 17134
rect 17155 17102 17190 17134
rect 17224 17102 17259 17134
rect 17180 17100 17190 17102
rect 17256 17100 17259 17102
rect 17293 17102 17328 17134
rect 17362 17102 17397 17134
rect 17431 17102 17466 17134
rect 17500 17102 17535 17134
rect 17569 17102 17604 17134
rect 17293 17100 17298 17102
rect 17362 17100 17374 17102
rect 17431 17100 17450 17102
rect 17500 17100 17526 17102
rect 17569 17100 17602 17102
rect 17638 17100 17673 17134
rect 17707 17102 17742 17134
rect 17776 17102 17811 17134
rect 17845 17102 17880 17134
rect 17914 17102 17949 17134
rect 17983 17102 18018 17134
rect 17712 17100 17742 17102
rect 17788 17100 17811 17102
rect 17864 17100 17880 17102
rect 17940 17100 17949 17102
rect 18016 17100 18018 17102
rect 18052 17100 18086 17134
rect 646 17032 714 17066
rect 16407 17068 17146 17100
rect 17180 17068 17222 17100
rect 17256 17068 17298 17100
rect 17332 17068 17374 17100
rect 17408 17068 17450 17100
rect 17484 17068 17526 17100
rect 17560 17068 17602 17100
rect 17636 17068 17678 17100
rect 17712 17068 17754 17100
rect 17788 17068 17830 17100
rect 17864 17068 17906 17100
rect 17940 17068 17982 17100
rect 18016 17068 18086 17100
rect 16407 17066 18086 17068
rect 646 17031 782 17032
rect 680 17028 782 17031
rect 712 16997 782 17028
rect 646 16994 678 16997
rect 712 16994 714 16997
rect 646 16963 714 16994
rect 748 16988 782 16997
rect 748 16963 750 16988
rect 13464 17032 13499 17034
rect 13533 17032 13568 17034
rect 13602 17032 13637 17034
rect 13671 17032 13706 17034
rect 13740 17032 13775 17034
rect 13809 17032 13844 17034
rect 13878 17032 13913 17034
rect 13947 17032 13982 17034
rect 14016 17032 14051 17034
rect 14085 17032 14120 17034
rect 14154 17032 14189 17034
rect 14223 17032 14258 17034
rect 14292 17032 14327 17034
rect 14361 17032 14396 17034
rect 14430 17032 14465 17034
rect 14499 17032 14534 17034
rect 14568 17032 14603 17034
rect 14637 17032 14672 17034
rect 14706 17032 14741 17034
rect 14775 17032 14810 17034
rect 14844 17032 14879 17034
rect 14913 17032 14948 17034
rect 14982 17032 15017 17034
rect 15051 17032 15086 17034
rect 15120 17032 15155 17034
rect 15189 17032 15224 17034
rect 15258 17032 15293 17034
rect 15327 17032 15362 17034
rect 15396 17032 15431 17034
rect 15465 17032 15500 17034
rect 15534 17032 15569 17034
rect 15603 17032 15638 17034
rect 15672 17032 15707 17034
rect 15741 17032 15776 17034
rect 15810 17032 15845 17034
rect 15879 17032 15914 17034
rect 15948 17032 15983 17034
rect 16017 17032 16052 17034
rect 16086 17032 16121 17034
rect 16155 17032 16190 17034
rect 16224 17032 16259 17034
rect 16293 17032 16328 17034
rect 16362 17032 16397 17034
rect 16431 17032 16466 17066
rect 16500 17032 16535 17066
rect 16569 17032 16604 17066
rect 16638 17032 16673 17066
rect 16707 17032 16742 17066
rect 16776 17032 16811 17066
rect 16845 17032 16880 17066
rect 16914 17032 16949 17066
rect 16983 17032 17018 17066
rect 17052 17032 17087 17066
rect 17121 17032 17156 17066
rect 17190 17032 17225 17066
rect 17259 17032 17294 17066
rect 17328 17032 17363 17066
rect 17397 17032 17432 17066
rect 17466 17032 17501 17066
rect 17535 17032 17570 17066
rect 17604 17032 17639 17066
rect 17673 17032 17708 17066
rect 17742 17032 17777 17066
rect 17811 17032 17846 17066
rect 17880 17032 17915 17066
rect 17949 17032 17984 17066
rect 18018 17032 18086 17066
rect 13396 17030 17984 17032
rect 13396 16998 17146 17030
rect 17180 16998 17218 17030
rect 17252 16998 17291 17030
rect 17325 16998 17364 17030
rect 17398 16998 17437 17030
rect 17471 16998 17510 17030
rect 17544 16998 17583 17030
rect 17617 16998 17656 17030
rect 17690 16998 17729 17030
rect 17763 16998 17802 17030
rect 17836 16998 17875 17030
rect 17909 16998 17948 17030
rect 17982 16998 17984 17030
rect 13396 16973 13431 16998
rect 13465 16973 13500 16998
rect 13534 16973 13569 16998
rect 13603 16973 13638 16998
rect 13672 16973 13707 16998
rect 13741 16973 13776 16998
rect 13810 16973 13845 16998
rect 13879 16973 13914 16998
rect 13948 16973 13983 16998
rect 14017 16973 14052 16998
rect 14086 16973 14121 16998
rect 14155 16973 14190 16998
rect 14224 16973 14259 16998
rect 14293 16973 14328 16998
rect 14362 16973 14397 16998
rect 14431 16973 14466 16998
rect 14500 16973 14535 16998
rect 14569 16973 14604 16998
rect 14638 16973 14673 16998
rect 14707 16973 14742 16998
rect 14776 16973 14811 16998
rect 14845 16973 14880 16998
rect 14914 16973 14949 16998
rect 14983 16973 15018 16998
rect 15052 16973 15087 16998
rect 15121 16973 15156 16998
rect 15190 16973 15225 16998
rect 15199 16964 15225 16973
rect 15259 16964 15294 16998
rect 15328 16964 15363 16998
rect 15397 16964 15432 16998
rect 15466 16964 15501 16998
rect 15535 16964 15570 16998
rect 15604 16964 15639 16998
rect 15673 16964 15708 16998
rect 15742 16964 15777 16998
rect 15811 16964 15846 16998
rect 15880 16964 15915 16998
rect 15949 16964 15984 16998
rect 16018 16964 16053 16998
rect 16087 16964 16122 16998
rect 16156 16964 16191 16998
rect 16225 16964 16260 16998
rect 16294 16964 16329 16998
rect 16363 16964 16398 16998
rect 16432 16964 16467 16998
rect 16501 16964 16536 16998
rect 16570 16964 16605 16998
rect 16639 16964 16674 16998
rect 16708 16964 16743 16998
rect 16777 16964 16812 16998
rect 16846 16964 16881 16998
rect 16915 16964 16950 16998
rect 16984 16964 17019 16998
rect 17053 16964 17088 16998
rect 17122 16996 17146 16998
rect 17191 16996 17218 16998
rect 17260 16996 17291 16998
rect 17122 16964 17157 16996
rect 17191 16964 17226 16996
rect 17260 16964 17295 16996
rect 17329 16964 17364 16998
rect 17398 16964 17433 16998
rect 17471 16996 17502 16998
rect 17544 16996 17571 16998
rect 17617 16996 17640 16998
rect 17690 16996 17709 16998
rect 17763 16996 17778 16998
rect 17836 16996 17847 16998
rect 17909 16996 17916 16998
rect 17467 16964 17502 16996
rect 17536 16964 17571 16996
rect 17605 16964 17640 16996
rect 17674 16964 17709 16996
rect 17743 16964 17778 16996
rect 17812 16964 17847 16996
rect 17881 16964 17916 16996
rect 646 16962 750 16963
rect 680 16955 750 16962
rect 712 16954 750 16955
rect 784 16954 816 16964
rect 712 16929 816 16954
rect 712 16928 782 16929
rect 646 16921 678 16928
rect 712 16921 714 16928
rect 646 16894 714 16921
rect 748 16908 782 16928
rect 748 16894 750 16908
rect 646 16893 750 16894
rect 680 16882 750 16893
rect 712 16874 750 16882
rect 784 16874 816 16895
rect 712 16860 816 16874
rect 712 16859 782 16860
rect 646 16848 678 16859
rect 712 16848 714 16859
rect 646 16825 714 16848
rect 748 16828 782 16859
rect 748 16825 750 16828
rect 646 16824 750 16825
rect 680 16808 750 16824
rect 712 16794 750 16808
rect 784 16794 816 16826
rect 712 16791 816 16794
rect 712 16790 782 16791
rect 646 16774 678 16790
rect 712 16774 714 16790
rect 646 16756 714 16774
rect 748 16757 782 16790
rect 748 16756 816 16757
rect 646 16755 816 16756
rect 680 16748 816 16755
rect 680 16734 750 16748
rect 712 16721 750 16734
rect 784 16722 816 16748
rect 646 16700 678 16721
rect 712 16700 714 16721
rect 646 16687 714 16700
rect 748 16714 750 16721
rect 748 16688 782 16714
rect 748 16687 816 16688
rect 646 16686 816 16687
rect 680 16667 816 16686
rect 680 16660 750 16667
rect 712 16652 750 16660
rect 784 16653 816 16667
rect 646 16626 678 16652
rect 712 16626 714 16652
rect 646 16618 714 16626
rect 748 16633 750 16652
rect 748 16619 782 16633
rect 748 16618 816 16619
rect 646 16617 816 16618
rect 680 16586 816 16617
rect 712 16583 750 16586
rect 784 16584 816 16586
rect 646 16552 678 16583
rect 712 16552 714 16583
rect 646 16549 714 16552
rect 748 16552 750 16583
rect 748 16550 782 16552
rect 748 16549 816 16550
rect 646 16548 816 16549
rect 680 16515 816 16548
rect 680 16514 782 16515
rect 646 16480 714 16514
rect 748 16481 782 16514
rect 748 16480 816 16481
rect 646 16479 816 16480
rect 680 16446 816 16479
rect 680 16445 782 16446
rect 646 16411 714 16445
rect 748 16412 782 16445
rect 748 16411 816 16412
rect 646 16410 816 16411
rect 680 16377 816 16410
rect 3301 16962 3339 16964
rect 3267 16916 3373 16962
rect 3301 16882 3339 16916
rect 3267 16836 3373 16882
rect 3301 16802 3339 16836
rect 3267 16756 3373 16802
rect 3301 16722 3339 16756
rect 3267 16676 3373 16722
rect 3301 16642 3339 16676
rect 3267 16596 3373 16642
rect 3301 16562 3339 16596
rect 3267 16515 3373 16562
rect 3301 16481 3339 16515
rect 3267 16434 3373 16481
rect 3301 16400 3339 16434
rect 5643 16962 5681 16964
rect 5609 16916 5715 16962
rect 5643 16882 5681 16916
rect 5609 16836 5715 16882
rect 5643 16802 5681 16836
rect 5609 16756 5715 16802
rect 5643 16722 5681 16756
rect 5609 16676 5715 16722
rect 5643 16642 5681 16676
rect 5609 16596 5715 16642
rect 5643 16562 5681 16596
rect 5609 16515 5715 16562
rect 5643 16481 5681 16515
rect 5609 16434 5715 16481
rect 5643 16400 5681 16434
rect 7951 16916 8057 16962
rect 7985 16882 8023 16916
rect 7951 16836 8057 16882
rect 7985 16802 8023 16836
rect 7951 16756 8057 16802
rect 7985 16722 8023 16756
rect 7951 16676 8057 16722
rect 7985 16642 8023 16676
rect 7951 16596 8057 16642
rect 7985 16562 8023 16596
rect 7951 16515 8057 16562
rect 7985 16481 8023 16515
rect 7951 16434 8057 16481
rect 7985 16400 8023 16434
rect 10293 16916 10399 16962
rect 10327 16882 10365 16916
rect 10293 16836 10399 16882
rect 10327 16802 10365 16836
rect 10293 16756 10399 16802
rect 10327 16722 10365 16756
rect 10431 16939 10476 16964
rect 10510 16939 10549 16964
rect 10583 16939 10622 16964
rect 10656 16939 10695 16964
rect 10729 16939 10768 16964
rect 10802 16939 10841 16964
rect 10875 16939 10914 16964
rect 10948 16939 10987 16964
rect 11021 16939 11060 16964
rect 11094 16939 11133 16964
rect 10431 16930 11133 16939
rect 15199 16930 15628 16964
rect 10431 16901 10494 16930
rect 10528 16901 10563 16930
rect 10597 16901 10632 16930
rect 10666 16901 10701 16930
rect 10735 16901 10770 16930
rect 10431 16867 10476 16901
rect 10528 16896 10549 16901
rect 10597 16896 10622 16901
rect 10666 16896 10695 16901
rect 10735 16896 10768 16901
rect 10804 16896 10839 16930
rect 10873 16901 10908 16930
rect 10942 16901 10977 16930
rect 11011 16901 11046 16930
rect 11080 16901 11115 16930
rect 10875 16896 10908 16901
rect 10948 16896 10977 16901
rect 11021 16896 11046 16901
rect 11094 16896 11115 16901
rect 10510 16867 10549 16896
rect 10583 16867 10622 16896
rect 10656 16867 10695 16896
rect 10729 16867 10768 16896
rect 10802 16867 10841 16896
rect 10875 16867 10914 16896
rect 10948 16867 10987 16896
rect 11021 16867 11060 16896
rect 11094 16867 11133 16896
rect 10431 16862 14496 16867
rect 10431 16828 10494 16862
rect 10528 16828 10563 16862
rect 10597 16828 10632 16862
rect 10666 16828 10701 16862
rect 10735 16828 10770 16862
rect 10804 16828 10839 16862
rect 10873 16828 10908 16862
rect 10942 16828 10977 16862
rect 11011 16828 11046 16862
rect 11080 16828 11115 16862
rect 11149 16828 11184 16862
rect 11218 16828 11253 16862
rect 11287 16828 11322 16862
rect 11356 16828 11391 16862
rect 11425 16828 11460 16862
rect 11494 16828 11529 16862
rect 11563 16828 11598 16862
rect 11632 16828 11667 16862
rect 11701 16828 11736 16862
rect 11770 16828 11805 16862
rect 11839 16828 11874 16862
rect 11908 16828 11943 16862
rect 11977 16828 12012 16862
rect 12046 16828 12081 16862
rect 12115 16828 12150 16862
rect 12184 16828 12219 16862
rect 12253 16828 12288 16862
rect 12322 16828 12357 16862
rect 12391 16828 12426 16862
rect 12460 16828 12495 16862
rect 12529 16828 12564 16862
rect 12598 16828 12633 16862
rect 12667 16828 12702 16862
rect 12736 16828 12771 16862
rect 12805 16828 12840 16862
rect 12874 16828 12909 16862
rect 12943 16828 12978 16862
rect 13012 16828 13047 16862
rect 13081 16828 13116 16862
rect 13150 16828 13185 16862
rect 13219 16828 13254 16862
rect 13288 16828 13323 16862
rect 13357 16828 13392 16862
rect 13426 16828 13461 16862
rect 13495 16828 13530 16862
rect 13564 16828 13599 16862
rect 13633 16828 13668 16862
rect 13702 16828 13737 16862
rect 13771 16828 13806 16862
rect 13840 16828 13875 16862
rect 13909 16828 13944 16862
rect 13978 16828 14013 16862
rect 14047 16828 14082 16862
rect 14116 16828 14151 16862
rect 14185 16828 14220 16862
rect 14254 16828 14289 16862
rect 14323 16828 14358 16862
rect 14392 16828 14427 16862
rect 14461 16828 14496 16862
rect 10431 16794 14496 16828
rect 10431 16760 10494 16794
rect 10528 16760 10563 16794
rect 10597 16760 10632 16794
rect 10666 16760 10701 16794
rect 10735 16760 10770 16794
rect 10804 16760 10839 16794
rect 10873 16760 10908 16794
rect 10942 16760 10977 16794
rect 11011 16760 11046 16794
rect 11080 16760 11115 16794
rect 11149 16760 11184 16794
rect 11218 16760 11253 16794
rect 11287 16760 11322 16794
rect 11356 16760 11391 16794
rect 11425 16760 11460 16794
rect 11494 16760 11529 16794
rect 11563 16760 11598 16794
rect 11632 16760 11667 16794
rect 11701 16760 11736 16794
rect 11770 16760 11805 16794
rect 11839 16760 11874 16794
rect 11908 16760 11943 16794
rect 11977 16760 12012 16794
rect 12046 16760 12081 16794
rect 12115 16760 12150 16794
rect 12184 16760 12219 16794
rect 12253 16760 12288 16794
rect 12322 16760 12357 16794
rect 12391 16760 12426 16794
rect 12460 16760 12495 16794
rect 12529 16760 12564 16794
rect 12598 16760 12633 16794
rect 12667 16760 12702 16794
rect 12736 16760 12771 16794
rect 12805 16760 12840 16794
rect 12874 16760 12909 16794
rect 12943 16760 12978 16794
rect 13012 16760 13047 16794
rect 13081 16760 13116 16794
rect 13150 16760 13185 16794
rect 13219 16760 13254 16794
rect 13288 16760 13323 16794
rect 13357 16760 13392 16794
rect 13426 16760 13461 16794
rect 13495 16760 13530 16794
rect 13564 16760 13599 16794
rect 13633 16760 13668 16794
rect 13702 16760 13737 16794
rect 13771 16760 13806 16794
rect 13840 16760 13875 16794
rect 13909 16760 13944 16794
rect 13978 16760 14013 16794
rect 14047 16760 14082 16794
rect 14116 16760 14151 16794
rect 14185 16760 14220 16794
rect 14254 16760 14289 16794
rect 14323 16760 14358 16794
rect 14392 16760 14427 16794
rect 14461 16760 14496 16794
rect 15210 16760 15260 16930
rect 15430 16928 15628 16930
rect 15430 16904 15634 16928
rect 15430 16870 15464 16904
rect 15498 16870 15532 16904
rect 15566 16870 15600 16904
rect 15430 16832 15634 16870
rect 15430 16798 15464 16832
rect 15498 16798 15532 16832
rect 15566 16798 15600 16832
rect 10431 16744 15260 16760
rect 10293 16676 10399 16722
rect 10327 16642 10365 16676
rect 10293 16596 10399 16642
rect 10327 16562 10365 16596
rect 10293 16515 10399 16562
rect 10327 16481 10365 16515
rect 10293 16434 10399 16481
rect 10327 16400 10365 16434
rect 15430 16760 15634 16798
rect 15430 16726 15464 16760
rect 15498 16726 15532 16760
rect 15566 16726 15600 16760
rect 15430 16688 15634 16726
rect 15430 16654 15464 16688
rect 15498 16654 15532 16688
rect 15566 16654 15600 16688
rect 15430 16616 15634 16654
rect 15430 16582 15464 16616
rect 15498 16582 15532 16616
rect 15566 16582 15600 16616
rect 15430 16544 15634 16582
rect 15430 16510 15464 16544
rect 15498 16510 15532 16544
rect 15566 16510 15600 16544
rect 15430 16472 15634 16510
rect 15430 16438 15464 16472
rect 15498 16438 15532 16472
rect 15566 16438 15600 16472
rect 680 16376 782 16377
rect 646 16342 714 16376
rect 748 16343 782 16376
rect 748 16342 816 16343
rect 646 16341 816 16342
rect 680 16308 816 16341
rect 680 16307 782 16308
rect 748 16274 782 16307
rect 748 16239 816 16274
rect 12718 16315 15075 16377
rect 12718 16281 14969 16315
rect 15003 16281 15041 16315
rect 12718 16263 15075 16281
rect 15142 16347 15162 16381
rect 15196 16347 15208 16381
rect 15142 16309 15208 16347
rect 15142 16275 15162 16309
rect 15196 16275 15208 16309
rect 12718 16205 14935 16263
rect 15142 16235 15208 16275
rect 10209 15385 10405 16136
rect 12718 15900 12914 16205
rect 15003 16195 15041 16229
rect 12752 15866 12914 15900
rect 12718 15803 12914 15866
rect 12752 15769 12914 15803
rect 12718 15706 12914 15769
rect 12752 15672 12914 15706
rect 12718 15656 12914 15672
rect 15041 15916 15075 16195
rect 15142 16201 15162 16235
rect 15196 16201 15208 16235
rect 15142 16163 15208 16201
rect 15142 16129 15162 16163
rect 15196 16129 15208 16163
rect 15041 15900 15108 15916
rect 15041 15866 15074 15900
rect 15041 15803 15108 15866
rect 15041 15769 15074 15803
rect 15041 15706 15108 15769
rect 15041 15672 15074 15706
rect 15041 15656 15108 15672
rect 14982 15412 15108 15428
rect 10209 14948 10530 15385
rect 14982 15378 15074 15412
rect 14982 15315 15108 15378
rect 14982 15281 15074 15315
rect 12752 15118 12914 15232
rect 14982 15218 15108 15281
rect 14982 15184 15074 15218
rect 14982 15168 15108 15184
rect 12752 14948 14917 15118
rect 3301 14880 3339 14914
rect 3267 14838 3373 14880
rect 3301 14804 3339 14838
rect 3267 14761 3373 14804
rect 3301 14727 3339 14761
rect 3267 14684 3373 14727
rect 7985 14880 8023 14914
rect 7951 14838 8057 14880
rect 7985 14804 8023 14838
rect 7951 14761 8057 14804
rect 7985 14727 8023 14761
rect 3301 14650 3339 14684
rect 3267 14607 3373 14650
rect 3301 14573 3339 14607
rect 3267 14530 3373 14573
rect 3301 14496 3339 14530
rect 3267 14453 3373 14496
rect 3301 14419 3339 14453
rect 3267 14376 3373 14419
rect 3301 14342 3339 14376
rect 3267 14299 3373 14342
rect 3301 14265 3339 14299
rect 3267 14222 3373 14265
rect 3301 14188 3339 14222
rect 3267 14145 3373 14188
rect 3301 14111 3339 14145
rect 3267 14068 3373 14111
rect 3301 14034 3339 14068
rect 3267 13991 3373 14034
rect 3301 13957 3339 13991
rect 3267 13914 3373 13957
rect 3301 13880 3339 13914
rect 5643 14683 5681 14717
rect 5609 14644 5715 14683
rect 5643 14610 5681 14644
rect 5609 14571 5715 14610
rect 5643 14537 5681 14571
rect 5609 14498 5715 14537
rect 5643 14464 5681 14498
rect 5609 14425 5715 14464
rect 5643 14391 5681 14425
rect 5609 14352 5715 14391
rect 5643 14318 5681 14352
rect 5609 14279 5715 14318
rect 5643 14245 5681 14279
rect 5609 14206 5715 14245
rect 5643 14172 5681 14206
rect 5609 14133 5715 14172
rect 5643 14099 5681 14133
rect 5609 14060 5715 14099
rect 5643 14026 5681 14060
rect 5609 13987 5715 14026
rect 5643 13953 5681 13987
rect 5609 13914 5715 13953
rect 5643 13880 5681 13914
rect 7951 14684 8057 14727
rect 12716 14880 12754 14914
rect 12682 14838 12788 14880
rect 12716 14804 12754 14838
rect 12682 14761 12788 14804
rect 12716 14727 12754 14761
rect 7985 14650 8023 14684
rect 7951 14607 8057 14650
rect 7985 14573 8023 14607
rect 7951 14530 8057 14573
rect 7985 14496 8023 14530
rect 7951 14453 8057 14496
rect 7985 14419 8023 14453
rect 7951 14376 8057 14419
rect 7985 14342 8023 14376
rect 7951 14299 8057 14342
rect 7985 14265 8023 14299
rect 7951 14222 8057 14265
rect 7985 14188 8023 14222
rect 7951 14145 8057 14188
rect 7985 14111 8023 14145
rect 7951 14068 8057 14111
rect 7985 14034 8023 14068
rect 7951 13991 8057 14034
rect 7985 13957 8023 13991
rect 7951 13914 8057 13957
rect 7985 13880 8023 13914
rect 10327 14683 10365 14717
rect 10293 14644 10399 14683
rect 10327 14610 10365 14644
rect 10293 14571 10399 14610
rect 10327 14537 10365 14571
rect 10293 14498 10399 14537
rect 10327 14464 10365 14498
rect 10293 14425 10399 14464
rect 10327 14391 10365 14425
rect 10293 14352 10399 14391
rect 10327 14318 10365 14352
rect 10293 14279 10399 14318
rect 10327 14245 10365 14279
rect 10293 14206 10399 14245
rect 10327 14172 10365 14206
rect 10293 14133 10399 14172
rect 10327 14099 10365 14133
rect 10293 14060 10399 14099
rect 10327 14026 10365 14060
rect 10293 13987 10399 14026
rect 10327 13953 10365 13987
rect 10293 13914 10399 13953
rect 10327 13880 10365 13914
rect 12682 14684 12788 14727
rect 12854 14833 14917 14948
rect 14982 14976 15088 15168
rect 14982 14942 14986 14976
rect 15020 14942 15088 14976
rect 14982 14904 15088 14942
rect 14982 14870 14986 14904
rect 15020 14870 15088 14904
rect 15142 14910 15208 16129
rect 15142 14876 15159 14910
rect 15193 14876 15208 14910
rect 15142 14838 15208 14876
rect 12854 14707 15088 14833
rect 12716 14650 12754 14684
rect 12682 14607 12788 14650
rect 12716 14573 12754 14607
rect 12682 14530 12788 14573
rect 12716 14496 12754 14530
rect 12682 14453 12788 14496
rect 12716 14419 12754 14453
rect 12682 14376 12788 14419
rect 12716 14342 12754 14376
rect 12682 14299 12788 14342
rect 12716 14265 12754 14299
rect 12682 14222 12788 14265
rect 12716 14188 12754 14222
rect 12682 14145 12788 14188
rect 14982 14643 15088 14707
rect 14982 14609 14986 14643
rect 15020 14609 15088 14643
rect 14982 14571 15088 14609
rect 14982 14537 14986 14571
rect 15020 14537 15088 14571
rect 14982 14172 15088 14537
rect 12716 14111 12754 14145
rect 12682 14068 12788 14111
rect 12716 14034 12754 14068
rect 12682 13991 12788 14034
rect 12716 13957 12754 13991
rect 12682 13914 12788 13957
rect 12716 13880 12754 13914
rect 12854 14002 15088 14172
rect 15142 14804 15159 14838
rect 15193 14804 15208 14838
rect 15142 14637 15208 14804
rect 15142 14603 15159 14637
rect 15193 14603 15208 14637
rect 15142 14565 15208 14603
rect 15142 14531 15159 14565
rect 15193 14531 15208 14565
rect 12854 13846 13024 14002
rect 10346 13562 10376 13846
rect 12718 13782 13024 13846
rect 14982 13830 15108 13846
rect 14982 13796 15074 13830
rect 12718 13366 12914 13782
rect 14982 13733 15108 13796
rect 14982 13699 15074 13733
rect 14982 13636 15108 13699
rect 14982 13602 15074 13636
rect 14982 13586 15108 13602
rect 12983 13138 14929 13154
rect 14982 13138 15075 13586
rect 15142 13154 15208 14531
rect 15430 16400 15634 16438
rect 15430 16366 15464 16400
rect 15498 16366 15532 16400
rect 15566 16366 15600 16400
rect 15430 16328 15634 16366
rect 15430 16294 15464 16328
rect 15498 16294 15532 16328
rect 15566 16294 15600 16328
rect 15430 16255 15634 16294
rect 15430 16221 15464 16255
rect 15498 16221 15532 16255
rect 15566 16221 15600 16255
rect 15430 16197 15634 16221
rect 17916 16598 18020 16624
rect 17916 16593 18052 16598
rect 17916 16589 17948 16593
rect 17982 16590 18052 16593
rect 17982 16589 18086 16590
rect 17982 16559 17984 16589
rect 17950 16555 17984 16559
rect 18018 16559 18086 16589
rect 18018 16555 18020 16559
rect 18054 16556 18086 16559
rect 17916 16525 18020 16555
rect 17916 16522 18052 16525
rect 17916 16520 18086 16522
rect 17982 16486 17984 16520
rect 18018 16488 18086 16520
rect 18018 16486 18052 16488
rect 17916 16452 18020 16486
rect 18054 16452 18086 16454
rect 17916 16451 18086 16452
rect 17950 16447 17984 16451
rect 17982 16417 17984 16447
rect 18018 16420 18086 16451
rect 18018 16417 18052 16420
rect 17916 16413 17948 16417
rect 17982 16413 18052 16417
rect 17916 16382 18020 16413
rect 17950 16374 17984 16382
rect 17982 16348 17984 16374
rect 18018 16379 18020 16382
rect 18054 16379 18086 16386
rect 18018 16352 18086 16379
rect 18018 16348 18052 16352
rect 17916 16340 17948 16348
rect 17982 16340 18052 16348
rect 17916 16313 18020 16340
rect 17950 16301 17984 16313
rect 17982 16279 17984 16301
rect 18018 16306 18020 16313
rect 18054 16306 18086 16318
rect 18018 16284 18086 16306
rect 18018 16279 18052 16284
rect 17916 16267 17948 16279
rect 17982 16267 18052 16279
rect 17916 16244 18020 16267
rect 17950 16228 17984 16244
rect 17982 16210 17984 16228
rect 18018 16233 18020 16244
rect 18054 16233 18086 16250
rect 18018 16216 18086 16233
rect 18018 16210 18052 16216
rect 17916 16194 17948 16210
rect 17982 16194 18052 16210
rect 17916 16175 18020 16194
rect 17950 16155 17984 16175
rect 17982 16141 17984 16155
rect 18018 16160 18020 16175
rect 18054 16160 18086 16182
rect 18018 16148 18086 16160
rect 18018 16141 18052 16148
rect 17916 16121 17948 16141
rect 17982 16121 18052 16141
rect 17916 16106 18020 16121
rect 17950 16082 17984 16106
rect 15260 14771 15396 14788
rect 15260 14753 15430 14771
rect 15294 14719 15328 14753
rect 15362 14719 15396 14753
rect 15260 14698 15396 14719
rect 15260 14684 15430 14698
rect 15294 14650 15328 14684
rect 15362 14650 15396 14684
rect 15260 14624 15396 14650
rect 15260 14615 15430 14624
rect 15294 14581 15328 14615
rect 15362 14581 15396 14615
rect 15260 14550 15396 14581
rect 15260 14546 15430 14550
rect 15294 14512 15328 14546
rect 15362 14512 15396 14546
rect 15260 14510 15430 14512
rect 15260 14477 15396 14510
rect 15294 14443 15328 14477
rect 15362 14443 15396 14477
rect 15260 14436 15430 14443
rect 15260 14408 15396 14436
rect 15294 14374 15328 14408
rect 15362 14374 15396 14408
rect 15260 14362 15430 14374
rect 15260 14350 15396 14362
rect 15242 13188 15348 14299
rect 15396 14288 15430 14306
rect 15396 14214 15430 14235
rect 15396 14140 15430 14164
rect 15396 14066 15430 14093
rect 15396 13992 15430 14022
rect 15396 13918 15430 13951
rect 15396 13844 15430 13880
rect 15396 13772 15430 13809
rect 15396 13701 15430 13736
rect 15396 13630 15430 13662
rect 15396 13559 15430 13588
rect 15396 13488 15430 13514
rect 15396 13417 15430 13440
rect 15396 13346 15430 13366
rect 15396 13275 15430 13292
rect 15396 13217 15430 13218
rect 15479 16065 15672 16081
rect 15479 16031 15638 16065
rect 15479 15968 15672 16031
rect 15479 15934 15638 15968
rect 15479 15871 15672 15934
rect 15479 15837 15638 15871
rect 15479 15821 15672 15837
rect 17982 16072 17984 16082
rect 18018 16087 18020 16106
rect 18054 16087 18086 16114
rect 18018 16080 18086 16087
rect 18018 16072 18052 16080
rect 17916 16048 17948 16072
rect 17982 16048 18052 16072
rect 17916 16037 18020 16048
rect 17950 16009 17984 16037
rect 17982 16003 17984 16009
rect 18018 16014 18020 16037
rect 18054 16014 18086 16046
rect 18018 16012 18086 16014
rect 18018 16003 18052 16012
rect 17916 15975 17948 16003
rect 17982 15978 18052 16003
rect 17982 15975 18086 15978
rect 17916 15968 18020 15975
rect 17950 15936 17984 15968
rect 17982 15934 17984 15936
rect 18018 15941 18020 15968
rect 18054 15944 18086 15975
rect 18018 15934 18052 15941
rect 17916 15902 17948 15934
rect 17982 15910 18052 15934
rect 17982 15902 18086 15910
rect 17916 15899 18020 15902
rect 17950 15865 17984 15899
rect 18018 15868 18020 15899
rect 18054 15876 18086 15902
rect 18018 15865 18052 15868
rect 17916 15863 18052 15865
rect 17916 15830 17948 15863
rect 17982 15842 18052 15863
rect 17982 15830 18086 15842
rect 17982 15829 17984 15830
rect 12983 13104 12985 13138
rect 13019 13104 14823 13138
rect 14857 13104 14895 13138
rect 15003 13104 15041 13138
rect 15123 13138 15229 13154
rect 15157 13104 15195 13138
rect 12983 13088 14929 13104
rect 15123 13088 15229 13104
rect 15263 13043 15348 13188
rect 15479 13183 15585 15821
rect 17950 15796 17984 15829
rect 18018 15829 18086 15830
rect 18018 15796 18020 15829
rect 18054 15808 18086 15829
rect 17916 15795 18020 15796
rect 17916 15790 18052 15795
rect 17916 15761 17948 15790
rect 17982 15774 18052 15790
rect 17982 15761 18086 15774
rect 17982 15756 17984 15761
rect 17950 15727 17984 15756
rect 18018 15756 18086 15761
rect 18018 15727 18020 15756
rect 18054 15740 18086 15756
rect 17916 15722 18020 15727
rect 17916 15717 18052 15722
rect 17916 15692 17948 15717
rect 17982 15706 18052 15717
rect 17982 15692 18086 15706
rect 17982 15683 17984 15692
rect 17950 15658 17984 15683
rect 18018 15683 18086 15692
rect 18018 15658 18020 15683
rect 18054 15672 18086 15683
rect 17916 15649 18020 15658
rect 17916 15644 18052 15649
rect 17916 15623 17948 15644
rect 17982 15638 18052 15644
rect 17982 15623 18086 15638
rect 17982 15610 17984 15623
rect 17950 15589 17984 15610
rect 18018 15610 18086 15623
rect 18018 15589 18020 15610
rect 18054 15604 18086 15610
rect 17916 15576 18020 15589
rect 17916 15571 18052 15576
rect 17916 15554 17948 15571
rect 17982 15570 18052 15571
rect 17982 15554 18086 15570
rect 17982 15537 17984 15554
rect 17950 15520 17984 15537
rect 18018 15537 18086 15554
rect 18018 15520 18020 15537
rect 18054 15536 18086 15537
rect 17916 15503 18020 15520
rect 17916 15502 18052 15503
rect 17916 15498 18086 15502
rect 17916 15485 17948 15498
rect 17982 15485 18086 15498
rect 17982 15464 17984 15485
rect 17950 15451 17984 15464
rect 18018 15468 18086 15485
rect 18018 15464 18052 15468
rect 18018 15451 18020 15464
rect 17916 15430 18020 15451
rect 18054 15430 18086 15434
rect 17916 15425 18086 15430
rect 17916 15416 17948 15425
rect 17982 15416 18086 15425
rect 17982 15391 17984 15416
rect 17950 15382 17984 15391
rect 18018 15400 18086 15416
rect 18018 15391 18052 15400
rect 18018 15382 18020 15391
rect 17916 15357 18020 15382
rect 18054 15357 18086 15366
rect 17916 15352 18086 15357
rect 17916 15347 17948 15352
rect 17982 15347 18086 15352
rect 17982 15318 17984 15347
rect 17950 15313 17984 15318
rect 18018 15332 18086 15347
rect 18018 15318 18052 15332
rect 18018 15313 18020 15318
rect 17916 15284 18020 15313
rect 18054 15284 18086 15298
rect 17916 15279 18086 15284
rect 17916 15278 17948 15279
rect 17982 15278 18086 15279
rect 17982 15245 17984 15278
rect 17950 15244 17984 15245
rect 18018 15264 18086 15278
rect 18018 15245 18052 15264
rect 18018 15244 18020 15245
rect 17916 15211 18020 15244
rect 18054 15211 18086 15230
rect 17916 15209 18086 15211
rect 17950 15206 17984 15209
rect 17982 15175 17984 15206
rect 18018 15196 18086 15209
rect 18018 15175 18052 15196
rect 17916 15172 17948 15175
rect 17982 15172 18052 15175
rect 17916 15140 18020 15172
rect 17950 15133 17984 15140
rect 17982 15106 17984 15133
rect 18018 15138 18020 15140
rect 18054 15138 18086 15162
rect 18018 15128 18086 15138
rect 18018 15106 18052 15128
rect 17916 15099 17948 15106
rect 17982 15099 18052 15106
rect 17916 15071 18020 15099
rect 17950 15060 17984 15071
rect 17982 15037 17984 15060
rect 18018 15065 18020 15071
rect 18054 15065 18086 15094
rect 18018 15060 18086 15065
rect 18018 15037 18052 15060
rect 17916 15026 17948 15037
rect 17982 15026 18052 15037
rect 17916 15002 18020 15026
rect 17950 14987 17984 15002
rect 15275 13009 15313 13043
rect 15347 13009 15348 13043
rect 15387 13077 15585 13183
rect 15619 14969 15692 14985
rect 15619 14935 15638 14969
rect 15672 14935 15692 14969
rect 15619 14872 15692 14935
rect 15619 14838 15638 14872
rect 15672 14838 15692 14872
rect 15619 14775 15692 14838
rect 15619 14741 15638 14775
rect 15672 14741 15692 14775
rect 15619 13607 15692 14741
rect 15619 13573 15638 13607
rect 15672 13573 15692 13607
rect 15619 13510 15692 13573
rect 15619 13476 15638 13510
rect 15672 13476 15692 13510
rect 15619 13413 15692 13476
rect 15619 13379 15638 13413
rect 15672 13379 15692 13413
rect 15387 13043 15499 13077
rect 15619 13043 15692 13379
rect 15421 13009 15459 13043
rect 15493 13009 15499 13043
rect 15567 13009 15605 13043
rect 15639 13009 15692 13043
rect 17982 14968 17984 14987
rect 18018 14992 18020 15002
rect 18054 14992 18086 15026
rect 18018 14968 18052 14992
rect 17916 14953 17948 14968
rect 17982 14958 18052 14968
rect 17982 14953 18086 14958
rect 17916 14933 18020 14953
rect 17950 14914 17984 14933
rect 17982 14899 17984 14914
rect 18018 14919 18020 14933
rect 18054 14924 18086 14953
rect 18018 14899 18052 14919
rect 17916 14880 17948 14899
rect 17982 14890 18052 14899
rect 17982 14880 18086 14890
rect 17916 14864 18020 14880
rect 17950 14841 17984 14864
rect 17982 14830 17984 14841
rect 18018 14846 18020 14864
rect 18054 14856 18086 14880
rect 18018 14830 18052 14846
rect 17916 14807 17948 14830
rect 17982 14822 18052 14830
rect 17982 14807 18086 14822
rect 17916 14795 18020 14807
rect 17950 14768 17984 14795
rect 17982 14761 17984 14768
rect 18018 14773 18020 14795
rect 18054 14788 18086 14807
rect 18018 14761 18052 14773
rect 17916 14734 17948 14761
rect 17982 14754 18052 14761
rect 17982 14734 18086 14754
rect 17916 14726 18020 14734
rect 17950 14695 17984 14726
rect 17982 14692 17984 14695
rect 18018 14700 18020 14726
rect 18054 14720 18086 14734
rect 18018 14692 18052 14700
rect 17916 14661 17948 14692
rect 17982 14686 18052 14692
rect 17982 14661 18086 14686
rect 17916 14657 18020 14661
rect 17950 14623 17984 14657
rect 18018 14627 18020 14657
rect 18054 14652 18086 14661
rect 18018 14623 18052 14627
rect 17916 14622 18052 14623
rect 17916 14588 17948 14622
rect 17982 14618 18052 14622
rect 17982 14588 18086 14618
rect 17950 14554 17984 14588
rect 18018 14554 18020 14588
rect 18054 14584 18086 14588
rect 17916 14550 18052 14554
rect 17916 14549 18086 14550
rect 17916 14519 17948 14549
rect 17982 14519 18086 14549
rect 17982 14515 17984 14519
rect 17950 14485 17984 14515
rect 18018 14516 18086 14519
rect 18018 14515 18052 14516
rect 18018 14485 18020 14515
rect 17916 14481 18020 14485
rect 18054 14481 18086 14482
rect 17916 14476 18086 14481
rect 17916 14450 17948 14476
rect 17982 14450 18086 14476
rect 17982 14442 17984 14450
rect 17950 14416 17984 14442
rect 18018 14448 18086 14450
rect 18018 14442 18052 14448
rect 18018 14416 18020 14442
rect 17916 14408 18020 14416
rect 18054 14408 18086 14414
rect 17916 14403 18086 14408
rect 17916 14381 17948 14403
rect 17982 14381 18086 14403
rect 17982 14369 17984 14381
rect 17950 14347 17984 14369
rect 18018 14380 18086 14381
rect 18018 14369 18052 14380
rect 18018 14347 18020 14369
rect 17916 14335 18020 14347
rect 18054 14335 18086 14346
rect 17916 14330 18086 14335
rect 17916 14312 17948 14330
rect 17982 14312 18086 14330
rect 17982 14296 17984 14312
rect 17950 14278 17984 14296
rect 18018 14296 18052 14312
rect 18018 14278 18020 14296
rect 17916 14262 18020 14278
rect 18054 14262 18086 14278
rect 17916 14257 18086 14262
rect 17916 14243 17948 14257
rect 17982 14243 18086 14257
rect 17982 14223 17984 14243
rect 17950 14209 17984 14223
rect 18018 14223 18052 14243
rect 18018 14209 18020 14223
rect 17916 14189 18020 14209
rect 18054 14189 18086 14209
rect 17916 14184 18086 14189
rect 17916 14174 17948 14184
rect 17982 14174 18086 14184
rect 17982 14150 17984 14174
rect 17950 14140 17984 14150
rect 18018 14150 18052 14174
rect 18018 14140 18020 14150
rect 17916 14116 18020 14140
rect 18054 14116 18086 14140
rect 17916 14111 18086 14116
rect 17916 14105 17948 14111
rect 17982 14105 18086 14111
rect 17982 14077 17984 14105
rect 17950 14071 17984 14077
rect 18018 14077 18052 14105
rect 18018 14071 18020 14077
rect 17916 14043 18020 14071
rect 18054 14043 18086 14071
rect 17916 14038 18086 14043
rect 17916 14036 17948 14038
rect 17982 14036 18086 14038
rect 17982 14004 17984 14036
rect 17950 14002 17984 14004
rect 18018 14004 18052 14036
rect 18018 14002 18020 14004
rect 17916 13970 18020 14002
rect 18054 13970 18086 14002
rect 17916 13967 18086 13970
rect 17950 13965 17984 13967
rect 17982 13933 17984 13965
rect 18018 13933 18052 13967
rect 17916 13931 17948 13933
rect 17982 13931 18086 13933
rect 17916 13898 18020 13931
rect 18054 13898 18086 13931
rect 17950 13892 17984 13898
rect 17982 13864 17984 13892
rect 18018 13897 18020 13898
rect 18018 13864 18052 13897
rect 17916 13858 17948 13864
rect 17982 13858 18086 13864
rect 17916 13829 18020 13858
rect 18054 13829 18086 13858
rect 17950 13819 17984 13829
rect 17982 13795 17984 13819
rect 18018 13824 18020 13829
rect 18018 13795 18052 13824
rect 17916 13785 17948 13795
rect 17982 13785 18086 13795
rect 17916 13760 18020 13785
rect 18054 13760 18086 13785
rect 17950 13746 17984 13760
rect 17982 13726 17984 13746
rect 18018 13751 18020 13760
rect 18018 13726 18052 13751
rect 17916 13712 17948 13726
rect 17982 13712 18086 13726
rect 17916 13691 18020 13712
rect 18054 13691 18086 13712
rect 17950 13673 17984 13691
rect 17982 13657 17984 13673
rect 18018 13678 18020 13691
rect 18018 13657 18052 13678
rect 17916 13639 17948 13657
rect 17982 13639 18086 13657
rect 17916 13622 18020 13639
rect 18054 13622 18086 13639
rect 17950 13600 17984 13622
rect 17982 13588 17984 13600
rect 18018 13605 18020 13622
rect 18018 13588 18052 13605
rect 17916 13566 17948 13588
rect 17982 13566 18086 13588
rect 17916 13553 18020 13566
rect 18054 13553 18086 13566
rect 17950 13527 17984 13553
rect 17982 13519 17984 13527
rect 18018 13532 18020 13553
rect 18018 13519 18052 13532
rect 17916 13493 17948 13519
rect 17982 13493 18086 13519
rect 17916 13484 18020 13493
rect 18054 13484 18086 13493
rect 17950 13454 17984 13484
rect 17982 13450 17984 13454
rect 18018 13459 18020 13484
rect 18018 13450 18052 13459
rect 17916 13420 17948 13450
rect 17982 13420 18086 13450
rect 17916 13415 18020 13420
rect 18054 13415 18086 13420
rect 17950 13381 17984 13415
rect 18018 13386 18020 13415
rect 18018 13381 18052 13386
rect 17916 13347 17948 13381
rect 17982 13347 18086 13381
rect 17916 13346 18020 13347
rect 18054 13346 18086 13347
rect 17950 13312 17984 13346
rect 18018 13313 18020 13346
rect 18018 13312 18052 13313
rect 17916 13308 18086 13312
rect 17916 13277 17948 13308
rect 17982 13277 18086 13308
rect 17982 13274 17984 13277
rect 17950 13243 17984 13274
rect 18018 13274 18052 13277
rect 18018 13243 18020 13274
rect 17916 13240 18020 13243
rect 18054 13240 18086 13243
rect 17916 13235 18086 13240
rect 17916 13208 17948 13235
rect 17982 13208 18086 13235
rect 17982 13201 17984 13208
rect 17950 13174 17984 13201
rect 18018 13201 18052 13208
rect 18018 13174 18020 13201
rect 17916 13167 18020 13174
rect 18054 13167 18086 13174
rect 17916 13162 18086 13167
rect 17916 13139 17948 13162
rect 17982 13139 18086 13162
rect 17982 13128 17984 13139
rect 17950 13105 17984 13128
rect 18018 13128 18052 13139
rect 18018 13105 18020 13128
rect 17916 13094 18020 13105
rect 18054 13094 18086 13105
rect 17916 13089 18086 13094
rect 17916 13070 17948 13089
rect 17982 13070 18086 13089
rect 17982 13055 17984 13070
rect 17950 13036 17984 13055
rect 18018 13055 18052 13070
rect 18018 13036 18020 13055
rect 17916 13021 18020 13036
rect 18054 13021 18086 13036
rect 17916 13016 18086 13021
rect 17916 13001 17948 13016
rect 17982 13001 18086 13016
rect 17982 12982 17984 13001
rect 816 12943 851 12975
rect 885 12943 920 12975
rect 954 12943 989 12975
rect 1023 12943 1058 12975
rect 1092 12943 1127 12975
rect 1161 12943 1196 12975
rect 1230 12943 1265 12975
rect 1299 12943 1334 12975
rect 1368 12943 1403 12975
rect 1437 12943 1472 12975
rect 1506 12943 1541 12975
rect 1575 12943 1610 12975
rect 1644 12943 1679 12975
rect 1713 12943 1748 12975
rect 1782 12943 1817 12975
rect 1851 12943 1886 12975
rect 1920 12943 1955 12975
rect 1989 12943 2024 12975
rect 2058 12943 2093 12975
rect 2127 12943 2162 12975
rect 2196 12943 2231 12975
rect 2265 12943 2300 12975
rect 2334 12943 2369 12975
rect 2403 12943 2438 12975
rect 17840 12967 17916 12975
rect 17950 12967 17984 12982
rect 18018 12982 18052 13001
rect 18018 12967 18020 12982
rect 17840 12948 18020 12967
rect 18054 12948 18086 12967
rect 17840 12943 18086 12948
rect 816 12941 829 12943
rect 748 12921 752 12941
rect 786 12921 829 12941
rect 748 12907 829 12921
rect 646 12881 714 12907
rect 646 12847 680 12881
rect 748 12881 783 12907
rect 748 12873 752 12881
rect 817 12873 829 12907
rect 17840 12909 17875 12943
rect 17909 12932 17948 12943
rect 17982 12932 18086 12943
rect 17909 12909 17916 12932
rect 17982 12909 17984 12932
rect 714 12847 752 12873
rect 786 12847 829 12873
rect 646 12839 829 12847
rect 646 12805 680 12839
rect 714 12805 749 12839
rect 783 12805 818 12839
rect 17840 12898 17916 12909
rect 17950 12898 17984 12909
rect 18018 12909 18052 12932
rect 18018 12898 18020 12909
rect 17840 12875 18020 12898
rect 18054 12875 18086 12898
rect 17840 12871 18086 12875
rect 17866 12837 17906 12871
rect 17940 12863 18086 12871
rect 852 12805 887 12837
rect 921 12805 956 12837
rect 990 12805 1025 12837
rect 1059 12805 1094 12837
rect 1128 12805 1163 12837
rect 1197 12805 1232 12837
rect 1266 12805 1301 12837
rect 1335 12805 1370 12837
rect 1404 12805 1439 12837
rect 1473 12805 1508 12837
rect 1542 12805 1577 12837
rect 1611 12805 1646 12837
rect 1680 12805 1715 12837
rect 1749 12805 1784 12837
rect 1818 12805 1853 12837
rect 1887 12805 1922 12837
rect 1956 12805 1991 12837
rect 2025 12805 2060 12837
rect 2094 12805 2129 12837
rect 2163 12805 2198 12837
rect 2232 12805 2267 12837
rect 2301 12805 2336 12837
rect 2370 12805 2405 12837
rect 2439 12805 2474 12837
rect 2508 12805 2543 12837
rect 2577 12805 2612 12837
rect 2646 12805 2681 12837
rect 2715 12805 2750 12837
rect 2784 12805 2819 12837
rect 2853 12805 2888 12837
rect 2922 12805 2957 12837
rect 2991 12805 3026 12837
rect 3060 12805 3095 12837
rect 3129 12805 3164 12837
rect 3198 12805 3233 12837
rect 3267 12805 3302 12837
rect 3336 12805 3371 12837
rect 3405 12805 3440 12837
rect 3474 12805 3509 12837
rect 3543 12805 3578 12837
rect 3612 12805 3647 12837
rect 3681 12805 3716 12837
rect 3750 12805 3785 12837
rect 3819 12805 3854 12837
rect 3888 12805 3923 12837
rect 3957 12805 3992 12837
rect 4026 12805 4061 12837
rect 4095 12805 4130 12837
rect 4164 12805 4199 12837
rect 4233 12805 4268 12837
rect 4302 12805 4337 12837
rect 4371 12805 4406 12837
rect 4440 12805 4475 12837
rect 4509 12805 4544 12837
rect 4578 12805 4613 12837
rect 4647 12805 4682 12837
rect 17840 12829 17916 12837
rect 17950 12829 17984 12863
rect 18018 12829 18052 12863
rect 17840 12805 18086 12829
rect 18239 15688 18307 15723
rect 18273 15686 18307 15688
rect 18305 15655 18307 15686
rect 18239 15652 18271 15654
rect 18305 15652 18375 15655
rect 18239 15620 18343 15652
rect 18239 15619 18307 15620
rect 18273 15613 18307 15619
rect 18305 15586 18307 15613
rect 18341 15618 18343 15620
rect 18377 15618 18409 15621
rect 18341 15586 18409 15618
rect 18239 15579 18271 15585
rect 18305 15579 18375 15586
rect 18239 15551 18343 15579
rect 18239 15550 18307 15551
rect 18273 15540 18307 15550
rect 18305 15517 18307 15540
rect 18341 15545 18343 15551
rect 18377 15545 18409 15552
rect 18341 15517 18409 15545
rect 18239 15506 18271 15516
rect 18305 15506 18375 15517
rect 18239 15482 18343 15506
rect 18239 15481 18307 15482
rect 18273 15467 18307 15481
rect 18305 15448 18307 15467
rect 18341 15472 18343 15482
rect 18377 15472 18409 15483
rect 18341 15448 18409 15472
rect 18239 15433 18271 15447
rect 18305 15433 18375 15448
rect 18239 15413 18343 15433
rect 18239 15412 18307 15413
rect 18273 15394 18307 15412
rect 18305 15379 18307 15394
rect 18341 15399 18343 15413
rect 18377 15399 18409 15414
rect 18341 15379 18409 15399
rect 18239 15360 18271 15378
rect 18305 15360 18375 15379
rect 18239 15344 18343 15360
rect 18239 15343 18307 15344
rect 18273 15321 18307 15343
rect 18305 15310 18307 15321
rect 18341 15326 18343 15344
rect 18377 15326 18409 15345
rect 18341 15310 18409 15326
rect 18239 15287 18271 15309
rect 18305 15287 18375 15310
rect 18239 15275 18343 15287
rect 18239 15274 18307 15275
rect 18273 15248 18307 15274
rect 18305 15241 18307 15248
rect 18341 15253 18343 15275
rect 18377 15253 18409 15276
rect 18341 15241 18409 15253
rect 18239 15214 18271 15240
rect 18305 15214 18375 15241
rect 18239 15206 18343 15214
rect 18239 15205 18307 15206
rect 18273 15175 18307 15205
rect 18305 15172 18307 15175
rect 18341 15180 18343 15206
rect 18377 15180 18409 15207
rect 18341 15172 18409 15180
rect 18239 15141 18271 15171
rect 18305 15141 18375 15172
rect 18239 15137 18343 15141
rect 18239 15136 18307 15137
rect 18273 15103 18307 15136
rect 18341 15107 18343 15137
rect 18377 15107 18409 15138
rect 18341 15103 18409 15107
rect 18273 15102 18375 15103
rect 18239 15068 18271 15102
rect 18305 15069 18375 15102
rect 18305 15068 18409 15069
rect 18239 15067 18307 15068
rect 18273 15034 18307 15067
rect 18341 15034 18343 15068
rect 18377 15034 18409 15068
rect 18273 15033 18375 15034
rect 18239 15029 18375 15033
rect 18239 14998 18271 15029
rect 18305 15000 18375 15029
rect 18305 14999 18409 15000
rect 18305 14995 18307 14999
rect 18273 14965 18307 14995
rect 18341 14995 18409 14999
rect 18341 14965 18343 14995
rect 18377 14965 18409 14995
rect 18273 14964 18343 14965
rect 18239 14961 18343 14964
rect 18239 14956 18375 14961
rect 18239 14929 18271 14956
rect 18305 14931 18375 14956
rect 18305 14930 18409 14931
rect 18305 14922 18307 14930
rect 18273 14896 18307 14922
rect 18341 14922 18409 14930
rect 18341 14896 18343 14922
rect 18377 14896 18409 14922
rect 18273 14895 18343 14896
rect 18239 14888 18343 14895
rect 18239 14883 18375 14888
rect 18239 14860 18271 14883
rect 18305 14862 18375 14883
rect 18305 14861 18409 14862
rect 18305 14849 18307 14861
rect 18273 14827 18307 14849
rect 18341 14849 18409 14861
rect 18341 14827 18343 14849
rect 18377 14827 18409 14849
rect 18273 14826 18343 14827
rect 18239 14815 18343 14826
rect 18239 14810 18375 14815
rect 18239 14791 18271 14810
rect 18305 14793 18375 14810
rect 18305 14792 18409 14793
rect 18305 14776 18307 14792
rect 18273 14758 18307 14776
rect 18341 14776 18409 14792
rect 18341 14758 18343 14776
rect 18377 14758 18409 14776
rect 18273 14757 18343 14758
rect 18239 14742 18343 14757
rect 18239 14737 18375 14742
rect 18239 14722 18271 14737
rect 18305 14724 18375 14737
rect 18305 14723 18409 14724
rect 18305 14703 18307 14723
rect 18273 14689 18307 14703
rect 18341 14703 18409 14723
rect 18341 14689 18343 14703
rect 18377 14689 18409 14703
rect 18273 14688 18343 14689
rect 18239 14669 18343 14688
rect 18239 14664 18375 14669
rect 18239 14653 18271 14664
rect 18305 14655 18375 14664
rect 18305 14654 18409 14655
rect 18305 14630 18307 14654
rect 18273 14620 18307 14630
rect 18341 14630 18409 14654
rect 18341 14620 18343 14630
rect 18377 14620 18409 14630
rect 18273 14619 18343 14620
rect 18239 14596 18343 14619
rect 18239 14591 18375 14596
rect 18239 14584 18271 14591
rect 18305 14586 18375 14591
rect 18305 14585 18409 14586
rect 18305 14557 18307 14585
rect 18273 14551 18307 14557
rect 18341 14557 18409 14585
rect 18341 14551 18343 14557
rect 18377 14551 18409 14557
rect 18273 14550 18343 14551
rect 18239 14523 18343 14550
rect 18239 14518 18375 14523
rect 18239 14515 18271 14518
rect 18305 14517 18375 14518
rect 18305 14516 18409 14517
rect 18305 14484 18307 14516
rect 18273 14482 18307 14484
rect 18341 14484 18409 14516
rect 18341 14482 18343 14484
rect 18377 14482 18409 14484
rect 18273 14481 18343 14482
rect 18239 14450 18343 14481
rect 18239 14448 18375 14450
rect 18239 14447 18409 14448
rect 18239 14446 18307 14447
rect 18273 14445 18307 14446
rect 18305 14413 18307 14445
rect 18341 14413 18409 14447
rect 18239 14411 18271 14412
rect 18305 14411 18375 14413
rect 18239 14378 18343 14411
rect 18239 14377 18307 14378
rect 18273 14372 18307 14377
rect 18305 14344 18307 14372
rect 18341 14377 18343 14378
rect 18377 14377 18409 14379
rect 18341 14344 18409 14377
rect 18239 14338 18271 14343
rect 18305 14338 18375 14344
rect 18239 14309 18343 14338
rect 18239 14308 18307 14309
rect 18273 14299 18307 14308
rect 18305 14275 18307 14299
rect 18341 14304 18343 14309
rect 18377 14304 18409 14310
rect 18341 14275 18409 14304
rect 18239 14265 18271 14274
rect 18305 14265 18375 14275
rect 18239 14240 18343 14265
rect 18239 14239 18307 14240
rect 18273 14226 18307 14239
rect 18305 14206 18307 14226
rect 18341 14231 18343 14240
rect 18377 14231 18409 14241
rect 18341 14206 18409 14231
rect 18239 14192 18271 14205
rect 18305 14192 18375 14206
rect 18239 14171 18343 14192
rect 18239 14170 18307 14171
rect 18273 14153 18307 14170
rect 18305 14137 18307 14153
rect 18341 14158 18343 14171
rect 18377 14158 18409 14172
rect 18341 14137 18409 14158
rect 18239 14119 18271 14136
rect 18305 14119 18375 14137
rect 18239 14102 18343 14119
rect 18239 14101 18307 14102
rect 18273 14080 18307 14101
rect 18305 14068 18307 14080
rect 18341 14085 18343 14102
rect 18377 14085 18409 14103
rect 18341 14068 18409 14085
rect 18239 14046 18271 14067
rect 18305 14046 18375 14068
rect 18239 14033 18343 14046
rect 18239 14032 18307 14033
rect 18273 14007 18307 14032
rect 18305 13999 18307 14007
rect 18341 14012 18343 14033
rect 18377 14012 18409 14034
rect 18341 13999 18409 14012
rect 18239 13973 18271 13998
rect 18305 13973 18375 13999
rect 18239 13964 18343 13973
rect 18239 13963 18307 13964
rect 18273 13934 18307 13963
rect 18305 13930 18307 13934
rect 18341 13939 18343 13964
rect 18377 13939 18409 13965
rect 18341 13930 18409 13939
rect 18239 13900 18271 13929
rect 18305 13900 18375 13930
rect 18239 13895 18343 13900
rect 18239 13894 18307 13895
rect 18273 13861 18307 13894
rect 18341 13866 18343 13895
rect 18377 13866 18409 13896
rect 18341 13861 18409 13866
rect 18239 13827 18271 13860
rect 18305 13827 18375 13861
rect 18239 13826 18343 13827
rect 18239 13825 18307 13826
rect 18273 13792 18307 13825
rect 18341 13793 18343 13826
rect 18377 13793 18409 13827
rect 18341 13792 18409 13793
rect 18273 13791 18375 13792
rect 18239 13788 18375 13791
rect 18239 13756 18271 13788
rect 18305 13758 18375 13788
rect 18305 13757 18409 13758
rect 18305 13754 18307 13757
rect 18273 13723 18307 13754
rect 18341 13754 18409 13757
rect 18341 13723 18343 13754
rect 18377 13723 18409 13754
rect 18273 13722 18343 13723
rect 18239 13720 18343 13722
rect 18239 13715 18375 13720
rect 18239 13687 18271 13715
rect 18305 13689 18375 13715
rect 18305 13688 18409 13689
rect 18305 13681 18307 13688
rect 18273 13654 18307 13681
rect 18341 13681 18409 13688
rect 18341 13654 18343 13681
rect 18377 13654 18409 13681
rect 18273 13653 18343 13654
rect 18239 13647 18343 13653
rect 18239 13642 18375 13647
rect 18239 13618 18271 13642
rect 18305 13620 18375 13642
rect 18305 13619 18409 13620
rect 18305 13608 18307 13619
rect 18273 13585 18307 13608
rect 18341 13608 18409 13619
rect 18341 13585 18343 13608
rect 18377 13585 18409 13608
rect 18273 13584 18343 13585
rect 18239 13574 18343 13584
rect 18239 13569 18375 13574
rect 18239 13549 18271 13569
rect 18305 13551 18375 13569
rect 18305 13550 18409 13551
rect 18305 13535 18307 13550
rect 18273 13516 18307 13535
rect 18341 13535 18409 13550
rect 18341 13516 18343 13535
rect 18377 13516 18409 13535
rect 18273 13515 18343 13516
rect 18239 13501 18343 13515
rect 18239 13496 18375 13501
rect 18239 13480 18271 13496
rect 18305 13482 18375 13496
rect 18305 13481 18409 13482
rect 18305 13462 18307 13481
rect 18273 13447 18307 13462
rect 18341 13462 18409 13481
rect 18341 13447 18343 13462
rect 18377 13447 18409 13462
rect 18273 13446 18343 13447
rect 18239 13428 18343 13446
rect 18239 13423 18375 13428
rect 18239 13411 18271 13423
rect 18305 13413 18375 13423
rect 18305 13412 18409 13413
rect 18305 13389 18307 13412
rect 18273 13378 18307 13389
rect 18341 13389 18409 13412
rect 18341 13378 18343 13389
rect 18377 13378 18409 13389
rect 18273 13377 18343 13378
rect 18239 13355 18343 13377
rect 18239 13350 18375 13355
rect 18239 13342 18271 13350
rect 18305 13344 18375 13350
rect 18305 13343 18409 13344
rect 18305 13316 18307 13343
rect 18273 13309 18307 13316
rect 18341 13316 18409 13343
rect 18341 13309 18343 13316
rect 18377 13309 18409 13316
rect 18273 13308 18343 13309
rect 18239 13282 18343 13308
rect 18239 13277 18375 13282
rect 18239 13273 18271 13277
rect 18305 13275 18375 13277
rect 18305 13274 18409 13275
rect 18305 13243 18307 13274
rect 18273 13240 18307 13243
rect 18341 13243 18409 13274
rect 18341 13240 18343 13243
rect 18377 13240 18409 13243
rect 18273 13239 18343 13240
rect 18239 13209 18343 13239
rect 18239 13206 18375 13209
rect 18239 13205 18409 13206
rect 18239 13204 18307 13205
rect 18305 13171 18307 13204
rect 18341 13171 18409 13205
rect 18305 13170 18375 13171
rect 18239 13136 18343 13170
rect 18377 13136 18409 13137
rect 18239 13135 18307 13136
rect 18273 13131 18307 13135
rect 18305 13102 18307 13131
rect 18341 13102 18409 13136
rect 18239 13097 18271 13101
rect 18305 13097 18375 13102
rect 18239 13067 18343 13097
rect 18239 13066 18307 13067
rect 18273 13058 18307 13066
rect 18305 13033 18307 13058
rect 18341 13063 18343 13067
rect 18377 13063 18409 13068
rect 18341 13033 18409 13063
rect 18239 13024 18271 13032
rect 18305 13024 18375 13033
rect 18239 12998 18343 13024
rect 18239 12997 18307 12998
rect 18273 12985 18307 12997
rect 18305 12964 18307 12985
rect 18341 12990 18343 12998
rect 18377 12990 18409 12999
rect 18341 12964 18409 12990
rect 18239 12951 18271 12963
rect 18305 12951 18375 12964
rect 18239 12929 18343 12951
rect 18239 12928 18307 12929
rect 18273 12912 18307 12928
rect 18305 12895 18307 12912
rect 18341 12917 18343 12929
rect 18377 12917 18409 12930
rect 18341 12895 18409 12917
rect 18239 12878 18271 12894
rect 18305 12878 18375 12895
rect 18239 12860 18343 12878
rect 18239 12859 18307 12860
rect 18273 12839 18307 12859
rect 18305 12826 18307 12839
rect 18341 12844 18343 12860
rect 18377 12844 18409 12861
rect 18341 12826 18409 12844
rect 18239 12805 18271 12825
rect 18305 12805 18375 12826
rect 323 12759 391 12794
rect 357 12755 391 12759
rect 323 12721 357 12725
rect 323 12689 391 12721
rect 357 12682 391 12689
rect 323 12648 357 12655
rect 18239 12791 18343 12805
rect 18239 12790 18307 12791
rect 18273 12766 18307 12790
rect 18305 12757 18307 12766
rect 18341 12771 18343 12791
rect 18377 12771 18409 12792
rect 18341 12757 18409 12771
rect 18239 12732 18271 12756
rect 18305 12732 18375 12757
rect 18239 12722 18343 12732
rect 18239 12721 18307 12722
rect 18273 12693 18307 12721
rect 18305 12688 18307 12693
rect 18341 12698 18343 12722
rect 18377 12698 18409 12723
rect 18341 12688 18409 12698
rect 18239 12659 18271 12687
rect 18305 12659 18375 12688
rect 18239 12653 18343 12659
rect 18239 12652 18307 12653
rect 323 12620 391 12648
rect 357 12618 391 12620
rect 493 12618 528 12652
rect 562 12618 597 12652
rect 631 12618 666 12652
rect 700 12618 735 12652
rect 769 12618 804 12652
rect 838 12618 873 12652
rect 907 12618 942 12652
rect 976 12618 1011 12652
rect 1045 12618 1080 12652
rect 1114 12618 1149 12652
rect 1183 12618 1218 12652
rect 1252 12618 1287 12652
rect 1321 12618 1356 12652
rect 1390 12618 1425 12652
rect 1459 12618 1494 12652
rect 1528 12618 1563 12652
rect 1597 12618 1632 12652
rect 1666 12618 1701 12652
rect 1735 12618 1770 12652
rect 1804 12618 1839 12652
rect 1873 12618 1908 12652
rect 1942 12618 1977 12652
rect 2011 12618 2046 12652
rect 2080 12618 2115 12652
rect 2149 12618 2184 12652
rect 2218 12618 2253 12652
rect 2287 12618 2322 12652
rect 2356 12618 2391 12652
rect 2425 12618 2460 12652
rect 2494 12618 2529 12652
rect 2563 12618 2598 12652
rect 2632 12623 2667 12652
rect 357 12609 2529 12618
rect 323 12575 357 12586
rect 391 12584 429 12609
rect 463 12589 2529 12609
rect 2563 12589 2602 12618
rect 2636 12589 2667 12623
rect 463 12584 2667 12589
rect 323 12550 391 12575
rect 425 12575 429 12584
rect 425 12550 460 12575
rect 494 12550 529 12584
rect 563 12550 598 12584
rect 632 12550 667 12584
rect 701 12550 736 12584
rect 770 12550 805 12584
rect 839 12550 874 12584
rect 908 12550 943 12584
rect 977 12550 1012 12584
rect 1046 12550 1081 12584
rect 1115 12550 1150 12584
rect 1184 12550 1219 12584
rect 1253 12550 1288 12584
rect 1322 12550 1357 12584
rect 1391 12550 1426 12584
rect 1460 12550 1495 12584
rect 1529 12550 1564 12584
rect 1598 12550 1633 12584
rect 1667 12550 1702 12584
rect 1736 12550 1771 12584
rect 1805 12550 1840 12584
rect 1874 12550 1909 12584
rect 1943 12550 1978 12584
rect 2012 12550 2047 12584
rect 2081 12550 2116 12584
rect 2150 12550 2185 12584
rect 2219 12550 2254 12584
rect 2288 12550 2323 12584
rect 2357 12550 2392 12584
rect 2426 12550 2461 12584
rect 2495 12551 2530 12584
rect 2495 12550 2529 12551
rect 2564 12550 2599 12584
rect 323 12536 2529 12550
rect 323 12482 357 12536
rect 391 12516 429 12536
rect 463 12517 2529 12536
rect 2563 12517 2599 12550
rect 18273 12620 18307 12652
rect 18305 12619 18307 12620
rect 18341 12625 18343 12653
rect 18377 12625 18409 12654
rect 18341 12619 18409 12625
rect 18305 12586 18375 12619
rect 18273 12584 18343 12586
rect 18341 12552 18343 12584
rect 18377 12552 18409 12585
rect 18341 12550 18409 12552
rect 463 12516 2599 12517
rect 391 12482 426 12516
rect 463 12502 495 12516
rect 460 12482 495 12502
rect 529 12482 564 12516
rect 598 12482 633 12516
rect 667 12482 702 12516
rect 736 12482 771 12516
rect 805 12482 840 12516
rect 874 12482 909 12516
rect 943 12482 978 12516
rect 1012 12482 1047 12516
rect 1081 12482 1116 12516
rect 1150 12482 1185 12516
rect 1219 12482 1254 12516
rect 1288 12482 1323 12516
rect 1357 12482 1392 12516
rect 1426 12482 1461 12516
rect 1495 12482 1530 12516
rect 1564 12482 1599 12516
rect 1633 12482 1668 12516
rect 1702 12482 1737 12516
rect 1771 12482 1806 12516
rect 1840 12482 1875 12516
rect 1909 12482 1944 12516
rect 1978 12482 2013 12516
rect 2047 12482 2082 12516
rect 2116 12482 2151 12516
rect 2185 12482 2220 12516
rect 2254 12482 2289 12516
rect 2323 12482 2358 12516
rect 2392 12482 2427 12516
rect 2461 12482 2496 12516
rect 2530 12482 2565 12516
rect 18307 12516 18375 12550
rect 18307 12482 18409 12516
rect 0 12253 170 12285
rect 18609 12318 18677 12353
rect 18643 12285 18677 12318
rect 18643 12284 18745 12285
rect 18609 12253 18745 12284
rect 0 12251 18745 12253
rect 0 12250 18779 12251
rect 0 12249 18677 12250
rect 0 12215 18124 12249
rect 18158 12215 18194 12249
rect 18228 12215 18264 12249
rect 18298 12215 18333 12249
rect 18367 12215 18402 12249
rect 18436 12215 18471 12249
rect 18505 12215 18540 12249
rect 18574 12215 18609 12249
rect 18643 12216 18677 12249
rect 18711 12216 18779 12250
rect 18643 12215 18745 12216
rect 0 12182 18745 12215
rect 0 12181 18779 12182
rect 0 12147 18124 12181
rect 18158 12147 18194 12181
rect 18228 12147 18263 12181
rect 18297 12147 18332 12181
rect 18366 12147 18401 12181
rect 18435 12147 18470 12181
rect 18504 12147 18539 12181
rect 18573 12147 18608 12181
rect 18642 12147 18677 12181
rect 18711 12147 18779 12181
rect 0 12113 18745 12147
rect 0 12079 18124 12113
rect 18158 12079 18197 12113
rect 18231 12079 18270 12113
rect 18304 12079 18343 12113
rect 18377 12079 18416 12113
rect 18450 12079 18489 12113
rect 18523 12079 18562 12113
rect 18596 12079 18635 12113
rect 18669 12079 18779 12113
rect 11972 7691 12142 12079
rect 17920 7691 18090 12079
rect 11972 7659 18090 7691
rect 11972 7625 17016 7659
rect 17050 7625 18090 7659
rect 11972 7521 18090 7625
rect 10135 3692 10237 3726
rect 14555 3694 14590 3726
rect 14624 3694 14659 3726
rect 14693 3694 14728 3726
rect 14762 3694 14797 3726
rect 14831 3694 14866 3726
rect 14900 3694 14935 3726
rect 14969 3694 15004 3726
rect 15038 3694 15073 3726
rect 10169 3658 10237 3692
rect 10135 3656 10203 3658
rect 10135 3622 10167 3656
rect 10201 3624 10203 3656
rect 10201 3622 10271 3624
rect 10135 3617 10239 3622
rect 10169 3588 10239 3617
rect 14555 3692 14559 3694
rect 14624 3692 14632 3694
rect 14693 3692 14705 3694
rect 14762 3692 14778 3694
rect 14831 3692 14851 3694
rect 14900 3692 14924 3694
rect 14969 3692 14997 3694
rect 15038 3692 15070 3694
rect 15107 3692 15142 3726
rect 15176 3694 15211 3726
rect 15245 3694 15280 3726
rect 15314 3694 15349 3726
rect 15383 3694 15418 3726
rect 15452 3694 15487 3726
rect 15521 3694 15556 3726
rect 15590 3694 15625 3726
rect 15659 3694 15694 3726
rect 15728 3694 15763 3726
rect 15177 3692 15211 3694
rect 15250 3692 15280 3694
rect 15323 3692 15349 3694
rect 15396 3692 15418 3694
rect 15469 3692 15487 3694
rect 15542 3692 15556 3694
rect 15615 3692 15625 3694
rect 15688 3692 15694 3694
rect 15761 3692 15763 3694
rect 15797 3692 15831 3726
rect 14521 3660 14559 3692
rect 14593 3660 14632 3692
rect 14666 3660 14705 3692
rect 14739 3660 14778 3692
rect 14812 3660 14851 3692
rect 14885 3660 14924 3692
rect 14958 3660 14997 3692
rect 15031 3660 15070 3692
rect 15104 3660 15143 3692
rect 15177 3660 15216 3692
rect 15250 3660 15289 3692
rect 15323 3660 15362 3692
rect 15396 3660 15435 3692
rect 15469 3660 15508 3692
rect 15542 3660 15581 3692
rect 15615 3660 15654 3692
rect 15688 3660 15727 3692
rect 15761 3660 15831 3692
rect 14521 3658 15831 3660
rect 14521 3624 14556 3658
rect 14590 3624 14625 3658
rect 14659 3624 14694 3658
rect 14728 3624 14763 3658
rect 14797 3624 14832 3658
rect 14866 3624 14901 3658
rect 14935 3624 14970 3658
rect 15004 3624 15039 3658
rect 15073 3624 15108 3658
rect 15142 3624 15177 3658
rect 15211 3624 15246 3658
rect 15280 3624 15315 3658
rect 15349 3624 15384 3658
rect 15418 3624 15453 3658
rect 15487 3624 15522 3658
rect 15556 3624 15591 3658
rect 15625 3624 15660 3658
rect 15694 3624 15729 3658
rect 15763 3624 15831 3658
rect 14453 3622 15797 3624
rect 14486 3590 14525 3622
rect 14559 3590 14598 3622
rect 14632 3590 14671 3622
rect 14705 3590 14744 3622
rect 14778 3590 14817 3622
rect 14851 3590 14890 3622
rect 14924 3590 14963 3622
rect 14997 3590 15036 3622
rect 15070 3590 15109 3622
rect 15143 3590 15182 3622
rect 15216 3590 15255 3622
rect 15289 3590 15328 3622
rect 15362 3590 15401 3622
rect 15435 3590 15474 3622
rect 15508 3590 15547 3622
rect 15581 3590 15620 3622
rect 15654 3590 15693 3622
rect 15727 3590 15797 3622
rect 14486 3588 14488 3590
rect 10169 3587 10271 3588
rect 10169 3583 10203 3587
rect 10135 3576 10203 3583
rect 10135 3543 10167 3576
rect 10201 3553 10203 3576
rect 10237 3556 10271 3587
rect 14453 3556 14488 3588
rect 14522 3588 14525 3590
rect 14591 3588 14598 3590
rect 14660 3588 14671 3590
rect 14729 3588 14744 3590
rect 14798 3588 14817 3590
rect 14867 3588 14890 3590
rect 14936 3588 14963 3590
rect 15005 3588 15036 3590
rect 14522 3556 14557 3588
rect 14591 3556 14626 3588
rect 14660 3556 14695 3588
rect 14729 3556 14764 3588
rect 14798 3556 14833 3588
rect 14867 3556 14902 3588
rect 14936 3556 14971 3588
rect 15005 3556 15040 3588
rect 15074 3556 15109 3590
rect 15143 3556 15178 3590
rect 15216 3588 15247 3590
rect 15289 3588 15316 3590
rect 15362 3588 15385 3590
rect 15435 3588 15454 3590
rect 15508 3588 15523 3590
rect 15581 3588 15592 3590
rect 15654 3588 15661 3590
rect 15727 3589 15831 3590
rect 15727 3588 15729 3589
rect 15212 3556 15247 3588
rect 15281 3556 15316 3588
rect 15350 3556 15385 3588
rect 15419 3556 15454 3588
rect 15488 3556 15523 3588
rect 15557 3556 15592 3588
rect 15626 3556 15661 3588
rect 15695 3556 15729 3588
rect 10237 3553 10305 3556
rect 10201 3546 10305 3553
rect 10201 3542 10239 3546
rect 10169 3516 10239 3542
rect 10273 3519 10305 3546
rect 10169 3509 10203 3516
rect 10135 3497 10203 3509
rect 10135 3469 10167 3497
rect 10201 3482 10203 3497
rect 10237 3512 10239 3516
rect 10237 3485 10271 3512
rect 10237 3482 10305 3485
rect 10201 3470 10305 3482
rect 10201 3463 10239 3470
rect 10169 3445 10239 3463
rect 10273 3448 10305 3470
rect 10169 3435 10203 3445
rect 10135 3418 10203 3435
rect 10135 3395 10167 3418
rect 10201 3411 10203 3418
rect 10237 3436 10239 3445
rect 10237 3414 10271 3436
rect 10237 3411 10305 3414
rect 10201 3394 10305 3411
rect 15661 3555 15729 3556
rect 15763 3582 15831 3589
rect 15763 3555 15765 3582
rect 15799 3556 15831 3582
rect 15661 3550 15765 3555
rect 15661 3521 15693 3550
rect 15727 3548 15765 3550
rect 15727 3522 15797 3548
rect 15727 3520 15831 3522
rect 15727 3516 15729 3520
rect 15695 3487 15729 3516
rect 15661 3486 15729 3487
rect 15763 3509 15831 3520
rect 15763 3486 15765 3509
rect 15799 3488 15831 3509
rect 15661 3478 15765 3486
rect 15661 3452 15693 3478
rect 15727 3475 15765 3478
rect 15727 3454 15797 3475
rect 15727 3451 15831 3454
rect 15727 3444 15729 3451
rect 15695 3418 15729 3444
rect 15661 3417 15729 3418
rect 15763 3436 15831 3451
rect 15763 3417 15765 3436
rect 15799 3420 15831 3436
rect 15661 3406 15765 3417
rect 10201 3384 10239 3394
rect 10169 3374 10239 3384
rect 10273 3377 10305 3394
rect 10169 3361 10203 3374
rect 10135 3340 10203 3361
rect 10237 3360 10239 3374
rect 10237 3343 10271 3360
rect 10237 3340 10305 3343
rect 10135 3339 10305 3340
rect 10135 3321 10167 3339
rect 10201 3319 10305 3339
rect 10201 3305 10239 3319
rect 10273 3306 10305 3319
rect 10169 3303 10239 3305
rect 10169 3287 10203 3303
rect 10135 3269 10203 3287
rect 10237 3285 10239 3303
rect 10237 3272 10271 3285
rect 10237 3269 10305 3272
rect 10135 3260 10305 3269
rect 10135 3247 10167 3260
rect 10201 3244 10305 3260
rect 10201 3232 10239 3244
rect 10273 3235 10305 3244
rect 10201 3226 10203 3232
rect 10169 3213 10203 3226
rect 10135 3198 10203 3213
rect 10237 3210 10239 3232
rect 10237 3201 10271 3210
rect 10237 3198 10305 3201
rect 10135 3181 10305 3198
rect 10135 3173 10167 3181
rect 10201 3169 10305 3181
rect 10201 3161 10239 3169
rect 10273 3164 10305 3169
rect 10201 3147 10203 3161
rect 10169 3139 10203 3147
rect 10135 3127 10203 3139
rect 10237 3135 10239 3161
rect 10237 3130 10271 3135
rect 10237 3127 10305 3130
rect 10135 3102 10305 3127
rect 10135 3099 10167 3102
rect 10201 3094 10305 3102
rect 10201 3091 10239 3094
rect 10273 3093 10305 3094
rect 10201 3068 10203 3091
rect 10169 3065 10203 3068
rect 10135 3057 10203 3065
rect 10237 3060 10239 3091
rect 10237 3059 10271 3060
rect 10237 3057 10305 3059
rect 10135 3025 10305 3057
rect 10169 3023 10305 3025
rect 10201 3022 10305 3023
rect 10201 3021 10271 3022
rect 10135 2989 10167 2991
rect 10201 2989 10203 3021
rect 10135 2987 10203 2989
rect 10237 3019 10271 3021
rect 10237 2987 10239 3019
rect 10135 2985 10239 2987
rect 10273 2985 10305 2988
rect 10135 2951 10305 2985
rect 10169 2944 10203 2951
rect 10201 2917 10203 2944
rect 10237 2944 10271 2951
rect 10237 2917 10239 2944
rect 10135 2910 10167 2917
rect 10201 2910 10239 2917
rect 10273 2910 10305 2917
rect 10135 236 10305 2910
rect 10491 3380 10737 3404
rect 10525 3346 10559 3380
rect 10593 3346 10627 3380
rect 10661 3373 10737 3380
rect 12267 3373 12301 3404
rect 12335 3373 12369 3404
rect 12403 3373 12437 3404
rect 12471 3373 12505 3404
rect 12539 3373 12573 3404
rect 12607 3373 12641 3404
rect 12675 3373 12709 3404
rect 12743 3373 12777 3404
rect 12811 3373 12845 3404
rect 12879 3373 12913 3404
rect 12947 3373 12981 3404
rect 13015 3373 13049 3404
rect 13083 3373 13117 3404
rect 13151 3373 13185 3404
rect 13219 3373 13253 3404
rect 13287 3373 13321 3404
rect 13355 3373 13389 3404
rect 13423 3373 13457 3404
rect 13491 3373 13525 3404
rect 13559 3373 13593 3404
rect 13627 3373 13661 3404
rect 10491 3335 10633 3346
rect 10491 3310 10523 3335
rect 10557 3311 10633 3335
rect 10557 3301 10559 3311
rect 10525 3277 10559 3301
rect 10593 3301 10627 3311
rect 10593 3277 10595 3301
rect 13653 3339 13657 3373
rect 13695 3370 13729 3404
rect 13763 3370 13797 3404
rect 13831 3373 13865 3404
rect 13899 3373 13933 3404
rect 13967 3373 14001 3404
rect 14035 3373 14069 3404
rect 14103 3373 14137 3404
rect 14171 3373 14205 3404
rect 14239 3373 14273 3404
rect 13835 3370 13865 3373
rect 13907 3370 13933 3373
rect 13979 3370 14001 3373
rect 14052 3370 14069 3373
rect 14125 3370 14137 3373
rect 14198 3370 14205 3373
rect 14271 3370 14273 3373
rect 14307 3373 14341 3404
rect 14375 3373 14409 3404
rect 14443 3373 14477 3404
rect 14511 3373 14545 3404
rect 14579 3373 14613 3404
rect 14647 3373 14682 3404
rect 14716 3373 14751 3404
rect 14307 3370 14310 3373
rect 14375 3370 14383 3373
rect 14443 3370 14456 3373
rect 14511 3370 14529 3373
rect 14579 3370 14602 3373
rect 14647 3370 14675 3373
rect 14716 3370 14748 3373
rect 14785 3370 14820 3404
rect 14854 3373 14889 3404
rect 14923 3373 14958 3404
rect 14992 3373 15027 3404
rect 15061 3373 15096 3404
rect 15130 3373 15165 3404
rect 15199 3373 15234 3404
rect 15268 3373 15303 3404
rect 15337 3373 15372 3404
rect 15406 3373 15441 3404
rect 14855 3370 14889 3373
rect 14928 3370 14958 3373
rect 15001 3370 15027 3373
rect 15074 3370 15096 3373
rect 15147 3370 15165 3373
rect 15220 3370 15234 3373
rect 15293 3370 15303 3373
rect 15366 3370 15372 3373
rect 15439 3370 15441 3373
rect 15475 3370 15509 3404
rect 13691 3339 13729 3370
rect 13763 3339 13801 3370
rect 13835 3339 13873 3370
rect 13907 3339 13945 3370
rect 13979 3339 14018 3370
rect 14052 3339 14091 3370
rect 14125 3339 14164 3370
rect 14198 3339 14237 3370
rect 14271 3339 14310 3370
rect 14344 3339 14383 3370
rect 14417 3339 14456 3370
rect 14490 3339 14529 3370
rect 14563 3339 14602 3370
rect 14636 3339 14675 3370
rect 14709 3339 14748 3370
rect 14782 3339 14821 3370
rect 14855 3339 14894 3370
rect 14928 3339 14967 3370
rect 15001 3339 15040 3370
rect 15074 3339 15113 3370
rect 15147 3339 15186 3370
rect 15220 3339 15259 3370
rect 15293 3339 15332 3370
rect 15366 3339 15405 3370
rect 15439 3339 15509 3370
rect 13653 3336 15509 3339
rect 13653 3302 13682 3336
rect 13716 3302 13751 3336
rect 13785 3302 13820 3336
rect 13854 3302 13889 3336
rect 13923 3302 13958 3336
rect 13992 3302 14027 3336
rect 14061 3302 14096 3336
rect 14130 3302 14165 3336
rect 14199 3302 14234 3336
rect 14268 3302 14303 3336
rect 14337 3302 14372 3336
rect 14406 3302 14441 3336
rect 14475 3302 14510 3336
rect 14544 3302 14579 3336
rect 14613 3302 14648 3336
rect 14682 3302 14717 3336
rect 14751 3302 14786 3336
rect 14820 3302 14855 3336
rect 14889 3302 14924 3336
rect 14958 3302 14993 3336
rect 15027 3302 15062 3336
rect 15096 3302 15131 3336
rect 15165 3302 15200 3336
rect 15234 3302 15269 3336
rect 15303 3302 15338 3336
rect 15372 3302 15407 3336
rect 15441 3302 15509 3336
rect 10525 3276 10595 3277
rect 10491 3267 10595 3276
rect 10629 3267 10633 3277
rect 13653 3301 15509 3302
rect 13653 3268 13692 3301
rect 13726 3268 13765 3301
rect 13799 3268 13838 3301
rect 13872 3268 13911 3301
rect 13945 3268 13984 3301
rect 14018 3268 14057 3301
rect 14091 3268 14130 3301
rect 14164 3268 14203 3301
rect 14237 3268 14276 3301
rect 14310 3268 14349 3301
rect 14383 3268 14422 3301
rect 14456 3268 14495 3301
rect 14529 3268 14568 3301
rect 14602 3268 14641 3301
rect 14675 3268 14714 3301
rect 14748 3268 14787 3301
rect 14821 3268 14860 3301
rect 14894 3268 14933 3301
rect 14967 3268 15006 3301
rect 15040 3268 15079 3301
rect 15113 3268 15152 3301
rect 15186 3268 15225 3301
rect 15259 3268 15298 3301
rect 15332 3268 15371 3301
rect 15405 3300 15509 3301
rect 13653 3267 13683 3268
rect 13726 3267 13752 3268
rect 13799 3267 13821 3268
rect 13872 3267 13890 3268
rect 13945 3267 13959 3268
rect 14018 3267 14028 3268
rect 14091 3267 14097 3268
rect 14164 3267 14166 3268
rect 10491 3262 10737 3267
rect 10491 3240 10523 3262
rect 10557 3242 10737 3262
rect 10557 3228 10559 3242
rect 10525 3208 10559 3228
rect 10593 3227 10627 3242
rect 10661 3234 10737 3242
rect 12199 3234 12234 3267
rect 12268 3234 12303 3267
rect 12337 3234 12372 3267
rect 12406 3234 12441 3267
rect 12475 3234 12510 3267
rect 12544 3234 12579 3267
rect 12613 3234 12648 3267
rect 12682 3234 12717 3267
rect 12751 3234 12786 3267
rect 12820 3234 12855 3267
rect 12889 3234 12924 3267
rect 12958 3234 12993 3267
rect 13027 3234 13062 3267
rect 13096 3234 13131 3267
rect 13165 3234 13200 3267
rect 13234 3234 13269 3267
rect 13303 3234 13338 3267
rect 13372 3234 13407 3267
rect 13441 3234 13476 3267
rect 13510 3234 13545 3267
rect 13579 3234 13614 3267
rect 13648 3234 13683 3267
rect 13717 3234 13752 3267
rect 13786 3234 13821 3267
rect 13855 3234 13890 3267
rect 13924 3234 13959 3267
rect 13993 3234 14028 3267
rect 14062 3234 14097 3267
rect 14131 3234 14166 3267
rect 14200 3267 14203 3268
rect 14269 3267 14276 3268
rect 14338 3267 14349 3268
rect 14407 3267 14422 3268
rect 14476 3267 14495 3268
rect 14545 3267 14568 3268
rect 14614 3267 14641 3268
rect 14683 3267 14714 3268
rect 14200 3234 14235 3267
rect 14269 3234 14304 3267
rect 14338 3234 14373 3267
rect 14407 3234 14442 3267
rect 14476 3234 14511 3267
rect 14545 3234 14580 3267
rect 14614 3234 14649 3267
rect 14683 3234 14718 3267
rect 14752 3234 14787 3268
rect 14821 3234 14856 3268
rect 14894 3267 14925 3268
rect 14967 3267 14994 3268
rect 15040 3267 15063 3268
rect 15113 3267 15132 3268
rect 15186 3267 15201 3268
rect 15259 3267 15270 3268
rect 15332 3267 15339 3268
rect 15405 3267 15475 3300
rect 14890 3234 14925 3267
rect 14959 3234 14994 3267
rect 15028 3234 15063 3267
rect 15097 3234 15132 3267
rect 15166 3234 15201 3267
rect 15235 3234 15270 3267
rect 15304 3234 15339 3267
rect 15373 3234 15407 3267
rect 10593 3208 10595 3227
rect 10525 3206 10595 3208
rect 10491 3193 10595 3206
rect 10629 3193 10661 3208
rect 10491 3189 10661 3193
rect 10491 3170 10523 3189
rect 10557 3173 10661 3189
rect 10557 3155 10559 3173
rect 10525 3139 10559 3155
rect 10593 3153 10627 3173
rect 10593 3139 10595 3153
rect 10525 3136 10595 3139
rect 10491 3119 10595 3136
rect 10629 3119 10661 3139
rect 10491 3116 10661 3119
rect 10491 3100 10523 3116
rect 10557 3104 10661 3116
rect 10557 3082 10559 3104
rect 10525 3070 10559 3082
rect 10593 3079 10627 3104
rect 10593 3070 10595 3079
rect 10525 3066 10595 3070
rect 10491 3045 10595 3066
rect 10629 3045 10661 3070
rect 10491 3043 10661 3045
rect 10491 3030 10523 3043
rect 10557 3035 10661 3043
rect 10557 3009 10559 3035
rect 10525 3001 10559 3009
rect 10593 3005 10627 3035
rect 10593 3001 10595 3005
rect 10525 2996 10595 3001
rect 10491 2971 10595 2996
rect 10629 2971 10661 3001
rect 10491 2970 10661 2971
rect 10491 2960 10523 2970
rect 10557 2966 10661 2970
rect 10557 2936 10559 2966
rect 10525 2932 10559 2936
rect 10593 2932 10627 2966
rect 10525 2931 10661 2932
rect 10525 2926 10595 2931
rect 10491 2898 10595 2926
rect 10491 2890 10523 2898
rect 10557 2897 10595 2898
rect 10629 2897 10661 2931
rect 10557 2864 10559 2897
rect 10525 2863 10559 2864
rect 10593 2863 10627 2897
rect 10525 2857 10661 2863
rect 10525 2856 10595 2857
rect 10491 2828 10595 2856
rect 10629 2828 10661 2857
rect 10491 2826 10559 2828
rect 10491 2820 10523 2826
rect 10557 2794 10559 2826
rect 10593 2823 10595 2828
rect 10593 2794 10627 2823
rect 10557 2792 10661 2794
rect 10525 2786 10661 2792
rect 10491 2783 10661 2786
rect 10491 2759 10595 2783
rect 10629 2759 10661 2783
rect 10491 2754 10559 2759
rect 10491 2750 10523 2754
rect 10557 2725 10559 2754
rect 10593 2749 10595 2759
rect 10593 2725 10627 2749
rect 10557 2720 10661 2725
rect 10525 2716 10661 2720
rect 10491 2709 10661 2716
rect 10491 2690 10595 2709
rect 10629 2690 10661 2709
rect 10491 2682 10559 2690
rect 10491 2680 10523 2682
rect 10557 2656 10559 2682
rect 10593 2675 10595 2690
rect 10593 2656 10627 2675
rect 10557 2648 10661 2656
rect 10525 2646 10661 2648
rect 10491 2636 10661 2646
rect 10491 2621 10595 2636
rect 10629 2621 10661 2636
rect 10491 2610 10559 2621
rect 10557 2587 10559 2610
rect 10593 2602 10595 2621
rect 10593 2587 10627 2602
rect 10557 2576 10661 2587
rect 10491 2563 10661 2576
rect 10491 2552 10595 2563
rect 10629 2552 10661 2563
rect 10491 2540 10559 2552
rect 10525 2538 10559 2540
rect 10557 2518 10559 2538
rect 10593 2529 10595 2552
rect 10593 2518 10627 2529
rect 10491 2504 10523 2506
rect 10557 2504 10661 2518
rect 10491 2490 10661 2504
rect 10491 2483 10595 2490
rect 10629 2483 10661 2490
rect 10491 2470 10559 2483
rect 10525 2466 10559 2470
rect 10557 2449 10559 2466
rect 10593 2456 10595 2483
rect 10593 2449 10627 2456
rect 10491 2432 10523 2436
rect 10557 2432 10661 2449
rect 10491 2417 10661 2432
rect 10491 2414 10595 2417
rect 10629 2414 10661 2417
rect 10491 2400 10559 2414
rect 10525 2394 10559 2400
rect 10557 2380 10559 2394
rect 10593 2383 10595 2414
rect 15339 3233 15407 3234
rect 15441 3266 15475 3267
rect 15441 3261 15509 3266
rect 15441 3233 15443 3261
rect 15339 3228 15443 3233
rect 15477 3231 15509 3261
rect 15339 3199 15371 3228
rect 15405 3227 15443 3228
rect 15405 3198 15475 3227
rect 15405 3194 15407 3198
rect 15373 3165 15407 3194
rect 15339 3164 15407 3165
rect 15441 3197 15475 3198
rect 15441 3188 15509 3197
rect 15441 3164 15443 3188
rect 15339 3155 15443 3164
rect 15477 3162 15509 3188
rect 15339 3130 15371 3155
rect 15405 3154 15443 3155
rect 15405 3129 15475 3154
rect 15405 3121 15407 3129
rect 15373 3096 15407 3121
rect 15339 3095 15407 3096
rect 15441 3128 15475 3129
rect 15441 3115 15509 3128
rect 15441 3095 15443 3115
rect 15339 3082 15443 3095
rect 15477 3093 15509 3115
rect 15339 3061 15371 3082
rect 15405 3081 15443 3082
rect 15405 3060 15475 3081
rect 15405 3048 15407 3060
rect 15373 3027 15407 3048
rect 15339 3026 15407 3027
rect 15441 3059 15475 3060
rect 15441 3042 15509 3059
rect 15441 3026 15443 3042
rect 15339 3009 15443 3026
rect 15477 3024 15509 3042
rect 15339 2992 15371 3009
rect 15405 3008 15443 3009
rect 15405 2991 15475 3008
rect 15405 2975 15407 2991
rect 15373 2958 15407 2975
rect 15339 2957 15407 2958
rect 15441 2990 15475 2991
rect 15441 2969 15509 2990
rect 15441 2957 15443 2969
rect 15339 2936 15443 2957
rect 15477 2955 15509 2969
rect 15339 2923 15371 2936
rect 15405 2935 15443 2936
rect 15405 2922 15475 2935
rect 15405 2902 15407 2922
rect 15373 2889 15407 2902
rect 15339 2888 15407 2889
rect 15441 2921 15475 2922
rect 15441 2896 15509 2921
rect 15441 2888 15443 2896
rect 15339 2863 15443 2888
rect 15477 2886 15509 2896
rect 15339 2854 15371 2863
rect 15405 2862 15443 2863
rect 15405 2853 15475 2862
rect 15405 2829 15407 2853
rect 15373 2820 15407 2829
rect 15339 2819 15407 2820
rect 15441 2852 15475 2853
rect 15441 2823 15509 2852
rect 15441 2819 15443 2823
rect 15339 2790 15443 2819
rect 15477 2817 15509 2823
rect 15339 2785 15371 2790
rect 15405 2789 15443 2790
rect 15405 2784 15475 2789
rect 15405 2756 15407 2784
rect 15373 2751 15407 2756
rect 15339 2750 15407 2751
rect 15441 2783 15475 2784
rect 15441 2750 15509 2783
rect 15339 2717 15443 2750
rect 15477 2748 15509 2750
rect 15339 2716 15371 2717
rect 15405 2716 15443 2717
rect 15405 2715 15475 2716
rect 15405 2683 15407 2715
rect 15373 2682 15407 2683
rect 15339 2681 15407 2682
rect 15441 2714 15475 2715
rect 15441 2681 15509 2714
rect 15339 2679 15509 2681
rect 15339 2677 15475 2679
rect 15339 2647 15443 2677
rect 15373 2646 15443 2647
rect 15373 2644 15407 2646
rect 15339 2610 15371 2613
rect 15405 2612 15407 2644
rect 15441 2643 15443 2646
rect 15477 2643 15509 2645
rect 15441 2612 15509 2643
rect 15405 2610 15509 2612
rect 15339 2604 15475 2610
rect 15339 2578 15443 2604
rect 15373 2577 15443 2578
rect 15373 2571 15407 2577
rect 15339 2537 15371 2544
rect 15405 2543 15407 2571
rect 15441 2570 15443 2577
rect 15477 2570 15509 2576
rect 15441 2543 15509 2570
rect 15405 2541 15509 2543
rect 15405 2537 15475 2541
rect 15339 2531 15475 2537
rect 15339 2509 15443 2531
rect 15373 2508 15443 2509
rect 15373 2498 15407 2508
rect 15339 2464 15371 2475
rect 15405 2474 15407 2498
rect 15441 2497 15443 2508
rect 15477 2497 15509 2507
rect 15441 2474 15509 2497
rect 15405 2472 15509 2474
rect 15405 2464 15475 2472
rect 15339 2458 15475 2464
rect 15339 2440 15443 2458
rect 15373 2439 15443 2440
rect 15373 2425 15407 2439
rect 10593 2380 10627 2383
rect 10491 2360 10523 2366
rect 10557 2360 10661 2380
rect 10491 2345 10661 2360
rect 10491 2330 10559 2345
rect 10525 2322 10559 2330
rect 10557 2311 10559 2322
rect 10593 2344 10627 2345
rect 10593 2311 10595 2344
rect 10557 2310 10595 2311
rect 10629 2310 10661 2311
rect 10491 2288 10523 2296
rect 10557 2288 10661 2310
rect 10491 2276 10661 2288
rect 10491 2260 10559 2276
rect 10525 2250 10559 2260
rect 10557 2242 10559 2250
rect 10593 2271 10627 2276
rect 10593 2242 10595 2271
rect 10557 2237 10595 2242
rect 10629 2237 10661 2242
rect 10491 2216 10523 2226
rect 10557 2216 10661 2237
rect 10491 2207 10661 2216
rect 10491 2190 10559 2207
rect 10525 2178 10559 2190
rect 10557 2173 10559 2178
rect 10593 2198 10627 2207
rect 10593 2173 10595 2198
rect 10557 2164 10595 2173
rect 10629 2164 10661 2173
rect 10491 2144 10523 2156
rect 10557 2144 10661 2164
rect 10491 2138 10661 2144
rect 10491 2120 10559 2138
rect 10525 2106 10559 2120
rect 10557 2104 10559 2106
rect 10593 2125 10627 2138
rect 10593 2104 10595 2125
rect 10557 2091 10595 2104
rect 10629 2091 10661 2104
rect 10491 2072 10523 2086
rect 10557 2072 10661 2091
rect 10491 2069 10661 2072
rect 10491 2050 10559 2069
rect 10525 2035 10559 2050
rect 10593 2052 10627 2069
rect 10593 2035 10595 2052
rect 10525 2034 10595 2035
rect 10557 2018 10595 2034
rect 10629 2018 10661 2035
rect 10491 2000 10523 2016
rect 10557 2000 10661 2018
rect 10491 1980 10559 2000
rect 10525 1966 10559 1980
rect 10593 1979 10627 2000
rect 10593 1966 10595 1979
rect 10525 1962 10595 1966
rect 10491 1928 10523 1946
rect 10557 1945 10595 1962
rect 10629 1945 10661 1966
rect 10557 1931 10661 1945
rect 10557 1928 10559 1931
rect 10491 1910 10559 1928
rect 10525 1897 10559 1910
rect 10593 1906 10627 1931
rect 10593 1897 10595 1906
rect 10525 1890 10595 1897
rect 10491 1856 10523 1876
rect 10557 1872 10595 1890
rect 10629 1872 10661 1897
rect 10557 1862 10661 1872
rect 10557 1856 10559 1862
rect 10491 1840 10559 1856
rect 10525 1828 10559 1840
rect 10593 1833 10627 1862
rect 10593 1828 10595 1833
rect 10525 1818 10595 1828
rect 10491 1784 10523 1806
rect 10557 1799 10595 1818
rect 10629 1799 10661 1828
rect 10557 1793 10661 1799
rect 10557 1784 10559 1793
rect 10491 1770 10559 1784
rect 10525 1759 10559 1770
rect 10593 1760 10627 1793
rect 10593 1759 10595 1760
rect 10525 1746 10595 1759
rect 10491 1712 10523 1736
rect 10557 1726 10595 1746
rect 10629 1726 10661 1759
rect 10557 1724 10661 1726
rect 10557 1712 10559 1724
rect 10491 1701 10559 1712
rect 10525 1690 10559 1701
rect 10593 1690 10627 1724
rect 10525 1687 10661 1690
rect 10525 1674 10595 1687
rect 10491 1640 10523 1667
rect 10557 1655 10595 1674
rect 10629 1655 10661 1687
rect 10557 1640 10559 1655
rect 10491 1632 10559 1640
rect 10525 1621 10559 1632
rect 10593 1653 10595 1655
rect 10593 1621 10627 1653
rect 10525 1614 10661 1621
rect 10525 1602 10595 1614
rect 10491 1568 10523 1598
rect 10557 1586 10595 1602
rect 10629 1586 10661 1614
rect 10557 1568 10559 1586
rect 10491 1563 10559 1568
rect 10525 1552 10559 1563
rect 10593 1580 10595 1586
rect 10593 1552 10627 1580
rect 10525 1541 10661 1552
rect 10525 1530 10595 1541
rect 10491 1496 10523 1529
rect 10557 1517 10595 1530
rect 10629 1517 10661 1541
rect 10709 2330 10743 2372
rect 10709 2253 10743 2296
rect 10709 2176 10743 2219
rect 10709 2099 10743 2142
rect 15257 2330 15291 2372
rect 15257 2253 15291 2296
rect 15257 2176 15291 2219
rect 10709 2022 10743 2065
rect 15257 2099 15291 2142
rect 15257 2022 15291 2065
rect 10709 1945 10743 1988
rect 10709 1868 10743 1911
rect 15257 1945 15291 1988
rect 10709 1791 10743 1834
rect 15257 1868 15291 1911
rect 10709 1714 10743 1757
rect 10709 1637 10743 1680
rect 10709 1560 10743 1603
rect 15257 1791 15291 1834
rect 15257 1714 15291 1757
rect 15257 1637 15291 1680
rect 15257 1560 15291 1603
rect 15339 2391 15371 2406
rect 15405 2405 15407 2425
rect 15441 2424 15443 2439
rect 15477 2424 15509 2438
rect 15441 2405 15509 2424
rect 15405 2403 15509 2405
rect 15405 2391 15475 2403
rect 15339 2385 15475 2391
rect 15339 2371 15443 2385
rect 15373 2370 15443 2371
rect 15373 2352 15407 2370
rect 15339 2318 15371 2337
rect 15405 2336 15407 2352
rect 15441 2351 15443 2370
rect 15477 2351 15509 2369
rect 15441 2336 15509 2351
rect 15405 2334 15509 2336
rect 15405 2318 15475 2334
rect 15339 2312 15475 2318
rect 15339 2302 15443 2312
rect 15373 2301 15443 2302
rect 15373 2279 15407 2301
rect 15339 2245 15371 2268
rect 15405 2267 15407 2279
rect 15441 2278 15443 2301
rect 15477 2278 15509 2300
rect 15441 2267 15509 2278
rect 15405 2265 15509 2267
rect 15405 2245 15475 2265
rect 15339 2239 15475 2245
rect 15339 2233 15443 2239
rect 15373 2232 15443 2233
rect 15373 2206 15407 2232
rect 15339 2172 15371 2199
rect 15405 2198 15407 2206
rect 15441 2205 15443 2232
rect 15477 2205 15509 2231
rect 15441 2198 15509 2205
rect 15405 2196 15509 2198
rect 15405 2172 15475 2196
rect 15339 2166 15475 2172
rect 15339 2164 15443 2166
rect 15373 2163 15443 2164
rect 15373 2133 15407 2163
rect 15339 2099 15371 2130
rect 15405 2129 15407 2133
rect 15441 2132 15443 2163
rect 15477 2132 15509 2162
rect 15441 2129 15509 2132
rect 15405 2127 15509 2129
rect 15405 2099 15475 2127
rect 15339 2095 15475 2099
rect 15373 2094 15475 2095
rect 15373 2061 15407 2094
rect 15339 2060 15407 2061
rect 15441 2093 15475 2094
rect 15441 2060 15443 2093
rect 15339 2026 15371 2060
rect 15405 2059 15443 2060
rect 15477 2059 15509 2093
rect 15405 2058 15509 2059
rect 15405 2026 15475 2058
rect 15373 2025 15475 2026
rect 15373 1992 15407 2025
rect 15339 1991 15407 1992
rect 15441 2024 15475 2025
rect 15441 2020 15509 2024
rect 15441 1991 15443 2020
rect 15339 1987 15443 1991
rect 15477 1989 15509 2020
rect 15339 1957 15371 1987
rect 15405 1986 15443 1987
rect 15405 1956 15475 1986
rect 15405 1953 15407 1956
rect 15373 1923 15407 1953
rect 15339 1922 15407 1923
rect 15441 1955 15475 1956
rect 15441 1947 15509 1955
rect 15441 1922 15443 1947
rect 15339 1914 15443 1922
rect 15477 1920 15509 1947
rect 15339 1888 15371 1914
rect 15405 1913 15443 1914
rect 15405 1887 15475 1913
rect 15405 1880 15407 1887
rect 15373 1854 15407 1880
rect 15339 1853 15407 1854
rect 15441 1886 15475 1887
rect 15441 1874 15509 1886
rect 15441 1853 15443 1874
rect 15339 1841 15443 1853
rect 15477 1851 15509 1874
rect 15339 1818 15371 1841
rect 15405 1840 15443 1841
rect 15405 1818 15475 1840
rect 15405 1807 15407 1818
rect 15373 1784 15407 1807
rect 15441 1817 15475 1818
rect 15441 1801 15509 1817
rect 15441 1784 15443 1801
rect 15339 1768 15443 1784
rect 15477 1782 15509 1801
rect 15339 1748 15371 1768
rect 15405 1767 15443 1768
rect 15405 1749 15475 1767
rect 15405 1734 15407 1749
rect 15373 1715 15407 1734
rect 15441 1748 15475 1749
rect 15441 1728 15509 1748
rect 15441 1715 15443 1728
rect 15373 1714 15443 1715
rect 15339 1695 15443 1714
rect 15477 1713 15509 1728
rect 15339 1678 15371 1695
rect 15405 1694 15443 1695
rect 15405 1680 15475 1694
rect 15405 1661 15407 1680
rect 15373 1646 15407 1661
rect 15441 1679 15475 1680
rect 15441 1655 15509 1679
rect 15441 1646 15443 1655
rect 15373 1644 15443 1646
rect 15477 1644 15509 1655
rect 15339 1622 15443 1644
rect 15339 1608 15371 1622
rect 15405 1621 15443 1622
rect 15405 1610 15475 1621
rect 15405 1588 15407 1610
rect 15373 1576 15407 1588
rect 15441 1582 15509 1610
rect 15441 1576 15443 1582
rect 15373 1574 15443 1576
rect 15477 1575 15509 1582
rect 15339 1549 15443 1574
rect 15339 1538 15371 1549
rect 15405 1548 15443 1549
rect 15405 1541 15475 1548
rect 15405 1540 15509 1541
rect 10557 1496 10559 1517
rect 10491 1494 10559 1496
rect 10525 1483 10559 1494
rect 10593 1507 10595 1517
rect 10593 1483 10627 1507
rect 10525 1468 10661 1483
rect 10525 1460 10595 1468
rect 10491 1458 10595 1460
rect 10491 1425 10523 1458
rect 10557 1448 10595 1458
rect 10629 1448 10661 1468
rect 10557 1424 10559 1448
rect 10525 1414 10559 1424
rect 10593 1434 10595 1448
rect 10593 1414 10627 1434
rect 10525 1395 10661 1414
rect 10525 1391 10595 1395
rect 10491 1386 10595 1391
rect 10491 1356 10523 1386
rect 10557 1379 10595 1386
rect 10629 1379 10661 1395
rect 10557 1352 10559 1379
rect 10525 1345 10559 1352
rect 10593 1361 10595 1379
rect 10593 1345 10627 1361
rect 10525 1322 10661 1345
rect 10491 1314 10595 1322
rect 10491 1287 10523 1314
rect 10557 1310 10595 1314
rect 10629 1310 10661 1322
rect 10557 1280 10559 1310
rect 10525 1253 10559 1280
rect 10491 1242 10559 1253
rect 10491 1218 10523 1242
rect 10557 1208 10559 1242
rect 10525 1184 10559 1208
rect 10491 1170 10559 1184
rect 10491 1149 10523 1170
rect 10557 1136 10559 1170
rect 10525 1115 10559 1136
rect 10491 1098 10559 1115
rect 10491 1080 10523 1098
rect 10557 1064 10559 1098
rect 10525 1046 10559 1064
rect 10491 1026 10559 1046
rect 10491 1011 10523 1026
rect 10557 992 10559 1026
rect 10525 977 10559 992
rect 10491 954 10559 977
rect 10491 942 10523 954
rect 10557 920 10559 954
rect 10525 908 10559 920
rect 10491 882 10559 908
rect 10491 873 10523 882
rect 10557 848 10559 882
rect 10525 839 10559 848
rect 10491 810 10559 839
rect 10491 804 10523 810
rect 10557 776 10559 810
rect 10525 770 10559 776
rect 10491 738 10559 770
rect 10491 735 10523 738
rect 10557 704 10559 738
rect 10525 701 10559 704
rect 10491 666 10559 701
rect 10525 665 10559 666
rect 15405 1515 15407 1540
rect 15373 1506 15407 1515
rect 15441 1509 15509 1540
rect 15441 1506 15443 1509
rect 15477 1506 15509 1509
rect 15373 1504 15443 1506
rect 15339 1476 15443 1504
rect 15339 1468 15371 1476
rect 15405 1475 15443 1476
rect 15405 1472 15475 1475
rect 15405 1470 15509 1472
rect 15405 1442 15407 1470
rect 15373 1436 15407 1442
rect 15441 1436 15509 1470
rect 15373 1434 15443 1436
rect 15339 1403 15443 1434
rect 15339 1398 15371 1403
rect 15405 1402 15443 1403
rect 15405 1400 15509 1402
rect 15405 1369 15407 1400
rect 15373 1366 15407 1369
rect 15441 1366 15509 1400
rect 15373 1364 15475 1366
rect 15339 1363 15475 1364
rect 15339 1330 15443 1363
rect 15339 1328 15371 1330
rect 15405 1296 15407 1330
rect 15441 1329 15443 1330
rect 15477 1329 15509 1332
rect 15441 1296 15509 1329
rect 15373 1294 15475 1296
rect 15339 1290 15475 1294
rect 15339 1260 15443 1290
rect 15339 1258 15407 1260
rect 15373 1257 15407 1258
rect 15405 1226 15407 1257
rect 15441 1256 15443 1260
rect 15477 1256 15509 1262
rect 15441 1226 15509 1256
rect 15339 1223 15371 1224
rect 15405 1223 15475 1226
rect 15339 1217 15475 1223
rect 15339 1190 15443 1217
rect 15339 1188 15407 1190
rect 15373 1183 15407 1188
rect 15405 1156 15407 1183
rect 15441 1183 15443 1190
rect 15477 1183 15509 1192
rect 15441 1156 15509 1183
rect 15339 1149 15371 1154
rect 15405 1149 15475 1156
rect 15339 1144 15475 1149
rect 15339 1120 15443 1144
rect 15339 1118 15407 1120
rect 15373 1109 15407 1118
rect 15405 1086 15407 1109
rect 15441 1110 15443 1120
rect 15477 1110 15509 1122
rect 15441 1086 15509 1110
rect 15339 1075 15371 1084
rect 15405 1075 15475 1086
rect 15339 1071 15475 1075
rect 15339 1050 15443 1071
rect 15339 1048 15407 1050
rect 15373 1035 15407 1048
rect 15405 1016 15407 1035
rect 15441 1037 15443 1050
rect 15477 1037 15509 1052
rect 15441 1016 15509 1037
rect 15339 1001 15371 1014
rect 15405 1001 15475 1016
rect 15339 998 15475 1001
rect 15339 980 15443 998
rect 15339 978 15407 980
rect 15373 961 15407 978
rect 15405 946 15407 961
rect 15441 964 15443 980
rect 15477 964 15509 982
rect 15441 946 15509 964
rect 15339 927 15371 944
rect 15405 927 15475 946
rect 15339 925 15475 927
rect 15339 910 15443 925
rect 15339 908 15407 910
rect 15373 887 15407 908
rect 15405 876 15407 887
rect 15441 891 15443 910
rect 15477 891 15509 912
rect 15441 876 15509 891
rect 15339 853 15371 874
rect 15405 853 15475 876
rect 15339 852 15475 853
rect 15339 840 15443 852
rect 15339 838 15407 840
rect 15373 813 15407 838
rect 15405 806 15407 813
rect 15441 818 15443 840
rect 15477 818 15509 842
rect 15441 806 15509 818
rect 15339 779 15371 804
rect 15405 779 15475 806
rect 15339 770 15443 779
rect 15339 768 15407 770
rect 15373 739 15407 768
rect 15405 736 15407 739
rect 15441 745 15443 770
rect 15477 745 15509 772
rect 15441 736 15509 745
rect 15339 705 15371 734
rect 15405 705 15475 736
rect 15339 700 15443 705
rect 15339 698 15407 700
rect 10661 665 10696 698
rect 10730 665 10765 698
rect 10799 665 10834 698
rect 10868 665 10903 698
rect 10937 665 10972 698
rect 11006 665 11041 698
rect 10525 632 10529 665
rect 10661 664 10675 665
rect 10730 664 10748 665
rect 10799 664 10821 665
rect 10868 664 10894 665
rect 10937 664 10967 665
rect 11006 664 11040 665
rect 11075 664 11110 698
rect 11144 665 11179 698
rect 11213 665 11248 698
rect 11282 665 11317 698
rect 11351 665 11386 698
rect 11420 665 11455 698
rect 11489 665 11524 698
rect 11558 665 11593 698
rect 11627 665 11662 698
rect 11147 664 11179 665
rect 11220 664 11248 665
rect 11293 664 11317 665
rect 11366 664 11386 665
rect 11439 664 11455 665
rect 11512 664 11524 665
rect 11585 664 11593 665
rect 11658 664 11662 665
rect 11696 665 11731 698
rect 11696 664 11697 665
rect 10491 631 10529 632
rect 10563 631 10602 664
rect 10636 631 10675 664
rect 10709 631 10748 664
rect 10782 631 10821 664
rect 10855 631 10894 664
rect 10928 631 10967 664
rect 11001 631 11040 664
rect 11074 631 11113 664
rect 11147 631 11186 664
rect 11220 631 11259 664
rect 11293 631 11332 664
rect 11366 631 11405 664
rect 11439 631 11478 664
rect 11512 631 11551 664
rect 11585 631 11624 664
rect 11658 631 11697 664
rect 11765 665 11800 698
rect 11834 665 11869 698
rect 11903 665 11938 698
rect 11972 665 12007 698
rect 15373 666 15407 698
rect 15441 671 15443 700
rect 15477 671 15509 702
rect 15441 666 15509 671
rect 15373 665 15475 666
rect 11765 664 11770 665
rect 11834 664 11843 665
rect 11903 664 11915 665
rect 11972 664 11987 665
rect 11731 631 11770 664
rect 11804 631 11843 664
rect 11877 631 11915 664
rect 11949 631 11987 664
rect 15405 632 15475 665
rect 15405 631 15509 632
rect 10491 630 12007 631
rect 10491 596 10559 630
rect 10593 596 10628 630
rect 10662 596 10697 630
rect 10731 596 10766 630
rect 10800 596 10835 630
rect 10869 596 10904 630
rect 10938 596 10973 630
rect 11007 596 11042 630
rect 11076 596 11111 630
rect 11145 596 11180 630
rect 11214 596 11249 630
rect 11283 596 11318 630
rect 11352 596 11387 630
rect 11421 596 11456 630
rect 11490 596 11525 630
rect 11559 596 11594 630
rect 11628 596 11663 630
rect 11697 596 11732 630
rect 11766 596 11801 630
rect 11835 596 11870 630
rect 11904 596 11939 630
rect 10491 593 11939 596
rect 10491 562 10529 593
rect 10563 562 10602 593
rect 10636 562 10675 593
rect 10709 562 10748 593
rect 10782 562 10821 593
rect 10855 562 10894 593
rect 10928 562 10967 593
rect 11001 562 11040 593
rect 11074 562 11113 593
rect 11147 562 11186 593
rect 11220 562 11259 593
rect 11293 562 11332 593
rect 11366 562 11405 593
rect 11439 562 11478 593
rect 11512 562 11551 593
rect 11585 562 11624 593
rect 11658 562 11697 593
rect 11731 562 11770 593
rect 11804 562 11843 593
rect 11877 562 11916 593
rect 10491 528 10525 562
rect 10563 559 10594 562
rect 10636 559 10663 562
rect 10709 559 10732 562
rect 10782 559 10801 562
rect 10855 559 10870 562
rect 10928 559 10939 562
rect 11001 559 11008 562
rect 11074 559 11077 562
rect 10559 528 10594 559
rect 10628 528 10663 559
rect 10697 528 10732 559
rect 10766 528 10801 559
rect 10835 528 10870 559
rect 10904 528 10939 559
rect 10973 528 11008 559
rect 11042 528 11077 559
rect 11111 559 11113 562
rect 11180 559 11186 562
rect 11249 559 11259 562
rect 11318 559 11332 562
rect 11387 559 11405 562
rect 11456 559 11478 562
rect 11525 559 11551 562
rect 11594 559 11624 562
rect 11663 559 11697 562
rect 11111 528 11146 559
rect 11180 528 11215 559
rect 11249 528 11284 559
rect 11318 528 11353 559
rect 11387 528 11422 559
rect 11456 528 11491 559
rect 11525 528 11560 559
rect 11594 528 11629 559
rect 11663 528 11698 559
rect 11732 528 11767 562
rect 11804 559 11836 562
rect 11877 559 11905 562
rect 15373 630 15443 631
rect 15441 597 15443 630
rect 15477 597 15509 631
rect 15441 596 15509 597
rect 15407 562 15475 596
rect 11801 528 11836 559
rect 11870 528 11905 559
rect 15407 528 15509 562
rect 15661 3383 15693 3406
rect 15727 3402 15765 3406
rect 15727 3386 15797 3402
rect 15727 3382 15831 3386
rect 15727 3372 15729 3382
rect 15695 3349 15729 3372
rect 15661 3348 15729 3349
rect 15763 3363 15831 3382
rect 15763 3348 15765 3363
rect 15799 3352 15831 3363
rect 15661 3334 15765 3348
rect 15661 3314 15693 3334
rect 15727 3329 15765 3334
rect 15727 3318 15797 3329
rect 15727 3313 15831 3318
rect 15727 3300 15729 3313
rect 15695 3280 15729 3300
rect 15661 3279 15729 3280
rect 15763 3290 15831 3313
rect 15763 3279 15765 3290
rect 15799 3284 15831 3290
rect 15661 3262 15765 3279
rect 15661 3245 15693 3262
rect 15727 3256 15765 3262
rect 15727 3250 15797 3256
rect 15727 3244 15831 3250
rect 15727 3228 15729 3244
rect 15695 3211 15729 3228
rect 15661 3210 15729 3211
rect 15763 3217 15831 3244
rect 15763 3210 15765 3217
rect 15799 3216 15831 3217
rect 15661 3190 15765 3210
rect 15661 3176 15693 3190
rect 15727 3183 15765 3190
rect 15727 3182 15797 3183
rect 15727 3175 15831 3182
rect 15727 3156 15729 3175
rect 15695 3142 15729 3156
rect 15661 3141 15729 3142
rect 15763 3148 15831 3175
rect 15763 3144 15797 3148
rect 15763 3141 15765 3144
rect 15661 3118 15765 3141
rect 15661 3107 15693 3118
rect 15727 3110 15765 3118
rect 15799 3110 15831 3114
rect 15727 3106 15831 3110
rect 15727 3084 15729 3106
rect 15695 3073 15729 3084
rect 15661 3072 15729 3073
rect 15763 3080 15831 3106
rect 15763 3072 15797 3080
rect 15661 3071 15797 3072
rect 15661 3046 15765 3071
rect 15661 3038 15693 3046
rect 15727 3037 15765 3046
rect 15799 3037 15831 3046
rect 15727 3012 15729 3037
rect 15695 3004 15729 3012
rect 15661 3003 15729 3004
rect 15763 3012 15831 3037
rect 15763 3003 15797 3012
rect 15661 2998 15797 3003
rect 15661 2974 15765 2998
rect 15661 2969 15693 2974
rect 15727 2968 15765 2974
rect 15727 2940 15729 2968
rect 15695 2935 15729 2940
rect 15661 2934 15729 2935
rect 15763 2964 15765 2968
rect 15799 2964 15831 2978
rect 15763 2944 15831 2964
rect 15763 2934 15797 2944
rect 15661 2925 15797 2934
rect 15661 2902 15765 2925
rect 15661 2900 15693 2902
rect 15727 2899 15765 2902
rect 15727 2868 15729 2899
rect 15695 2866 15729 2868
rect 15661 2865 15729 2866
rect 15763 2891 15765 2899
rect 15799 2891 15831 2910
rect 15763 2876 15831 2891
rect 15763 2865 15797 2876
rect 15661 2852 15797 2865
rect 15661 2831 15765 2852
rect 15695 2830 15765 2831
rect 15661 2796 15693 2797
rect 15727 2796 15729 2830
rect 15763 2818 15765 2830
rect 15799 2818 15831 2842
rect 15763 2808 15831 2818
rect 15763 2796 15797 2808
rect 15661 2779 15797 2796
rect 15661 2762 15765 2779
rect 15695 2761 15765 2762
rect 15695 2758 15729 2761
rect 15661 2724 15693 2728
rect 15727 2727 15729 2758
rect 15763 2745 15765 2761
rect 15799 2745 15831 2774
rect 15763 2740 15831 2745
rect 15763 2727 15797 2740
rect 15727 2724 15797 2727
rect 15661 2706 15797 2724
rect 15661 2693 15765 2706
rect 15695 2692 15765 2693
rect 15695 2686 15729 2692
rect 15661 2652 15693 2659
rect 15727 2658 15729 2686
rect 15763 2672 15765 2692
rect 15799 2672 15831 2706
rect 15763 2658 15797 2672
rect 15727 2652 15797 2658
rect 15661 2638 15797 2652
rect 15661 2633 15831 2638
rect 15661 2624 15765 2633
rect 15695 2623 15765 2624
rect 15695 2614 15729 2623
rect 15661 2580 15693 2590
rect 15727 2589 15729 2614
rect 15763 2599 15765 2623
rect 15799 2604 15831 2633
rect 15763 2589 15797 2599
rect 15727 2580 15797 2589
rect 15661 2570 15797 2580
rect 15661 2560 15831 2570
rect 15661 2555 15765 2560
rect 15695 2554 15765 2555
rect 15695 2542 15729 2554
rect 15661 2508 15693 2521
rect 15727 2520 15729 2542
rect 15763 2526 15765 2554
rect 15799 2536 15831 2560
rect 15763 2520 15797 2526
rect 15727 2508 15797 2520
rect 15661 2502 15797 2508
rect 15661 2487 15831 2502
rect 15661 2486 15765 2487
rect 15695 2485 15765 2486
rect 15695 2469 15729 2485
rect 15661 2435 15693 2452
rect 15727 2451 15729 2469
rect 15763 2453 15765 2485
rect 15799 2468 15831 2487
rect 15763 2451 15797 2453
rect 15727 2435 15797 2451
rect 15661 2434 15797 2435
rect 15661 2417 15831 2434
rect 15695 2416 15831 2417
rect 15695 2396 15729 2416
rect 15661 2362 15693 2383
rect 15727 2382 15729 2396
rect 15763 2414 15831 2416
rect 15763 2382 15765 2414
rect 15799 2400 15831 2414
rect 15727 2380 15765 2382
rect 15727 2366 15797 2380
rect 15727 2362 15831 2366
rect 15661 2348 15831 2362
rect 15695 2347 15831 2348
rect 15695 2323 15729 2347
rect 15661 2289 15693 2314
rect 15727 2313 15729 2323
rect 15763 2341 15831 2347
rect 15763 2313 15765 2341
rect 15799 2331 15831 2341
rect 15727 2307 15765 2313
rect 15727 2297 15797 2307
rect 15727 2289 15831 2297
rect 15661 2279 15831 2289
rect 15695 2278 15831 2279
rect 15695 2250 15729 2278
rect 15661 2216 15693 2245
rect 15727 2244 15729 2250
rect 15763 2268 15831 2278
rect 15763 2244 15765 2268
rect 15799 2262 15831 2268
rect 15727 2234 15765 2244
rect 15727 2228 15797 2234
rect 15727 2216 15831 2228
rect 15661 2210 15831 2216
rect 15695 2209 15831 2210
rect 15695 2177 15729 2209
rect 15661 2143 15693 2176
rect 15727 2175 15729 2177
rect 15763 2195 15831 2209
rect 15763 2175 15765 2195
rect 15799 2193 15831 2195
rect 15727 2161 15765 2175
rect 15727 2159 15797 2161
rect 15727 2143 15831 2159
rect 15661 2141 15831 2143
rect 15695 2140 15831 2141
rect 15695 2107 15729 2140
rect 15661 2106 15729 2107
rect 15763 2124 15831 2140
rect 15763 2122 15797 2124
rect 15763 2106 15765 2122
rect 15661 2104 15765 2106
rect 15661 2072 15693 2104
rect 15727 2088 15765 2104
rect 15799 2088 15831 2090
rect 15727 2071 15831 2088
rect 15727 2070 15729 2071
rect 15695 2038 15729 2070
rect 15661 2037 15729 2038
rect 15763 2055 15831 2071
rect 15763 2049 15797 2055
rect 15763 2037 15765 2049
rect 15661 2031 15765 2037
rect 15661 2003 15693 2031
rect 15727 2015 15765 2031
rect 15799 2015 15831 2021
rect 15727 2002 15831 2015
rect 15727 1997 15729 2002
rect 15695 1969 15729 1997
rect 15661 1968 15729 1969
rect 15763 1986 15831 2002
rect 15763 1976 15797 1986
rect 15763 1968 15765 1976
rect 15661 1958 15765 1968
rect 15661 1934 15693 1958
rect 15727 1942 15765 1958
rect 15799 1942 15831 1952
rect 15727 1933 15831 1942
rect 15727 1924 15729 1933
rect 15695 1900 15729 1924
rect 15661 1899 15729 1900
rect 15763 1917 15831 1933
rect 15763 1903 15797 1917
rect 15763 1899 15765 1903
rect 15661 1885 15765 1899
rect 15661 1865 15693 1885
rect 15727 1869 15765 1885
rect 15799 1869 15831 1883
rect 15727 1864 15831 1869
rect 15727 1851 15729 1864
rect 15695 1831 15729 1851
rect 15661 1830 15729 1831
rect 15763 1848 15831 1864
rect 15763 1830 15797 1848
rect 15661 1812 15765 1830
rect 15661 1796 15693 1812
rect 15727 1796 15765 1812
rect 15799 1796 15831 1814
rect 15727 1795 15831 1796
rect 15727 1778 15729 1795
rect 15695 1762 15729 1778
rect 15661 1761 15729 1762
rect 15763 1779 15831 1795
rect 15763 1761 15797 1779
rect 15661 1757 15797 1761
rect 15661 1739 15765 1757
rect 15661 1727 15693 1739
rect 15727 1726 15765 1739
rect 15727 1705 15729 1726
rect 15695 1693 15729 1705
rect 15661 1692 15729 1693
rect 15763 1723 15765 1726
rect 15799 1723 15831 1745
rect 15763 1710 15831 1723
rect 15763 1692 15797 1710
rect 15661 1684 15797 1692
rect 15661 1666 15765 1684
rect 15661 1658 15693 1666
rect 15727 1657 15765 1666
rect 15727 1632 15729 1657
rect 15695 1624 15729 1632
rect 15661 1623 15729 1624
rect 15763 1650 15765 1657
rect 15799 1650 15831 1676
rect 15763 1641 15831 1650
rect 15763 1623 15797 1641
rect 15661 1610 15797 1623
rect 15661 1593 15765 1610
rect 15661 1589 15693 1593
rect 15727 1588 15765 1593
rect 15727 1559 15729 1588
rect 15695 1555 15729 1559
rect 15661 1554 15729 1555
rect 15763 1576 15765 1588
rect 15799 1576 15831 1607
rect 15763 1572 15831 1576
rect 15763 1554 15797 1572
rect 15661 1538 15797 1554
rect 15661 1536 15831 1538
rect 15661 1520 15765 1536
rect 15727 1519 15765 1520
rect 15727 1486 15729 1519
rect 15661 1485 15729 1486
rect 15763 1502 15765 1519
rect 15799 1503 15831 1536
rect 15763 1485 15797 1502
rect 15661 1469 15797 1485
rect 15661 1462 15831 1469
rect 15661 1450 15765 1462
rect 15695 1447 15729 1450
rect 15727 1416 15729 1447
rect 15763 1428 15765 1450
rect 15799 1434 15831 1462
rect 15763 1416 15797 1428
rect 15661 1413 15693 1416
rect 15727 1413 15797 1416
rect 15661 1400 15797 1413
rect 15661 1388 15831 1400
rect 15661 1380 15765 1388
rect 15695 1374 15729 1380
rect 15727 1346 15729 1374
rect 15763 1354 15765 1380
rect 15799 1365 15831 1388
rect 15763 1346 15797 1354
rect 15661 1340 15693 1346
rect 15727 1340 15797 1346
rect 15661 1331 15797 1340
rect 15661 1314 15831 1331
rect 15661 1310 15765 1314
rect 15695 1301 15729 1310
rect 15727 1276 15729 1301
rect 15763 1280 15765 1310
rect 15799 1296 15831 1314
rect 15763 1276 15797 1280
rect 15661 1267 15693 1276
rect 15727 1267 15797 1276
rect 15661 1262 15797 1267
rect 15661 1240 15831 1262
rect 15695 1228 15729 1240
rect 15727 1206 15729 1228
rect 15763 1206 15765 1240
rect 15799 1227 15831 1240
rect 15661 1194 15693 1206
rect 15727 1194 15797 1206
rect 15661 1193 15797 1194
rect 15661 1170 15831 1193
rect 15695 1155 15729 1170
rect 15727 1136 15729 1155
rect 15763 1166 15831 1170
rect 15763 1136 15765 1166
rect 15799 1158 15831 1166
rect 15661 1121 15693 1136
rect 15727 1132 15765 1136
rect 15727 1124 15797 1132
rect 15727 1121 15831 1124
rect 15661 1100 15831 1121
rect 15695 1082 15729 1100
rect 15727 1066 15729 1082
rect 15763 1092 15831 1100
rect 15763 1066 15765 1092
rect 15799 1089 15831 1092
rect 15661 1048 15693 1066
rect 15727 1058 15765 1066
rect 15727 1055 15797 1058
rect 15727 1048 15831 1055
rect 15661 1030 15831 1048
rect 15695 1009 15729 1030
rect 15727 996 15729 1009
rect 15763 1020 15831 1030
rect 15763 1018 15797 1020
rect 15763 996 15765 1018
rect 15661 975 15693 996
rect 15727 984 15765 996
rect 15799 984 15831 986
rect 15727 975 15831 984
rect 15661 960 15831 975
rect 15695 936 15729 960
rect 15727 926 15729 936
rect 15763 951 15831 960
rect 15763 944 15797 951
rect 15763 926 15765 944
rect 15661 902 15693 926
rect 15727 910 15765 926
rect 15799 910 15831 917
rect 15727 902 15831 910
rect 15661 890 15831 902
rect 15695 863 15729 890
rect 15727 856 15729 863
rect 15763 882 15831 890
rect 15763 870 15797 882
rect 15763 856 15765 870
rect 15661 829 15693 856
rect 15727 836 15765 856
rect 15799 836 15831 848
rect 15727 829 15831 836
rect 15661 820 15831 829
rect 15695 790 15729 820
rect 15727 786 15729 790
rect 15763 813 15831 820
rect 15763 796 15797 813
rect 15763 786 15765 796
rect 15661 756 15693 786
rect 15727 762 15765 786
rect 15799 762 15831 779
rect 15727 756 15831 762
rect 15661 750 15831 756
rect 15695 717 15729 750
rect 15727 716 15729 717
rect 15763 744 15831 750
rect 15763 722 15797 744
rect 15763 716 15765 722
rect 15661 683 15693 716
rect 15727 688 15765 716
rect 15799 688 15831 710
rect 15727 683 15831 688
rect 15661 680 15831 683
rect 15695 646 15729 680
rect 15763 675 15831 680
rect 15763 648 15797 675
rect 15763 646 15765 648
rect 15661 644 15765 646
rect 15661 610 15693 644
rect 15727 614 15765 644
rect 15799 614 15831 641
rect 15727 610 15831 614
rect 15695 576 15729 610
rect 15763 606 15831 610
rect 15763 576 15797 606
rect 15661 574 15797 576
rect 15661 571 15765 574
rect 15661 540 15693 571
rect 15727 540 15765 571
rect 15799 540 15831 572
rect 15727 537 15729 540
rect 15695 506 15729 537
rect 15763 537 15831 540
rect 15763 506 15797 537
rect 15661 503 15797 506
rect 15661 500 15831 503
rect 15661 498 15765 500
rect 15661 470 15693 498
rect 15727 470 15765 498
rect 15727 464 15729 470
rect 15695 436 15729 464
rect 15763 466 15765 470
rect 15799 468 15831 500
rect 15763 436 15797 466
rect 15661 434 15797 436
rect 15661 426 15831 434
rect 15661 425 15765 426
rect 10809 399 10915 415
rect 10845 365 10881 399
rect 10809 349 10915 365
rect 12951 399 13057 415
rect 12985 365 13021 399
rect 12951 349 13057 365
rect 15661 400 15693 425
rect 15727 400 15765 425
rect 15727 391 15729 400
rect 15695 366 15729 391
rect 15763 392 15765 400
rect 15799 399 15831 426
rect 15763 366 15797 392
rect 15661 365 15797 366
rect 15661 352 15831 365
rect 15661 330 15693 352
rect 15727 330 15765 352
rect 15799 330 15831 352
rect 15727 318 15729 330
rect 15695 296 15729 318
rect 15763 318 15765 330
rect 15763 296 15797 318
rect 15661 236 15831 296
rect 10135 66 15831 236
<< viali >>
rect 393 17391 425 17425
rect 425 17391 427 17425
rect 466 17391 500 17425
rect 539 17391 573 17425
rect 612 17391 646 17425
rect 685 17391 719 17425
rect 758 17391 792 17425
rect 831 17391 865 17425
rect 904 17391 938 17425
rect 977 17391 1011 17425
rect 1050 17391 1084 17425
rect 1123 17391 1157 17425
rect 1196 17391 1230 17425
rect 1269 17391 1303 17425
rect 1342 17391 1376 17425
rect 1415 17391 1449 17425
rect 1488 17391 1522 17425
rect 1561 17391 1595 17425
rect 1634 17391 1668 17425
rect 1707 17391 1741 17425
rect 1780 17391 1814 17425
rect 1853 17391 1887 17425
rect 1926 17391 1960 17425
rect 1999 17391 2033 17425
rect 2072 17391 2106 17425
rect 2145 17391 2179 17425
rect 2218 17391 2252 17425
rect 2291 17391 2325 17425
rect 2364 17391 2398 17425
rect 2437 17391 2471 17425
rect 2510 17391 2544 17425
rect 2583 17391 2617 17425
rect 2656 17391 2690 17425
rect 2729 17391 2763 17425
rect 2802 17391 2836 17425
rect 2875 17391 2909 17425
rect 2948 17391 2982 17425
rect 3021 17391 3055 17425
rect 3094 17391 3128 17425
rect 3167 17391 3201 17425
rect 3240 17391 3274 17425
rect 3313 17391 3347 17425
rect 3386 17391 3420 17425
rect 3459 17391 3493 17425
rect 3532 17391 3566 17425
rect 3605 17391 3639 17425
rect 3678 17391 3712 17425
rect 3751 17391 3785 17425
rect 3824 17391 3858 17425
rect 3897 17391 3931 17425
rect 3970 17391 4004 17425
rect 4043 17391 4077 17425
rect 4116 17391 4150 17425
rect 4189 17391 4223 17425
rect 4262 17391 4296 17425
rect 4335 17391 4369 17425
rect 4408 17391 4442 17425
rect 4481 17391 4515 17425
rect 4554 17391 4588 17425
rect 4627 17391 4661 17425
rect 4700 17391 4734 17425
rect 4773 17423 16167 17425
rect 16167 17423 16202 17425
rect 16202 17423 16236 17425
rect 16236 17423 16271 17425
rect 16271 17423 16305 17425
rect 16305 17423 16340 17425
rect 16340 17423 16374 17425
rect 16374 17423 16409 17425
rect 16409 17423 16443 17425
rect 16443 17423 16478 17425
rect 16478 17423 16512 17425
rect 16512 17423 16543 17425
rect 16963 17423 16995 17425
rect 16995 17423 16997 17425
rect 17037 17423 17064 17425
rect 17064 17423 17071 17425
rect 17111 17423 17133 17425
rect 17133 17423 17145 17425
rect 17185 17423 17202 17425
rect 17202 17423 17219 17425
rect 17259 17423 17271 17425
rect 17271 17423 17293 17425
rect 17333 17423 17340 17425
rect 17340 17423 17367 17425
rect 17407 17423 17409 17425
rect 17409 17423 17441 17425
rect 17481 17423 17513 17425
rect 17513 17423 17515 17425
rect 17555 17423 17582 17425
rect 17582 17423 17589 17425
rect 17630 17423 17651 17425
rect 17651 17423 17664 17425
rect 17705 17423 17720 17425
rect 17720 17423 17739 17425
rect 17780 17423 17789 17425
rect 17789 17423 17814 17425
rect 17855 17423 17858 17425
rect 17858 17423 17889 17425
rect 17930 17423 17961 17425
rect 17961 17423 17964 17425
rect 18005 17423 18030 17425
rect 18030 17423 18039 17425
rect 18080 17423 18099 17425
rect 18099 17423 18114 17425
rect 18155 17423 18168 17425
rect 18168 17423 18189 17425
rect 18230 17423 18237 17425
rect 18237 17423 18264 17425
rect 18305 17423 18306 17425
rect 18306 17423 18339 17425
rect 4773 17355 16133 17423
rect 16133 17389 16543 17423
rect 16963 17391 16997 17423
rect 17037 17391 17071 17423
rect 17111 17391 17145 17423
rect 17185 17391 17219 17423
rect 17259 17391 17293 17423
rect 17333 17391 17367 17423
rect 17407 17391 17441 17423
rect 17481 17391 17515 17423
rect 17555 17391 17589 17423
rect 17630 17391 17664 17423
rect 17705 17391 17739 17423
rect 17780 17391 17814 17423
rect 17855 17391 17889 17423
rect 17930 17391 17964 17423
rect 18005 17391 18039 17423
rect 18080 17391 18114 17423
rect 18155 17391 18189 17423
rect 18230 17391 18264 17423
rect 18305 17391 18339 17423
rect 16133 17355 16168 17389
rect 16168 17355 16202 17389
rect 16202 17355 16237 17389
rect 16237 17355 16271 17389
rect 16271 17355 16306 17389
rect 16306 17355 16340 17389
rect 16340 17355 16375 17389
rect 16375 17355 16409 17389
rect 16409 17355 16444 17389
rect 16444 17355 16478 17389
rect 16478 17355 16513 17389
rect 16513 17355 16543 17389
rect 355 17285 389 17309
rect 427 17319 459 17353
rect 459 17319 461 17353
rect 500 17319 534 17353
rect 573 17319 607 17353
rect 646 17319 680 17353
rect 719 17319 753 17353
rect 792 17319 826 17353
rect 865 17319 899 17353
rect 938 17319 972 17353
rect 1011 17319 1045 17353
rect 1084 17319 1118 17353
rect 1157 17319 1191 17353
rect 1230 17319 1264 17353
rect 1303 17319 1337 17353
rect 1376 17319 1410 17353
rect 1449 17319 1483 17353
rect 1522 17319 1556 17353
rect 1595 17319 1629 17353
rect 1668 17319 1702 17353
rect 1741 17319 1775 17353
rect 1814 17319 1848 17353
rect 1887 17319 1921 17353
rect 1960 17319 1994 17353
rect 2033 17319 2067 17353
rect 2106 17319 2140 17353
rect 2179 17319 2213 17353
rect 2252 17319 2286 17353
rect 2325 17319 2359 17353
rect 2397 17319 2431 17353
rect 2469 17319 2503 17353
rect 2541 17319 2575 17353
rect 2613 17319 2647 17353
rect 2685 17319 2719 17353
rect 2757 17319 2791 17353
rect 2829 17319 2863 17353
rect 2901 17319 2935 17353
rect 2973 17319 3007 17353
rect 3045 17319 3079 17353
rect 3117 17319 3151 17353
rect 3189 17319 3223 17353
rect 3261 17319 3295 17353
rect 3333 17319 3367 17353
rect 3405 17319 3439 17353
rect 3477 17319 3511 17353
rect 3549 17319 3583 17353
rect 3621 17319 3655 17353
rect 3693 17319 3727 17353
rect 3765 17319 3799 17353
rect 3837 17319 3871 17353
rect 3909 17319 3943 17353
rect 3981 17319 4015 17353
rect 4053 17319 4087 17353
rect 4125 17319 4159 17353
rect 4197 17319 4231 17353
rect 4269 17319 4303 17353
rect 4341 17319 4375 17353
rect 4413 17319 4447 17353
rect 4485 17319 4519 17353
rect 4557 17319 4591 17353
rect 4629 17319 4663 17353
rect 4701 17319 4735 17353
rect 4773 17319 16065 17355
rect 16065 17321 16543 17355
rect 16065 17319 16100 17321
rect 16100 17319 16134 17321
rect 16134 17319 16169 17321
rect 16169 17319 16203 17321
rect 16203 17319 16238 17321
rect 16238 17319 16272 17321
rect 16272 17319 16307 17321
rect 16307 17319 16341 17321
rect 16341 17319 16376 17321
rect 16376 17319 16410 17321
rect 16410 17319 16445 17321
rect 16445 17319 16479 17321
rect 16479 17319 16514 17321
rect 16514 17319 16543 17321
rect 16963 17319 16997 17353
rect 17035 17321 17069 17353
rect 17107 17321 17141 17353
rect 17179 17321 17213 17353
rect 17251 17321 17285 17353
rect 17323 17321 17357 17353
rect 17395 17321 17429 17353
rect 17468 17321 17502 17353
rect 17541 17321 17575 17353
rect 17614 17321 17648 17353
rect 17687 17321 17721 17353
rect 17760 17321 17794 17353
rect 17833 17321 17867 17353
rect 17906 17321 17940 17353
rect 17979 17321 18013 17353
rect 18052 17321 18086 17353
rect 18125 17321 18159 17353
rect 18198 17321 18232 17353
rect 18271 17321 18305 17353
rect 17035 17319 17066 17321
rect 17066 17319 17069 17321
rect 17107 17319 17135 17321
rect 17135 17319 17141 17321
rect 17179 17319 17204 17321
rect 17204 17319 17213 17321
rect 17251 17319 17273 17321
rect 17273 17319 17285 17321
rect 17323 17319 17342 17321
rect 17342 17319 17357 17321
rect 17395 17319 17411 17321
rect 17411 17319 17429 17321
rect 17468 17319 17480 17321
rect 17480 17319 17502 17321
rect 17541 17319 17549 17321
rect 17549 17319 17575 17321
rect 17614 17319 17618 17321
rect 17618 17319 17648 17321
rect 17687 17319 17721 17321
rect 17760 17319 17790 17321
rect 17790 17319 17794 17321
rect 17833 17319 17859 17321
rect 17859 17319 17867 17321
rect 17906 17319 17928 17321
rect 17928 17319 17940 17321
rect 17979 17319 17997 17321
rect 17997 17319 18013 17321
rect 18052 17319 18066 17321
rect 18066 17319 18086 17321
rect 18125 17319 18135 17321
rect 18135 17319 18159 17321
rect 18198 17319 18204 17321
rect 18204 17319 18232 17321
rect 18271 17319 18305 17321
rect 355 17275 357 17285
rect 357 17275 389 17285
rect 427 17252 461 17280
rect 355 17216 389 17234
rect 427 17246 459 17252
rect 459 17246 461 17252
rect 355 17200 357 17216
rect 357 17200 389 17216
rect 427 17183 461 17207
rect 355 17147 389 17158
rect 427 17173 459 17183
rect 459 17173 461 17183
rect 355 17124 357 17147
rect 357 17124 389 17147
rect 716 17134 750 17140
rect 789 17134 823 17140
rect 862 17134 896 17140
rect 935 17134 969 17140
rect 1008 17134 1042 17140
rect 1081 17134 1115 17140
rect 1154 17134 1188 17140
rect 1227 17134 1261 17140
rect 1300 17134 1334 17140
rect 1373 17134 1407 17140
rect 1446 17134 1480 17140
rect 1519 17134 1553 17140
rect 1592 17134 1626 17140
rect 1665 17134 1699 17140
rect 1738 17134 1772 17140
rect 1811 17134 1845 17140
rect 1884 17134 1918 17140
rect 1957 17134 1991 17140
rect 2030 17134 2064 17140
rect 2103 17134 2137 17140
rect 2176 17134 2210 17140
rect 2249 17134 2283 17140
rect 2322 17134 2356 17140
rect 2395 17134 2429 17140
rect 2468 17134 2502 17140
rect 2541 17134 2575 17140
rect 2614 17134 2648 17140
rect 2687 17134 2721 17140
rect 2760 17134 2794 17140
rect 2833 17134 2867 17140
rect 2906 17134 2940 17140
rect 2979 17134 3013 17140
rect 3052 17134 3086 17140
rect 3125 17134 3159 17140
rect 3197 17134 3231 17140
rect 3269 17134 3303 17140
rect 3341 17134 3375 17140
rect 3413 17134 3447 17140
rect 3485 17134 3519 17140
rect 3557 17134 3591 17140
rect 3629 17134 3663 17140
rect 3701 17134 3735 17140
rect 3773 17134 3807 17140
rect 3845 17134 3879 17140
rect 3917 17134 3951 17140
rect 3989 17134 4023 17140
rect 4061 17134 4095 17140
rect 4133 17134 4167 17140
rect 4205 17134 4239 17140
rect 4277 17134 4311 17140
rect 4349 17134 4383 17140
rect 4421 17134 4455 17140
rect 4493 17134 4527 17140
rect 4565 17134 4599 17140
rect 4637 17134 4671 17140
rect 4709 17134 4743 17140
rect 4781 17134 4815 17140
rect 4853 17134 4887 17140
rect 4925 17134 4959 17140
rect 4997 17134 5031 17140
rect 5069 17134 5103 17140
rect 5141 17134 5175 17140
rect 5213 17134 5247 17140
rect 5285 17134 5319 17140
rect 5357 17134 5391 17140
rect 5429 17134 5463 17140
rect 5501 17134 5535 17140
rect 5573 17134 5607 17140
rect 5645 17134 5679 17140
rect 5717 17134 5751 17140
rect 5789 17134 5823 17140
rect 5861 17134 5895 17140
rect 5933 17134 16407 17140
rect 427 17114 461 17134
rect 355 17078 389 17082
rect 427 17100 459 17114
rect 459 17100 461 17114
rect 355 17048 357 17078
rect 357 17048 389 17078
rect 427 17045 461 17061
rect 427 17027 459 17045
rect 459 17027 461 17045
rect 355 16975 357 17006
rect 357 16975 389 17006
rect 427 16976 461 16988
rect 355 16972 389 16975
rect 427 16954 459 16976
rect 459 16954 461 16976
rect 355 16906 357 16930
rect 357 16906 389 16930
rect 427 16907 461 16915
rect 355 16896 389 16906
rect 427 16881 459 16907
rect 459 16881 461 16907
rect 355 16837 357 16854
rect 357 16837 389 16854
rect 427 16838 461 16842
rect 355 16820 389 16837
rect 427 16808 459 16838
rect 459 16808 461 16838
rect 355 16768 357 16778
rect 357 16768 389 16778
rect 355 16744 389 16768
rect 427 16735 461 16769
rect 355 16699 357 16702
rect 357 16699 389 16702
rect 355 16668 389 16699
rect 427 16662 461 16696
rect 355 16595 389 16626
rect 355 16592 357 16595
rect 357 16592 389 16595
rect 427 16588 461 16622
rect 355 16526 389 16550
rect 355 16516 357 16526
rect 357 16516 389 16526
rect 427 16514 461 16548
rect 355 16457 389 16474
rect 355 16440 357 16457
rect 357 16440 389 16457
rect 427 16440 461 16474
rect 357 15813 391 15847
rect 429 15813 463 15847
rect 357 15739 391 15773
rect 429 15739 463 15773
rect 357 15665 391 15699
rect 429 15665 463 15699
rect 357 15591 391 15625
rect 429 15591 463 15625
rect 357 15517 391 15551
rect 429 15517 463 15551
rect 357 15443 391 15477
rect 429 15443 463 15477
rect 357 15369 391 15403
rect 429 15369 463 15403
rect 357 15295 391 15329
rect 429 15295 463 15329
rect 357 15221 391 15255
rect 429 15221 463 15255
rect 357 15147 391 15181
rect 429 15147 463 15181
rect 357 15073 391 15107
rect 429 15073 463 15107
rect 357 14999 391 15033
rect 429 14999 463 15033
rect 357 14925 391 14959
rect 429 14925 463 14959
rect 357 14851 391 14885
rect 429 14851 463 14885
rect 357 14777 391 14811
rect 429 14777 463 14811
rect 357 14703 391 14737
rect 429 14703 463 14737
rect 357 14629 391 14663
rect 429 14629 463 14663
rect 357 14555 391 14589
rect 429 14555 463 14589
rect 357 14481 391 14515
rect 429 14481 463 14515
rect 357 14407 391 14441
rect 429 14407 463 14441
rect 357 14333 391 14367
rect 429 14333 463 14367
rect 357 14259 391 14293
rect 429 14259 463 14293
rect 357 14185 391 14219
rect 429 14185 463 14219
rect 357 14111 391 14145
rect 429 14111 463 14145
rect 357 14037 391 14071
rect 429 14037 463 14071
rect 357 13963 391 13997
rect 429 13963 463 13997
rect 357 13889 391 13923
rect 429 13889 463 13923
rect 357 13816 391 13850
rect 429 13845 459 13850
rect 459 13845 463 13850
rect 429 13816 463 13845
rect 357 13743 391 13777
rect 429 13776 459 13777
rect 459 13776 463 13777
rect 429 13743 463 13776
rect 357 13670 391 13704
rect 429 13672 463 13704
rect 429 13670 463 13672
rect 357 13597 391 13631
rect 429 13597 463 13631
rect 357 13524 391 13558
rect 429 13524 463 13558
rect 357 13451 391 13485
rect 429 13451 463 13485
rect 357 13378 391 13412
rect 429 13378 463 13412
rect 357 13305 391 13339
rect 429 13305 463 13339
rect 357 13232 391 13266
rect 429 13232 463 13266
rect 357 13159 391 13193
rect 429 13159 463 13193
rect 357 13086 391 13120
rect 429 13086 463 13120
rect 357 13013 391 13047
rect 429 13013 463 13047
rect 357 12940 391 12974
rect 429 12940 463 12974
rect 357 12867 391 12901
rect 429 12867 463 12901
rect 357 12794 391 12828
rect 429 12794 463 12828
rect 716 17106 748 17134
rect 748 17106 750 17134
rect 789 17106 823 17134
rect 862 17106 896 17134
rect 935 17106 969 17134
rect 1008 17106 1042 17134
rect 1081 17106 1115 17134
rect 1154 17106 1188 17134
rect 1227 17106 1261 17134
rect 1300 17106 1334 17134
rect 1373 17106 1407 17134
rect 1446 17106 1480 17134
rect 1519 17106 1553 17134
rect 1592 17106 1626 17134
rect 1665 17106 1699 17134
rect 1738 17106 1772 17134
rect 1811 17106 1845 17134
rect 1884 17106 1918 17134
rect 1957 17106 1991 17134
rect 2030 17106 2064 17134
rect 2103 17106 2137 17134
rect 2176 17106 2210 17134
rect 2249 17106 2283 17134
rect 2322 17106 2356 17134
rect 2395 17106 2429 17134
rect 2468 17106 2502 17134
rect 2541 17106 2575 17134
rect 2614 17106 2648 17134
rect 2687 17106 2721 17134
rect 2760 17106 2794 17134
rect 2833 17106 2867 17134
rect 2906 17106 2940 17134
rect 2979 17106 3013 17134
rect 3052 17106 3086 17134
rect 3125 17106 3159 17134
rect 3197 17106 3231 17134
rect 3269 17106 3303 17134
rect 3341 17106 3375 17134
rect 3413 17106 3447 17134
rect 3485 17106 3519 17134
rect 3557 17106 3591 17134
rect 3629 17106 3663 17134
rect 3701 17106 3735 17134
rect 3773 17106 3807 17134
rect 3845 17106 3879 17134
rect 3917 17106 3951 17134
rect 3989 17106 4023 17134
rect 4061 17106 4095 17134
rect 4133 17106 4167 17134
rect 4205 17106 4239 17134
rect 4277 17106 4311 17134
rect 4349 17106 4383 17134
rect 4421 17106 4455 17134
rect 4493 17106 4527 17134
rect 4565 17106 4599 17134
rect 4637 17106 4671 17134
rect 4709 17106 4743 17134
rect 4781 17106 4815 17134
rect 4853 17106 4887 17134
rect 4925 17106 4959 17134
rect 4997 17106 5031 17134
rect 5069 17106 5103 17134
rect 5141 17106 5175 17134
rect 5213 17106 5247 17134
rect 5285 17106 5319 17134
rect 5357 17106 5391 17134
rect 5429 17106 5463 17134
rect 5501 17106 5535 17134
rect 5573 17106 5607 17134
rect 5645 17106 5679 17134
rect 5717 17106 5751 17134
rect 5789 17106 5823 17134
rect 5861 17106 5895 17134
rect 5933 17100 13498 17134
rect 13498 17100 13533 17134
rect 13533 17100 13567 17134
rect 13567 17100 13602 17134
rect 13602 17100 13636 17134
rect 13636 17100 13671 17134
rect 13671 17100 13705 17134
rect 13705 17100 13740 17134
rect 13740 17100 13774 17134
rect 13774 17100 13809 17134
rect 13809 17100 13843 17134
rect 13843 17100 13878 17134
rect 13878 17100 13912 17134
rect 13912 17100 13947 17134
rect 13947 17100 13981 17134
rect 13981 17100 14016 17134
rect 14016 17100 14050 17134
rect 14050 17100 14085 17134
rect 14085 17100 14119 17134
rect 14119 17100 14154 17134
rect 14154 17100 14188 17134
rect 14188 17100 14223 17134
rect 14223 17100 14257 17134
rect 14257 17100 14292 17134
rect 14292 17100 14326 17134
rect 14326 17100 14361 17134
rect 14361 17100 14395 17134
rect 14395 17100 14430 17134
rect 14430 17100 14464 17134
rect 14464 17100 14499 17134
rect 14499 17100 14533 17134
rect 14533 17100 14568 17134
rect 14568 17100 14602 17134
rect 14602 17100 14637 17134
rect 14637 17100 14671 17134
rect 14671 17100 14706 17134
rect 14706 17100 14740 17134
rect 14740 17100 14775 17134
rect 14775 17100 14809 17134
rect 14809 17100 14844 17134
rect 14844 17100 14878 17134
rect 14878 17100 14913 17134
rect 14913 17100 14947 17134
rect 14947 17100 14982 17134
rect 14982 17100 15016 17134
rect 15016 17100 15051 17134
rect 15051 17100 15085 17134
rect 15085 17100 15120 17134
rect 15120 17100 15154 17134
rect 15154 17100 15189 17134
rect 15189 17100 15223 17134
rect 15223 17100 15258 17134
rect 15258 17100 15292 17134
rect 15292 17100 15327 17134
rect 15327 17100 15361 17134
rect 15361 17100 15396 17134
rect 15396 17100 15430 17134
rect 15430 17100 15465 17134
rect 15465 17100 15499 17134
rect 15499 17100 15534 17134
rect 15534 17100 15568 17134
rect 15568 17100 15603 17134
rect 15603 17100 15637 17134
rect 15637 17100 15672 17134
rect 15672 17100 15706 17134
rect 15706 17100 15741 17134
rect 15741 17100 15775 17134
rect 15775 17100 15810 17134
rect 15810 17100 15844 17134
rect 15844 17100 15879 17134
rect 15879 17100 15913 17134
rect 15913 17100 15948 17134
rect 15948 17100 15982 17134
rect 15982 17100 16017 17134
rect 16017 17100 16051 17134
rect 16051 17100 16086 17134
rect 16086 17100 16120 17134
rect 16120 17100 16155 17134
rect 16155 17100 16189 17134
rect 16189 17100 16224 17134
rect 16224 17100 16258 17134
rect 16258 17100 16293 17134
rect 16293 17100 16327 17134
rect 16327 17100 16362 17134
rect 16362 17100 16396 17134
rect 16396 17100 16407 17134
rect 17146 17100 17155 17102
rect 17155 17100 17180 17102
rect 17222 17100 17224 17102
rect 17224 17100 17256 17102
rect 17298 17100 17328 17102
rect 17328 17100 17332 17102
rect 17374 17100 17397 17102
rect 17397 17100 17408 17102
rect 17450 17100 17466 17102
rect 17466 17100 17484 17102
rect 17526 17100 17535 17102
rect 17535 17100 17560 17102
rect 17602 17100 17604 17102
rect 17604 17100 17636 17102
rect 17678 17100 17707 17102
rect 17707 17100 17712 17102
rect 17754 17100 17776 17102
rect 17776 17100 17788 17102
rect 17830 17100 17845 17102
rect 17845 17100 17864 17102
rect 17906 17100 17914 17102
rect 17914 17100 17940 17102
rect 17982 17100 17983 17102
rect 17983 17100 18016 17102
rect 750 17034 784 17068
rect 823 17034 857 17068
rect 896 17034 930 17068
rect 969 17034 1003 17068
rect 1042 17034 1076 17068
rect 1115 17034 1149 17068
rect 1188 17034 1222 17068
rect 1261 17034 1295 17068
rect 1334 17034 1368 17068
rect 1407 17034 1441 17068
rect 1480 17034 1514 17068
rect 1553 17034 1587 17068
rect 1626 17034 1660 17068
rect 1699 17034 1733 17068
rect 1772 17034 1806 17068
rect 1845 17034 1879 17068
rect 1918 17034 1952 17068
rect 1991 17034 2025 17068
rect 2064 17034 2098 17068
rect 2137 17034 2171 17068
rect 2210 17034 2244 17068
rect 2283 17034 2317 17068
rect 2356 17034 2390 17068
rect 2429 17034 2463 17068
rect 2502 17034 2536 17068
rect 2575 17034 2609 17068
rect 2648 17034 2682 17068
rect 2721 17034 2755 17068
rect 2794 17034 2828 17068
rect 2867 17034 2901 17068
rect 2940 17034 2974 17068
rect 3013 17034 3047 17068
rect 3086 17034 3120 17068
rect 3159 17034 3193 17068
rect 3232 17034 3266 17068
rect 3305 17034 3339 17068
rect 3378 17034 3412 17068
rect 3451 17034 3485 17068
rect 3524 17034 3558 17068
rect 3597 17034 3631 17068
rect 3670 17034 3704 17068
rect 3743 17034 3777 17068
rect 3816 17034 3850 17068
rect 3889 17034 3923 17068
rect 3962 17034 3996 17068
rect 4035 17034 4069 17068
rect 4108 17034 4142 17068
rect 4181 17034 4215 17068
rect 4254 17034 4288 17068
rect 4327 17034 4361 17068
rect 4400 17034 4434 17068
rect 4473 17034 4507 17068
rect 4546 17034 4580 17068
rect 4619 17034 4653 17068
rect 4692 17034 4726 17068
rect 4765 17034 4799 17068
rect 4838 17034 4872 17068
rect 4911 17034 4945 17068
rect 4984 17034 5018 17068
rect 5057 17034 5091 17068
rect 5130 17034 5164 17068
rect 5203 17034 5237 17068
rect 5276 17034 5310 17068
rect 5349 17034 5383 17068
rect 5422 17034 5456 17068
rect 5495 17034 5529 17068
rect 5568 17034 5602 17068
rect 5641 17034 5675 17068
rect 5714 17034 5748 17068
rect 5787 17034 5821 17068
rect 5860 17034 5894 17068
rect 5933 17034 13464 17100
rect 13464 17066 16407 17100
rect 17146 17068 17180 17100
rect 17222 17068 17256 17100
rect 17298 17068 17332 17100
rect 17374 17068 17408 17100
rect 17450 17068 17484 17100
rect 17526 17068 17560 17100
rect 17602 17068 17636 17100
rect 17678 17068 17712 17100
rect 17754 17068 17788 17100
rect 17830 17068 17864 17100
rect 17906 17068 17940 17100
rect 17982 17068 18016 17100
rect 13464 17034 13499 17066
rect 13499 17034 13533 17066
rect 13533 17034 13568 17066
rect 13568 17034 13602 17066
rect 13602 17034 13637 17066
rect 13637 17034 13671 17066
rect 13671 17034 13706 17066
rect 13706 17034 13740 17066
rect 13740 17034 13775 17066
rect 13775 17034 13809 17066
rect 13809 17034 13844 17066
rect 13844 17034 13878 17066
rect 13878 17034 13913 17066
rect 13913 17034 13947 17066
rect 13947 17034 13982 17066
rect 13982 17034 14016 17066
rect 14016 17034 14051 17066
rect 14051 17034 14085 17066
rect 14085 17034 14120 17066
rect 14120 17034 14154 17066
rect 14154 17034 14189 17066
rect 14189 17034 14223 17066
rect 14223 17034 14258 17066
rect 14258 17034 14292 17066
rect 14292 17034 14327 17066
rect 14327 17034 14361 17066
rect 14361 17034 14396 17066
rect 14396 17034 14430 17066
rect 14430 17034 14465 17066
rect 14465 17034 14499 17066
rect 14499 17034 14534 17066
rect 14534 17034 14568 17066
rect 14568 17034 14603 17066
rect 14603 17034 14637 17066
rect 14637 17034 14672 17066
rect 14672 17034 14706 17066
rect 14706 17034 14741 17066
rect 14741 17034 14775 17066
rect 14775 17034 14810 17066
rect 14810 17034 14844 17066
rect 14844 17034 14879 17066
rect 14879 17034 14913 17066
rect 14913 17034 14948 17066
rect 14948 17034 14982 17066
rect 14982 17034 15017 17066
rect 15017 17034 15051 17066
rect 15051 17034 15086 17066
rect 15086 17034 15120 17066
rect 15120 17034 15155 17066
rect 15155 17034 15189 17066
rect 15189 17034 15224 17066
rect 15224 17034 15258 17066
rect 15258 17034 15293 17066
rect 15293 17034 15327 17066
rect 15327 17034 15362 17066
rect 15362 17034 15396 17066
rect 15396 17034 15431 17066
rect 15431 17034 15465 17066
rect 15465 17034 15500 17066
rect 15500 17034 15534 17066
rect 15534 17034 15569 17066
rect 15569 17034 15603 17066
rect 15603 17034 15638 17066
rect 15638 17034 15672 17066
rect 15672 17034 15707 17066
rect 15707 17034 15741 17066
rect 15741 17034 15776 17066
rect 15776 17034 15810 17066
rect 15810 17034 15845 17066
rect 15845 17034 15879 17066
rect 15879 17034 15914 17066
rect 15914 17034 15948 17066
rect 15948 17034 15983 17066
rect 15983 17034 16017 17066
rect 16017 17034 16052 17066
rect 16052 17034 16086 17066
rect 16086 17034 16121 17066
rect 16121 17034 16155 17066
rect 16155 17034 16190 17066
rect 16190 17034 16224 17066
rect 16224 17034 16259 17066
rect 16259 17034 16293 17066
rect 16293 17034 16328 17066
rect 16328 17034 16362 17066
rect 16362 17034 16397 17066
rect 16397 17034 16407 17066
rect 678 16997 680 17028
rect 680 16997 712 17028
rect 678 16994 712 16997
rect 750 16964 782 16988
rect 782 16964 784 16988
rect 3267 16964 3301 16996
rect 3339 16964 3373 16996
rect 5609 16964 5643 16996
rect 5681 16964 5715 16996
rect 7951 16964 8057 17034
rect 10293 16964 10399 17034
rect 17146 16998 17180 17030
rect 17218 16998 17252 17030
rect 17291 16998 17325 17030
rect 17364 16998 17398 17030
rect 17437 16998 17471 17030
rect 17510 16998 17544 17030
rect 17583 16998 17617 17030
rect 17656 16998 17690 17030
rect 17729 16998 17763 17030
rect 17802 16998 17836 17030
rect 17875 16998 17909 17030
rect 17948 16998 17982 17030
rect 10476 16964 10510 16973
rect 10549 16964 10583 16973
rect 10622 16964 10656 16973
rect 10695 16964 10729 16973
rect 10768 16964 10802 16973
rect 10841 16964 10875 16973
rect 10914 16964 10948 16973
rect 10987 16964 11021 16973
rect 11060 16964 11094 16973
rect 11133 16964 13396 16973
rect 13396 16964 13431 16973
rect 13431 16964 13465 16973
rect 13465 16964 13500 16973
rect 13500 16964 13534 16973
rect 13534 16964 13569 16973
rect 13569 16964 13603 16973
rect 13603 16964 13638 16973
rect 13638 16964 13672 16973
rect 13672 16964 13707 16973
rect 13707 16964 13741 16973
rect 13741 16964 13776 16973
rect 13776 16964 13810 16973
rect 13810 16964 13845 16973
rect 13845 16964 13879 16973
rect 13879 16964 13914 16973
rect 13914 16964 13948 16973
rect 13948 16964 13983 16973
rect 13983 16964 14017 16973
rect 14017 16964 14052 16973
rect 14052 16964 14086 16973
rect 14086 16964 14121 16973
rect 14121 16964 14155 16973
rect 14155 16964 14190 16973
rect 14190 16964 14224 16973
rect 14224 16964 14259 16973
rect 14259 16964 14293 16973
rect 14293 16964 14328 16973
rect 14328 16964 14362 16973
rect 14362 16964 14397 16973
rect 14397 16964 14431 16973
rect 14431 16964 14466 16973
rect 14466 16964 14500 16973
rect 14500 16964 14535 16973
rect 14535 16964 14569 16973
rect 14569 16964 14604 16973
rect 14604 16964 14638 16973
rect 14638 16964 14673 16973
rect 14673 16964 14707 16973
rect 14707 16964 14742 16973
rect 14742 16964 14776 16973
rect 14776 16964 14811 16973
rect 14811 16964 14845 16973
rect 14845 16964 14880 16973
rect 14880 16964 14914 16973
rect 14914 16964 14949 16973
rect 14949 16964 14983 16973
rect 14983 16964 15018 16973
rect 15018 16964 15052 16973
rect 15052 16964 15087 16973
rect 15087 16964 15121 16973
rect 15121 16964 15156 16973
rect 15156 16964 15190 16973
rect 15190 16964 15199 16973
rect 17146 16996 17157 16998
rect 17157 16996 17180 16998
rect 17218 16996 17226 16998
rect 17226 16996 17252 16998
rect 17291 16996 17295 16998
rect 17295 16996 17325 16998
rect 17364 16996 17398 16998
rect 17437 16996 17467 16998
rect 17467 16996 17471 16998
rect 17510 16996 17536 16998
rect 17536 16996 17544 16998
rect 17583 16996 17605 16998
rect 17605 16996 17617 16998
rect 17656 16996 17674 16998
rect 17674 16996 17690 16998
rect 17729 16996 17743 16998
rect 17743 16996 17763 16998
rect 17802 16996 17812 16998
rect 17812 16996 17836 16998
rect 17875 16996 17881 16998
rect 17881 16996 17909 16998
rect 17948 16996 17982 16998
rect 678 16928 680 16955
rect 680 16928 712 16955
rect 750 16954 784 16964
rect 678 16921 712 16928
rect 750 16895 782 16908
rect 782 16895 784 16908
rect 678 16859 680 16882
rect 680 16859 712 16882
rect 750 16874 784 16895
rect 678 16848 712 16859
rect 750 16826 782 16828
rect 782 16826 784 16828
rect 678 16790 680 16808
rect 680 16790 712 16808
rect 750 16794 784 16826
rect 678 16774 712 16790
rect 678 16721 680 16734
rect 680 16721 712 16734
rect 750 16722 784 16748
rect 678 16700 712 16721
rect 750 16714 782 16722
rect 782 16714 784 16722
rect 678 16652 680 16660
rect 680 16652 712 16660
rect 750 16653 784 16667
rect 678 16626 712 16652
rect 750 16633 782 16653
rect 782 16633 784 16653
rect 678 16583 680 16586
rect 680 16583 712 16586
rect 750 16584 784 16586
rect 678 16552 712 16583
rect 750 16552 782 16584
rect 782 16552 784 16584
rect 3267 16962 3301 16964
rect 3339 16962 3373 16964
rect 3267 16882 3301 16916
rect 3339 16882 3373 16916
rect 3267 16802 3301 16836
rect 3339 16802 3373 16836
rect 3267 16722 3301 16756
rect 3339 16722 3373 16756
rect 3267 16642 3301 16676
rect 3339 16642 3373 16676
rect 3267 16562 3301 16596
rect 3339 16562 3373 16596
rect 3267 16481 3301 16515
rect 3339 16481 3373 16515
rect 3267 16400 3301 16434
rect 3339 16400 3373 16434
rect 5609 16962 5643 16964
rect 5681 16962 5715 16964
rect 5609 16882 5643 16916
rect 5681 16882 5715 16916
rect 5609 16802 5643 16836
rect 5681 16802 5715 16836
rect 5609 16722 5643 16756
rect 5681 16722 5715 16756
rect 5609 16642 5643 16676
rect 5681 16642 5715 16676
rect 5609 16562 5643 16596
rect 5681 16562 5715 16596
rect 5609 16481 5643 16515
rect 5681 16481 5715 16515
rect 5609 16400 5643 16434
rect 5681 16400 5715 16434
rect 7951 16962 8057 16964
rect 7951 16882 7985 16916
rect 8023 16882 8057 16916
rect 7951 16802 7985 16836
rect 8023 16802 8057 16836
rect 7951 16722 7985 16756
rect 8023 16722 8057 16756
rect 7951 16642 7985 16676
rect 8023 16642 8057 16676
rect 7951 16562 7985 16596
rect 8023 16562 8057 16596
rect 7951 16481 7985 16515
rect 8023 16481 8057 16515
rect 7951 16400 7985 16434
rect 8023 16400 8057 16434
rect 10293 16962 10399 16964
rect 10293 16882 10327 16916
rect 10365 16882 10399 16916
rect 10293 16802 10327 16836
rect 10365 16802 10399 16836
rect 10293 16722 10327 16756
rect 10365 16722 10399 16756
rect 10476 16939 10510 16964
rect 10549 16939 10583 16964
rect 10622 16939 10656 16964
rect 10695 16939 10729 16964
rect 10768 16939 10802 16964
rect 10841 16939 10875 16964
rect 10914 16939 10948 16964
rect 10987 16939 11021 16964
rect 11060 16939 11094 16964
rect 11133 16930 15199 16964
rect 10476 16896 10494 16901
rect 10494 16896 10510 16901
rect 10549 16896 10563 16901
rect 10563 16896 10583 16901
rect 10622 16896 10632 16901
rect 10632 16896 10656 16901
rect 10695 16896 10701 16901
rect 10701 16896 10729 16901
rect 10768 16896 10770 16901
rect 10770 16896 10802 16901
rect 10841 16896 10873 16901
rect 10873 16896 10875 16901
rect 10914 16896 10942 16901
rect 10942 16896 10948 16901
rect 10987 16896 11011 16901
rect 11011 16896 11021 16901
rect 11060 16896 11080 16901
rect 11080 16896 11094 16901
rect 11133 16896 11149 16930
rect 11149 16896 11184 16930
rect 11184 16896 11218 16930
rect 11218 16896 11253 16930
rect 11253 16896 11287 16930
rect 11287 16896 11322 16930
rect 11322 16896 11356 16930
rect 11356 16896 11391 16930
rect 11391 16896 11425 16930
rect 11425 16896 11460 16930
rect 11460 16896 11494 16930
rect 11494 16896 11529 16930
rect 11529 16896 11563 16930
rect 11563 16896 11598 16930
rect 11598 16896 11632 16930
rect 11632 16896 11667 16930
rect 11667 16896 11701 16930
rect 11701 16896 11736 16930
rect 11736 16896 11770 16930
rect 11770 16896 11805 16930
rect 11805 16896 11839 16930
rect 11839 16896 11874 16930
rect 11874 16896 11908 16930
rect 11908 16896 11943 16930
rect 11943 16896 11977 16930
rect 11977 16896 12012 16930
rect 12012 16896 12046 16930
rect 12046 16896 12081 16930
rect 12081 16896 12115 16930
rect 12115 16896 12150 16930
rect 12150 16896 12184 16930
rect 12184 16896 12219 16930
rect 12219 16896 12253 16930
rect 12253 16896 12288 16930
rect 12288 16896 12322 16930
rect 12322 16896 12357 16930
rect 12357 16896 12391 16930
rect 12391 16896 12426 16930
rect 12426 16896 12460 16930
rect 12460 16896 12495 16930
rect 12495 16896 12529 16930
rect 12529 16896 12564 16930
rect 12564 16896 12598 16930
rect 12598 16896 12633 16930
rect 12633 16896 12667 16930
rect 12667 16896 12702 16930
rect 12702 16896 12736 16930
rect 12736 16896 12771 16930
rect 12771 16896 12805 16930
rect 12805 16896 12840 16930
rect 12840 16896 12874 16930
rect 12874 16896 12909 16930
rect 12909 16896 12943 16930
rect 12943 16896 12978 16930
rect 12978 16896 13012 16930
rect 13012 16896 13047 16930
rect 13047 16896 13081 16930
rect 13081 16896 13116 16930
rect 13116 16896 13150 16930
rect 13150 16896 13185 16930
rect 13185 16896 13219 16930
rect 13219 16896 13254 16930
rect 13254 16896 13288 16930
rect 13288 16896 13323 16930
rect 13323 16896 13357 16930
rect 13357 16896 13392 16930
rect 13392 16896 13426 16930
rect 13426 16896 13461 16930
rect 13461 16896 13495 16930
rect 13495 16896 13530 16930
rect 13530 16896 13564 16930
rect 13564 16896 13599 16930
rect 13599 16896 13633 16930
rect 13633 16896 13668 16930
rect 13668 16896 13702 16930
rect 13702 16896 13737 16930
rect 13737 16896 13771 16930
rect 13771 16896 13806 16930
rect 13806 16896 13840 16930
rect 13840 16896 13875 16930
rect 13875 16896 13909 16930
rect 13909 16896 13944 16930
rect 13944 16896 13978 16930
rect 13978 16896 14013 16930
rect 14013 16896 14047 16930
rect 14047 16896 14082 16930
rect 14082 16896 14116 16930
rect 14116 16896 14151 16930
rect 14151 16896 14185 16930
rect 14185 16896 14220 16930
rect 14220 16896 14254 16930
rect 14254 16896 14289 16930
rect 14289 16896 14323 16930
rect 14323 16896 14358 16930
rect 14358 16896 14392 16930
rect 14392 16896 14427 16930
rect 14427 16896 14461 16930
rect 14461 16896 14496 16930
rect 10476 16867 10510 16896
rect 10549 16867 10583 16896
rect 10622 16867 10656 16896
rect 10695 16867 10729 16896
rect 10768 16867 10802 16896
rect 10841 16867 10875 16896
rect 10914 16867 10948 16896
rect 10987 16867 11021 16896
rect 11060 16867 11094 16896
rect 11133 16867 14496 16896
rect 14496 16867 15199 16930
rect 15396 16888 15430 16922
rect 15396 16815 15430 16849
rect 10293 16642 10327 16676
rect 10365 16642 10399 16676
rect 10293 16562 10327 16596
rect 10365 16562 10399 16596
rect 10293 16481 10327 16515
rect 10365 16481 10399 16515
rect 10293 16400 10327 16434
rect 10365 16400 10399 16434
rect 15396 16742 15430 16776
rect 15396 16669 15430 16703
rect 15396 16596 15430 16630
rect 15396 16523 15430 16557
rect 15396 16450 15430 16484
rect 14969 16281 15003 16315
rect 15041 16281 15075 16315
rect 15162 16347 15196 16381
rect 15162 16275 15196 16309
rect 14969 16195 15003 16229
rect 15041 16195 15075 16229
rect 15162 16201 15196 16235
rect 15162 16129 15196 16163
rect 680 14712 714 14746
rect 752 14712 786 14746
rect 680 14637 714 14671
rect 752 14637 786 14671
rect 680 14562 714 14596
rect 752 14562 786 14596
rect 680 14487 714 14521
rect 752 14487 786 14521
rect 680 14412 714 14446
rect 752 14412 786 14446
rect 680 14337 714 14371
rect 752 14337 786 14371
rect 680 14262 714 14296
rect 752 14262 786 14296
rect 680 14187 714 14221
rect 752 14187 786 14221
rect 680 14112 714 14146
rect 752 14112 786 14146
rect 680 14037 714 14071
rect 752 14037 786 14071
rect 680 13962 714 13996
rect 752 13962 786 13996
rect 680 13887 714 13921
rect 752 13887 786 13921
rect 3267 14880 3301 14914
rect 3339 14880 3373 14914
rect 3267 14804 3301 14838
rect 3339 14804 3373 14838
rect 3267 14727 3301 14761
rect 3339 14727 3373 14761
rect 7951 14880 7985 14914
rect 8023 14880 8057 14914
rect 7951 14804 7985 14838
rect 8023 14804 8057 14838
rect 7951 14727 7985 14761
rect 8023 14727 8057 14761
rect 3267 14650 3301 14684
rect 3339 14650 3373 14684
rect 3267 14573 3301 14607
rect 3339 14573 3373 14607
rect 3267 14496 3301 14530
rect 3339 14496 3373 14530
rect 3267 14419 3301 14453
rect 3339 14419 3373 14453
rect 3267 14342 3301 14376
rect 3339 14342 3373 14376
rect 3267 14265 3301 14299
rect 3339 14265 3373 14299
rect 3267 14188 3301 14222
rect 3339 14188 3373 14222
rect 3267 14111 3301 14145
rect 3339 14111 3373 14145
rect 3267 14034 3301 14068
rect 3339 14034 3373 14068
rect 3267 13957 3301 13991
rect 3339 13957 3373 13991
rect 3267 13880 3301 13914
rect 3339 13880 3373 13914
rect 5609 14683 5643 14717
rect 5681 14683 5715 14717
rect 5609 14610 5643 14644
rect 5681 14610 5715 14644
rect 5609 14537 5643 14571
rect 5681 14537 5715 14571
rect 5609 14464 5643 14498
rect 5681 14464 5715 14498
rect 5609 14391 5643 14425
rect 5681 14391 5715 14425
rect 5609 14318 5643 14352
rect 5681 14318 5715 14352
rect 5609 14245 5643 14279
rect 5681 14245 5715 14279
rect 5609 14172 5643 14206
rect 5681 14172 5715 14206
rect 5609 14099 5643 14133
rect 5681 14099 5715 14133
rect 5609 14026 5643 14060
rect 5681 14026 5715 14060
rect 5609 13953 5643 13987
rect 5681 13953 5715 13987
rect 5609 13880 5643 13914
rect 5681 13880 5715 13914
rect 12682 14880 12716 14914
rect 12754 14880 12788 14914
rect 12682 14804 12716 14838
rect 12754 14804 12788 14838
rect 12682 14727 12716 14761
rect 12754 14727 12788 14761
rect 7951 14650 7985 14684
rect 8023 14650 8057 14684
rect 7951 14573 7985 14607
rect 8023 14573 8057 14607
rect 7951 14496 7985 14530
rect 8023 14496 8057 14530
rect 7951 14419 7985 14453
rect 8023 14419 8057 14453
rect 7951 14342 7985 14376
rect 8023 14342 8057 14376
rect 7951 14265 7985 14299
rect 8023 14265 8057 14299
rect 7951 14188 7985 14222
rect 8023 14188 8057 14222
rect 7951 14111 7985 14145
rect 8023 14111 8057 14145
rect 7951 14034 7985 14068
rect 8023 14034 8057 14068
rect 7951 13957 7985 13991
rect 8023 13957 8057 13991
rect 7951 13880 7985 13914
rect 8023 13880 8057 13914
rect 10293 14683 10327 14717
rect 10365 14683 10399 14717
rect 10293 14610 10327 14644
rect 10365 14610 10399 14644
rect 10293 14537 10327 14571
rect 10365 14537 10399 14571
rect 10293 14464 10327 14498
rect 10365 14464 10399 14498
rect 10293 14391 10327 14425
rect 10365 14391 10399 14425
rect 10293 14318 10327 14352
rect 10365 14318 10399 14352
rect 10293 14245 10327 14279
rect 10365 14245 10399 14279
rect 10293 14172 10327 14206
rect 10365 14172 10399 14206
rect 10293 14099 10327 14133
rect 10365 14099 10399 14133
rect 10293 14026 10327 14060
rect 10365 14026 10399 14060
rect 10293 13953 10327 13987
rect 10365 13953 10399 13987
rect 10293 13880 10327 13914
rect 10365 13880 10399 13914
rect 14986 14942 15020 14976
rect 14986 14870 15020 14904
rect 15159 14876 15193 14910
rect 12682 14650 12716 14684
rect 12754 14650 12788 14684
rect 12682 14573 12716 14607
rect 12754 14573 12788 14607
rect 12682 14496 12716 14530
rect 12754 14496 12788 14530
rect 12682 14419 12716 14453
rect 12754 14419 12788 14453
rect 12682 14342 12716 14376
rect 12754 14342 12788 14376
rect 12682 14265 12716 14299
rect 12754 14265 12788 14299
rect 12682 14188 12716 14222
rect 12754 14188 12788 14222
rect 14986 14609 15020 14643
rect 14986 14537 15020 14571
rect 12682 14111 12716 14145
rect 12754 14111 12788 14145
rect 12682 14034 12716 14068
rect 12754 14034 12788 14068
rect 12682 13957 12716 13991
rect 12754 13957 12788 13991
rect 12682 13880 12716 13914
rect 12754 13880 12788 13914
rect 15159 14804 15193 14838
rect 15159 14603 15193 14637
rect 15159 14531 15193 14565
rect 680 13812 714 13846
rect 752 13812 786 13846
rect 680 13737 714 13771
rect 752 13737 786 13771
rect 680 13662 714 13696
rect 752 13662 786 13696
rect 680 13587 714 13621
rect 752 13587 786 13621
rect 680 13513 714 13547
rect 752 13513 786 13547
rect 680 13439 714 13473
rect 752 13439 786 13473
rect 680 13365 714 13399
rect 752 13365 786 13399
rect 680 13291 714 13325
rect 752 13291 786 13325
rect 680 13217 714 13251
rect 752 13217 786 13251
rect 680 13143 714 13177
rect 752 13143 786 13177
rect 680 13069 714 13103
rect 752 13069 786 13103
rect 15396 16377 15430 16411
rect 15396 16304 15430 16338
rect 15396 16231 15430 16265
rect 17948 16924 18054 16992
rect 18020 16886 18054 16920
rect 17948 16851 17982 16885
rect 18020 16814 18054 16848
rect 17948 16778 17982 16812
rect 18020 16742 18054 16776
rect 17948 16705 17982 16739
rect 18020 16670 18054 16704
rect 17948 16632 17982 16666
rect 18020 16624 18054 16632
rect 18020 16598 18052 16624
rect 18052 16598 18054 16624
rect 17948 16589 17982 16593
rect 17948 16559 17950 16589
rect 17950 16559 17982 16589
rect 18020 16556 18054 16559
rect 18020 16525 18052 16556
rect 18052 16525 18054 16556
rect 17948 16486 17950 16520
rect 17950 16486 17982 16520
rect 18020 16454 18052 16486
rect 18052 16454 18054 16486
rect 18020 16452 18054 16454
rect 17948 16417 17950 16447
rect 17950 16417 17982 16447
rect 17948 16413 17982 16417
rect 18020 16386 18052 16413
rect 18052 16386 18054 16413
rect 17948 16348 17950 16374
rect 17950 16348 17982 16374
rect 18020 16379 18054 16386
rect 17948 16340 17982 16348
rect 18020 16318 18052 16340
rect 18052 16318 18054 16340
rect 17948 16279 17950 16301
rect 17950 16279 17982 16301
rect 18020 16306 18054 16318
rect 17948 16267 17982 16279
rect 18020 16250 18052 16267
rect 18052 16250 18054 16267
rect 17948 16210 17950 16228
rect 17950 16210 17982 16228
rect 18020 16233 18054 16250
rect 15396 16158 15430 16192
rect 15396 16085 15430 16119
rect 17948 16194 17982 16210
rect 18020 16182 18052 16194
rect 18052 16182 18054 16194
rect 17948 16141 17950 16155
rect 17950 16141 17982 16155
rect 18020 16160 18054 16182
rect 17948 16121 17982 16141
rect 18020 16114 18052 16121
rect 18052 16114 18054 16121
rect 15396 16012 15430 16046
rect 15396 15939 15430 15973
rect 15396 15866 15430 15900
rect 15396 15793 15430 15827
rect 15396 15720 15430 15754
rect 15396 15647 15430 15681
rect 15396 15574 15430 15608
rect 15396 15501 15430 15535
rect 15396 15428 15430 15462
rect 15396 15355 15430 15389
rect 15396 15282 15430 15316
rect 15396 15209 15430 15243
rect 15396 15136 15430 15170
rect 15396 15063 15430 15097
rect 15396 14990 15430 15024
rect 15396 14917 15430 14951
rect 15396 14844 15430 14878
rect 15396 14788 15430 14805
rect 15396 14771 15430 14788
rect 15396 14719 15430 14732
rect 15396 14698 15430 14719
rect 15396 14650 15430 14658
rect 15396 14624 15430 14650
rect 15396 14581 15430 14584
rect 15396 14550 15430 14581
rect 15396 14477 15430 14510
rect 15396 14476 15430 14477
rect 15396 14408 15430 14436
rect 15396 14402 15430 14408
rect 15396 14340 15430 14362
rect 15396 14328 15430 14340
rect 15396 14269 15430 14288
rect 15396 14254 15430 14269
rect 15396 14198 15430 14214
rect 15396 14180 15430 14198
rect 15396 14127 15430 14140
rect 15396 14106 15430 14127
rect 15396 14056 15430 14066
rect 15396 14032 15430 14056
rect 15396 13985 15430 13992
rect 15396 13958 15430 13985
rect 15396 13914 15430 13918
rect 15396 13884 15430 13914
rect 15396 13843 15430 13844
rect 15396 13810 15430 13843
rect 15396 13738 15430 13770
rect 15396 13736 15430 13738
rect 15396 13667 15430 13696
rect 15396 13662 15430 13667
rect 15396 13596 15430 13622
rect 15396 13588 15430 13596
rect 15396 13525 15430 13548
rect 15396 13514 15430 13525
rect 15396 13454 15430 13474
rect 15396 13440 15430 13454
rect 15396 13383 15430 13400
rect 15396 13366 15430 13383
rect 15396 13312 15430 13326
rect 15396 13292 15430 13312
rect 15396 13241 15430 13252
rect 15396 13218 15430 13241
rect 17948 16072 17950 16082
rect 17950 16072 17982 16082
rect 18020 16087 18054 16114
rect 17948 16048 17982 16072
rect 18020 16046 18052 16048
rect 18052 16046 18054 16048
rect 17948 16003 17950 16009
rect 17950 16003 17982 16009
rect 18020 16014 18054 16046
rect 17948 15975 17982 16003
rect 17948 15934 17950 15936
rect 17950 15934 17982 15936
rect 18020 15944 18054 15975
rect 18020 15941 18052 15944
rect 18052 15941 18054 15944
rect 17948 15902 17982 15934
rect 18020 15876 18054 15902
rect 18020 15868 18052 15876
rect 18052 15868 18054 15876
rect 17948 15830 17982 15863
rect 17948 15829 17950 15830
rect 17950 15829 17982 15830
rect 14823 13104 14857 13138
rect 14895 13104 14929 13138
rect 14969 13104 15003 13138
rect 15041 13104 15075 13138
rect 15123 13104 15157 13138
rect 15195 13104 15229 13138
rect 18020 15808 18054 15829
rect 18020 15795 18052 15808
rect 18052 15795 18054 15808
rect 17948 15761 17982 15790
rect 17948 15756 17950 15761
rect 17950 15756 17982 15761
rect 18020 15740 18054 15756
rect 18020 15722 18052 15740
rect 18052 15722 18054 15740
rect 17948 15692 17982 15717
rect 17948 15683 17950 15692
rect 17950 15683 17982 15692
rect 18020 15672 18054 15683
rect 18020 15649 18052 15672
rect 18052 15649 18054 15672
rect 17948 15623 17982 15644
rect 17948 15610 17950 15623
rect 17950 15610 17982 15623
rect 18020 15604 18054 15610
rect 18020 15576 18052 15604
rect 18052 15576 18054 15604
rect 17948 15554 17982 15571
rect 17948 15537 17950 15554
rect 17950 15537 17982 15554
rect 18020 15536 18054 15537
rect 18020 15503 18052 15536
rect 18052 15503 18054 15536
rect 17948 15485 17982 15498
rect 17948 15464 17950 15485
rect 17950 15464 17982 15485
rect 18020 15434 18052 15464
rect 18052 15434 18054 15464
rect 18020 15430 18054 15434
rect 17948 15416 17982 15425
rect 17948 15391 17950 15416
rect 17950 15391 17982 15416
rect 18020 15366 18052 15391
rect 18052 15366 18054 15391
rect 18020 15357 18054 15366
rect 17948 15347 17982 15352
rect 17948 15318 17950 15347
rect 17950 15318 17982 15347
rect 18020 15298 18052 15318
rect 18052 15298 18054 15318
rect 18020 15284 18054 15298
rect 17948 15278 17982 15279
rect 17948 15245 17950 15278
rect 17950 15245 17982 15278
rect 18020 15230 18052 15245
rect 18052 15230 18054 15245
rect 18020 15211 18054 15230
rect 17948 15175 17950 15206
rect 17950 15175 17982 15206
rect 17948 15172 17982 15175
rect 18020 15162 18052 15172
rect 18052 15162 18054 15172
rect 17948 15106 17950 15133
rect 17950 15106 17982 15133
rect 18020 15138 18054 15162
rect 17948 15099 17982 15106
rect 18020 15094 18052 15099
rect 18052 15094 18054 15099
rect 17948 15037 17950 15060
rect 17950 15037 17982 15060
rect 18020 15065 18054 15094
rect 17948 15026 17982 15037
rect 680 12995 714 13029
rect 752 12995 786 13029
rect 15241 13009 15275 13043
rect 15313 13009 15347 13043
rect 15387 13009 15421 13043
rect 15459 13009 15493 13043
rect 15533 13009 15567 13043
rect 15605 13009 15639 13043
rect 17948 14968 17950 14987
rect 17950 14968 17982 14987
rect 18020 14992 18054 15026
rect 17948 14953 17982 14968
rect 17948 14899 17950 14914
rect 17950 14899 17982 14914
rect 18020 14924 18054 14953
rect 18020 14919 18052 14924
rect 18052 14919 18054 14924
rect 17948 14880 17982 14899
rect 17948 14830 17950 14841
rect 17950 14830 17982 14841
rect 18020 14856 18054 14880
rect 18020 14846 18052 14856
rect 18052 14846 18054 14856
rect 17948 14807 17982 14830
rect 17948 14761 17950 14768
rect 17950 14761 17982 14768
rect 18020 14788 18054 14807
rect 18020 14773 18052 14788
rect 18052 14773 18054 14788
rect 17948 14734 17982 14761
rect 17948 14692 17950 14695
rect 17950 14692 17982 14695
rect 18020 14720 18054 14734
rect 18020 14700 18052 14720
rect 18052 14700 18054 14720
rect 17948 14661 17982 14692
rect 18020 14652 18054 14661
rect 18020 14627 18052 14652
rect 18052 14627 18054 14652
rect 17948 14588 17982 14622
rect 18020 14584 18054 14588
rect 18020 14554 18052 14584
rect 18052 14554 18054 14584
rect 17948 14519 17982 14549
rect 17948 14515 17950 14519
rect 17950 14515 17982 14519
rect 18020 14482 18052 14515
rect 18052 14482 18054 14515
rect 18020 14481 18054 14482
rect 17948 14450 17982 14476
rect 17948 14442 17950 14450
rect 17950 14442 17982 14450
rect 18020 14414 18052 14442
rect 18052 14414 18054 14442
rect 18020 14408 18054 14414
rect 17948 14381 17982 14403
rect 17948 14369 17950 14381
rect 17950 14369 17982 14381
rect 18020 14346 18052 14369
rect 18052 14346 18054 14369
rect 18020 14335 18054 14346
rect 17948 14312 17982 14330
rect 17948 14296 17950 14312
rect 17950 14296 17982 14312
rect 18020 14278 18052 14296
rect 18052 14278 18054 14296
rect 18020 14262 18054 14278
rect 17948 14243 17982 14257
rect 17948 14223 17950 14243
rect 17950 14223 17982 14243
rect 18020 14209 18052 14223
rect 18052 14209 18054 14223
rect 18020 14189 18054 14209
rect 17948 14174 17982 14184
rect 17948 14150 17950 14174
rect 17950 14150 17982 14174
rect 18020 14140 18052 14150
rect 18052 14140 18054 14150
rect 18020 14116 18054 14140
rect 17948 14105 17982 14111
rect 17948 14077 17950 14105
rect 17950 14077 17982 14105
rect 18020 14071 18052 14077
rect 18052 14071 18054 14077
rect 18020 14043 18054 14071
rect 17948 14036 17982 14038
rect 17948 14004 17950 14036
rect 17950 14004 17982 14036
rect 18020 14002 18052 14004
rect 18052 14002 18054 14004
rect 18020 13970 18054 14002
rect 17948 13933 17950 13965
rect 17950 13933 17982 13965
rect 17948 13931 17982 13933
rect 18020 13898 18054 13931
rect 17948 13864 17950 13892
rect 17950 13864 17982 13892
rect 18020 13897 18052 13898
rect 18052 13897 18054 13898
rect 17948 13858 17982 13864
rect 18020 13829 18054 13858
rect 17948 13795 17950 13819
rect 17950 13795 17982 13819
rect 18020 13824 18052 13829
rect 18052 13824 18054 13829
rect 17948 13785 17982 13795
rect 18020 13760 18054 13785
rect 17948 13726 17950 13746
rect 17950 13726 17982 13746
rect 18020 13751 18052 13760
rect 18052 13751 18054 13760
rect 17948 13712 17982 13726
rect 18020 13691 18054 13712
rect 17948 13657 17950 13673
rect 17950 13657 17982 13673
rect 18020 13678 18052 13691
rect 18052 13678 18054 13691
rect 17948 13639 17982 13657
rect 18020 13622 18054 13639
rect 17948 13588 17950 13600
rect 17950 13588 17982 13600
rect 18020 13605 18052 13622
rect 18052 13605 18054 13622
rect 17948 13566 17982 13588
rect 18020 13553 18054 13566
rect 17948 13519 17950 13527
rect 17950 13519 17982 13527
rect 18020 13532 18052 13553
rect 18052 13532 18054 13553
rect 17948 13493 17982 13519
rect 18020 13484 18054 13493
rect 17948 13450 17950 13454
rect 17950 13450 17982 13454
rect 18020 13459 18052 13484
rect 18052 13459 18054 13484
rect 17948 13420 17982 13450
rect 18020 13415 18054 13420
rect 18020 13386 18052 13415
rect 18052 13386 18054 13415
rect 17948 13347 17982 13381
rect 18020 13346 18054 13347
rect 18020 13313 18052 13346
rect 18052 13313 18054 13346
rect 17948 13277 17982 13308
rect 17948 13274 17950 13277
rect 17950 13274 17982 13277
rect 18020 13243 18052 13274
rect 18052 13243 18054 13274
rect 18020 13240 18054 13243
rect 17948 13208 17982 13235
rect 17948 13201 17950 13208
rect 17950 13201 17982 13208
rect 18020 13174 18052 13201
rect 18052 13174 18054 13201
rect 18020 13167 18054 13174
rect 17948 13139 17982 13162
rect 17948 13128 17950 13139
rect 17950 13128 17982 13139
rect 18020 13105 18052 13128
rect 18052 13105 18054 13128
rect 18020 13094 18054 13105
rect 17948 13070 17982 13089
rect 17948 13055 17950 13070
rect 17950 13055 17982 13070
rect 18020 13036 18052 13055
rect 18052 13036 18054 13055
rect 18020 13021 18054 13036
rect 17948 13001 17982 13016
rect 17948 12982 17950 13001
rect 17950 12982 17982 13001
rect 680 12921 714 12955
rect 752 12941 786 12955
rect 18020 12967 18052 12982
rect 18052 12967 18054 12982
rect 18020 12948 18054 12967
rect 829 12941 851 12943
rect 851 12941 885 12943
rect 885 12941 920 12943
rect 920 12941 954 12943
rect 954 12941 989 12943
rect 989 12941 1023 12943
rect 1023 12941 1058 12943
rect 1058 12941 1092 12943
rect 1092 12941 1127 12943
rect 1127 12941 1161 12943
rect 1161 12941 1196 12943
rect 1196 12941 1230 12943
rect 1230 12941 1265 12943
rect 1265 12941 1299 12943
rect 1299 12941 1334 12943
rect 1334 12941 1368 12943
rect 1368 12941 1403 12943
rect 1403 12941 1437 12943
rect 1437 12941 1472 12943
rect 1472 12941 1506 12943
rect 1506 12941 1541 12943
rect 1541 12941 1575 12943
rect 1575 12941 1610 12943
rect 1610 12941 1644 12943
rect 1644 12941 1679 12943
rect 1679 12941 1713 12943
rect 1713 12941 1748 12943
rect 1748 12941 1782 12943
rect 1782 12941 1817 12943
rect 1817 12941 1851 12943
rect 1851 12941 1886 12943
rect 1886 12941 1920 12943
rect 1920 12941 1955 12943
rect 1955 12941 1989 12943
rect 1989 12941 2024 12943
rect 2024 12941 2058 12943
rect 2058 12941 2093 12943
rect 2093 12941 2127 12943
rect 2127 12941 2162 12943
rect 2162 12941 2196 12943
rect 2196 12941 2231 12943
rect 2231 12941 2265 12943
rect 2265 12941 2300 12943
rect 2300 12941 2334 12943
rect 2334 12941 2369 12943
rect 2369 12941 2403 12943
rect 2403 12941 2438 12943
rect 752 12921 786 12941
rect 829 12907 2438 12941
rect 680 12847 714 12881
rect 752 12873 783 12881
rect 783 12873 786 12881
rect 829 12873 852 12907
rect 852 12873 886 12907
rect 886 12873 921 12907
rect 921 12873 955 12907
rect 955 12873 990 12907
rect 990 12873 1024 12907
rect 1024 12873 1059 12907
rect 1059 12873 1093 12907
rect 1093 12873 1128 12907
rect 1128 12873 1162 12907
rect 1162 12873 1197 12907
rect 1197 12873 1231 12907
rect 1231 12873 1266 12907
rect 1266 12873 1300 12907
rect 1300 12873 1335 12907
rect 1335 12873 1369 12907
rect 1369 12873 1404 12907
rect 1404 12873 1438 12907
rect 1438 12873 1473 12907
rect 1473 12873 1507 12907
rect 1507 12873 1542 12907
rect 1542 12873 1576 12907
rect 1576 12873 1611 12907
rect 1611 12873 1645 12907
rect 1645 12873 1680 12907
rect 1680 12873 1714 12907
rect 1714 12873 1749 12907
rect 1749 12873 1783 12907
rect 1783 12873 1818 12907
rect 1818 12873 1852 12907
rect 1852 12873 1887 12907
rect 1887 12873 1921 12907
rect 1921 12873 1956 12907
rect 1956 12873 1990 12907
rect 1990 12873 2025 12907
rect 2025 12873 2059 12907
rect 2059 12873 2094 12907
rect 2094 12873 2128 12907
rect 2128 12873 2163 12907
rect 2163 12873 2197 12907
rect 2197 12873 2232 12907
rect 2232 12873 2266 12907
rect 2266 12873 2301 12907
rect 2301 12873 2335 12907
rect 2335 12873 2370 12907
rect 2370 12873 2404 12907
rect 2404 12873 2438 12907
rect 2438 12873 12311 12943
rect 12350 12909 12384 12943
rect 12423 12909 12457 12943
rect 12496 12909 12530 12943
rect 12569 12909 12603 12943
rect 12642 12909 12676 12943
rect 12715 12909 12749 12943
rect 12788 12909 12822 12943
rect 12861 12909 12895 12943
rect 12934 12909 12968 12943
rect 13007 12909 13041 12943
rect 13080 12909 13114 12943
rect 13153 12909 13187 12943
rect 13226 12909 13260 12943
rect 13299 12909 13333 12943
rect 13372 12909 13406 12943
rect 13445 12909 13479 12943
rect 13518 12909 13552 12943
rect 13591 12909 13625 12943
rect 13664 12909 13698 12943
rect 13737 12909 13771 12943
rect 13810 12909 13844 12943
rect 13883 12909 13917 12943
rect 13956 12909 13990 12943
rect 14029 12909 14063 12943
rect 14102 12909 14136 12943
rect 14175 12909 14209 12943
rect 14248 12909 14282 12943
rect 14321 12909 14355 12943
rect 14394 12909 14428 12943
rect 14467 12909 14501 12943
rect 14540 12909 14574 12943
rect 15752 12909 15786 12943
rect 15826 12909 15860 12943
rect 15900 12909 15934 12943
rect 15974 12909 16008 12943
rect 16048 12909 16082 12943
rect 16122 12909 16156 12943
rect 16196 12909 16230 12943
rect 16269 12909 16303 12943
rect 16342 12909 16376 12943
rect 16415 12909 16449 12943
rect 16488 12909 16522 12943
rect 16561 12909 16595 12943
rect 16634 12909 16668 12943
rect 16707 12909 16741 12943
rect 16780 12909 16814 12943
rect 16853 12909 16887 12943
rect 16926 12909 16960 12943
rect 16999 12909 17033 12943
rect 17072 12909 17106 12943
rect 17145 12909 17179 12943
rect 17218 12909 17252 12943
rect 17291 12909 17325 12943
rect 17364 12909 17398 12943
rect 17437 12909 17471 12943
rect 17510 12909 17544 12943
rect 17583 12909 17617 12943
rect 17656 12909 17690 12943
rect 17729 12909 17763 12943
rect 17802 12909 17836 12943
rect 17875 12909 17909 12943
rect 17948 12932 17982 12943
rect 17948 12909 17950 12932
rect 17950 12909 17982 12932
rect 752 12847 786 12873
rect 829 12839 4682 12873
rect 829 12837 852 12839
rect 852 12837 887 12839
rect 887 12837 921 12839
rect 921 12837 956 12839
rect 956 12837 990 12839
rect 990 12837 1025 12839
rect 1025 12837 1059 12839
rect 1059 12837 1094 12839
rect 1094 12837 1128 12839
rect 1128 12837 1163 12839
rect 1163 12837 1197 12839
rect 1197 12837 1232 12839
rect 1232 12837 1266 12839
rect 1266 12837 1301 12839
rect 1301 12837 1335 12839
rect 1335 12837 1370 12839
rect 1370 12837 1404 12839
rect 1404 12837 1439 12839
rect 1439 12837 1473 12839
rect 1473 12837 1508 12839
rect 1508 12837 1542 12839
rect 1542 12837 1577 12839
rect 1577 12837 1611 12839
rect 1611 12837 1646 12839
rect 1646 12837 1680 12839
rect 1680 12837 1715 12839
rect 1715 12837 1749 12839
rect 1749 12837 1784 12839
rect 1784 12837 1818 12839
rect 1818 12837 1853 12839
rect 1853 12837 1887 12839
rect 1887 12837 1922 12839
rect 1922 12837 1956 12839
rect 1956 12837 1991 12839
rect 1991 12837 2025 12839
rect 2025 12837 2060 12839
rect 2060 12837 2094 12839
rect 2094 12837 2129 12839
rect 2129 12837 2163 12839
rect 2163 12837 2198 12839
rect 2198 12837 2232 12839
rect 2232 12837 2267 12839
rect 2267 12837 2301 12839
rect 2301 12837 2336 12839
rect 2336 12837 2370 12839
rect 2370 12837 2405 12839
rect 2405 12837 2439 12839
rect 2439 12837 2474 12839
rect 2474 12837 2508 12839
rect 2508 12837 2543 12839
rect 2543 12837 2577 12839
rect 2577 12837 2612 12839
rect 2612 12837 2646 12839
rect 2646 12837 2681 12839
rect 2681 12837 2715 12839
rect 2715 12837 2750 12839
rect 2750 12837 2784 12839
rect 2784 12837 2819 12839
rect 2819 12837 2853 12839
rect 2853 12837 2888 12839
rect 2888 12837 2922 12839
rect 2922 12837 2957 12839
rect 2957 12837 2991 12839
rect 2991 12837 3026 12839
rect 3026 12837 3060 12839
rect 3060 12837 3095 12839
rect 3095 12837 3129 12839
rect 3129 12837 3164 12839
rect 3164 12837 3198 12839
rect 3198 12837 3233 12839
rect 3233 12837 3267 12839
rect 3267 12837 3302 12839
rect 3302 12837 3336 12839
rect 3336 12837 3371 12839
rect 3371 12837 3405 12839
rect 3405 12837 3440 12839
rect 3440 12837 3474 12839
rect 3474 12837 3509 12839
rect 3509 12837 3543 12839
rect 3543 12837 3578 12839
rect 3578 12837 3612 12839
rect 3612 12837 3647 12839
rect 3647 12837 3681 12839
rect 3681 12837 3716 12839
rect 3716 12837 3750 12839
rect 3750 12837 3785 12839
rect 3785 12837 3819 12839
rect 3819 12837 3854 12839
rect 3854 12837 3888 12839
rect 3888 12837 3923 12839
rect 3923 12837 3957 12839
rect 3957 12837 3992 12839
rect 3992 12837 4026 12839
rect 4026 12837 4061 12839
rect 4061 12837 4095 12839
rect 4095 12837 4130 12839
rect 4130 12837 4164 12839
rect 4164 12837 4199 12839
rect 4199 12837 4233 12839
rect 4233 12837 4268 12839
rect 4268 12837 4302 12839
rect 4302 12837 4337 12839
rect 4337 12837 4371 12839
rect 4371 12837 4406 12839
rect 4406 12837 4440 12839
rect 4440 12837 4475 12839
rect 4475 12837 4509 12839
rect 4509 12837 4544 12839
rect 4544 12837 4578 12839
rect 4578 12837 4613 12839
rect 4613 12837 4647 12839
rect 4647 12837 4682 12839
rect 4682 12837 12311 12873
rect 18020 12898 18052 12909
rect 18052 12898 18054 12909
rect 18020 12875 18054 12898
rect 12350 12837 12384 12871
rect 12423 12837 12457 12871
rect 12496 12837 12530 12871
rect 12569 12837 12603 12871
rect 12642 12837 12676 12871
rect 12715 12837 12749 12871
rect 12788 12837 12822 12871
rect 12861 12837 12895 12871
rect 12934 12837 12968 12871
rect 13007 12837 13041 12871
rect 13080 12837 13114 12871
rect 13153 12837 13187 12871
rect 13226 12837 13260 12871
rect 13299 12837 13333 12871
rect 13372 12837 13406 12871
rect 13445 12837 13479 12871
rect 13518 12837 13552 12871
rect 13591 12837 13625 12871
rect 13664 12837 13698 12871
rect 13737 12837 13771 12871
rect 13810 12837 13844 12871
rect 13883 12837 13917 12871
rect 13956 12837 13990 12871
rect 14029 12837 14063 12871
rect 14102 12837 14136 12871
rect 14175 12837 14209 12871
rect 14248 12837 14282 12871
rect 14321 12837 14355 12871
rect 14394 12837 14428 12871
rect 14467 12837 14501 12871
rect 14540 12837 14574 12871
rect 15752 12837 15786 12871
rect 15827 12837 15861 12871
rect 15902 12837 15936 12871
rect 15977 12837 16011 12871
rect 16052 12837 16086 12871
rect 16127 12837 16161 12871
rect 16202 12837 16236 12871
rect 16277 12837 16311 12871
rect 16352 12837 16386 12871
rect 16426 12837 16460 12871
rect 16500 12837 16534 12871
rect 16574 12837 16608 12871
rect 16648 12837 16682 12871
rect 16722 12837 16756 12871
rect 16796 12837 16830 12871
rect 16870 12837 16904 12871
rect 16944 12837 16978 12871
rect 17018 12837 17052 12871
rect 17092 12837 17126 12871
rect 17166 12837 17200 12871
rect 17240 12837 17274 12871
rect 17314 12837 17348 12871
rect 17388 12837 17422 12871
rect 17462 12837 17496 12871
rect 17536 12837 17570 12871
rect 17610 12837 17644 12871
rect 17684 12837 17718 12871
rect 17758 12837 17792 12871
rect 17832 12837 17840 12871
rect 17840 12837 17866 12871
rect 17906 12863 17940 12871
rect 17906 12837 17916 12863
rect 17916 12837 17940 12863
rect 18271 16455 18377 17315
rect 18343 16417 18377 16451
rect 18271 16382 18305 16416
rect 18343 16345 18377 16379
rect 18271 16309 18305 16343
rect 18343 16273 18377 16307
rect 18271 16236 18305 16270
rect 18343 16201 18377 16235
rect 18271 16163 18305 16197
rect 18343 16129 18377 16163
rect 18271 16090 18305 16124
rect 18343 16056 18377 16090
rect 18271 16017 18305 16051
rect 18343 15983 18377 16017
rect 18271 15944 18305 15978
rect 18343 15910 18377 15944
rect 18271 15871 18305 15905
rect 18343 15837 18377 15871
rect 18271 15798 18305 15832
rect 18343 15764 18377 15798
rect 18271 15725 18305 15759
rect 18343 15691 18377 15725
rect 18271 15654 18273 15686
rect 18273 15654 18305 15686
rect 18271 15652 18305 15654
rect 18343 15621 18375 15652
rect 18375 15621 18377 15652
rect 18271 15585 18273 15613
rect 18273 15585 18305 15613
rect 18343 15618 18377 15621
rect 18271 15579 18305 15585
rect 18343 15552 18375 15579
rect 18375 15552 18377 15579
rect 18271 15516 18273 15540
rect 18273 15516 18305 15540
rect 18343 15545 18377 15552
rect 18271 15506 18305 15516
rect 18343 15483 18375 15506
rect 18375 15483 18377 15506
rect 18271 15447 18273 15467
rect 18273 15447 18305 15467
rect 18343 15472 18377 15483
rect 18271 15433 18305 15447
rect 18343 15414 18375 15433
rect 18375 15414 18377 15433
rect 18271 15378 18273 15394
rect 18273 15378 18305 15394
rect 18343 15399 18377 15414
rect 18271 15360 18305 15378
rect 18343 15345 18375 15360
rect 18375 15345 18377 15360
rect 18271 15309 18273 15321
rect 18273 15309 18305 15321
rect 18343 15326 18377 15345
rect 18271 15287 18305 15309
rect 18343 15276 18375 15287
rect 18375 15276 18377 15287
rect 18271 15240 18273 15248
rect 18273 15240 18305 15248
rect 18343 15253 18377 15276
rect 18271 15214 18305 15240
rect 18343 15207 18375 15214
rect 18375 15207 18377 15214
rect 18271 15171 18273 15175
rect 18273 15171 18305 15175
rect 18343 15180 18377 15207
rect 18271 15141 18305 15171
rect 18343 15138 18375 15141
rect 18375 15138 18377 15141
rect 18343 15107 18377 15138
rect 18271 15068 18305 15102
rect 18343 15034 18377 15068
rect 18271 14998 18305 15029
rect 18271 14995 18273 14998
rect 18273 14995 18305 14998
rect 18343 14965 18377 14995
rect 18343 14961 18375 14965
rect 18375 14961 18377 14965
rect 18271 14929 18305 14956
rect 18271 14922 18273 14929
rect 18273 14922 18305 14929
rect 18343 14896 18377 14922
rect 18343 14888 18375 14896
rect 18375 14888 18377 14896
rect 18271 14860 18305 14883
rect 18271 14849 18273 14860
rect 18273 14849 18305 14860
rect 18343 14827 18377 14849
rect 18343 14815 18375 14827
rect 18375 14815 18377 14827
rect 18271 14791 18305 14810
rect 18271 14776 18273 14791
rect 18273 14776 18305 14791
rect 18343 14758 18377 14776
rect 18343 14742 18375 14758
rect 18375 14742 18377 14758
rect 18271 14722 18305 14737
rect 18271 14703 18273 14722
rect 18273 14703 18305 14722
rect 18343 14689 18377 14703
rect 18343 14669 18375 14689
rect 18375 14669 18377 14689
rect 18271 14653 18305 14664
rect 18271 14630 18273 14653
rect 18273 14630 18305 14653
rect 18343 14620 18377 14630
rect 18343 14596 18375 14620
rect 18375 14596 18377 14620
rect 18271 14584 18305 14591
rect 18271 14557 18273 14584
rect 18273 14557 18305 14584
rect 18343 14551 18377 14557
rect 18343 14523 18375 14551
rect 18375 14523 18377 14551
rect 18271 14515 18305 14518
rect 18271 14484 18273 14515
rect 18273 14484 18305 14515
rect 18343 14482 18377 14484
rect 18343 14450 18375 14482
rect 18375 14450 18377 14482
rect 18271 14412 18273 14445
rect 18273 14412 18305 14445
rect 18271 14411 18305 14412
rect 18343 14379 18375 14411
rect 18375 14379 18377 14411
rect 18271 14343 18273 14372
rect 18273 14343 18305 14372
rect 18343 14377 18377 14379
rect 18271 14338 18305 14343
rect 18343 14310 18375 14338
rect 18375 14310 18377 14338
rect 18271 14274 18273 14299
rect 18273 14274 18305 14299
rect 18343 14304 18377 14310
rect 18271 14265 18305 14274
rect 18343 14241 18375 14265
rect 18375 14241 18377 14265
rect 18271 14205 18273 14226
rect 18273 14205 18305 14226
rect 18343 14231 18377 14241
rect 18271 14192 18305 14205
rect 18343 14172 18375 14192
rect 18375 14172 18377 14192
rect 18271 14136 18273 14153
rect 18273 14136 18305 14153
rect 18343 14158 18377 14172
rect 18271 14119 18305 14136
rect 18343 14103 18375 14119
rect 18375 14103 18377 14119
rect 18271 14067 18273 14080
rect 18273 14067 18305 14080
rect 18343 14085 18377 14103
rect 18271 14046 18305 14067
rect 18343 14034 18375 14046
rect 18375 14034 18377 14046
rect 18271 13998 18273 14007
rect 18273 13998 18305 14007
rect 18343 14012 18377 14034
rect 18271 13973 18305 13998
rect 18343 13965 18375 13973
rect 18375 13965 18377 13973
rect 18271 13929 18273 13934
rect 18273 13929 18305 13934
rect 18343 13939 18377 13965
rect 18271 13900 18305 13929
rect 18343 13896 18375 13900
rect 18375 13896 18377 13900
rect 18343 13866 18377 13896
rect 18271 13860 18273 13861
rect 18273 13860 18305 13861
rect 18271 13827 18305 13860
rect 18343 13793 18377 13827
rect 18271 13756 18305 13788
rect 18271 13754 18273 13756
rect 18273 13754 18305 13756
rect 18343 13723 18377 13754
rect 18343 13720 18375 13723
rect 18375 13720 18377 13723
rect 18271 13687 18305 13715
rect 18271 13681 18273 13687
rect 18273 13681 18305 13687
rect 18343 13654 18377 13681
rect 18343 13647 18375 13654
rect 18375 13647 18377 13654
rect 18271 13618 18305 13642
rect 18271 13608 18273 13618
rect 18273 13608 18305 13618
rect 18343 13585 18377 13608
rect 18343 13574 18375 13585
rect 18375 13574 18377 13585
rect 18271 13549 18305 13569
rect 18271 13535 18273 13549
rect 18273 13535 18305 13549
rect 18343 13516 18377 13535
rect 18343 13501 18375 13516
rect 18375 13501 18377 13516
rect 18271 13480 18305 13496
rect 18271 13462 18273 13480
rect 18273 13462 18305 13480
rect 18343 13447 18377 13462
rect 18343 13428 18375 13447
rect 18375 13428 18377 13447
rect 18271 13411 18305 13423
rect 18271 13389 18273 13411
rect 18273 13389 18305 13411
rect 18343 13378 18377 13389
rect 18343 13355 18375 13378
rect 18375 13355 18377 13378
rect 18271 13342 18305 13350
rect 18271 13316 18273 13342
rect 18273 13316 18305 13342
rect 18343 13309 18377 13316
rect 18343 13282 18375 13309
rect 18375 13282 18377 13309
rect 18271 13273 18305 13277
rect 18271 13243 18273 13273
rect 18273 13243 18305 13273
rect 18343 13240 18377 13243
rect 18343 13209 18375 13240
rect 18375 13209 18377 13240
rect 18271 13170 18273 13204
rect 18273 13170 18305 13204
rect 18343 13137 18375 13170
rect 18375 13137 18377 13170
rect 18343 13136 18377 13137
rect 18271 13101 18273 13131
rect 18273 13101 18305 13131
rect 18271 13097 18305 13101
rect 18343 13068 18375 13097
rect 18375 13068 18377 13097
rect 18271 13032 18273 13058
rect 18273 13032 18305 13058
rect 18343 13063 18377 13068
rect 18271 13024 18305 13032
rect 18343 12999 18375 13024
rect 18375 12999 18377 13024
rect 18271 12963 18273 12985
rect 18273 12963 18305 12985
rect 18343 12990 18377 12999
rect 18271 12951 18305 12963
rect 18343 12930 18375 12951
rect 18375 12930 18377 12951
rect 18271 12894 18273 12912
rect 18273 12894 18305 12912
rect 18343 12917 18377 12930
rect 18271 12878 18305 12894
rect 18343 12861 18375 12878
rect 18375 12861 18377 12878
rect 18271 12825 18273 12839
rect 18273 12825 18305 12839
rect 18343 12844 18377 12861
rect 18271 12805 18305 12825
rect 357 12721 391 12755
rect 429 12721 463 12755
rect 357 12648 391 12682
rect 429 12648 463 12682
rect 18343 12792 18375 12805
rect 18375 12792 18377 12805
rect 18271 12756 18273 12766
rect 18273 12756 18305 12766
rect 18343 12771 18377 12792
rect 18271 12732 18305 12756
rect 18343 12723 18375 12732
rect 18375 12723 18377 12732
rect 18271 12687 18273 12693
rect 18273 12687 18305 12693
rect 18343 12698 18377 12723
rect 18271 12659 18305 12687
rect 18343 12654 18375 12659
rect 18375 12654 18377 12659
rect 2529 12618 2563 12623
rect 2602 12618 2632 12623
rect 2632 12618 2636 12623
rect 357 12575 391 12609
rect 429 12584 463 12609
rect 2529 12589 2563 12618
rect 2602 12589 2636 12618
rect 2675 12589 2709 12623
rect 2748 12589 2782 12623
rect 2821 12589 2855 12623
rect 2894 12589 2928 12623
rect 2967 12589 3001 12623
rect 3040 12589 3074 12623
rect 3113 12589 3147 12623
rect 3186 12589 3220 12623
rect 3259 12589 3293 12623
rect 3332 12589 3366 12623
rect 3405 12589 3439 12623
rect 3478 12589 3512 12623
rect 3551 12589 3585 12623
rect 3624 12589 3658 12623
rect 3697 12589 3731 12623
rect 429 12575 460 12584
rect 460 12575 463 12584
rect 2529 12550 2530 12551
rect 2530 12550 2563 12551
rect 357 12516 391 12536
rect 429 12516 463 12536
rect 2529 12517 2563 12550
rect 2602 12517 2636 12551
rect 2675 12517 2709 12551
rect 2748 12517 2782 12551
rect 2821 12517 2855 12551
rect 2894 12517 2928 12551
rect 2967 12517 3001 12551
rect 3040 12517 3074 12551
rect 3113 12517 3147 12551
rect 3186 12517 3220 12551
rect 3259 12517 3293 12551
rect 3332 12517 3366 12551
rect 3405 12517 3439 12551
rect 3478 12517 3512 12551
rect 3551 12517 3585 12551
rect 3624 12517 3658 12551
rect 3697 12517 3731 12551
rect 3770 12517 4236 12623
rect 6663 12589 6697 12623
rect 6736 12589 6770 12623
rect 6809 12589 6843 12623
rect 6882 12589 6916 12623
rect 6955 12589 6989 12623
rect 7028 12589 7062 12623
rect 7101 12589 7135 12623
rect 7174 12589 7208 12623
rect 7247 12589 7281 12623
rect 7320 12589 7354 12623
rect 7393 12589 7427 12623
rect 7466 12589 7500 12623
rect 7539 12589 7573 12623
rect 7612 12589 7646 12623
rect 7685 12589 7719 12623
rect 7758 12589 7792 12623
rect 7831 12589 7865 12623
rect 6663 12517 6697 12551
rect 6736 12517 6770 12551
rect 6809 12517 6843 12551
rect 6882 12517 6916 12551
rect 6955 12517 6989 12551
rect 7028 12517 7062 12551
rect 7101 12517 7135 12551
rect 7174 12517 7208 12551
rect 7247 12517 7281 12551
rect 7320 12517 7354 12551
rect 7393 12517 7427 12551
rect 7466 12517 7500 12551
rect 7539 12517 7573 12551
rect 7612 12517 7646 12551
rect 7685 12517 7719 12551
rect 7758 12517 7792 12551
rect 7831 12517 7865 12551
rect 7904 12517 8370 12623
rect 10790 12589 10824 12623
rect 10864 12589 10898 12623
rect 10938 12589 10972 12623
rect 11012 12589 11046 12623
rect 11086 12589 11120 12623
rect 11160 12589 11194 12623
rect 11233 12589 11267 12623
rect 11306 12589 11340 12623
rect 11379 12589 11413 12623
rect 11452 12589 11486 12623
rect 11525 12589 11559 12623
rect 11598 12589 11632 12623
rect 11671 12589 11705 12623
rect 11744 12589 11778 12623
rect 11817 12589 11851 12623
rect 11890 12589 11924 12623
rect 11963 12589 11997 12623
rect 12036 12589 12070 12623
rect 12109 12589 12143 12623
rect 12182 12589 12216 12623
rect 12255 12589 12289 12623
rect 12328 12589 12362 12623
rect 12401 12589 12435 12623
rect 12474 12589 12508 12623
rect 12547 12589 12581 12623
rect 12620 12589 12654 12623
rect 12693 12589 12727 12623
rect 12766 12589 12800 12623
rect 12839 12589 12873 12623
rect 12912 12589 12946 12623
rect 12985 12589 13019 12623
rect 13058 12589 13092 12623
rect 13131 12589 13165 12623
rect 13204 12589 13238 12623
rect 13277 12589 13311 12623
rect 13350 12589 13384 12623
rect 13423 12589 13457 12623
rect 13496 12589 13530 12623
rect 13569 12589 13603 12623
rect 13642 12589 13676 12623
rect 13715 12589 13749 12623
rect 13788 12589 13822 12623
rect 13861 12589 13895 12623
rect 13934 12589 13968 12623
rect 14007 12589 14041 12623
rect 14080 12589 14114 12623
rect 14153 12589 14187 12623
rect 14226 12589 14260 12623
rect 14299 12589 14333 12623
rect 14372 12589 14406 12623
rect 14445 12589 14479 12623
rect 14518 12589 14552 12623
rect 14591 12589 14625 12623
rect 14664 12589 14698 12623
rect 16036 12586 16070 12620
rect 16109 12586 16143 12620
rect 16182 12586 16216 12620
rect 16255 12586 16289 12620
rect 16327 12586 16361 12620
rect 16399 12586 16433 12620
rect 16471 12586 16505 12620
rect 16543 12586 16577 12620
rect 16615 12586 16649 12620
rect 16687 12586 16721 12620
rect 16759 12586 16793 12620
rect 16831 12586 16865 12620
rect 16903 12586 16937 12620
rect 16975 12586 17009 12620
rect 17047 12586 17081 12620
rect 17119 12586 17153 12620
rect 17191 12586 17225 12620
rect 17263 12586 17297 12620
rect 17335 12586 17369 12620
rect 17407 12586 17441 12620
rect 17479 12586 17513 12620
rect 17551 12586 17585 12620
rect 17623 12586 17657 12620
rect 17695 12586 17729 12620
rect 17767 12586 17801 12620
rect 17839 12586 17873 12620
rect 17911 12586 17945 12620
rect 17983 12586 18017 12620
rect 18055 12586 18089 12620
rect 18127 12586 18161 12620
rect 18199 12586 18233 12620
rect 18271 12586 18273 12620
rect 18273 12586 18305 12620
rect 18343 12625 18377 12654
rect 18343 12585 18375 12586
rect 18375 12585 18377 12586
rect 18343 12552 18377 12585
rect 10790 12517 10824 12551
rect 10864 12517 10898 12551
rect 10938 12517 10972 12551
rect 11012 12517 11046 12551
rect 11086 12517 11120 12551
rect 11160 12517 11194 12551
rect 11233 12517 11267 12551
rect 11306 12517 11340 12551
rect 11379 12517 11413 12551
rect 11452 12517 11486 12551
rect 11525 12517 11559 12551
rect 11598 12517 11632 12551
rect 11671 12517 11705 12551
rect 11744 12517 11778 12551
rect 11817 12517 11851 12551
rect 11890 12517 11924 12551
rect 11963 12517 11997 12551
rect 12036 12517 12070 12551
rect 12109 12517 12143 12551
rect 12182 12517 12216 12551
rect 12255 12517 12289 12551
rect 12328 12517 12362 12551
rect 12401 12517 12435 12551
rect 12474 12517 12508 12551
rect 12547 12517 12581 12551
rect 12620 12517 12654 12551
rect 12693 12517 12727 12551
rect 12766 12517 12800 12551
rect 12839 12517 12873 12551
rect 12912 12517 12946 12551
rect 12985 12517 13019 12551
rect 13058 12517 13092 12551
rect 13131 12517 13165 12551
rect 13204 12517 13238 12551
rect 13277 12517 13311 12551
rect 13350 12517 13384 12551
rect 13423 12517 13457 12551
rect 13496 12517 13530 12551
rect 13569 12517 13603 12551
rect 13642 12517 13676 12551
rect 13715 12517 13749 12551
rect 13788 12517 13822 12551
rect 13861 12517 13895 12551
rect 13934 12517 13968 12551
rect 14007 12517 14041 12551
rect 14080 12517 14114 12551
rect 14153 12517 14187 12551
rect 14226 12517 14260 12551
rect 14299 12517 14333 12551
rect 14372 12517 14406 12551
rect 14445 12517 14479 12551
rect 14518 12517 14552 12551
rect 14591 12517 14625 12551
rect 14664 12517 14698 12551
rect 357 12502 391 12516
rect 429 12502 460 12516
rect 460 12502 463 12516
rect 16036 12514 16070 12548
rect 16110 12514 16144 12548
rect 16184 12514 16218 12548
rect 16258 12514 16292 12548
rect 16332 12514 16366 12548
rect 16406 12514 16440 12548
rect 16479 12514 16513 12548
rect 16552 12514 16586 12548
rect 16625 12514 16659 12548
rect 16698 12514 16732 12548
rect 16771 12514 16805 12548
rect 16844 12514 16878 12548
rect 16917 12514 16951 12548
rect 16990 12514 17024 12548
rect 17063 12514 17097 12548
rect 17136 12514 17170 12548
rect 17209 12514 17243 12548
rect 17282 12514 17316 12548
rect 17355 12514 17389 12548
rect 17428 12514 17462 12548
rect 17501 12514 17535 12548
rect 17574 12514 17608 12548
rect 17647 12514 17681 12548
rect 17720 12514 17754 12548
rect 17793 12514 17827 12548
rect 17866 12514 17900 12548
rect 17939 12514 17973 12548
rect 18012 12514 18046 12548
rect 18085 12514 18119 12548
rect 18158 12514 18192 12548
rect 18231 12514 18265 12548
rect 17016 7625 17050 7659
rect 10167 3622 10201 3656
rect 10239 3588 10271 3622
rect 10271 3588 10273 3622
rect 10277 3588 11785 3694
rect 11789 3660 11823 3694
rect 11861 3660 11895 3694
rect 11933 3660 11967 3694
rect 12005 3660 12039 3694
rect 12077 3660 12111 3694
rect 12150 3660 12184 3694
rect 12223 3660 12257 3694
rect 12296 3660 12330 3694
rect 12369 3660 12403 3694
rect 12442 3660 12476 3694
rect 12515 3660 12549 3694
rect 12588 3660 12622 3694
rect 12661 3660 12695 3694
rect 12734 3660 12768 3694
rect 12807 3660 12841 3694
rect 12880 3660 12914 3694
rect 12953 3660 12987 3694
rect 13026 3660 13060 3694
rect 13099 3660 13133 3694
rect 13172 3660 13206 3694
rect 13245 3660 13279 3694
rect 13318 3660 13352 3694
rect 13391 3660 13425 3694
rect 13464 3660 13498 3694
rect 13537 3660 13571 3694
rect 13610 3660 13644 3694
rect 13683 3660 13717 3694
rect 13756 3660 13790 3694
rect 13829 3660 13863 3694
rect 13902 3660 13936 3694
rect 13975 3660 14009 3694
rect 14048 3660 14082 3694
rect 14121 3660 14155 3694
rect 14194 3660 14228 3694
rect 14267 3660 14301 3694
rect 14340 3660 14374 3694
rect 14413 3660 14447 3694
rect 14486 3660 14520 3694
rect 14559 3692 14590 3694
rect 14590 3692 14593 3694
rect 14632 3692 14659 3694
rect 14659 3692 14666 3694
rect 14705 3692 14728 3694
rect 14728 3692 14739 3694
rect 14778 3692 14797 3694
rect 14797 3692 14812 3694
rect 14851 3692 14866 3694
rect 14866 3692 14885 3694
rect 14924 3692 14935 3694
rect 14935 3692 14958 3694
rect 14997 3692 15004 3694
rect 15004 3692 15031 3694
rect 15070 3692 15073 3694
rect 15073 3692 15104 3694
rect 15143 3692 15176 3694
rect 15176 3692 15177 3694
rect 15216 3692 15245 3694
rect 15245 3692 15250 3694
rect 15289 3692 15314 3694
rect 15314 3692 15323 3694
rect 15362 3692 15383 3694
rect 15383 3692 15396 3694
rect 15435 3692 15452 3694
rect 15452 3692 15469 3694
rect 15508 3692 15521 3694
rect 15521 3692 15542 3694
rect 15581 3692 15590 3694
rect 15590 3692 15615 3694
rect 15654 3692 15659 3694
rect 15659 3692 15688 3694
rect 15727 3692 15728 3694
rect 15728 3692 15761 3694
rect 14559 3660 14593 3692
rect 14632 3660 14666 3692
rect 14705 3660 14739 3692
rect 14778 3660 14812 3692
rect 14851 3660 14885 3692
rect 14924 3660 14958 3692
rect 14997 3660 15031 3692
rect 15070 3660 15104 3692
rect 15143 3660 15177 3692
rect 15216 3660 15250 3692
rect 15289 3660 15323 3692
rect 15362 3660 15396 3692
rect 15435 3660 15469 3692
rect 15508 3660 15542 3692
rect 15581 3660 15615 3692
rect 15654 3660 15688 3692
rect 15727 3660 15761 3692
rect 11824 3588 11858 3622
rect 11897 3588 11931 3622
rect 11970 3588 12004 3622
rect 12043 3588 12077 3622
rect 12116 3588 12150 3622
rect 12189 3588 12223 3622
rect 12262 3588 12296 3622
rect 12335 3588 12369 3622
rect 12408 3588 12442 3622
rect 12481 3588 12515 3622
rect 12554 3588 12588 3622
rect 12627 3588 12661 3622
rect 12700 3588 12734 3622
rect 12773 3588 12807 3622
rect 12846 3588 12880 3622
rect 12919 3588 12953 3622
rect 12992 3588 13026 3622
rect 13065 3588 13099 3622
rect 13138 3588 13172 3622
rect 13211 3588 13245 3622
rect 13284 3588 13318 3622
rect 13357 3588 13391 3622
rect 13430 3588 13464 3622
rect 13503 3588 13537 3622
rect 13576 3588 13610 3622
rect 13649 3588 13683 3622
rect 13722 3588 13756 3622
rect 13795 3588 13829 3622
rect 13868 3588 13902 3622
rect 13941 3588 13975 3622
rect 14014 3588 14048 3622
rect 14087 3588 14121 3622
rect 14160 3588 14194 3622
rect 14233 3588 14267 3622
rect 14306 3588 14340 3622
rect 14379 3588 14413 3622
rect 14452 3588 14453 3622
rect 14453 3588 14486 3622
rect 14525 3590 14559 3622
rect 14598 3590 14632 3622
rect 14671 3590 14705 3622
rect 14744 3590 14778 3622
rect 14817 3590 14851 3622
rect 14890 3590 14924 3622
rect 14963 3590 14997 3622
rect 15036 3590 15070 3622
rect 15109 3590 15143 3622
rect 15182 3590 15216 3622
rect 15255 3590 15289 3622
rect 15328 3590 15362 3622
rect 15401 3590 15435 3622
rect 15474 3590 15508 3622
rect 15547 3590 15581 3622
rect 15620 3590 15654 3622
rect 15693 3590 15727 3622
rect 10167 3543 10201 3576
rect 14525 3588 14557 3590
rect 14557 3588 14559 3590
rect 14598 3588 14626 3590
rect 14626 3588 14632 3590
rect 14671 3588 14695 3590
rect 14695 3588 14705 3590
rect 14744 3588 14764 3590
rect 14764 3588 14778 3590
rect 14817 3588 14833 3590
rect 14833 3588 14851 3590
rect 14890 3588 14902 3590
rect 14902 3588 14924 3590
rect 14963 3588 14971 3590
rect 14971 3588 14997 3590
rect 15036 3588 15040 3590
rect 15040 3588 15070 3590
rect 15109 3588 15143 3590
rect 15182 3588 15212 3590
rect 15212 3588 15216 3590
rect 15255 3588 15281 3590
rect 15281 3588 15289 3590
rect 15328 3588 15350 3590
rect 15350 3588 15362 3590
rect 15401 3588 15419 3590
rect 15419 3588 15435 3590
rect 15474 3588 15488 3590
rect 15488 3588 15508 3590
rect 15547 3588 15557 3590
rect 15557 3588 15581 3590
rect 15620 3588 15626 3590
rect 15626 3588 15654 3590
rect 15693 3588 15695 3590
rect 15695 3588 15727 3590
rect 10167 3542 10169 3543
rect 10169 3542 10201 3543
rect 10239 3519 10273 3546
rect 10167 3469 10201 3497
rect 10239 3512 10271 3519
rect 10271 3512 10273 3519
rect 10167 3463 10169 3469
rect 10169 3463 10201 3469
rect 10239 3448 10273 3470
rect 10167 3395 10201 3418
rect 10239 3436 10271 3448
rect 10271 3436 10273 3448
rect 10167 3384 10169 3395
rect 10169 3384 10201 3395
rect 15765 3556 15799 3582
rect 15693 3521 15727 3550
rect 15765 3548 15797 3556
rect 15797 3548 15799 3556
rect 15693 3516 15695 3521
rect 15695 3516 15727 3521
rect 15765 3488 15799 3509
rect 15693 3452 15727 3478
rect 15765 3475 15797 3488
rect 15797 3475 15799 3488
rect 15693 3444 15695 3452
rect 15695 3444 15727 3452
rect 15765 3420 15799 3436
rect 10239 3377 10273 3394
rect 10239 3360 10271 3377
rect 10271 3360 10273 3377
rect 10167 3321 10201 3339
rect 10167 3305 10169 3321
rect 10169 3305 10201 3321
rect 10239 3306 10273 3319
rect 10239 3285 10271 3306
rect 10271 3285 10273 3306
rect 10167 3247 10201 3260
rect 10167 3226 10169 3247
rect 10169 3226 10201 3247
rect 10239 3235 10273 3244
rect 10239 3210 10271 3235
rect 10271 3210 10273 3235
rect 10167 3173 10201 3181
rect 10167 3147 10169 3173
rect 10169 3147 10201 3173
rect 10239 3164 10273 3169
rect 10239 3135 10271 3164
rect 10271 3135 10273 3164
rect 10167 3099 10201 3102
rect 10167 3068 10169 3099
rect 10169 3068 10201 3099
rect 10239 3093 10273 3094
rect 10239 3060 10271 3093
rect 10271 3060 10273 3093
rect 10167 2991 10169 3023
rect 10169 2991 10201 3023
rect 10167 2989 10201 2991
rect 10239 2988 10271 3019
rect 10271 2988 10273 3019
rect 10239 2985 10273 2988
rect 10167 2917 10169 2944
rect 10169 2917 10201 2944
rect 10239 2917 10271 2944
rect 10271 2917 10273 2944
rect 10167 2910 10201 2917
rect 10239 2910 10273 2917
rect 10633 3346 10661 3373
rect 10661 3346 10737 3373
rect 10523 3310 10557 3335
rect 10633 3311 10737 3346
rect 10523 3301 10525 3310
rect 10525 3301 10557 3310
rect 10595 3277 10627 3301
rect 10627 3277 10629 3301
rect 10633 3277 10661 3311
rect 10661 3277 10737 3311
rect 10737 3302 12267 3373
rect 12267 3370 12301 3373
rect 12301 3370 12335 3373
rect 12335 3370 12369 3373
rect 12369 3370 12403 3373
rect 12403 3370 12437 3373
rect 12437 3370 12471 3373
rect 12471 3370 12505 3373
rect 12505 3370 12539 3373
rect 12539 3370 12573 3373
rect 12573 3370 12607 3373
rect 12607 3370 12641 3373
rect 12641 3370 12675 3373
rect 12675 3370 12709 3373
rect 12709 3370 12743 3373
rect 12743 3370 12777 3373
rect 12777 3370 12811 3373
rect 12811 3370 12845 3373
rect 12845 3370 12879 3373
rect 12879 3370 12913 3373
rect 12913 3370 12947 3373
rect 12947 3370 12981 3373
rect 12981 3370 13015 3373
rect 13015 3370 13049 3373
rect 13049 3370 13083 3373
rect 13083 3370 13117 3373
rect 13117 3370 13151 3373
rect 13151 3370 13185 3373
rect 13185 3370 13219 3373
rect 13219 3370 13253 3373
rect 13253 3370 13287 3373
rect 13287 3370 13321 3373
rect 13321 3370 13355 3373
rect 13355 3370 13389 3373
rect 13389 3370 13423 3373
rect 13423 3370 13457 3373
rect 13457 3370 13491 3373
rect 13491 3370 13525 3373
rect 13525 3370 13559 3373
rect 13559 3370 13593 3373
rect 13593 3370 13627 3373
rect 13627 3370 13653 3373
rect 12267 3336 13653 3370
rect 13657 3370 13661 3373
rect 13661 3370 13691 3373
rect 13729 3370 13763 3373
rect 13801 3370 13831 3373
rect 13831 3370 13835 3373
rect 13873 3370 13899 3373
rect 13899 3370 13907 3373
rect 13945 3370 13967 3373
rect 13967 3370 13979 3373
rect 14018 3370 14035 3373
rect 14035 3370 14052 3373
rect 14091 3370 14103 3373
rect 14103 3370 14125 3373
rect 14164 3370 14171 3373
rect 14171 3370 14198 3373
rect 14237 3370 14239 3373
rect 14239 3370 14271 3373
rect 14310 3370 14341 3373
rect 14341 3370 14344 3373
rect 14383 3370 14409 3373
rect 14409 3370 14417 3373
rect 14456 3370 14477 3373
rect 14477 3370 14490 3373
rect 14529 3370 14545 3373
rect 14545 3370 14563 3373
rect 14602 3370 14613 3373
rect 14613 3370 14636 3373
rect 14675 3370 14682 3373
rect 14682 3370 14709 3373
rect 14748 3370 14751 3373
rect 14751 3370 14782 3373
rect 14821 3370 14854 3373
rect 14854 3370 14855 3373
rect 14894 3370 14923 3373
rect 14923 3370 14928 3373
rect 14967 3370 14992 3373
rect 14992 3370 15001 3373
rect 15040 3370 15061 3373
rect 15061 3370 15074 3373
rect 15113 3370 15130 3373
rect 15130 3370 15147 3373
rect 15186 3370 15199 3373
rect 15199 3370 15220 3373
rect 15259 3370 15268 3373
rect 15268 3370 15293 3373
rect 15332 3370 15337 3373
rect 15337 3370 15366 3373
rect 15405 3370 15406 3373
rect 15406 3370 15439 3373
rect 13657 3339 13691 3370
rect 13729 3339 13763 3370
rect 13801 3339 13835 3370
rect 13873 3339 13907 3370
rect 13945 3339 13979 3370
rect 14018 3339 14052 3370
rect 14091 3339 14125 3370
rect 14164 3339 14198 3370
rect 14237 3339 14271 3370
rect 14310 3339 14344 3370
rect 14383 3339 14417 3370
rect 14456 3339 14490 3370
rect 14529 3339 14563 3370
rect 14602 3339 14636 3370
rect 14675 3339 14709 3370
rect 14748 3339 14782 3370
rect 14821 3339 14855 3370
rect 14894 3339 14928 3370
rect 14967 3339 15001 3370
rect 15040 3339 15074 3370
rect 15113 3339 15147 3370
rect 15186 3339 15220 3370
rect 15259 3339 15293 3370
rect 15332 3339 15366 3370
rect 15405 3339 15439 3370
rect 12267 3302 12302 3336
rect 12302 3302 12336 3336
rect 12336 3302 12371 3336
rect 12371 3302 12405 3336
rect 12405 3302 12440 3336
rect 12440 3302 12474 3336
rect 12474 3302 12509 3336
rect 12509 3302 12543 3336
rect 12543 3302 12578 3336
rect 12578 3302 12612 3336
rect 12612 3302 12647 3336
rect 12647 3302 12681 3336
rect 12681 3302 12716 3336
rect 12716 3302 12750 3336
rect 12750 3302 12785 3336
rect 12785 3302 12819 3336
rect 12819 3302 12854 3336
rect 12854 3302 12888 3336
rect 12888 3302 12923 3336
rect 12923 3302 12957 3336
rect 12957 3302 12992 3336
rect 12992 3302 13026 3336
rect 13026 3302 13061 3336
rect 13061 3302 13095 3336
rect 13095 3302 13130 3336
rect 13130 3302 13164 3336
rect 13164 3302 13199 3336
rect 13199 3302 13233 3336
rect 13233 3302 13268 3336
rect 13268 3302 13302 3336
rect 13302 3302 13337 3336
rect 13337 3302 13371 3336
rect 13371 3302 13406 3336
rect 13406 3302 13440 3336
rect 13440 3302 13475 3336
rect 13475 3302 13509 3336
rect 13509 3302 13544 3336
rect 13544 3302 13578 3336
rect 13578 3302 13613 3336
rect 13613 3302 13647 3336
rect 13647 3302 13653 3336
rect 10595 3267 10629 3277
rect 10633 3267 10737 3277
rect 10737 3267 12199 3302
rect 12199 3268 13653 3302
rect 13692 3268 13726 3301
rect 13765 3268 13799 3301
rect 13838 3268 13872 3301
rect 13911 3268 13945 3301
rect 13984 3268 14018 3301
rect 14057 3268 14091 3301
rect 14130 3268 14164 3301
rect 14203 3268 14237 3301
rect 14276 3268 14310 3301
rect 14349 3268 14383 3301
rect 14422 3268 14456 3301
rect 14495 3268 14529 3301
rect 14568 3268 14602 3301
rect 14641 3268 14675 3301
rect 14714 3268 14748 3301
rect 14787 3268 14821 3301
rect 14860 3268 14894 3301
rect 14933 3268 14967 3301
rect 15006 3268 15040 3301
rect 15079 3268 15113 3301
rect 15152 3268 15186 3301
rect 15225 3268 15259 3301
rect 15298 3268 15332 3301
rect 15371 3268 15405 3301
rect 12199 3267 12234 3268
rect 12234 3267 12268 3268
rect 12268 3267 12303 3268
rect 12303 3267 12337 3268
rect 12337 3267 12372 3268
rect 12372 3267 12406 3268
rect 12406 3267 12441 3268
rect 12441 3267 12475 3268
rect 12475 3267 12510 3268
rect 12510 3267 12544 3268
rect 12544 3267 12579 3268
rect 12579 3267 12613 3268
rect 12613 3267 12648 3268
rect 12648 3267 12682 3268
rect 12682 3267 12717 3268
rect 12717 3267 12751 3268
rect 12751 3267 12786 3268
rect 12786 3267 12820 3268
rect 12820 3267 12855 3268
rect 12855 3267 12889 3268
rect 12889 3267 12924 3268
rect 12924 3267 12958 3268
rect 12958 3267 12993 3268
rect 12993 3267 13027 3268
rect 13027 3267 13062 3268
rect 13062 3267 13096 3268
rect 13096 3267 13131 3268
rect 13131 3267 13165 3268
rect 13165 3267 13200 3268
rect 13200 3267 13234 3268
rect 13234 3267 13269 3268
rect 13269 3267 13303 3268
rect 13303 3267 13338 3268
rect 13338 3267 13372 3268
rect 13372 3267 13407 3268
rect 13407 3267 13441 3268
rect 13441 3267 13476 3268
rect 13476 3267 13510 3268
rect 13510 3267 13545 3268
rect 13545 3267 13579 3268
rect 13579 3267 13614 3268
rect 13614 3267 13648 3268
rect 13648 3267 13653 3268
rect 13692 3267 13717 3268
rect 13717 3267 13726 3268
rect 13765 3267 13786 3268
rect 13786 3267 13799 3268
rect 13838 3267 13855 3268
rect 13855 3267 13872 3268
rect 13911 3267 13924 3268
rect 13924 3267 13945 3268
rect 13984 3267 13993 3268
rect 13993 3267 14018 3268
rect 14057 3267 14062 3268
rect 14062 3267 14091 3268
rect 14130 3267 14131 3268
rect 14131 3267 14164 3268
rect 10523 3240 10557 3262
rect 10523 3228 10525 3240
rect 10525 3228 10557 3240
rect 14203 3267 14235 3268
rect 14235 3267 14237 3268
rect 14276 3267 14304 3268
rect 14304 3267 14310 3268
rect 14349 3267 14373 3268
rect 14373 3267 14383 3268
rect 14422 3267 14442 3268
rect 14442 3267 14456 3268
rect 14495 3267 14511 3268
rect 14511 3267 14529 3268
rect 14568 3267 14580 3268
rect 14580 3267 14602 3268
rect 14641 3267 14649 3268
rect 14649 3267 14675 3268
rect 14714 3267 14718 3268
rect 14718 3267 14748 3268
rect 14787 3267 14821 3268
rect 14860 3267 14890 3268
rect 14890 3267 14894 3268
rect 14933 3267 14959 3268
rect 14959 3267 14967 3268
rect 15006 3267 15028 3268
rect 15028 3267 15040 3268
rect 15079 3267 15097 3268
rect 15097 3267 15113 3268
rect 15152 3267 15166 3268
rect 15166 3267 15186 3268
rect 15225 3267 15235 3268
rect 15235 3267 15259 3268
rect 15298 3267 15304 3268
rect 15304 3267 15332 3268
rect 15371 3267 15373 3268
rect 15373 3267 15405 3268
rect 10595 3208 10627 3227
rect 10627 3208 10629 3227
rect 10595 3193 10629 3208
rect 10523 3170 10557 3189
rect 10523 3155 10525 3170
rect 10525 3155 10557 3170
rect 10595 3139 10627 3153
rect 10627 3139 10629 3153
rect 10595 3119 10629 3139
rect 10523 3100 10557 3116
rect 10523 3082 10525 3100
rect 10525 3082 10557 3100
rect 10595 3070 10627 3079
rect 10627 3070 10629 3079
rect 10595 3045 10629 3070
rect 10523 3030 10557 3043
rect 10523 3009 10525 3030
rect 10525 3009 10557 3030
rect 10595 3001 10627 3005
rect 10627 3001 10629 3005
rect 10595 2971 10629 3001
rect 10523 2960 10557 2970
rect 10523 2936 10525 2960
rect 10525 2936 10557 2960
rect 10523 2890 10557 2898
rect 10595 2897 10629 2931
rect 10523 2864 10525 2890
rect 10525 2864 10557 2890
rect 10595 2828 10629 2857
rect 10523 2820 10557 2826
rect 10523 2792 10525 2820
rect 10525 2792 10557 2820
rect 10595 2823 10627 2828
rect 10627 2823 10629 2828
rect 10595 2759 10629 2783
rect 10523 2750 10557 2754
rect 10523 2720 10525 2750
rect 10525 2720 10557 2750
rect 10595 2749 10627 2759
rect 10627 2749 10629 2759
rect 10595 2690 10629 2709
rect 10523 2680 10557 2682
rect 10523 2648 10525 2680
rect 10525 2648 10557 2680
rect 10595 2675 10627 2690
rect 10627 2675 10629 2690
rect 10595 2621 10629 2636
rect 10523 2576 10525 2610
rect 10525 2576 10557 2610
rect 10595 2602 10627 2621
rect 10627 2602 10629 2621
rect 10595 2552 10629 2563
rect 10523 2506 10525 2538
rect 10525 2506 10557 2538
rect 10595 2529 10627 2552
rect 10627 2529 10629 2552
rect 10523 2504 10557 2506
rect 10595 2483 10629 2490
rect 10523 2436 10525 2466
rect 10525 2436 10557 2466
rect 10595 2456 10627 2483
rect 10627 2456 10629 2483
rect 10523 2432 10557 2436
rect 10595 2414 10629 2417
rect 10523 2366 10525 2394
rect 10525 2366 10557 2394
rect 10595 2383 10627 2414
rect 10627 2383 10629 2414
rect 15443 3231 15477 3261
rect 15371 3199 15405 3228
rect 15443 3227 15475 3231
rect 15475 3227 15477 3231
rect 15371 3194 15373 3199
rect 15373 3194 15405 3199
rect 15443 3162 15477 3188
rect 15371 3130 15405 3155
rect 15443 3154 15475 3162
rect 15475 3154 15477 3162
rect 15371 3121 15373 3130
rect 15373 3121 15405 3130
rect 15443 3093 15477 3115
rect 15371 3061 15405 3082
rect 15443 3081 15475 3093
rect 15475 3081 15477 3093
rect 15371 3048 15373 3061
rect 15373 3048 15405 3061
rect 15443 3024 15477 3042
rect 15371 2992 15405 3009
rect 15443 3008 15475 3024
rect 15475 3008 15477 3024
rect 15371 2975 15373 2992
rect 15373 2975 15405 2992
rect 15443 2955 15477 2969
rect 15371 2923 15405 2936
rect 15443 2935 15475 2955
rect 15475 2935 15477 2955
rect 15371 2902 15373 2923
rect 15373 2902 15405 2923
rect 15443 2886 15477 2896
rect 15371 2854 15405 2863
rect 15443 2862 15475 2886
rect 15475 2862 15477 2886
rect 15371 2829 15373 2854
rect 15373 2829 15405 2854
rect 15443 2817 15477 2823
rect 15371 2785 15405 2790
rect 15443 2789 15475 2817
rect 15475 2789 15477 2817
rect 15371 2756 15373 2785
rect 15373 2756 15405 2785
rect 15443 2748 15477 2750
rect 15371 2716 15405 2717
rect 15443 2716 15475 2748
rect 15475 2716 15477 2748
rect 15371 2683 15373 2716
rect 15373 2683 15405 2716
rect 15371 2613 15373 2644
rect 15373 2613 15405 2644
rect 15371 2610 15405 2613
rect 15443 2645 15475 2677
rect 15475 2645 15477 2677
rect 15443 2643 15477 2645
rect 15371 2544 15373 2571
rect 15373 2544 15405 2571
rect 15371 2537 15405 2544
rect 15443 2576 15475 2604
rect 15475 2576 15477 2604
rect 15443 2570 15477 2576
rect 15371 2475 15373 2498
rect 15373 2475 15405 2498
rect 15371 2464 15405 2475
rect 15443 2507 15475 2531
rect 15475 2507 15477 2531
rect 15443 2497 15477 2507
rect 15371 2406 15373 2425
rect 15373 2406 15405 2425
rect 10523 2360 10557 2366
rect 10523 2296 10525 2322
rect 10525 2296 10557 2322
rect 10595 2311 10627 2344
rect 10627 2311 10629 2344
rect 10595 2310 10629 2311
rect 10523 2288 10557 2296
rect 10523 2226 10525 2250
rect 10525 2226 10557 2250
rect 10595 2242 10627 2271
rect 10627 2242 10629 2271
rect 10595 2237 10629 2242
rect 10523 2216 10557 2226
rect 10523 2156 10525 2178
rect 10525 2156 10557 2178
rect 10595 2173 10627 2198
rect 10627 2173 10629 2198
rect 10595 2164 10629 2173
rect 10523 2144 10557 2156
rect 10523 2086 10525 2106
rect 10525 2086 10557 2106
rect 10595 2104 10627 2125
rect 10627 2104 10629 2125
rect 10595 2091 10629 2104
rect 10523 2072 10557 2086
rect 10595 2035 10627 2052
rect 10627 2035 10629 2052
rect 10523 2016 10525 2034
rect 10525 2016 10557 2034
rect 10595 2018 10629 2035
rect 10523 2000 10557 2016
rect 10595 1966 10627 1979
rect 10627 1966 10629 1979
rect 10523 1946 10525 1962
rect 10525 1946 10557 1962
rect 10523 1928 10557 1946
rect 10595 1945 10629 1966
rect 10595 1897 10627 1906
rect 10627 1897 10629 1906
rect 10523 1876 10525 1890
rect 10525 1876 10557 1890
rect 10523 1856 10557 1876
rect 10595 1872 10629 1897
rect 10595 1828 10627 1833
rect 10627 1828 10629 1833
rect 10523 1806 10525 1818
rect 10525 1806 10557 1818
rect 10523 1784 10557 1806
rect 10595 1799 10629 1828
rect 10595 1759 10627 1760
rect 10627 1759 10629 1760
rect 10523 1736 10525 1746
rect 10525 1736 10557 1746
rect 10523 1712 10557 1736
rect 10595 1726 10629 1759
rect 10523 1667 10525 1674
rect 10525 1667 10557 1674
rect 10523 1640 10557 1667
rect 10595 1655 10629 1687
rect 10595 1653 10627 1655
rect 10627 1653 10629 1655
rect 10523 1598 10525 1602
rect 10525 1598 10557 1602
rect 10523 1568 10557 1598
rect 10595 1586 10629 1614
rect 10595 1580 10627 1586
rect 10627 1580 10629 1586
rect 10523 1529 10525 1530
rect 10525 1529 10557 1530
rect 10523 1496 10557 1529
rect 10595 1517 10629 1541
rect 10709 2372 10743 2406
rect 10709 2296 10743 2330
rect 10709 2219 10743 2253
rect 10709 2142 10743 2176
rect 15257 2372 15291 2406
rect 15257 2296 15291 2330
rect 15257 2219 15291 2253
rect 15257 2142 15291 2176
rect 10709 2065 10743 2099
rect 10709 1988 10743 2022
rect 12951 2012 13057 2118
rect 15257 2065 15291 2099
rect 10709 1911 10743 1945
rect 15257 1988 15291 2022
rect 15257 1911 15291 1945
rect 10709 1834 10743 1868
rect 12951 1801 13057 1907
rect 15257 1834 15291 1868
rect 10709 1757 10743 1791
rect 10709 1680 10743 1714
rect 10709 1603 10743 1637
rect 10709 1526 10743 1560
rect 15257 1757 15291 1791
rect 15257 1680 15291 1714
rect 15257 1603 15291 1637
rect 15257 1526 15291 1560
rect 15371 2391 15405 2406
rect 15443 2438 15475 2458
rect 15475 2438 15477 2458
rect 15443 2424 15477 2438
rect 15371 2337 15373 2352
rect 15373 2337 15405 2352
rect 15371 2318 15405 2337
rect 15443 2369 15475 2385
rect 15475 2369 15477 2385
rect 15443 2351 15477 2369
rect 15371 2268 15373 2279
rect 15373 2268 15405 2279
rect 15371 2245 15405 2268
rect 15443 2300 15475 2312
rect 15475 2300 15477 2312
rect 15443 2278 15477 2300
rect 15371 2199 15373 2206
rect 15373 2199 15405 2206
rect 15371 2172 15405 2199
rect 15443 2231 15475 2239
rect 15475 2231 15477 2239
rect 15443 2205 15477 2231
rect 15371 2130 15373 2133
rect 15373 2130 15405 2133
rect 15371 2099 15405 2130
rect 15443 2162 15475 2166
rect 15475 2162 15477 2166
rect 15443 2132 15477 2162
rect 15371 2026 15405 2060
rect 15443 2059 15477 2093
rect 15443 1989 15477 2020
rect 15371 1957 15405 1987
rect 15443 1986 15475 1989
rect 15475 1986 15477 1989
rect 15371 1953 15373 1957
rect 15373 1953 15405 1957
rect 15443 1920 15477 1947
rect 15371 1888 15405 1914
rect 15443 1913 15475 1920
rect 15475 1913 15477 1920
rect 15371 1880 15373 1888
rect 15373 1880 15405 1888
rect 15443 1851 15477 1874
rect 15371 1818 15405 1841
rect 15443 1840 15475 1851
rect 15475 1840 15477 1851
rect 15371 1807 15373 1818
rect 15373 1807 15405 1818
rect 15443 1782 15477 1801
rect 15371 1748 15405 1768
rect 15443 1767 15475 1782
rect 15475 1767 15477 1782
rect 15371 1734 15373 1748
rect 15373 1734 15405 1748
rect 15443 1713 15477 1728
rect 15371 1678 15405 1695
rect 15443 1694 15475 1713
rect 15475 1694 15477 1713
rect 15371 1661 15373 1678
rect 15373 1661 15405 1678
rect 15443 1644 15477 1655
rect 15371 1608 15405 1622
rect 15443 1621 15475 1644
rect 15475 1621 15477 1644
rect 15371 1588 15373 1608
rect 15373 1588 15405 1608
rect 15443 1575 15477 1582
rect 15371 1538 15405 1549
rect 15443 1548 15475 1575
rect 15475 1548 15477 1575
rect 10595 1507 10627 1517
rect 10627 1507 10629 1517
rect 10523 1425 10557 1458
rect 10595 1448 10629 1468
rect 10523 1424 10525 1425
rect 10525 1424 10557 1425
rect 10595 1434 10627 1448
rect 10627 1434 10629 1448
rect 10523 1356 10557 1386
rect 10595 1379 10629 1395
rect 10523 1352 10525 1356
rect 10525 1352 10557 1356
rect 10595 1361 10627 1379
rect 10627 1361 10629 1379
rect 10523 1287 10557 1314
rect 10595 1310 10629 1322
rect 10523 1280 10525 1287
rect 10525 1280 10557 1287
rect 10595 1288 10629 1310
rect 10523 1218 10557 1242
rect 10523 1208 10525 1218
rect 10525 1208 10557 1218
rect 10595 1215 10629 1249
rect 10523 1149 10557 1170
rect 10523 1136 10525 1149
rect 10525 1136 10557 1149
rect 10595 1142 10629 1176
rect 10523 1080 10557 1098
rect 10523 1064 10525 1080
rect 10525 1064 10557 1080
rect 10595 1069 10629 1103
rect 10523 1011 10557 1026
rect 10523 992 10525 1011
rect 10525 992 10557 1011
rect 10595 996 10629 1030
rect 10523 942 10557 954
rect 10523 920 10525 942
rect 10525 920 10557 942
rect 10595 923 10629 957
rect 10523 873 10557 882
rect 10523 848 10525 873
rect 10525 848 10557 873
rect 10595 850 10629 884
rect 10523 804 10557 810
rect 10523 776 10525 804
rect 10525 776 10557 804
rect 10595 777 10629 811
rect 10523 735 10557 738
rect 10523 704 10525 735
rect 10525 704 10557 735
rect 10595 704 10629 738
rect 15371 1515 15373 1538
rect 15373 1515 15405 1538
rect 15443 1506 15477 1509
rect 15371 1468 15405 1476
rect 15443 1475 15475 1506
rect 15475 1475 15477 1506
rect 15371 1442 15373 1468
rect 15373 1442 15405 1468
rect 15371 1398 15405 1403
rect 15443 1402 15475 1436
rect 15475 1402 15477 1436
rect 15371 1369 15373 1398
rect 15373 1369 15405 1398
rect 15443 1332 15475 1363
rect 15475 1332 15477 1363
rect 15371 1328 15405 1330
rect 15371 1296 15373 1328
rect 15373 1296 15405 1328
rect 15443 1329 15477 1332
rect 15443 1262 15475 1290
rect 15475 1262 15477 1290
rect 15371 1224 15373 1257
rect 15373 1224 15405 1257
rect 15443 1256 15477 1262
rect 15371 1223 15405 1224
rect 15443 1192 15475 1217
rect 15475 1192 15477 1217
rect 15371 1154 15373 1183
rect 15373 1154 15405 1183
rect 15443 1183 15477 1192
rect 15371 1149 15405 1154
rect 15443 1122 15475 1144
rect 15475 1122 15477 1144
rect 15371 1084 15373 1109
rect 15373 1084 15405 1109
rect 15443 1110 15477 1122
rect 15371 1075 15405 1084
rect 15443 1052 15475 1071
rect 15475 1052 15477 1071
rect 15371 1014 15373 1035
rect 15373 1014 15405 1035
rect 15443 1037 15477 1052
rect 15371 1001 15405 1014
rect 15443 982 15475 998
rect 15475 982 15477 998
rect 15371 944 15373 961
rect 15373 944 15405 961
rect 15443 964 15477 982
rect 15371 927 15405 944
rect 15443 912 15475 925
rect 15475 912 15477 925
rect 15371 874 15373 887
rect 15373 874 15405 887
rect 15443 891 15477 912
rect 15371 853 15405 874
rect 15443 842 15475 852
rect 15475 842 15477 852
rect 15371 804 15373 813
rect 15373 804 15405 813
rect 15443 818 15477 842
rect 15371 779 15405 804
rect 15443 772 15475 779
rect 15475 772 15477 779
rect 15371 734 15373 739
rect 15373 734 15405 739
rect 15443 745 15477 772
rect 15371 705 15405 734
rect 15443 702 15475 705
rect 15475 702 15477 705
rect 10529 664 10559 665
rect 10559 664 10563 665
rect 10602 664 10636 665
rect 10675 664 10696 665
rect 10696 664 10709 665
rect 10748 664 10765 665
rect 10765 664 10782 665
rect 10821 664 10834 665
rect 10834 664 10855 665
rect 10894 664 10903 665
rect 10903 664 10928 665
rect 10967 664 10972 665
rect 10972 664 11001 665
rect 11040 664 11041 665
rect 11041 664 11074 665
rect 11113 664 11144 665
rect 11144 664 11147 665
rect 11186 664 11213 665
rect 11213 664 11220 665
rect 11259 664 11282 665
rect 11282 664 11293 665
rect 11332 664 11351 665
rect 11351 664 11366 665
rect 11405 664 11420 665
rect 11420 664 11439 665
rect 11478 664 11489 665
rect 11489 664 11512 665
rect 11551 664 11558 665
rect 11558 664 11585 665
rect 11624 664 11627 665
rect 11627 664 11658 665
rect 10529 631 10563 664
rect 10602 631 10636 664
rect 10675 631 10709 664
rect 10748 631 10782 664
rect 10821 631 10855 664
rect 10894 631 10928 664
rect 10967 631 11001 664
rect 11040 631 11074 664
rect 11113 631 11147 664
rect 11186 631 11220 664
rect 11259 631 11293 664
rect 11332 631 11366 664
rect 11405 631 11439 664
rect 11478 631 11512 664
rect 11551 631 11585 664
rect 11624 631 11658 664
rect 11697 631 11731 665
rect 15443 671 15477 702
rect 11770 664 11800 665
rect 11800 664 11804 665
rect 11843 664 11869 665
rect 11869 664 11877 665
rect 11915 664 11938 665
rect 11938 664 11949 665
rect 11770 631 11804 664
rect 11843 631 11877 664
rect 11915 631 11949 664
rect 11987 631 12007 665
rect 12007 631 12021 665
rect 12059 631 12093 665
rect 12131 631 12165 665
rect 12203 631 12237 665
rect 12275 631 12309 665
rect 12347 631 12381 665
rect 12419 631 12453 665
rect 12491 631 12525 665
rect 12563 631 12597 665
rect 12635 631 12669 665
rect 12707 631 12741 665
rect 12779 631 12813 665
rect 12851 631 12885 665
rect 12923 631 12957 665
rect 12995 631 13029 665
rect 13067 631 13101 665
rect 13139 631 13173 665
rect 13211 631 13245 665
rect 13283 631 13317 665
rect 13355 631 13389 665
rect 13427 631 13461 665
rect 13499 631 13533 665
rect 13571 631 13605 665
rect 13643 631 13677 665
rect 13715 631 13749 665
rect 13787 631 13821 665
rect 13859 631 13893 665
rect 13931 631 13965 665
rect 14003 631 14037 665
rect 14075 631 14109 665
rect 14147 631 14181 665
rect 14219 631 14253 665
rect 14291 631 15367 665
rect 15371 631 15373 665
rect 15373 631 15405 665
rect 10529 562 10563 593
rect 10602 562 10636 593
rect 10675 562 10709 593
rect 10748 562 10782 593
rect 10821 562 10855 593
rect 10894 562 10928 593
rect 10967 562 11001 593
rect 11040 562 11074 593
rect 11113 562 11147 593
rect 11186 562 11220 593
rect 11259 562 11293 593
rect 11332 562 11366 593
rect 11405 562 11439 593
rect 11478 562 11512 593
rect 11551 562 11585 593
rect 11624 562 11658 593
rect 11697 562 11731 593
rect 11770 562 11804 593
rect 11843 562 11877 593
rect 11916 562 11939 593
rect 11939 562 11950 593
rect 10529 559 10559 562
rect 10559 559 10563 562
rect 10602 559 10628 562
rect 10628 559 10636 562
rect 10675 559 10697 562
rect 10697 559 10709 562
rect 10748 559 10766 562
rect 10766 559 10782 562
rect 10821 559 10835 562
rect 10835 559 10855 562
rect 10894 559 10904 562
rect 10904 559 10928 562
rect 10967 559 10973 562
rect 10973 559 11001 562
rect 11040 559 11042 562
rect 11042 559 11074 562
rect 11113 559 11146 562
rect 11146 559 11147 562
rect 11186 559 11215 562
rect 11215 559 11220 562
rect 11259 559 11284 562
rect 11284 559 11293 562
rect 11332 559 11353 562
rect 11353 559 11366 562
rect 11405 559 11422 562
rect 11422 559 11439 562
rect 11478 559 11491 562
rect 11491 559 11512 562
rect 11551 559 11560 562
rect 11560 559 11585 562
rect 11624 559 11629 562
rect 11629 559 11658 562
rect 11697 559 11698 562
rect 11698 559 11731 562
rect 11770 559 11801 562
rect 11801 559 11804 562
rect 11843 559 11870 562
rect 11870 559 11877 562
rect 11916 559 11950 562
rect 11989 559 12023 593
rect 12062 559 12096 593
rect 12135 559 12169 593
rect 12208 559 12242 593
rect 12281 559 12315 593
rect 12354 559 12388 593
rect 12427 559 12461 593
rect 12500 559 12534 593
rect 12573 559 12607 593
rect 12646 559 12680 593
rect 12719 559 12753 593
rect 12792 559 12826 593
rect 12865 559 12899 593
rect 12938 559 12972 593
rect 13011 559 13045 593
rect 13084 559 13118 593
rect 13157 559 13191 593
rect 13230 559 13264 593
rect 13303 559 13337 593
rect 13376 559 13410 593
rect 13449 559 13483 593
rect 13522 559 13556 593
rect 13595 559 13629 593
rect 13668 559 13702 593
rect 13741 559 13775 593
rect 13814 559 13848 593
rect 13887 559 13921 593
rect 13960 559 13994 593
rect 14033 559 14067 593
rect 14106 559 14140 593
rect 14179 559 14213 593
rect 14252 559 14286 593
rect 14325 559 15367 631
rect 15443 597 15477 631
rect 15693 3383 15727 3406
rect 15765 3402 15797 3420
rect 15797 3402 15799 3420
rect 15693 3372 15695 3383
rect 15695 3372 15727 3383
rect 15765 3352 15799 3363
rect 15693 3314 15727 3334
rect 15765 3329 15797 3352
rect 15797 3329 15799 3352
rect 15693 3300 15695 3314
rect 15695 3300 15727 3314
rect 15765 3284 15799 3290
rect 15693 3245 15727 3262
rect 15765 3256 15797 3284
rect 15797 3256 15799 3284
rect 15693 3228 15695 3245
rect 15695 3228 15727 3245
rect 15765 3216 15799 3217
rect 15693 3176 15727 3190
rect 15765 3183 15797 3216
rect 15797 3183 15799 3216
rect 15693 3156 15695 3176
rect 15695 3156 15727 3176
rect 15693 3107 15727 3118
rect 15765 3114 15797 3144
rect 15797 3114 15799 3144
rect 15765 3110 15799 3114
rect 15693 3084 15695 3107
rect 15695 3084 15727 3107
rect 15765 3046 15797 3071
rect 15797 3046 15799 3071
rect 15693 3038 15727 3046
rect 15693 3012 15695 3038
rect 15695 3012 15727 3038
rect 15765 3037 15799 3046
rect 15765 2978 15797 2998
rect 15797 2978 15799 2998
rect 15693 2969 15727 2974
rect 15693 2940 15695 2969
rect 15695 2940 15727 2969
rect 15765 2964 15799 2978
rect 15765 2910 15797 2925
rect 15797 2910 15799 2925
rect 15693 2900 15727 2902
rect 15693 2868 15695 2900
rect 15695 2868 15727 2900
rect 15765 2891 15799 2910
rect 15765 2842 15797 2852
rect 15797 2842 15799 2852
rect 15693 2797 15695 2830
rect 15695 2797 15727 2830
rect 15693 2796 15727 2797
rect 15765 2818 15799 2842
rect 15765 2774 15797 2779
rect 15797 2774 15799 2779
rect 15693 2728 15695 2758
rect 15695 2728 15727 2758
rect 15693 2724 15727 2728
rect 15765 2745 15799 2774
rect 15693 2659 15695 2686
rect 15695 2659 15727 2686
rect 15693 2652 15727 2659
rect 15765 2672 15799 2706
rect 15693 2590 15695 2614
rect 15695 2590 15727 2614
rect 15693 2580 15727 2590
rect 15765 2604 15799 2633
rect 15765 2599 15797 2604
rect 15797 2599 15799 2604
rect 15693 2521 15695 2542
rect 15695 2521 15727 2542
rect 15693 2508 15727 2521
rect 15765 2536 15799 2560
rect 15765 2526 15797 2536
rect 15797 2526 15799 2536
rect 15693 2452 15695 2469
rect 15695 2452 15727 2469
rect 15693 2435 15727 2452
rect 15765 2468 15799 2487
rect 15765 2453 15797 2468
rect 15797 2453 15799 2468
rect 15693 2383 15695 2396
rect 15695 2383 15727 2396
rect 15693 2362 15727 2383
rect 15765 2400 15799 2414
rect 15765 2380 15797 2400
rect 15797 2380 15799 2400
rect 15693 2314 15695 2323
rect 15695 2314 15727 2323
rect 15693 2289 15727 2314
rect 15765 2331 15799 2341
rect 15765 2307 15797 2331
rect 15797 2307 15799 2331
rect 15693 2245 15695 2250
rect 15695 2245 15727 2250
rect 15693 2216 15727 2245
rect 15765 2262 15799 2268
rect 15765 2234 15797 2262
rect 15797 2234 15799 2262
rect 15693 2176 15695 2177
rect 15695 2176 15727 2177
rect 15693 2143 15727 2176
rect 15765 2193 15799 2195
rect 15765 2161 15797 2193
rect 15797 2161 15799 2193
rect 15693 2072 15727 2104
rect 15765 2090 15797 2122
rect 15797 2090 15799 2122
rect 15765 2088 15799 2090
rect 15693 2070 15695 2072
rect 15695 2070 15727 2072
rect 15693 2003 15727 2031
rect 15765 2021 15797 2049
rect 15797 2021 15799 2049
rect 15765 2015 15799 2021
rect 15693 1997 15695 2003
rect 15695 1997 15727 2003
rect 15693 1934 15727 1958
rect 15765 1952 15797 1976
rect 15797 1952 15799 1976
rect 15765 1942 15799 1952
rect 15693 1924 15695 1934
rect 15695 1924 15727 1934
rect 15693 1865 15727 1885
rect 15765 1883 15797 1903
rect 15797 1883 15799 1903
rect 15765 1869 15799 1883
rect 15693 1851 15695 1865
rect 15695 1851 15727 1865
rect 15765 1814 15797 1830
rect 15797 1814 15799 1830
rect 15693 1796 15727 1812
rect 15765 1796 15799 1814
rect 15693 1778 15695 1796
rect 15695 1778 15727 1796
rect 15765 1745 15797 1757
rect 15797 1745 15799 1757
rect 15693 1727 15727 1739
rect 15693 1705 15695 1727
rect 15695 1705 15727 1727
rect 15765 1723 15799 1745
rect 15765 1676 15797 1684
rect 15797 1676 15799 1684
rect 15693 1658 15727 1666
rect 15693 1632 15695 1658
rect 15695 1632 15727 1658
rect 15765 1650 15799 1676
rect 15765 1607 15797 1610
rect 15797 1607 15799 1610
rect 15693 1589 15727 1593
rect 15693 1559 15695 1589
rect 15695 1559 15727 1589
rect 15765 1576 15799 1607
rect 15693 1486 15695 1520
rect 15695 1486 15727 1520
rect 15765 1503 15799 1536
rect 15765 1502 15797 1503
rect 15797 1502 15799 1503
rect 15693 1416 15695 1447
rect 15695 1416 15727 1447
rect 15765 1434 15799 1462
rect 15765 1428 15797 1434
rect 15797 1428 15799 1434
rect 15693 1413 15727 1416
rect 15693 1346 15695 1374
rect 15695 1346 15727 1374
rect 15765 1365 15799 1388
rect 15765 1354 15797 1365
rect 15797 1354 15799 1365
rect 15693 1340 15727 1346
rect 15693 1276 15695 1301
rect 15695 1276 15727 1301
rect 15765 1296 15799 1314
rect 15765 1280 15797 1296
rect 15797 1280 15799 1296
rect 15693 1267 15727 1276
rect 15693 1206 15695 1228
rect 15695 1206 15727 1228
rect 15765 1227 15799 1240
rect 15765 1206 15797 1227
rect 15797 1206 15799 1227
rect 15693 1194 15727 1206
rect 15693 1136 15695 1155
rect 15695 1136 15727 1155
rect 15765 1158 15799 1166
rect 15693 1121 15727 1136
rect 15765 1132 15797 1158
rect 15797 1132 15799 1158
rect 15693 1066 15695 1082
rect 15695 1066 15727 1082
rect 15765 1089 15799 1092
rect 15693 1048 15727 1066
rect 15765 1058 15797 1089
rect 15797 1058 15799 1089
rect 15693 996 15695 1009
rect 15695 996 15727 1009
rect 15693 975 15727 996
rect 15765 986 15797 1018
rect 15797 986 15799 1018
rect 15765 984 15799 986
rect 15693 926 15695 936
rect 15695 926 15727 936
rect 15693 902 15727 926
rect 15765 917 15797 944
rect 15797 917 15799 944
rect 15765 910 15799 917
rect 15693 856 15695 863
rect 15695 856 15727 863
rect 15693 829 15727 856
rect 15765 848 15797 870
rect 15797 848 15799 870
rect 15765 836 15799 848
rect 15693 786 15695 790
rect 15695 786 15727 790
rect 15693 756 15727 786
rect 15765 779 15797 796
rect 15797 779 15799 796
rect 15765 762 15799 779
rect 15693 716 15695 717
rect 15695 716 15727 717
rect 15693 683 15727 716
rect 15765 710 15797 722
rect 15797 710 15799 722
rect 15765 688 15799 710
rect 15693 610 15727 644
rect 15765 641 15797 648
rect 15797 641 15799 648
rect 15765 614 15799 641
rect 15765 572 15797 574
rect 15797 572 15799 574
rect 15693 540 15727 571
rect 15765 540 15799 572
rect 15693 537 15695 540
rect 15695 537 15727 540
rect 15693 470 15727 498
rect 15693 464 15695 470
rect 15695 464 15727 470
rect 15765 468 15799 500
rect 15765 466 15797 468
rect 15797 466 15799 468
rect 10809 365 10811 399
rect 10811 365 10843 399
rect 10881 365 10915 399
rect 12951 365 12985 399
rect 13023 365 13055 399
rect 13055 365 13057 399
rect 15693 400 15727 425
rect 15693 391 15695 400
rect 15695 391 15727 400
rect 15765 399 15799 426
rect 15765 392 15797 399
rect 15797 392 15799 399
rect 15693 330 15727 352
rect 15765 330 15799 352
rect 15693 318 15695 330
rect 15695 318 15727 330
rect 15765 318 15797 330
rect 15797 318 15799 330
<< metal1 >>
rect 349 17425 16555 17431
rect 349 17391 393 17425
rect 427 17391 466 17425
rect 500 17391 539 17425
rect 573 17391 612 17425
rect 646 17391 685 17425
rect 719 17391 758 17425
rect 792 17391 831 17425
rect 865 17391 904 17425
rect 938 17391 977 17425
rect 1011 17391 1050 17425
rect 1084 17391 1123 17425
rect 1157 17391 1196 17425
rect 1230 17391 1269 17425
rect 1303 17391 1342 17425
rect 1376 17391 1415 17425
rect 1449 17391 1488 17425
rect 1522 17391 1561 17425
rect 1595 17391 1634 17425
rect 1668 17391 1707 17425
rect 1741 17391 1780 17425
rect 1814 17391 1853 17425
rect 1887 17391 1926 17425
rect 1960 17391 1999 17425
rect 2033 17391 2072 17425
rect 2106 17391 2145 17425
rect 2179 17391 2218 17425
rect 2252 17391 2291 17425
rect 2325 17391 2364 17425
rect 2398 17391 2437 17425
rect 2471 17391 2510 17425
rect 2544 17391 2583 17425
rect 2617 17391 2656 17425
rect 2690 17391 2729 17425
rect 2763 17391 2802 17425
rect 2836 17391 2875 17425
rect 2909 17391 2948 17425
rect 2982 17391 3021 17425
rect 3055 17391 3094 17425
rect 3128 17391 3167 17425
rect 3201 17391 3240 17425
rect 3274 17391 3313 17425
rect 3347 17391 3386 17425
rect 3420 17391 3459 17425
rect 3493 17391 3532 17425
rect 3566 17391 3605 17425
rect 3639 17391 3678 17425
rect 3712 17391 3751 17425
rect 3785 17391 3824 17425
rect 3858 17391 3897 17425
rect 3931 17391 3970 17425
rect 4004 17391 4043 17425
rect 4077 17391 4116 17425
rect 4150 17391 4189 17425
rect 4223 17391 4262 17425
rect 4296 17391 4335 17425
rect 4369 17391 4408 17425
rect 4442 17391 4481 17425
rect 4515 17391 4554 17425
rect 4588 17391 4627 17425
rect 4661 17391 4700 17425
rect 4734 17391 4773 17425
rect 349 17353 4773 17391
rect 349 17319 427 17353
rect 461 17319 500 17353
rect 534 17319 573 17353
rect 607 17319 646 17353
rect 680 17319 719 17353
rect 753 17319 792 17353
rect 826 17319 865 17353
rect 899 17319 938 17353
rect 972 17319 1011 17353
rect 1045 17319 1084 17353
rect 1118 17319 1157 17353
rect 1191 17319 1230 17353
rect 1264 17319 1303 17353
rect 1337 17319 1376 17353
rect 1410 17319 1449 17353
rect 1483 17319 1522 17353
rect 1556 17319 1595 17353
rect 1629 17319 1668 17353
rect 1702 17319 1741 17353
rect 1775 17319 1814 17353
rect 1848 17319 1887 17353
rect 1921 17319 1960 17353
rect 1994 17319 2033 17353
rect 2067 17319 2106 17353
rect 2140 17319 2179 17353
rect 2213 17319 2252 17353
rect 2286 17319 2325 17353
rect 2359 17319 2397 17353
rect 2431 17319 2469 17353
rect 2503 17319 2541 17353
rect 2575 17319 2613 17353
rect 2647 17319 2685 17353
rect 2719 17319 2757 17353
rect 2791 17319 2829 17353
rect 2863 17319 2901 17353
rect 2935 17319 2973 17353
rect 3007 17319 3045 17353
rect 3079 17319 3117 17353
rect 3151 17319 3189 17353
rect 3223 17319 3261 17353
rect 3295 17319 3333 17353
rect 3367 17319 3405 17353
rect 3439 17319 3477 17353
rect 3511 17319 3549 17353
rect 3583 17319 3621 17353
rect 3655 17319 3693 17353
rect 3727 17319 3765 17353
rect 3799 17319 3837 17353
rect 3871 17319 3909 17353
rect 3943 17319 3981 17353
rect 4015 17319 4053 17353
rect 4087 17319 4125 17353
rect 4159 17319 4197 17353
rect 4231 17319 4269 17353
rect 4303 17319 4341 17353
rect 4375 17319 4413 17353
rect 4447 17319 4485 17353
rect 4519 17319 4557 17353
rect 4591 17319 4629 17353
rect 4663 17319 4701 17353
rect 4735 17319 4773 17353
rect 16543 17319 16555 17425
rect 349 17313 16555 17319
rect 16951 17425 18383 17431
rect 16951 17391 16963 17425
rect 16997 17391 17037 17425
rect 17071 17391 17111 17425
rect 17145 17391 17185 17425
rect 17219 17391 17259 17425
rect 17293 17391 17333 17425
rect 17367 17391 17407 17425
rect 17441 17391 17481 17425
rect 17515 17391 17555 17425
rect 17589 17391 17630 17425
rect 17664 17391 17705 17425
rect 17739 17391 17780 17425
rect 17814 17391 17855 17425
rect 17889 17391 17930 17425
rect 17964 17391 18005 17425
rect 18039 17391 18080 17425
rect 18114 17391 18155 17425
rect 18189 17391 18230 17425
rect 18264 17391 18305 17425
rect 18339 17391 18383 17425
rect 16951 17353 18383 17391
rect 16951 17319 16963 17353
rect 16997 17319 17035 17353
rect 17069 17319 17107 17353
rect 17141 17319 17179 17353
rect 17213 17319 17251 17353
rect 17285 17319 17323 17353
rect 17357 17319 17395 17353
rect 17429 17319 17468 17353
rect 17502 17319 17541 17353
rect 17575 17319 17614 17353
rect 17648 17319 17687 17353
rect 17721 17319 17760 17353
rect 17794 17319 17833 17353
rect 17867 17319 17906 17353
rect 17940 17319 17979 17353
rect 18013 17319 18052 17353
rect 18086 17319 18125 17353
rect 18159 17319 18198 17353
rect 18232 17319 18271 17353
rect 18305 17319 18383 17353
rect 16951 17315 18383 17319
rect 16951 17313 18271 17315
rect 349 17309 467 17313
rect 349 17275 355 17309
rect 389 17280 467 17309
tri 18240 17288 18265 17313 ne
rect 389 17275 427 17280
rect 349 17246 427 17275
rect 461 17246 467 17280
rect 349 17234 467 17246
rect 349 17200 355 17234
rect 389 17207 467 17234
rect 389 17200 427 17207
rect 349 17173 427 17200
rect 461 17173 467 17207
rect 349 17158 467 17173
rect 349 17124 355 17158
rect 389 17134 467 17158
rect 389 17124 427 17134
rect 349 17100 427 17124
rect 461 17100 467 17134
rect 349 17082 467 17100
rect 349 17048 355 17082
rect 389 17061 467 17082
rect 389 17048 427 17061
rect 349 17027 427 17048
rect 461 17027 467 17061
rect 349 17006 467 17027
rect 349 16972 355 17006
rect 389 16988 467 17006
rect 389 16972 427 16988
rect 349 16954 427 16972
rect 461 16954 467 16988
rect 349 16930 467 16954
rect -184 16434 -60 16907
rect 349 16896 355 16930
rect 389 16915 467 16930
rect 389 16896 427 16915
rect 349 16881 427 16896
rect 461 16881 467 16915
rect 349 16854 467 16881
rect 349 16820 355 16854
rect 389 16842 467 16854
rect 389 16820 427 16842
rect 349 16808 427 16820
rect 461 16808 467 16842
rect 349 16778 467 16808
rect 349 16744 355 16778
rect 389 16769 467 16778
rect 389 16744 427 16769
rect 349 16735 427 16744
rect 461 16735 467 16769
rect 349 16702 467 16735
rect 349 16668 355 16702
rect 389 16696 467 16702
rect 389 16668 427 16696
rect 349 16662 427 16668
rect 461 16662 467 16696
rect 349 16626 467 16662
rect 349 16592 355 16626
rect 389 16622 467 16626
rect 389 16592 427 16622
rect 349 16588 427 16592
rect 461 16588 467 16622
rect 349 16550 467 16588
rect 349 16516 355 16550
rect 389 16548 467 16550
rect 389 16516 427 16548
rect 349 16514 427 16516
rect 461 16514 467 16548
rect 672 17140 16419 17146
rect 672 17106 716 17140
rect 750 17106 789 17140
rect 823 17106 862 17140
rect 896 17106 935 17140
rect 969 17106 1008 17140
rect 1042 17106 1081 17140
rect 1115 17106 1154 17140
rect 1188 17106 1227 17140
rect 1261 17106 1300 17140
rect 1334 17106 1373 17140
rect 1407 17106 1446 17140
rect 1480 17106 1519 17140
rect 1553 17106 1592 17140
rect 1626 17106 1665 17140
rect 1699 17106 1738 17140
rect 1772 17106 1811 17140
rect 1845 17106 1884 17140
rect 1918 17106 1957 17140
rect 1991 17106 2030 17140
rect 2064 17106 2103 17140
rect 2137 17106 2176 17140
rect 2210 17106 2249 17140
rect 2283 17106 2322 17140
rect 2356 17106 2395 17140
rect 2429 17106 2468 17140
rect 2502 17106 2541 17140
rect 2575 17106 2614 17140
rect 2648 17106 2687 17140
rect 2721 17106 2760 17140
rect 2794 17106 2833 17140
rect 2867 17106 2906 17140
rect 2940 17106 2979 17140
rect 3013 17106 3052 17140
rect 3086 17106 3125 17140
rect 3159 17106 3197 17140
rect 3231 17106 3269 17140
rect 3303 17106 3341 17140
rect 3375 17106 3413 17140
rect 3447 17106 3485 17140
rect 3519 17106 3557 17140
rect 3591 17106 3629 17140
rect 3663 17106 3701 17140
rect 3735 17106 3773 17140
rect 3807 17106 3845 17140
rect 3879 17106 3917 17140
rect 3951 17106 3989 17140
rect 4023 17106 4061 17140
rect 4095 17106 4133 17140
rect 4167 17106 4205 17140
rect 4239 17106 4277 17140
rect 4311 17106 4349 17140
rect 4383 17106 4421 17140
rect 4455 17106 4493 17140
rect 4527 17106 4565 17140
rect 4599 17106 4637 17140
rect 4671 17106 4709 17140
rect 4743 17106 4781 17140
rect 4815 17106 4853 17140
rect 4887 17106 4925 17140
rect 4959 17106 4997 17140
rect 5031 17106 5069 17140
rect 5103 17106 5141 17140
rect 5175 17106 5213 17140
rect 5247 17106 5285 17140
rect 5319 17106 5357 17140
rect 5391 17106 5429 17140
rect 5463 17106 5501 17140
rect 5535 17106 5573 17140
rect 5607 17106 5645 17140
rect 5679 17106 5717 17140
rect 5751 17106 5789 17140
rect 5823 17106 5861 17140
rect 5895 17106 5933 17140
rect 672 17068 5933 17106
rect 672 17034 750 17068
rect 784 17034 823 17068
rect 857 17034 896 17068
rect 930 17034 969 17068
rect 1003 17034 1042 17068
rect 1076 17034 1115 17068
rect 1149 17034 1188 17068
rect 1222 17034 1261 17068
rect 1295 17034 1334 17068
rect 1368 17034 1407 17068
rect 1441 17034 1480 17068
rect 1514 17034 1553 17068
rect 1587 17034 1626 17068
rect 1660 17034 1699 17068
rect 1733 17034 1772 17068
rect 1806 17034 1845 17068
rect 1879 17034 1918 17068
rect 1952 17034 1991 17068
rect 2025 17034 2064 17068
rect 2098 17034 2137 17068
rect 2171 17034 2210 17068
rect 2244 17034 2283 17068
rect 2317 17034 2356 17068
rect 2390 17034 2429 17068
rect 2463 17034 2502 17068
rect 2536 17034 2575 17068
rect 2609 17034 2648 17068
rect 2682 17034 2721 17068
rect 2755 17034 2794 17068
rect 2828 17034 2867 17068
rect 2901 17034 2940 17068
rect 2974 17034 3013 17068
rect 3047 17034 3086 17068
rect 3120 17034 3159 17068
rect 3193 17034 3232 17068
rect 3266 17034 3305 17068
rect 3339 17034 3378 17068
rect 3412 17034 3451 17068
rect 3485 17034 3524 17068
rect 3558 17034 3597 17068
rect 3631 17034 3670 17068
rect 3704 17034 3743 17068
rect 3777 17034 3816 17068
rect 3850 17034 3889 17068
rect 3923 17034 3962 17068
rect 3996 17034 4035 17068
rect 4069 17034 4108 17068
rect 4142 17034 4181 17068
rect 4215 17034 4254 17068
rect 4288 17034 4327 17068
rect 4361 17034 4400 17068
rect 4434 17034 4473 17068
rect 4507 17034 4546 17068
rect 4580 17034 4619 17068
rect 4653 17034 4692 17068
rect 4726 17034 4765 17068
rect 4799 17034 4838 17068
rect 4872 17034 4911 17068
rect 4945 17034 4984 17068
rect 5018 17034 5057 17068
rect 5091 17034 5130 17068
rect 5164 17034 5203 17068
rect 5237 17034 5276 17068
rect 5310 17034 5349 17068
rect 5383 17034 5422 17068
rect 5456 17034 5495 17068
rect 5529 17034 5568 17068
rect 5602 17034 5641 17068
rect 5675 17034 5714 17068
rect 5748 17034 5787 17068
rect 5821 17034 5860 17068
rect 5894 17034 5933 17068
rect 16407 17034 16419 17140
rect 672 17028 7951 17034
rect 672 16994 678 17028
rect 712 16994 790 17028
tri 3188 16996 3220 17028 ne
rect 3220 16996 3420 17028
tri 3420 16996 3452 17028 nw
tri 5530 16996 5562 17028 ne
rect 5562 16996 5728 17028
rect 672 16988 790 16994
rect 672 16955 750 16988
rect 672 16921 678 16955
rect 712 16954 750 16955
rect 784 16954 790 16988
tri 3220 16962 3254 16996 ne
rect 3254 16962 3267 16996
rect 3301 16962 3339 16996
rect 3373 16962 3386 16996
tri 3386 16962 3420 16996 nw
tri 5562 16962 5596 16996 ne
rect 5596 16962 5609 16996
rect 5643 16962 5681 16996
rect 5715 16962 5728 16996
tri 5728 16962 5794 17028 nw
tri 7872 16962 7938 17028 ne
rect 7938 16962 7951 17028
rect 8057 17028 10293 17034
rect 8057 16962 8070 17028
tri 8070 16962 8136 17028 nw
tri 10214 16962 10280 17028 ne
rect 10280 16962 10293 17028
rect 10399 17028 16419 17034
rect 17134 17102 18060 17108
rect 17134 17068 17146 17102
rect 17180 17068 17222 17102
rect 17256 17068 17298 17102
rect 17332 17068 17374 17102
rect 17408 17068 17450 17102
rect 17484 17068 17526 17102
rect 17560 17068 17602 17102
rect 17636 17068 17678 17102
rect 17712 17068 17754 17102
rect 17788 17068 17830 17102
rect 17864 17068 17906 17102
rect 17940 17068 17982 17102
rect 18016 17068 18060 17102
rect 17134 17030 18060 17068
rect 10399 16996 15749 17028
tri 15749 16996 15781 17028 nw
rect 17134 16996 17146 17030
rect 17180 16996 17218 17030
rect 17252 16996 17291 17030
rect 17325 16996 17364 17030
rect 17398 16996 17437 17030
rect 17471 16996 17510 17030
rect 17544 16996 17583 17030
rect 17617 16996 17656 17030
rect 17690 16996 17729 17030
rect 17763 16996 17802 17030
rect 17836 16996 17875 17030
rect 17909 16996 17948 17030
rect 17982 16996 18060 17030
rect 10399 16992 15745 16996
tri 15745 16992 15749 16996 nw
rect 17134 16992 18060 16996
rect 10399 16973 15677 16992
rect 10399 16962 10476 16973
tri 3254 16955 3261 16962 ne
rect 712 16921 790 16954
rect 672 16908 790 16921
rect 672 16882 750 16908
rect 672 16848 678 16882
rect 712 16874 750 16882
rect 784 16874 790 16908
rect 712 16848 790 16874
rect 672 16828 790 16848
rect 672 16808 750 16828
rect 672 16774 678 16808
rect 712 16794 750 16808
rect 784 16794 790 16828
rect 712 16774 790 16794
rect 672 16748 790 16774
rect 672 16734 750 16748
rect 672 16700 678 16734
rect 712 16714 750 16734
rect 784 16714 790 16748
rect 712 16700 790 16714
rect 672 16667 790 16700
rect 672 16660 750 16667
rect 672 16626 678 16660
rect 712 16633 750 16660
rect 784 16633 790 16667
rect 712 16626 790 16633
rect 672 16586 790 16626
rect 672 16552 678 16586
rect 712 16552 750 16586
rect 784 16552 790 16586
rect 672 16540 790 16552
rect 3261 16916 3379 16962
tri 3379 16955 3386 16962 nw
tri 5596 16955 5603 16962 ne
rect 3261 16882 3267 16916
rect 3301 16882 3339 16916
rect 3373 16882 3379 16916
rect 3261 16836 3379 16882
rect 3261 16802 3267 16836
rect 3301 16802 3339 16836
rect 3373 16802 3379 16836
rect 3261 16756 3379 16802
rect 3261 16722 3267 16756
rect 3301 16722 3339 16756
rect 3373 16722 3379 16756
rect 3261 16676 3379 16722
rect 3261 16642 3267 16676
rect 3301 16642 3339 16676
rect 3373 16642 3379 16676
rect 3261 16596 3379 16642
rect 3261 16562 3267 16596
rect 3301 16562 3339 16596
rect 3373 16562 3379 16596
rect 349 16474 467 16514
rect 349 16440 355 16474
rect 389 16440 427 16474
rect 461 16440 467 16474
rect 3261 16515 3379 16562
rect 3261 16481 3267 16515
rect 3301 16481 3339 16515
rect 3373 16481 3379 16515
tri -60 16434 -58 16436 sw
rect -184 16400 -58 16434
tri -58 16400 -24 16434 sw
rect 349 16428 467 16440
tri 1213 16434 1220 16441 se
rect 1220 16434 3078 16441
tri 3078 16434 3085 16441 sw
rect 3261 16434 3379 16481
rect 5603 16916 5721 16962
tri 5721 16955 5728 16962 nw
tri 7938 16955 7945 16962 ne
rect 5603 16882 5609 16916
rect 5643 16882 5681 16916
rect 5715 16882 5721 16916
rect 5603 16836 5721 16882
rect 5603 16802 5609 16836
rect 5643 16802 5681 16836
rect 5715 16802 5721 16836
rect 5603 16756 5721 16802
rect 5603 16722 5609 16756
rect 5643 16722 5681 16756
rect 5715 16722 5721 16756
rect 5603 16676 5721 16722
rect 5603 16642 5609 16676
rect 5643 16642 5681 16676
rect 5715 16642 5721 16676
rect 5603 16596 5721 16642
rect 5603 16562 5609 16596
rect 5643 16562 5681 16596
rect 5715 16562 5721 16596
rect 5603 16515 5721 16562
rect 5603 16481 5609 16515
rect 5643 16481 5681 16515
rect 5715 16481 5721 16515
tri 3555 16434 3562 16441 se
rect 3562 16434 5420 16441
tri 5420 16434 5427 16441 sw
rect 5603 16434 5721 16481
rect 7945 16916 8063 16962
tri 8063 16955 8070 16962 nw
tri 10280 16955 10287 16962 ne
rect 7945 16882 7951 16916
rect 7985 16882 8023 16916
rect 8057 16882 8063 16916
rect 7945 16836 8063 16882
rect 7945 16802 7951 16836
rect 7985 16802 8023 16836
rect 8057 16802 8063 16836
rect 7945 16756 8063 16802
rect 7945 16722 7951 16756
rect 7985 16722 8023 16756
rect 8057 16722 8063 16756
rect 7945 16676 8063 16722
rect 7945 16642 7951 16676
rect 7985 16642 8023 16676
rect 8057 16642 8063 16676
rect 7945 16596 8063 16642
rect 7945 16562 7951 16596
rect 7985 16562 8023 16596
rect 8057 16562 8063 16596
rect 7945 16515 8063 16562
rect 7945 16481 7951 16515
rect 7985 16481 8023 16515
rect 8057 16481 8063 16515
tri 5897 16434 5904 16441 se
rect 5904 16434 7762 16441
tri 7762 16434 7769 16441 sw
rect 7945 16434 8063 16481
rect 10287 16939 10476 16962
rect 10510 16939 10549 16973
rect 10583 16939 10622 16973
rect 10656 16939 10695 16973
rect 10729 16939 10768 16973
rect 10802 16939 10841 16973
rect 10875 16939 10914 16973
rect 10948 16939 10987 16973
rect 11021 16939 11060 16973
rect 11094 16939 11133 16973
rect 10287 16916 11133 16939
rect 10287 16882 10293 16916
rect 10327 16882 10365 16916
rect 10399 16901 11133 16916
rect 10399 16882 10476 16901
rect 10287 16867 10476 16882
rect 10510 16867 10549 16901
rect 10583 16867 10622 16901
rect 10656 16867 10695 16901
rect 10729 16867 10768 16901
rect 10802 16867 10841 16901
rect 10875 16867 10914 16901
rect 10948 16867 10987 16901
rect 11021 16867 11060 16901
rect 11094 16867 11133 16901
rect 15199 16924 15677 16973
tri 15677 16924 15745 16992 nw
rect 17134 16990 17948 16992
rect 17942 16924 17948 16990
rect 18054 16924 18060 16992
rect 15199 16922 15673 16924
rect 15199 16888 15396 16922
rect 15430 16920 15673 16922
tri 15673 16920 15677 16924 nw
rect 17942 16920 18060 16924
rect 15430 16888 15639 16920
rect 15199 16886 15639 16888
tri 15639 16886 15673 16920 nw
rect 17942 16886 18020 16920
rect 18054 16886 18060 16920
rect 15199 16885 15638 16886
tri 15638 16885 15639 16886 nw
rect 17942 16885 18060 16886
rect 15199 16867 15628 16885
tri 15628 16875 15638 16885 nw
rect 10287 16849 15628 16867
rect 10287 16836 15396 16849
rect 10287 16802 10293 16836
rect 10327 16802 10365 16836
rect 10399 16815 15396 16836
rect 15430 16815 15628 16849
rect 10399 16812 15628 16815
rect 10399 16802 10419 16812
rect 10287 16778 10419 16802
tri 10419 16778 10453 16812 nw
tri 15055 16778 15089 16812 ne
rect 15089 16778 15628 16812
rect 10287 16776 10417 16778
tri 10417 16776 10419 16778 nw
tri 15089 16776 15091 16778 ne
rect 15091 16776 15628 16778
rect 10287 16756 10405 16776
tri 10405 16764 10417 16776 nw
tri 15091 16764 15103 16776 ne
rect 15103 16764 15396 16776
rect 10287 16722 10293 16756
rect 10327 16722 10365 16756
rect 10399 16722 10405 16756
tri 15103 16743 15124 16764 ne
rect 15124 16743 15396 16764
rect 10287 16676 10405 16722
rect 10287 16642 10293 16676
rect 10327 16642 10365 16676
rect 10399 16642 10405 16676
rect 10287 16596 10405 16642
rect 10287 16562 10293 16596
rect 10327 16562 10365 16596
rect 10399 16562 10405 16596
rect 10287 16515 10405 16562
rect 10287 16481 10293 16515
rect 10327 16481 10365 16515
rect 10399 16481 10405 16515
tri 8239 16434 8246 16441 se
rect 8246 16434 10104 16441
tri 10104 16434 10111 16441 sw
rect 10287 16434 10405 16481
tri 1207 16428 1213 16434 se
rect 1213 16428 3085 16434
tri 1179 16400 1207 16428 se
rect 1207 16400 3085 16428
tri 3085 16400 3119 16434 sw
rect 3261 16400 3267 16434
rect 3301 16400 3339 16434
rect 3373 16400 3379 16434
tri 3521 16400 3555 16434 se
rect 3555 16400 5427 16434
tri 5427 16400 5461 16434 sw
rect 5603 16400 5609 16434
rect 5643 16400 5681 16434
rect 5715 16400 5721 16434
tri 5863 16400 5897 16434 se
rect 5897 16400 7769 16434
tri 7769 16400 7803 16434 sw
rect 7945 16400 7951 16434
rect 7985 16400 8023 16434
rect 8057 16400 8063 16434
tri 8205 16400 8239 16434 se
rect 8239 16400 10111 16434
tri 10111 16400 10145 16434 sw
rect 10287 16400 10293 16434
rect 10327 16400 10365 16434
rect 10399 16400 10405 16434
rect -184 16381 -24 16400
tri -24 16381 -5 16400 sw
tri 1160 16381 1179 16400 se
rect 1179 16381 3119 16400
tri 3119 16381 3138 16400 sw
rect 3261 16388 3379 16400
tri 3509 16388 3521 16400 se
rect 3521 16388 5461 16400
tri 3502 16381 3509 16388 se
rect 3509 16381 5461 16388
tri 5461 16381 5480 16400 sw
rect 5603 16388 5721 16400
tri 5851 16388 5863 16400 se
rect 5863 16388 7803 16400
tri 5844 16381 5851 16388 se
rect 5851 16381 7803 16388
tri 7803 16381 7822 16400 sw
rect 7945 16388 8063 16400
tri 8193 16388 8205 16400 se
rect 8205 16388 10145 16400
tri 8186 16381 8193 16388 se
rect 8193 16381 10145 16388
tri 10145 16381 10164 16400 sw
rect 10287 16388 10405 16400
rect -184 16351 -5 16381
tri -5 16351 25 16381 sw
tri 1130 16351 1160 16381 se
rect 1160 16351 3138 16381
rect -184 16347 969 16351
tri 969 16347 973 16351 sw
tri 1126 16347 1130 16351 se
rect 1130 16347 3138 16351
tri 3138 16347 3172 16381 sw
tri 3468 16347 3502 16381 se
rect 3502 16347 5480 16381
tri 5480 16347 5514 16381 sw
tri 5810 16347 5844 16381 se
rect 5844 16347 7822 16381
tri 7822 16347 7856 16381 sw
tri 8152 16347 8186 16381 se
rect 8186 16347 10164 16381
tri 10164 16347 10198 16381 sw
rect -184 16340 973 16347
tri 973 16340 980 16347 sw
tri 1119 16340 1126 16347 se
rect 1126 16340 3172 16347
tri 3172 16340 3179 16347 sw
tri 3461 16340 3468 16347 se
rect 3468 16340 5514 16347
tri 5514 16340 5521 16347 sw
tri 5803 16340 5810 16347 se
rect 5810 16340 7856 16347
tri 7856 16340 7863 16347 sw
tri 8145 16340 8152 16347 se
rect 8152 16340 10198 16347
tri 10198 16340 10205 16347 sw
rect -184 16338 980 16340
tri 980 16338 982 16340 sw
tri 1117 16338 1119 16340 se
rect 1119 16338 3179 16340
tri 3179 16338 3181 16340 sw
tri 3459 16338 3461 16340 se
rect 3461 16338 5521 16340
tri 5521 16338 5523 16340 sw
tri 5801 16338 5803 16340 se
rect 5803 16338 7863 16340
tri 7863 16338 7865 16340 sw
tri 8143 16338 8145 16340 se
rect 8145 16338 10205 16340
tri 10205 16338 10207 16340 sw
rect -184 16315 982 16338
tri 982 16315 1005 16338 sw
tri 1094 16315 1117 16338 se
rect 1117 16315 3181 16338
tri 3181 16315 3204 16338 sw
tri 3436 16315 3459 16338 se
rect 3459 16315 5523 16338
tri 5523 16315 5546 16338 sw
tri 5778 16315 5801 16338 se
rect 5801 16315 7865 16338
tri 7865 16315 7888 16338 sw
tri 8120 16315 8143 16338 se
rect 8143 16315 10207 16338
tri 10207 16315 10230 16338 sw
rect -184 16302 1005 16315
tri 1005 16302 1018 16315 sw
tri 1081 16302 1094 16315 se
rect 1094 16302 3204 16315
rect -184 16299 3204 16302
tri 3204 16299 3220 16315 sw
tri 3420 16299 3436 16315 se
rect 3436 16299 5546 16315
tri 5546 16299 5562 16315 sw
tri 5762 16299 5778 16315 se
rect 5778 16299 7888 16315
tri 7888 16299 7904 16315 sw
tri 8104 16299 8120 16315 se
rect 8120 16299 10230 16315
rect -184 16281 10230 16299
tri 10230 16281 10264 16315 sw
rect -184 16275 10264 16281
tri 10264 16275 10270 16281 sw
rect -184 16269 10270 16275
tri 10270 16269 10276 16275 sw
rect -184 16267 10276 16269
tri 10276 16267 10278 16269 sw
rect -184 16265 10278 16267
tri 10278 16265 10280 16267 sw
rect -184 16235 10280 16265
tri 10280 16235 10310 16265 sw
rect -184 16229 10310 16235
tri 10310 16229 10316 16235 sw
rect -184 16195 10316 16229
tri 10316 16195 10350 16229 sw
rect -184 16194 10350 16195
tri 10350 16194 10351 16195 sw
rect -184 16192 10351 16194
tri 10351 16192 10353 16194 sw
rect 10651 16193 14861 16743
tri 15124 16742 15125 16743 ne
rect 15125 16742 15396 16743
rect 15430 16742 15628 16776
tri 15125 16739 15128 16742 ne
rect 15128 16739 15628 16742
tri 15128 16705 15162 16739 ne
rect 15162 16705 15628 16739
tri 15162 16704 15163 16705 ne
rect 15163 16704 15628 16705
tri 15163 16703 15164 16704 ne
rect 15164 16703 15628 16704
tri 15164 16669 15198 16703 ne
rect 15198 16669 15396 16703
rect 15430 16669 15628 16703
tri 15198 16666 15201 16669 ne
rect 15201 16666 15628 16669
tri 15201 16632 15235 16666 ne
rect 15235 16632 15628 16666
tri 15235 16630 15237 16632 ne
rect 15237 16630 15628 16632
tri 15237 16596 15271 16630 ne
rect 15271 16596 15396 16630
rect 15430 16596 15628 16630
tri 15271 16593 15274 16596 ne
rect 15274 16593 15628 16596
tri 15274 16559 15308 16593 ne
rect 15308 16559 15628 16593
tri 15308 16557 15310 16559 ne
rect 15310 16557 15628 16559
tri 15310 16523 15344 16557 ne
rect 15344 16523 15396 16557
rect 15430 16523 15628 16557
tri 15344 16520 15347 16523 ne
rect 15347 16520 15628 16523
tri 15347 16486 15381 16520 ne
rect 15381 16486 15628 16520
tri 15381 16484 15383 16486 ne
rect 15383 16484 15628 16486
tri 15383 16477 15390 16484 ne
tri 15004 16450 15027 16473 se
rect 15027 16450 15079 16473
tri 15001 16447 15004 16450 se
rect 15004 16447 15079 16450
tri 14967 16413 15001 16447 se
rect 15001 16415 15079 16447
rect 15080 16416 15081 16472
rect 15117 16416 15118 16472
rect 15119 16415 15354 16473
rect 15001 16413 15077 16415
tri 15077 16413 15079 16415 nw
tri 15223 16413 15225 16415 ne
rect 15225 16413 15354 16415
tri 14965 16411 14967 16413 se
rect 14967 16411 15075 16413
tri 15075 16411 15077 16413 nw
tri 15225 16411 15227 16413 ne
rect 15227 16411 15354 16413
tri 14963 16409 14965 16411 se
rect 14965 16409 15054 16411
rect 14963 16347 15054 16409
tri 15054 16390 15075 16411 nw
tri 15227 16390 15248 16411 ne
rect 15248 16390 15354 16411
tri 15248 16387 15251 16390 ne
rect 15251 16387 15354 16390
rect 15150 16381 15208 16387
tri 15144 16352 15150 16358 se
rect 15150 16352 15162 16381
tri 15054 16347 15059 16352 sw
tri 15139 16347 15144 16352 se
rect 15144 16347 15162 16352
rect 15196 16347 15208 16381
tri 15251 16377 15261 16387 ne
rect 15261 16377 15354 16387
tri 15261 16375 15263 16377 ne
rect 14963 16340 15059 16347
tri 15059 16340 15066 16347 sw
tri 15132 16340 15139 16347 se
rect 15139 16340 15208 16347
rect 14963 16338 15066 16340
tri 15066 16338 15068 16340 sw
tri 15130 16338 15132 16340 se
rect 15132 16338 15208 16340
rect 14963 16327 15068 16338
tri 15068 16327 15079 16338 sw
tri 15119 16327 15130 16338 se
rect 15130 16327 15208 16338
rect 14963 16315 15079 16327
rect 15081 16326 15117 16327
rect 14963 16281 14969 16315
rect 15003 16281 15041 16315
rect 15075 16281 15079 16315
rect 14963 16269 15079 16281
rect 15080 16270 15118 16326
rect 15119 16309 15208 16327
rect 15119 16275 15162 16309
rect 15196 16275 15208 16309
rect 15081 16269 15117 16270
rect 15119 16269 15208 16275
rect -184 16163 10353 16192
tri 10353 16163 10382 16192 sw
rect 10652 16191 14860 16192
rect 14963 16229 15079 16241
rect 15081 16240 15117 16241
rect 14963 16195 14969 16229
rect 15003 16195 15041 16229
rect 15075 16195 15079 16229
rect 14963 16183 15079 16195
rect 15080 16184 15118 16240
rect 15119 16235 15208 16241
rect 15119 16201 15162 16235
rect 15196 16201 15208 16235
rect 15081 16183 15117 16184
rect 15119 16183 15208 16201
rect 14963 16163 15059 16183
tri 15059 16163 15079 16183 nw
tri 15119 16163 15139 16183 ne
rect 15139 16163 15208 16183
rect -184 16138 10382 16163
tri -184 16129 -175 16138 ne
rect -175 16129 10382 16138
tri 10382 16129 10416 16163 sw
rect 10652 16134 14860 16135
tri 10647 16129 10651 16133 se
rect 10651 16129 14861 16133
tri 14861 16129 14865 16133 sw
tri -175 16121 -167 16129 ne
rect -167 16121 10416 16129
tri 10416 16121 10424 16129 sw
tri 10639 16121 10647 16129 se
rect 10647 16121 14865 16129
tri 14865 16121 14873 16129 sw
tri -167 16119 -165 16121 ne
rect -165 16119 10424 16121
tri 10424 16119 10426 16121 sw
tri 10637 16119 10639 16121 se
rect 10639 16119 14873 16121
tri 14873 16119 14875 16121 sw
rect 14963 16119 15054 16163
tri 15054 16158 15059 16163 nw
tri 15139 16158 15144 16163 ne
rect 15144 16158 15162 16163
tri 15144 16152 15150 16158 ne
rect 15150 16129 15162 16158
rect 15196 16129 15208 16163
rect 15150 16123 15208 16129
tri 15251 16123 15263 16135 se
rect 15263 16123 15354 16377
tri 15249 16121 15251 16123 se
rect 15251 16121 15354 16123
tri 15248 16120 15249 16121 se
rect 15249 16120 15354 16121
tri 15054 16119 15055 16120 sw
tri 15247 16119 15248 16120 se
rect 15248 16119 15354 16120
tri -165 16085 -131 16119 ne
rect -131 16085 10426 16119
tri 10426 16085 10460 16119 sw
tri 10603 16085 10637 16119 se
rect 10637 16101 14875 16119
tri 14875 16101 14893 16119 sw
rect 14963 16101 15055 16119
rect 10637 16085 14893 16101
tri 14893 16085 14909 16101 sw
tri 14963 16085 14979 16101 ne
rect 14979 16095 15055 16101
tri 15055 16095 15079 16119 sw
tri 15223 16095 15247 16119 se
rect 15247 16095 15354 16119
rect 14979 16085 15079 16095
tri -131 16082 -128 16085 ne
rect -128 16082 10460 16085
tri 10460 16082 10463 16085 sw
tri 10600 16082 10603 16085 se
rect 10603 16082 14909 16085
tri 14909 16082 14912 16085 sw
tri 14979 16082 14982 16085 ne
rect 14982 16082 15079 16085
tri -128 16048 -94 16082 ne
rect -94 16048 14912 16082
tri 14912 16048 14946 16082 sw
tri 14982 16048 15016 16082 ne
rect 15016 16048 15079 16082
tri -94 16046 -92 16048 ne
rect -92 16046 14946 16048
tri 14946 16046 14948 16048 sw
tri 15016 16046 15018 16048 ne
rect 15018 16046 15079 16048
tri -92 16012 -58 16046 ne
rect -58 16037 14948 16046
tri 14948 16037 14957 16046 sw
tri 15018 16037 15027 16046 ne
rect 15027 16037 15079 16046
rect 15080 16038 15081 16094
rect 15117 16038 15118 16094
rect 15119 16037 15354 16095
rect -58 16012 14957 16037
tri 14957 16012 14982 16037 sw
tri 15223 16012 15248 16037 ne
tri -58 16009 -55 16012 ne
rect -55 16009 14982 16012
tri 14982 16009 14985 16012 sw
tri -55 15975 -21 16009 ne
rect -21 15975 14985 16009
tri 14985 15975 15019 16009 sw
tri -21 15973 -19 15975 ne
rect -19 15973 15019 15975
tri 15019 15973 15021 15975 sw
tri -19 15939 15 15973 ne
rect 15 15939 15021 15973
tri 15021 15939 15055 15973 sw
tri 15 15936 18 15939 ne
rect 18 15936 15055 15939
tri 15055 15936 15058 15939 sw
tri 18 15915 39 15936 ne
rect 39 15915 15058 15936
tri 535 15902 548 15915 ne
rect 548 15902 15058 15915
tri 15058 15902 15092 15936 sw
tri 548 15900 550 15902 ne
rect 550 15900 15092 15902
tri 15092 15900 15094 15902 sw
tri 550 15866 584 15900 ne
rect 584 15875 15094 15900
tri 15094 15875 15119 15900 sw
rect 584 15874 15119 15875
rect 584 15866 1240 15874
tri 1240 15866 1248 15874 nw
tri 5315 15866 5323 15874 ne
rect 5323 15866 6001 15874
tri 6001 15866 6009 15874 nw
tri 9999 15866 10007 15874 ne
rect 10007 15866 10731 15874
tri 10731 15866 10739 15874 nw
tri 14849 15866 14857 15874 ne
rect 14857 15866 15119 15874
tri 584 15863 587 15866 ne
rect 587 15863 1237 15866
tri 1237 15863 1240 15866 nw
tri 5323 15863 5326 15866 ne
rect 5326 15863 5998 15866
tri 5998 15863 6001 15866 nw
tri 10007 15863 10010 15866 ne
rect 10010 15863 10728 15866
tri 10728 15863 10731 15866 nw
tri 14857 15863 14860 15866 ne
rect 14860 15863 15119 15866
tri 587 15859 591 15863 ne
rect 591 15859 1203 15863
rect 351 15847 469 15859
rect 351 15813 357 15847
rect 391 15813 429 15847
rect 463 15813 469 15847
tri 591 15829 621 15859 ne
rect 621 15829 1203 15859
tri 1203 15829 1237 15863 nw
tri 5326 15829 5360 15863 ne
rect 5360 15829 5964 15863
tri 5964 15829 5998 15863 nw
tri 10010 15829 10044 15863 ne
rect 10044 15829 10694 15863
tri 10694 15829 10728 15863 nw
tri 14860 15829 14894 15863 ne
rect 14894 15829 15119 15863
tri 621 15827 623 15829 ne
rect 623 15827 1201 15829
tri 1201 15827 1203 15829 nw
tri 5360 15827 5362 15829 ne
rect 5362 15827 5962 15829
tri 5962 15827 5964 15829 nw
tri 10044 15827 10046 15829 ne
rect 10046 15827 10692 15829
tri 10692 15827 10694 15829 nw
tri 14894 15827 14896 15829 ne
rect 14896 15827 15119 15829
rect 351 15773 469 15813
tri 623 15793 657 15827 ne
rect 657 15793 1167 15827
tri 1167 15793 1201 15827 nw
tri 5362 15818 5371 15827 ne
rect 5371 15818 5928 15827
tri 657 15790 660 15793 ne
rect 660 15790 1164 15793
tri 1164 15790 1167 15793 nw
rect 351 15739 357 15773
rect 391 15739 429 15773
rect 463 15739 469 15773
tri 660 15762 688 15790 ne
rect 351 15699 469 15739
rect 351 15665 357 15699
rect 391 15665 429 15699
rect 463 15665 469 15699
rect 351 15625 469 15665
rect 351 15591 357 15625
rect 391 15591 429 15625
rect 463 15591 469 15625
rect 351 15551 469 15591
rect 351 15517 357 15551
rect 391 15517 429 15551
rect 463 15517 469 15551
rect 351 15477 469 15517
rect 351 15443 357 15477
rect 391 15443 429 15477
rect 463 15443 469 15477
rect 351 15403 469 15443
rect 351 15369 357 15403
rect 391 15369 429 15403
rect 463 15369 469 15403
rect 351 15329 469 15369
rect 351 15295 357 15329
rect 391 15295 429 15329
rect 463 15295 469 15329
rect 351 15255 469 15295
rect 688 15756 1130 15790
tri 1130 15756 1164 15790 nw
rect 688 15754 1128 15756
tri 1128 15754 1130 15756 nw
rect 688 15720 1094 15754
tri 1094 15720 1128 15754 nw
rect 688 15355 1092 15720
tri 1092 15718 1094 15720 nw
tri 1092 15355 1114 15377 sw
rect 688 15352 1114 15355
tri 1114 15352 1117 15355 sw
rect 688 15318 1117 15352
tri 1117 15318 1151 15352 sw
rect 688 15316 1151 15318
tri 1151 15316 1153 15318 sw
rect 688 15282 1153 15316
tri 1153 15282 1187 15316 sw
rect 688 15281 1187 15282
tri 1187 15281 1188 15282 sw
tri 688 15279 690 15281 ne
rect 690 15279 1188 15281
tri 1188 15279 1190 15281 sw
rect 351 15221 357 15255
rect 391 15221 429 15255
rect 463 15221 469 15255
tri 690 15245 724 15279 ne
rect 724 15245 1190 15279
tri 1190 15245 1224 15279 sw
rect 2842 15266 3798 15818
tri 5371 15793 5396 15818 ne
rect 5396 15793 5928 15818
tri 5928 15793 5962 15827 nw
tri 10046 15818 10055 15827 ne
rect 10055 15818 10658 15827
tri 5396 15790 5399 15793 ne
rect 5399 15790 5925 15793
tri 5925 15790 5928 15793 nw
tri 5399 15756 5433 15790 ne
rect 5433 15756 5891 15790
tri 5891 15756 5925 15790 nw
tri 5433 15754 5435 15756 ne
rect 5435 15754 5889 15756
tri 5889 15754 5891 15756 nw
tri 5435 15729 5460 15754 ne
tri 5452 15355 5460 15363 se
rect 5460 15355 5864 15754
tri 5864 15729 5889 15754 nw
tri 5864 15355 5872 15363 sw
tri 5449 15352 5452 15355 se
rect 5452 15352 5872 15355
tri 5872 15352 5875 15355 sw
tri 5415 15318 5449 15352 se
rect 5449 15318 5875 15352
tri 5875 15318 5909 15352 sw
tri 5413 15316 5415 15318 se
rect 5415 15316 5909 15318
tri 5909 15316 5911 15318 sw
tri 5379 15282 5413 15316 se
rect 5413 15282 5911 15316
tri 5911 15282 5945 15316 sw
tri 5376 15279 5379 15282 se
rect 5379 15279 5945 15282
tri 5945 15279 5948 15282 sw
tri 2842 15245 2863 15266 ne
rect 2863 15245 3777 15266
tri 3777 15245 3798 15266 nw
tri 5342 15245 5376 15279 se
rect 5376 15245 5948 15279
tri 5948 15245 5982 15279 sw
rect 7526 15266 8482 15818
tri 10055 15793 10080 15818 ne
rect 10080 15793 10658 15818
tri 10658 15793 10692 15827 nw
tri 14896 15818 14905 15827 ne
rect 14905 15818 15119 15827
tri 10080 15790 10083 15793 ne
rect 10083 15790 10655 15793
tri 10655 15790 10658 15793 nw
tri 10083 15756 10117 15790 ne
rect 10117 15756 10621 15790
tri 10621 15756 10655 15790 nw
tri 10117 15754 10119 15756 ne
rect 10119 15754 10619 15756
tri 10619 15754 10621 15756 nw
tri 10119 15729 10144 15754 ne
tri 10136 15355 10144 15363 se
rect 10144 15355 10595 15754
tri 10595 15730 10619 15754 nw
tri 10133 15352 10136 15355 se
rect 10136 15352 10595 15355
tri 10595 15352 10597 15354 sw
tri 10099 15318 10133 15352 se
rect 10133 15318 10597 15352
tri 10597 15318 10631 15352 sw
tri 10097 15316 10099 15318 se
rect 10099 15316 10631 15318
tri 10631 15316 10633 15318 sw
tri 10063 15282 10097 15316 se
rect 10097 15282 10633 15316
tri 10633 15282 10667 15316 sw
rect 12257 15307 13213 15818
tri 14905 15806 14917 15818 ne
rect 12257 15282 13188 15307
tri 13188 15282 13213 15307 nw
tri 14910 15282 14917 15289 se
rect 14917 15282 15119 15818
tri 10060 15279 10063 15282 se
rect 10063 15279 10667 15282
tri 10667 15279 10670 15282 sw
rect 12257 15279 13185 15282
tri 13185 15279 13188 15282 nw
tri 14907 15279 14910 15282 se
rect 14910 15279 15119 15282
tri 7526 15245 7547 15266 ne
rect 7547 15245 8461 15266
tri 8461 15245 8482 15266 nw
tri 10026 15245 10060 15279 se
rect 10060 15245 10670 15279
tri 10670 15245 10704 15279 sw
rect 12257 15266 13151 15279
tri 12257 15245 12278 15266 ne
rect 12278 15245 13151 15266
tri 13151 15245 13185 15279 nw
tri 14873 15245 14907 15279 se
rect 14907 15245 15119 15279
tri 724 15243 726 15245 ne
rect 726 15243 1224 15245
tri 1224 15243 1226 15245 sw
tri 2863 15243 2865 15245 ne
rect 2865 15243 3775 15245
tri 3775 15243 3777 15245 nw
tri 5340 15243 5342 15245 se
rect 5342 15243 5982 15245
tri 5982 15243 5984 15245 sw
tri 7547 15243 7549 15245 ne
rect 7549 15243 8459 15245
tri 8459 15243 8461 15245 nw
tri 10024 15243 10026 15245 se
rect 10026 15243 10704 15245
tri 10704 15243 10706 15245 sw
tri 12278 15243 12280 15245 ne
rect 12280 15243 13149 15245
tri 13149 15243 13151 15245 nw
tri 14871 15243 14873 15245 se
rect 14873 15243 15119 15245
rect 351 15181 469 15221
tri 726 15209 760 15243 ne
rect 760 15210 1226 15243
tri 1226 15210 1259 15243 sw
tri 2865 15210 2898 15243 ne
rect 2898 15210 3742 15243
tri 3742 15210 3775 15243 nw
tri 5307 15210 5340 15243 se
rect 5340 15210 5984 15243
tri 5984 15210 6017 15243 sw
tri 7549 15210 7582 15243 ne
rect 7582 15210 8426 15243
tri 8426 15210 8459 15243 nw
tri 9991 15210 10024 15243 se
rect 10024 15210 10706 15243
tri 10706 15210 10739 15243 sw
tri 12280 15210 12313 15243 ne
rect 12313 15210 13116 15243
tri 13116 15210 13149 15243 nw
tri 14838 15210 14871 15243 se
rect 14871 15211 15119 15243
rect 14871 15210 15118 15211
tri 15118 15210 15119 15211 nw
rect 760 15209 2818 15210
tri 2818 15209 2819 15210 sw
tri 2898 15209 2899 15210 ne
rect 2899 15209 3741 15210
tri 3741 15209 3742 15210 nw
tri 3821 15209 3822 15210 se
rect 3822 15209 7502 15210
tri 7502 15209 7503 15210 sw
tri 7582 15209 7583 15210 ne
rect 7583 15209 8425 15210
tri 8425 15209 8426 15210 nw
tri 8505 15209 8506 15210 se
rect 8506 15209 12186 15210
tri 12186 15209 12187 15210 sw
tri 12313 15209 12314 15210 ne
rect 12314 15209 13115 15210
tri 13115 15209 13116 15210 nw
tri 13195 15209 13196 15210 se
rect 13196 15209 15117 15210
tri 15117 15209 15118 15210 nw
tri 760 15206 763 15209 ne
rect 763 15206 2819 15209
tri 2819 15206 2822 15209 sw
tri 2899 15206 2902 15209 ne
rect 2902 15206 3738 15209
tri 3738 15206 3741 15209 nw
tri 3818 15206 3821 15209 se
rect 3821 15206 7503 15209
tri 7503 15206 7506 15209 sw
tri 7583 15206 7586 15209 ne
rect 7586 15206 8422 15209
tri 8422 15206 8425 15209 nw
tri 8502 15206 8505 15209 se
rect 8505 15206 12187 15209
tri 12187 15206 12190 15209 sw
tri 12314 15206 12317 15209 ne
rect 12317 15206 13112 15209
tri 13112 15206 13115 15209 nw
tri 13192 15206 13195 15209 se
rect 13195 15206 15114 15209
tri 15114 15206 15117 15209 nw
rect 351 15147 357 15181
rect 391 15147 429 15181
rect 463 15147 469 15181
tri 763 15172 797 15206 ne
rect 797 15172 2822 15206
tri 2822 15172 2856 15206 sw
tri 2902 15172 2936 15206 ne
rect 2936 15172 3704 15206
tri 3704 15172 3738 15206 nw
tri 3784 15172 3818 15206 se
rect 3818 15172 7506 15206
tri 7506 15172 7540 15206 sw
tri 7586 15172 7620 15206 ne
rect 7620 15172 8388 15206
tri 8388 15172 8422 15206 nw
tri 8468 15172 8502 15206 se
rect 8502 15172 12190 15206
tri 12190 15172 12224 15206 sw
tri 12317 15172 12351 15206 ne
rect 12351 15172 13078 15206
tri 13078 15172 13112 15206 nw
tri 13158 15172 13192 15206 se
rect 13192 15172 15080 15206
tri 15080 15172 15114 15206 nw
tri 797 15170 799 15172 ne
rect 799 15170 2856 15172
tri 2856 15170 2858 15172 sw
tri 2936 15170 2938 15172 ne
rect 2938 15170 3702 15172
tri 3702 15170 3704 15172 nw
tri 3782 15170 3784 15172 se
rect 3784 15170 7540 15172
tri 7540 15170 7542 15172 sw
tri 7620 15170 7622 15172 ne
rect 7622 15170 8386 15172
tri 8386 15170 8388 15172 nw
tri 8466 15170 8468 15172 se
rect 8468 15170 12224 15172
tri 12224 15170 12226 15172 sw
tri 12351 15170 12353 15172 ne
rect 12353 15170 13076 15172
tri 13076 15170 13078 15172 nw
tri 13156 15170 13158 15172 se
rect 13158 15170 15078 15172
tri 15078 15170 15080 15172 nw
rect 351 15107 469 15147
tri 799 15136 833 15170 ne
rect 833 15136 2858 15170
tri 2858 15136 2892 15170 sw
tri 2938 15136 2972 15170 ne
rect 2972 15136 3668 15170
tri 3668 15136 3702 15170 nw
tri 3748 15136 3782 15170 se
rect 3782 15136 7542 15170
tri 7542 15136 7576 15170 sw
tri 7622 15136 7656 15170 ne
rect 7656 15136 8352 15170
tri 8352 15136 8386 15170 nw
tri 8432 15136 8466 15170 se
rect 8466 15136 12226 15170
tri 12226 15136 12260 15170 sw
tri 12353 15136 12387 15170 ne
rect 12387 15136 13042 15170
tri 13042 15136 13076 15170 nw
tri 13122 15136 13156 15170 se
rect 13156 15136 15044 15170
tri 15044 15136 15078 15170 nw
tri 833 15133 836 15136 ne
rect 836 15133 2892 15136
tri 2892 15133 2895 15136 sw
tri 2972 15133 2975 15136 ne
rect 2975 15133 3665 15136
tri 3665 15133 3668 15136 nw
tri 3745 15133 3748 15136 se
rect 3748 15133 7576 15136
tri 7576 15133 7579 15136 sw
tri 7656 15133 7659 15136 ne
rect 7659 15133 8349 15136
tri 8349 15133 8352 15136 nw
tri 8429 15133 8432 15136 se
rect 8432 15133 12260 15136
tri 12260 15133 12263 15136 sw
tri 12387 15133 12390 15136 ne
rect 12390 15133 13039 15136
tri 13039 15133 13042 15136 nw
tri 13119 15133 13122 15136 se
rect 13122 15133 15041 15136
tri 15041 15133 15044 15136 nw
rect 351 15073 357 15107
rect 391 15073 429 15107
rect 463 15073 469 15107
tri 836 15099 870 15133 ne
rect 870 15130 2895 15133
tri 2895 15130 2898 15133 sw
tri 2975 15130 2978 15133 ne
rect 2978 15130 3662 15133
tri 3662 15130 3665 15133 nw
tri 3742 15130 3745 15133 se
rect 3745 15130 7579 15133
tri 7579 15130 7582 15133 sw
tri 7659 15130 7662 15133 ne
rect 7662 15130 8346 15133
tri 8346 15130 8349 15133 nw
tri 8426 15130 8429 15133 se
rect 8429 15130 12263 15133
rect 870 15126 2898 15130
tri 2898 15126 2902 15130 sw
tri 2978 15126 2982 15130 ne
rect 2982 15126 3658 15130
tri 3658 15126 3662 15130 nw
tri 3738 15126 3742 15130 se
rect 3742 15126 7582 15130
tri 7582 15126 7586 15130 sw
tri 7662 15126 7666 15130 ne
rect 7666 15126 8342 15130
tri 8342 15126 8346 15130 nw
tri 8422 15126 8426 15130 se
rect 8426 15126 12263 15130
rect 870 15099 2902 15126
tri 2902 15099 2929 15126 sw
tri 2982 15099 3009 15126 ne
rect 3009 15099 3631 15126
tri 3631 15099 3658 15126 nw
tri 3711 15099 3738 15126 se
rect 3738 15099 7586 15126
tri 7586 15099 7613 15126 sw
tri 7666 15099 7693 15126 ne
rect 7693 15099 8315 15126
tri 8315 15099 8342 15126 nw
tri 8395 15099 8422 15126 se
rect 8422 15099 12263 15126
tri 12263 15099 12297 15133 sw
tri 12390 15099 12424 15133 ne
rect 12424 15130 13036 15133
tri 13036 15130 13039 15133 nw
tri 13116 15130 13119 15133 se
rect 13119 15130 15007 15133
rect 12424 15129 13035 15130
tri 13035 15129 13036 15130 nw
tri 13115 15129 13116 15130 se
rect 13116 15129 15007 15130
rect 12424 15099 13005 15129
tri 13005 15099 13035 15129 nw
tri 13085 15099 13115 15129 se
rect 13115 15099 15007 15129
tri 15007 15099 15041 15133 nw
tri 870 15097 872 15099 ne
rect 872 15097 2929 15099
tri 2929 15097 2931 15099 sw
tri 3009 15097 3011 15099 ne
rect 3011 15097 3629 15099
tri 3629 15097 3631 15099 nw
tri 3709 15097 3711 15099 se
rect 3711 15097 7613 15099
tri 7613 15097 7615 15099 sw
tri 7693 15097 7695 15099 ne
rect 7695 15097 8313 15099
tri 8313 15097 8315 15099 nw
tri 8393 15097 8395 15099 se
rect 8395 15097 12297 15099
tri 12297 15097 12299 15099 sw
tri 12424 15097 12426 15099 ne
rect 12426 15097 13003 15099
tri 13003 15097 13005 15099 nw
tri 13083 15097 13085 15099 se
rect 13085 15097 15005 15099
tri 15005 15097 15007 15099 nw
rect 351 15033 469 15073
tri 872 15063 906 15097 ne
rect 906 15063 2931 15097
tri 2931 15063 2965 15097 sw
tri 3011 15063 3045 15097 ne
rect 3045 15063 3595 15097
tri 3595 15063 3629 15097 nw
tri 3675 15063 3709 15097 se
rect 3709 15063 7615 15097
tri 7615 15063 7649 15097 sw
tri 7695 15063 7729 15097 ne
rect 7729 15063 8279 15097
tri 8279 15063 8313 15097 nw
tri 8359 15063 8393 15097 se
rect 8393 15083 12299 15097
tri 12299 15083 12313 15097 sw
tri 12426 15083 12440 15097 ne
rect 12440 15083 12969 15097
rect 8393 15063 12313 15083
tri 12313 15063 12333 15083 sw
tri 12440 15063 12460 15083 ne
rect 12460 15063 12969 15083
tri 12969 15063 13003 15097 nw
tri 13049 15063 13083 15097 se
rect 13083 15063 14971 15097
tri 14971 15063 15005 15097 nw
tri 15234 15063 15248 15077 se
rect 15248 15063 15354 16037
tri 906 15060 909 15063 ne
rect 909 15060 2965 15063
tri 2965 15060 2968 15063 sw
tri 3045 15060 3048 15063 ne
rect 3048 15060 3592 15063
tri 3592 15060 3595 15063 nw
tri 3672 15060 3675 15063 se
rect 3675 15060 7649 15063
tri 7649 15060 7652 15063 sw
tri 7729 15060 7732 15063 ne
rect 7732 15060 8276 15063
tri 8276 15060 8279 15063 nw
tri 8356 15060 8359 15063 se
rect 8359 15060 12333 15063
tri 12333 15060 12336 15063 sw
tri 12460 15060 12463 15063 ne
rect 12463 15060 12966 15063
tri 12966 15060 12969 15063 nw
tri 13046 15060 13049 15063 se
rect 13049 15060 14968 15063
tri 14968 15060 14971 15063 nw
tri 15231 15060 15234 15063 se
rect 15234 15060 15354 15063
rect 351 14999 357 15033
rect 391 14999 429 15033
rect 463 14999 469 15033
tri 909 15026 943 15060 ne
rect 943 15046 2968 15060
tri 2968 15046 2982 15060 sw
tri 3048 15046 3062 15060 ne
rect 3062 15046 3578 15060
tri 3578 15046 3592 15060 nw
tri 3658 15046 3672 15060 se
rect 3672 15046 7652 15060
tri 7652 15046 7666 15060 sw
tri 7732 15046 7746 15060 ne
rect 7746 15046 8262 15060
tri 8262 15046 8276 15060 nw
tri 8342 15046 8356 15060 se
rect 8356 15046 12336 15060
rect 943 15026 2982 15046
tri 2982 15026 3002 15046 sw
tri 3062 15026 3082 15046 ne
rect 3082 15026 3558 15046
tri 3558 15026 3578 15046 nw
tri 3638 15026 3658 15046 se
rect 3658 15026 7666 15046
tri 7666 15026 7686 15046 sw
tri 7746 15026 7766 15046 ne
rect 7766 15026 8242 15046
tri 8242 15026 8262 15046 nw
tri 8322 15026 8342 15046 se
rect 8342 15026 12336 15046
tri 12336 15026 12370 15060 sw
tri 12463 15026 12497 15060 ne
rect 12497 15049 12955 15060
tri 12955 15049 12966 15060 nw
tri 13038 15052 13046 15060 se
rect 13046 15052 14960 15060
tri 14960 15052 14968 15060 nw
tri 15223 15052 15231 15060 se
rect 15231 15052 15354 15060
tri 13035 15049 13038 15052 se
rect 13038 15049 14934 15052
rect 12497 15026 12937 15049
tri 12937 15031 12955 15049 nw
tri 943 15024 945 15026 ne
rect 945 15024 3002 15026
tri 3002 15024 3004 15026 sw
tri 3082 15024 3084 15026 ne
rect 3084 15024 3556 15026
tri 3556 15024 3558 15026 nw
tri 3636 15024 3638 15026 se
rect 3638 15024 7686 15026
tri 7686 15024 7688 15026 sw
tri 7766 15024 7768 15026 ne
rect 7768 15024 8240 15026
tri 8240 15024 8242 15026 nw
tri 8320 15024 8322 15026 se
rect 8322 15024 12370 15026
tri 12370 15024 12372 15026 sw
tri 12497 15024 12499 15026 ne
rect 12499 15024 12937 15026
rect 351 14959 469 14999
tri 945 14990 979 15024 ne
rect 979 14990 3004 15024
tri 3004 14990 3038 15024 sw
tri 3084 14990 3118 15024 ne
tri 979 14987 982 14990 ne
rect 982 14987 3038 14990
tri 3038 14987 3041 14990 sw
tri 982 14976 993 14987 ne
rect 993 14976 3041 14987
tri 3041 14976 3052 14987 sw
rect 351 14925 357 14959
rect 391 14925 429 14959
rect 463 14925 469 14959
tri 993 14942 1027 14976 ne
rect 1027 14966 3052 14976
tri 3052 14966 3062 14976 sw
rect 1027 14942 3062 14966
rect 351 14885 469 14925
tri 1027 14917 1052 14942 ne
rect 1052 14917 3062 14942
tri 1052 14914 1055 14917 ne
rect 1055 14914 3062 14917
rect 351 14851 357 14885
rect 391 14851 429 14885
rect 463 14851 469 14885
tri 1055 14880 1089 14914 ne
rect 1089 14880 3062 14914
tri 1089 14870 1099 14880 ne
rect 1099 14870 3062 14880
rect 351 14811 469 14851
tri 1099 14844 1125 14870 ne
rect 1125 14844 3062 14870
tri 1125 14841 1128 14844 ne
rect 1128 14841 3062 14844
tri 1128 14838 1131 14841 ne
rect 1131 14838 3062 14841
rect 351 14777 357 14811
rect 391 14777 429 14811
rect 463 14777 469 14811
tri 1131 14804 1165 14838 ne
rect 1165 14804 3062 14838
tri 1165 14781 1188 14804 ne
rect 1188 14781 3062 14804
rect 351 14737 469 14777
tri 1188 14771 1198 14781 ne
rect 1198 14771 3062 14781
tri 1198 14768 1201 14771 ne
rect 1201 14768 3062 14771
tri 1201 14761 1208 14768 ne
rect 1208 14761 3062 14768
tri 1208 14758 1211 14761 ne
rect 1211 14758 3062 14761
rect 351 14703 357 14737
rect 391 14703 429 14737
rect 463 14703 469 14737
rect 351 14663 469 14703
rect 351 14629 357 14663
rect 391 14629 429 14663
rect 463 14629 469 14663
rect 351 14589 469 14629
rect 351 14555 357 14589
rect 391 14555 429 14589
rect 463 14555 469 14589
rect 351 14515 469 14555
rect 351 14481 357 14515
rect 391 14481 429 14515
rect 463 14481 469 14515
rect 351 14441 469 14481
rect 351 14407 357 14441
rect 391 14407 429 14441
rect 463 14407 469 14441
rect 351 14367 469 14407
rect 351 14333 357 14367
rect 391 14333 429 14367
rect 463 14333 469 14367
rect 351 14293 469 14333
rect 351 14259 357 14293
rect 391 14259 429 14293
rect 463 14259 469 14293
rect 351 14219 469 14259
rect 351 14185 357 14219
rect 391 14185 429 14219
rect 463 14185 469 14219
rect 351 14145 469 14185
rect 351 14111 357 14145
rect 391 14111 429 14145
rect 463 14111 469 14145
rect 351 14071 469 14111
rect 351 14037 357 14071
rect 391 14037 429 14071
rect 463 14037 469 14071
rect 351 13997 469 14037
rect 351 13963 357 13997
rect 391 13963 429 13997
rect 463 13963 469 13997
rect 351 13923 469 13963
rect 351 13889 357 13923
rect 391 13889 429 13923
rect 463 13889 469 13923
rect 351 13850 469 13889
rect 351 13816 357 13850
rect 391 13816 429 13850
rect 463 13816 469 13850
rect 351 13777 469 13816
rect 351 13743 357 13777
rect 391 13743 429 13777
rect 463 13743 469 13777
rect 351 13704 469 13743
rect 351 13670 357 13704
rect 391 13670 429 13704
rect 463 13670 469 13704
rect 351 13631 469 13670
rect 351 13597 357 13631
rect 391 13597 429 13631
rect 463 13597 469 13631
rect 351 13558 469 13597
rect 351 13524 357 13558
rect 391 13524 429 13558
rect 463 13524 469 13558
rect 351 13485 469 13524
rect 351 13451 357 13485
rect 391 13451 429 13485
rect 463 13451 469 13485
rect 351 13412 469 13451
rect 351 13378 357 13412
rect 391 13378 429 13412
rect 463 13378 469 13412
rect 351 13339 469 13378
rect 351 13305 357 13339
rect 391 13305 429 13339
rect 463 13305 469 13339
rect 351 13266 469 13305
rect 351 13232 357 13266
rect 391 13232 429 13266
rect 463 13232 469 13266
rect 351 13193 469 13232
rect 351 13159 357 13193
rect 391 13159 429 13193
rect 463 13159 469 13193
rect 351 13120 469 13159
rect 351 13086 357 13120
rect 391 13086 429 13120
rect 463 13086 469 13120
rect 351 13047 469 13086
rect 351 13013 357 13047
rect 391 13013 429 13047
rect 463 13013 469 13047
rect 351 12974 469 13013
rect 351 12940 357 12974
rect 391 12940 429 12974
rect 463 12940 469 12974
rect 351 12901 469 12940
rect 351 12867 357 12901
rect 391 12867 429 12901
rect 463 12867 469 12901
rect 351 12828 469 12867
rect 351 12794 357 12828
rect 391 12794 429 12828
rect 463 12794 469 12828
rect 351 12755 469 12794
rect 351 12721 357 12755
rect 391 12721 429 12755
rect 463 12721 469 12755
rect 351 12682 469 12721
rect 351 12648 357 12682
rect 391 12648 429 12682
rect 463 12648 469 12682
rect 351 12609 469 12648
rect 351 12575 357 12609
rect 391 12575 429 12609
rect 463 12575 469 12609
rect 351 12536 469 12575
rect 674 14746 792 14758
rect 674 14712 680 14746
rect 714 14712 752 14746
rect 786 14712 792 14746
tri 1211 14733 1236 14758 ne
rect 1236 14733 3062 14758
rect 3118 14914 3522 15024
tri 3522 14990 3556 15024 nw
tri 3602 14990 3636 15024 se
rect 3636 14990 7688 15024
tri 7688 14990 7722 15024 sw
tri 7768 14990 7802 15024 ne
tri 3599 14987 3602 14990 se
rect 3602 14987 7722 14990
tri 7722 14987 7725 14990 sw
tri 3588 14976 3599 14987 se
rect 3599 14976 7725 14987
tri 7725 14976 7736 14987 sw
rect 3118 14880 3267 14914
rect 3301 14880 3339 14914
rect 3373 14880 3522 14914
rect 3118 14838 3522 14880
rect 3118 14804 3267 14838
rect 3301 14804 3339 14838
rect 3373 14804 3522 14838
rect 3118 14761 3522 14804
rect 674 14671 792 14712
rect 674 14637 680 14671
rect 714 14637 752 14671
rect 786 14637 792 14671
rect 674 14596 792 14637
rect 674 14562 680 14596
rect 714 14562 752 14596
rect 786 14562 792 14596
rect 674 14521 792 14562
rect 674 14487 680 14521
rect 714 14487 752 14521
rect 786 14487 792 14521
rect 674 14446 792 14487
rect 674 14412 680 14446
rect 714 14412 752 14446
rect 786 14412 792 14446
rect 674 14371 792 14412
rect 674 14337 680 14371
rect 714 14337 752 14371
rect 786 14337 792 14371
rect 674 14296 792 14337
rect 674 14262 680 14296
rect 714 14262 752 14296
rect 786 14262 792 14296
rect 674 14221 792 14262
rect 674 14187 680 14221
rect 714 14187 752 14221
rect 786 14187 792 14221
rect 674 14150 792 14187
rect 3118 14727 3267 14761
rect 3301 14727 3339 14761
rect 3373 14727 3522 14761
tri 3578 14966 3588 14976 se
rect 3588 14966 7736 14976
tri 7736 14966 7746 14976 sw
rect 3578 14785 7746 14966
rect 3578 14771 5442 14785
tri 5442 14771 5456 14785 nw
tri 5868 14771 5882 14785 ne
rect 5882 14771 7746 14785
rect 3578 14768 5439 14771
tri 5439 14768 5442 14771 nw
tri 5882 14768 5885 14771 ne
rect 5885 14768 7746 14771
rect 3578 14761 5432 14768
tri 5432 14761 5439 14768 nw
tri 5885 14761 5892 14768 ne
rect 5892 14761 7746 14768
rect 3578 14733 5404 14761
tri 5404 14733 5432 14761 nw
tri 5892 14733 5920 14761 ne
rect 5920 14733 7746 14761
rect 7802 14914 8206 15024
tri 8206 14990 8240 15024 nw
tri 8286 14990 8320 15024 se
rect 8320 14990 12372 15024
tri 12372 14990 12406 15024 sw
tri 12499 14990 12533 15024 ne
tri 8283 14987 8286 14990 se
rect 8286 14987 12406 14990
tri 12406 14987 12409 14990 sw
tri 8272 14976 8283 14987 se
rect 8283 14976 12409 14987
tri 12409 14976 12420 14987 sw
rect 7802 14880 7951 14914
rect 7985 14880 8023 14914
rect 8057 14880 8206 14914
rect 7802 14838 8206 14880
rect 7802 14804 7951 14838
rect 7985 14804 8023 14838
rect 8057 14804 8206 14838
rect 7802 14761 8206 14804
rect 3118 14684 3522 14727
rect 3118 14650 3267 14684
rect 3301 14650 3339 14684
rect 3373 14650 3522 14684
rect 3118 14607 3522 14650
rect 3118 14573 3267 14607
rect 3301 14573 3339 14607
rect 3373 14573 3522 14607
rect 3118 14530 3522 14573
rect 3118 14496 3267 14530
rect 3301 14496 3339 14530
rect 3373 14496 3522 14530
rect 3118 14453 3522 14496
rect 3118 14419 3267 14453
rect 3301 14419 3339 14453
rect 3373 14419 3522 14453
rect 3118 14376 3522 14419
rect 3118 14342 3267 14376
rect 3301 14342 3339 14376
rect 3373 14342 3522 14376
rect 3118 14299 3522 14342
rect 3118 14265 3267 14299
rect 3301 14265 3339 14299
rect 3373 14265 3522 14299
rect 3118 14222 3522 14265
rect 3118 14188 3267 14222
rect 3301 14188 3339 14222
rect 3373 14188 3522 14222
tri 792 14150 799 14157 sw
rect 674 14146 799 14150
rect 674 14112 680 14146
rect 714 14112 752 14146
rect 786 14145 799 14146
tri 799 14145 804 14150 sw
rect 3118 14145 3522 14188
rect 786 14112 804 14145
rect 674 14111 804 14112
tri 804 14111 838 14145 sw
rect 3118 14111 3267 14145
rect 3301 14111 3339 14145
rect 3373 14133 3522 14145
rect 5603 14717 5721 14729
rect 5603 14683 5609 14717
rect 5643 14683 5681 14717
rect 5715 14683 5721 14717
rect 5603 14644 5721 14683
rect 5603 14610 5609 14644
rect 5643 14610 5681 14644
rect 5715 14610 5721 14644
rect 5603 14571 5721 14610
rect 5603 14537 5609 14571
rect 5643 14537 5681 14571
rect 5715 14537 5721 14571
rect 5603 14498 5721 14537
rect 5603 14464 5609 14498
rect 5643 14464 5681 14498
rect 5715 14464 5721 14498
rect 5603 14425 5721 14464
rect 5603 14391 5609 14425
rect 5643 14391 5681 14425
rect 5715 14391 5721 14425
rect 5603 14352 5721 14391
rect 5603 14318 5609 14352
rect 5643 14318 5681 14352
rect 5715 14318 5721 14352
rect 5603 14279 5721 14318
rect 5603 14245 5609 14279
rect 5643 14245 5681 14279
rect 5715 14245 5721 14279
rect 5603 14206 5721 14245
rect 5603 14172 5609 14206
rect 5643 14172 5681 14206
rect 5715 14172 5721 14206
tri 3522 14133 3533 14144 sw
rect 5603 14133 5721 14172
rect 7802 14727 7951 14761
rect 7985 14727 8023 14761
rect 8057 14727 8206 14761
tri 8262 14966 8272 14976 se
rect 8272 14966 12420 14976
tri 12420 14966 12430 14976 sw
rect 8262 14942 12430 14966
tri 12430 14942 12454 14966 sw
rect 8262 14919 12454 14942
tri 12454 14919 12477 14942 sw
rect 8262 14785 12477 14919
rect 8262 14771 10126 14785
tri 10126 14771 10140 14785 nw
tri 10599 14771 10613 14785 ne
rect 10613 14771 12477 14785
rect 8262 14768 10123 14771
tri 10123 14768 10126 14771 nw
tri 10613 14768 10616 14771 ne
rect 10616 14768 12477 14771
rect 8262 14761 10116 14768
tri 10116 14761 10123 14768 nw
tri 10616 14761 10623 14768 ne
rect 10623 14761 12477 14768
rect 8262 14733 10088 14761
tri 10088 14733 10116 14761 nw
tri 10623 14733 10651 14761 ne
rect 10651 14733 12477 14761
rect 12533 14914 12937 15024
rect 12533 14880 12682 14914
rect 12716 14880 12754 14914
rect 12788 14880 12937 14914
rect 12533 14838 12937 14880
rect 12533 14804 12682 14838
rect 12716 14804 12754 14838
rect 12788 14804 12937 14838
rect 12533 14761 12937 14804
rect 13035 15026 14934 15049
tri 14934 15026 14960 15052 nw
tri 15014 15026 15040 15052 se
rect 15040 15026 15092 15052
rect 15094 15051 15130 15052
rect 13035 15024 14932 15026
tri 14932 15024 14934 15026 nw
tri 15012 15024 15014 15026 se
rect 15014 15024 15092 15026
rect 13035 14990 14898 15024
tri 14898 14990 14932 15024 nw
tri 14980 14992 15012 15024 se
rect 15012 14994 15092 15024
rect 15093 14995 15131 15051
rect 15094 14994 15130 14995
rect 15132 14994 15354 15052
rect 15012 14992 15074 14994
rect 14980 14990 15074 14992
tri 15074 14990 15078 14994 nw
tri 15223 14990 15227 14994 ne
rect 15227 14990 15354 14994
rect 13035 14987 14895 14990
tri 14895 14987 14898 14990 nw
rect 14980 14987 15071 14990
tri 15071 14987 15074 14990 nw
tri 15227 14987 15230 14990 ne
rect 15230 14987 15354 14990
rect 13035 14976 14884 14987
tri 14884 14976 14895 14987 nw
rect 14980 14976 15053 14987
rect 13035 14953 14861 14976
tri 14861 14953 14884 14976 nw
rect 13036 14951 14860 14952
rect 13035 14895 14861 14951
rect 13036 14894 14860 14895
rect 13035 14841 14861 14893
rect 14980 14942 14986 14976
rect 15020 14942 15053 14976
tri 15053 14969 15071 14987 nw
tri 15230 14969 15248 14987 ne
rect 15248 14969 15354 14987
tri 15248 14955 15262 14969 ne
rect 14980 14917 15053 14942
tri 15053 14917 15077 14941 sw
rect 14980 14916 15077 14917
tri 15077 14916 15078 14917 sw
rect 14980 14904 15078 14916
rect 14980 14870 14986 14904
rect 15020 14870 15078 14904
rect 14980 14858 15078 14870
rect 15079 14859 15080 14915
rect 15116 14859 15117 14915
rect 15118 14910 15205 14916
rect 15118 14876 15159 14910
rect 15193 14876 15205 14910
rect 15118 14858 15205 14876
tri 15117 14844 15131 14858 ne
rect 15131 14844 15205 14858
tri 15131 14841 15134 14844 ne
rect 15134 14841 15205 14844
rect 13035 14776 13079 14841
tri 15134 14838 15137 14841 ne
rect 15137 14838 15205 14841
tri 15137 14828 15147 14838 ne
rect 15147 14804 15159 14838
rect 15193 14804 15205 14838
rect 15147 14798 15205 14804
rect 7802 14684 8206 14727
rect 7802 14650 7951 14684
rect 7985 14650 8023 14684
rect 8057 14650 8206 14684
rect 7802 14607 8206 14650
rect 7802 14573 7951 14607
rect 7985 14573 8023 14607
rect 8057 14573 8206 14607
rect 7802 14530 8206 14573
rect 7802 14496 7951 14530
rect 7985 14496 8023 14530
rect 8057 14496 8206 14530
rect 7802 14453 8206 14496
rect 7802 14419 7951 14453
rect 7985 14419 8023 14453
rect 8057 14419 8206 14453
rect 7802 14376 8206 14419
rect 7802 14342 7951 14376
rect 7985 14342 8023 14376
rect 8057 14342 8206 14376
rect 7802 14299 8206 14342
rect 7802 14265 7951 14299
rect 7985 14265 8023 14299
rect 8057 14265 8206 14299
rect 7802 14222 8206 14265
rect 7802 14188 7951 14222
rect 7985 14188 8023 14222
rect 8057 14188 8206 14222
rect 7802 14145 8206 14188
rect 3373 14111 3533 14133
rect 674 14099 838 14111
tri 838 14099 850 14111 sw
rect 3118 14099 3533 14111
tri 3533 14099 3567 14133 sw
rect 5603 14099 5609 14133
rect 5643 14099 5681 14133
rect 5715 14099 5721 14133
tri 7769 14111 7802 14144 se
rect 7802 14111 7951 14145
rect 7985 14111 8023 14145
rect 8057 14133 8206 14145
rect 10287 14717 10405 14729
rect 10287 14683 10293 14717
rect 10327 14683 10365 14717
rect 10399 14683 10405 14717
rect 10287 14644 10405 14683
rect 10287 14610 10293 14644
rect 10327 14610 10365 14644
rect 10399 14610 10405 14644
rect 10287 14571 10405 14610
rect 10287 14537 10293 14571
rect 10327 14537 10365 14571
rect 10399 14537 10405 14571
rect 10287 14498 10405 14537
rect 10287 14464 10293 14498
rect 10327 14464 10365 14498
rect 10399 14464 10405 14498
rect 10287 14425 10405 14464
rect 10287 14391 10293 14425
rect 10327 14391 10365 14425
rect 10399 14391 10405 14425
rect 10287 14352 10405 14391
rect 10287 14318 10293 14352
rect 10327 14318 10365 14352
rect 10399 14318 10405 14352
rect 10287 14279 10405 14318
rect 10287 14245 10293 14279
rect 10327 14245 10365 14279
rect 10399 14245 10405 14279
rect 10287 14206 10405 14245
rect 10287 14172 10293 14206
rect 10327 14172 10365 14206
rect 10399 14172 10405 14206
tri 8206 14133 8217 14144 sw
rect 10287 14133 10405 14172
rect 8057 14111 8217 14133
tri 7757 14099 7769 14111 se
rect 7769 14099 8217 14111
tri 8217 14099 8251 14133 sw
rect 10287 14099 10293 14133
rect 10327 14099 10365 14133
rect 10399 14099 10405 14133
rect 674 14077 850 14099
tri 850 14077 872 14099 sw
tri 3103 14077 3118 14092 se
rect 3118 14077 3567 14099
tri 3567 14077 3589 14099 sw
rect 674 14071 872 14077
rect 674 14037 680 14071
rect 714 14037 752 14071
rect 786 14068 872 14071
tri 872 14068 881 14077 sw
tri 3094 14068 3103 14077 se
rect 3103 14068 3589 14077
tri 3589 14068 3598 14077 sw
tri 5600 14068 5603 14071 se
rect 5603 14068 5721 14099
tri 7735 14077 7757 14099 se
rect 7757 14077 8251 14099
tri 8251 14077 8273 14099 sw
tri 7728 14070 7735 14077 se
rect 7735 14070 8273 14077
tri 5721 14068 5723 14070 sw
tri 7726 14068 7728 14070 se
rect 7728 14068 8273 14070
tri 8273 14068 8282 14077 sw
tri 10284 14068 10287 14071 se
rect 10287 14068 10405 14099
rect 12533 14727 12682 14761
rect 12716 14727 12754 14761
rect 12788 14727 12937 14761
rect 12533 14684 12937 14727
rect 12533 14650 12682 14684
rect 12716 14650 12754 14684
rect 12788 14650 12937 14684
rect 12533 14607 12937 14650
rect 12533 14573 12682 14607
rect 12716 14573 12754 14607
rect 12788 14573 12937 14607
rect 12533 14530 12937 14573
rect 12533 14496 12682 14530
rect 12716 14496 12754 14530
rect 12788 14496 12937 14530
rect 12533 14453 12937 14496
rect 12533 14419 12682 14453
rect 12716 14419 12754 14453
rect 12788 14419 12937 14453
rect 14980 14643 15026 14655
rect 14980 14609 14986 14643
rect 15020 14609 15026 14643
rect 15147 14637 15205 14643
rect 14980 14603 15026 14609
tri 15026 14603 15058 14635 sw
tri 15138 14603 15147 14612 se
rect 15147 14603 15159 14637
rect 15193 14603 15205 14637
rect 14980 14588 15058 14603
tri 15058 14588 15073 14603 sw
tri 15123 14588 15138 14603 se
rect 15138 14588 15205 14603
rect 14980 14584 15073 14588
tri 15073 14584 15077 14588 sw
tri 15119 14584 15123 14588 se
rect 15123 14584 15205 14588
rect 14980 14583 15077 14584
tri 15077 14583 15078 14584 sw
tri 15118 14583 15119 14584 se
rect 15119 14583 15205 14584
rect 14980 14571 15078 14583
rect 14980 14537 14986 14571
rect 15020 14537 15078 14571
rect 14980 14525 15078 14537
rect 15079 14526 15080 14582
rect 15116 14526 15117 14582
rect 15118 14565 15205 14583
rect 15118 14531 15159 14565
rect 15193 14531 15205 14565
rect 15118 14525 15205 14531
rect 14980 14515 15068 14525
tri 15068 14515 15078 14525 nw
rect 14980 14510 15063 14515
tri 15063 14510 15068 14515 nw
rect 14980 14449 15053 14510
tri 15053 14500 15063 14510 nw
tri 15252 14476 15262 14486 se
rect 15262 14476 15354 14969
tri 15248 14472 15252 14476 se
rect 15252 14472 15354 14476
tri 14980 14442 14987 14449 ne
rect 14987 14447 15053 14449
tri 15053 14447 15078 14472 sw
tri 15223 14447 15248 14472 se
rect 15248 14447 15354 14472
rect 14987 14442 15092 14447
rect 15094 14446 15130 14447
tri 14987 14436 14993 14442 ne
rect 14993 14436 15092 14442
rect 12533 14376 12937 14419
tri 14993 14402 15027 14436 ne
rect 15027 14402 15092 14436
tri 15027 14389 15040 14402 ne
rect 15040 14389 15092 14402
rect 15093 14390 15131 14446
rect 15094 14389 15130 14390
rect 15132 14389 15354 14447
rect 12533 14342 12682 14376
rect 12716 14342 12754 14376
rect 12788 14342 12937 14376
tri 15211 14369 15231 14389 ne
rect 15231 14369 15354 14389
tri 15231 14364 15236 14369 ne
rect 12533 14299 12937 14342
rect 12533 14265 12682 14299
rect 12716 14265 12754 14299
rect 12788 14265 12937 14299
rect 12533 14222 12937 14265
rect 12533 14188 12682 14222
rect 12716 14188 12754 14222
rect 12788 14188 12937 14222
rect 12533 14180 12937 14188
tri 12937 14180 12965 14208 sw
rect 12533 14150 12965 14180
tri 12965 14150 12995 14180 sw
rect 12533 14145 12995 14150
rect 12533 14111 12682 14145
rect 12716 14111 12754 14145
rect 12788 14140 12995 14145
tri 12995 14140 13005 14150 sw
rect 12788 14111 13005 14140
rect 12533 14106 13005 14111
tri 13005 14106 13039 14140 sw
tri 12518 14077 12533 14092 se
rect 12533 14077 13039 14106
tri 13039 14077 13068 14106 sw
tri 12510 14069 12518 14077 se
rect 12518 14069 13068 14077
tri 10405 14068 10406 14069 sw
tri 12509 14068 12510 14069 se
rect 12510 14068 13068 14069
rect 786 14037 881 14068
rect 674 14034 881 14037
tri 881 14034 915 14068 sw
tri 3060 14034 3094 14068 se
rect 3094 14034 3267 14068
rect 3301 14034 3339 14068
rect 3373 14060 3598 14068
tri 3598 14060 3606 14068 sw
tri 5592 14060 5600 14068 se
rect 5600 14060 5723 14068
rect 3373 14034 3606 14060
rect 674 14026 915 14034
tri 915 14026 923 14034 sw
tri 3052 14026 3060 14034 se
rect 3060 14026 3606 14034
tri 3606 14026 3640 14060 sw
tri 5558 14026 5592 14060 se
rect 5592 14026 5609 14060
rect 5643 14026 5681 14060
rect 5715 14034 5723 14060
tri 5723 14034 5757 14068 sw
tri 7692 14034 7726 14068 se
rect 7726 14034 7951 14068
rect 7985 14034 8023 14068
rect 8057 14060 8282 14068
tri 8282 14060 8290 14068 sw
tri 10276 14060 10284 14068 se
rect 10284 14060 10406 14068
rect 8057 14034 8290 14060
rect 5715 14026 5757 14034
tri 5757 14026 5765 14034 sw
tri 7684 14026 7692 14034 se
rect 7692 14026 8290 14034
tri 8290 14026 8324 14060 sw
tri 10242 14026 10276 14060 se
rect 10276 14026 10293 14060
rect 10327 14026 10365 14060
rect 10399 14034 10406 14060
tri 10406 14034 10440 14068 sw
tri 12475 14034 12509 14068 se
rect 12509 14034 12682 14068
rect 12716 14034 12754 14068
rect 12788 14066 13068 14068
tri 13068 14066 13079 14077 sw
rect 12788 14049 13079 14066
tri 13079 14049 13096 14066 sw
rect 12788 14034 15113 14049
rect 10399 14032 10440 14034
tri 10440 14032 10442 14034 sw
tri 12473 14032 12475 14034 se
rect 12475 14032 15113 14034
tri 15113 14032 15130 14049 sw
rect 15236 14037 15354 14369
rect 15390 16450 15396 16484
rect 15430 16450 15628 16484
rect 15390 16411 15628 16450
rect 15390 16377 15396 16411
rect 15430 16377 15628 16411
rect 15390 16338 15628 16377
rect 15390 16304 15396 16338
rect 15430 16304 15628 16338
rect 15390 16265 15628 16304
rect 15390 16231 15396 16265
rect 15430 16231 15628 16265
rect 15390 16212 15628 16231
rect 15390 16194 15610 16212
tri 15610 16194 15628 16212 nw
rect 17942 16851 17948 16885
rect 17982 16851 18060 16885
rect 17942 16848 18060 16851
rect 17942 16814 18020 16848
rect 18054 16814 18060 16848
rect 17942 16812 18060 16814
rect 17942 16778 17948 16812
rect 17982 16778 18060 16812
rect 17942 16776 18060 16778
rect 17942 16742 18020 16776
rect 18054 16742 18060 16776
rect 17942 16739 18060 16742
rect 17942 16705 17948 16739
rect 17982 16705 18060 16739
rect 17942 16704 18060 16705
rect 17942 16670 18020 16704
rect 18054 16670 18060 16704
rect 17942 16666 18060 16670
rect 17942 16632 17948 16666
rect 17982 16632 18060 16666
rect 17942 16598 18020 16632
rect 18054 16598 18060 16632
rect 17942 16593 18060 16598
rect 17942 16559 17948 16593
rect 17982 16559 18060 16593
rect 17942 16525 18020 16559
rect 18054 16525 18060 16559
rect 17942 16520 18060 16525
rect 17942 16486 17948 16520
rect 17982 16486 18060 16520
rect 17942 16452 18020 16486
rect 18054 16452 18060 16486
rect 17942 16447 18060 16452
rect 17942 16413 17948 16447
rect 17982 16413 18060 16447
rect 17942 16379 18020 16413
rect 18054 16379 18060 16413
rect 17942 16374 18060 16379
rect 17942 16340 17948 16374
rect 17982 16340 18060 16374
rect 17942 16306 18020 16340
rect 18054 16306 18060 16340
rect 17942 16301 18060 16306
rect 17942 16267 17948 16301
rect 17982 16267 18060 16301
rect 17942 16233 18020 16267
rect 18054 16233 18060 16267
rect 17942 16228 18060 16233
rect 17942 16194 17948 16228
rect 17982 16194 18060 16228
rect 15390 16192 15576 16194
rect 15390 16158 15396 16192
rect 15430 16160 15576 16192
tri 15576 16160 15610 16194 nw
rect 17942 16160 18020 16194
rect 18054 16160 18060 16194
rect 15430 16158 15571 16160
rect 15390 16155 15571 16158
tri 15571 16155 15576 16160 nw
rect 17942 16155 18060 16160
rect 15390 16121 15537 16155
tri 15537 16121 15571 16155 nw
rect 17942 16121 17948 16155
rect 17982 16121 18060 16155
rect 15390 16119 15503 16121
rect 15390 16085 15396 16119
rect 15430 16087 15503 16119
tri 15503 16087 15537 16121 nw
rect 17942 16087 18020 16121
rect 18054 16087 18060 16121
rect 15430 16085 15498 16087
rect 15390 16046 15498 16085
tri 15498 16082 15503 16087 nw
rect 17942 16082 18060 16087
rect 15390 16012 15396 16046
rect 15430 16012 15498 16046
rect 15390 15973 15498 16012
rect 17942 16048 17948 16082
rect 17982 16048 18060 16082
rect 17942 16014 18020 16048
rect 18054 16014 18060 16048
rect 17942 16009 18060 16014
rect 15390 15939 15396 15973
rect 15430 15939 15498 15973
rect 15390 15900 15498 15939
rect 15390 15866 15396 15900
rect 15430 15866 15498 15900
rect 15390 15827 15498 15866
rect 15390 15793 15396 15827
rect 15430 15793 15498 15827
rect 15390 15754 15498 15793
rect 15390 15720 15396 15754
rect 15430 15720 15498 15754
rect 15390 15681 15498 15720
rect 15390 15647 15396 15681
rect 15430 15647 15498 15681
rect 15390 15608 15498 15647
rect 15390 15574 15396 15608
rect 15430 15574 15498 15608
rect 15390 15535 15498 15574
rect 15390 15501 15396 15535
rect 15430 15501 15498 15535
rect 15390 15462 15498 15501
rect 15390 15428 15396 15462
rect 15430 15428 15498 15462
rect 15390 15389 15498 15428
rect 15390 15355 15396 15389
rect 15430 15355 15498 15389
rect 15390 15316 15498 15355
rect 15390 15282 15396 15316
rect 15430 15282 15498 15316
rect 15390 15243 15498 15282
rect 15390 15209 15396 15243
rect 15430 15209 15498 15243
rect 15390 15170 15498 15209
rect 15390 15136 15396 15170
rect 15430 15136 15498 15170
rect 15390 15097 15498 15136
rect 15390 15063 15396 15097
rect 15430 15063 15498 15097
rect 15390 15024 15498 15063
rect 15390 14990 15396 15024
rect 15430 14990 15498 15024
rect 15390 14951 15498 14990
rect 15390 14917 15396 14951
rect 15430 14917 15498 14951
rect 15390 14878 15498 14917
rect 15390 14844 15396 14878
rect 15430 14844 15498 14878
rect 15390 14805 15498 14844
rect 15390 14771 15396 14805
rect 15430 14771 15498 14805
rect 15390 14732 15498 14771
rect 15390 14698 15396 14732
rect 15430 14698 15498 14732
rect 15390 14658 15498 14698
rect 15390 14624 15396 14658
rect 15430 14624 15498 14658
rect 15390 14584 15498 14624
rect 15390 14550 15396 14584
rect 15430 14550 15498 14584
rect 15390 14510 15498 14550
rect 15390 14476 15396 14510
rect 15430 14476 15498 14510
rect 15390 14436 15498 14476
rect 15390 14402 15396 14436
rect 15430 14402 15498 14436
rect 15390 14362 15498 14402
rect 15390 14328 15396 14362
rect 15430 14328 15498 14362
rect 15390 14288 15498 14328
rect 15390 14254 15396 14288
rect 15430 14254 15498 14288
rect 15390 14214 15498 14254
rect 15390 14180 15396 14214
rect 15430 14180 15498 14214
rect 15390 14140 15498 14180
rect 15390 14106 15396 14140
rect 15430 14106 15498 14140
rect 15390 14066 15498 14106
rect 15390 14032 15396 14066
rect 15430 14032 15498 14066
rect 10399 14026 10442 14032
rect 674 14004 923 14026
tri 923 14004 945 14026 sw
tri 3030 14004 3052 14026 se
rect 3052 14004 3640 14026
tri 3640 14004 3662 14026 sw
tri 5536 14004 5558 14026 se
rect 5558 14004 5765 14026
tri 5765 14004 5787 14026 sw
tri 7662 14004 7684 14026 se
rect 7684 14004 8324 14026
tri 8324 14004 8346 14026 sw
tri 10220 14004 10242 14026 se
rect 10242 14004 10442 14026
tri 10442 14004 10470 14032 sw
tri 12445 14004 12473 14032 se
rect 12473 14004 15130 14032
tri 15130 14004 15158 14032 sw
tri 15388 14004 15390 14006 se
rect 15390 14004 15498 14032
rect 674 13996 945 14004
rect 674 13962 680 13996
rect 714 13962 752 13996
rect 786 13992 945 13996
tri 945 13992 957 14004 sw
tri 3018 13992 3030 14004 se
rect 3030 13992 3662 14004
tri 3662 13992 3674 14004 sw
tri 5524 13992 5536 14004 se
rect 5536 13992 5787 14004
tri 5787 13992 5799 14004 sw
tri 7650 13992 7662 14004 se
rect 7662 13992 8346 14004
tri 8346 13992 8358 14004 sw
tri 10208 13992 10220 14004 se
rect 10220 13992 10470 14004
tri 10470 13992 10482 14004 sw
tri 12433 13992 12445 14004 se
rect 12445 13992 15158 14004
tri 15158 13992 15170 14004 sw
tri 15376 13992 15388 14004 se
rect 15388 13992 15498 14004
rect 786 13991 957 13992
tri 957 13991 958 13992 sw
tri 3017 13991 3018 13992 se
rect 3018 13991 3674 13992
tri 3674 13991 3675 13992 sw
tri 5523 13991 5524 13992 se
rect 5524 13991 5799 13992
tri 5799 13991 5800 13992 sw
tri 7649 13991 7650 13992 se
rect 7650 13991 8358 13992
tri 8358 13991 8359 13992 sw
tri 10207 13991 10208 13992 se
rect 10208 13991 10482 13992
tri 10482 13991 10483 13992 sw
tri 12432 13991 12433 13992 se
rect 12433 13991 15170 13992
rect 786 13962 958 13991
rect 674 13957 958 13962
tri 958 13957 992 13991 sw
tri 2983 13957 3017 13991 se
rect 3017 13957 3267 13991
rect 3301 13957 3339 13991
rect 3373 13987 3675 13991
tri 3675 13987 3679 13991 sw
tri 5519 13987 5523 13991 se
rect 5523 13987 5800 13991
rect 3373 13957 3679 13987
rect 674 13953 992 13957
tri 992 13953 996 13957 sw
tri 2979 13953 2983 13957 se
rect 2983 13953 3679 13957
tri 3679 13953 3713 13987 sw
tri 5485 13953 5519 13987 se
rect 5519 13953 5609 13987
rect 5643 13953 5681 13987
rect 5715 13957 5800 13987
tri 5800 13957 5834 13991 sw
tri 7615 13957 7649 13991 se
rect 7649 13957 7951 13991
rect 7985 13957 8023 13991
rect 8057 13987 8359 13991
tri 8359 13987 8363 13991 sw
tri 10203 13987 10207 13991 se
rect 10207 13987 10483 13991
rect 8057 13957 8363 13987
rect 5715 13953 5834 13957
tri 5834 13953 5838 13957 sw
tri 7611 13953 7615 13957 se
rect 7615 13953 8363 13957
tri 8363 13953 8397 13987 sw
tri 10169 13953 10203 13987 se
rect 10203 13953 10293 13987
rect 10327 13953 10365 13987
rect 10399 13957 10483 13987
tri 10483 13957 10517 13991 sw
tri 12398 13957 12432 13991 se
rect 12432 13957 12682 13991
rect 12716 13957 12754 13991
rect 12788 13981 15170 13991
tri 15170 13981 15181 13992 sw
tri 15365 13981 15376 13992 se
rect 15376 13981 15396 13992
rect 12788 13958 15396 13981
rect 15430 13958 15498 13992
rect 15554 15431 17675 15983
rect 17942 15975 17948 16009
rect 17982 15975 18060 16009
rect 17942 15941 18020 15975
rect 18054 15941 18060 15975
rect 17942 15936 18060 15941
rect 17942 15902 17948 15936
rect 17982 15902 18060 15936
rect 17942 15868 18020 15902
rect 18054 15868 18060 15902
rect 17942 15863 18060 15868
rect 17942 15829 17948 15863
rect 17982 15829 18060 15863
rect 17942 15795 18020 15829
rect 18054 15795 18060 15829
rect 17942 15790 18060 15795
rect 17942 15756 17948 15790
rect 17982 15756 18060 15790
rect 17942 15722 18020 15756
rect 18054 15722 18060 15756
rect 17942 15717 18060 15722
rect 17942 15683 17948 15717
rect 17982 15683 18060 15717
rect 17942 15649 18020 15683
rect 18054 15649 18060 15683
rect 17942 15644 18060 15649
rect 17942 15610 17948 15644
rect 17982 15610 18060 15644
rect 17942 15576 18020 15610
rect 18054 15576 18060 15610
rect 17942 15571 18060 15576
rect 17942 15537 17948 15571
rect 17982 15537 18060 15571
tri 17917 15503 17942 15528 se
rect 17942 15503 18020 15537
rect 18054 15503 18060 15537
tri 17912 15498 17917 15503 se
rect 17917 15498 18060 15503
tri 17878 15464 17912 15498 se
rect 17912 15464 17948 15498
rect 17982 15464 18060 15498
tri 17845 15431 17878 15464 se
rect 17878 15431 18020 15464
rect 15554 15430 15938 15431
tri 15938 15430 15939 15431 nw
tri 17844 15430 17845 15431 se
rect 17845 15430 18020 15431
rect 18054 15430 18060 15464
rect 15554 15425 15933 15430
tri 15933 15425 15938 15430 nw
tri 17839 15425 17844 15430 se
rect 17844 15425 18060 15430
rect 15554 15391 15899 15425
tri 15899 15391 15933 15425 nw
tri 17805 15391 17839 15425 se
rect 17839 15391 17948 15425
rect 17982 15391 18060 15425
rect 15554 15357 15865 15391
tri 15865 15357 15899 15391 nw
tri 17789 15375 17805 15391 se
rect 17805 15375 18020 15391
tri 15945 15357 15963 15375 se
rect 15963 15357 18020 15375
rect 18054 15357 18060 15391
rect 15554 15352 15860 15357
tri 15860 15352 15865 15357 nw
tri 15940 15352 15945 15357 se
rect 15945 15352 18060 15357
rect 15554 15351 15859 15352
tri 15859 15351 15860 15352 nw
tri 15939 15351 15940 15352 se
rect 15940 15351 17948 15352
rect 15554 15318 15826 15351
tri 15826 15318 15859 15351 nw
tri 15906 15318 15939 15351 se
rect 15939 15318 17948 15351
rect 17982 15318 18060 15352
rect 15554 14588 15793 15318
tri 15793 15285 15826 15318 nw
tri 15873 15285 15906 15318 se
rect 15906 15285 18020 15318
tri 15872 15284 15873 15285 se
rect 15873 15284 18020 15285
rect 18054 15284 18060 15318
tri 15867 15279 15872 15284 se
rect 15872 15279 18060 15284
tri 15849 15261 15867 15279 se
rect 15867 15261 17948 15279
rect 15849 15245 17948 15261
rect 17982 15245 18060 15279
rect 15849 15211 18020 15245
rect 18054 15211 18060 15245
rect 15849 15206 18060 15211
rect 15849 15172 17948 15206
rect 17982 15172 18060 15206
rect 15849 15138 18020 15172
rect 18054 15138 18060 15172
rect 15849 15133 18060 15138
rect 15849 15099 17948 15133
rect 17982 15099 18060 15133
rect 15849 15065 18020 15099
rect 18054 15065 18060 15099
rect 15849 15060 18060 15065
rect 15849 15026 17948 15060
rect 17982 15026 18060 15060
rect 15849 14992 18020 15026
rect 18054 14992 18060 15026
rect 15849 14987 18060 14992
rect 15849 14953 17948 14987
rect 17982 14953 18060 14987
rect 15849 14919 18020 14953
rect 18054 14919 18060 14953
rect 15849 14914 18060 14919
rect 15849 14880 17948 14914
rect 17982 14880 18060 14914
rect 15849 14846 18020 14880
rect 18054 14846 18060 14880
rect 15849 14841 18060 14846
rect 15849 14807 17948 14841
rect 17982 14807 18060 14841
rect 15849 14773 18020 14807
rect 18054 14773 18060 14807
rect 15849 14768 18060 14773
rect 15849 14734 17948 14768
rect 17982 14734 18060 14768
rect 15849 14700 18020 14734
rect 18054 14700 18060 14734
rect 15849 14695 18060 14700
rect 15849 14661 17948 14695
rect 17982 14661 18060 14695
rect 15849 14644 18020 14661
tri 17561 14627 17578 14644 ne
rect 17578 14627 18020 14644
rect 18054 14627 18060 14661
tri 17578 14622 17583 14627 ne
rect 17583 14622 18060 14627
tri 17583 14596 17609 14622 ne
rect 17609 14596 17948 14622
tri 15793 14588 15801 14596 sw
tri 17609 14588 17617 14596 ne
rect 17617 14588 17948 14596
rect 17982 14588 18060 14622
rect 15554 14554 15801 14588
tri 15801 14554 15835 14588 sw
tri 17617 14554 17651 14588 ne
rect 17651 14554 18020 14588
rect 18054 14554 18060 14588
rect 15554 14549 15835 14554
tri 15835 14549 15840 14554 sw
tri 17651 14549 17656 14554 ne
rect 17656 14549 18060 14554
rect 15554 14515 15840 14549
tri 15840 14515 15874 14549 sw
tri 17656 14515 17690 14549 ne
rect 17690 14515 17948 14549
rect 17982 14515 18060 14549
rect 15554 14481 15874 14515
tri 15874 14481 15908 14515 sw
tri 17690 14481 17724 14515 ne
rect 17724 14481 18020 14515
rect 18054 14481 18060 14515
rect 15554 14476 15908 14481
tri 15908 14476 15913 14481 sw
tri 17724 14476 17729 14481 ne
rect 17729 14476 18060 14481
rect 15554 14450 15913 14476
tri 15913 14450 15939 14476 sw
tri 17729 14474 17731 14476 ne
rect 15554 14442 17628 14450
tri 17628 14442 17636 14450 sw
rect 17731 14442 17948 14476
rect 17982 14442 18060 14476
rect 15554 14408 17636 14442
tri 17636 14408 17670 14442 sw
rect 17731 14408 18020 14442
rect 18054 14408 18060 14442
rect 15554 14403 17670 14408
tri 17670 14403 17675 14408 sw
rect 15554 13976 17675 14403
tri 15554 13970 15560 13976 ne
rect 15560 13970 17675 13976
tri 15560 13965 15565 13970 ne
rect 15565 13965 17675 13970
rect 12788 13957 15498 13958
rect 10399 13953 10517 13957
rect 674 13939 996 13953
tri 996 13939 1010 13953 sw
tri 2965 13939 2979 13953 se
rect 2979 13939 3713 13953
tri 3713 13939 3727 13953 sw
tri 5471 13939 5485 13953 se
rect 5485 13939 5838 13953
tri 5838 13939 5852 13953 sw
tri 7597 13939 7611 13953 se
rect 7611 13939 8397 13953
tri 8397 13939 8411 13953 sw
tri 10155 13939 10169 13953 se
rect 10169 13939 10517 13953
tri 10517 13939 10535 13957 sw
tri 12380 13939 12398 13957 se
rect 12398 13939 15498 13957
tri 15565 13952 15578 13965 ne
rect 15578 13952 17675 13965
rect 674 13931 15498 13939
tri 15498 13931 15519 13952 sw
tri 15578 13931 15599 13952 ne
rect 15599 13945 17675 13952
rect 15599 13931 17661 13945
tri 17661 13931 17675 13945 nw
rect 17731 14403 18060 14408
rect 17731 14369 17948 14403
rect 17982 14369 18060 14403
rect 17731 14335 18020 14369
rect 18054 14335 18060 14369
rect 17731 14330 18060 14335
rect 17731 14296 17948 14330
rect 17982 14296 18060 14330
rect 17731 14262 18020 14296
rect 18054 14262 18060 14296
rect 17731 14257 18060 14262
rect 17731 14223 17948 14257
rect 17982 14223 18060 14257
rect 17731 14189 18020 14223
rect 18054 14189 18060 14223
rect 17731 14184 18060 14189
rect 17731 14150 17948 14184
rect 17982 14150 18060 14184
rect 17731 14116 18020 14150
rect 18054 14116 18060 14150
rect 17731 14111 18060 14116
rect 17731 14077 17948 14111
rect 17982 14077 18060 14111
rect 17731 14043 18020 14077
rect 18054 14043 18060 14077
rect 17731 14038 18060 14043
rect 17731 14004 17948 14038
rect 17982 14004 18060 14038
rect 17731 13970 18020 14004
rect 18054 13970 18060 14004
rect 17731 13965 18060 13970
rect 17731 13931 17948 13965
rect 17982 13931 18060 13965
rect 674 13921 15519 13931
rect 674 13887 680 13921
rect 714 13887 752 13921
rect 786 13918 15519 13921
rect 786 13914 15396 13918
rect 786 13887 3267 13914
rect 674 13880 3267 13887
rect 3301 13880 3339 13914
rect 3373 13880 5609 13914
rect 5643 13880 5681 13914
rect 5715 13880 7951 13914
rect 7985 13880 8023 13914
rect 8057 13880 10293 13914
rect 10327 13880 10365 13914
rect 10399 13880 12682 13914
rect 12716 13880 12754 13914
rect 12788 13884 15396 13914
rect 15430 13898 15519 13918
tri 15519 13898 15552 13931 sw
tri 15599 13898 15632 13931 ne
rect 15632 13898 17628 13931
tri 17628 13898 17661 13931 nw
rect 15430 13897 15552 13898
tri 15552 13897 15553 13898 sw
rect 17731 13897 18020 13931
rect 18054 13897 18060 13931
rect 15430 13892 15553 13897
tri 15553 13892 15558 13897 sw
rect 17731 13892 18060 13897
rect 15430 13884 15558 13892
rect 12788 13880 15558 13884
rect 674 13858 15558 13880
tri 15558 13858 15592 13892 sw
tri 17714 13858 17731 13875 se
rect 17731 13858 17948 13892
rect 17982 13858 18060 13892
rect 674 13846 15592 13858
rect 674 13812 680 13846
rect 714 13812 752 13846
rect 786 13844 15592 13846
rect 786 13812 15396 13844
rect 674 13810 15396 13812
rect 15430 13824 15592 13844
tri 15592 13824 15626 13858 sw
tri 17680 13824 17714 13858 se
rect 17714 13824 18020 13858
rect 18054 13824 18060 13858
rect 15430 13819 15626 13824
tri 15626 13819 15631 13824 sw
tri 17675 13819 17680 13824 se
rect 17680 13819 18060 13824
rect 15430 13810 15631 13819
rect 674 13785 15631 13810
tri 15631 13785 15665 13819 sw
tri 17641 13785 17675 13819 se
rect 17675 13785 17948 13819
rect 17982 13785 18060 13819
rect 674 13771 15665 13785
rect 674 13737 680 13771
rect 714 13737 752 13771
rect 786 13770 15665 13771
rect 786 13737 15396 13770
rect 674 13736 15396 13737
rect 15430 13751 15665 13770
tri 15665 13751 15699 13785 sw
tri 17607 13751 17641 13785 se
rect 17641 13751 18020 13785
rect 18054 13751 18060 13785
rect 15430 13746 15699 13751
tri 15699 13746 15704 13751 sw
tri 17602 13746 17607 13751 se
rect 17607 13746 18060 13751
rect 15430 13736 15704 13746
rect 674 13733 15704 13736
tri 15704 13733 15717 13746 sw
tri 17589 13733 17602 13746 se
rect 17602 13733 17948 13746
rect 674 13712 17948 13733
rect 17982 13712 18060 13746
rect 674 13696 18020 13712
rect 674 13662 680 13696
rect 714 13662 752 13696
rect 786 13662 15396 13696
rect 15430 13678 18020 13696
rect 18054 13678 18060 13712
rect 15430 13673 18060 13678
rect 15430 13662 17948 13673
rect 674 13639 17948 13662
rect 17982 13639 18060 13673
rect 674 13622 18020 13639
rect 674 13621 15396 13622
rect 674 13587 680 13621
rect 714 13587 752 13621
rect 786 13588 15396 13621
rect 15430 13605 18020 13622
rect 18054 13605 18060 13639
rect 15430 13600 18060 13605
rect 15430 13588 17948 13600
rect 786 13587 17948 13588
rect 674 13566 17948 13587
rect 17982 13566 18060 13600
rect 674 13548 18020 13566
rect 674 13547 15396 13548
rect 674 13513 680 13547
rect 714 13513 752 13547
rect 786 13514 15396 13547
rect 15430 13532 18020 13548
rect 18054 13532 18060 13566
rect 15430 13527 18060 13532
rect 15430 13514 17948 13527
rect 786 13513 17948 13514
rect 674 13493 17948 13513
rect 17982 13493 18060 13527
rect 674 13474 18020 13493
rect 674 13473 15396 13474
rect 674 13439 680 13473
rect 714 13439 752 13473
rect 786 13440 15396 13473
rect 15430 13459 18020 13474
rect 18054 13459 18060 13493
rect 15430 13454 18060 13459
rect 15430 13440 17948 13454
rect 786 13439 17948 13440
rect 674 13420 17948 13439
rect 17982 13420 18060 13454
rect 674 13400 18020 13420
rect 674 13399 15396 13400
rect 674 13365 680 13399
rect 714 13365 752 13399
rect 786 13366 15396 13399
rect 15430 13386 18020 13400
rect 18054 13386 18060 13420
rect 15430 13381 18060 13386
rect 15430 13366 17948 13381
rect 786 13365 17948 13366
rect 674 13347 17948 13365
rect 17982 13347 18060 13381
rect 674 13326 18020 13347
rect 674 13325 15396 13326
rect 674 13291 680 13325
rect 714 13291 752 13325
rect 786 13292 15396 13325
rect 15430 13313 18020 13326
rect 18054 13313 18060 13347
rect 15430 13308 18060 13313
rect 15430 13292 17948 13308
rect 786 13291 17948 13292
rect 674 13274 17948 13291
rect 17982 13274 18060 13308
rect 674 13252 18020 13274
rect 674 13251 15396 13252
rect 674 13217 680 13251
rect 714 13217 752 13251
rect 786 13218 15396 13251
rect 15430 13240 18020 13252
rect 18054 13240 18060 13274
rect 15430 13235 18060 13240
rect 15430 13218 17948 13235
rect 786 13217 17948 13218
rect 674 13206 17948 13217
rect 674 13201 14728 13206
tri 14728 13201 14733 13206 nw
tri 15574 13201 15579 13206 ne
rect 15579 13201 17948 13206
rect 17982 13201 18060 13235
rect 674 13177 14694 13201
rect 674 13143 680 13177
rect 714 13143 752 13177
rect 786 13167 14694 13177
tri 14694 13167 14728 13201 nw
tri 15579 13167 15613 13201 ne
rect 15613 13167 18020 13201
rect 18054 13167 18060 13201
rect 786 13162 14689 13167
tri 14689 13162 14694 13167 nw
tri 15613 13162 15618 13167 ne
rect 15618 13162 18060 13167
rect 786 13143 14665 13162
rect 674 13138 14665 13143
tri 14665 13138 14689 13162 nw
tri 15618 13150 15630 13162 ne
rect 15630 13150 17948 13162
rect 14817 13138 14935 13150
rect 674 13104 14631 13138
tri 14631 13104 14665 13138 nw
rect 14817 13104 14823 13138
rect 14857 13104 14895 13138
rect 14929 13104 14935 13138
rect 674 13103 14621 13104
rect 674 13069 680 13103
rect 714 13069 752 13103
rect 786 13094 14621 13103
tri 14621 13094 14631 13104 nw
rect 786 13089 14616 13094
tri 14616 13089 14621 13094 nw
rect 786 13069 14586 13089
rect 674 13029 14586 13069
tri 14586 13059 14616 13089 nw
rect 674 12995 680 13029
rect 714 12995 752 13029
rect 786 12995 14586 13029
rect 674 12955 14586 12995
rect 674 12921 680 12955
rect 714 12921 752 12955
rect 786 12943 14586 12955
rect 786 12921 829 12943
rect 674 12881 829 12921
rect 674 12847 680 12881
rect 714 12847 752 12881
rect 786 12847 829 12881
rect 674 12837 829 12847
rect 12311 12909 12350 12943
rect 12384 12909 12423 12943
rect 12457 12909 12496 12943
rect 12530 12909 12569 12943
rect 12603 12909 12642 12943
rect 12676 12909 12715 12943
rect 12749 12909 12788 12943
rect 12822 12909 12861 12943
rect 12895 12909 12934 12943
rect 12968 12909 13007 12943
rect 13041 12909 13080 12943
rect 13114 12909 13153 12943
rect 13187 12909 13226 12943
rect 13260 12909 13299 12943
rect 13333 12909 13372 12943
rect 13406 12909 13445 12943
rect 13479 12909 13518 12943
rect 13552 12909 13591 12943
rect 13625 12909 13664 12943
rect 13698 12909 13737 12943
rect 13771 12909 13810 12943
rect 13844 12909 13883 12943
rect 13917 12909 13956 12943
rect 13990 12909 14029 12943
rect 14063 12909 14102 12943
rect 14136 12909 14175 12943
rect 14209 12909 14248 12943
rect 14282 12909 14321 12943
rect 14355 12909 14394 12943
rect 14428 12909 14467 12943
rect 14501 12909 14540 12943
rect 14574 12909 14586 12943
rect 12311 12871 14586 12909
rect 12311 12837 12350 12871
rect 12384 12837 12423 12871
rect 12457 12837 12496 12871
rect 12530 12837 12569 12871
rect 12603 12837 12642 12871
rect 12676 12837 12715 12871
rect 12749 12837 12788 12871
rect 12822 12837 12861 12871
rect 12895 12837 12934 12871
rect 12968 12837 13007 12871
rect 13041 12837 13080 12871
rect 13114 12837 13153 12871
rect 13187 12837 13226 12871
rect 13260 12837 13299 12871
rect 13333 12837 13372 12871
rect 13406 12837 13445 12871
rect 13479 12837 13518 12871
rect 13552 12837 13591 12871
rect 13625 12837 13664 12871
rect 13698 12837 13737 12871
rect 13771 12837 13810 12871
rect 13844 12837 13883 12871
rect 13917 12837 13956 12871
rect 13990 12837 14029 12871
rect 14063 12837 14102 12871
rect 14136 12837 14175 12871
rect 14209 12837 14248 12871
rect 14282 12837 14321 12871
rect 14355 12837 14394 12871
rect 14428 12837 14467 12871
rect 14501 12837 14540 12871
rect 14574 12837 14586 12871
rect 674 12737 14586 12837
rect 674 12732 10769 12737
tri 10769 12732 10774 12737 nw
rect 674 12717 10735 12732
rect 674 12698 2490 12717
tri 2490 12698 2509 12717 nw
tri 4318 12698 4337 12717 ne
rect 4337 12698 6613 12717
tri 6613 12698 6632 12717 nw
tri 8441 12698 8460 12717 ne
rect 8460 12698 10735 12717
tri 10735 12698 10769 12732 nw
rect 674 12693 2485 12698
tri 2485 12693 2490 12698 nw
tri 4337 12693 4342 12698 ne
rect 4342 12693 6608 12698
tri 6608 12693 6613 12698 nw
tri 8460 12693 8465 12698 ne
rect 8465 12693 10730 12698
tri 10730 12693 10735 12698 nw
rect 674 12659 2451 12693
tri 2451 12659 2485 12693 nw
tri 4342 12659 4376 12693 ne
rect 4376 12659 6574 12693
tri 6574 12659 6608 12693 nw
tri 8465 12659 8499 12693 ne
rect 8499 12659 10696 12693
tri 10696 12659 10730 12693 nw
rect 674 12625 2417 12659
tri 2417 12625 2451 12659 nw
tri 4376 12629 4406 12659 ne
rect 4406 12629 6540 12659
rect 674 12623 2415 12625
tri 2415 12623 2417 12625 nw
rect 2517 12623 4252 12629
tri 4406 12625 4410 12629 ne
rect 4410 12625 6540 12629
tri 6540 12625 6574 12659 nw
tri 8499 12629 8529 12659 ne
rect 8529 12629 10662 12659
tri 4410 12623 4412 12625 ne
rect 4412 12623 6538 12625
tri 6538 12623 6540 12625 nw
rect 6646 12623 8382 12629
tri 8529 12625 8533 12629 ne
rect 8533 12625 10662 12629
tri 10662 12625 10696 12659 nw
tri 8533 12623 8535 12625 ne
rect 8535 12623 10660 12625
tri 10660 12623 10662 12625 nw
rect 10778 12623 14710 12629
rect 674 12589 2381 12623
tri 2381 12589 2415 12623 nw
rect 2517 12589 2529 12623
rect 2563 12589 2602 12623
rect 2636 12589 2675 12623
rect 2709 12589 2748 12623
rect 2782 12589 2821 12623
rect 2855 12589 2894 12623
rect 2928 12589 2967 12623
rect 3001 12589 3040 12623
rect 3074 12589 3113 12623
rect 3147 12589 3186 12623
rect 3220 12589 3259 12623
rect 3293 12589 3332 12623
rect 3366 12589 3405 12623
rect 3439 12589 3478 12623
rect 3512 12589 3551 12623
rect 3585 12589 3624 12623
rect 3658 12589 3697 12623
rect 3731 12589 3770 12623
rect 674 12582 2344 12589
rect 674 12551 1221 12582
tri 1221 12551 1252 12582 nw
tri 1453 12551 1484 12582 ne
rect 1484 12551 2344 12582
tri 2344 12552 2381 12589 nw
rect 351 12502 357 12536
rect 391 12502 429 12536
rect 463 12502 469 12536
tri 651 12517 674 12540 se
rect 674 12517 1187 12551
tri 1187 12517 1221 12551 nw
tri 1484 12517 1518 12551 ne
rect 1518 12517 2344 12551
tri 648 12514 651 12517 se
rect 651 12514 1184 12517
tri 1184 12514 1187 12517 nw
tri 1518 12514 1521 12517 ne
rect 1521 12514 2344 12517
rect 351 12490 469 12502
tri 624 12490 648 12514 se
rect 648 12490 1107 12514
tri 556 12422 624 12490 se
rect 624 12422 1107 12490
tri 1107 12437 1184 12514 nw
tri 1521 12437 1598 12514 ne
rect 360 12257 1107 12422
rect 1598 12285 2344 12514
rect 2517 12551 3770 12589
rect 2517 12517 2529 12551
rect 2563 12517 2602 12551
rect 2636 12517 2675 12551
rect 2709 12517 2748 12551
rect 2782 12517 2821 12551
rect 2855 12517 2894 12551
rect 2928 12517 2967 12551
rect 3001 12517 3040 12551
rect 3074 12517 3113 12551
rect 3147 12517 3186 12551
rect 3220 12517 3259 12551
rect 3293 12517 3332 12551
rect 3366 12517 3405 12551
rect 3439 12517 3478 12551
rect 3512 12517 3551 12551
rect 3585 12517 3624 12551
rect 3658 12517 3697 12551
rect 3731 12517 3770 12551
rect 4236 12517 4252 12623
tri 4412 12589 4446 12623 ne
rect 4446 12589 6504 12623
tri 6504 12589 6538 12623 nw
rect 6646 12589 6663 12623
rect 6697 12589 6736 12623
rect 6770 12589 6809 12623
rect 6843 12589 6882 12623
rect 6916 12589 6955 12623
rect 6989 12589 7028 12623
rect 7062 12589 7101 12623
rect 7135 12589 7174 12623
rect 7208 12589 7247 12623
rect 7281 12589 7320 12623
rect 7354 12589 7393 12623
rect 7427 12589 7466 12623
rect 7500 12589 7539 12623
rect 7573 12589 7612 12623
rect 7646 12589 7685 12623
rect 7719 12589 7758 12623
rect 7792 12589 7831 12623
rect 7865 12589 7904 12623
tri 4446 12552 4483 12589 ne
rect 4483 12582 6467 12589
rect 2517 12257 4252 12517
rect 4483 12551 5343 12582
tri 5343 12551 5374 12582 nw
tri 5576 12551 5607 12582 ne
rect 5607 12551 6467 12582
tri 6467 12552 6504 12589 nw
rect 4483 12517 5309 12551
tri 5309 12517 5343 12551 nw
tri 5607 12517 5641 12551 ne
rect 5641 12517 6467 12551
rect 4483 12514 5306 12517
tri 5306 12514 5309 12517 nw
tri 5641 12514 5644 12517 ne
rect 5644 12514 6467 12517
rect 4483 12285 5229 12514
tri 5229 12437 5306 12514 nw
tri 5644 12437 5721 12514 ne
rect 5721 12285 6467 12514
rect 6646 12551 7904 12589
rect 6646 12517 6663 12551
rect 6697 12517 6736 12551
rect 6770 12517 6809 12551
rect 6843 12517 6882 12551
rect 6916 12517 6955 12551
rect 6989 12517 7028 12551
rect 7062 12517 7101 12551
rect 7135 12517 7174 12551
rect 7208 12517 7247 12551
rect 7281 12517 7320 12551
rect 7354 12517 7393 12551
rect 7427 12517 7466 12551
rect 7500 12517 7539 12551
rect 7573 12517 7612 12551
rect 7646 12517 7685 12551
rect 7719 12517 7758 12551
rect 7792 12517 7831 12551
rect 7865 12517 7904 12551
rect 8370 12517 8382 12623
tri 8535 12589 8569 12623 ne
rect 8569 12589 10626 12623
tri 10626 12589 10660 12623 nw
rect 10778 12589 10790 12623
rect 10824 12589 10864 12623
rect 10898 12589 10938 12623
rect 10972 12589 11012 12623
rect 11046 12589 11086 12623
rect 11120 12589 11160 12623
rect 11194 12589 11233 12623
rect 11267 12589 11306 12623
rect 11340 12589 11379 12623
rect 11413 12589 11452 12623
rect 11486 12589 11525 12623
rect 11559 12589 11598 12623
rect 11632 12589 11671 12623
rect 11705 12589 11744 12623
rect 11778 12589 11817 12623
rect 11851 12589 11890 12623
rect 11924 12589 11963 12623
rect 11997 12589 12036 12623
rect 12070 12589 12109 12623
rect 12143 12589 12182 12623
rect 12216 12589 12255 12623
rect 12289 12589 12328 12623
rect 12362 12589 12401 12623
rect 12435 12589 12474 12623
rect 12508 12589 12547 12623
rect 12581 12589 12620 12623
rect 12654 12589 12693 12623
rect 12727 12589 12766 12623
rect 12800 12589 12839 12623
rect 12873 12589 12912 12623
rect 12946 12589 12985 12623
rect 13019 12589 13058 12623
rect 13092 12589 13131 12623
rect 13165 12589 13204 12623
rect 13238 12589 13277 12623
rect 13311 12589 13350 12623
rect 13384 12589 13423 12623
rect 13457 12589 13496 12623
rect 13530 12589 13569 12623
rect 13603 12589 13642 12623
rect 13676 12589 13715 12623
rect 13749 12589 13788 12623
rect 13822 12589 13861 12623
rect 13895 12589 13934 12623
rect 13968 12589 14007 12623
rect 14041 12589 14080 12623
rect 14114 12589 14153 12623
rect 14187 12589 14226 12623
rect 14260 12589 14299 12623
rect 14333 12589 14372 12623
rect 14406 12589 14445 12623
rect 14479 12589 14518 12623
rect 14552 12589 14591 12623
rect 14625 12589 14664 12623
rect 14698 12589 14710 12623
tri 8569 12586 8572 12589 ne
rect 8572 12586 10623 12589
tri 10623 12586 10626 12589 nw
tri 8572 12553 8605 12586 ne
rect 8605 12582 10589 12586
rect 6646 12257 8382 12517
rect 8605 12552 9467 12582
tri 9467 12552 9497 12582 nw
tri 9698 12552 9728 12582 ne
rect 9728 12552 10589 12582
tri 10589 12552 10623 12586 nw
rect 8605 12551 9466 12552
tri 9466 12551 9467 12552 nw
tri 9728 12551 9729 12552 ne
rect 9729 12551 10589 12552
rect 8605 12517 9432 12551
tri 9432 12517 9466 12551 nw
tri 9729 12517 9763 12551 ne
rect 9763 12517 10589 12551
rect 8605 12514 9429 12517
tri 9429 12514 9432 12517 nw
tri 9763 12514 9766 12517 ne
rect 9766 12514 10589 12517
rect 8605 12285 9352 12514
tri 9352 12437 9429 12514 nw
tri 9766 12437 9843 12514 ne
rect 9843 12285 10589 12514
rect 10778 12551 14710 12589
rect 10778 12517 10790 12551
rect 10824 12517 10864 12551
rect 10898 12517 10938 12551
rect 10972 12517 11012 12551
rect 11046 12517 11086 12551
rect 11120 12517 11160 12551
rect 11194 12517 11233 12551
rect 11267 12517 11306 12551
rect 11340 12517 11379 12551
rect 11413 12517 11452 12551
rect 11486 12517 11525 12551
rect 11559 12517 11598 12551
rect 11632 12517 11671 12551
rect 11705 12517 11744 12551
rect 11778 12517 11817 12551
rect 11851 12517 11890 12551
rect 11924 12517 11963 12551
rect 11997 12517 12036 12551
rect 12070 12517 12109 12551
rect 12143 12517 12182 12551
rect 12216 12517 12255 12551
rect 12289 12517 12328 12551
rect 12362 12517 12401 12551
rect 12435 12517 12474 12551
rect 12508 12517 12547 12551
rect 12581 12517 12620 12551
rect 12654 12517 12693 12551
rect 12727 12517 12766 12551
rect 12800 12517 12839 12551
rect 12873 12517 12912 12551
rect 12946 12517 12985 12551
rect 13019 12517 13058 12551
rect 13092 12517 13131 12551
rect 13165 12517 13204 12551
rect 13238 12517 13277 12551
rect 13311 12517 13350 12551
rect 13384 12517 13423 12551
rect 13457 12517 13496 12551
rect 13530 12517 13569 12551
rect 13603 12517 13642 12551
rect 13676 12517 13715 12551
rect 13749 12517 13788 12551
rect 13822 12517 13861 12551
rect 13895 12517 13934 12551
rect 13968 12517 14007 12551
rect 14041 12517 14080 12551
rect 14114 12517 14153 12551
rect 14187 12517 14226 12551
rect 14260 12517 14299 12551
rect 14333 12517 14372 12551
rect 14406 12517 14445 12551
rect 14479 12517 14518 12551
rect 14552 12517 14591 12551
rect 14625 12517 14664 12551
rect 14698 12517 14710 12551
rect 10778 12511 14710 12517
rect 10778 12257 11739 12511
tri 11739 12486 11764 12511 nw
rect 14817 12329 14935 13104
rect 14963 13138 15079 13150
rect 15081 13149 15117 13150
rect 14963 13104 14969 13138
rect 15003 13104 15041 13138
rect 15075 13104 15079 13138
rect 14963 13092 15079 13104
rect 15080 13093 15118 13149
rect 15119 13138 15235 13150
rect 15119 13104 15123 13138
rect 15157 13104 15195 13138
rect 15229 13104 15235 13138
tri 15630 13128 15652 13150 ne
rect 15652 13128 17948 13150
rect 17982 13128 18060 13162
rect 15081 13092 15117 13093
rect 15119 13092 15235 13104
tri 15652 13094 15686 13128 ne
rect 15686 13094 18020 13128
rect 18054 13094 18060 13128
tri 15686 13092 15688 13094 ne
rect 15688 13092 18060 13094
rect 14963 13089 15076 13092
tri 15076 13089 15079 13092 nw
tri 15688 13089 15691 13092 ne
rect 15691 13089 18060 13092
rect 14963 13014 15054 13089
tri 15054 13067 15076 13089 nw
tri 15691 13067 15713 13089 ne
rect 15713 13067 17948 13089
tri 15713 13055 15725 13067 ne
rect 15725 13055 17948 13067
rect 17982 13055 18060 13089
tri 15223 13043 15235 13055 se
rect 15235 13043 15353 13055
tri 15219 13039 15223 13043 se
rect 15223 13039 15241 13043
tri 15054 13014 15079 13039 sw
tri 15194 13014 15219 13039 se
rect 15219 13014 15241 13039
rect 14963 12956 15079 13014
rect 15080 12957 15081 13013
rect 15117 12957 15118 13013
rect 15119 13009 15241 13014
rect 15275 13009 15313 13043
rect 15347 13009 15353 13043
rect 15119 12956 15353 13009
tri 15210 12948 15218 12956 ne
rect 15218 12948 15353 12956
tri 15218 12943 15223 12948 ne
rect 15223 12943 15353 12948
tri 15223 12931 15235 12943 ne
rect 15235 12329 15353 12943
rect 15381 13043 15499 13055
rect 15381 13009 15387 13043
rect 15421 13009 15459 13043
rect 15493 13009 15499 13043
rect 15381 12329 15499 13009
rect 15527 13043 15645 13055
tri 15725 13044 15736 13055 ne
rect 15527 13009 15533 13043
rect 15567 13009 15605 13043
rect 15639 13009 15645 13043
rect 15527 12329 15645 13009
rect 15736 13021 18020 13055
rect 18054 13021 18060 13055
rect 15736 13016 18060 13021
rect 15736 12982 17948 13016
rect 17982 12982 18060 13016
rect 15736 12948 18020 12982
rect 18054 12948 18060 12982
rect 15736 12943 18060 12948
rect 15736 12909 15752 12943
rect 15786 12909 15826 12943
rect 15860 12909 15900 12943
rect 15934 12909 15974 12943
rect 16008 12909 16048 12943
rect 16082 12909 16122 12943
rect 16156 12909 16196 12943
rect 16230 12909 16269 12943
rect 16303 12909 16342 12943
rect 16376 12909 16415 12943
rect 16449 12909 16488 12943
rect 16522 12909 16561 12943
rect 16595 12909 16634 12943
rect 16668 12909 16707 12943
rect 16741 12909 16780 12943
rect 16814 12909 16853 12943
rect 16887 12909 16926 12943
rect 16960 12909 16999 12943
rect 17033 12909 17072 12943
rect 17106 12909 17145 12943
rect 17179 12909 17218 12943
rect 17252 12909 17291 12943
rect 17325 12909 17364 12943
rect 17398 12909 17437 12943
rect 17471 12909 17510 12943
rect 17544 12909 17583 12943
rect 17617 12909 17656 12943
rect 17690 12909 17729 12943
rect 17763 12909 17802 12943
rect 17836 12909 17875 12943
rect 17909 12909 17948 12943
rect 17982 12909 18060 12943
rect 15736 12875 18020 12909
rect 18054 12875 18060 12909
rect 15736 12871 18060 12875
rect 15736 12837 15752 12871
rect 15786 12837 15827 12871
rect 15861 12837 15902 12871
rect 15936 12837 15977 12871
rect 16011 12837 16052 12871
rect 16086 12837 16127 12871
rect 16161 12837 16202 12871
rect 16236 12837 16277 12871
rect 16311 12837 16352 12871
rect 16386 12837 16426 12871
rect 16460 12837 16500 12871
rect 16534 12837 16574 12871
rect 16608 12837 16648 12871
rect 16682 12837 16722 12871
rect 16756 12837 16796 12871
rect 16830 12837 16870 12871
rect 16904 12837 16944 12871
rect 16978 12837 17018 12871
rect 17052 12837 17092 12871
rect 17126 12837 17166 12871
rect 17200 12837 17240 12871
rect 17274 12837 17314 12871
rect 17348 12837 17388 12871
rect 17422 12837 17462 12871
rect 17496 12837 17536 12871
rect 17570 12837 17610 12871
rect 17644 12837 17684 12871
rect 17718 12837 17758 12871
rect 17792 12837 17832 12871
rect 17866 12837 17906 12871
rect 17940 12837 18060 12871
rect 15736 12831 18060 12837
rect 18265 16455 18271 17313
rect 18377 16455 18383 17315
rect 18265 16451 18383 16455
rect 18265 16417 18343 16451
rect 18377 16417 18383 16451
rect 18265 16416 18383 16417
rect 18265 16382 18271 16416
rect 18305 16382 18383 16416
rect 18265 16379 18383 16382
rect 18265 16345 18343 16379
rect 18377 16345 18383 16379
rect 18265 16343 18383 16345
rect 18265 16309 18271 16343
rect 18305 16309 18383 16343
rect 18265 16307 18383 16309
rect 18265 16273 18343 16307
rect 18377 16273 18383 16307
rect 18265 16270 18383 16273
rect 18265 16236 18271 16270
rect 18305 16236 18383 16270
rect 18265 16235 18383 16236
rect 18265 16201 18343 16235
rect 18377 16201 18383 16235
rect 18265 16197 18383 16201
rect 18265 16163 18271 16197
rect 18305 16163 18383 16197
rect 18265 16129 18343 16163
rect 18377 16129 18383 16163
rect 18265 16124 18383 16129
rect 18265 16090 18271 16124
rect 18305 16090 18383 16124
rect 18265 16056 18343 16090
rect 18377 16056 18383 16090
rect 18265 16051 18383 16056
rect 18265 16017 18271 16051
rect 18305 16017 18383 16051
rect 18265 15983 18343 16017
rect 18377 15983 18383 16017
rect 18265 15978 18383 15983
rect 18265 15944 18271 15978
rect 18305 15944 18383 15978
rect 18265 15910 18343 15944
rect 18377 15910 18383 15944
rect 18265 15905 18383 15910
rect 18265 15871 18271 15905
rect 18305 15871 18383 15905
rect 18265 15837 18343 15871
rect 18377 15837 18383 15871
rect 18265 15832 18383 15837
rect 18265 15798 18271 15832
rect 18305 15798 18383 15832
rect 18265 15764 18343 15798
rect 18377 15764 18383 15798
rect 18265 15759 18383 15764
rect 18265 15725 18271 15759
rect 18305 15725 18383 15759
rect 18265 15691 18343 15725
rect 18377 15691 18383 15725
rect 18265 15686 18383 15691
rect 18265 15652 18271 15686
rect 18305 15652 18383 15686
rect 18265 15618 18343 15652
rect 18377 15618 18383 15652
rect 18265 15613 18383 15618
rect 18265 15579 18271 15613
rect 18305 15579 18383 15613
rect 18265 15545 18343 15579
rect 18377 15545 18383 15579
rect 18265 15540 18383 15545
rect 18265 15506 18271 15540
rect 18305 15506 18383 15540
rect 18265 15472 18343 15506
rect 18377 15472 18383 15506
rect 18265 15467 18383 15472
rect 18265 15433 18271 15467
rect 18305 15433 18383 15467
rect 18265 15399 18343 15433
rect 18377 15399 18383 15433
rect 18265 15394 18383 15399
rect 18265 15360 18271 15394
rect 18305 15360 18383 15394
rect 18265 15326 18343 15360
rect 18377 15326 18383 15360
rect 18265 15321 18383 15326
rect 18265 15287 18271 15321
rect 18305 15287 18383 15321
rect 18265 15253 18343 15287
rect 18377 15253 18383 15287
rect 18265 15248 18383 15253
rect 18265 15214 18271 15248
rect 18305 15214 18383 15248
rect 18265 15180 18343 15214
rect 18377 15180 18383 15214
rect 18265 15175 18383 15180
rect 18265 15141 18271 15175
rect 18305 15141 18383 15175
rect 18265 15107 18343 15141
rect 18377 15107 18383 15141
rect 18265 15102 18383 15107
rect 18265 15068 18271 15102
rect 18305 15068 18383 15102
rect 18265 15034 18343 15068
rect 18377 15034 18383 15068
rect 18265 15029 18383 15034
rect 18265 14995 18271 15029
rect 18305 14995 18383 15029
rect 18265 14961 18343 14995
rect 18377 14961 18383 14995
rect 18265 14956 18383 14961
rect 18265 14922 18271 14956
rect 18305 14922 18383 14956
rect 18265 14888 18343 14922
rect 18377 14888 18383 14922
rect 18265 14883 18383 14888
rect 18265 14849 18271 14883
rect 18305 14849 18383 14883
rect 18265 14815 18343 14849
rect 18377 14815 18383 14849
rect 18265 14810 18383 14815
rect 18265 14776 18271 14810
rect 18305 14776 18383 14810
rect 18265 14742 18343 14776
rect 18377 14742 18383 14776
rect 18265 14737 18383 14742
rect 18265 14703 18271 14737
rect 18305 14703 18383 14737
rect 18265 14669 18343 14703
rect 18377 14669 18383 14703
rect 18265 14664 18383 14669
rect 18265 14630 18271 14664
rect 18305 14630 18383 14664
rect 18265 14596 18343 14630
rect 18377 14596 18383 14630
rect 18265 14591 18383 14596
rect 18265 14557 18271 14591
rect 18305 14557 18383 14591
rect 18265 14523 18343 14557
rect 18377 14523 18383 14557
rect 18265 14518 18383 14523
rect 18265 14484 18271 14518
rect 18305 14484 18383 14518
rect 18265 14450 18343 14484
rect 18377 14450 18383 14484
rect 18265 14445 18383 14450
rect 18265 14411 18271 14445
rect 18305 14411 18383 14445
rect 18265 14377 18343 14411
rect 18377 14377 18383 14411
rect 18265 14372 18383 14377
rect 18265 14338 18271 14372
rect 18305 14338 18383 14372
rect 18265 14304 18343 14338
rect 18377 14304 18383 14338
rect 18265 14299 18383 14304
rect 18265 14265 18271 14299
rect 18305 14265 18383 14299
rect 18265 14231 18343 14265
rect 18377 14231 18383 14265
rect 18265 14226 18383 14231
rect 18265 14192 18271 14226
rect 18305 14192 18383 14226
rect 18265 14158 18343 14192
rect 18377 14158 18383 14192
rect 18265 14153 18383 14158
rect 18265 14119 18271 14153
rect 18305 14119 18383 14153
rect 18265 14085 18343 14119
rect 18377 14085 18383 14119
rect 18265 14080 18383 14085
rect 18265 14046 18271 14080
rect 18305 14046 18383 14080
rect 18265 14012 18343 14046
rect 18377 14012 18383 14046
rect 18265 14007 18383 14012
rect 18265 13973 18271 14007
rect 18305 13973 18383 14007
rect 18265 13939 18343 13973
rect 18377 13939 18383 13973
rect 18265 13934 18383 13939
rect 18265 13900 18271 13934
rect 18305 13900 18383 13934
rect 18265 13866 18343 13900
rect 18377 13866 18383 13900
rect 18265 13861 18383 13866
rect 18265 13827 18271 13861
rect 18305 13827 18383 13861
rect 18265 13793 18343 13827
rect 18377 13793 18383 13827
rect 18265 13788 18383 13793
rect 18265 13754 18271 13788
rect 18305 13754 18383 13788
rect 18265 13720 18343 13754
rect 18377 13720 18383 13754
rect 18265 13715 18383 13720
rect 18265 13681 18271 13715
rect 18305 13681 18383 13715
rect 18265 13647 18343 13681
rect 18377 13647 18383 13681
rect 18265 13642 18383 13647
rect 18265 13608 18271 13642
rect 18305 13608 18383 13642
rect 18265 13574 18343 13608
rect 18377 13574 18383 13608
rect 18265 13569 18383 13574
rect 18265 13535 18271 13569
rect 18305 13535 18383 13569
rect 18265 13501 18343 13535
rect 18377 13501 18383 13535
rect 18265 13496 18383 13501
rect 18265 13462 18271 13496
rect 18305 13462 18383 13496
rect 18265 13428 18343 13462
rect 18377 13428 18383 13462
rect 18265 13423 18383 13428
rect 18265 13389 18271 13423
rect 18305 13389 18383 13423
rect 18265 13355 18343 13389
rect 18377 13355 18383 13389
rect 18265 13350 18383 13355
rect 18265 13316 18271 13350
rect 18305 13316 18383 13350
rect 18265 13282 18343 13316
rect 18377 13282 18383 13316
rect 18265 13277 18383 13282
rect 18265 13243 18271 13277
rect 18305 13243 18383 13277
rect 18265 13209 18343 13243
rect 18377 13209 18383 13243
rect 18265 13204 18383 13209
rect 18265 13170 18271 13204
rect 18305 13170 18383 13204
rect 18265 13136 18343 13170
rect 18377 13136 18383 13170
rect 18265 13131 18383 13136
rect 18265 13097 18271 13131
rect 18305 13097 18383 13131
rect 18265 13063 18343 13097
rect 18377 13063 18383 13097
rect 18265 13058 18383 13063
rect 18265 13024 18271 13058
rect 18305 13024 18383 13058
rect 18265 12990 18343 13024
rect 18377 12990 18383 13024
rect 18265 12985 18383 12990
rect 18265 12951 18271 12985
rect 18305 12951 18383 12985
rect 18265 12917 18343 12951
rect 18377 12917 18383 12951
rect 18265 12912 18383 12917
rect 18265 12878 18271 12912
rect 18305 12878 18383 12912
rect 18265 12844 18343 12878
rect 18377 12844 18383 12878
rect 18265 12839 18383 12844
rect 18265 12805 18271 12839
rect 18305 12805 18383 12839
rect 18265 12771 18343 12805
rect 18377 12771 18383 12805
rect 18265 12766 18383 12771
rect 18265 12732 18271 12766
rect 18305 12732 18383 12766
rect 18265 12698 18343 12732
rect 18377 12698 18383 12732
rect 18265 12693 18383 12698
rect 18265 12659 18271 12693
rect 18305 12659 18383 12693
tri 18240 12626 18265 12651 se
rect 18265 12626 18343 12659
rect 16024 12625 18343 12626
rect 18377 12625 18383 12659
rect 16024 12620 18383 12625
rect 16024 12586 16036 12620
rect 16070 12586 16109 12620
rect 16143 12586 16182 12620
rect 16216 12586 16255 12620
rect 16289 12586 16327 12620
rect 16361 12586 16399 12620
rect 16433 12586 16471 12620
rect 16505 12586 16543 12620
rect 16577 12586 16615 12620
rect 16649 12586 16687 12620
rect 16721 12586 16759 12620
rect 16793 12586 16831 12620
rect 16865 12586 16903 12620
rect 16937 12586 16975 12620
rect 17009 12586 17047 12620
rect 17081 12586 17119 12620
rect 17153 12586 17191 12620
rect 17225 12586 17263 12620
rect 17297 12586 17335 12620
rect 17369 12586 17407 12620
rect 17441 12586 17479 12620
rect 17513 12586 17551 12620
rect 17585 12586 17623 12620
rect 17657 12586 17695 12620
rect 17729 12586 17767 12620
rect 17801 12586 17839 12620
rect 17873 12586 17911 12620
rect 17945 12586 17983 12620
rect 18017 12586 18055 12620
rect 18089 12586 18127 12620
rect 18161 12586 18199 12620
rect 18233 12586 18271 12620
rect 18305 12586 18383 12620
rect 16024 12552 18343 12586
rect 18377 12552 18383 12586
rect 16024 12548 18383 12552
rect 16024 12514 16036 12548
rect 16070 12514 16110 12548
rect 16144 12514 16184 12548
rect 16218 12514 16258 12548
rect 16292 12514 16332 12548
rect 16366 12514 16406 12548
rect 16440 12514 16479 12548
rect 16513 12514 16552 12548
rect 16586 12514 16625 12548
rect 16659 12514 16698 12548
rect 16732 12514 16771 12548
rect 16805 12514 16844 12548
rect 16878 12514 16917 12548
rect 16951 12514 16990 12548
rect 17024 12514 17063 12548
rect 17097 12514 17136 12548
rect 17170 12514 17209 12548
rect 17243 12514 17282 12548
rect 17316 12514 17355 12548
rect 17389 12514 17428 12548
rect 17462 12514 17501 12548
rect 17535 12514 17574 12548
rect 17608 12514 17647 12548
rect 17681 12514 17720 12548
rect 17754 12514 17793 12548
rect 17827 12514 17866 12548
rect 17900 12514 17939 12548
rect 17973 12514 18012 12548
rect 18046 12514 18085 12548
rect 18119 12514 18158 12548
rect 18192 12514 18231 12548
rect 18265 12514 18383 12548
rect 16024 12508 18383 12514
rect 17004 7659 17062 7665
rect 17004 7625 17016 7659
rect 17050 7625 17062 7659
rect 17004 7619 17062 7625
rect 10161 3694 15805 3700
rect 10161 3656 10277 3694
rect 10161 3622 10167 3656
rect 10201 3622 10277 3656
rect 10161 3588 10239 3622
rect 10273 3588 10277 3622
rect 11785 3660 11789 3694
rect 11823 3660 11861 3694
rect 11895 3660 11933 3694
rect 11967 3660 12005 3694
rect 12039 3660 12077 3694
rect 12111 3660 12150 3694
rect 12184 3660 12223 3694
rect 12257 3660 12296 3694
rect 12330 3660 12369 3694
rect 12403 3660 12442 3694
rect 12476 3660 12515 3694
rect 12549 3660 12588 3694
rect 12622 3660 12661 3694
rect 12695 3660 12734 3694
rect 12768 3660 12807 3694
rect 12841 3660 12880 3694
rect 12914 3660 12953 3694
rect 12987 3660 13026 3694
rect 13060 3660 13099 3694
rect 13133 3660 13172 3694
rect 13206 3660 13245 3694
rect 13279 3660 13318 3694
rect 13352 3660 13391 3694
rect 13425 3660 13464 3694
rect 13498 3660 13537 3694
rect 13571 3660 13610 3694
rect 13644 3660 13683 3694
rect 13717 3660 13756 3694
rect 13790 3660 13829 3694
rect 13863 3660 13902 3694
rect 13936 3660 13975 3694
rect 14009 3660 14048 3694
rect 14082 3660 14121 3694
rect 14155 3660 14194 3694
rect 14228 3660 14267 3694
rect 14301 3660 14340 3694
rect 14374 3660 14413 3694
rect 14447 3660 14486 3694
rect 14520 3660 14559 3694
rect 14593 3660 14632 3694
rect 14666 3660 14705 3694
rect 14739 3660 14778 3694
rect 14812 3660 14851 3694
rect 14885 3660 14924 3694
rect 14958 3660 14997 3694
rect 15031 3660 15070 3694
rect 15104 3660 15143 3694
rect 15177 3660 15216 3694
rect 15250 3660 15289 3694
rect 15323 3660 15362 3694
rect 15396 3660 15435 3694
rect 15469 3660 15508 3694
rect 15542 3660 15581 3694
rect 15615 3660 15654 3694
rect 15688 3660 15727 3694
rect 15761 3660 15805 3694
rect 11785 3622 15805 3660
rect 11785 3588 11824 3622
rect 11858 3588 11897 3622
rect 11931 3588 11970 3622
rect 12004 3588 12043 3622
rect 12077 3588 12116 3622
rect 12150 3588 12189 3622
rect 12223 3588 12262 3622
rect 12296 3588 12335 3622
rect 12369 3588 12408 3622
rect 12442 3588 12481 3622
rect 12515 3588 12554 3622
rect 12588 3588 12627 3622
rect 12661 3588 12700 3622
rect 12734 3588 12773 3622
rect 12807 3588 12846 3622
rect 12880 3588 12919 3622
rect 12953 3588 12992 3622
rect 13026 3588 13065 3622
rect 13099 3588 13138 3622
rect 13172 3588 13211 3622
rect 13245 3588 13284 3622
rect 13318 3588 13357 3622
rect 13391 3588 13430 3622
rect 13464 3588 13503 3622
rect 13537 3588 13576 3622
rect 13610 3588 13649 3622
rect 13683 3588 13722 3622
rect 13756 3588 13795 3622
rect 13829 3588 13868 3622
rect 13902 3588 13941 3622
rect 13975 3588 14014 3622
rect 14048 3588 14087 3622
rect 14121 3588 14160 3622
rect 14194 3588 14233 3622
rect 14267 3588 14306 3622
rect 14340 3588 14379 3622
rect 14413 3588 14452 3622
rect 14486 3588 14525 3622
rect 14559 3588 14598 3622
rect 14632 3588 14671 3622
rect 14705 3588 14744 3622
rect 14778 3588 14817 3622
rect 14851 3588 14890 3622
rect 14924 3588 14963 3622
rect 14997 3588 15036 3622
rect 15070 3588 15109 3622
rect 15143 3588 15182 3622
rect 15216 3588 15255 3622
rect 15289 3588 15328 3622
rect 15362 3588 15401 3622
rect 15435 3588 15474 3622
rect 15508 3588 15547 3622
rect 15581 3588 15620 3622
rect 15654 3588 15693 3622
rect 15727 3588 15805 3622
rect 10161 3582 15805 3588
rect 10161 3576 10350 3582
rect 10161 3542 10167 3576
rect 10201 3550 10350 3576
tri 10350 3550 10382 3582 nw
tri 15662 3557 15687 3582 ne
rect 15687 3550 15765 3582
rect 10201 3546 10316 3550
rect 10201 3542 10239 3546
rect 10161 3512 10239 3542
rect 10273 3516 10316 3546
tri 10316 3516 10350 3550 nw
rect 15687 3516 15693 3550
rect 15727 3548 15765 3550
rect 15799 3548 15805 3582
rect 15727 3516 15805 3548
rect 10273 3512 10309 3516
rect 10161 3509 10309 3512
tri 10309 3509 10316 3516 nw
rect 15687 3509 15805 3516
rect 10161 3497 10279 3509
rect 10161 3463 10167 3497
rect 10201 3470 10279 3497
tri 10279 3479 10309 3509 nw
rect 10201 3463 10239 3470
rect 10161 3436 10239 3463
rect 10273 3436 10279 3470
rect 10161 3418 10279 3436
rect 10161 3384 10167 3418
rect 10201 3394 10279 3418
rect 10201 3384 10239 3394
rect 10161 3360 10239 3384
rect 10273 3360 10279 3394
rect 15687 3478 15765 3509
rect 15687 3444 15693 3478
rect 15727 3475 15765 3478
rect 15799 3475 15805 3509
rect 15727 3444 15805 3475
rect 15687 3436 15805 3444
rect 15687 3406 15765 3436
rect 10161 3339 10279 3360
rect 10161 3305 10167 3339
rect 10201 3319 10279 3339
rect 10201 3305 10239 3319
rect 10161 3285 10239 3305
rect 10273 3285 10279 3319
rect 10161 3260 10279 3285
rect 10161 3226 10167 3260
rect 10201 3244 10279 3260
rect 10201 3226 10239 3244
rect 10161 3210 10239 3226
rect 10273 3210 10279 3244
rect 10161 3181 10279 3210
rect 10161 3147 10167 3181
rect 10201 3169 10279 3181
rect 10201 3147 10239 3169
rect 10161 3135 10239 3147
rect 10273 3135 10279 3169
rect 10161 3102 10279 3135
rect 10161 3068 10167 3102
rect 10201 3094 10279 3102
rect 10201 3068 10239 3094
rect 10161 3060 10239 3068
rect 10273 3060 10279 3094
rect 10161 3023 10279 3060
rect 10161 2989 10167 3023
rect 10201 3019 10279 3023
rect 10201 2989 10239 3019
rect 10161 2985 10239 2989
rect 10273 2985 10279 3019
tri 10145 2944 10161 2960 se
rect 10161 2944 10279 2985
tri 10111 2910 10145 2944 se
rect 10145 2910 10167 2944
rect 10201 2910 10239 2944
rect 10273 2910 10279 2944
tri 10099 2898 10111 2910 se
rect 10111 2898 10279 2910
tri 10065 2864 10099 2898 se
rect 10099 2864 10279 2898
tri 10064 2863 10065 2864 se
rect 10065 2863 10279 2864
rect 10064 2826 10279 2863
rect 10517 3373 15483 3379
rect 10517 3335 10633 3373
rect 10517 3301 10523 3335
rect 10557 3301 10633 3335
rect 10517 3267 10595 3301
rect 10629 3267 10633 3301
rect 13653 3339 13657 3373
rect 13691 3339 13729 3373
rect 13763 3339 13801 3373
rect 13835 3339 13873 3373
rect 13907 3339 13945 3373
rect 13979 3339 14018 3373
rect 14052 3339 14091 3373
rect 14125 3339 14164 3373
rect 14198 3339 14237 3373
rect 14271 3339 14310 3373
rect 14344 3339 14383 3373
rect 14417 3339 14456 3373
rect 14490 3339 14529 3373
rect 14563 3339 14602 3373
rect 14636 3339 14675 3373
rect 14709 3339 14748 3373
rect 14782 3339 14821 3373
rect 14855 3339 14894 3373
rect 14928 3339 14967 3373
rect 15001 3339 15040 3373
rect 15074 3339 15113 3373
rect 15147 3339 15186 3373
rect 15220 3339 15259 3373
rect 15293 3339 15332 3373
rect 15366 3339 15405 3373
rect 15439 3339 15483 3373
rect 13653 3301 15483 3339
rect 13653 3267 13692 3301
rect 13726 3267 13765 3301
rect 13799 3267 13838 3301
rect 13872 3267 13911 3301
rect 13945 3267 13984 3301
rect 14018 3267 14057 3301
rect 14091 3267 14130 3301
rect 14164 3267 14203 3301
rect 14237 3267 14276 3301
rect 14310 3267 14349 3301
rect 14383 3267 14422 3301
rect 14456 3267 14495 3301
rect 14529 3267 14568 3301
rect 14602 3267 14641 3301
rect 14675 3267 14714 3301
rect 14748 3267 14787 3301
rect 14821 3267 14860 3301
rect 14894 3267 14933 3301
rect 14967 3267 15006 3301
rect 15040 3267 15079 3301
rect 15113 3267 15152 3301
rect 15186 3267 15225 3301
rect 15259 3267 15298 3301
rect 15332 3267 15371 3301
rect 15405 3267 15483 3301
rect 10517 3262 15483 3267
rect 10517 3228 10523 3262
rect 10557 3261 15483 3262
rect 10557 3228 10706 3261
tri 10706 3228 10739 3261 nw
tri 15299 3233 15327 3261 ne
rect 15327 3233 15443 3261
rect 10517 3227 10672 3228
rect 10517 3193 10595 3227
rect 10629 3194 10672 3227
tri 10672 3194 10706 3228 nw
rect 10629 3193 10668 3194
rect 10517 3190 10668 3193
tri 10668 3190 10672 3194 nw
rect 10517 3189 10666 3190
rect 10517 3155 10523 3189
rect 10557 3188 10666 3189
tri 10666 3188 10668 3190 nw
rect 10557 3155 10635 3188
tri 10635 3157 10666 3188 nw
rect 10517 3153 10635 3155
rect 10517 3119 10595 3153
rect 10629 3119 10635 3153
rect 10517 3116 10635 3119
rect 10517 3082 10523 3116
rect 10557 3082 10635 3116
rect 10517 3079 10635 3082
rect 10517 3045 10595 3079
rect 10629 3045 10635 3079
rect 10517 3043 10635 3045
rect 10517 3009 10523 3043
rect 10557 3009 10635 3043
rect 10517 3005 10635 3009
rect 10517 2971 10595 3005
rect 10629 2971 10635 3005
rect 10517 2970 10635 2971
rect 10517 2936 10523 2970
rect 10557 2936 10635 2970
rect 10517 2931 10635 2936
rect 10517 2898 10595 2931
rect 10517 2864 10523 2898
rect 10557 2897 10595 2898
rect 10629 2897 10635 2931
rect 10557 2864 10635 2897
rect 10517 2857 10635 2864
tri 10279 2826 10289 2836 sw
rect 10517 2826 10595 2857
rect 10064 2792 10289 2826
tri 10289 2792 10323 2826 sw
rect 10517 2792 10523 2826
rect 10557 2823 10595 2826
rect 10629 2823 10635 2857
rect 10557 2792 10635 2823
rect 10064 2790 10323 2792
tri 10323 2790 10325 2792 sw
rect 10064 2783 10325 2790
tri 10325 2783 10332 2790 sw
rect 10517 2783 10635 2792
rect 10064 2765 10332 2783
tri 10332 2765 10350 2783 sw
rect 10064 2713 10350 2765
rect 10517 2754 10595 2783
rect 10517 2720 10523 2754
rect 10557 2749 10595 2754
rect 10629 2749 10635 2783
rect 10557 2720 10635 2749
rect 10517 2709 10635 2720
rect 10517 2682 10595 2709
rect 10517 2648 10523 2682
rect 10557 2675 10595 2682
rect 10629 2675 10635 2709
rect 10836 2681 15164 3233
tri 15327 3228 15332 3233 ne
rect 15332 3228 15443 3233
tri 15332 3195 15365 3228 ne
rect 15365 3194 15371 3228
rect 15405 3227 15443 3228
rect 15477 3227 15483 3261
rect 15405 3194 15483 3227
rect 15365 3188 15483 3194
rect 15365 3155 15443 3188
rect 15365 3121 15371 3155
rect 15405 3154 15443 3155
rect 15477 3154 15483 3188
rect 15405 3121 15483 3154
rect 15365 3115 15483 3121
rect 15365 3082 15443 3115
rect 15365 3048 15371 3082
rect 15405 3081 15443 3082
rect 15477 3081 15483 3115
rect 15405 3048 15483 3081
rect 15365 3042 15483 3048
rect 15365 3009 15443 3042
rect 15365 2975 15371 3009
rect 15405 3008 15443 3009
rect 15477 3008 15483 3042
rect 15405 2975 15483 3008
rect 15365 2969 15483 2975
rect 15365 2936 15443 2969
rect 15365 2902 15371 2936
rect 15405 2935 15443 2936
rect 15477 2935 15483 2969
rect 15405 2902 15483 2935
rect 15365 2896 15483 2902
rect 15365 2863 15443 2896
rect 15365 2829 15371 2863
rect 15405 2862 15443 2863
rect 15477 2862 15483 2896
rect 15405 2829 15483 2862
rect 15365 2823 15483 2829
rect 15365 2790 15443 2823
rect 15365 2756 15371 2790
rect 15405 2789 15443 2790
rect 15477 2789 15483 2823
rect 15405 2756 15483 2789
rect 15365 2750 15483 2756
rect 15365 2717 15443 2750
rect 15365 2683 15371 2717
rect 15405 2716 15443 2717
rect 15477 2716 15483 2750
rect 15405 2683 15483 2716
rect 10557 2648 10635 2675
rect 10517 2636 10635 2648
rect 10517 2610 10595 2636
rect 10517 2576 10523 2610
rect 10557 2602 10595 2610
rect 10629 2602 10635 2636
rect 10557 2576 10635 2602
rect 10517 2563 10635 2576
rect 10517 2538 10595 2563
rect 10517 2504 10523 2538
rect 10557 2529 10595 2538
rect 10629 2529 10635 2563
rect 10557 2504 10635 2529
rect 10517 2490 10635 2504
rect 10517 2466 10595 2490
rect 10517 2432 10523 2466
rect 10557 2456 10595 2466
rect 10629 2456 10635 2490
rect 10557 2432 10635 2456
rect 10517 2417 10635 2432
rect 15365 2677 15483 2683
rect 15365 2644 15443 2677
rect 15365 2610 15371 2644
rect 15405 2643 15443 2644
rect 15477 2643 15483 2677
rect 15405 2610 15483 2643
rect 15365 2604 15483 2610
rect 15365 2571 15443 2604
rect 15365 2537 15371 2571
rect 15405 2570 15443 2571
rect 15477 2570 15483 2604
rect 15405 2537 15483 2570
rect 15365 2531 15483 2537
rect 15365 2498 15443 2531
rect 15365 2464 15371 2498
rect 15405 2497 15443 2498
rect 15477 2497 15483 2531
rect 15405 2464 15483 2497
rect 15365 2458 15483 2464
rect 15365 2425 15443 2458
rect 10517 2394 10595 2417
rect 10517 2360 10523 2394
rect 10557 2383 10595 2394
rect 10629 2383 10635 2417
rect 10557 2360 10635 2383
rect 10517 2344 10635 2360
rect 10517 2322 10595 2344
rect 10517 2288 10523 2322
rect 10557 2310 10595 2322
rect 10629 2310 10635 2344
rect 10557 2288 10635 2310
rect 10517 2271 10635 2288
rect 10517 2250 10595 2271
rect 10517 2216 10523 2250
rect 10557 2237 10595 2250
rect 10629 2237 10635 2271
rect 10557 2216 10635 2237
rect 10517 2198 10635 2216
rect 10517 2178 10595 2198
rect 10517 2144 10523 2178
rect 10557 2164 10595 2178
rect 10629 2164 10635 2198
rect 10557 2144 10635 2164
rect 10517 2125 10635 2144
rect 10517 2106 10595 2125
rect 10517 2072 10523 2106
rect 10557 2091 10595 2106
rect 10629 2091 10635 2125
rect 10557 2072 10635 2091
rect 10517 2052 10635 2072
rect 10517 2034 10595 2052
rect 10517 2000 10523 2034
rect 10557 2018 10595 2034
rect 10629 2018 10635 2052
rect 10557 2000 10635 2018
rect 10517 1979 10635 2000
rect 10517 1962 10595 1979
rect 10517 1928 10523 1962
rect 10557 1945 10595 1962
rect 10629 1945 10635 1979
rect 10557 1928 10635 1945
rect 10517 1906 10635 1928
rect 10517 1890 10595 1906
rect 10517 1856 10523 1890
rect 10557 1872 10595 1890
rect 10629 1872 10635 1906
rect 10557 1856 10635 1872
rect 10517 1833 10635 1856
rect 10517 1818 10595 1833
rect 10517 1784 10523 1818
rect 10557 1799 10595 1818
rect 10629 1799 10635 1833
rect 10557 1784 10635 1799
rect 10517 1760 10635 1784
rect 10517 1746 10595 1760
rect 10517 1712 10523 1746
rect 10557 1726 10595 1746
rect 10629 1726 10635 1760
rect 10557 1712 10635 1726
rect 10517 1687 10635 1712
rect 10517 1674 10595 1687
rect 10517 1640 10523 1674
rect 10557 1653 10595 1674
rect 10629 1653 10635 1687
rect 10557 1640 10635 1653
rect 10517 1614 10635 1640
rect 10517 1602 10595 1614
rect 10517 1568 10523 1602
rect 10557 1580 10595 1602
rect 10629 1580 10635 1614
rect 10557 1568 10635 1580
rect 10517 1541 10635 1568
rect 10517 1530 10595 1541
rect 10517 1496 10523 1530
rect 10557 1507 10595 1530
rect 10629 1507 10635 1541
rect 10703 2406 10749 2418
rect 10703 2372 10709 2406
rect 10743 2372 10749 2406
rect 10703 2330 10749 2372
rect 15251 2406 15297 2418
rect 15251 2372 15257 2406
rect 15291 2372 15297 2406
rect 10703 2296 10709 2330
rect 10743 2296 10749 2330
rect 10703 2253 10749 2296
rect 10703 2219 10709 2253
rect 10743 2219 10749 2253
rect 10703 2176 10749 2219
rect 10703 2142 10709 2176
rect 10743 2142 10749 2176
rect 12946 2336 14989 2342
rect 12946 2220 14873 2336
rect 12946 2214 14989 2220
rect 15251 2330 15297 2372
rect 15251 2296 15257 2330
rect 15291 2296 15297 2330
rect 15251 2253 15297 2296
rect 15251 2219 15257 2253
rect 15291 2219 15297 2253
rect 12946 2206 13079 2214
tri 13079 2206 13087 2214 nw
tri 10749 2142 10762 2155 sw
tri 12933 2142 12946 2155 se
rect 12946 2142 13062 2206
tri 13062 2189 13079 2206 nw
rect 15251 2176 15297 2219
tri 13062 2142 13075 2155 sw
tri 15238 2142 15251 2155 se
rect 15251 2142 15257 2176
rect 15291 2142 15297 2176
rect 10703 2133 10762 2142
tri 10762 2133 10771 2142 sw
tri 12924 2133 12933 2142 se
rect 12933 2133 13075 2142
tri 13075 2133 13084 2142 sw
tri 15229 2133 15238 2142 se
rect 15238 2133 15297 2142
rect 10703 2130 10771 2133
tri 10771 2130 10774 2133 sw
tri 12921 2130 12924 2133 se
rect 12924 2130 13084 2133
tri 13084 2130 13087 2133 sw
tri 15226 2130 15229 2133 se
rect 15229 2130 15297 2133
rect 10703 2099 12726 2130
rect 12728 2129 12764 2130
rect 10703 2065 10709 2099
rect 10743 2065 12726 2099
rect 10703 2022 12726 2065
rect 10703 1988 10709 2022
rect 10743 1997 12726 2022
rect 12727 1998 12765 2129
rect 12766 2118 13242 2130
rect 13244 2129 13280 2130
rect 12766 2012 12951 2118
rect 13057 2012 13242 2118
rect 12728 1997 12764 1998
rect 12766 1997 13242 2012
rect 13243 1998 13281 2129
rect 13282 2099 15297 2130
rect 13282 2065 15257 2099
rect 15291 2065 15297 2099
rect 13282 2022 15297 2065
rect 13244 1997 13280 1998
rect 13282 1997 15257 2022
rect 10743 1988 12705 1997
tri 12705 1988 12714 1997 nw
tri 13294 1988 13303 1997 ne
rect 13303 1988 15257 1997
rect 15291 1988 15297 2022
rect 10703 1987 12704 1988
tri 12704 1987 12705 1988 nw
tri 13303 1987 13304 1988 ne
rect 13304 1987 15297 1988
rect 10703 1945 12689 1987
tri 12689 1972 12704 1987 nw
tri 13304 1972 13319 1987 ne
rect 10703 1911 10709 1945
rect 10743 1919 12689 1945
rect 13319 1945 15297 1987
tri 12689 1919 12714 1944 sw
tri 13294 1919 13319 1944 se
rect 13319 1919 15257 1945
rect 10743 1911 12726 1919
rect 10703 1868 12726 1911
rect 10703 1834 10709 1868
rect 10743 1834 12726 1868
rect 10703 1791 12726 1834
rect 10703 1757 10709 1791
rect 10743 1786 12726 1791
rect 12727 1787 12728 1918
rect 12764 1787 12765 1918
rect 12766 1908 13242 1919
rect 12766 1792 12946 1908
rect 13062 1792 13242 1908
rect 12766 1786 13242 1792
rect 13243 1787 13244 1918
rect 13280 1787 13281 1918
rect 13282 1911 15257 1919
rect 15291 1911 15297 1945
rect 13282 1868 15297 1911
rect 13282 1834 15257 1868
rect 15291 1834 15297 1868
rect 13282 1791 15297 1834
rect 13282 1786 15257 1791
rect 10743 1757 10749 1786
tri 10749 1761 10774 1786 nw
tri 15226 1761 15251 1786 ne
rect 10703 1714 10749 1757
rect 10703 1680 10709 1714
rect 10743 1680 10749 1714
rect 10703 1637 10749 1680
rect 10703 1603 10709 1637
rect 10743 1603 10749 1637
rect 10703 1560 10749 1603
rect 10703 1526 10709 1560
rect 10743 1526 10749 1560
rect 10703 1514 10749 1526
rect 15251 1757 15257 1786
rect 15291 1757 15297 1791
rect 15251 1714 15297 1757
rect 15251 1680 15257 1714
rect 15291 1680 15297 1714
rect 15251 1637 15297 1680
rect 15251 1603 15257 1637
rect 15291 1603 15297 1637
rect 15251 1560 15297 1603
rect 15251 1526 15257 1560
rect 15291 1526 15297 1560
rect 15251 1514 15297 1526
rect 15365 2391 15371 2425
rect 15405 2424 15443 2425
rect 15477 2424 15483 2458
rect 15405 2391 15483 2424
rect 15365 2385 15483 2391
rect 15365 2352 15443 2385
rect 15365 2318 15371 2352
rect 15405 2351 15443 2352
rect 15477 2351 15483 2385
rect 15405 2318 15483 2351
rect 15365 2312 15483 2318
rect 15365 2279 15443 2312
rect 15365 2245 15371 2279
rect 15405 2278 15443 2279
rect 15477 2278 15483 2312
rect 15405 2245 15483 2278
rect 15365 2239 15483 2245
rect 15365 2206 15443 2239
rect 15365 2172 15371 2206
rect 15405 2205 15443 2206
rect 15477 2205 15483 2239
rect 15405 2172 15483 2205
rect 15365 2166 15483 2172
rect 15365 2133 15443 2166
rect 15365 2099 15371 2133
rect 15405 2132 15443 2133
rect 15477 2132 15483 2166
rect 15405 2099 15483 2132
rect 15365 2093 15483 2099
rect 15365 2060 15443 2093
rect 15365 2026 15371 2060
rect 15405 2059 15443 2060
rect 15477 2059 15483 2093
rect 15405 2026 15483 2059
rect 15365 2020 15483 2026
rect 15365 1987 15443 2020
rect 15365 1953 15371 1987
rect 15405 1986 15443 1987
rect 15477 1986 15483 2020
rect 15405 1953 15483 1986
rect 15365 1947 15483 1953
rect 15365 1914 15443 1947
rect 15365 1880 15371 1914
rect 15405 1913 15443 1914
rect 15477 1913 15483 1947
rect 15405 1880 15483 1913
rect 15365 1874 15483 1880
rect 15365 1841 15443 1874
rect 15365 1807 15371 1841
rect 15405 1840 15443 1841
rect 15477 1840 15483 1874
rect 15405 1807 15483 1840
rect 15365 1801 15483 1807
rect 15365 1768 15443 1801
rect 15365 1734 15371 1768
rect 15405 1767 15443 1768
rect 15477 1767 15483 1801
rect 15405 1734 15483 1767
rect 15365 1728 15483 1734
rect 15365 1695 15443 1728
rect 15365 1661 15371 1695
rect 15405 1694 15443 1695
rect 15477 1694 15483 1728
rect 15405 1661 15483 1694
rect 15365 1655 15483 1661
rect 15365 1622 15443 1655
rect 15365 1588 15371 1622
rect 15405 1621 15443 1622
rect 15477 1621 15483 1655
rect 15405 1588 15483 1621
rect 15365 1582 15483 1588
rect 15365 1549 15443 1582
rect 15365 1515 15371 1549
rect 15405 1548 15443 1549
rect 15477 1548 15483 1582
rect 15405 1515 15483 1548
rect 10557 1496 10635 1507
rect 10517 1468 10635 1496
rect 10517 1458 10595 1468
rect 10517 1424 10523 1458
rect 10557 1434 10595 1458
rect 10629 1434 10635 1468
rect 10557 1424 10635 1434
rect 10517 1395 10635 1424
rect 10517 1386 10595 1395
rect 10517 1352 10523 1386
rect 10557 1361 10595 1386
rect 10629 1361 10635 1395
rect 10557 1352 10635 1361
rect 10517 1322 10635 1352
rect 10517 1314 10595 1322
rect 10517 1280 10523 1314
rect 10557 1288 10595 1314
rect 10629 1288 10635 1322
rect 10557 1280 10635 1288
rect 10517 1249 10635 1280
rect 15365 1509 15483 1515
rect 15365 1476 15443 1509
rect 15365 1442 15371 1476
rect 15405 1475 15443 1476
rect 15477 1475 15483 1509
rect 15405 1442 15483 1475
rect 15365 1436 15483 1442
rect 15365 1403 15443 1436
rect 15365 1369 15371 1403
rect 15405 1402 15443 1403
rect 15477 1402 15483 1436
rect 15405 1369 15483 1402
rect 15365 1363 15483 1369
rect 15365 1330 15443 1363
rect 15365 1296 15371 1330
rect 15405 1329 15443 1330
rect 15477 1329 15483 1363
rect 15405 1296 15483 1329
rect 15365 1290 15483 1296
rect 15365 1257 15443 1290
rect 10517 1242 10595 1249
rect 10517 1208 10523 1242
rect 10557 1215 10595 1242
rect 10629 1215 10635 1249
rect 10557 1208 10635 1215
rect 10517 1176 10635 1208
rect 10517 1170 10595 1176
rect 10517 1136 10523 1170
rect 10557 1142 10595 1170
rect 10629 1142 10635 1176
rect 10557 1136 10635 1142
rect 10517 1103 10635 1136
rect 10517 1098 10595 1103
rect 10517 1064 10523 1098
rect 10557 1069 10595 1098
rect 10629 1069 10635 1103
rect 10557 1064 10635 1069
rect 10517 1030 10635 1064
rect 10517 1026 10595 1030
rect 10517 992 10523 1026
rect 10557 996 10595 1026
rect 10629 996 10635 1030
rect 10557 992 10635 996
rect 10517 957 10635 992
rect 10517 954 10595 957
rect 10517 920 10523 954
rect 10557 923 10595 954
rect 10629 923 10635 957
rect 10557 920 10635 923
rect 10517 884 10635 920
rect 10517 882 10595 884
rect 10517 848 10523 882
rect 10557 850 10595 882
rect 10629 850 10635 884
rect 10557 848 10635 850
rect 10517 811 10635 848
rect 10517 810 10595 811
rect 10517 776 10523 810
rect 10557 777 10595 810
rect 10629 777 10635 811
rect 10557 776 10635 777
rect 10517 738 10635 776
rect 10517 704 10523 738
rect 10557 704 10595 738
rect 10629 704 10635 738
rect 10517 671 10635 704
rect 10836 699 15164 1251
rect 15365 1223 15371 1257
rect 15405 1256 15443 1257
rect 15477 1256 15483 1290
rect 15405 1223 15483 1256
rect 15365 1217 15483 1223
rect 15365 1183 15443 1217
rect 15477 1183 15483 1217
rect 15365 1149 15371 1183
rect 15405 1149 15483 1183
rect 15365 1144 15483 1149
rect 15365 1110 15443 1144
rect 15477 1110 15483 1144
rect 15365 1109 15483 1110
rect 15365 1075 15371 1109
rect 15405 1075 15483 1109
rect 15365 1071 15483 1075
rect 15365 1037 15443 1071
rect 15477 1037 15483 1071
rect 15365 1035 15483 1037
rect 15365 1001 15371 1035
rect 15405 1001 15483 1035
rect 15365 998 15483 1001
rect 15365 964 15443 998
rect 15477 964 15483 998
rect 15365 961 15483 964
rect 15365 927 15371 961
rect 15405 927 15483 961
rect 15365 925 15483 927
rect 15365 891 15443 925
rect 15477 891 15483 925
rect 15365 887 15483 891
rect 15365 853 15371 887
rect 15405 853 15483 887
rect 15365 852 15483 853
rect 15365 818 15443 852
rect 15477 818 15483 852
rect 15365 813 15483 818
rect 15365 779 15371 813
rect 15405 779 15483 813
rect 15365 745 15443 779
rect 15477 745 15483 779
rect 15365 739 15483 745
rect 15365 705 15371 739
rect 15405 705 15483 739
tri 10635 671 10660 696 sw
tri 15340 671 15365 696 se
rect 15365 671 15443 705
rect 15477 671 15483 705
rect 10517 665 15483 671
rect 10517 631 10529 665
rect 10563 631 10602 665
rect 10636 631 10675 665
rect 10709 631 10748 665
rect 10782 631 10821 665
rect 10855 631 10894 665
rect 10928 631 10967 665
rect 11001 631 11040 665
rect 11074 631 11113 665
rect 11147 631 11186 665
rect 11220 631 11259 665
rect 11293 631 11332 665
rect 11366 631 11405 665
rect 11439 631 11478 665
rect 11512 631 11551 665
rect 11585 631 11624 665
rect 11658 631 11697 665
rect 11731 631 11770 665
rect 11804 631 11843 665
rect 11877 631 11915 665
rect 11949 631 11987 665
rect 12021 631 12059 665
rect 12093 631 12131 665
rect 12165 631 12203 665
rect 12237 631 12275 665
rect 12309 631 12347 665
rect 12381 631 12419 665
rect 12453 631 12491 665
rect 12525 631 12563 665
rect 12597 631 12635 665
rect 12669 631 12707 665
rect 12741 631 12779 665
rect 12813 631 12851 665
rect 12885 631 12923 665
rect 12957 631 12995 665
rect 13029 631 13067 665
rect 13101 631 13139 665
rect 13173 631 13211 665
rect 13245 631 13283 665
rect 13317 631 13355 665
rect 13389 631 13427 665
rect 13461 631 13499 665
rect 13533 631 13571 665
rect 13605 631 13643 665
rect 13677 631 13715 665
rect 13749 631 13787 665
rect 13821 631 13859 665
rect 13893 631 13931 665
rect 13965 631 14003 665
rect 14037 631 14075 665
rect 14109 631 14147 665
rect 14181 631 14219 665
rect 14253 631 14291 665
rect 15367 631 15371 665
rect 15405 631 15483 665
rect 10517 593 14325 631
rect 10517 559 10529 593
rect 10563 559 10602 593
rect 10636 559 10675 593
rect 10709 559 10748 593
rect 10782 559 10821 593
rect 10855 559 10894 593
rect 10928 559 10967 593
rect 11001 559 11040 593
rect 11074 559 11113 593
rect 11147 559 11186 593
rect 11220 559 11259 593
rect 11293 559 11332 593
rect 11366 559 11405 593
rect 11439 559 11478 593
rect 11512 559 11551 593
rect 11585 559 11624 593
rect 11658 559 11697 593
rect 11731 559 11770 593
rect 11804 559 11843 593
rect 11877 559 11916 593
rect 11950 559 11989 593
rect 12023 559 12062 593
rect 12096 559 12135 593
rect 12169 559 12208 593
rect 12242 559 12281 593
rect 12315 559 12354 593
rect 12388 559 12427 593
rect 12461 559 12500 593
rect 12534 559 12573 593
rect 12607 559 12646 593
rect 12680 559 12719 593
rect 12753 559 12792 593
rect 12826 559 12865 593
rect 12899 559 12938 593
rect 12972 559 13011 593
rect 13045 559 13084 593
rect 13118 559 13157 593
rect 13191 559 13230 593
rect 13264 559 13303 593
rect 13337 559 13376 593
rect 13410 559 13449 593
rect 13483 559 13522 593
rect 13556 559 13595 593
rect 13629 559 13668 593
rect 13702 559 13741 593
rect 13775 559 13814 593
rect 13848 559 13887 593
rect 13921 559 13960 593
rect 13994 559 14033 593
rect 14067 559 14106 593
rect 14140 559 14179 593
rect 14213 559 14252 593
rect 14286 559 14325 593
rect 15367 597 15443 631
rect 15477 597 15483 631
rect 15367 559 15483 597
rect 10517 553 15483 559
rect 15687 3372 15693 3406
rect 15727 3402 15765 3406
rect 15799 3402 15805 3436
rect 15727 3372 15805 3402
rect 15687 3363 15805 3372
rect 15687 3334 15765 3363
rect 15687 3300 15693 3334
rect 15727 3329 15765 3334
rect 15799 3329 15805 3363
rect 15727 3300 15805 3329
rect 15687 3290 15805 3300
rect 15687 3262 15765 3290
rect 15687 3228 15693 3262
rect 15727 3256 15765 3262
rect 15799 3256 15805 3290
rect 15727 3228 15805 3256
rect 15687 3217 15805 3228
rect 15687 3190 15765 3217
rect 15687 3156 15693 3190
rect 15727 3183 15765 3190
rect 15799 3183 15805 3217
rect 15727 3156 15805 3183
rect 15687 3144 15805 3156
rect 15687 3118 15765 3144
rect 15687 3084 15693 3118
rect 15727 3110 15765 3118
rect 15799 3110 15805 3144
rect 15727 3084 15805 3110
rect 15687 3071 15805 3084
rect 15687 3046 15765 3071
rect 15687 3012 15693 3046
rect 15727 3037 15765 3046
rect 15799 3037 15805 3071
rect 15727 3012 15805 3037
rect 15687 2998 15805 3012
rect 15687 2974 15765 2998
rect 15687 2940 15693 2974
rect 15727 2964 15765 2974
rect 15799 2964 15805 2998
rect 15727 2940 15805 2964
rect 15687 2925 15805 2940
rect 15687 2902 15765 2925
rect 15687 2868 15693 2902
rect 15727 2891 15765 2902
rect 15799 2891 15805 2925
rect 15727 2868 15805 2891
rect 15687 2852 15805 2868
rect 15687 2830 15765 2852
rect 15687 2796 15693 2830
rect 15727 2818 15765 2830
rect 15799 2818 15805 2852
rect 15727 2796 15805 2818
rect 15687 2779 15805 2796
rect 15687 2758 15765 2779
rect 15687 2724 15693 2758
rect 15727 2745 15765 2758
rect 15799 2745 15805 2779
rect 15727 2724 15805 2745
rect 15687 2706 15805 2724
rect 15687 2686 15765 2706
rect 15687 2652 15693 2686
rect 15727 2672 15765 2686
rect 15799 2672 15805 2706
rect 15727 2652 15805 2672
rect 15687 2633 15805 2652
rect 15687 2614 15765 2633
rect 15687 2580 15693 2614
rect 15727 2599 15765 2614
rect 15799 2599 15805 2633
rect 15727 2580 15805 2599
rect 15687 2560 15805 2580
rect 15687 2542 15765 2560
rect 15687 2508 15693 2542
rect 15727 2526 15765 2542
rect 15799 2526 15805 2560
rect 15727 2508 15805 2526
rect 15687 2487 15805 2508
rect 15687 2469 15765 2487
rect 15687 2435 15693 2469
rect 15727 2453 15765 2469
rect 15799 2453 15805 2487
rect 15727 2435 15805 2453
rect 15687 2414 15805 2435
rect 15687 2396 15765 2414
rect 15687 2362 15693 2396
rect 15727 2380 15765 2396
rect 15799 2380 15805 2414
rect 15727 2362 15805 2380
rect 15687 2341 15805 2362
rect 15687 2323 15765 2341
rect 15687 2289 15693 2323
rect 15727 2307 15765 2323
rect 15799 2307 15805 2341
rect 15727 2289 15805 2307
rect 15687 2268 15805 2289
rect 15687 2250 15765 2268
rect 15687 2216 15693 2250
rect 15727 2234 15765 2250
rect 15799 2234 15805 2268
rect 15727 2216 15805 2234
rect 15687 2195 15805 2216
rect 15687 2177 15765 2195
rect 15687 2143 15693 2177
rect 15727 2161 15765 2177
rect 15799 2161 15805 2195
rect 15727 2143 15805 2161
rect 15687 2122 15805 2143
rect 15687 2104 15765 2122
rect 15687 2070 15693 2104
rect 15727 2088 15765 2104
rect 15799 2088 15805 2122
rect 15727 2070 15805 2088
rect 15687 2049 15805 2070
rect 15687 2031 15765 2049
rect 15687 1997 15693 2031
rect 15727 2015 15765 2031
rect 15799 2015 15805 2049
rect 15727 1997 15805 2015
rect 15687 1976 15805 1997
rect 15687 1958 15765 1976
rect 15687 1924 15693 1958
rect 15727 1942 15765 1958
rect 15799 1942 15805 1976
rect 15727 1924 15805 1942
rect 15687 1903 15805 1924
rect 15687 1885 15765 1903
rect 15687 1851 15693 1885
rect 15727 1869 15765 1885
rect 15799 1869 15805 1903
rect 15727 1851 15805 1869
rect 15687 1830 15805 1851
rect 15687 1812 15765 1830
rect 15687 1778 15693 1812
rect 15727 1796 15765 1812
rect 15799 1796 15805 1830
rect 15727 1778 15805 1796
rect 15687 1757 15805 1778
rect 15687 1739 15765 1757
rect 15687 1705 15693 1739
rect 15727 1723 15765 1739
rect 15799 1723 15805 1757
rect 15727 1705 15805 1723
rect 15687 1684 15805 1705
rect 15687 1666 15765 1684
rect 15687 1632 15693 1666
rect 15727 1650 15765 1666
rect 15799 1650 15805 1684
rect 15727 1632 15805 1650
rect 15687 1610 15805 1632
rect 15687 1593 15765 1610
rect 15687 1559 15693 1593
rect 15727 1576 15765 1593
rect 15799 1576 15805 1610
rect 15727 1559 15805 1576
rect 15687 1536 15805 1559
rect 15687 1520 15765 1536
rect 15687 1486 15693 1520
rect 15727 1502 15765 1520
rect 15799 1502 15805 1536
rect 15727 1486 15805 1502
rect 15687 1462 15805 1486
rect 15687 1447 15765 1462
rect 15687 1413 15693 1447
rect 15727 1428 15765 1447
rect 15799 1428 15805 1462
rect 15727 1413 15805 1428
rect 15687 1388 15805 1413
rect 15687 1374 15765 1388
rect 15687 1340 15693 1374
rect 15727 1354 15765 1374
rect 15799 1354 15805 1388
rect 15727 1340 15805 1354
rect 15687 1314 15805 1340
rect 15687 1301 15765 1314
rect 15687 1267 15693 1301
rect 15727 1280 15765 1301
rect 15799 1280 15805 1314
rect 15727 1267 15805 1280
rect 15687 1240 15805 1267
rect 15687 1228 15765 1240
rect 15687 1194 15693 1228
rect 15727 1206 15765 1228
rect 15799 1206 15805 1240
rect 15727 1194 15805 1206
rect 15687 1166 15805 1194
rect 15687 1155 15765 1166
rect 15687 1121 15693 1155
rect 15727 1132 15765 1155
rect 15799 1132 15805 1166
rect 15727 1121 15805 1132
rect 15687 1092 15805 1121
rect 15687 1082 15765 1092
rect 15687 1048 15693 1082
rect 15727 1058 15765 1082
rect 15799 1058 15805 1092
rect 15727 1048 15805 1058
rect 15687 1018 15805 1048
rect 15687 1009 15765 1018
rect 15687 975 15693 1009
rect 15727 984 15765 1009
rect 15799 984 15805 1018
rect 15727 975 15805 984
rect 15687 944 15805 975
rect 15687 936 15765 944
rect 15687 902 15693 936
rect 15727 910 15765 936
rect 15799 910 15805 944
rect 15727 902 15805 910
rect 15687 870 15805 902
rect 15687 863 15765 870
rect 15687 829 15693 863
rect 15727 836 15765 863
rect 15799 836 15805 870
rect 15727 829 15805 836
rect 15687 796 15805 829
rect 15687 790 15765 796
rect 15687 756 15693 790
rect 15727 762 15765 790
rect 15799 762 15805 796
rect 15727 756 15805 762
rect 15687 722 15805 756
rect 15687 717 15765 722
rect 15687 683 15693 717
rect 15727 688 15765 717
rect 15799 688 15805 722
rect 15727 683 15805 688
rect 15687 648 15805 683
rect 15687 644 15765 648
rect 15687 610 15693 644
rect 15727 614 15765 644
rect 15799 614 15805 648
rect 15727 610 15805 614
rect 15687 574 15805 610
rect 15687 571 15765 574
tri 10778 537 10794 553 ne
rect 10794 537 10930 553
tri 10930 537 10946 553 nw
rect 15687 537 15693 571
rect 15727 540 15765 571
rect 15799 540 15805 574
rect 15727 537 15805 540
tri 10794 528 10803 537 ne
rect 10803 399 10921 537
tri 10921 528 10930 537 nw
rect 15687 500 15805 537
rect 15687 498 15765 500
rect 15687 464 15693 498
rect 15727 466 15765 498
rect 15799 466 15805 500
rect 15727 464 15805 466
rect 15687 426 15805 464
rect 15687 425 15765 426
rect 10803 365 10809 399
rect 10843 365 10881 399
rect 10915 365 10921 399
rect 10803 353 10921 365
rect 12945 408 13063 414
rect 12945 356 12946 408
rect 12998 356 13010 408
rect 13062 356 13063 408
rect 12945 350 13063 356
rect 15687 391 15693 425
rect 15727 392 15765 425
rect 15799 392 15805 426
rect 15727 391 15805 392
rect 15687 352 15805 391
rect 15687 318 15693 352
rect 15727 318 15765 352
rect 15799 318 15805 352
rect 15687 286 15805 318
<< rmetal1 >>
rect 15079 16472 15081 16473
rect 15079 16416 15080 16472
rect 15079 16415 15081 16416
rect 15117 16472 15119 16473
rect 15118 16416 15119 16472
rect 15117 16415 15119 16416
rect 15079 16326 15081 16327
rect 15117 16326 15119 16327
rect 15079 16270 15080 16326
rect 15118 16270 15119 16326
rect 15079 16269 15081 16270
rect 15117 16269 15119 16270
rect 10651 16192 14861 16193
rect 10651 16191 10652 16192
rect 14860 16191 14861 16192
rect 15079 16240 15081 16241
rect 15117 16240 15119 16241
rect 15079 16184 15080 16240
rect 15118 16184 15119 16240
rect 15079 16183 15081 16184
rect 15117 16183 15119 16184
rect 10651 16134 10652 16135
rect 14860 16134 14861 16135
rect 10651 16133 14861 16134
rect 15079 16094 15081 16095
rect 15079 16038 15080 16094
rect 15079 16037 15081 16038
rect 15117 16094 15119 16095
rect 15118 16038 15119 16094
rect 15117 16037 15119 16038
rect 15092 15051 15094 15052
rect 15130 15051 15132 15052
rect 15092 14995 15093 15051
rect 15131 14995 15132 15051
rect 15092 14994 15094 14995
rect 15130 14994 15132 14995
rect 13035 14952 14861 14953
rect 13035 14951 13036 14952
rect 14860 14951 14861 14952
rect 13035 14894 13036 14895
rect 14860 14894 14861 14895
rect 13035 14893 14861 14894
rect 15078 14915 15080 14916
rect 15078 14859 15079 14915
rect 15078 14858 15080 14859
rect 15116 14915 15118 14916
rect 15117 14859 15118 14915
rect 15116 14858 15118 14859
rect 15078 14582 15080 14583
rect 15078 14526 15079 14582
rect 15078 14525 15080 14526
rect 15116 14582 15118 14583
rect 15117 14526 15118 14582
rect 15116 14525 15118 14526
rect 15092 14446 15094 14447
rect 15130 14446 15132 14447
rect 15092 14390 15093 14446
rect 15131 14390 15132 14446
rect 15092 14389 15094 14390
rect 15130 14389 15132 14390
rect 15079 13149 15081 13150
rect 15117 13149 15119 13150
rect 15079 13093 15080 13149
rect 15118 13093 15119 13149
rect 15079 13092 15081 13093
rect 15117 13092 15119 13093
rect 15079 13013 15081 13014
rect 15079 12957 15080 13013
rect 15079 12956 15081 12957
rect 15117 13013 15119 13014
rect 15118 12957 15119 13013
rect 15117 12956 15119 12957
rect 12726 2129 12728 2130
rect 12764 2129 12766 2130
rect 12726 1998 12727 2129
rect 12765 1998 12766 2129
rect 13242 2129 13244 2130
rect 13280 2129 13282 2130
rect 12726 1997 12728 1998
rect 12764 1997 12766 1998
rect 13242 1998 13243 2129
rect 13281 1998 13282 2129
rect 13242 1997 13244 1998
rect 13280 1997 13282 1998
rect 12726 1918 12728 1919
rect 12726 1787 12727 1918
rect 12726 1786 12728 1787
rect 12764 1918 12766 1919
rect 12765 1787 12766 1918
rect 13242 1918 13244 1919
rect 12764 1786 12766 1787
rect 13242 1787 13243 1918
rect 13242 1786 13244 1787
rect 13280 1918 13282 1919
rect 13281 1787 13282 1918
rect 13280 1786 13282 1787
<< via1 >>
rect 14873 2220 14989 2336
rect 12946 1907 13062 1908
rect 12946 1801 12951 1907
rect 12951 1801 13057 1907
rect 13057 1801 13062 1907
rect 12946 1792 13062 1801
rect 12946 399 12998 408
rect 12946 365 12951 399
rect 12951 365 12985 399
rect 12985 365 12998 399
rect 12946 356 12998 365
rect 13010 399 13062 408
rect 13010 365 13023 399
rect 13023 365 13057 399
rect 13057 365 13062 399
rect 13010 356 13062 365
<< metal2 >>
rect 14873 2336 14989 3430
rect 15017 3191 15145 3430
rect 14873 2214 14989 2220
rect 12946 1908 13062 1919
rect 10844 695 12895 1249
rect 12946 408 13062 1792
rect 13397 695 15155 1249
rect 12998 356 13010 408
rect 12946 350 13062 356
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 -1 15075 -1 0 16315
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform -1 0 15193 0 1 14804
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform -1 0 15193 0 -1 14637
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 0 1 15533 1 0 13009
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform 0 1 15387 1 0 13009
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform 0 1 15241 1 0 13009
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1704896540
transform 0 1 10809 1 0 365
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1704896540
transform 0 1 12951 1 0 365
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1704896540
transform 0 -1 14929 1 0 13104
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1704896540
transform 0 -1 15075 1 0 13104
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1704896540
transform 0 -1 15229 1 0 13104
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1704896540
transform 0 -1 15075 1 0 16195
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1704896540
transform 1 0 15162 0 -1 16381
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1704896540
transform 1 0 15162 0 1 16129
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 1 14986 1 0 14537
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 1 14986 1 0 14870
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1704896540
transform 0 1 12951 1 0 2012
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_1
timestamp 1704896540
transform 0 1 12951 1 0 1801
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform 1 0 17016 0 1 7625
box 0 0 1 1
use L1M1_CDNS_524688791851562  L1M1_CDNS_524688791851562_0
timestamp 1704896540
transform 0 1 15242 1 0 14049
box -12 -6 262 112
use L1M1_CDNS_524688791851586  L1M1_CDNS_524688791851586_0
timestamp 1704896540
transform 1 0 15492 0 1 16220
box -12 -6 118 760
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1704896540
transform 0 1 14873 1 0 2214
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1704896540
transform 0 1 12946 1 0 1786
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform 0 1 12946 1 0 350
box 0 0 1 1
use M1M2_CDNS_524688791851589  M1M2_CDNS_524688791851589_0
timestamp 1704896540
transform 1 0 15017 0 1 2691
box 0 0 128 500
use M1M2_CDNS_524688791851590  M1M2_CDNS_524688791851590_0
timestamp 1704896540
transform 1 0 10847 0 1 730
box 0 0 2048 500
use M1M2_CDNS_524688791851591  M1M2_CDNS_524688791851591_0
timestamp 1704896540
transform -1 0 15155 0 1 730
box 0 0 1728 500
use M2M3_CDNS_524688791851587  M2M3_CDNS_524688791851587_0
timestamp 1704896540
transform 1 0 10844 0 1 695
box -5 0 1981 554
use M2M3_CDNS_524688791851588  M2M3_CDNS_524688791851588_0
timestamp 1704896540
transform 1 0 13397 0 1 695
box -5 0 1741 554
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform -1 0 13035 0 1 13088
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform -1 0 10861 0 1 349
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_2
timestamp 1704896540
transform 1 0 15179 0 1 13088
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_3
timestamp 1704896540
transform 1 0 13005 0 1 349
box 0 0 1 1
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_0
timestamp 1704896540
transform 1 0 13087 0 -1 13171
box -50 0 2090 100
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_1
timestamp 1704896540
transform 1 0 10913 0 -1 432
box -50 0 2090 100
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_0
timestamp 1704896540
transform 0 -1 12620 -1 0 16694
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_1
timestamp 1704896540
transform 0 1 12892 -1 0 14608
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_2
timestamp 1704896540
transform 0 1 12892 -1 0 16694
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_3
timestamp 1704896540
transform 0 1 15706 -1 0 16859
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_4
timestamp 1704896540
transform 0 1 15706 -1 0 14401
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_5
timestamp 1704896540
transform 0 1 12892 1 0 14390
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative10_09_6
timestamp 1704896540
transform 0 1 15706 1 0 13947
box -49 -82 1428 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x2  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x2_0
timestamp 1704896540
transform 1 0 10421 0 -1 16963
box -45 1145 2425 3987
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3_0
timestamp 1704896540
transform 1 0 1006 0 -1 16963
box -91 -27 2425 4014
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3_1
timestamp 1704896540
transform 1 0 3348 0 -1 16963
box -91 -27 2425 4014
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3_2
timestamp 1704896540
transform 1 0 5690 0 -1 16963
box -91 -27 2425 4014
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_2x3_3
timestamp 1704896540
transform 1 0 8032 0 -1 16963
box -91 -27 2425 4014
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_4  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_4_0
timestamp 1704896540
transform 0 -1 12892 -1 0 2964
box -269 -87 2265 2199
use sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_4  sky130_fd_io__sio_pudrvr_reg_pu_nhvnative_10_4_1
timestamp 1704896540
transform 0 1 13108 -1 0 2964
box -269 -87 2265 2199
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1704896540
transform -1 0 15170 0 1 14858
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1704896540
transform -1 0 15170 0 -1 14583
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_2
timestamp 1704896540
transform 1 0 15027 0 -1 13014
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_3
timestamp 1704896540
transform 1 0 15027 0 -1 16095
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_4
timestamp 1704896540
transform 1 0 15027 0 1 16415
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851592  sky130_fd_io__tk_em1o_CDNS_524688791851592_0
timestamp 1704896540
transform -1 0 12818 0 1 1786
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851592  sky130_fd_io__tk_em1o_CDNS_524688791851592_1
timestamp 1704896540
transform 1 0 13190 0 1 1786
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851593  sky130_fd_io__tk_em1o_CDNS_524688791851593_0
timestamp 1704896540
transform 0 1 10651 -1 0 16245
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_0
timestamp 1704896540
transform -1 0 15171 0 1 16269
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_1
timestamp 1704896540
transform -1 0 15171 0 -1 13150
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_2
timestamp 1704896540
transform -1 0 15171 0 -1 16241
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_3
timestamp 1704896540
transform 1 0 15040 0 -1 14447
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_4
timestamp 1704896540
transform 1 0 15040 0 1 14994
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851594  sky130_fd_io__tk_em1s_CDNS_524688791851594_0
timestamp 1704896540
transform 0 -1 14861 1 0 14841
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851595  sky130_fd_io__tk_em1s_CDNS_524688791851595_0
timestamp 1704896540
transform -1 0 12818 0 1 1997
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851595  sky130_fd_io__tk_em1s_CDNS_524688791851595_1
timestamp 1704896540
transform 1 0 13190 0 1 1997
box 0 0 1 1
<< labels >>
flabel comment s 15437 12341 15437 12341 0 FreeSans 200 0 0 0 vref_int
flabel comment s 15586 12338 15586 12338 0 FreeSans 200 0 0 0 drvhi_h
flabel comment s 15288 12340 15288 12340 0 FreeSans 200 0 0 0 vref_nng
flabel comment s 14874 12343 14874 12343 0 FreeSans 200 0 0 0 vgnd_io
flabel comment s 13982 13711 13982 13711 0 FreeSans 500 0 0 0 M<3>
flabel comment s 13875 15324 13875 15324 0 FreeSans 500 0 0 0 M<2>
flabel comment s 13963 15811 13963 15811 0 FreeSans 500 0 0 0 M<0>
flabel comment s 11547 15821 11547 15821 0 FreeSans 500 0 0 0 M<1>
<< properties >>
string GDS_END 95585724
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94937402
string path 393.650 6.150 393.650 91.025 255.500 91.025 255.500 71.675 
<< end >>
