magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect -43 3357 9951 6465
rect -43 3087 11273 3357
rect 7547 -53 11273 3087
<< nwell >>
rect -124 6186 10031 6546
rect -124 3367 237 6186
rect 7523 3367 7827 6186
rect -124 3007 7827 3367
rect 7466 227 7827 3007
rect 9671 3437 10031 6186
rect 10431 3898 13597 6479
rect 9671 3133 11353 3437
rect 11049 227 11353 3133
rect 12473 3272 13467 3440
rect 12473 3076 12670 3272
rect 13299 3076 13467 3272
rect 12473 2908 13467 3076
rect 7466 -133 11353 227
<< pwell >>
rect 13949 6662 14125 7362
rect 297 6040 7463 6126
rect 297 3514 383 6040
rect 4809 3514 4975 6040
rect 6535 3514 6621 6040
rect 7377 3514 7463 6040
rect 297 3428 7463 3514
rect 7887 6040 9611 6126
rect 7887 781 7973 6040
rect 9525 3073 9611 6040
rect 9525 2987 10989 3073
rect 7887 695 10079 781
rect 7887 373 7973 695
rect 10903 373 10989 2987
rect 7887 287 10989 373
rect 13667 2758 14125 6662
rect 11413 1370 14125 2758
<< nsubdiff >>
rect 12540 3247 12574 3373
rect 12608 3339 12740 3373
rect 12774 3339 12808 3373
rect 12842 3339 12876 3373
rect 12910 3339 12944 3373
rect 12978 3339 13012 3373
rect 13046 3339 13080 3373
rect 13114 3339 13148 3373
rect 13182 3339 13216 3373
rect 13250 3339 13284 3373
rect 13318 3339 13400 3373
rect 13366 3271 13400 3305
rect 12540 3179 12574 3213
rect 12540 3111 12574 3145
rect 13366 3203 13400 3237
rect 13366 3135 13400 3169
rect 12540 3043 12574 3077
rect 12540 2975 12652 3009
rect 12686 2975 12720 3009
rect 12754 2975 12788 3009
rect 12822 2975 12856 3009
rect 12890 2975 12924 3009
rect 12958 2975 12992 3009
rect 13026 2975 13060 3009
rect 13094 2975 13128 3009
rect 13162 2975 13196 3009
rect 13230 2975 13264 3009
rect 13298 2975 13332 3009
rect 13366 2975 13400 3101
<< mvpsubdiff >>
rect 13975 6636 14099 7336
rect 13693 6602 14099 6636
rect 323 6066 449 6100
rect 483 6066 517 6100
rect 551 6066 585 6100
rect 619 6066 653 6100
rect 687 6066 721 6100
rect 755 6066 789 6100
rect 823 6066 857 6100
rect 891 6066 925 6100
rect 959 6066 993 6100
rect 1027 6066 1061 6100
rect 1095 6066 1129 6100
rect 1163 6066 1197 6100
rect 1231 6066 1265 6100
rect 1299 6066 1333 6100
rect 1367 6066 1401 6100
rect 1435 6066 1469 6100
rect 1503 6066 1537 6100
rect 1571 6066 1605 6100
rect 1639 6066 1673 6100
rect 1707 6066 1741 6100
rect 1775 6066 1809 6100
rect 1843 6066 1877 6100
rect 1911 6066 1945 6100
rect 1979 6066 2013 6100
rect 2047 6066 2081 6100
rect 2115 6066 2149 6100
rect 2183 6066 2217 6100
rect 2251 6066 2285 6100
rect 2319 6066 2353 6100
rect 2387 6066 2421 6100
rect 2455 6066 2489 6100
rect 2523 6066 2557 6100
rect 2591 6066 2625 6100
rect 2659 6066 2693 6100
rect 2727 6066 2761 6100
rect 2795 6066 2829 6100
rect 2863 6066 2897 6100
rect 2931 6066 2965 6100
rect 2999 6066 3033 6100
rect 3067 6066 3101 6100
rect 3135 6066 3169 6100
rect 3203 6066 3237 6100
rect 3271 6066 3305 6100
rect 3339 6066 3373 6100
rect 3407 6066 3441 6100
rect 3475 6066 3509 6100
rect 3543 6066 3577 6100
rect 3611 6066 3645 6100
rect 3679 6066 3713 6100
rect 3747 6066 3781 6100
rect 3815 6066 3849 6100
rect 3883 6066 3917 6100
rect 3951 6066 3985 6100
rect 4019 6066 4053 6100
rect 4087 6066 4121 6100
rect 4155 6066 4189 6100
rect 4223 6066 4257 6100
rect 4291 6066 4325 6100
rect 4359 6066 4393 6100
rect 4427 6066 4461 6100
rect 4495 6066 4529 6100
rect 4563 6066 4597 6100
rect 4631 6066 4665 6100
rect 4699 6066 4733 6100
rect 4767 6066 4801 6100
rect 4835 6066 4989 6100
rect 5023 6066 5057 6100
rect 5091 6066 5125 6100
rect 5159 6066 5193 6100
rect 5227 6066 5261 6100
rect 5295 6066 5329 6100
rect 5363 6066 5397 6100
rect 5431 6066 5465 6100
rect 5499 6066 5533 6100
rect 5567 6066 5601 6100
rect 5635 6066 5669 6100
rect 5703 6066 5737 6100
rect 5771 6066 5805 6100
rect 5839 6066 5873 6100
rect 5907 6066 5941 6100
rect 5975 6066 6009 6100
rect 6043 6066 6077 6100
rect 6111 6066 6145 6100
rect 6179 6066 6213 6100
rect 6247 6066 6281 6100
rect 6315 6066 6349 6100
rect 6383 6066 6417 6100
rect 6451 6066 6485 6100
rect 6519 6066 6553 6100
rect 6587 6066 6621 6100
rect 6655 6066 6689 6100
rect 6723 6066 6757 6100
rect 6791 6066 6825 6100
rect 6859 6066 6893 6100
rect 6927 6066 6961 6100
rect 6995 6066 7029 6100
rect 7063 6066 7097 6100
rect 7131 6066 7165 6100
rect 7199 6066 7233 6100
rect 7267 6066 7301 6100
rect 7335 6066 7369 6100
rect 323 5998 357 6032
rect 323 5930 357 5964
rect 323 5862 357 5896
rect 4835 6032 4915 6066
rect 4835 5998 4949 6032
rect 4835 5970 4915 5998
rect 4869 5964 4915 5970
rect 4869 5936 4949 5964
rect 4835 5930 4949 5936
rect 4835 5902 4915 5930
rect 323 5794 357 5828
rect 4869 5896 4915 5902
rect 4869 5868 4949 5896
rect 4835 5862 4949 5868
rect 4835 5834 4915 5862
rect 323 5726 357 5760
rect 323 5658 357 5692
rect 323 5590 357 5624
rect 323 5522 357 5556
rect 323 5454 357 5488
rect 323 5386 357 5420
rect 323 5318 357 5352
rect 323 5250 357 5284
rect 323 5182 357 5216
rect 323 5114 357 5148
rect 323 5046 357 5080
rect 323 4978 357 5012
rect 323 4910 357 4944
rect 323 4842 357 4876
rect 323 4774 357 4808
rect 323 4706 357 4740
rect 323 4638 357 4672
rect 323 4570 357 4604
rect 323 4502 357 4536
rect 323 4434 357 4468
rect 323 4366 357 4400
rect 323 4298 357 4332
rect 323 4230 357 4264
rect 323 4162 357 4196
rect 323 4094 357 4128
rect 323 4026 357 4060
rect 323 3958 357 3992
rect 323 3890 357 3924
rect 323 3822 357 3856
rect 323 3754 357 3788
rect 4869 5828 4915 5834
rect 4869 5800 4949 5828
rect 4835 5794 4949 5800
rect 4835 5766 4915 5794
rect 4869 5760 4915 5766
rect 4869 5732 4949 5760
rect 4835 5726 4949 5732
rect 4835 5698 4915 5726
rect 4869 5692 4915 5698
rect 4869 5664 4949 5692
rect 4835 5658 4949 5664
rect 4835 5630 4915 5658
rect 4869 5624 4915 5630
rect 4869 5596 4949 5624
rect 4835 5590 4949 5596
rect 4835 5562 4915 5590
rect 4869 5556 4915 5562
rect 4869 5528 4949 5556
rect 4835 5522 4949 5528
rect 4835 5494 4915 5522
rect 4869 5488 4915 5494
rect 4869 5460 4949 5488
rect 4835 5454 4949 5460
rect 4835 5426 4915 5454
rect 4869 5420 4915 5426
rect 4869 5392 4949 5420
rect 4835 5386 4949 5392
rect 4835 5358 4915 5386
rect 4869 5352 4915 5358
rect 4869 5324 4949 5352
rect 4835 5318 4949 5324
rect 4835 5290 4915 5318
rect 4869 5284 4915 5290
rect 4869 5256 4949 5284
rect 4835 5250 4949 5256
rect 4835 5222 4915 5250
rect 4869 5216 4915 5222
rect 4869 5188 4949 5216
rect 4835 5182 4949 5188
rect 4835 5154 4915 5182
rect 4869 5148 4915 5154
rect 4869 5120 4949 5148
rect 4835 5114 4949 5120
rect 4835 5086 4915 5114
rect 4869 5080 4915 5086
rect 4869 5052 4949 5080
rect 4835 5046 4949 5052
rect 4835 5018 4915 5046
rect 4869 5012 4915 5018
rect 4869 4984 4949 5012
rect 4835 4978 4949 4984
rect 4835 4950 4915 4978
rect 4869 4944 4915 4950
rect 4869 4916 4949 4944
rect 4835 4910 4949 4916
rect 4835 4882 4915 4910
rect 4869 4876 4915 4882
rect 4869 4848 4949 4876
rect 4835 4842 4949 4848
rect 4835 4814 4915 4842
rect 4869 4808 4915 4814
rect 4869 4780 4949 4808
rect 4835 4774 4949 4780
rect 4835 4746 4915 4774
rect 4869 4740 4915 4746
rect 4869 4712 4949 4740
rect 4835 4706 4949 4712
rect 4835 4678 4915 4706
rect 4869 4672 4915 4678
rect 4869 4644 4949 4672
rect 4835 4638 4949 4644
rect 4835 4610 4915 4638
rect 4869 4604 4915 4610
rect 4869 4576 4949 4604
rect 4835 4570 4949 4576
rect 4835 4542 4915 4570
rect 4869 4536 4915 4542
rect 4869 4508 4949 4536
rect 4835 4502 4949 4508
rect 4835 4474 4915 4502
rect 4869 4468 4915 4474
rect 4869 4440 4949 4468
rect 4835 4434 4949 4440
rect 4835 4406 4915 4434
rect 4869 4400 4915 4406
rect 4869 4372 4949 4400
rect 4835 4366 4949 4372
rect 4835 4338 4915 4366
rect 4869 4332 4915 4338
rect 4869 4304 4949 4332
rect 4835 4298 4949 4304
rect 4835 4270 4915 4298
rect 4869 4264 4915 4270
rect 4869 4236 4949 4264
rect 4835 4230 4949 4236
rect 4835 4202 4915 4230
rect 4869 4196 4915 4202
rect 4869 4168 4949 4196
rect 4835 4162 4949 4168
rect 4835 4134 4915 4162
rect 4869 4128 4915 4134
rect 4869 4100 4949 4128
rect 4835 4094 4949 4100
rect 4835 4066 4915 4094
rect 4869 4060 4915 4066
rect 4869 4032 4949 4060
rect 4835 4026 4949 4032
rect 4835 3998 4915 4026
rect 4869 3992 4915 3998
rect 4869 3964 4949 3992
rect 4835 3958 4949 3964
rect 4835 3930 4915 3958
rect 4869 3924 4915 3930
rect 4869 3896 4949 3924
rect 4835 3890 4949 3896
rect 4835 3862 4915 3890
rect 4869 3856 4915 3862
rect 4869 3828 4949 3856
rect 4835 3822 4949 3828
rect 4835 3794 4915 3822
rect 4869 3788 4915 3794
rect 4869 3760 4949 3788
rect 4835 3754 4949 3760
rect 323 3686 357 3720
rect 4835 3726 4915 3754
rect 4869 3720 4915 3726
rect 4869 3692 4949 3720
rect 4835 3686 4949 3692
rect 323 3618 357 3652
rect 323 3454 357 3584
rect 4835 3658 4915 3686
rect 4869 3652 4915 3658
rect 4869 3624 4949 3652
rect 4835 3618 4949 3624
rect 4835 3590 4915 3618
rect 4869 3584 4915 3590
rect 4869 3556 4949 3584
rect 4835 3522 4949 3556
rect 4869 3488 4949 3522
rect 6561 5990 6595 6066
rect 6561 5922 6595 5956
rect 6561 5854 6595 5888
rect 6561 5786 6595 5820
rect 6561 5718 6595 5752
rect 6561 5650 6595 5684
rect 6561 5582 6595 5616
rect 6561 5514 6595 5548
rect 6561 5446 6595 5480
rect 6561 5378 6595 5412
rect 6561 5310 6595 5344
rect 6561 5242 6595 5276
rect 6561 5174 6595 5208
rect 6561 5106 6595 5140
rect 6561 5038 6595 5072
rect 6561 4970 6595 5004
rect 6561 4902 6595 4936
rect 6561 4834 6595 4868
rect 6561 4766 6595 4800
rect 6561 4698 6595 4732
rect 6561 4630 6595 4664
rect 6561 4562 6595 4596
rect 6561 4494 6595 4528
rect 6561 4426 6595 4460
rect 6561 4357 6595 4392
rect 6561 4288 6595 4323
rect 6561 4219 6595 4254
rect 6561 4150 6595 4185
rect 6561 4081 6595 4116
rect 6561 4012 6595 4047
rect 6561 3943 6595 3978
rect 6561 3874 6595 3909
rect 7403 5970 7437 6100
rect 7403 5902 7437 5936
rect 7403 5834 7437 5868
rect 7403 5766 7437 5800
rect 7403 5698 7437 5732
rect 7403 5630 7437 5664
rect 7403 5562 7437 5596
rect 7403 5494 7437 5528
rect 7403 5426 7437 5460
rect 7403 5358 7437 5392
rect 7403 5290 7437 5324
rect 7403 5222 7437 5256
rect 7403 5154 7437 5188
rect 7403 5086 7437 5120
rect 7403 5018 7437 5052
rect 7403 4950 7437 4984
rect 7403 4882 7437 4916
rect 7403 4814 7437 4848
rect 7403 4746 7437 4780
rect 7403 4678 7437 4712
rect 7403 4610 7437 4644
rect 7403 4542 7437 4576
rect 7403 4474 7437 4508
rect 7403 4406 7437 4440
rect 7403 4338 7437 4372
rect 7403 4270 7437 4304
rect 7403 4202 7437 4236
rect 7403 4134 7437 4168
rect 7403 4066 7437 4100
rect 7403 3998 7437 4032
rect 7403 3930 7437 3964
rect 6561 3805 6595 3840
rect 6561 3736 6595 3771
rect 7403 3862 7437 3896
rect 7403 3794 7437 3828
rect 6561 3667 6595 3702
rect 6561 3598 6595 3633
rect 6561 3488 6595 3564
rect 7403 3726 7437 3760
rect 7403 3658 7437 3692
rect 7403 3590 7437 3624
rect 7403 3522 7437 3556
rect 391 3454 425 3488
rect 459 3454 493 3488
rect 527 3454 561 3488
rect 595 3454 629 3488
rect 663 3454 697 3488
rect 731 3454 765 3488
rect 799 3454 833 3488
rect 867 3454 901 3488
rect 935 3454 969 3488
rect 1003 3454 1037 3488
rect 1071 3454 1105 3488
rect 1139 3454 1173 3488
rect 1207 3454 1241 3488
rect 1275 3454 1309 3488
rect 1343 3454 1377 3488
rect 1411 3454 1445 3488
rect 1479 3454 1513 3488
rect 1547 3454 1581 3488
rect 1615 3454 1649 3488
rect 1683 3454 1717 3488
rect 1751 3454 1785 3488
rect 1819 3454 1853 3488
rect 1887 3454 1921 3488
rect 1955 3454 1989 3488
rect 2023 3454 2057 3488
rect 2091 3454 2125 3488
rect 2159 3454 2193 3488
rect 2227 3454 2261 3488
rect 2295 3454 2329 3488
rect 2363 3454 2397 3488
rect 2431 3454 2465 3488
rect 2499 3454 2533 3488
rect 2567 3454 2601 3488
rect 2635 3454 2669 3488
rect 2703 3454 2737 3488
rect 2771 3454 2805 3488
rect 2839 3454 2873 3488
rect 2907 3454 2941 3488
rect 2975 3454 3009 3488
rect 3043 3454 3077 3488
rect 3111 3454 3145 3488
rect 3179 3454 3213 3488
rect 3247 3454 3281 3488
rect 3315 3454 3349 3488
rect 3383 3454 3417 3488
rect 3451 3454 3485 3488
rect 3519 3454 3553 3488
rect 3587 3454 3621 3488
rect 3655 3454 3689 3488
rect 3723 3454 3757 3488
rect 3791 3454 3825 3488
rect 3859 3454 3893 3488
rect 3927 3454 3961 3488
rect 3995 3454 4029 3488
rect 4063 3454 4097 3488
rect 4131 3454 4165 3488
rect 4199 3454 4233 3488
rect 4267 3454 4301 3488
rect 4335 3454 4369 3488
rect 4403 3454 4437 3488
rect 4471 3454 4505 3488
rect 4539 3454 4573 3488
rect 4607 3454 4641 3488
rect 4675 3454 4709 3488
rect 4743 3454 4949 3488
rect 4983 3454 5017 3488
rect 5051 3454 5085 3488
rect 5119 3454 5153 3488
rect 5187 3454 5221 3488
rect 5255 3454 5289 3488
rect 5323 3454 5357 3488
rect 5391 3454 5425 3488
rect 5459 3454 5493 3488
rect 5527 3454 5561 3488
rect 5595 3454 5629 3488
rect 5663 3454 5697 3488
rect 5731 3454 5765 3488
rect 5799 3454 5833 3488
rect 5867 3454 5901 3488
rect 5935 3454 5969 3488
rect 6003 3454 6037 3488
rect 6071 3454 6105 3488
rect 6139 3454 6173 3488
rect 6207 3454 6241 3488
rect 6275 3454 6309 3488
rect 6343 3454 6377 3488
rect 6411 3454 6445 3488
rect 6479 3454 6513 3488
rect 6547 3454 6581 3488
rect 6615 3454 6649 3488
rect 6683 3454 6717 3488
rect 6751 3454 6785 3488
rect 6819 3454 6853 3488
rect 6887 3454 6921 3488
rect 6955 3454 6989 3488
rect 7023 3454 7057 3488
rect 7091 3454 7125 3488
rect 7159 3454 7193 3488
rect 7227 3454 7261 3488
rect 7295 3454 7329 3488
rect 7363 3454 7437 3488
rect 7913 6066 7997 6100
rect 8031 6066 8065 6100
rect 8099 6066 8133 6100
rect 8167 6066 8201 6100
rect 8235 6066 8269 6100
rect 8303 6066 8337 6100
rect 8371 6066 8405 6100
rect 8439 6066 8473 6100
rect 8507 6066 8541 6100
rect 8575 6066 8701 6100
rect 8735 6066 8769 6100
rect 8803 6066 8837 6100
rect 8871 6066 8905 6100
rect 8939 6066 8973 6100
rect 9007 6066 9041 6100
rect 9075 6066 9109 6100
rect 9143 6066 9177 6100
rect 9211 6066 9245 6100
rect 9279 6066 9313 6100
rect 9347 6066 9381 6100
rect 9415 6066 9449 6100
rect 9483 6066 9517 6100
rect 7913 5998 7947 6032
rect 7913 5930 7947 5964
rect 9551 6005 9585 6100
rect 7913 5862 7947 5896
rect 7913 5794 7947 5828
rect 7913 5726 7947 5760
rect 7913 5658 7947 5692
rect 7913 5590 7947 5624
rect 7913 5522 7947 5556
rect 7913 5454 7947 5488
rect 7913 5386 7947 5420
rect 9551 5937 9585 5971
rect 9551 5869 9585 5903
rect 9551 5801 9585 5835
rect 9551 5733 9585 5767
rect 9551 5665 9585 5699
rect 9551 5597 9585 5631
rect 9551 5529 9585 5563
rect 9551 5461 9585 5495
rect 7913 5318 7947 5352
rect 9551 5393 9585 5427
rect 7913 5250 7947 5284
rect 7913 5182 7947 5216
rect 7913 5114 7947 5148
rect 7913 5046 7947 5080
rect 7913 4978 7947 5012
rect 7913 4910 7947 4944
rect 7913 4842 7947 4876
rect 7913 4774 7947 4808
rect 7913 4706 7947 4740
rect 7913 4638 7947 4672
rect 7913 4570 7947 4604
rect 7913 4502 7947 4536
rect 7913 4434 7947 4468
rect 7913 4366 7947 4400
rect 9551 5325 9585 5359
rect 9551 5257 9585 5291
rect 9551 5189 9585 5223
rect 9551 5121 9585 5155
rect 9551 5053 9585 5087
rect 9551 4985 9585 5019
rect 9551 4917 9585 4951
rect 9551 4849 9585 4883
rect 9551 4781 9585 4815
rect 9551 4713 9585 4747
rect 9551 4645 9585 4679
rect 9551 4577 9585 4611
rect 9551 4509 9585 4543
rect 9551 4441 9585 4475
rect 7913 4298 7947 4332
rect 7913 4230 7947 4264
rect 9551 4373 9585 4407
rect 9551 4305 9585 4339
rect 7913 4162 7947 4196
rect 7913 4094 7947 4128
rect 7913 4026 7947 4060
rect 7913 3958 7947 3992
rect 9551 4237 9585 4271
rect 9551 4169 9585 4203
rect 9551 4101 9585 4135
rect 9551 4033 9585 4067
rect 9551 3965 9585 3999
rect 7913 3890 7947 3924
rect 7913 3822 7947 3856
rect 7913 3754 7947 3788
rect 7913 3686 7947 3720
rect 7913 3618 7947 3652
rect 9551 3897 9585 3931
rect 9551 3829 9585 3863
rect 9551 3761 9585 3795
rect 9551 3693 9585 3727
rect 9551 3625 9585 3659
rect 7913 3550 7947 3584
rect 7913 3482 7947 3516
rect 9551 3557 9585 3591
rect 9551 3489 9585 3523
rect 7913 3414 7947 3448
rect 7913 3346 7947 3380
rect 9551 3421 9585 3455
rect 7913 3278 7947 3312
rect 7913 3210 7947 3244
rect 9551 3353 9585 3387
rect 9551 3285 9585 3319
rect 9551 3217 9585 3251
rect 7913 3142 7947 3176
rect 7913 3074 7947 3108
rect 7913 3006 7947 3040
rect 9551 3149 9585 3183
rect 9551 3081 9585 3115
rect 9551 3013 9619 3047
rect 9653 3013 9687 3047
rect 9721 3013 9755 3047
rect 9789 3013 9823 3047
rect 9857 3013 9891 3047
rect 9925 3013 9959 3047
rect 9993 3013 10027 3047
rect 10061 3013 10095 3047
rect 10129 3013 10163 3047
rect 10197 3013 10231 3047
rect 10265 3013 10299 3047
rect 10333 3013 10367 3047
rect 10401 3013 10435 3047
rect 10469 3013 10503 3047
rect 10537 3013 10571 3047
rect 10605 3013 10639 3047
rect 10673 3013 10707 3047
rect 10741 3013 10775 3047
rect 10809 3013 10843 3047
rect 10877 3013 10963 3047
rect 7913 2938 7947 2972
rect 7913 2870 7947 2904
rect 10929 2945 10963 2979
rect 10929 2877 10963 2911
rect 7913 2802 7947 2836
rect 7913 2734 7947 2768
rect 7913 2666 7947 2700
rect 7913 2598 7947 2632
rect 7913 2530 7947 2564
rect 7913 2462 7947 2496
rect 7913 2394 7947 2428
rect 7913 2326 7947 2360
rect 7913 2258 7947 2292
rect 7913 2190 7947 2224
rect 7913 2122 7947 2156
rect 7913 2054 7947 2088
rect 7913 1986 7947 2020
rect 7913 1918 7947 1952
rect 7913 1850 7947 1884
rect 7913 1782 7947 1816
rect 7913 1714 7947 1748
rect 7913 1646 7947 1680
rect 7913 1578 7947 1612
rect 7913 1510 7947 1544
rect 7913 1442 7947 1476
rect 7913 1374 7947 1408
rect 7913 1306 7947 1340
rect 7913 1238 7947 1272
rect 7913 1170 7947 1204
rect 7913 1102 7947 1136
rect 7913 1034 7947 1068
rect 7913 966 7947 1000
rect 7913 898 7947 932
rect 7913 830 7947 864
rect 7913 755 7947 796
rect 10929 2809 10963 2843
rect 10929 2741 10963 2775
rect 10929 2673 10963 2707
rect 10929 2605 10963 2639
rect 10929 2537 10963 2571
rect 10929 2469 10963 2503
rect 10929 2401 10963 2435
rect 10929 2333 10963 2367
rect 10929 2265 10963 2299
rect 10929 2197 10963 2231
rect 10929 2129 10963 2163
rect 10929 2061 10963 2095
rect 10929 1993 10963 2027
rect 10929 1925 10963 1959
rect 10929 1857 10963 1891
rect 10929 1789 10963 1823
rect 10929 1721 10963 1755
rect 10929 1653 10963 1687
rect 10929 1585 10963 1619
rect 10929 1517 10963 1551
rect 10929 1449 10963 1483
rect 10929 1381 10963 1415
rect 10929 1313 10963 1347
rect 10929 1245 10963 1279
rect 10929 1177 10963 1211
rect 10929 1109 10963 1143
rect 10929 1041 10963 1075
rect 10929 973 10963 1007
rect 10929 905 10963 939
rect 10929 837 10963 871
rect 7913 721 7937 755
rect 7971 721 8005 755
rect 8039 721 8073 755
rect 8107 721 8141 755
rect 8175 721 8209 755
rect 8243 721 8277 755
rect 8311 721 8345 755
rect 8379 721 8413 755
rect 8447 721 8481 755
rect 8515 721 8549 755
rect 8583 721 8617 755
rect 8651 721 8685 755
rect 8719 721 8753 755
rect 8787 721 8822 755
rect 8856 721 8891 755
rect 8925 721 8960 755
rect 8994 721 9029 755
rect 9063 721 9098 755
rect 9132 721 9167 755
rect 9201 721 9236 755
rect 9270 721 9305 755
rect 9339 721 9374 755
rect 9408 721 9443 755
rect 9477 721 9512 755
rect 9546 721 9581 755
rect 9615 721 9650 755
rect 9684 721 9719 755
rect 9753 721 9788 755
rect 9822 721 9857 755
rect 9891 721 9926 755
rect 9960 721 9995 755
rect 10029 721 10053 755
rect 7913 687 7947 721
rect 7913 619 7947 653
rect 7913 551 7947 585
rect 7913 483 7947 517
rect 7913 415 7947 449
rect 7913 347 7947 381
rect 10929 687 10963 803
rect 10929 619 10963 653
rect 10929 551 10963 585
rect 10929 483 10963 517
rect 10929 415 10963 449
rect 10929 347 10963 381
rect 7913 313 7937 347
rect 7971 313 8006 347
rect 8040 313 8075 347
rect 8109 313 8144 347
rect 8178 313 8213 347
rect 8247 313 8282 347
rect 8316 313 8351 347
rect 8385 313 8420 347
rect 8454 313 8489 347
rect 8523 313 8558 347
rect 8592 313 8627 347
rect 8661 313 8696 347
rect 8730 313 8765 347
rect 8799 313 8834 347
rect 8868 313 8903 347
rect 8937 313 8972 347
rect 9006 313 9041 347
rect 9075 313 9110 347
rect 9144 313 9179 347
rect 9213 313 9248 347
rect 9282 313 9317 347
rect 9351 313 9386 347
rect 9420 313 9455 347
rect 9489 313 9524 347
rect 9558 313 9593 347
rect 9627 313 9662 347
rect 9696 313 9731 347
rect 9765 313 9800 347
rect 9834 313 9869 347
rect 9903 313 9938 347
rect 9972 313 10007 347
rect 10041 313 10076 347
rect 10110 313 10145 347
rect 10179 313 10214 347
rect 10248 313 10283 347
rect 10317 313 10352 347
rect 10386 313 10421 347
rect 10455 313 10490 347
rect 10524 313 10559 347
rect 10593 313 10628 347
rect 10662 313 10697 347
rect 10731 313 10766 347
rect 10800 313 10835 347
rect 10869 313 10905 347
rect 10939 313 10963 347
rect 13693 3032 13709 6602
rect 14083 3032 14099 6602
rect 13693 2997 14099 3032
rect 13693 2963 13709 2997
rect 13743 2963 13777 2997
rect 13811 2963 13845 2997
rect 13879 2963 13913 2997
rect 13947 2963 13981 2997
rect 14015 2963 14049 2997
rect 14083 2963 14099 2997
rect 13693 2928 14099 2963
rect 13693 2894 13709 2928
rect 13743 2894 13777 2928
rect 13811 2894 13845 2928
rect 13879 2894 13913 2928
rect 13947 2894 13981 2928
rect 14015 2894 14049 2928
rect 14083 2894 14099 2928
rect 13693 2859 14099 2894
rect 13693 2825 13709 2859
rect 13743 2825 13777 2859
rect 13811 2825 13845 2859
rect 13879 2825 13913 2859
rect 13947 2825 13981 2859
rect 14015 2825 14049 2859
rect 14083 2825 14099 2859
rect 13693 2790 14099 2825
rect 13693 2756 13709 2790
rect 13743 2756 13777 2790
rect 13811 2756 13845 2790
rect 13879 2756 13913 2790
rect 13947 2756 13981 2790
rect 14015 2756 14049 2790
rect 14083 2756 14099 2790
rect 13693 2732 14099 2756
rect 11439 2695 14099 2732
rect 11439 2661 11476 2695
rect 11510 2661 11546 2695
rect 11580 2661 11616 2695
rect 11650 2661 11686 2695
rect 11720 2661 11756 2695
rect 11790 2661 11826 2695
rect 11860 2661 11896 2695
rect 11930 2661 11966 2695
rect 12000 2661 12036 2695
rect 12070 2661 12106 2695
rect 12140 2661 12176 2695
rect 12210 2661 12246 2695
rect 12280 2661 12316 2695
rect 12350 2661 12385 2695
rect 12419 2661 12454 2695
rect 12488 2661 12523 2695
rect 12557 2661 12592 2695
rect 12626 2661 12661 2695
rect 12695 2661 12730 2695
rect 12764 2661 12799 2695
rect 12833 2661 12868 2695
rect 12902 2661 12937 2695
rect 12971 2661 13006 2695
rect 13040 2661 13075 2695
rect 13109 2661 13144 2695
rect 13178 2661 13213 2695
rect 13247 2661 13282 2695
rect 13316 2661 13351 2695
rect 13385 2661 13420 2695
rect 13454 2661 13489 2695
rect 13523 2661 13558 2695
rect 13592 2661 13627 2695
rect 13661 2661 13696 2695
rect 13730 2661 13765 2695
rect 13799 2661 13834 2695
rect 13868 2661 13903 2695
rect 13937 2661 13972 2695
rect 14006 2661 14041 2695
rect 14075 2661 14099 2695
rect 11439 2627 14099 2661
rect 11439 2593 11476 2627
rect 11510 2593 11546 2627
rect 11580 2593 11616 2627
rect 11650 2593 11686 2627
rect 11720 2593 11756 2627
rect 11790 2593 11826 2627
rect 11860 2593 11896 2627
rect 11930 2593 11966 2627
rect 12000 2593 12036 2627
rect 12070 2593 12106 2627
rect 12140 2593 12176 2627
rect 12210 2593 12246 2627
rect 12280 2593 12316 2627
rect 12350 2593 12385 2627
rect 12419 2593 12454 2627
rect 12488 2593 12523 2627
rect 12557 2593 12592 2627
rect 12626 2593 12661 2627
rect 12695 2593 12730 2627
rect 12764 2593 12799 2627
rect 12833 2593 12868 2627
rect 12902 2593 12937 2627
rect 12971 2593 13006 2627
rect 13040 2593 13075 2627
rect 13109 2593 13144 2627
rect 13178 2593 13213 2627
rect 13247 2593 13282 2627
rect 13316 2593 13351 2627
rect 13385 2593 13420 2627
rect 13454 2593 13489 2627
rect 13523 2593 13558 2627
rect 13592 2593 13627 2627
rect 13661 2593 13696 2627
rect 13730 2593 13765 2627
rect 13799 2593 13834 2627
rect 13868 2593 13903 2627
rect 13937 2593 13972 2627
rect 14006 2593 14041 2627
rect 14075 2593 14099 2627
rect 11439 2559 14099 2593
rect 11439 2525 11476 2559
rect 11510 2525 11546 2559
rect 11580 2525 11616 2559
rect 11650 2525 11686 2559
rect 11720 2525 11756 2559
rect 11790 2525 11826 2559
rect 11860 2525 11896 2559
rect 11930 2525 11966 2559
rect 12000 2525 12036 2559
rect 12070 2525 12106 2559
rect 12140 2525 12176 2559
rect 12210 2525 12246 2559
rect 12280 2525 12316 2559
rect 12350 2525 12385 2559
rect 12419 2525 12454 2559
rect 12488 2525 12523 2559
rect 12557 2525 12592 2559
rect 12626 2525 12661 2559
rect 12695 2525 12730 2559
rect 12764 2525 12799 2559
rect 12833 2525 12868 2559
rect 12902 2525 12937 2559
rect 12971 2525 13006 2559
rect 13040 2525 13075 2559
rect 13109 2525 13144 2559
rect 13178 2525 13213 2559
rect 13247 2525 13282 2559
rect 13316 2525 13351 2559
rect 13385 2525 13420 2559
rect 13454 2525 13489 2559
rect 13523 2525 13558 2559
rect 13592 2525 13627 2559
rect 13661 2525 13696 2559
rect 13730 2525 13765 2559
rect 13799 2525 13834 2559
rect 13868 2525 13903 2559
rect 13937 2525 13972 2559
rect 14006 2525 14041 2559
rect 14075 2525 14099 2559
rect 11439 2491 14099 2525
rect 11439 2457 11476 2491
rect 11510 2457 11546 2491
rect 11580 2457 11616 2491
rect 11650 2457 11686 2491
rect 11720 2457 11756 2491
rect 11790 2457 11826 2491
rect 11860 2457 11896 2491
rect 11930 2457 11966 2491
rect 12000 2457 12036 2491
rect 12070 2457 12106 2491
rect 12140 2457 12176 2491
rect 12210 2457 12246 2491
rect 12280 2457 12316 2491
rect 12350 2457 12385 2491
rect 12419 2457 12454 2491
rect 12488 2457 12523 2491
rect 12557 2457 12592 2491
rect 12626 2457 12661 2491
rect 12695 2457 12730 2491
rect 12764 2457 12799 2491
rect 12833 2457 12868 2491
rect 12902 2457 12937 2491
rect 12971 2457 13006 2491
rect 13040 2457 13075 2491
rect 13109 2457 13144 2491
rect 13178 2457 13213 2491
rect 13247 2457 13282 2491
rect 13316 2457 13351 2491
rect 13385 2457 13420 2491
rect 13454 2457 13489 2491
rect 13523 2457 13558 2491
rect 13592 2457 13627 2491
rect 13661 2457 13696 2491
rect 13730 2457 13765 2491
rect 13799 2457 13834 2491
rect 13868 2457 13903 2491
rect 13937 2457 13972 2491
rect 14006 2457 14041 2491
rect 14075 2457 14099 2491
rect 11439 2423 14099 2457
rect 11439 2389 11476 2423
rect 11510 2389 11546 2423
rect 11580 2389 11616 2423
rect 11650 2389 11686 2423
rect 11720 2389 11756 2423
rect 11790 2389 11826 2423
rect 11860 2389 11896 2423
rect 11930 2389 11966 2423
rect 12000 2389 12036 2423
rect 12070 2389 12106 2423
rect 12140 2389 12176 2423
rect 12210 2389 12246 2423
rect 12280 2389 12316 2423
rect 12350 2389 12385 2423
rect 12419 2389 12454 2423
rect 12488 2389 12523 2423
rect 12557 2389 12592 2423
rect 12626 2389 12661 2423
rect 12695 2389 12730 2423
rect 12764 2389 12799 2423
rect 12833 2389 12868 2423
rect 12902 2389 12937 2423
rect 12971 2389 13006 2423
rect 13040 2389 13075 2423
rect 13109 2389 13144 2423
rect 13178 2389 13213 2423
rect 13247 2389 13282 2423
rect 13316 2389 13351 2423
rect 13385 2389 13420 2423
rect 13454 2389 13489 2423
rect 13523 2389 13558 2423
rect 13592 2389 13627 2423
rect 13661 2389 13696 2423
rect 13730 2389 13765 2423
rect 13799 2389 13834 2423
rect 13868 2389 13903 2423
rect 13937 2389 13972 2423
rect 14006 2389 14041 2423
rect 14075 2389 14099 2423
rect 11439 2355 14099 2389
rect 11439 2321 11476 2355
rect 11510 2321 11546 2355
rect 11580 2321 11616 2355
rect 11650 2321 11686 2355
rect 11720 2321 11756 2355
rect 11790 2321 11826 2355
rect 11860 2321 11896 2355
rect 11930 2321 11966 2355
rect 12000 2321 12036 2355
rect 12070 2321 12106 2355
rect 12140 2321 12176 2355
rect 12210 2321 12246 2355
rect 12280 2321 12316 2355
rect 12350 2321 12385 2355
rect 12419 2321 12454 2355
rect 12488 2321 12523 2355
rect 12557 2321 12592 2355
rect 12626 2321 12661 2355
rect 12695 2321 12730 2355
rect 12764 2321 12799 2355
rect 12833 2321 12868 2355
rect 12902 2321 12937 2355
rect 12971 2321 13006 2355
rect 13040 2321 13075 2355
rect 13109 2321 13144 2355
rect 13178 2321 13213 2355
rect 13247 2321 13282 2355
rect 13316 2321 13351 2355
rect 13385 2321 13420 2355
rect 13454 2321 13489 2355
rect 13523 2321 13558 2355
rect 13592 2321 13627 2355
rect 13661 2321 13696 2355
rect 13730 2321 13765 2355
rect 13799 2321 13834 2355
rect 13868 2321 13903 2355
rect 13937 2321 13972 2355
rect 14006 2321 14041 2355
rect 14075 2321 14099 2355
rect 11439 2287 14099 2321
rect 11439 2253 11476 2287
rect 11510 2253 11546 2287
rect 11580 2253 11616 2287
rect 11650 2253 11686 2287
rect 11720 2253 11756 2287
rect 11790 2253 11826 2287
rect 11860 2253 11896 2287
rect 11930 2253 11966 2287
rect 12000 2253 12036 2287
rect 12070 2253 12106 2287
rect 12140 2253 12176 2287
rect 12210 2253 12246 2287
rect 12280 2253 12316 2287
rect 12350 2253 12385 2287
rect 12419 2253 12454 2287
rect 12488 2253 12523 2287
rect 12557 2253 12592 2287
rect 12626 2253 12661 2287
rect 12695 2253 12730 2287
rect 12764 2253 12799 2287
rect 12833 2253 12868 2287
rect 12902 2253 12937 2287
rect 12971 2253 13006 2287
rect 13040 2253 13075 2287
rect 13109 2253 13144 2287
rect 13178 2253 13213 2287
rect 13247 2253 13282 2287
rect 13316 2253 13351 2287
rect 13385 2253 13420 2287
rect 13454 2253 13489 2287
rect 13523 2253 13558 2287
rect 13592 2253 13627 2287
rect 13661 2253 13696 2287
rect 13730 2253 13765 2287
rect 13799 2253 13834 2287
rect 13868 2253 13903 2287
rect 13937 2253 13972 2287
rect 14006 2253 14041 2287
rect 14075 2253 14099 2287
rect 11439 2219 14099 2253
rect 11439 2185 11476 2219
rect 11510 2185 11546 2219
rect 11580 2185 11616 2219
rect 11650 2185 11686 2219
rect 11720 2185 11756 2219
rect 11790 2185 11826 2219
rect 11860 2185 11896 2219
rect 11930 2185 11966 2219
rect 12000 2185 12036 2219
rect 12070 2185 12106 2219
rect 12140 2185 12176 2219
rect 12210 2185 12246 2219
rect 12280 2185 12316 2219
rect 12350 2185 12385 2219
rect 12419 2185 12454 2219
rect 12488 2185 12523 2219
rect 12557 2185 12592 2219
rect 12626 2185 12661 2219
rect 12695 2185 12730 2219
rect 12764 2185 12799 2219
rect 12833 2185 12868 2219
rect 12902 2185 12937 2219
rect 12971 2185 13006 2219
rect 13040 2185 13075 2219
rect 13109 2185 13144 2219
rect 13178 2185 13213 2219
rect 13247 2185 13282 2219
rect 13316 2185 13351 2219
rect 13385 2185 13420 2219
rect 13454 2185 13489 2219
rect 13523 2185 13558 2219
rect 13592 2185 13627 2219
rect 13661 2185 13696 2219
rect 13730 2185 13765 2219
rect 13799 2185 13834 2219
rect 13868 2185 13903 2219
rect 13937 2185 13972 2219
rect 14006 2185 14041 2219
rect 14075 2185 14099 2219
rect 11439 2151 14099 2185
rect 11439 2117 11476 2151
rect 11510 2117 11546 2151
rect 11580 2117 11616 2151
rect 11650 2117 11686 2151
rect 11720 2117 11756 2151
rect 11790 2117 11826 2151
rect 11860 2117 11896 2151
rect 11930 2117 11966 2151
rect 12000 2117 12036 2151
rect 12070 2117 12106 2151
rect 12140 2117 12176 2151
rect 12210 2117 12246 2151
rect 12280 2117 12316 2151
rect 12350 2117 12385 2151
rect 12419 2117 12454 2151
rect 12488 2117 12523 2151
rect 12557 2117 12592 2151
rect 12626 2117 12661 2151
rect 12695 2117 12730 2151
rect 12764 2117 12799 2151
rect 12833 2117 12868 2151
rect 12902 2117 12937 2151
rect 12971 2117 13006 2151
rect 13040 2117 13075 2151
rect 13109 2117 13144 2151
rect 13178 2117 13213 2151
rect 13247 2117 13282 2151
rect 13316 2117 13351 2151
rect 13385 2117 13420 2151
rect 13454 2117 13489 2151
rect 13523 2117 13558 2151
rect 13592 2117 13627 2151
rect 13661 2117 13696 2151
rect 13730 2117 13765 2151
rect 13799 2117 13834 2151
rect 13868 2117 13903 2151
rect 13937 2117 13972 2151
rect 14006 2117 14041 2151
rect 14075 2117 14099 2151
rect 11439 2083 14099 2117
rect 11439 2049 11476 2083
rect 11510 2049 11546 2083
rect 11580 2049 11616 2083
rect 11650 2049 11686 2083
rect 11720 2049 11756 2083
rect 11790 2049 11826 2083
rect 11860 2049 11896 2083
rect 11930 2049 11966 2083
rect 12000 2049 12036 2083
rect 12070 2049 12106 2083
rect 12140 2049 12176 2083
rect 12210 2049 12246 2083
rect 12280 2049 12316 2083
rect 12350 2049 12385 2083
rect 12419 2049 12454 2083
rect 12488 2049 12523 2083
rect 12557 2049 12592 2083
rect 12626 2049 12661 2083
rect 12695 2049 12730 2083
rect 12764 2049 12799 2083
rect 12833 2049 12868 2083
rect 12902 2049 12937 2083
rect 12971 2049 13006 2083
rect 13040 2049 13075 2083
rect 13109 2049 13144 2083
rect 13178 2049 13213 2083
rect 13247 2049 13282 2083
rect 13316 2049 13351 2083
rect 13385 2049 13420 2083
rect 13454 2049 13489 2083
rect 13523 2049 13558 2083
rect 13592 2049 13627 2083
rect 13661 2049 13696 2083
rect 13730 2049 13765 2083
rect 13799 2049 13834 2083
rect 13868 2049 13903 2083
rect 13937 2049 13972 2083
rect 14006 2049 14041 2083
rect 14075 2049 14099 2083
rect 11439 2015 14099 2049
rect 11439 1981 11476 2015
rect 11510 1981 11546 2015
rect 11580 1981 11616 2015
rect 11650 1981 11686 2015
rect 11720 1981 11756 2015
rect 11790 1981 11826 2015
rect 11860 1981 11896 2015
rect 11930 1981 11966 2015
rect 12000 1981 12036 2015
rect 12070 1981 12106 2015
rect 12140 1981 12176 2015
rect 12210 1981 12246 2015
rect 12280 1981 12316 2015
rect 12350 1981 12385 2015
rect 12419 1981 12454 2015
rect 12488 1981 12523 2015
rect 12557 1981 12592 2015
rect 12626 1981 12661 2015
rect 12695 1981 12730 2015
rect 12764 1981 12799 2015
rect 12833 1981 12868 2015
rect 12902 1981 12937 2015
rect 12971 1981 13006 2015
rect 13040 1981 13075 2015
rect 13109 1981 13144 2015
rect 13178 1981 13213 2015
rect 13247 1981 13282 2015
rect 13316 1981 13351 2015
rect 13385 1981 13420 2015
rect 13454 1981 13489 2015
rect 13523 1981 13558 2015
rect 13592 1981 13627 2015
rect 13661 1981 13696 2015
rect 13730 1981 13765 2015
rect 13799 1981 13834 2015
rect 13868 1981 13903 2015
rect 13937 1981 13972 2015
rect 14006 1981 14041 2015
rect 14075 1981 14099 2015
rect 11439 1947 14099 1981
rect 11439 1913 11476 1947
rect 11510 1913 11546 1947
rect 11580 1913 11616 1947
rect 11650 1913 11686 1947
rect 11720 1913 11756 1947
rect 11790 1913 11826 1947
rect 11860 1913 11896 1947
rect 11930 1913 11966 1947
rect 12000 1913 12036 1947
rect 12070 1913 12106 1947
rect 12140 1913 12176 1947
rect 12210 1913 12246 1947
rect 12280 1913 12316 1947
rect 12350 1913 12385 1947
rect 12419 1913 12454 1947
rect 12488 1913 12523 1947
rect 12557 1913 12592 1947
rect 12626 1913 12661 1947
rect 12695 1913 12730 1947
rect 12764 1913 12799 1947
rect 12833 1913 12868 1947
rect 12902 1913 12937 1947
rect 12971 1913 13006 1947
rect 13040 1913 13075 1947
rect 13109 1913 13144 1947
rect 13178 1913 13213 1947
rect 13247 1913 13282 1947
rect 13316 1913 13351 1947
rect 13385 1913 13420 1947
rect 13454 1913 13489 1947
rect 13523 1913 13558 1947
rect 13592 1913 13627 1947
rect 13661 1913 13696 1947
rect 13730 1913 13765 1947
rect 13799 1913 13834 1947
rect 13868 1913 13903 1947
rect 13937 1913 13972 1947
rect 14006 1913 14041 1947
rect 14075 1913 14099 1947
rect 11439 1879 14099 1913
rect 11439 1845 11476 1879
rect 11510 1845 11546 1879
rect 11580 1845 11616 1879
rect 11650 1845 11686 1879
rect 11720 1845 11756 1879
rect 11790 1845 11826 1879
rect 11860 1845 11896 1879
rect 11930 1845 11966 1879
rect 12000 1845 12036 1879
rect 12070 1845 12106 1879
rect 12140 1845 12176 1879
rect 12210 1845 12246 1879
rect 12280 1845 12316 1879
rect 12350 1845 12385 1879
rect 12419 1845 12454 1879
rect 12488 1845 12523 1879
rect 12557 1845 12592 1879
rect 12626 1845 12661 1879
rect 12695 1845 12730 1879
rect 12764 1845 12799 1879
rect 12833 1845 12868 1879
rect 12902 1845 12937 1879
rect 12971 1845 13006 1879
rect 13040 1845 13075 1879
rect 13109 1845 13144 1879
rect 13178 1845 13213 1879
rect 13247 1845 13282 1879
rect 13316 1845 13351 1879
rect 13385 1845 13420 1879
rect 13454 1845 13489 1879
rect 13523 1845 13558 1879
rect 13592 1845 13627 1879
rect 13661 1845 13696 1879
rect 13730 1845 13765 1879
rect 13799 1845 13834 1879
rect 13868 1845 13903 1879
rect 13937 1845 13972 1879
rect 14006 1845 14041 1879
rect 14075 1845 14099 1879
rect 11439 1811 14099 1845
rect 11439 1777 11476 1811
rect 11510 1777 11546 1811
rect 11580 1777 11616 1811
rect 11650 1777 11686 1811
rect 11720 1777 11756 1811
rect 11790 1777 11826 1811
rect 11860 1777 11896 1811
rect 11930 1777 11966 1811
rect 12000 1777 12036 1811
rect 12070 1777 12106 1811
rect 12140 1777 12176 1811
rect 12210 1777 12246 1811
rect 12280 1777 12316 1811
rect 12350 1777 12385 1811
rect 12419 1777 12454 1811
rect 12488 1777 12523 1811
rect 12557 1777 12592 1811
rect 12626 1777 12661 1811
rect 12695 1777 12730 1811
rect 12764 1777 12799 1811
rect 12833 1777 12868 1811
rect 12902 1777 12937 1811
rect 12971 1777 13006 1811
rect 13040 1777 13075 1811
rect 13109 1777 13144 1811
rect 13178 1777 13213 1811
rect 13247 1777 13282 1811
rect 13316 1777 13351 1811
rect 13385 1777 13420 1811
rect 13454 1777 13489 1811
rect 13523 1777 13558 1811
rect 13592 1777 13627 1811
rect 13661 1777 13696 1811
rect 13730 1777 13765 1811
rect 13799 1777 13834 1811
rect 13868 1777 13903 1811
rect 13937 1777 13972 1811
rect 14006 1777 14041 1811
rect 14075 1777 14099 1811
rect 11439 1743 14099 1777
rect 11439 1709 11476 1743
rect 11510 1709 11546 1743
rect 11580 1709 11616 1743
rect 11650 1709 11686 1743
rect 11720 1709 11756 1743
rect 11790 1709 11826 1743
rect 11860 1709 11896 1743
rect 11930 1709 11966 1743
rect 12000 1709 12036 1743
rect 12070 1709 12106 1743
rect 12140 1709 12176 1743
rect 12210 1709 12246 1743
rect 12280 1709 12316 1743
rect 12350 1709 12385 1743
rect 12419 1709 12454 1743
rect 12488 1709 12523 1743
rect 12557 1709 12592 1743
rect 12626 1709 12661 1743
rect 12695 1709 12730 1743
rect 12764 1709 12799 1743
rect 12833 1709 12868 1743
rect 12902 1709 12937 1743
rect 12971 1709 13006 1743
rect 13040 1709 13075 1743
rect 13109 1709 13144 1743
rect 13178 1709 13213 1743
rect 13247 1709 13282 1743
rect 13316 1709 13351 1743
rect 13385 1709 13420 1743
rect 13454 1709 13489 1743
rect 13523 1709 13558 1743
rect 13592 1709 13627 1743
rect 13661 1709 13696 1743
rect 13730 1709 13765 1743
rect 13799 1709 13834 1743
rect 13868 1709 13903 1743
rect 13937 1709 13972 1743
rect 14006 1709 14041 1743
rect 14075 1709 14099 1743
rect 11439 1675 14099 1709
rect 11439 1641 11476 1675
rect 11510 1641 11546 1675
rect 11580 1641 11616 1675
rect 11650 1641 11686 1675
rect 11720 1641 11756 1675
rect 11790 1641 11826 1675
rect 11860 1641 11896 1675
rect 11930 1641 11966 1675
rect 12000 1641 12036 1675
rect 12070 1641 12106 1675
rect 12140 1641 12176 1675
rect 12210 1641 12246 1675
rect 12280 1641 12316 1675
rect 12350 1641 12385 1675
rect 12419 1641 12454 1675
rect 12488 1641 12523 1675
rect 12557 1641 12592 1675
rect 12626 1641 12661 1675
rect 12695 1641 12730 1675
rect 12764 1641 12799 1675
rect 12833 1641 12868 1675
rect 12902 1641 12937 1675
rect 12971 1641 13006 1675
rect 13040 1641 13075 1675
rect 13109 1641 13144 1675
rect 13178 1641 13213 1675
rect 13247 1641 13282 1675
rect 13316 1641 13351 1675
rect 13385 1641 13420 1675
rect 13454 1641 13489 1675
rect 13523 1641 13558 1675
rect 13592 1641 13627 1675
rect 13661 1641 13696 1675
rect 13730 1641 13765 1675
rect 13799 1641 13834 1675
rect 13868 1641 13903 1675
rect 13937 1641 13972 1675
rect 14006 1641 14041 1675
rect 14075 1641 14099 1675
rect 11439 1566 14099 1641
rect 11439 1532 12957 1566
rect 12991 1532 13030 1566
rect 13064 1532 13103 1566
rect 13137 1532 13176 1566
rect 13210 1532 13249 1566
rect 13283 1532 13321 1566
rect 13355 1532 13393 1566
rect 13427 1532 13465 1566
rect 13499 1532 13537 1566
rect 13571 1532 13609 1566
rect 13643 1532 13681 1566
rect 13715 1532 13753 1566
rect 13787 1532 13825 1566
rect 13859 1532 13897 1566
rect 13931 1532 13969 1566
rect 14003 1532 14041 1566
rect 14075 1532 14099 1566
rect 11439 1498 14099 1532
rect 11439 1464 12957 1498
rect 12991 1464 13030 1498
rect 13064 1464 13103 1498
rect 13137 1464 13176 1498
rect 13210 1464 13249 1498
rect 13283 1464 13321 1498
rect 13355 1464 13393 1498
rect 13427 1464 13465 1498
rect 13499 1464 13537 1498
rect 13571 1464 13609 1498
rect 13643 1464 13681 1498
rect 13715 1464 13753 1498
rect 13787 1464 13825 1498
rect 13859 1464 13897 1498
rect 13931 1464 13969 1498
rect 14003 1464 14041 1498
rect 14075 1464 14099 1498
rect 11439 1430 14099 1464
rect 11439 1396 12957 1430
rect 12991 1396 13030 1430
rect 13064 1396 13103 1430
rect 13137 1396 13176 1430
rect 13210 1396 13249 1430
rect 13283 1396 13321 1430
rect 13355 1396 13393 1430
rect 13427 1396 13465 1430
rect 13499 1396 13537 1430
rect 13571 1396 13609 1430
rect 13643 1396 13681 1430
rect 13715 1396 13753 1430
rect 13787 1396 13825 1430
rect 13859 1396 13897 1430
rect 13931 1396 13969 1430
rect 14003 1396 14041 1430
rect 14075 1396 14099 1430
<< mvnsubdiff >>
rect 0 6389 123 6423
rect 157 6389 191 6423
rect 34 6355 191 6389
rect 102 6321 191 6355
rect 2061 6389 2129 6423
rect 2163 6389 2198 6423
rect 2232 6389 2267 6423
rect 2301 6389 2336 6423
rect 2370 6389 2405 6423
rect 2439 6389 2474 6423
rect 2508 6389 2543 6423
rect 2577 6389 2612 6423
rect 2646 6389 2681 6423
rect 2715 6389 2750 6423
rect 2784 6389 2819 6423
rect 2853 6389 2888 6423
rect 2922 6389 2957 6423
rect 2991 6389 3026 6423
rect 3060 6389 3095 6423
rect 3129 6389 3164 6423
rect 3198 6389 3233 6423
rect 3267 6389 3302 6423
rect 3336 6389 3371 6423
rect 3405 6389 3440 6423
rect 3474 6389 3509 6423
rect 3543 6389 3578 6423
rect 3612 6389 3647 6423
rect 3681 6389 3716 6423
rect 3750 6389 3785 6423
rect 3819 6389 3854 6423
rect 3888 6389 3923 6423
rect 3957 6389 3992 6423
rect 4026 6389 4061 6423
rect 4095 6389 4130 6423
rect 4164 6389 4199 6423
rect 4233 6389 4268 6423
rect 4302 6389 4337 6423
rect 4371 6389 4406 6423
rect 4440 6389 4475 6423
rect 4509 6389 4544 6423
rect 4578 6389 4613 6423
rect 4647 6389 4682 6423
rect 4716 6389 4751 6423
rect 4785 6389 4820 6423
rect 4854 6389 4889 6423
rect 4923 6389 4958 6423
rect 4992 6389 5027 6423
rect 5061 6389 5096 6423
rect 5130 6389 5165 6423
rect 5199 6389 5234 6423
rect 5268 6389 5303 6423
rect 5337 6389 5372 6423
rect 5406 6389 5441 6423
rect 5475 6389 5510 6423
rect 5544 6389 5579 6423
rect 5613 6389 5648 6423
rect 5682 6389 5717 6423
rect 5751 6389 5786 6423
rect 5820 6389 5855 6423
rect 5889 6389 5924 6423
rect 2061 6355 5924 6389
rect 7658 6389 7794 6423
rect 7658 6355 7726 6389
rect 7760 6355 7794 6389
rect 2061 6321 2129 6355
rect 2163 6321 2198 6355
rect 2232 6321 2267 6355
rect 2301 6321 2336 6355
rect 2370 6321 2405 6355
rect 2439 6321 2474 6355
rect 2508 6321 2543 6355
rect 2577 6321 2612 6355
rect 2646 6321 2681 6355
rect 2715 6321 2750 6355
rect 2784 6321 2819 6355
rect 2853 6321 2888 6355
rect 2922 6321 2957 6355
rect 2991 6321 3026 6355
rect 3060 6321 3095 6355
rect 3129 6321 3164 6355
rect 3198 6321 3233 6355
rect 3267 6321 3302 6355
rect 3336 6321 3371 6355
rect 3405 6321 3440 6355
rect 3474 6321 3509 6355
rect 3543 6321 3578 6355
rect 7692 6321 7794 6355
rect 9732 6389 9766 6423
rect 9800 6389 9908 6423
rect 9732 6355 9874 6389
rect 9732 6321 9806 6355
rect 102 6287 259 6321
rect 170 6253 259 6287
rect 2061 6287 3578 6321
rect 2061 6253 2129 6287
rect 2163 6253 2198 6287
rect 2232 6253 2267 6287
rect 2301 6253 2336 6287
rect 2370 6253 2405 6287
rect 2439 6253 2474 6287
rect 2508 6253 2543 6287
rect 2577 6253 2612 6287
rect 2646 6253 2681 6287
rect 2715 6253 2750 6287
rect 2784 6253 2819 6287
rect 2853 6253 2888 6287
rect 2922 6253 2957 6287
rect 2991 6253 3026 6287
rect 3060 6253 3095 6287
rect 3129 6253 3164 6287
rect 3198 6253 3233 6287
rect 3267 6253 3302 6287
rect 3336 6253 3371 6287
rect 3405 6253 3440 6287
rect 3474 6253 3509 6287
rect 3543 6253 3578 6287
rect 7624 6320 7794 6321
rect 7624 6286 7726 6320
rect 7624 6253 7658 6286
rect 7590 6252 7658 6253
rect 7692 6253 7726 6286
rect 9664 6287 9806 6321
rect 9664 6253 9738 6287
rect 7692 6252 7760 6253
rect 7590 6218 7726 6252
rect 7624 6217 7760 6218
rect 7624 6184 7658 6217
rect 7590 6183 7658 6184
rect 7692 6184 7760 6217
rect 7692 6183 7726 6184
rect 7590 6150 7726 6183
rect 7590 6149 7760 6150
rect 7624 6148 7760 6149
rect 7624 6115 7658 6148
rect 7590 6114 7658 6115
rect 7692 6116 7760 6148
rect 7692 6114 7726 6116
rect 7590 6082 7726 6114
rect 7590 6080 7760 6082
rect 7624 6079 7760 6080
rect 7624 6046 7658 6079
rect 7590 6045 7658 6046
rect 7692 6048 7760 6079
rect 7692 6045 7726 6048
rect 7590 6014 7726 6045
rect 7590 6011 7760 6014
rect 7624 6010 7760 6011
rect 7624 5977 7658 6010
rect 7590 5976 7658 5977
rect 7692 5980 7760 6010
rect 7692 5976 7726 5980
rect 7590 5946 7726 5976
rect 7590 5942 7760 5946
rect 7624 5941 7760 5942
rect 7624 5908 7658 5941
rect 7590 5907 7658 5908
rect 7692 5912 7760 5941
rect 7692 5907 7726 5912
rect 7590 5878 7726 5907
rect 7590 5873 7760 5878
rect 7624 5872 7760 5873
rect 7624 5839 7658 5872
rect 7590 5838 7658 5839
rect 7692 5844 7760 5872
rect 7692 5838 7726 5844
rect 7590 5810 7726 5838
rect 7590 5804 7760 5810
rect 7624 5803 7760 5804
rect 7624 5770 7658 5803
rect 7590 5769 7658 5770
rect 7692 5776 7760 5803
rect 7692 5769 7726 5776
rect 7590 5742 7726 5769
rect 7590 5735 7760 5742
rect 7624 5734 7760 5735
rect 7624 5701 7658 5734
rect 7590 5700 7658 5701
rect 7692 5708 7760 5734
rect 7692 5700 7726 5708
rect 7590 5674 7726 5700
rect 7590 5666 7760 5674
rect 7624 5665 7760 5666
rect 7624 5632 7658 5665
rect 7590 5631 7658 5632
rect 7692 5640 7760 5665
rect 7692 5631 7726 5640
rect 7590 5606 7726 5631
rect 7590 5597 7760 5606
rect 7624 5596 7760 5597
rect 7624 5563 7658 5596
rect 7590 5562 7658 5563
rect 7692 5572 7760 5596
rect 7692 5562 7726 5572
rect 7590 5538 7726 5562
rect 7590 5528 7760 5538
rect 7624 5527 7760 5528
rect 7624 5494 7658 5527
rect 7590 5493 7658 5494
rect 7692 5504 7760 5527
rect 7692 5493 7726 5504
rect 7590 5470 7726 5493
rect 7590 5459 7760 5470
rect 7624 5458 7760 5459
rect 7624 5425 7658 5458
rect 7590 5424 7658 5425
rect 7692 5436 7760 5458
rect 7692 5424 7726 5436
rect 7590 5402 7726 5424
rect 7590 5390 7760 5402
rect 7624 5389 7760 5390
rect 7624 5356 7658 5389
rect 7590 5355 7658 5356
rect 7692 5368 7760 5389
rect 7692 5355 7726 5368
rect 7590 5334 7726 5355
rect 7590 5321 7760 5334
rect 7624 5320 7760 5321
rect 7624 5287 7658 5320
rect 7590 5286 7658 5287
rect 7692 5300 7760 5320
rect 7692 5286 7726 5300
rect 7590 5266 7726 5286
rect 7590 5252 7760 5266
rect 7624 5251 7760 5252
rect 7624 5218 7658 5251
rect 7590 5217 7658 5218
rect 7692 5232 7760 5251
rect 7692 5217 7726 5232
rect 7590 5198 7726 5217
rect 7590 5183 7760 5198
rect 7624 5182 7760 5183
rect 7624 5149 7658 5182
rect 7590 5148 7658 5149
rect 7692 5164 7760 5182
rect 7692 5148 7726 5164
rect 7590 5130 7726 5148
rect 7590 5114 7760 5130
rect 7624 5113 7760 5114
rect 7624 5080 7658 5113
rect 7590 5079 7658 5080
rect 7692 5096 7760 5113
rect 7692 5079 7726 5096
rect 7590 5062 7726 5079
rect 7590 5045 7760 5062
rect 7624 5044 7760 5045
rect 7624 5011 7658 5044
rect 7590 5010 7658 5011
rect 7692 5028 7760 5044
rect 7692 5010 7726 5028
rect 7590 4994 7726 5010
rect 7590 4976 7760 4994
rect 7624 4975 7760 4976
rect 7624 4942 7658 4975
rect 7590 4941 7658 4942
rect 7692 4960 7760 4975
rect 7692 4941 7726 4960
rect 7590 4926 7726 4941
rect 7590 4907 7760 4926
rect 7624 4906 7760 4907
rect 7624 4873 7658 4906
rect 7590 4872 7658 4873
rect 7692 4892 7760 4906
rect 7692 4872 7726 4892
rect 7590 4858 7726 4872
rect 7590 4838 7760 4858
rect 7624 4837 7760 4838
rect 7624 4804 7658 4837
rect 7590 4803 7658 4804
rect 7692 4824 7760 4837
rect 7692 4803 7726 4824
rect 7590 4790 7726 4803
rect 7590 4769 7760 4790
rect 7624 4768 7760 4769
rect 7624 4735 7658 4768
rect 7590 4734 7658 4735
rect 7692 4756 7760 4768
rect 7692 4734 7726 4756
rect 7590 4722 7726 4734
rect 7590 4700 7760 4722
rect 7624 4699 7760 4700
rect 7624 4666 7658 4699
rect 7590 4665 7658 4666
rect 7692 4688 7760 4699
rect 7692 4665 7726 4688
rect 7590 4654 7726 4665
rect 7590 4631 7760 4654
rect 7624 4630 7760 4631
rect 7624 4597 7658 4630
rect 7590 4596 7658 4597
rect 7692 4620 7760 4630
rect 7692 4596 7726 4620
rect 7590 4586 7726 4596
rect 7590 4562 7760 4586
rect 7624 4561 7760 4562
rect 7624 4528 7658 4561
rect 7590 4527 7658 4528
rect 7692 4552 7760 4561
rect 7692 4527 7726 4552
rect 7590 4518 7726 4527
rect 7590 4493 7760 4518
rect 7624 4492 7760 4493
rect 7624 4459 7658 4492
rect 7590 4458 7658 4459
rect 7692 4484 7760 4492
rect 7692 4458 7726 4484
rect 7590 4450 7726 4458
rect 7590 4424 7760 4450
rect 7624 4423 7760 4424
rect 7624 4390 7658 4423
rect 7590 4389 7658 4390
rect 7692 4416 7760 4423
rect 7692 4389 7726 4416
rect 7590 4382 7726 4389
rect 7590 4355 7760 4382
rect 7624 4354 7760 4355
rect 7624 4321 7658 4354
rect 7590 4320 7658 4321
rect 7692 4348 7760 4354
rect 7692 4320 7726 4348
rect 7590 4314 7726 4320
rect 7590 4286 7760 4314
rect 7624 4285 7760 4286
rect 7624 4252 7658 4285
rect 7590 4251 7658 4252
rect 7692 4280 7760 4285
rect 7692 4251 7726 4280
rect 7590 4246 7726 4251
rect 7590 4217 7760 4246
rect 7624 4216 7760 4217
rect 7624 4183 7658 4216
rect 7590 4182 7658 4183
rect 7692 4212 7760 4216
rect 7692 4182 7726 4212
rect 7590 4178 7726 4182
rect 7590 4148 7760 4178
rect 7624 4147 7760 4148
rect 7624 4114 7658 4147
rect 7590 4113 7658 4114
rect 7692 4144 7760 4147
rect 7692 4113 7726 4144
rect 7590 4110 7726 4113
rect 7590 4079 7760 4110
rect 7624 4078 7760 4079
rect 7624 4045 7658 4078
rect 7590 4044 7658 4045
rect 7692 4076 7760 4078
rect 7692 4044 7726 4076
rect 7590 4042 7726 4044
rect 7590 4010 7760 4042
rect 7624 4009 7760 4010
rect 7624 3976 7658 4009
rect 7590 3975 7658 3976
rect 7692 4008 7760 4009
rect 7692 3975 7726 4008
rect 7590 3974 7726 3975
rect 7590 3941 7760 3974
rect 7624 3940 7760 3941
rect 7624 3907 7658 3940
rect 7590 3872 7658 3907
rect 0 3261 68 3295
rect 0 3204 170 3261
rect 7590 3204 7760 3498
rect 0 3170 7760 3204
rect 7664 64 7760 3170
rect 10498 6378 10617 6412
rect 10651 6378 10685 6412
rect 10719 6378 10753 6412
rect 10787 6378 10821 6412
rect 10855 6378 10889 6412
rect 10923 6378 10957 6412
rect 10991 6378 11025 6412
rect 11059 6378 11093 6412
rect 11127 6378 11161 6412
rect 11195 6378 11229 6412
rect 11263 6378 11297 6412
rect 11331 6378 11365 6412
rect 11399 6378 11480 6412
rect 11514 6378 11548 6412
rect 11582 6378 11616 6412
rect 11650 6378 11684 6412
rect 11718 6378 11752 6412
rect 11786 6378 11820 6412
rect 11854 6378 11888 6412
rect 11922 6378 11956 6412
rect 11990 6378 12024 6412
rect 12058 6378 12092 6412
rect 12126 6378 12160 6412
rect 12194 6378 12228 6412
rect 12262 6378 12296 6412
rect 12330 6378 12364 6412
rect 12398 6378 12432 6412
rect 12466 6378 12500 6412
rect 12534 6378 12568 6412
rect 12602 6378 12636 6412
rect 12670 6378 12704 6412
rect 12738 6378 12772 6412
rect 12806 6378 12840 6412
rect 12874 6378 12908 6412
rect 12942 6378 12976 6412
rect 13010 6378 13044 6412
rect 13078 6378 13112 6412
rect 13146 6378 13258 6412
rect 13292 6378 13326 6412
rect 13360 6378 13394 6412
rect 13428 6378 13462 6412
rect 10498 6310 10532 6344
rect 13496 6328 13530 6412
rect 10498 6242 10532 6276
rect 13496 6260 13530 6294
rect 10498 6174 10532 6208
rect 10498 6106 10532 6140
rect 10498 6038 10532 6072
rect 10498 5970 10532 6004
rect 10498 5902 10532 5936
rect 10498 5834 10532 5868
rect 10498 5766 10532 5800
rect 10498 5698 10532 5732
rect 10498 5630 10532 5664
rect 10498 5562 10532 5596
rect 10498 5494 10532 5528
rect 13496 6192 13530 6226
rect 13496 6124 13530 6158
rect 13496 6056 13530 6090
rect 13496 5988 13530 6022
rect 13496 5920 13530 5954
rect 13496 5852 13530 5886
rect 13496 5784 13530 5818
rect 13496 5716 13530 5750
rect 13496 5597 13530 5682
rect 13496 5529 13530 5563
rect 10498 5426 10532 5460
rect 13496 5461 13530 5495
rect 10498 5358 10532 5392
rect 10498 5290 10532 5324
rect 10498 5222 10532 5256
rect 10498 5154 10532 5188
rect 10498 5086 10532 5120
rect 10498 5018 10532 5052
rect 10498 4950 10532 4984
rect 10498 4882 10532 4916
rect 10498 4814 10532 4848
rect 13496 5393 13530 5427
rect 13496 5325 13530 5359
rect 13496 5257 13530 5291
rect 13496 5189 13530 5223
rect 13496 5121 13530 5155
rect 13496 5053 13530 5087
rect 13496 4985 13530 5019
rect 13496 4917 13530 4951
rect 13496 4849 13530 4883
rect 10498 4746 10532 4780
rect 13496 4781 13530 4815
rect 10498 4678 10532 4712
rect 10498 4610 10532 4644
rect 10498 4542 10532 4576
rect 10498 4474 10532 4508
rect 10498 4406 10532 4440
rect 10498 4338 10532 4372
rect 10498 4270 10532 4304
rect 10498 4202 10532 4236
rect 10498 4134 10532 4168
rect 10498 3965 10532 4100
rect 13496 4713 13530 4747
rect 13496 4645 13530 4679
rect 13496 4577 13530 4611
rect 13496 4509 13530 4543
rect 13496 4441 13530 4475
rect 13496 4373 13530 4407
rect 13496 4305 13530 4339
rect 13496 4237 13530 4271
rect 13496 4169 13530 4203
rect 13496 4101 13530 4135
rect 13496 4033 13530 4067
rect 10566 3965 10600 3999
rect 10634 3965 10668 3999
rect 10702 3965 10736 3999
rect 10770 3965 10804 3999
rect 10838 3965 10872 3999
rect 10906 3965 10940 3999
rect 10974 3965 11008 3999
rect 11042 3965 11076 3999
rect 11110 3965 11144 3999
rect 11178 3965 11212 3999
rect 11246 3965 11280 3999
rect 11314 3965 11348 3999
rect 11382 3965 11416 3999
rect 11450 3965 11484 3999
rect 11518 3965 11552 3999
rect 11586 3965 11620 3999
rect 11654 3965 11688 3999
rect 11722 3965 11756 3999
rect 11790 3965 11824 3999
rect 11858 3965 11892 3999
rect 11926 3965 11960 3999
rect 11994 3965 12028 3999
rect 12062 3965 12096 3999
rect 12130 3965 12164 3999
rect 12198 3965 12232 3999
rect 12266 3965 12300 3999
rect 12334 3965 12368 3999
rect 12402 3965 12436 3999
rect 12470 3965 12504 3999
rect 12538 3965 12572 3999
rect 12606 3965 12640 3999
rect 12674 3965 12708 3999
rect 12742 3965 12776 3999
rect 12810 3965 12844 3999
rect 12878 3965 12912 3999
rect 12946 3965 12980 3999
rect 13014 3965 13048 3999
rect 13082 3965 13116 3999
rect 13150 3965 13184 3999
rect 13218 3965 13252 3999
rect 13286 3965 13320 3999
rect 13354 3965 13388 3999
rect 13422 3965 13530 3999
rect 11132 3336 11166 3370
rect 11200 3336 11286 3370
rect 11132 3302 11252 3336
rect 9840 3261 9942 3295
rect 11132 3268 11184 3302
rect 9738 3200 9942 3261
rect 11064 3234 11184 3268
rect 11064 3200 11116 3234
rect 11116 106 11252 140
rect 11116 64 11286 106
rect 7664 30 11286 64
<< nsubdiffcont >>
rect 12574 3339 12608 3373
rect 12740 3339 12774 3373
rect 12808 3339 12842 3373
rect 12876 3339 12910 3373
rect 12944 3339 12978 3373
rect 13012 3339 13046 3373
rect 13080 3339 13114 3373
rect 13148 3339 13182 3373
rect 13216 3339 13250 3373
rect 13284 3339 13318 3373
rect 13366 3305 13400 3339
rect 12540 3213 12574 3247
rect 12540 3145 12574 3179
rect 13366 3237 13400 3271
rect 13366 3169 13400 3203
rect 12540 3077 12574 3111
rect 12540 3009 12574 3043
rect 13366 3101 13400 3135
rect 12652 2975 12686 3009
rect 12720 2975 12754 3009
rect 12788 2975 12822 3009
rect 12856 2975 12890 3009
rect 12924 2975 12958 3009
rect 12992 2975 13026 3009
rect 13060 2975 13094 3009
rect 13128 2975 13162 3009
rect 13196 2975 13230 3009
rect 13264 2975 13298 3009
rect 13332 2975 13366 3009
<< mvpsubdiffcont >>
rect 449 6066 483 6100
rect 517 6066 551 6100
rect 585 6066 619 6100
rect 653 6066 687 6100
rect 721 6066 755 6100
rect 789 6066 823 6100
rect 857 6066 891 6100
rect 925 6066 959 6100
rect 993 6066 1027 6100
rect 1061 6066 1095 6100
rect 1129 6066 1163 6100
rect 1197 6066 1231 6100
rect 1265 6066 1299 6100
rect 1333 6066 1367 6100
rect 1401 6066 1435 6100
rect 1469 6066 1503 6100
rect 1537 6066 1571 6100
rect 1605 6066 1639 6100
rect 1673 6066 1707 6100
rect 1741 6066 1775 6100
rect 1809 6066 1843 6100
rect 1877 6066 1911 6100
rect 1945 6066 1979 6100
rect 2013 6066 2047 6100
rect 2081 6066 2115 6100
rect 2149 6066 2183 6100
rect 2217 6066 2251 6100
rect 2285 6066 2319 6100
rect 2353 6066 2387 6100
rect 2421 6066 2455 6100
rect 2489 6066 2523 6100
rect 2557 6066 2591 6100
rect 2625 6066 2659 6100
rect 2693 6066 2727 6100
rect 2761 6066 2795 6100
rect 2829 6066 2863 6100
rect 2897 6066 2931 6100
rect 2965 6066 2999 6100
rect 3033 6066 3067 6100
rect 3101 6066 3135 6100
rect 3169 6066 3203 6100
rect 3237 6066 3271 6100
rect 3305 6066 3339 6100
rect 3373 6066 3407 6100
rect 3441 6066 3475 6100
rect 3509 6066 3543 6100
rect 3577 6066 3611 6100
rect 3645 6066 3679 6100
rect 3713 6066 3747 6100
rect 3781 6066 3815 6100
rect 3849 6066 3883 6100
rect 3917 6066 3951 6100
rect 3985 6066 4019 6100
rect 4053 6066 4087 6100
rect 4121 6066 4155 6100
rect 4189 6066 4223 6100
rect 4257 6066 4291 6100
rect 4325 6066 4359 6100
rect 4393 6066 4427 6100
rect 4461 6066 4495 6100
rect 4529 6066 4563 6100
rect 4597 6066 4631 6100
rect 4665 6066 4699 6100
rect 4733 6066 4767 6100
rect 4801 6066 4835 6100
rect 4989 6066 5023 6100
rect 5057 6066 5091 6100
rect 5125 6066 5159 6100
rect 5193 6066 5227 6100
rect 5261 6066 5295 6100
rect 5329 6066 5363 6100
rect 5397 6066 5431 6100
rect 5465 6066 5499 6100
rect 5533 6066 5567 6100
rect 5601 6066 5635 6100
rect 5669 6066 5703 6100
rect 5737 6066 5771 6100
rect 5805 6066 5839 6100
rect 5873 6066 5907 6100
rect 5941 6066 5975 6100
rect 6009 6066 6043 6100
rect 6077 6066 6111 6100
rect 6145 6066 6179 6100
rect 6213 6066 6247 6100
rect 6281 6066 6315 6100
rect 6349 6066 6383 6100
rect 6417 6066 6451 6100
rect 6485 6066 6519 6100
rect 6553 6066 6587 6100
rect 6621 6066 6655 6100
rect 6689 6066 6723 6100
rect 6757 6066 6791 6100
rect 6825 6066 6859 6100
rect 6893 6066 6927 6100
rect 6961 6066 6995 6100
rect 7029 6066 7063 6100
rect 7097 6066 7131 6100
rect 7165 6066 7199 6100
rect 7233 6066 7267 6100
rect 7301 6066 7335 6100
rect 7369 6066 7403 6100
rect 323 6032 357 6066
rect 323 5964 357 5998
rect 323 5896 357 5930
rect 4915 6032 4949 6066
rect 4835 5936 4869 5970
rect 4915 5964 4949 5998
rect 323 5828 357 5862
rect 4835 5868 4869 5902
rect 4915 5896 4949 5930
rect 323 5760 357 5794
rect 323 5692 357 5726
rect 323 5624 357 5658
rect 323 5556 357 5590
rect 323 5488 357 5522
rect 323 5420 357 5454
rect 323 5352 357 5386
rect 323 5284 357 5318
rect 323 5216 357 5250
rect 323 5148 357 5182
rect 323 5080 357 5114
rect 323 5012 357 5046
rect 323 4944 357 4978
rect 323 4876 357 4910
rect 323 4808 357 4842
rect 323 4740 357 4774
rect 323 4672 357 4706
rect 323 4604 357 4638
rect 323 4536 357 4570
rect 323 4468 357 4502
rect 323 4400 357 4434
rect 323 4332 357 4366
rect 323 4264 357 4298
rect 323 4196 357 4230
rect 323 4128 357 4162
rect 323 4060 357 4094
rect 323 3992 357 4026
rect 323 3924 357 3958
rect 323 3856 357 3890
rect 323 3788 357 3822
rect 323 3720 357 3754
rect 4835 5800 4869 5834
rect 4915 5828 4949 5862
rect 4835 5732 4869 5766
rect 4915 5760 4949 5794
rect 4835 5664 4869 5698
rect 4915 5692 4949 5726
rect 4835 5596 4869 5630
rect 4915 5624 4949 5658
rect 4835 5528 4869 5562
rect 4915 5556 4949 5590
rect 4835 5460 4869 5494
rect 4915 5488 4949 5522
rect 4835 5392 4869 5426
rect 4915 5420 4949 5454
rect 4835 5324 4869 5358
rect 4915 5352 4949 5386
rect 4835 5256 4869 5290
rect 4915 5284 4949 5318
rect 4835 5188 4869 5222
rect 4915 5216 4949 5250
rect 4835 5120 4869 5154
rect 4915 5148 4949 5182
rect 4835 5052 4869 5086
rect 4915 5080 4949 5114
rect 4835 4984 4869 5018
rect 4915 5012 4949 5046
rect 4835 4916 4869 4950
rect 4915 4944 4949 4978
rect 4835 4848 4869 4882
rect 4915 4876 4949 4910
rect 4835 4780 4869 4814
rect 4915 4808 4949 4842
rect 4835 4712 4869 4746
rect 4915 4740 4949 4774
rect 4835 4644 4869 4678
rect 4915 4672 4949 4706
rect 4835 4576 4869 4610
rect 4915 4604 4949 4638
rect 4835 4508 4869 4542
rect 4915 4536 4949 4570
rect 4835 4440 4869 4474
rect 4915 4468 4949 4502
rect 4835 4372 4869 4406
rect 4915 4400 4949 4434
rect 4835 4304 4869 4338
rect 4915 4332 4949 4366
rect 4835 4236 4869 4270
rect 4915 4264 4949 4298
rect 4835 4168 4869 4202
rect 4915 4196 4949 4230
rect 4835 4100 4869 4134
rect 4915 4128 4949 4162
rect 4835 4032 4869 4066
rect 4915 4060 4949 4094
rect 4835 3964 4869 3998
rect 4915 3992 4949 4026
rect 4835 3896 4869 3930
rect 4915 3924 4949 3958
rect 4835 3828 4869 3862
rect 4915 3856 4949 3890
rect 4835 3760 4869 3794
rect 4915 3788 4949 3822
rect 323 3652 357 3686
rect 4835 3692 4869 3726
rect 4915 3720 4949 3754
rect 323 3584 357 3618
rect 4835 3624 4869 3658
rect 4915 3652 4949 3686
rect 4835 3556 4869 3590
rect 4915 3584 4949 3618
rect 4835 3488 4869 3522
rect 6561 5956 6595 5990
rect 6561 5888 6595 5922
rect 6561 5820 6595 5854
rect 6561 5752 6595 5786
rect 6561 5684 6595 5718
rect 6561 5616 6595 5650
rect 6561 5548 6595 5582
rect 6561 5480 6595 5514
rect 6561 5412 6595 5446
rect 6561 5344 6595 5378
rect 6561 5276 6595 5310
rect 6561 5208 6595 5242
rect 6561 5140 6595 5174
rect 6561 5072 6595 5106
rect 6561 5004 6595 5038
rect 6561 4936 6595 4970
rect 6561 4868 6595 4902
rect 6561 4800 6595 4834
rect 6561 4732 6595 4766
rect 6561 4664 6595 4698
rect 6561 4596 6595 4630
rect 6561 4528 6595 4562
rect 6561 4460 6595 4494
rect 6561 4392 6595 4426
rect 6561 4323 6595 4357
rect 6561 4254 6595 4288
rect 6561 4185 6595 4219
rect 6561 4116 6595 4150
rect 6561 4047 6595 4081
rect 6561 3978 6595 4012
rect 6561 3909 6595 3943
rect 6561 3840 6595 3874
rect 7403 5936 7437 5970
rect 7403 5868 7437 5902
rect 7403 5800 7437 5834
rect 7403 5732 7437 5766
rect 7403 5664 7437 5698
rect 7403 5596 7437 5630
rect 7403 5528 7437 5562
rect 7403 5460 7437 5494
rect 7403 5392 7437 5426
rect 7403 5324 7437 5358
rect 7403 5256 7437 5290
rect 7403 5188 7437 5222
rect 7403 5120 7437 5154
rect 7403 5052 7437 5086
rect 7403 4984 7437 5018
rect 7403 4916 7437 4950
rect 7403 4848 7437 4882
rect 7403 4780 7437 4814
rect 7403 4712 7437 4746
rect 7403 4644 7437 4678
rect 7403 4576 7437 4610
rect 7403 4508 7437 4542
rect 7403 4440 7437 4474
rect 7403 4372 7437 4406
rect 7403 4304 7437 4338
rect 7403 4236 7437 4270
rect 7403 4168 7437 4202
rect 7403 4100 7437 4134
rect 7403 4032 7437 4066
rect 7403 3964 7437 3998
rect 7403 3896 7437 3930
rect 6561 3771 6595 3805
rect 7403 3828 7437 3862
rect 6561 3702 6595 3736
rect 6561 3633 6595 3667
rect 6561 3564 6595 3598
rect 7403 3760 7437 3794
rect 7403 3692 7437 3726
rect 7403 3624 7437 3658
rect 7403 3556 7437 3590
rect 7403 3488 7437 3522
rect 357 3454 391 3488
rect 425 3454 459 3488
rect 493 3454 527 3488
rect 561 3454 595 3488
rect 629 3454 663 3488
rect 697 3454 731 3488
rect 765 3454 799 3488
rect 833 3454 867 3488
rect 901 3454 935 3488
rect 969 3454 1003 3488
rect 1037 3454 1071 3488
rect 1105 3454 1139 3488
rect 1173 3454 1207 3488
rect 1241 3454 1275 3488
rect 1309 3454 1343 3488
rect 1377 3454 1411 3488
rect 1445 3454 1479 3488
rect 1513 3454 1547 3488
rect 1581 3454 1615 3488
rect 1649 3454 1683 3488
rect 1717 3454 1751 3488
rect 1785 3454 1819 3488
rect 1853 3454 1887 3488
rect 1921 3454 1955 3488
rect 1989 3454 2023 3488
rect 2057 3454 2091 3488
rect 2125 3454 2159 3488
rect 2193 3454 2227 3488
rect 2261 3454 2295 3488
rect 2329 3454 2363 3488
rect 2397 3454 2431 3488
rect 2465 3454 2499 3488
rect 2533 3454 2567 3488
rect 2601 3454 2635 3488
rect 2669 3454 2703 3488
rect 2737 3454 2771 3488
rect 2805 3454 2839 3488
rect 2873 3454 2907 3488
rect 2941 3454 2975 3488
rect 3009 3454 3043 3488
rect 3077 3454 3111 3488
rect 3145 3454 3179 3488
rect 3213 3454 3247 3488
rect 3281 3454 3315 3488
rect 3349 3454 3383 3488
rect 3417 3454 3451 3488
rect 3485 3454 3519 3488
rect 3553 3454 3587 3488
rect 3621 3454 3655 3488
rect 3689 3454 3723 3488
rect 3757 3454 3791 3488
rect 3825 3454 3859 3488
rect 3893 3454 3927 3488
rect 3961 3454 3995 3488
rect 4029 3454 4063 3488
rect 4097 3454 4131 3488
rect 4165 3454 4199 3488
rect 4233 3454 4267 3488
rect 4301 3454 4335 3488
rect 4369 3454 4403 3488
rect 4437 3454 4471 3488
rect 4505 3454 4539 3488
rect 4573 3454 4607 3488
rect 4641 3454 4675 3488
rect 4709 3454 4743 3488
rect 4949 3454 4983 3488
rect 5017 3454 5051 3488
rect 5085 3454 5119 3488
rect 5153 3454 5187 3488
rect 5221 3454 5255 3488
rect 5289 3454 5323 3488
rect 5357 3454 5391 3488
rect 5425 3454 5459 3488
rect 5493 3454 5527 3488
rect 5561 3454 5595 3488
rect 5629 3454 5663 3488
rect 5697 3454 5731 3488
rect 5765 3454 5799 3488
rect 5833 3454 5867 3488
rect 5901 3454 5935 3488
rect 5969 3454 6003 3488
rect 6037 3454 6071 3488
rect 6105 3454 6139 3488
rect 6173 3454 6207 3488
rect 6241 3454 6275 3488
rect 6309 3454 6343 3488
rect 6377 3454 6411 3488
rect 6445 3454 6479 3488
rect 6513 3454 6547 3488
rect 6581 3454 6615 3488
rect 6649 3454 6683 3488
rect 6717 3454 6751 3488
rect 6785 3454 6819 3488
rect 6853 3454 6887 3488
rect 6921 3454 6955 3488
rect 6989 3454 7023 3488
rect 7057 3454 7091 3488
rect 7125 3454 7159 3488
rect 7193 3454 7227 3488
rect 7261 3454 7295 3488
rect 7329 3454 7363 3488
rect 7997 6066 8031 6100
rect 8065 6066 8099 6100
rect 8133 6066 8167 6100
rect 8201 6066 8235 6100
rect 8269 6066 8303 6100
rect 8337 6066 8371 6100
rect 8405 6066 8439 6100
rect 8473 6066 8507 6100
rect 8541 6066 8575 6100
rect 8701 6066 8735 6100
rect 8769 6066 8803 6100
rect 8837 6066 8871 6100
rect 8905 6066 8939 6100
rect 8973 6066 9007 6100
rect 9041 6066 9075 6100
rect 9109 6066 9143 6100
rect 9177 6066 9211 6100
rect 9245 6066 9279 6100
rect 9313 6066 9347 6100
rect 9381 6066 9415 6100
rect 9449 6066 9483 6100
rect 9517 6066 9551 6100
rect 7913 6032 7947 6066
rect 7913 5964 7947 5998
rect 9551 5971 9585 6005
rect 7913 5896 7947 5930
rect 7913 5828 7947 5862
rect 7913 5760 7947 5794
rect 7913 5692 7947 5726
rect 7913 5624 7947 5658
rect 7913 5556 7947 5590
rect 7913 5488 7947 5522
rect 7913 5420 7947 5454
rect 9551 5903 9585 5937
rect 9551 5835 9585 5869
rect 9551 5767 9585 5801
rect 9551 5699 9585 5733
rect 9551 5631 9585 5665
rect 9551 5563 9585 5597
rect 9551 5495 9585 5529
rect 9551 5427 9585 5461
rect 7913 5352 7947 5386
rect 9551 5359 9585 5393
rect 7913 5284 7947 5318
rect 7913 5216 7947 5250
rect 7913 5148 7947 5182
rect 7913 5080 7947 5114
rect 7913 5012 7947 5046
rect 7913 4944 7947 4978
rect 7913 4876 7947 4910
rect 7913 4808 7947 4842
rect 7913 4740 7947 4774
rect 7913 4672 7947 4706
rect 7913 4604 7947 4638
rect 7913 4536 7947 4570
rect 7913 4468 7947 4502
rect 7913 4400 7947 4434
rect 9551 5291 9585 5325
rect 9551 5223 9585 5257
rect 9551 5155 9585 5189
rect 9551 5087 9585 5121
rect 9551 5019 9585 5053
rect 9551 4951 9585 4985
rect 9551 4883 9585 4917
rect 9551 4815 9585 4849
rect 9551 4747 9585 4781
rect 9551 4679 9585 4713
rect 9551 4611 9585 4645
rect 9551 4543 9585 4577
rect 9551 4475 9585 4509
rect 9551 4407 9585 4441
rect 7913 4332 7947 4366
rect 7913 4264 7947 4298
rect 9551 4339 9585 4373
rect 9551 4271 9585 4305
rect 7913 4196 7947 4230
rect 7913 4128 7947 4162
rect 7913 4060 7947 4094
rect 7913 3992 7947 4026
rect 7913 3924 7947 3958
rect 9551 4203 9585 4237
rect 9551 4135 9585 4169
rect 9551 4067 9585 4101
rect 9551 3999 9585 4033
rect 9551 3931 9585 3965
rect 7913 3856 7947 3890
rect 7913 3788 7947 3822
rect 7913 3720 7947 3754
rect 7913 3652 7947 3686
rect 7913 3584 7947 3618
rect 9551 3863 9585 3897
rect 9551 3795 9585 3829
rect 9551 3727 9585 3761
rect 9551 3659 9585 3693
rect 7913 3516 7947 3550
rect 7913 3448 7947 3482
rect 9551 3591 9585 3625
rect 9551 3523 9585 3557
rect 7913 3380 7947 3414
rect 9551 3455 9585 3489
rect 9551 3387 9585 3421
rect 7913 3312 7947 3346
rect 7913 3244 7947 3278
rect 7913 3176 7947 3210
rect 9551 3319 9585 3353
rect 9551 3251 9585 3285
rect 7913 3108 7947 3142
rect 7913 3040 7947 3074
rect 9551 3183 9585 3217
rect 9551 3115 9585 3149
rect 9551 3047 9585 3081
rect 9619 3013 9653 3047
rect 9687 3013 9721 3047
rect 9755 3013 9789 3047
rect 9823 3013 9857 3047
rect 9891 3013 9925 3047
rect 9959 3013 9993 3047
rect 10027 3013 10061 3047
rect 10095 3013 10129 3047
rect 10163 3013 10197 3047
rect 10231 3013 10265 3047
rect 10299 3013 10333 3047
rect 10367 3013 10401 3047
rect 10435 3013 10469 3047
rect 10503 3013 10537 3047
rect 10571 3013 10605 3047
rect 10639 3013 10673 3047
rect 10707 3013 10741 3047
rect 10775 3013 10809 3047
rect 10843 3013 10877 3047
rect 7913 2972 7947 3006
rect 7913 2904 7947 2938
rect 7913 2836 7947 2870
rect 10929 2979 10963 3013
rect 10929 2911 10963 2945
rect 7913 2768 7947 2802
rect 7913 2700 7947 2734
rect 7913 2632 7947 2666
rect 7913 2564 7947 2598
rect 7913 2496 7947 2530
rect 7913 2428 7947 2462
rect 7913 2360 7947 2394
rect 7913 2292 7947 2326
rect 7913 2224 7947 2258
rect 7913 2156 7947 2190
rect 7913 2088 7947 2122
rect 7913 2020 7947 2054
rect 7913 1952 7947 1986
rect 7913 1884 7947 1918
rect 7913 1816 7947 1850
rect 7913 1748 7947 1782
rect 7913 1680 7947 1714
rect 7913 1612 7947 1646
rect 7913 1544 7947 1578
rect 7913 1476 7947 1510
rect 7913 1408 7947 1442
rect 7913 1340 7947 1374
rect 7913 1272 7947 1306
rect 7913 1204 7947 1238
rect 7913 1136 7947 1170
rect 7913 1068 7947 1102
rect 7913 1000 7947 1034
rect 7913 932 7947 966
rect 7913 864 7947 898
rect 7913 796 7947 830
rect 10929 2843 10963 2877
rect 10929 2775 10963 2809
rect 10929 2707 10963 2741
rect 10929 2639 10963 2673
rect 10929 2571 10963 2605
rect 10929 2503 10963 2537
rect 10929 2435 10963 2469
rect 10929 2367 10963 2401
rect 10929 2299 10963 2333
rect 10929 2231 10963 2265
rect 10929 2163 10963 2197
rect 10929 2095 10963 2129
rect 10929 2027 10963 2061
rect 10929 1959 10963 1993
rect 10929 1891 10963 1925
rect 10929 1823 10963 1857
rect 10929 1755 10963 1789
rect 10929 1687 10963 1721
rect 10929 1619 10963 1653
rect 10929 1551 10963 1585
rect 10929 1483 10963 1517
rect 10929 1415 10963 1449
rect 10929 1347 10963 1381
rect 10929 1279 10963 1313
rect 10929 1211 10963 1245
rect 10929 1143 10963 1177
rect 10929 1075 10963 1109
rect 10929 1007 10963 1041
rect 10929 939 10963 973
rect 10929 871 10963 905
rect 10929 803 10963 837
rect 7937 721 7971 755
rect 8005 721 8039 755
rect 8073 721 8107 755
rect 8141 721 8175 755
rect 8209 721 8243 755
rect 8277 721 8311 755
rect 8345 721 8379 755
rect 8413 721 8447 755
rect 8481 721 8515 755
rect 8549 721 8583 755
rect 8617 721 8651 755
rect 8685 721 8719 755
rect 8753 721 8787 755
rect 8822 721 8856 755
rect 8891 721 8925 755
rect 8960 721 8994 755
rect 9029 721 9063 755
rect 9098 721 9132 755
rect 9167 721 9201 755
rect 9236 721 9270 755
rect 9305 721 9339 755
rect 9374 721 9408 755
rect 9443 721 9477 755
rect 9512 721 9546 755
rect 9581 721 9615 755
rect 9650 721 9684 755
rect 9719 721 9753 755
rect 9788 721 9822 755
rect 9857 721 9891 755
rect 9926 721 9960 755
rect 9995 721 10029 755
rect 7913 653 7947 687
rect 7913 585 7947 619
rect 7913 517 7947 551
rect 7913 449 7947 483
rect 7913 381 7947 415
rect 10929 653 10963 687
rect 10929 585 10963 619
rect 10929 517 10963 551
rect 10929 449 10963 483
rect 10929 381 10963 415
rect 7937 313 7971 347
rect 8006 313 8040 347
rect 8075 313 8109 347
rect 8144 313 8178 347
rect 8213 313 8247 347
rect 8282 313 8316 347
rect 8351 313 8385 347
rect 8420 313 8454 347
rect 8489 313 8523 347
rect 8558 313 8592 347
rect 8627 313 8661 347
rect 8696 313 8730 347
rect 8765 313 8799 347
rect 8834 313 8868 347
rect 8903 313 8937 347
rect 8972 313 9006 347
rect 9041 313 9075 347
rect 9110 313 9144 347
rect 9179 313 9213 347
rect 9248 313 9282 347
rect 9317 313 9351 347
rect 9386 313 9420 347
rect 9455 313 9489 347
rect 9524 313 9558 347
rect 9593 313 9627 347
rect 9662 313 9696 347
rect 9731 313 9765 347
rect 9800 313 9834 347
rect 9869 313 9903 347
rect 9938 313 9972 347
rect 10007 313 10041 347
rect 10076 313 10110 347
rect 10145 313 10179 347
rect 10214 313 10248 347
rect 10283 313 10317 347
rect 10352 313 10386 347
rect 10421 313 10455 347
rect 10490 313 10524 347
rect 10559 313 10593 347
rect 10628 313 10662 347
rect 10697 313 10731 347
rect 10766 313 10800 347
rect 10835 313 10869 347
rect 10905 313 10939 347
rect 13709 3032 14083 6602
rect 13709 2963 13743 2997
rect 13777 2963 13811 2997
rect 13845 2963 13879 2997
rect 13913 2963 13947 2997
rect 13981 2963 14015 2997
rect 14049 2963 14083 2997
rect 13709 2894 13743 2928
rect 13777 2894 13811 2928
rect 13845 2894 13879 2928
rect 13913 2894 13947 2928
rect 13981 2894 14015 2928
rect 14049 2894 14083 2928
rect 13709 2825 13743 2859
rect 13777 2825 13811 2859
rect 13845 2825 13879 2859
rect 13913 2825 13947 2859
rect 13981 2825 14015 2859
rect 14049 2825 14083 2859
rect 13709 2756 13743 2790
rect 13777 2756 13811 2790
rect 13845 2756 13879 2790
rect 13913 2756 13947 2790
rect 13981 2756 14015 2790
rect 14049 2756 14083 2790
rect 11476 2661 11510 2695
rect 11546 2661 11580 2695
rect 11616 2661 11650 2695
rect 11686 2661 11720 2695
rect 11756 2661 11790 2695
rect 11826 2661 11860 2695
rect 11896 2661 11930 2695
rect 11966 2661 12000 2695
rect 12036 2661 12070 2695
rect 12106 2661 12140 2695
rect 12176 2661 12210 2695
rect 12246 2661 12280 2695
rect 12316 2661 12350 2695
rect 12385 2661 12419 2695
rect 12454 2661 12488 2695
rect 12523 2661 12557 2695
rect 12592 2661 12626 2695
rect 12661 2661 12695 2695
rect 12730 2661 12764 2695
rect 12799 2661 12833 2695
rect 12868 2661 12902 2695
rect 12937 2661 12971 2695
rect 13006 2661 13040 2695
rect 13075 2661 13109 2695
rect 13144 2661 13178 2695
rect 13213 2661 13247 2695
rect 13282 2661 13316 2695
rect 13351 2661 13385 2695
rect 13420 2661 13454 2695
rect 13489 2661 13523 2695
rect 13558 2661 13592 2695
rect 13627 2661 13661 2695
rect 13696 2661 13730 2695
rect 13765 2661 13799 2695
rect 13834 2661 13868 2695
rect 13903 2661 13937 2695
rect 13972 2661 14006 2695
rect 14041 2661 14075 2695
rect 11476 2593 11510 2627
rect 11546 2593 11580 2627
rect 11616 2593 11650 2627
rect 11686 2593 11720 2627
rect 11756 2593 11790 2627
rect 11826 2593 11860 2627
rect 11896 2593 11930 2627
rect 11966 2593 12000 2627
rect 12036 2593 12070 2627
rect 12106 2593 12140 2627
rect 12176 2593 12210 2627
rect 12246 2593 12280 2627
rect 12316 2593 12350 2627
rect 12385 2593 12419 2627
rect 12454 2593 12488 2627
rect 12523 2593 12557 2627
rect 12592 2593 12626 2627
rect 12661 2593 12695 2627
rect 12730 2593 12764 2627
rect 12799 2593 12833 2627
rect 12868 2593 12902 2627
rect 12937 2593 12971 2627
rect 13006 2593 13040 2627
rect 13075 2593 13109 2627
rect 13144 2593 13178 2627
rect 13213 2593 13247 2627
rect 13282 2593 13316 2627
rect 13351 2593 13385 2627
rect 13420 2593 13454 2627
rect 13489 2593 13523 2627
rect 13558 2593 13592 2627
rect 13627 2593 13661 2627
rect 13696 2593 13730 2627
rect 13765 2593 13799 2627
rect 13834 2593 13868 2627
rect 13903 2593 13937 2627
rect 13972 2593 14006 2627
rect 14041 2593 14075 2627
rect 11476 2525 11510 2559
rect 11546 2525 11580 2559
rect 11616 2525 11650 2559
rect 11686 2525 11720 2559
rect 11756 2525 11790 2559
rect 11826 2525 11860 2559
rect 11896 2525 11930 2559
rect 11966 2525 12000 2559
rect 12036 2525 12070 2559
rect 12106 2525 12140 2559
rect 12176 2525 12210 2559
rect 12246 2525 12280 2559
rect 12316 2525 12350 2559
rect 12385 2525 12419 2559
rect 12454 2525 12488 2559
rect 12523 2525 12557 2559
rect 12592 2525 12626 2559
rect 12661 2525 12695 2559
rect 12730 2525 12764 2559
rect 12799 2525 12833 2559
rect 12868 2525 12902 2559
rect 12937 2525 12971 2559
rect 13006 2525 13040 2559
rect 13075 2525 13109 2559
rect 13144 2525 13178 2559
rect 13213 2525 13247 2559
rect 13282 2525 13316 2559
rect 13351 2525 13385 2559
rect 13420 2525 13454 2559
rect 13489 2525 13523 2559
rect 13558 2525 13592 2559
rect 13627 2525 13661 2559
rect 13696 2525 13730 2559
rect 13765 2525 13799 2559
rect 13834 2525 13868 2559
rect 13903 2525 13937 2559
rect 13972 2525 14006 2559
rect 14041 2525 14075 2559
rect 11476 2457 11510 2491
rect 11546 2457 11580 2491
rect 11616 2457 11650 2491
rect 11686 2457 11720 2491
rect 11756 2457 11790 2491
rect 11826 2457 11860 2491
rect 11896 2457 11930 2491
rect 11966 2457 12000 2491
rect 12036 2457 12070 2491
rect 12106 2457 12140 2491
rect 12176 2457 12210 2491
rect 12246 2457 12280 2491
rect 12316 2457 12350 2491
rect 12385 2457 12419 2491
rect 12454 2457 12488 2491
rect 12523 2457 12557 2491
rect 12592 2457 12626 2491
rect 12661 2457 12695 2491
rect 12730 2457 12764 2491
rect 12799 2457 12833 2491
rect 12868 2457 12902 2491
rect 12937 2457 12971 2491
rect 13006 2457 13040 2491
rect 13075 2457 13109 2491
rect 13144 2457 13178 2491
rect 13213 2457 13247 2491
rect 13282 2457 13316 2491
rect 13351 2457 13385 2491
rect 13420 2457 13454 2491
rect 13489 2457 13523 2491
rect 13558 2457 13592 2491
rect 13627 2457 13661 2491
rect 13696 2457 13730 2491
rect 13765 2457 13799 2491
rect 13834 2457 13868 2491
rect 13903 2457 13937 2491
rect 13972 2457 14006 2491
rect 14041 2457 14075 2491
rect 11476 2389 11510 2423
rect 11546 2389 11580 2423
rect 11616 2389 11650 2423
rect 11686 2389 11720 2423
rect 11756 2389 11790 2423
rect 11826 2389 11860 2423
rect 11896 2389 11930 2423
rect 11966 2389 12000 2423
rect 12036 2389 12070 2423
rect 12106 2389 12140 2423
rect 12176 2389 12210 2423
rect 12246 2389 12280 2423
rect 12316 2389 12350 2423
rect 12385 2389 12419 2423
rect 12454 2389 12488 2423
rect 12523 2389 12557 2423
rect 12592 2389 12626 2423
rect 12661 2389 12695 2423
rect 12730 2389 12764 2423
rect 12799 2389 12833 2423
rect 12868 2389 12902 2423
rect 12937 2389 12971 2423
rect 13006 2389 13040 2423
rect 13075 2389 13109 2423
rect 13144 2389 13178 2423
rect 13213 2389 13247 2423
rect 13282 2389 13316 2423
rect 13351 2389 13385 2423
rect 13420 2389 13454 2423
rect 13489 2389 13523 2423
rect 13558 2389 13592 2423
rect 13627 2389 13661 2423
rect 13696 2389 13730 2423
rect 13765 2389 13799 2423
rect 13834 2389 13868 2423
rect 13903 2389 13937 2423
rect 13972 2389 14006 2423
rect 14041 2389 14075 2423
rect 11476 2321 11510 2355
rect 11546 2321 11580 2355
rect 11616 2321 11650 2355
rect 11686 2321 11720 2355
rect 11756 2321 11790 2355
rect 11826 2321 11860 2355
rect 11896 2321 11930 2355
rect 11966 2321 12000 2355
rect 12036 2321 12070 2355
rect 12106 2321 12140 2355
rect 12176 2321 12210 2355
rect 12246 2321 12280 2355
rect 12316 2321 12350 2355
rect 12385 2321 12419 2355
rect 12454 2321 12488 2355
rect 12523 2321 12557 2355
rect 12592 2321 12626 2355
rect 12661 2321 12695 2355
rect 12730 2321 12764 2355
rect 12799 2321 12833 2355
rect 12868 2321 12902 2355
rect 12937 2321 12971 2355
rect 13006 2321 13040 2355
rect 13075 2321 13109 2355
rect 13144 2321 13178 2355
rect 13213 2321 13247 2355
rect 13282 2321 13316 2355
rect 13351 2321 13385 2355
rect 13420 2321 13454 2355
rect 13489 2321 13523 2355
rect 13558 2321 13592 2355
rect 13627 2321 13661 2355
rect 13696 2321 13730 2355
rect 13765 2321 13799 2355
rect 13834 2321 13868 2355
rect 13903 2321 13937 2355
rect 13972 2321 14006 2355
rect 14041 2321 14075 2355
rect 11476 2253 11510 2287
rect 11546 2253 11580 2287
rect 11616 2253 11650 2287
rect 11686 2253 11720 2287
rect 11756 2253 11790 2287
rect 11826 2253 11860 2287
rect 11896 2253 11930 2287
rect 11966 2253 12000 2287
rect 12036 2253 12070 2287
rect 12106 2253 12140 2287
rect 12176 2253 12210 2287
rect 12246 2253 12280 2287
rect 12316 2253 12350 2287
rect 12385 2253 12419 2287
rect 12454 2253 12488 2287
rect 12523 2253 12557 2287
rect 12592 2253 12626 2287
rect 12661 2253 12695 2287
rect 12730 2253 12764 2287
rect 12799 2253 12833 2287
rect 12868 2253 12902 2287
rect 12937 2253 12971 2287
rect 13006 2253 13040 2287
rect 13075 2253 13109 2287
rect 13144 2253 13178 2287
rect 13213 2253 13247 2287
rect 13282 2253 13316 2287
rect 13351 2253 13385 2287
rect 13420 2253 13454 2287
rect 13489 2253 13523 2287
rect 13558 2253 13592 2287
rect 13627 2253 13661 2287
rect 13696 2253 13730 2287
rect 13765 2253 13799 2287
rect 13834 2253 13868 2287
rect 13903 2253 13937 2287
rect 13972 2253 14006 2287
rect 14041 2253 14075 2287
rect 11476 2185 11510 2219
rect 11546 2185 11580 2219
rect 11616 2185 11650 2219
rect 11686 2185 11720 2219
rect 11756 2185 11790 2219
rect 11826 2185 11860 2219
rect 11896 2185 11930 2219
rect 11966 2185 12000 2219
rect 12036 2185 12070 2219
rect 12106 2185 12140 2219
rect 12176 2185 12210 2219
rect 12246 2185 12280 2219
rect 12316 2185 12350 2219
rect 12385 2185 12419 2219
rect 12454 2185 12488 2219
rect 12523 2185 12557 2219
rect 12592 2185 12626 2219
rect 12661 2185 12695 2219
rect 12730 2185 12764 2219
rect 12799 2185 12833 2219
rect 12868 2185 12902 2219
rect 12937 2185 12971 2219
rect 13006 2185 13040 2219
rect 13075 2185 13109 2219
rect 13144 2185 13178 2219
rect 13213 2185 13247 2219
rect 13282 2185 13316 2219
rect 13351 2185 13385 2219
rect 13420 2185 13454 2219
rect 13489 2185 13523 2219
rect 13558 2185 13592 2219
rect 13627 2185 13661 2219
rect 13696 2185 13730 2219
rect 13765 2185 13799 2219
rect 13834 2185 13868 2219
rect 13903 2185 13937 2219
rect 13972 2185 14006 2219
rect 14041 2185 14075 2219
rect 11476 2117 11510 2151
rect 11546 2117 11580 2151
rect 11616 2117 11650 2151
rect 11686 2117 11720 2151
rect 11756 2117 11790 2151
rect 11826 2117 11860 2151
rect 11896 2117 11930 2151
rect 11966 2117 12000 2151
rect 12036 2117 12070 2151
rect 12106 2117 12140 2151
rect 12176 2117 12210 2151
rect 12246 2117 12280 2151
rect 12316 2117 12350 2151
rect 12385 2117 12419 2151
rect 12454 2117 12488 2151
rect 12523 2117 12557 2151
rect 12592 2117 12626 2151
rect 12661 2117 12695 2151
rect 12730 2117 12764 2151
rect 12799 2117 12833 2151
rect 12868 2117 12902 2151
rect 12937 2117 12971 2151
rect 13006 2117 13040 2151
rect 13075 2117 13109 2151
rect 13144 2117 13178 2151
rect 13213 2117 13247 2151
rect 13282 2117 13316 2151
rect 13351 2117 13385 2151
rect 13420 2117 13454 2151
rect 13489 2117 13523 2151
rect 13558 2117 13592 2151
rect 13627 2117 13661 2151
rect 13696 2117 13730 2151
rect 13765 2117 13799 2151
rect 13834 2117 13868 2151
rect 13903 2117 13937 2151
rect 13972 2117 14006 2151
rect 14041 2117 14075 2151
rect 11476 2049 11510 2083
rect 11546 2049 11580 2083
rect 11616 2049 11650 2083
rect 11686 2049 11720 2083
rect 11756 2049 11790 2083
rect 11826 2049 11860 2083
rect 11896 2049 11930 2083
rect 11966 2049 12000 2083
rect 12036 2049 12070 2083
rect 12106 2049 12140 2083
rect 12176 2049 12210 2083
rect 12246 2049 12280 2083
rect 12316 2049 12350 2083
rect 12385 2049 12419 2083
rect 12454 2049 12488 2083
rect 12523 2049 12557 2083
rect 12592 2049 12626 2083
rect 12661 2049 12695 2083
rect 12730 2049 12764 2083
rect 12799 2049 12833 2083
rect 12868 2049 12902 2083
rect 12937 2049 12971 2083
rect 13006 2049 13040 2083
rect 13075 2049 13109 2083
rect 13144 2049 13178 2083
rect 13213 2049 13247 2083
rect 13282 2049 13316 2083
rect 13351 2049 13385 2083
rect 13420 2049 13454 2083
rect 13489 2049 13523 2083
rect 13558 2049 13592 2083
rect 13627 2049 13661 2083
rect 13696 2049 13730 2083
rect 13765 2049 13799 2083
rect 13834 2049 13868 2083
rect 13903 2049 13937 2083
rect 13972 2049 14006 2083
rect 14041 2049 14075 2083
rect 11476 1981 11510 2015
rect 11546 1981 11580 2015
rect 11616 1981 11650 2015
rect 11686 1981 11720 2015
rect 11756 1981 11790 2015
rect 11826 1981 11860 2015
rect 11896 1981 11930 2015
rect 11966 1981 12000 2015
rect 12036 1981 12070 2015
rect 12106 1981 12140 2015
rect 12176 1981 12210 2015
rect 12246 1981 12280 2015
rect 12316 1981 12350 2015
rect 12385 1981 12419 2015
rect 12454 1981 12488 2015
rect 12523 1981 12557 2015
rect 12592 1981 12626 2015
rect 12661 1981 12695 2015
rect 12730 1981 12764 2015
rect 12799 1981 12833 2015
rect 12868 1981 12902 2015
rect 12937 1981 12971 2015
rect 13006 1981 13040 2015
rect 13075 1981 13109 2015
rect 13144 1981 13178 2015
rect 13213 1981 13247 2015
rect 13282 1981 13316 2015
rect 13351 1981 13385 2015
rect 13420 1981 13454 2015
rect 13489 1981 13523 2015
rect 13558 1981 13592 2015
rect 13627 1981 13661 2015
rect 13696 1981 13730 2015
rect 13765 1981 13799 2015
rect 13834 1981 13868 2015
rect 13903 1981 13937 2015
rect 13972 1981 14006 2015
rect 14041 1981 14075 2015
rect 11476 1913 11510 1947
rect 11546 1913 11580 1947
rect 11616 1913 11650 1947
rect 11686 1913 11720 1947
rect 11756 1913 11790 1947
rect 11826 1913 11860 1947
rect 11896 1913 11930 1947
rect 11966 1913 12000 1947
rect 12036 1913 12070 1947
rect 12106 1913 12140 1947
rect 12176 1913 12210 1947
rect 12246 1913 12280 1947
rect 12316 1913 12350 1947
rect 12385 1913 12419 1947
rect 12454 1913 12488 1947
rect 12523 1913 12557 1947
rect 12592 1913 12626 1947
rect 12661 1913 12695 1947
rect 12730 1913 12764 1947
rect 12799 1913 12833 1947
rect 12868 1913 12902 1947
rect 12937 1913 12971 1947
rect 13006 1913 13040 1947
rect 13075 1913 13109 1947
rect 13144 1913 13178 1947
rect 13213 1913 13247 1947
rect 13282 1913 13316 1947
rect 13351 1913 13385 1947
rect 13420 1913 13454 1947
rect 13489 1913 13523 1947
rect 13558 1913 13592 1947
rect 13627 1913 13661 1947
rect 13696 1913 13730 1947
rect 13765 1913 13799 1947
rect 13834 1913 13868 1947
rect 13903 1913 13937 1947
rect 13972 1913 14006 1947
rect 14041 1913 14075 1947
rect 11476 1845 11510 1879
rect 11546 1845 11580 1879
rect 11616 1845 11650 1879
rect 11686 1845 11720 1879
rect 11756 1845 11790 1879
rect 11826 1845 11860 1879
rect 11896 1845 11930 1879
rect 11966 1845 12000 1879
rect 12036 1845 12070 1879
rect 12106 1845 12140 1879
rect 12176 1845 12210 1879
rect 12246 1845 12280 1879
rect 12316 1845 12350 1879
rect 12385 1845 12419 1879
rect 12454 1845 12488 1879
rect 12523 1845 12557 1879
rect 12592 1845 12626 1879
rect 12661 1845 12695 1879
rect 12730 1845 12764 1879
rect 12799 1845 12833 1879
rect 12868 1845 12902 1879
rect 12937 1845 12971 1879
rect 13006 1845 13040 1879
rect 13075 1845 13109 1879
rect 13144 1845 13178 1879
rect 13213 1845 13247 1879
rect 13282 1845 13316 1879
rect 13351 1845 13385 1879
rect 13420 1845 13454 1879
rect 13489 1845 13523 1879
rect 13558 1845 13592 1879
rect 13627 1845 13661 1879
rect 13696 1845 13730 1879
rect 13765 1845 13799 1879
rect 13834 1845 13868 1879
rect 13903 1845 13937 1879
rect 13972 1845 14006 1879
rect 14041 1845 14075 1879
rect 11476 1777 11510 1811
rect 11546 1777 11580 1811
rect 11616 1777 11650 1811
rect 11686 1777 11720 1811
rect 11756 1777 11790 1811
rect 11826 1777 11860 1811
rect 11896 1777 11930 1811
rect 11966 1777 12000 1811
rect 12036 1777 12070 1811
rect 12106 1777 12140 1811
rect 12176 1777 12210 1811
rect 12246 1777 12280 1811
rect 12316 1777 12350 1811
rect 12385 1777 12419 1811
rect 12454 1777 12488 1811
rect 12523 1777 12557 1811
rect 12592 1777 12626 1811
rect 12661 1777 12695 1811
rect 12730 1777 12764 1811
rect 12799 1777 12833 1811
rect 12868 1777 12902 1811
rect 12937 1777 12971 1811
rect 13006 1777 13040 1811
rect 13075 1777 13109 1811
rect 13144 1777 13178 1811
rect 13213 1777 13247 1811
rect 13282 1777 13316 1811
rect 13351 1777 13385 1811
rect 13420 1777 13454 1811
rect 13489 1777 13523 1811
rect 13558 1777 13592 1811
rect 13627 1777 13661 1811
rect 13696 1777 13730 1811
rect 13765 1777 13799 1811
rect 13834 1777 13868 1811
rect 13903 1777 13937 1811
rect 13972 1777 14006 1811
rect 14041 1777 14075 1811
rect 11476 1709 11510 1743
rect 11546 1709 11580 1743
rect 11616 1709 11650 1743
rect 11686 1709 11720 1743
rect 11756 1709 11790 1743
rect 11826 1709 11860 1743
rect 11896 1709 11930 1743
rect 11966 1709 12000 1743
rect 12036 1709 12070 1743
rect 12106 1709 12140 1743
rect 12176 1709 12210 1743
rect 12246 1709 12280 1743
rect 12316 1709 12350 1743
rect 12385 1709 12419 1743
rect 12454 1709 12488 1743
rect 12523 1709 12557 1743
rect 12592 1709 12626 1743
rect 12661 1709 12695 1743
rect 12730 1709 12764 1743
rect 12799 1709 12833 1743
rect 12868 1709 12902 1743
rect 12937 1709 12971 1743
rect 13006 1709 13040 1743
rect 13075 1709 13109 1743
rect 13144 1709 13178 1743
rect 13213 1709 13247 1743
rect 13282 1709 13316 1743
rect 13351 1709 13385 1743
rect 13420 1709 13454 1743
rect 13489 1709 13523 1743
rect 13558 1709 13592 1743
rect 13627 1709 13661 1743
rect 13696 1709 13730 1743
rect 13765 1709 13799 1743
rect 13834 1709 13868 1743
rect 13903 1709 13937 1743
rect 13972 1709 14006 1743
rect 14041 1709 14075 1743
rect 11476 1641 11510 1675
rect 11546 1641 11580 1675
rect 11616 1641 11650 1675
rect 11686 1641 11720 1675
rect 11756 1641 11790 1675
rect 11826 1641 11860 1675
rect 11896 1641 11930 1675
rect 11966 1641 12000 1675
rect 12036 1641 12070 1675
rect 12106 1641 12140 1675
rect 12176 1641 12210 1675
rect 12246 1641 12280 1675
rect 12316 1641 12350 1675
rect 12385 1641 12419 1675
rect 12454 1641 12488 1675
rect 12523 1641 12557 1675
rect 12592 1641 12626 1675
rect 12661 1641 12695 1675
rect 12730 1641 12764 1675
rect 12799 1641 12833 1675
rect 12868 1641 12902 1675
rect 12937 1641 12971 1675
rect 13006 1641 13040 1675
rect 13075 1641 13109 1675
rect 13144 1641 13178 1675
rect 13213 1641 13247 1675
rect 13282 1641 13316 1675
rect 13351 1641 13385 1675
rect 13420 1641 13454 1675
rect 13489 1641 13523 1675
rect 13558 1641 13592 1675
rect 13627 1641 13661 1675
rect 13696 1641 13730 1675
rect 13765 1641 13799 1675
rect 13834 1641 13868 1675
rect 13903 1641 13937 1675
rect 13972 1641 14006 1675
rect 14041 1641 14075 1675
rect 12957 1532 12991 1566
rect 13030 1532 13064 1566
rect 13103 1532 13137 1566
rect 13176 1532 13210 1566
rect 13249 1532 13283 1566
rect 13321 1532 13355 1566
rect 13393 1532 13427 1566
rect 13465 1532 13499 1566
rect 13537 1532 13571 1566
rect 13609 1532 13643 1566
rect 13681 1532 13715 1566
rect 13753 1532 13787 1566
rect 13825 1532 13859 1566
rect 13897 1532 13931 1566
rect 13969 1532 14003 1566
rect 14041 1532 14075 1566
rect 12957 1464 12991 1498
rect 13030 1464 13064 1498
rect 13103 1464 13137 1498
rect 13176 1464 13210 1498
rect 13249 1464 13283 1498
rect 13321 1464 13355 1498
rect 13393 1464 13427 1498
rect 13465 1464 13499 1498
rect 13537 1464 13571 1498
rect 13609 1464 13643 1498
rect 13681 1464 13715 1498
rect 13753 1464 13787 1498
rect 13825 1464 13859 1498
rect 13897 1464 13931 1498
rect 13969 1464 14003 1498
rect 14041 1464 14075 1498
rect 12957 1396 12991 1430
rect 13030 1396 13064 1430
rect 13103 1396 13137 1430
rect 13176 1396 13210 1430
rect 13249 1396 13283 1430
rect 13321 1396 13355 1430
rect 13393 1396 13427 1430
rect 13465 1396 13499 1430
rect 13537 1396 13571 1430
rect 13609 1396 13643 1430
rect 13681 1396 13715 1430
rect 13753 1396 13787 1430
rect 13825 1396 13859 1430
rect 13897 1396 13931 1430
rect 13969 1396 14003 1430
rect 14041 1396 14075 1430
<< mvnsubdiffcont >>
rect 123 6389 157 6423
rect 0 6355 34 6389
rect 0 6287 102 6355
rect 191 6321 2061 6423
rect 2129 6389 2163 6423
rect 2198 6389 2232 6423
rect 2267 6389 2301 6423
rect 2336 6389 2370 6423
rect 2405 6389 2439 6423
rect 2474 6389 2508 6423
rect 2543 6389 2577 6423
rect 2612 6389 2646 6423
rect 2681 6389 2715 6423
rect 2750 6389 2784 6423
rect 2819 6389 2853 6423
rect 2888 6389 2922 6423
rect 2957 6389 2991 6423
rect 3026 6389 3060 6423
rect 3095 6389 3129 6423
rect 3164 6389 3198 6423
rect 3233 6389 3267 6423
rect 3302 6389 3336 6423
rect 3371 6389 3405 6423
rect 3440 6389 3474 6423
rect 3509 6389 3543 6423
rect 3578 6389 3612 6423
rect 3647 6389 3681 6423
rect 3716 6389 3750 6423
rect 3785 6389 3819 6423
rect 3854 6389 3888 6423
rect 3923 6389 3957 6423
rect 3992 6389 4026 6423
rect 4061 6389 4095 6423
rect 4130 6389 4164 6423
rect 4199 6389 4233 6423
rect 4268 6389 4302 6423
rect 4337 6389 4371 6423
rect 4406 6389 4440 6423
rect 4475 6389 4509 6423
rect 4544 6389 4578 6423
rect 4613 6389 4647 6423
rect 4682 6389 4716 6423
rect 4751 6389 4785 6423
rect 4820 6389 4854 6423
rect 4889 6389 4923 6423
rect 4958 6389 4992 6423
rect 5027 6389 5061 6423
rect 5096 6389 5130 6423
rect 5165 6389 5199 6423
rect 5234 6389 5268 6423
rect 5303 6389 5337 6423
rect 5372 6389 5406 6423
rect 5441 6389 5475 6423
rect 5510 6389 5544 6423
rect 5579 6389 5613 6423
rect 5648 6389 5682 6423
rect 5717 6389 5751 6423
rect 5786 6389 5820 6423
rect 5855 6389 5889 6423
rect 5924 6355 7658 6423
rect 7726 6355 7760 6389
rect 2129 6321 2163 6355
rect 2198 6321 2232 6355
rect 2267 6321 2301 6355
rect 2336 6321 2370 6355
rect 2405 6321 2439 6355
rect 2474 6321 2508 6355
rect 2543 6321 2577 6355
rect 2612 6321 2646 6355
rect 2681 6321 2715 6355
rect 2750 6321 2784 6355
rect 2819 6321 2853 6355
rect 2888 6321 2922 6355
rect 2957 6321 2991 6355
rect 3026 6321 3060 6355
rect 3095 6321 3129 6355
rect 3164 6321 3198 6355
rect 3233 6321 3267 6355
rect 3302 6321 3336 6355
rect 3371 6321 3405 6355
rect 3440 6321 3474 6355
rect 3509 6321 3543 6355
rect 3578 6321 7692 6355
rect 7794 6321 9732 6423
rect 9766 6389 9800 6423
rect 9874 6355 9908 6389
rect 0 3295 170 6287
rect 259 6253 2061 6321
rect 2129 6253 2163 6287
rect 2198 6253 2232 6287
rect 2267 6253 2301 6287
rect 2336 6253 2370 6287
rect 2405 6253 2439 6287
rect 2474 6253 2508 6287
rect 2543 6253 2577 6287
rect 2612 6253 2646 6287
rect 2681 6253 2715 6287
rect 2750 6253 2784 6287
rect 2819 6253 2853 6287
rect 2888 6253 2922 6287
rect 2957 6253 2991 6287
rect 3026 6253 3060 6287
rect 3095 6253 3129 6287
rect 3164 6253 3198 6287
rect 3233 6253 3267 6287
rect 3302 6253 3336 6287
rect 3371 6253 3405 6287
rect 3440 6253 3474 6287
rect 3509 6253 3543 6287
rect 3578 6253 7624 6321
rect 7794 6320 9664 6321
rect 7658 6252 7692 6286
rect 7726 6253 9664 6320
rect 9806 6287 9908 6355
rect 7726 6218 7760 6252
rect 7590 6184 7624 6218
rect 7658 6183 7692 6217
rect 7726 6150 7760 6184
rect 7590 6115 7624 6149
rect 7658 6114 7692 6148
rect 7726 6082 7760 6116
rect 7590 6046 7624 6080
rect 7658 6045 7692 6079
rect 7726 6014 7760 6048
rect 7590 5977 7624 6011
rect 7658 5976 7692 6010
rect 7726 5946 7760 5980
rect 7590 5908 7624 5942
rect 7658 5907 7692 5941
rect 7726 5878 7760 5912
rect 7590 5839 7624 5873
rect 7658 5838 7692 5872
rect 7726 5810 7760 5844
rect 7590 5770 7624 5804
rect 7658 5769 7692 5803
rect 7726 5742 7760 5776
rect 7590 5701 7624 5735
rect 7658 5700 7692 5734
rect 7726 5674 7760 5708
rect 7590 5632 7624 5666
rect 7658 5631 7692 5665
rect 7726 5606 7760 5640
rect 7590 5563 7624 5597
rect 7658 5562 7692 5596
rect 7726 5538 7760 5572
rect 7590 5494 7624 5528
rect 7658 5493 7692 5527
rect 7726 5470 7760 5504
rect 7590 5425 7624 5459
rect 7658 5424 7692 5458
rect 7726 5402 7760 5436
rect 7590 5356 7624 5390
rect 7658 5355 7692 5389
rect 7726 5334 7760 5368
rect 7590 5287 7624 5321
rect 7658 5286 7692 5320
rect 7726 5266 7760 5300
rect 7590 5218 7624 5252
rect 7658 5217 7692 5251
rect 7726 5198 7760 5232
rect 7590 5149 7624 5183
rect 7658 5148 7692 5182
rect 7726 5130 7760 5164
rect 7590 5080 7624 5114
rect 7658 5079 7692 5113
rect 7726 5062 7760 5096
rect 7590 5011 7624 5045
rect 7658 5010 7692 5044
rect 7726 4994 7760 5028
rect 7590 4942 7624 4976
rect 7658 4941 7692 4975
rect 7726 4926 7760 4960
rect 7590 4873 7624 4907
rect 7658 4872 7692 4906
rect 7726 4858 7760 4892
rect 7590 4804 7624 4838
rect 7658 4803 7692 4837
rect 7726 4790 7760 4824
rect 7590 4735 7624 4769
rect 7658 4734 7692 4768
rect 7726 4722 7760 4756
rect 7590 4666 7624 4700
rect 7658 4665 7692 4699
rect 7726 4654 7760 4688
rect 7590 4597 7624 4631
rect 7658 4596 7692 4630
rect 7726 4586 7760 4620
rect 7590 4528 7624 4562
rect 7658 4527 7692 4561
rect 7726 4518 7760 4552
rect 7590 4459 7624 4493
rect 7658 4458 7692 4492
rect 7726 4450 7760 4484
rect 7590 4390 7624 4424
rect 7658 4389 7692 4423
rect 7726 4382 7760 4416
rect 7590 4321 7624 4355
rect 7658 4320 7692 4354
rect 7726 4314 7760 4348
rect 7590 4252 7624 4286
rect 7658 4251 7692 4285
rect 7726 4246 7760 4280
rect 7590 4183 7624 4217
rect 7658 4182 7692 4216
rect 7726 4178 7760 4212
rect 7590 4114 7624 4148
rect 7658 4113 7692 4147
rect 7726 4110 7760 4144
rect 7590 4045 7624 4079
rect 7658 4044 7692 4078
rect 7726 4042 7760 4076
rect 7590 3976 7624 4010
rect 7658 3975 7692 4009
rect 7726 3974 7760 4008
rect 7590 3907 7624 3941
rect 7658 3872 7760 3940
rect 7590 3498 7760 3872
rect 68 3261 170 3295
rect 9738 3370 9908 6287
rect 10617 6378 10651 6412
rect 10685 6378 10719 6412
rect 10753 6378 10787 6412
rect 10821 6378 10855 6412
rect 10889 6378 10923 6412
rect 10957 6378 10991 6412
rect 11025 6378 11059 6412
rect 11093 6378 11127 6412
rect 11161 6378 11195 6412
rect 11229 6378 11263 6412
rect 11297 6378 11331 6412
rect 11365 6378 11399 6412
rect 11480 6378 11514 6412
rect 11548 6378 11582 6412
rect 11616 6378 11650 6412
rect 11684 6378 11718 6412
rect 11752 6378 11786 6412
rect 11820 6378 11854 6412
rect 11888 6378 11922 6412
rect 11956 6378 11990 6412
rect 12024 6378 12058 6412
rect 12092 6378 12126 6412
rect 12160 6378 12194 6412
rect 12228 6378 12262 6412
rect 12296 6378 12330 6412
rect 12364 6378 12398 6412
rect 12432 6378 12466 6412
rect 12500 6378 12534 6412
rect 12568 6378 12602 6412
rect 12636 6378 12670 6412
rect 12704 6378 12738 6412
rect 12772 6378 12806 6412
rect 12840 6378 12874 6412
rect 12908 6378 12942 6412
rect 12976 6378 13010 6412
rect 13044 6378 13078 6412
rect 13112 6378 13146 6412
rect 13258 6378 13292 6412
rect 13326 6378 13360 6412
rect 13394 6378 13428 6412
rect 13462 6378 13496 6412
rect 10498 6344 10532 6378
rect 10498 6276 10532 6310
rect 13496 6294 13530 6328
rect 10498 6208 10532 6242
rect 13496 6226 13530 6260
rect 10498 6140 10532 6174
rect 10498 6072 10532 6106
rect 10498 6004 10532 6038
rect 10498 5936 10532 5970
rect 10498 5868 10532 5902
rect 10498 5800 10532 5834
rect 10498 5732 10532 5766
rect 10498 5664 10532 5698
rect 10498 5596 10532 5630
rect 10498 5528 10532 5562
rect 13496 6158 13530 6192
rect 13496 6090 13530 6124
rect 13496 6022 13530 6056
rect 13496 5954 13530 5988
rect 13496 5886 13530 5920
rect 13496 5818 13530 5852
rect 13496 5750 13530 5784
rect 13496 5682 13530 5716
rect 13496 5563 13530 5597
rect 10498 5460 10532 5494
rect 13496 5495 13530 5529
rect 10498 5392 10532 5426
rect 10498 5324 10532 5358
rect 10498 5256 10532 5290
rect 10498 5188 10532 5222
rect 10498 5120 10532 5154
rect 10498 5052 10532 5086
rect 10498 4984 10532 5018
rect 10498 4916 10532 4950
rect 10498 4848 10532 4882
rect 10498 4780 10532 4814
rect 13496 5427 13530 5461
rect 13496 5359 13530 5393
rect 13496 5291 13530 5325
rect 13496 5223 13530 5257
rect 13496 5155 13530 5189
rect 13496 5087 13530 5121
rect 13496 5019 13530 5053
rect 13496 4951 13530 4985
rect 13496 4883 13530 4917
rect 13496 4815 13530 4849
rect 10498 4712 10532 4746
rect 13496 4747 13530 4781
rect 10498 4644 10532 4678
rect 10498 4576 10532 4610
rect 10498 4508 10532 4542
rect 10498 4440 10532 4474
rect 10498 4372 10532 4406
rect 10498 4304 10532 4338
rect 10498 4236 10532 4270
rect 10498 4168 10532 4202
rect 10498 4100 10532 4134
rect 13496 4679 13530 4713
rect 13496 4611 13530 4645
rect 13496 4543 13530 4577
rect 13496 4475 13530 4509
rect 13496 4407 13530 4441
rect 13496 4339 13530 4373
rect 13496 4271 13530 4305
rect 13496 4203 13530 4237
rect 13496 4135 13530 4169
rect 13496 4067 13530 4101
rect 13496 3999 13530 4033
rect 10532 3965 10566 3999
rect 10600 3965 10634 3999
rect 10668 3965 10702 3999
rect 10736 3965 10770 3999
rect 10804 3965 10838 3999
rect 10872 3965 10906 3999
rect 10940 3965 10974 3999
rect 11008 3965 11042 3999
rect 11076 3965 11110 3999
rect 11144 3965 11178 3999
rect 11212 3965 11246 3999
rect 11280 3965 11314 3999
rect 11348 3965 11382 3999
rect 11416 3965 11450 3999
rect 11484 3965 11518 3999
rect 11552 3965 11586 3999
rect 11620 3965 11654 3999
rect 11688 3965 11722 3999
rect 11756 3965 11790 3999
rect 11824 3965 11858 3999
rect 11892 3965 11926 3999
rect 11960 3965 11994 3999
rect 12028 3965 12062 3999
rect 12096 3965 12130 3999
rect 12164 3965 12198 3999
rect 12232 3965 12266 3999
rect 12300 3965 12334 3999
rect 12368 3965 12402 3999
rect 12436 3965 12470 3999
rect 12504 3965 12538 3999
rect 12572 3965 12606 3999
rect 12640 3965 12674 3999
rect 12708 3965 12742 3999
rect 12776 3965 12810 3999
rect 12844 3965 12878 3999
rect 12912 3965 12946 3999
rect 12980 3965 13014 3999
rect 13048 3965 13082 3999
rect 13116 3965 13150 3999
rect 13184 3965 13218 3999
rect 13252 3965 13286 3999
rect 13320 3965 13354 3999
rect 13388 3965 13422 3999
rect 9738 3295 11132 3370
rect 11166 3336 11200 3370
rect 11252 3302 11286 3336
rect 9738 3261 9840 3295
rect 9942 3268 11132 3295
rect 9942 3200 11064 3268
rect 11184 3234 11286 3302
rect 11116 140 11286 3234
rect 11252 106 11286 140
<< poly >>
rect 2196 5859 2996 5875
rect 2196 5825 2212 5859
rect 2246 5825 2286 5859
rect 2320 5825 2360 5859
rect 2394 5825 2434 5859
rect 2468 5825 2508 5859
rect 2542 5825 2581 5859
rect 2615 5825 2654 5859
rect 2688 5825 2727 5859
rect 2761 5825 2800 5859
rect 2834 5825 2873 5859
rect 2907 5825 2946 5859
rect 2980 5825 2996 5859
rect 484 5803 2114 5809
rect 2196 5803 2996 5825
rect 3052 5859 4708 5875
rect 3052 5825 3068 5859
rect 3102 5825 3138 5859
rect 3172 5825 3208 5859
rect 3242 5825 3278 5859
rect 3312 5825 3347 5859
rect 3381 5825 3416 5859
rect 3450 5825 3485 5859
rect 3519 5825 3554 5859
rect 3588 5825 3623 5859
rect 3657 5825 3692 5859
rect 3726 5825 3761 5859
rect 3795 5825 3830 5859
rect 3864 5825 3899 5859
rect 3933 5825 3968 5859
rect 4002 5825 4037 5859
rect 4071 5825 4106 5859
rect 4140 5825 4175 5859
rect 4209 5825 4244 5859
rect 4278 5825 4313 5859
rect 4347 5825 4382 5859
rect 4416 5825 4451 5859
rect 4485 5825 4520 5859
rect 4554 5825 4589 5859
rect 4623 5825 4658 5859
rect 4692 5825 4708 5859
rect 3052 5803 4708 5825
rect 484 3729 2140 3751
rect 484 3695 523 3729
rect 557 3695 592 3729
rect 626 3695 661 3729
rect 695 3695 730 3729
rect 764 3695 799 3729
rect 833 3695 868 3729
rect 902 3695 937 3729
rect 971 3695 1006 3729
rect 1040 3695 1075 3729
rect 1109 3695 1143 3729
rect 1177 3695 1211 3729
rect 1245 3695 1380 3729
rect 1414 3695 1449 3729
rect 1483 3695 1518 3729
rect 1552 3695 1587 3729
rect 1621 3695 1656 3729
rect 1690 3695 1725 3729
rect 1759 3695 1794 3729
rect 1828 3695 1863 3729
rect 1897 3695 1931 3729
rect 1965 3695 1999 3729
rect 2033 3695 2067 3729
rect 2101 3695 2140 3729
rect 484 3679 2140 3695
rect 2196 3679 2996 3751
rect 3052 3729 4708 3751
rect 3052 3695 3091 3729
rect 3125 3695 3160 3729
rect 3194 3695 3229 3729
rect 3263 3695 3298 3729
rect 3332 3695 3367 3729
rect 3401 3695 3436 3729
rect 3470 3695 3505 3729
rect 3539 3695 3574 3729
rect 3608 3695 3643 3729
rect 3677 3695 3711 3729
rect 3745 3695 3779 3729
rect 3813 3695 3947 3729
rect 3981 3695 4016 3729
rect 4050 3695 4085 3729
rect 4119 3695 4154 3729
rect 4188 3695 4223 3729
rect 4257 3695 4292 3729
rect 4326 3695 4361 3729
rect 4395 3695 4430 3729
rect 4464 3695 4499 3729
rect 4533 3695 4567 3729
rect 4601 3695 4635 3729
rect 4669 3695 4708 3729
rect 3052 3679 4708 3695
rect 6750 3770 7276 3864
rect 8647 5397 8653 5939
rect 8761 5937 8833 5953
rect 8761 5903 8777 5937
rect 8811 5903 8833 5937
rect 8761 5869 8833 5903
rect 8761 5835 8777 5869
rect 8811 5835 8833 5869
rect 8761 5801 8833 5835
rect 8761 5767 8777 5801
rect 8811 5767 8833 5801
rect 8761 5733 8833 5767
rect 8761 5699 8777 5733
rect 8811 5699 8833 5733
rect 8761 5683 8833 5699
rect 8719 5515 8833 5531
rect 8719 5481 8777 5515
rect 8811 5481 8833 5515
rect 8719 5447 8833 5481
rect 8719 5413 8777 5447
rect 8811 5413 8833 5447
rect 8719 5397 8833 5413
rect 8647 5189 8719 5205
rect 8647 5155 8669 5189
rect 8703 5155 8719 5189
rect 8647 5121 8719 5155
rect 8647 5087 8669 5121
rect 8703 5087 8719 5121
rect 8647 5005 8719 5087
rect 8647 4933 8719 4949
rect 8647 4899 8669 4933
rect 8703 4899 8719 4933
rect 8647 4865 8719 4899
rect 8647 4831 8669 4865
rect 8703 4831 8719 4865
rect 8647 4653 8719 4831
rect 8827 4663 8833 5341
rect 8647 4581 8719 4597
rect 8761 4583 8833 4663
rect 8647 4547 8669 4581
rect 8703 4547 8719 4581
rect 8647 4513 8719 4547
rect 8647 4479 8669 4513
rect 8703 4479 8719 4513
rect 8647 4445 8719 4479
rect 8647 4411 8669 4445
rect 8703 4411 8719 4445
rect 8647 4397 8719 4411
rect 8653 4395 8719 4397
rect 8761 4511 8833 4527
rect 8761 4477 8777 4511
rect 8811 4477 8833 4511
rect 8761 4443 8833 4477
rect 8761 4409 8777 4443
rect 8811 4409 8833 4443
rect 8761 4393 8833 4409
rect 8761 4245 8833 4261
rect 8647 4212 8719 4231
rect 8647 4178 8669 4212
rect 8703 4178 8719 4212
rect 8647 4144 8719 4178
rect 8647 4110 8669 4144
rect 8703 4110 8719 4144
rect 8647 4076 8719 4110
rect 8647 4042 8669 4076
rect 8703 4042 8719 4076
rect 8647 4008 8719 4042
rect 8647 3974 8669 4008
rect 8703 3974 8719 4008
rect 8647 3935 8719 3974
rect 8761 4211 8777 4245
rect 8811 4211 8833 4245
rect 8761 4177 8833 4211
rect 8761 4143 8777 4177
rect 8811 4143 8833 4177
rect 8761 4109 8833 4143
rect 8761 4075 8777 4109
rect 8811 4075 8833 4109
rect 8761 4041 8833 4075
rect 8761 4007 8777 4041
rect 8811 4007 8833 4041
rect 8761 3965 8833 4007
rect 8647 3863 8719 3879
rect 8647 3829 8669 3863
rect 8703 3829 8719 3863
rect 8647 3795 8719 3829
rect 8647 3761 8669 3795
rect 8703 3761 8719 3795
rect 8647 3745 8719 3761
rect 8761 3799 8833 3909
rect 8761 3765 8777 3799
rect 8811 3765 8833 3799
rect 8761 3731 8833 3765
rect 8761 3697 8777 3731
rect 8811 3697 8833 3731
rect 8761 3663 8833 3697
rect 8761 3629 8777 3663
rect 8811 3629 8833 3663
rect 8761 3613 8833 3629
rect 8247 3577 8319 3593
rect 8247 3543 8269 3577
rect 8303 3543 8319 3577
rect 8247 3509 8319 3543
rect 8247 3475 8269 3509
rect 8303 3475 8319 3509
rect 8247 3459 8319 3475
rect 8361 3343 8427 3359
rect 8361 3309 8377 3343
rect 8411 3309 8427 3343
rect 8361 3293 8427 3309
rect 8361 3275 8433 3293
rect 8361 3241 8377 3275
rect 8411 3241 8433 3275
rect 8361 3193 8433 3241
rect 10659 6277 11211 6293
rect 10659 6243 10675 6277
rect 10709 6243 10743 6277
rect 10777 6243 10811 6277
rect 10845 6243 10879 6277
rect 10913 6243 10947 6277
rect 10981 6243 11211 6277
rect 10659 6221 11211 6243
rect 11945 6227 12281 6293
rect 11267 6221 12281 6227
rect 12568 6277 12702 6293
rect 12568 6243 12584 6277
rect 12618 6243 12652 6277
rect 12686 6243 12702 6277
rect 12568 6221 12702 6243
rect 12758 6277 13214 6293
rect 12758 6243 13096 6277
rect 13130 6243 13164 6277
rect 13198 6243 13214 6277
rect 12758 6221 13214 6243
rect 12003 5511 12137 5527
rect 12003 5477 12019 5511
rect 12053 5477 12087 5511
rect 12121 5477 12137 5511
rect 10629 5455 11851 5461
rect 12003 5455 12137 5477
rect 12186 5511 12320 5527
rect 12186 5477 12202 5511
rect 12236 5477 12270 5511
rect 12304 5477 12320 5511
rect 12186 5455 12320 5477
rect 12369 5511 12665 5527
rect 12369 5477 12385 5511
rect 12419 5477 12453 5511
rect 12487 5477 12521 5511
rect 12555 5477 12665 5511
rect 12369 5455 12665 5477
rect 12721 5455 13399 5461
rect 10659 4745 11851 4803
rect 10658 4087 13104 4093
rect 8060 2855 10778 2861
rect 12608 3234 12674 3250
rect 12608 3200 12624 3234
rect 12658 3232 12674 3234
rect 12658 3200 12680 3232
rect 12608 3166 12680 3200
rect 12608 3132 12624 3166
rect 12658 3132 12680 3166
rect 12608 3116 12680 3132
<< polycont >>
rect 2212 5825 2246 5859
rect 2286 5825 2320 5859
rect 2360 5825 2394 5859
rect 2434 5825 2468 5859
rect 2508 5825 2542 5859
rect 2581 5825 2615 5859
rect 2654 5825 2688 5859
rect 2727 5825 2761 5859
rect 2800 5825 2834 5859
rect 2873 5825 2907 5859
rect 2946 5825 2980 5859
rect 3068 5825 3102 5859
rect 3138 5825 3172 5859
rect 3208 5825 3242 5859
rect 3278 5825 3312 5859
rect 3347 5825 3381 5859
rect 3416 5825 3450 5859
rect 3485 5825 3519 5859
rect 3554 5825 3588 5859
rect 3623 5825 3657 5859
rect 3692 5825 3726 5859
rect 3761 5825 3795 5859
rect 3830 5825 3864 5859
rect 3899 5825 3933 5859
rect 3968 5825 4002 5859
rect 4037 5825 4071 5859
rect 4106 5825 4140 5859
rect 4175 5825 4209 5859
rect 4244 5825 4278 5859
rect 4313 5825 4347 5859
rect 4382 5825 4416 5859
rect 4451 5825 4485 5859
rect 4520 5825 4554 5859
rect 4589 5825 4623 5859
rect 4658 5825 4692 5859
rect 523 3695 557 3729
rect 592 3695 626 3729
rect 661 3695 695 3729
rect 730 3695 764 3729
rect 799 3695 833 3729
rect 868 3695 902 3729
rect 937 3695 971 3729
rect 1006 3695 1040 3729
rect 1075 3695 1109 3729
rect 1143 3695 1177 3729
rect 1211 3695 1245 3729
rect 1380 3695 1414 3729
rect 1449 3695 1483 3729
rect 1518 3695 1552 3729
rect 1587 3695 1621 3729
rect 1656 3695 1690 3729
rect 1725 3695 1759 3729
rect 1794 3695 1828 3729
rect 1863 3695 1897 3729
rect 1931 3695 1965 3729
rect 1999 3695 2033 3729
rect 2067 3695 2101 3729
rect 3091 3695 3125 3729
rect 3160 3695 3194 3729
rect 3229 3695 3263 3729
rect 3298 3695 3332 3729
rect 3367 3695 3401 3729
rect 3436 3695 3470 3729
rect 3505 3695 3539 3729
rect 3574 3695 3608 3729
rect 3643 3695 3677 3729
rect 3711 3695 3745 3729
rect 3779 3695 3813 3729
rect 3947 3695 3981 3729
rect 4016 3695 4050 3729
rect 4085 3695 4119 3729
rect 4154 3695 4188 3729
rect 4223 3695 4257 3729
rect 4292 3695 4326 3729
rect 4361 3695 4395 3729
rect 4430 3695 4464 3729
rect 4499 3695 4533 3729
rect 4567 3695 4601 3729
rect 4635 3695 4669 3729
rect 8777 5903 8811 5937
rect 8777 5835 8811 5869
rect 8777 5767 8811 5801
rect 8777 5699 8811 5733
rect 8777 5481 8811 5515
rect 8777 5413 8811 5447
rect 8669 5155 8703 5189
rect 8669 5087 8703 5121
rect 8669 4899 8703 4933
rect 8669 4831 8703 4865
rect 8669 4547 8703 4581
rect 8669 4479 8703 4513
rect 8669 4411 8703 4445
rect 8777 4477 8811 4511
rect 8777 4409 8811 4443
rect 8669 4178 8703 4212
rect 8669 4110 8703 4144
rect 8669 4042 8703 4076
rect 8669 3974 8703 4008
rect 8777 4211 8811 4245
rect 8777 4143 8811 4177
rect 8777 4075 8811 4109
rect 8777 4007 8811 4041
rect 8669 3829 8703 3863
rect 8669 3761 8703 3795
rect 8777 3765 8811 3799
rect 8777 3697 8811 3731
rect 8777 3629 8811 3663
rect 8269 3543 8303 3577
rect 8269 3475 8303 3509
rect 8377 3309 8411 3343
rect 8377 3241 8411 3275
rect 10675 6243 10709 6277
rect 10743 6243 10777 6277
rect 10811 6243 10845 6277
rect 10879 6243 10913 6277
rect 10947 6243 10981 6277
rect 12584 6243 12618 6277
rect 12652 6243 12686 6277
rect 13096 6243 13130 6277
rect 13164 6243 13198 6277
rect 12019 5477 12053 5511
rect 12087 5477 12121 5511
rect 12202 5477 12236 5511
rect 12270 5477 12304 5511
rect 12385 5477 12419 5511
rect 12453 5477 12487 5511
rect 12521 5477 12555 5511
rect 12624 3200 12658 3234
rect 12624 3132 12658 3166
<< locali >>
rect 13975 6636 14099 7336
rect 13693 6602 14099 6636
rect 0 6433 74 6467
rect 108 6433 146 6467
rect 180 6433 218 6467
rect 252 6433 290 6467
rect 324 6433 362 6467
rect 396 6433 434 6467
rect 468 6433 506 6467
rect 540 6433 578 6467
rect 612 6433 650 6467
rect 684 6433 722 6467
rect 756 6433 794 6467
rect 828 6433 866 6467
rect 900 6433 938 6467
rect 972 6433 1010 6467
rect 1044 6433 1082 6467
rect 1116 6433 1154 6467
rect 1188 6433 1226 6467
rect 1260 6433 1298 6467
rect 1332 6433 1370 6467
rect 1404 6433 1442 6467
rect 1476 6433 1514 6467
rect 1548 6433 1586 6467
rect 1620 6433 1658 6467
rect 1692 6433 1730 6467
rect 1764 6433 1802 6467
rect 1836 6433 1874 6467
rect 1908 6433 1946 6467
rect 1980 6433 2018 6467
rect 2052 6433 2090 6467
rect 2124 6433 2162 6467
rect 2196 6433 2234 6467
rect 2268 6433 2306 6467
rect 2340 6433 2378 6467
rect 2412 6433 2450 6467
rect 2484 6433 2522 6467
rect 2556 6433 2594 6467
rect 2628 6433 2666 6467
rect 2700 6433 2738 6467
rect 2772 6433 2810 6467
rect 2844 6433 2882 6467
rect 2916 6433 2954 6467
rect 2988 6433 3026 6467
rect 3060 6433 3098 6467
rect 3132 6433 3170 6467
rect 3204 6433 3242 6467
rect 3276 6433 3314 6467
rect 3348 6433 3386 6467
rect 3420 6433 3458 6467
rect 3492 6433 3530 6467
rect 3564 6433 3602 6467
rect 3636 6433 3674 6467
rect 3708 6433 3746 6467
rect 3780 6433 3818 6467
rect 3852 6433 3890 6467
rect 3924 6433 3962 6467
rect 3996 6433 4034 6467
rect 4068 6433 4106 6467
rect 4140 6433 4178 6467
rect 4212 6433 4250 6467
rect 4284 6433 4322 6467
rect 4356 6433 4394 6467
rect 4428 6433 4466 6467
rect 4500 6433 4538 6467
rect 4572 6433 4610 6467
rect 4644 6433 4682 6467
rect 4716 6433 4754 6467
rect 4788 6433 4826 6467
rect 4860 6433 4898 6467
rect 4932 6433 4971 6467
rect 5005 6433 5044 6467
rect 5078 6433 5117 6467
rect 5151 6433 5190 6467
rect 5224 6433 5263 6467
rect 5297 6433 5336 6467
rect 5370 6433 5409 6467
rect 5443 6433 5482 6467
rect 5516 6433 5555 6467
rect 5589 6433 5628 6467
rect 5662 6433 5701 6467
rect 5735 6433 5774 6467
rect 5808 6433 5847 6467
rect 5881 6433 5920 6467
rect 5954 6433 5993 6467
rect 6027 6433 6066 6467
rect 6100 6433 6139 6467
rect 6173 6433 6212 6467
rect 6246 6433 6285 6467
rect 6319 6433 6358 6467
rect 6392 6433 6431 6467
rect 6465 6433 6504 6467
rect 6538 6433 6577 6467
rect 6611 6433 6650 6467
rect 6684 6433 6723 6467
rect 6757 6433 6796 6467
rect 6830 6433 6869 6467
rect 6903 6433 6942 6467
rect 6976 6433 7015 6467
rect 7049 6433 7088 6467
rect 7122 6433 7161 6467
rect 7195 6433 7234 6467
rect 7268 6433 7307 6467
rect 7341 6433 7380 6467
rect 7414 6433 7453 6467
rect 7487 6433 7526 6467
rect 7560 6433 7599 6467
rect 7633 6433 7672 6467
rect 7706 6433 7745 6467
rect 7779 6433 7818 6467
rect 7852 6433 7891 6467
rect 7925 6433 7964 6467
rect 7998 6433 8037 6467
rect 8071 6433 8110 6467
rect 8144 6433 8183 6467
rect 8217 6433 8256 6467
rect 8290 6433 8329 6467
rect 8363 6433 8402 6467
rect 8436 6433 8475 6467
rect 8509 6433 8548 6467
rect 8582 6433 8621 6467
rect 8655 6433 8694 6467
rect 8728 6433 8767 6467
rect 8801 6433 8840 6467
rect 8874 6433 8913 6467
rect 8947 6433 8986 6467
rect 9020 6433 9059 6467
rect 9093 6433 9132 6467
rect 9166 6433 9205 6467
rect 9239 6433 9278 6467
rect 9312 6433 9351 6467
rect 9385 6433 9424 6467
rect 9458 6433 9497 6467
rect 9531 6433 9570 6467
rect 9604 6433 9643 6467
rect 9677 6433 9716 6467
rect 9750 6433 9789 6467
rect 9823 6433 9862 6467
rect 9896 6433 9908 6467
rect 0 6423 9908 6433
rect 0 6395 123 6423
rect 0 6389 68 6395
rect 34 6361 68 6389
rect 102 6389 123 6395
rect 157 6389 191 6423
rect 102 6361 191 6389
rect 34 6355 191 6361
rect 102 6321 191 6355
rect 2061 6389 2129 6423
rect 2163 6389 2198 6423
rect 2232 6389 2267 6423
rect 2301 6389 2336 6423
rect 2370 6389 2405 6423
rect 2439 6389 2474 6423
rect 2508 6389 2543 6423
rect 2577 6389 2612 6423
rect 2646 6389 2681 6423
rect 2715 6389 2750 6423
rect 2784 6389 2819 6423
rect 2853 6389 2888 6423
rect 2922 6389 2957 6423
rect 2991 6389 3026 6423
rect 3060 6389 3095 6423
rect 3129 6389 3164 6423
rect 3198 6389 3233 6423
rect 3267 6389 3302 6423
rect 3336 6389 3371 6423
rect 3405 6389 3440 6423
rect 3474 6389 3509 6423
rect 3543 6389 3578 6423
rect 3612 6389 3647 6423
rect 3681 6389 3716 6423
rect 3750 6389 3785 6423
rect 3819 6389 3854 6423
rect 3888 6389 3923 6423
rect 3957 6389 3992 6423
rect 4026 6389 4061 6423
rect 4095 6389 4130 6423
rect 4164 6389 4199 6423
rect 4233 6389 4268 6423
rect 4302 6389 4337 6423
rect 4371 6389 4406 6423
rect 4440 6389 4475 6423
rect 4509 6389 4544 6423
rect 4578 6389 4613 6423
rect 4647 6389 4682 6423
rect 4716 6389 4751 6423
rect 4785 6389 4820 6423
rect 4854 6389 4889 6423
rect 4923 6389 4958 6423
rect 4992 6389 5027 6423
rect 5061 6389 5096 6423
rect 5130 6389 5165 6423
rect 5199 6389 5234 6423
rect 5268 6389 5303 6423
rect 5337 6389 5372 6423
rect 5406 6389 5441 6423
rect 5475 6389 5510 6423
rect 5544 6389 5579 6423
rect 5613 6389 5648 6423
rect 5682 6389 5717 6423
rect 5751 6389 5786 6423
rect 5820 6389 5855 6423
rect 5889 6389 5924 6423
rect 2061 6355 5924 6389
rect 7658 6389 7794 6423
rect 7658 6355 7726 6389
rect 7760 6355 7794 6389
rect 2061 6321 2129 6355
rect 2163 6321 2198 6355
rect 2232 6321 2267 6355
rect 2301 6321 2336 6355
rect 2370 6321 2405 6355
rect 2439 6321 2474 6355
rect 2508 6321 2543 6355
rect 2577 6321 2612 6355
rect 2646 6321 2681 6355
rect 2715 6321 2750 6355
rect 2784 6321 2819 6355
rect 2853 6321 2888 6355
rect 2922 6321 2957 6355
rect 2991 6321 3026 6355
rect 3060 6321 3095 6355
rect 3129 6321 3164 6355
rect 3198 6321 3233 6355
rect 3267 6321 3302 6355
rect 3336 6321 3371 6355
rect 3405 6321 3440 6355
rect 3474 6321 3509 6355
rect 3543 6321 3578 6355
rect 7692 6321 7794 6355
rect 9732 6389 9766 6423
rect 9800 6389 9908 6423
rect 9732 6355 9874 6389
rect 9732 6321 9806 6355
rect 102 6287 259 6321
rect 170 6253 259 6287
rect 2061 6287 3578 6321
rect 2061 6253 2129 6287
rect 2163 6253 2198 6287
rect 2232 6253 2267 6287
rect 2301 6253 2336 6287
rect 2370 6253 2405 6287
rect 2439 6253 2474 6287
rect 2508 6253 2543 6287
rect 2577 6253 2612 6287
rect 2646 6253 2681 6287
rect 2715 6253 2750 6287
rect 2784 6253 2819 6287
rect 2853 6253 2888 6287
rect 2922 6253 2957 6287
rect 2991 6253 3026 6287
rect 3060 6253 3095 6287
rect 3129 6253 3164 6287
rect 3198 6253 3233 6287
rect 3267 6253 3302 6287
rect 3336 6253 3371 6287
rect 3405 6253 3440 6287
rect 3474 6253 3509 6287
rect 3543 6253 3578 6287
rect 7624 6320 7794 6321
rect 7624 6286 7726 6320
rect 7624 6253 7658 6286
rect 7590 6252 7658 6253
rect 7692 6253 7726 6286
rect 9664 6287 9806 6321
rect 9664 6253 9738 6287
rect 7692 6252 7760 6253
rect 7590 6218 7726 6252
rect 7624 6217 7760 6218
rect 7624 6184 7658 6217
rect 7590 6183 7658 6184
rect 7692 6184 7760 6217
rect 7692 6183 7726 6184
rect 7590 6150 7726 6183
rect 7590 6149 7760 6150
rect 7624 6148 7760 6149
rect 7624 6115 7658 6148
rect 7590 6114 7658 6115
rect 7692 6116 7760 6148
rect 7692 6114 7726 6116
rect 323 6094 395 6100
rect 357 6066 395 6094
rect 429 6066 449 6100
rect 507 6066 517 6100
rect 619 6066 629 6100
rect 687 6066 707 6100
rect 755 6066 784 6100
rect 823 6066 857 6100
rect 891 6066 925 6100
rect 984 6066 993 6100
rect 1095 6066 1104 6100
rect 1163 6066 1181 6100
rect 1231 6066 1258 6100
rect 1299 6066 1333 6100
rect 1369 6066 1401 6100
rect 1446 6066 1469 6100
rect 1522 6066 1537 6100
rect 1598 6066 1605 6100
rect 1639 6066 1640 6100
rect 1707 6066 1741 6100
rect 1775 6066 1806 6100
rect 1843 6066 1877 6100
rect 1917 6066 1945 6100
rect 1994 6066 2013 6100
rect 2071 6066 2081 6100
rect 2148 6066 2149 6100
rect 2183 6066 2191 6100
rect 2251 6066 2268 6100
rect 2319 6066 2344 6100
rect 2387 6066 2420 6100
rect 2455 6066 2489 6100
rect 2530 6066 2557 6100
rect 2591 6066 2625 6100
rect 2659 6066 2662 6100
rect 2727 6066 2739 6100
rect 2795 6066 2816 6100
rect 2863 6066 2893 6100
rect 2931 6066 2965 6100
rect 3004 6066 3033 6100
rect 3081 6066 3101 6100
rect 3158 6066 3169 6100
rect 3234 6066 3237 6100
rect 3271 6066 3276 6100
rect 3339 6066 3352 6100
rect 3407 6066 3441 6100
rect 3475 6066 3509 6100
rect 3552 6066 3577 6100
rect 3629 6066 3645 6100
rect 3705 6066 3713 6100
rect 3815 6066 3823 6100
rect 3883 6066 3899 6100
rect 3951 6066 3975 6100
rect 4019 6066 4051 6100
rect 4087 6066 4121 6100
rect 4161 6066 4189 6100
rect 4237 6066 4257 6100
rect 4291 6066 4325 6100
rect 4359 6066 4379 6100
rect 4427 6066 4455 6100
rect 4495 6066 4529 6100
rect 4565 6066 4597 6100
rect 4641 6066 4665 6100
rect 4717 6066 4733 6100
rect 4793 6066 4801 6100
rect 4835 6094 4987 6100
rect 4937 6066 4987 6094
rect 5023 6066 5057 6100
rect 5095 6066 5125 6100
rect 5169 6066 5193 6100
rect 5243 6066 5261 6100
rect 5317 6066 5329 6100
rect 5391 6066 5397 6100
rect 5499 6066 5505 6100
rect 5567 6066 5579 6100
rect 5635 6066 5652 6100
rect 5703 6066 5725 6100
rect 5771 6066 5798 6100
rect 5839 6066 5871 6100
rect 5907 6066 5941 6100
rect 5978 6066 6009 6100
rect 6051 6066 6077 6100
rect 6124 6066 6145 6100
rect 6197 6066 6213 6100
rect 6270 6066 6281 6100
rect 6343 6066 6349 6100
rect 6416 6066 6417 6100
rect 6451 6066 6455 6100
rect 6519 6066 6528 6100
rect 6587 6066 6601 6100
rect 6655 6066 6674 6100
rect 6723 6066 6747 6100
rect 6791 6066 6820 6100
rect 6859 6066 6893 6100
rect 6927 6066 6961 6100
rect 7000 6066 7029 6100
rect 7073 6066 7097 6100
rect 7146 6066 7165 6100
rect 7219 6066 7233 6100
rect 7292 6066 7301 6100
rect 7365 6066 7369 6100
rect 7403 6094 7437 6100
rect 323 6022 357 6032
rect 323 5950 357 5964
rect 323 5878 357 5896
rect 4937 5998 4949 6032
rect 4937 5930 4949 5964
rect 4937 5862 4949 5896
rect 323 5806 357 5828
rect 730 5825 781 5859
rect 815 5825 866 5859
rect 900 5825 952 5859
rect 986 5825 1038 5859
rect 1586 5825 1637 5859
rect 1671 5825 1722 5859
rect 1756 5825 1808 5859
rect 1842 5825 1894 5859
rect 2196 5825 2212 5859
rect 2246 5825 2286 5859
rect 2320 5825 2360 5859
rect 2394 5825 2408 5859
rect 2468 5825 2493 5859
rect 2542 5825 2578 5859
rect 2615 5825 2654 5859
rect 2698 5825 2727 5859
rect 2784 5825 2800 5859
rect 2834 5825 2873 5859
rect 2907 5825 2946 5859
rect 2980 5825 2996 5859
rect 3052 5825 3068 5859
rect 3102 5825 3138 5859
rect 3172 5825 3208 5859
rect 3242 5825 3264 5859
rect 3312 5825 3347 5859
rect 3383 5825 3416 5859
rect 3468 5825 3485 5859
rect 3519 5825 3520 5859
rect 3588 5825 3606 5859
rect 3657 5825 3692 5859
rect 3726 5825 3761 5859
rect 3795 5825 3830 5859
rect 3864 5825 3899 5859
rect 3933 5825 3968 5859
rect 4002 5825 4037 5859
rect 4071 5825 4106 5859
rect 4154 5825 4175 5859
rect 4239 5825 4244 5859
rect 4278 5825 4290 5859
rect 4347 5825 4376 5859
rect 4416 5825 4451 5859
rect 4496 5825 4520 5859
rect 4554 5825 4589 5859
rect 4623 5825 4658 5859
rect 4692 5825 4708 5859
rect 323 5734 357 5760
rect 4937 5794 4949 5828
rect 323 5662 357 5692
rect 323 5590 357 5624
rect 323 5522 357 5556
rect 323 5454 357 5484
rect 323 5386 357 5412
rect 323 5318 357 5340
rect 323 5250 357 5268
rect 323 5182 357 5196
rect 323 5114 357 5124
rect 323 5046 357 5052
rect 323 4978 357 4980
rect 323 4942 357 4944
rect 323 4870 357 4876
rect 323 4798 357 4808
rect 323 4726 357 4740
rect 323 4654 357 4672
rect 323 4582 357 4604
rect 323 4510 357 4536
rect 323 4438 357 4468
rect 323 4366 357 4400
rect 323 4298 357 4332
rect 323 4230 357 4260
rect 323 4162 357 4188
rect 323 4094 357 4116
rect 323 4026 357 4044
rect 323 3958 357 3971
rect 323 3890 357 3898
rect 323 3822 357 3825
rect 323 3786 357 3788
rect 439 5658 473 5697
rect 439 5585 473 5624
rect 439 5512 473 5551
rect 439 5439 473 5478
rect 439 5366 473 5405
rect 439 5293 473 5332
rect 439 5220 473 5259
rect 439 5147 473 5186
rect 439 5074 473 5113
rect 439 5001 473 5040
rect 439 4928 473 4967
rect 439 4855 473 4894
rect 439 4781 473 4821
rect 439 4707 473 4747
rect 439 4633 473 4673
rect 439 4559 473 4599
rect 439 4485 473 4525
rect 439 4411 473 4451
rect 439 4337 473 4377
rect 439 4263 473 4303
rect 439 4189 473 4229
rect 439 4115 473 4155
rect 439 4041 473 4081
rect 439 3967 473 4007
rect 439 3893 473 3933
rect 439 3819 473 3859
rect 1295 5658 1329 5697
rect 1295 5585 1329 5624
rect 1295 5512 1329 5551
rect 1295 5439 1329 5478
rect 1295 5366 1329 5405
rect 1295 5293 1329 5332
rect 1295 5220 1329 5259
rect 1295 5147 1329 5186
rect 1295 5074 1329 5113
rect 1295 5001 1329 5040
rect 1295 4928 1329 4967
rect 1295 4855 1329 4894
rect 1295 4781 1329 4821
rect 1295 4707 1329 4747
rect 1295 4633 1329 4673
rect 1295 4559 1329 4599
rect 1295 4485 1329 4525
rect 1295 4411 1329 4451
rect 1295 4337 1329 4377
rect 1295 4263 1329 4303
rect 1295 4189 1329 4229
rect 1295 4115 1329 4155
rect 1295 4041 1329 4081
rect 1295 3967 1329 4007
rect 1295 3893 1329 3933
rect 1295 3819 1329 3859
rect 2151 5658 2185 5697
rect 2151 5585 2185 5624
rect 2151 5512 2185 5551
rect 2151 5439 2185 5478
rect 2151 5366 2185 5405
rect 2151 5293 2185 5332
rect 2151 5220 2185 5259
rect 2151 5147 2185 5186
rect 2151 5074 2185 5113
rect 2151 5001 2185 5040
rect 2151 4928 2185 4967
rect 2151 4855 2185 4894
rect 2151 4781 2185 4821
rect 2151 4707 2185 4747
rect 2151 4633 2185 4673
rect 2151 4559 2185 4599
rect 2151 4485 2185 4525
rect 2151 4411 2185 4451
rect 2151 4337 2185 4377
rect 2151 4263 2185 4303
rect 2151 4189 2185 4229
rect 2151 4115 2185 4155
rect 2151 4041 2185 4081
rect 2151 3967 2185 4007
rect 2151 3893 2185 3933
rect 2151 3819 2185 3859
rect 3007 5658 3041 5697
rect 3007 5585 3041 5624
rect 3007 5512 3041 5551
rect 3007 5439 3041 5478
rect 3007 5366 3041 5405
rect 3007 5293 3041 5332
rect 3007 5220 3041 5259
rect 3007 5147 3041 5186
rect 3007 5074 3041 5113
rect 3007 5001 3041 5040
rect 3007 4928 3041 4967
rect 3007 4855 3041 4894
rect 3007 4781 3041 4821
rect 3007 4707 3041 4747
rect 3007 4633 3041 4673
rect 3007 4559 3041 4599
rect 3007 4485 3041 4525
rect 3007 4411 3041 4451
rect 3007 4337 3041 4377
rect 3007 4263 3041 4303
rect 3007 4189 3041 4229
rect 3007 4115 3041 4155
rect 3007 4041 3041 4081
rect 3007 3967 3041 4007
rect 3007 3893 3041 3933
rect 3007 3819 3041 3859
rect 3863 5658 3897 5697
rect 3863 5585 3897 5624
rect 3863 5512 3897 5551
rect 3863 5439 3897 5478
rect 3863 5366 3897 5405
rect 3863 5293 3897 5332
rect 3863 5220 3897 5259
rect 3863 5147 3897 5186
rect 3863 5074 3897 5113
rect 3863 5001 3897 5040
rect 3863 4928 3897 4967
rect 3863 4855 3897 4894
rect 3863 4781 3897 4821
rect 3863 4707 3897 4747
rect 3863 4633 3897 4673
rect 3863 4559 3897 4599
rect 3863 4485 3897 4525
rect 3863 4411 3897 4451
rect 3863 4337 3897 4377
rect 3863 4263 3897 4303
rect 3863 4189 3897 4229
rect 3863 4115 3897 4155
rect 3863 4041 3897 4081
rect 3863 3967 3897 4007
rect 3863 3893 3897 3933
rect 3863 3819 3897 3859
rect 4719 5658 4753 5697
rect 4719 5585 4753 5624
rect 4719 5512 4753 5551
rect 4719 5439 4753 5478
rect 4719 5366 4753 5405
rect 4719 5293 4753 5332
rect 4719 5220 4753 5259
rect 4719 5147 4753 5186
rect 4719 5074 4753 5113
rect 4719 5001 4753 5040
rect 4719 4928 4753 4967
rect 4719 4855 4753 4894
rect 4719 4781 4753 4821
rect 4719 4707 4753 4747
rect 4719 4633 4753 4673
rect 4719 4559 4753 4599
rect 4719 4485 4753 4525
rect 4719 4411 4753 4451
rect 4719 4337 4753 4377
rect 4719 4263 4753 4303
rect 4719 4189 4753 4229
rect 4719 4115 4753 4155
rect 4719 4041 4753 4081
rect 4719 3967 4753 4007
rect 4719 3893 4753 3933
rect 4719 3819 4753 3859
rect 4937 5726 4949 5760
rect 4937 5658 4949 5692
rect 4937 5590 4949 5624
rect 4937 5522 4949 5556
rect 4937 5454 4949 5488
rect 4937 5386 4949 5420
rect 4937 5318 4949 5352
rect 4937 5250 4949 5284
rect 4937 5182 4949 5216
rect 4937 5114 4949 5148
rect 4937 5046 4949 5080
rect 4937 4978 4949 5012
rect 4937 4910 4949 4944
rect 4937 4842 4949 4876
rect 4937 4774 4949 4808
rect 4937 4706 4949 4740
rect 4937 4638 4949 4672
rect 4937 4570 4949 4604
rect 4937 4502 4949 4536
rect 4937 4434 4949 4468
rect 4937 4366 4949 4400
rect 4937 4298 4949 4332
rect 4937 4230 4949 4264
rect 4937 4162 4949 4196
rect 4937 4094 4949 4128
rect 4937 4044 4949 4060
rect 4831 4032 4835 4044
rect 4869 4032 4949 4044
rect 4831 4026 4949 4032
rect 4831 4005 4915 4026
rect 4865 3998 4903 4005
rect 4869 3971 4903 3998
rect 4937 3971 4949 3992
rect 4831 3964 4835 3971
rect 4869 3964 4949 3971
rect 4831 3958 4949 3964
rect 4831 3932 4915 3958
rect 4865 3930 4903 3932
rect 4869 3898 4903 3930
rect 4937 3898 4949 3924
rect 4831 3896 4835 3898
rect 4869 3896 4949 3898
rect 4831 3890 4949 3896
rect 4831 3862 4915 3890
rect 4831 3859 4835 3862
rect 4869 3859 4915 3862
rect 4869 3828 4903 3859
rect 4865 3825 4903 3828
rect 4937 3825 4949 3856
rect 4831 3822 4949 3825
rect 4831 3794 4915 3822
rect 4831 3786 4835 3794
rect 4869 3788 4915 3794
rect 4869 3786 4949 3788
rect 4869 3760 4903 3786
rect 4865 3752 4903 3760
rect 4937 3754 4949 3786
rect 323 3713 357 3720
rect 507 3695 523 3729
rect 557 3695 592 3729
rect 626 3695 661 3729
rect 695 3695 696 3729
rect 764 3695 781 3729
rect 833 3695 866 3729
rect 902 3695 937 3729
rect 986 3695 1006 3729
rect 1072 3695 1075 3729
rect 1109 3695 1143 3729
rect 1177 3695 1211 3729
rect 1245 3695 1261 3729
rect 1364 3695 1380 3729
rect 1414 3695 1449 3729
rect 1483 3695 1518 3729
rect 1586 3695 1587 3729
rect 1621 3695 1637 3729
rect 1690 3695 1722 3729
rect 1759 3695 1794 3729
rect 1842 3695 1863 3729
rect 1928 3695 1931 3729
rect 1965 3695 1999 3729
rect 2033 3695 2067 3729
rect 2101 3695 2117 3729
rect 2442 3695 2493 3729
rect 2527 3695 2578 3729
rect 2612 3695 2664 3729
rect 2698 3695 2750 3729
rect 3075 3695 3091 3729
rect 3125 3695 3160 3729
rect 3194 3695 3229 3729
rect 3263 3695 3264 3729
rect 3332 3695 3349 3729
rect 3401 3695 3434 3729
rect 3470 3695 3505 3729
rect 3554 3695 3574 3729
rect 3640 3695 3643 3729
rect 3677 3695 3711 3729
rect 3745 3695 3779 3729
rect 3813 3695 3829 3729
rect 3931 3695 3947 3729
rect 3981 3695 4016 3729
rect 4050 3695 4085 3729
rect 4119 3695 4120 3729
rect 4188 3695 4205 3729
rect 4257 3695 4290 3729
rect 4326 3695 4361 3729
rect 4410 3695 4430 3729
rect 4496 3695 4499 3729
rect 4533 3695 4567 3729
rect 4601 3695 4635 3729
rect 4669 3695 4685 3729
rect 4831 3726 4915 3752
rect 4831 3713 4835 3726
rect 4869 3720 4915 3726
rect 4869 3713 4949 3720
rect 323 3640 357 3652
rect 323 3567 357 3584
rect 323 3494 357 3533
rect 4869 3692 4903 3713
rect 4865 3679 4903 3692
rect 4937 3686 4949 3713
rect 4831 3658 4915 3679
rect 4831 3640 4835 3658
rect 4869 3652 4915 3658
rect 4869 3640 4949 3652
rect 4869 3624 4903 3640
rect 4865 3606 4903 3624
rect 4937 3618 4949 3640
rect 4831 3590 4915 3606
rect 4831 3567 4835 3590
rect 4869 3584 4915 3590
rect 4869 3567 4949 3584
rect 4869 3556 4903 3567
rect 4865 3533 4903 3556
rect 4937 3533 4949 3567
rect 4831 3522 4949 3533
rect 4831 3494 4835 3522
rect 4869 3494 4949 3522
rect 4869 3488 4903 3494
rect 323 3454 357 3460
rect 391 3454 395 3488
rect 459 3454 468 3488
rect 527 3454 541 3488
rect 595 3454 614 3488
rect 663 3454 687 3488
rect 731 3454 760 3488
rect 799 3454 833 3488
rect 867 3454 901 3488
rect 940 3454 969 3488
rect 1013 3454 1037 3488
rect 1086 3454 1105 3488
rect 1159 3454 1173 3488
rect 1232 3454 1241 3488
rect 1305 3454 1309 3488
rect 1343 3454 1344 3488
rect 1411 3454 1417 3488
rect 1479 3454 1490 3488
rect 1547 3454 1563 3488
rect 1615 3454 1636 3488
rect 1683 3454 1709 3488
rect 1751 3454 1782 3488
rect 1819 3454 1853 3488
rect 1889 3454 1921 3488
rect 1962 3454 1989 3488
rect 2035 3454 2057 3488
rect 2108 3454 2125 3488
rect 2181 3454 2193 3488
rect 2254 3454 2261 3488
rect 2327 3454 2329 3488
rect 2363 3454 2366 3488
rect 2431 3454 2439 3488
rect 2499 3454 2512 3488
rect 2567 3454 2585 3488
rect 2635 3454 2658 3488
rect 2703 3454 2731 3488
rect 2771 3454 2804 3488
rect 2839 3454 2873 3488
rect 2911 3454 2941 3488
rect 2984 3454 3009 3488
rect 3057 3454 3077 3488
rect 3130 3454 3145 3488
rect 3203 3454 3213 3488
rect 3276 3454 3281 3488
rect 3383 3454 3388 3488
rect 3451 3454 3461 3488
rect 3519 3454 3534 3488
rect 3587 3454 3607 3488
rect 3655 3454 3679 3488
rect 3723 3454 3751 3488
rect 3791 3454 3823 3488
rect 3859 3454 3893 3488
rect 3929 3454 3961 3488
rect 4001 3454 4029 3488
rect 4073 3454 4097 3488
rect 4145 3454 4165 3488
rect 4217 3454 4233 3488
rect 4289 3454 4301 3488
rect 4361 3454 4369 3488
rect 4433 3454 4437 3488
rect 4539 3454 4543 3488
rect 4607 3454 4615 3488
rect 4675 3454 4687 3488
rect 4743 3454 4759 3488
rect 4793 3460 4831 3488
rect 4865 3460 4903 3488
rect 4937 3460 4949 3494
rect 6561 6028 6595 6066
rect 6561 5990 6595 5994
rect 6561 5955 6595 5956
rect 6561 5882 6595 5888
rect 7403 6018 7437 6060
rect 7590 6082 7726 6114
rect 7590 6080 7760 6082
rect 7624 6079 7760 6080
rect 7624 6046 7658 6079
rect 7590 6045 7658 6046
rect 7692 6048 7760 6079
rect 7692 6045 7726 6048
rect 7590 6014 7726 6045
rect 7590 6011 7760 6014
rect 7624 6010 7760 6011
rect 7403 5970 7437 5984
rect 7403 5902 7437 5908
rect 6561 5809 6595 5820
rect 6561 5736 6595 5752
rect 6561 5663 6595 5684
rect 6561 5590 6595 5616
rect 6561 5517 6595 5548
rect 6561 5446 6595 5480
rect 6561 5378 6595 5409
rect 6561 5310 6595 5335
rect 6561 5242 6595 5261
rect 6561 5174 6595 5187
rect 6561 5106 6595 5113
rect 6561 5038 6595 5039
rect 6561 4999 6595 5004
rect 6561 4925 6595 4936
rect 6561 4851 6595 4868
rect 6561 4777 6595 4800
rect 6561 4703 6595 4732
rect 6561 4630 6595 4664
rect 6561 4562 6595 4595
rect 6561 4494 6595 4521
rect 6561 4426 6595 4447
rect 6561 4357 6595 4373
rect 6561 4288 6595 4299
rect 6561 4219 6595 4225
rect 6561 4150 6595 4151
rect 6561 4111 6595 4116
rect 6561 4037 6595 4047
rect 6561 3963 6595 3978
rect 6705 5810 6739 5848
rect 6705 5738 6739 5776
rect 6705 5666 6739 5704
rect 6705 5594 6739 5632
rect 6705 5522 6739 5560
rect 6705 5450 6739 5488
rect 6705 5378 6739 5416
rect 6705 5306 6739 5344
rect 6705 5234 6739 5272
rect 6705 5162 6739 5200
rect 6705 5090 6739 5128
rect 6705 5018 6739 5056
rect 6705 4946 6739 4984
rect 6705 4874 6739 4912
rect 6705 4802 6739 4840
rect 6705 4730 6739 4768
rect 6705 4658 6739 4696
rect 6705 4586 6739 4624
rect 6705 4514 6739 4552
rect 6705 4442 6739 4480
rect 6705 4370 6739 4408
rect 6705 4298 6739 4336
rect 6705 4226 6739 4264
rect 6705 4154 6739 4192
rect 6705 4082 6739 4120
rect 6941 5809 6975 5848
rect 6941 5736 6975 5775
rect 6941 5663 6975 5702
rect 6941 5590 6975 5629
rect 6941 5517 6975 5556
rect 6941 5444 6975 5483
rect 6941 5371 6975 5410
rect 6941 5298 6975 5337
rect 6941 5225 6975 5264
rect 6941 5152 6975 5191
rect 6941 5079 6975 5118
rect 6941 5006 6975 5045
rect 6941 4933 6975 4972
rect 6941 4860 6975 4899
rect 6941 4787 6975 4826
rect 6941 4714 6975 4753
rect 6941 4641 6975 4680
rect 6941 4568 6975 4607
rect 6941 4495 6975 4534
rect 6941 4422 6975 4461
rect 6941 4349 6975 4388
rect 6941 4276 6975 4315
rect 6941 4203 6975 4242
rect 6941 4130 6975 4169
rect 7051 5809 7085 5848
rect 7051 5736 7085 5775
rect 7051 5663 7085 5702
rect 7051 5590 7085 5629
rect 7051 5517 7085 5556
rect 7051 5444 7085 5483
rect 7051 5371 7085 5410
rect 7051 5298 7085 5337
rect 7051 5225 7085 5264
rect 7051 5152 7085 5191
rect 7051 5079 7085 5118
rect 7051 5006 7085 5045
rect 7051 4933 7085 4972
rect 7051 4860 7085 4899
rect 7051 4787 7085 4826
rect 7051 4714 7085 4753
rect 7051 4641 7085 4680
rect 7051 4568 7085 4607
rect 7051 4495 7085 4534
rect 7051 4422 7085 4461
rect 7051 4349 7085 4388
rect 7051 4276 7085 4315
rect 7051 4203 7085 4242
rect 7051 4130 7085 4169
rect 7287 5809 7321 5848
rect 7287 5736 7321 5775
rect 7287 5663 7321 5702
rect 7287 5590 7321 5629
rect 7287 5517 7321 5556
rect 7287 5444 7321 5483
rect 7287 5371 7321 5410
rect 7287 5298 7321 5337
rect 7287 5225 7321 5264
rect 7287 5152 7321 5191
rect 7287 5079 7321 5118
rect 7287 5006 7321 5045
rect 7287 4933 7321 4972
rect 7287 4860 7321 4899
rect 7287 4787 7321 4826
rect 7287 4714 7321 4753
rect 7287 4641 7321 4680
rect 7287 4568 7321 4607
rect 7287 4495 7321 4534
rect 7287 4422 7321 4461
rect 7287 4349 7321 4388
rect 7287 4276 7321 4315
rect 7287 4203 7321 4242
rect 7287 4130 7321 4169
rect 7403 5866 7437 5868
rect 7403 5790 7437 5800
rect 7403 5714 7437 5732
rect 7403 5638 7437 5664
rect 7403 5562 7437 5596
rect 7403 5494 7437 5528
rect 7403 5426 7437 5452
rect 7403 5358 7437 5376
rect 7403 5290 7437 5300
rect 7403 5222 7437 5224
rect 7403 5182 7437 5188
rect 7403 5106 7437 5120
rect 7403 5029 7437 5052
rect 7403 4952 7437 4984
rect 7624 5977 7658 6010
rect 7692 6008 7760 6010
rect 7913 6107 7925 6141
rect 7959 6107 7998 6141
rect 8032 6107 8071 6141
rect 8105 6107 8144 6141
rect 8178 6107 8217 6141
rect 8251 6107 8290 6141
rect 8324 6107 8363 6141
rect 8397 6107 8436 6141
rect 8470 6107 8509 6141
rect 8543 6107 8582 6141
rect 8616 6107 8655 6141
rect 8689 6107 8728 6141
rect 8762 6107 8801 6141
rect 8835 6107 8874 6141
rect 8908 6107 8947 6141
rect 8981 6107 9021 6141
rect 9055 6107 9095 6141
rect 9129 6107 9169 6141
rect 9203 6107 9243 6141
rect 9277 6107 9317 6141
rect 9351 6107 9391 6141
rect 9425 6107 9465 6141
rect 9499 6107 9539 6141
rect 9573 6107 9585 6141
rect 7913 6100 9585 6107
rect 7913 6069 7997 6100
rect 7947 6066 7997 6069
rect 8031 6066 8065 6100
rect 8099 6066 8133 6100
rect 8167 6066 8201 6100
rect 8235 6066 8269 6100
rect 8303 6066 8337 6100
rect 8371 6066 8405 6100
rect 8439 6066 8473 6100
rect 8507 6066 8541 6100
rect 8575 6066 8701 6100
rect 8735 6066 8769 6100
rect 8803 6066 8837 6100
rect 8871 6066 8905 6100
rect 8939 6066 8973 6100
rect 9007 6066 9041 6100
rect 9075 6066 9109 6100
rect 9143 6066 9177 6100
rect 9211 6066 9245 6100
rect 9279 6066 9313 6100
rect 9347 6066 9381 6100
rect 9415 6066 9449 6100
rect 9483 6066 9517 6100
rect 7623 5976 7658 5977
rect 7695 5980 7733 6008
rect 7623 5974 7661 5976
rect 7695 5974 7726 5980
rect 7589 5946 7726 5974
rect 7760 5946 7767 5974
rect 7589 5942 7767 5946
rect 7589 5932 7590 5942
rect 7624 5941 7767 5942
rect 7624 5908 7658 5941
rect 7692 5932 7767 5941
rect 7623 5907 7658 5908
rect 7695 5912 7733 5932
rect 7623 5898 7661 5907
rect 7695 5898 7726 5912
rect 7589 5878 7726 5898
rect 7760 5878 7767 5898
rect 7589 5873 7767 5878
rect 7589 5856 7590 5873
rect 7624 5872 7767 5873
rect 7624 5839 7658 5872
rect 7692 5856 7767 5872
rect 7623 5838 7658 5839
rect 7695 5844 7733 5856
rect 7623 5822 7661 5838
rect 7695 5822 7726 5844
rect 7589 5810 7726 5822
rect 7760 5810 7767 5822
rect 7589 5804 7767 5810
rect 7589 5780 7590 5804
rect 7624 5803 7767 5804
rect 7624 5770 7658 5803
rect 7692 5780 7767 5803
rect 7623 5769 7658 5770
rect 7695 5776 7733 5780
rect 7623 5746 7661 5769
rect 7695 5746 7726 5776
rect 7589 5742 7726 5746
rect 7760 5742 7767 5746
rect 7589 5735 7767 5742
rect 7589 5704 7590 5735
rect 7624 5734 7767 5735
rect 7624 5701 7658 5734
rect 7692 5708 7767 5734
rect 7692 5704 7726 5708
rect 7760 5704 7767 5708
rect 7623 5700 7658 5701
rect 7623 5670 7661 5700
rect 7695 5674 7726 5704
rect 7695 5670 7733 5674
rect 7589 5666 7767 5670
rect 7589 5632 7590 5666
rect 7624 5665 7767 5666
rect 7624 5632 7658 5665
rect 7589 5631 7658 5632
rect 7692 5640 7767 5665
rect 7692 5631 7726 5640
rect 7589 5628 7726 5631
rect 7760 5628 7767 5640
rect 7623 5597 7661 5628
rect 7624 5596 7661 5597
rect 7695 5606 7726 5628
rect 7589 5563 7590 5594
rect 7624 5563 7658 5596
rect 7695 5594 7733 5606
rect 7589 5562 7658 5563
rect 7692 5572 7767 5594
rect 7692 5562 7726 5572
rect 7589 5552 7726 5562
rect 7760 5552 7767 5572
rect 7623 5528 7661 5552
rect 7624 5527 7661 5528
rect 7695 5538 7726 5552
rect 7589 5494 7590 5518
rect 7624 5494 7658 5527
rect 7695 5518 7733 5538
rect 7589 5493 7658 5494
rect 7692 5504 7767 5518
rect 7692 5493 7726 5504
rect 7589 5477 7726 5493
rect 7760 5477 7767 5504
rect 7623 5459 7661 5477
rect 7624 5458 7661 5459
rect 7695 5470 7726 5477
rect 7589 5425 7590 5443
rect 7624 5425 7658 5458
rect 7695 5443 7733 5470
rect 7589 5424 7658 5425
rect 7692 5436 7767 5443
rect 7692 5424 7726 5436
rect 7589 5402 7726 5424
rect 7760 5402 7767 5436
rect 7623 5390 7661 5402
rect 7624 5389 7661 5390
rect 7589 5356 7590 5368
rect 7624 5356 7658 5389
rect 7695 5368 7733 5402
rect 7589 5355 7658 5356
rect 7692 5355 7726 5368
rect 7589 5334 7726 5355
rect 7760 5334 7767 5368
rect 7589 5327 7767 5334
rect 7623 5321 7661 5327
rect 7624 5320 7661 5321
rect 7589 5287 7590 5293
rect 7624 5287 7658 5320
rect 7695 5300 7733 5327
rect 7695 5293 7726 5300
rect 7589 5286 7658 5287
rect 7692 5286 7726 5293
rect 7589 5266 7726 5286
rect 7760 5266 7767 5293
rect 7589 5252 7767 5266
rect 7624 5251 7661 5252
rect 7624 5218 7658 5251
rect 7695 5232 7733 5252
rect 7695 5218 7726 5232
rect 7589 5217 7658 5218
rect 7692 5217 7726 5218
rect 7589 5198 7726 5217
rect 7760 5198 7767 5218
rect 7589 5183 7767 5198
rect 7589 5177 7590 5183
rect 7624 5182 7767 5183
rect 7624 5149 7658 5182
rect 7692 5177 7767 5182
rect 7623 5148 7658 5149
rect 7695 5164 7733 5177
rect 7623 5143 7661 5148
rect 7695 5143 7726 5164
rect 7589 5130 7726 5143
rect 7760 5130 7767 5143
rect 7589 5114 7767 5130
rect 7589 5102 7590 5114
rect 7624 5113 7767 5114
rect 7624 5080 7658 5113
rect 7692 5102 7767 5113
rect 7623 5079 7658 5080
rect 7695 5096 7733 5102
rect 7623 5068 7661 5079
rect 7695 5068 7726 5096
rect 7589 5062 7726 5068
rect 7760 5062 7767 5068
rect 7589 5045 7767 5062
rect 7589 5027 7590 5045
rect 7624 5044 7767 5045
rect 7624 5011 7658 5044
rect 7692 5028 7767 5044
rect 7692 5027 7726 5028
rect 7760 5027 7767 5028
rect 7623 5010 7658 5011
rect 7623 4993 7661 5010
rect 7695 4994 7726 5027
rect 7695 4993 7733 4994
rect 7589 4976 7767 4993
rect 7589 4952 7590 4976
rect 7624 4975 7767 4976
rect 7624 4942 7658 4975
rect 7692 4960 7767 4975
rect 7692 4952 7726 4960
rect 7760 4952 7767 4960
rect 7623 4941 7658 4942
rect 7623 4918 7661 4941
rect 7695 4926 7726 4952
rect 7695 4918 7733 4926
rect 7913 5998 7947 6032
rect 9551 6005 9585 6100
rect 7913 5930 7947 5959
rect 7913 5862 7947 5883
rect 7913 5794 7947 5807
rect 7913 5726 7947 5731
rect 7913 5689 7947 5692
rect 7913 5613 7947 5624
rect 7913 5536 7947 5556
rect 7913 5459 7947 5488
rect 7913 5386 7947 5420
rect 7913 5318 7947 5348
rect 8015 5950 8027 5984
rect 8061 5950 8104 5984
rect 8138 5950 8181 5984
rect 8215 5950 8259 5984
rect 8015 5672 8049 5950
rect 8777 5937 8811 5953
rect 8967 5950 9013 5984
rect 9047 5950 9093 5984
rect 9127 5950 9174 5984
rect 9208 5950 9255 5984
rect 9289 5950 9336 5984
rect 9370 5950 9417 5984
rect 9551 5937 9585 5971
rect 8811 5873 8849 5907
rect 8777 5869 8811 5873
rect 8129 5794 8175 5828
rect 8209 5794 8255 5828
rect 8289 5794 8336 5828
rect 8370 5794 8417 5828
rect 8451 5794 8498 5828
rect 8532 5794 8579 5828
rect 8777 5801 8811 5835
rect 9551 5869 9585 5903
rect 8967 5794 9014 5828
rect 9048 5794 9095 5828
rect 9129 5794 9177 5828
rect 9211 5794 9259 5828
rect 9293 5794 9341 5828
rect 9375 5794 9423 5828
rect 9551 5801 9585 5835
rect 8777 5733 8811 5767
rect 8777 5683 8811 5699
rect 9551 5733 9585 5767
rect 8015 5638 8027 5672
rect 8061 5638 8107 5672
rect 8141 5638 8187 5672
rect 8221 5638 8268 5672
rect 8302 5638 8349 5672
rect 8898 5638 8943 5672
rect 8977 5638 9023 5672
rect 9057 5638 9103 5672
rect 9137 5638 9183 5672
rect 9217 5638 9263 5672
rect 9297 5638 9343 5672
rect 9377 5638 9423 5672
rect 9551 5665 9585 5699
rect 8015 5360 8049 5638
rect 9551 5597 9585 5631
rect 8129 5482 8175 5516
rect 8209 5482 8255 5516
rect 8289 5482 8336 5516
rect 8370 5482 8417 5516
rect 8451 5482 8498 5516
rect 8532 5482 8579 5516
rect 8669 5515 8811 5531
rect 8901 5528 8946 5562
rect 8980 5528 9025 5562
rect 9059 5528 9104 5562
rect 9138 5528 9183 5562
rect 9217 5528 9263 5562
rect 9297 5528 9343 5562
rect 9377 5528 9423 5562
rect 9551 5529 9585 5563
rect 8669 5484 8777 5515
rect 8669 5450 8681 5484
rect 8715 5450 8753 5484
rect 8787 5450 8811 5481
rect 8669 5447 8811 5450
rect 8669 5413 8777 5447
rect 8669 5397 8811 5413
rect 9551 5461 9585 5495
rect 9551 5393 9585 5427
rect 8015 5326 8027 5360
rect 8061 5326 8105 5360
rect 8139 5326 8184 5360
rect 8218 5326 8263 5360
rect 8297 5326 8342 5360
rect 8376 5326 8421 5360
rect 8455 5326 8500 5360
rect 8534 5326 8579 5360
rect 8896 5352 8937 5386
rect 8971 5352 9012 5386
rect 9046 5352 9087 5386
rect 9121 5352 9162 5386
rect 9196 5352 9237 5386
rect 9271 5352 9312 5386
rect 9346 5352 9387 5386
rect 9421 5352 9463 5386
rect 9497 5352 9539 5386
rect 9573 5352 9585 5359
rect 7913 5250 7947 5271
rect 9551 5325 9585 5352
rect 9551 5257 9585 5291
rect 8063 5216 8104 5250
rect 8138 5216 8179 5250
rect 8213 5216 8254 5250
rect 8288 5216 8330 5250
rect 8364 5216 8406 5250
rect 8440 5216 8482 5250
rect 10498 6378 10510 6412
rect 10544 6378 10584 6412
rect 10651 6378 10658 6412
rect 10719 6378 10732 6412
rect 10787 6378 10806 6412
rect 10855 6378 10880 6412
rect 10923 6378 10954 6412
rect 10991 6378 11025 6412
rect 11062 6378 11093 6412
rect 11136 6378 11161 6412
rect 11210 6378 11229 6412
rect 11284 6378 11297 6412
rect 11358 6378 11365 6412
rect 11432 6378 11472 6412
rect 11514 6378 11546 6412
rect 11582 6378 11616 6412
rect 11654 6378 11684 6412
rect 11728 6378 11752 6412
rect 11802 6378 11820 6412
rect 11876 6378 11888 6412
rect 11950 6378 11956 6412
rect 12058 6378 12064 6412
rect 12126 6378 12138 6412
rect 12194 6378 12212 6412
rect 12262 6378 12286 6412
rect 12330 6378 12360 6412
rect 12398 6378 12432 6412
rect 12468 6378 12500 6412
rect 12542 6378 12568 6412
rect 12615 6378 12636 6412
rect 12688 6378 12704 6412
rect 12761 6378 12772 6412
rect 12834 6378 12840 6412
rect 12907 6378 12908 6412
rect 12942 6378 12946 6412
rect 13010 6378 13019 6412
rect 13078 6378 13092 6412
rect 13146 6378 13165 6412
rect 13199 6378 13238 6412
rect 13292 6378 13311 6412
rect 13360 6378 13384 6412
rect 13428 6378 13462 6412
rect 10498 6310 10532 6344
rect 13496 6374 13530 6412
rect 10498 6242 10532 6276
rect 10659 6243 10675 6277
rect 10741 6243 10743 6277
rect 10777 6243 10779 6277
rect 10845 6243 10879 6277
rect 10913 6243 10947 6277
rect 10981 6243 10997 6277
rect 10498 6174 10532 6208
rect 13496 6328 13530 6340
rect 12008 6277 12050 6311
rect 13134 6277 13172 6280
rect 12013 6243 12051 6277
rect 12568 6243 12580 6277
rect 12618 6243 12652 6277
rect 12686 6243 12702 6277
rect 11046 6199 11080 6232
rect 11290 6192 11396 6243
rect 11324 6158 11362 6192
rect 10498 6106 10532 6140
rect 10498 6038 10532 6072
rect 10498 5970 10532 6004
rect 10498 5902 10532 5936
rect 10870 6024 10904 6062
rect 10870 5952 10904 5990
rect 11222 6024 11256 6062
rect 11222 5952 11256 5990
rect 10498 5834 10532 5868
rect 10498 5766 10532 5800
rect 10498 5698 10532 5732
rect 11588 5720 11622 5758
rect 11940 5720 11974 5758
rect 10498 5630 10532 5664
rect 10614 5618 10648 5657
rect 10870 5623 10904 5657
rect 11222 5623 11256 5657
rect 10498 5562 10532 5596
rect 10870 5589 11256 5623
rect 11764 5646 11798 5684
rect 10498 5494 10532 5528
rect 12008 5511 12050 6243
rect 13080 6243 13096 6277
rect 13134 6246 13164 6277
rect 13206 6246 13214 6277
rect 13130 6243 13164 6246
rect 13198 6243 13214 6246
rect 13496 6260 13530 6266
rect 13496 6152 13530 6158
rect 13496 6078 13530 6090
rect 12713 5983 12747 6021
rect 12713 5911 12747 5949
rect 12713 5839 12747 5877
rect 12292 5720 12326 5758
rect 12378 5720 12412 5758
rect 12713 5767 12747 5805
rect 13225 5983 13259 6021
rect 13225 5911 13259 5949
rect 13225 5839 13259 5877
rect 13225 5767 13259 5805
rect 13496 6005 13530 6022
rect 13496 5932 13530 5954
rect 13496 5859 13530 5886
rect 13496 5786 13530 5818
rect 12116 5646 12150 5684
rect 12378 5597 12412 5686
rect 13496 5716 13530 5750
rect 12286 5563 12412 5597
rect 12286 5511 12320 5563
rect 12537 5511 12571 5663
rect 12969 5511 13003 5657
rect 13496 5640 13530 5679
rect 13496 5597 13530 5606
rect 13496 5529 13530 5533
rect 12003 5477 12019 5511
rect 12053 5477 12087 5511
rect 12121 5477 12137 5511
rect 12186 5477 12202 5511
rect 12236 5477 12270 5511
rect 12304 5477 12320 5511
rect 12369 5478 12385 5511
rect 10498 5426 10532 5460
rect 12369 5444 12381 5478
rect 12419 5477 12453 5511
rect 12487 5477 12521 5511
rect 12555 5477 12571 5511
rect 12415 5444 12453 5477
rect 12487 5444 12571 5477
rect 13496 5494 13530 5495
rect 12852 5426 13238 5435
rect 10498 5358 10532 5392
rect 10498 5290 10532 5324
rect 7913 5182 7947 5194
rect 8634 5189 8672 5210
rect 8634 5176 8669 5189
rect 8927 5176 8974 5210
rect 9008 5176 9055 5210
rect 9089 5176 9136 5210
rect 9170 5176 9217 5210
rect 9251 5176 9297 5210
rect 9331 5176 9377 5210
rect 9551 5189 9585 5192
rect 7913 5114 7947 5117
rect 7913 5074 7947 5080
rect 8669 5121 8703 5155
rect 9551 5150 9585 5155
rect 8669 5071 8703 5087
rect 8896 5066 8941 5100
rect 8975 5066 9021 5100
rect 9055 5066 9101 5100
rect 9135 5066 9181 5100
rect 9215 5066 9261 5100
rect 9295 5066 9341 5100
rect 9375 5066 9421 5100
rect 9551 5073 9585 5087
rect 7913 4997 7947 5012
rect 9551 4996 9585 5019
rect 7947 4960 8029 4994
rect 8063 4960 8111 4994
rect 8145 4960 8192 4994
rect 8226 4960 8273 4994
rect 8307 4960 8354 4994
rect 8388 4960 8435 4994
rect 7403 4882 7437 4916
rect 7403 4814 7437 4848
rect 7403 4746 7437 4780
rect 7403 4708 7437 4712
rect 7403 4636 7437 4644
rect 7590 4907 7760 4918
rect 7624 4906 7760 4907
rect 7624 4873 7658 4906
rect 7590 4872 7658 4873
rect 7692 4892 7760 4906
rect 7692 4872 7726 4892
rect 7590 4858 7726 4872
rect 7590 4838 7760 4858
rect 7624 4837 7760 4838
rect 7624 4804 7658 4837
rect 7590 4803 7658 4804
rect 7692 4824 7760 4837
rect 7692 4803 7726 4824
rect 7590 4790 7726 4803
rect 7590 4769 7760 4790
rect 7624 4768 7760 4769
rect 7624 4735 7658 4768
rect 7590 4734 7658 4735
rect 7692 4756 7760 4768
rect 7692 4734 7726 4756
rect 7590 4722 7726 4734
rect 7590 4700 7760 4722
rect 7624 4699 7760 4700
rect 7624 4666 7658 4699
rect 7590 4665 7658 4666
rect 7692 4688 7760 4699
rect 7692 4665 7726 4688
rect 7590 4654 7726 4665
rect 7590 4634 7760 4654
rect 7913 4910 7947 4944
rect 8669 4933 8703 4949
rect 9551 4924 9585 4951
rect 8619 4887 8657 4921
rect 8691 4887 8703 4899
rect 8901 4890 8942 4924
rect 8976 4890 9017 4924
rect 9051 4890 9092 4924
rect 9126 4890 9167 4924
rect 9201 4890 9242 4924
rect 9276 4890 9317 4924
rect 9351 4890 9391 4924
rect 9425 4890 9465 4924
rect 9499 4890 9539 4924
rect 9573 4917 9585 4924
rect 9734 5151 9738 5192
rect 9908 5151 9912 5192
rect 9734 5076 9738 5117
rect 9908 5076 9912 5117
rect 9734 5001 9738 5042
rect 9908 5001 9912 5042
rect 9734 4927 9738 4967
rect 9908 4927 9912 4967
rect 10498 5222 10532 5256
rect 10770 5287 10804 5336
rect 10498 5154 10532 5188
rect 10498 5086 10532 5120
rect 10498 5018 10532 5052
rect 10498 4950 10532 4984
rect 7913 4842 7947 4876
rect 8669 4865 8703 4887
rect 7913 4774 7947 4808
rect 8063 4784 8111 4818
rect 8145 4784 8192 4818
rect 8226 4784 8273 4818
rect 8307 4784 8354 4818
rect 8388 4784 8435 4818
rect 8669 4815 8703 4831
rect 9551 4849 9585 4883
rect 9551 4781 9585 4815
rect 7913 4708 7947 4740
rect 8749 4714 8787 4748
rect 8952 4714 8991 4748
rect 9025 4714 9063 4748
rect 9097 4714 9135 4748
rect 9169 4714 9207 4748
rect 9241 4714 9279 4748
rect 9313 4714 9351 4748
rect 9551 4745 9585 4747
rect 10498 4882 10532 4916
rect 10498 4814 10532 4848
rect 10614 5129 10648 5178
rect 10614 5045 10648 5095
rect 10614 4961 10648 5011
rect 10770 5203 10804 5253
rect 11082 5287 11116 5336
rect 10770 5119 10804 5169
rect 10770 5035 10804 5085
rect 10926 5129 10960 5178
rect 10926 5045 10960 5095
rect 10614 4877 10648 4927
rect 10926 4961 10960 5011
rect 11082 5203 11116 5253
rect 11394 5287 11428 5336
rect 11082 5119 11116 5169
rect 11082 5035 11116 5085
rect 11238 5129 11272 5178
rect 11238 5045 11272 5095
rect 10926 4877 10960 4927
rect 11238 4961 11272 5011
rect 11394 5203 11428 5253
rect 11706 5287 11740 5336
rect 11394 5119 11428 5169
rect 11394 5035 11428 5085
rect 11550 5129 11584 5178
rect 11550 5045 11584 5095
rect 11238 4877 11272 4927
rect 11550 4961 11584 5011
rect 11706 5203 11740 5253
rect 11706 5119 11740 5169
rect 11706 5035 11740 5085
rect 11862 5288 11896 5336
rect 11862 5206 11896 5254
rect 11862 5124 11896 5172
rect 11862 5042 11896 5090
rect 11550 4877 11584 4927
rect 11862 4960 11896 5008
rect 11862 4877 11896 4926
rect 11972 5275 12006 5321
rect 11972 5195 12006 5241
rect 11972 5114 12006 5161
rect 11972 5033 12006 5080
rect 11972 4952 12006 4999
rect 11972 4871 12006 4918
rect 12324 5276 12358 5321
rect 12324 5197 12358 5242
rect 12324 5117 12358 5163
rect 12324 5037 12358 5083
rect 12324 4957 12358 5003
rect 12500 5324 12534 5362
rect 12886 5401 13205 5426
rect 12500 5252 12534 5290
rect 12500 5180 12534 5218
rect 12500 5108 12534 5146
rect 12500 5035 12534 5074
rect 12676 5276 12710 5321
rect 12676 5197 12710 5242
rect 12676 5117 12710 5163
rect 12676 5037 12710 5083
rect 12324 4877 12358 4923
rect 12676 4957 12710 5003
rect 12852 5348 12886 5392
rect 13204 5392 13205 5401
rect 13204 5367 13239 5392
rect 12852 5270 12886 5314
rect 12852 5192 12886 5236
rect 12852 5114 12886 5158
rect 12852 5035 12886 5080
rect 13028 5276 13062 5321
rect 13028 5197 13062 5242
rect 13028 5117 13062 5163
rect 13028 5037 13062 5083
rect 12676 4877 12710 4923
rect 13028 4957 13062 5003
rect 13205 5348 13239 5367
rect 13496 5421 13530 5427
rect 13205 5270 13239 5314
rect 13205 5192 13239 5236
rect 13205 5114 13239 5158
rect 13205 5035 13239 5080
rect 13380 5276 13414 5321
rect 13380 5197 13414 5242
rect 13380 5117 13414 5163
rect 13380 5037 13414 5083
rect 13028 4877 13062 4923
rect 13380 4957 13414 5003
rect 13380 4877 13414 4923
rect 13496 5348 13530 5359
rect 13496 5275 13530 5291
rect 13496 5202 13530 5223
rect 13496 5129 13530 5155
rect 13496 5056 13530 5087
rect 13496 4985 13530 5019
rect 13496 4917 13530 4949
rect 13496 4849 13530 4876
rect 10498 4746 10532 4780
rect 10770 4791 10804 4825
rect 11082 4791 11116 4825
rect 11394 4791 11428 4825
rect 11706 4791 11740 4825
rect 10770 4757 11740 4791
rect 13496 4781 13530 4803
rect 7913 4642 7947 4672
rect 9551 4658 9585 4679
rect 7913 4638 8029 4642
rect 7403 4564 7437 4576
rect 7403 4492 7437 4508
rect 7403 4420 7437 4440
rect 7403 4348 7437 4372
rect 7403 4276 7437 4304
rect 7403 4203 7437 4236
rect 7403 4134 7437 4168
rect 7947 4608 8029 4638
rect 8063 4608 8110 4642
rect 8144 4608 8191 4642
rect 8225 4608 8272 4642
rect 8306 4608 8353 4642
rect 8387 4608 8433 4642
rect 8467 4608 8513 4642
rect 7913 4570 7947 4602
rect 7913 4502 7947 4530
rect 7913 4434 7947 4458
rect 8669 4581 8703 4597
rect 9551 4577 9585 4611
rect 8669 4513 8703 4547
rect 8777 4538 8855 4572
rect 8901 4538 8948 4572
rect 8982 4538 9029 4572
rect 9063 4538 9110 4572
rect 9144 4538 9191 4572
rect 9225 4538 9271 4572
rect 9305 4538 9351 4572
rect 8777 4511 8811 4538
rect 8669 4451 8674 4479
rect 8669 4445 8708 4451
rect 8703 4413 8708 4445
rect 7913 4366 7947 4386
rect 8063 4352 8104 4386
rect 8138 4352 8179 4386
rect 8213 4352 8254 4386
rect 8288 4352 8328 4386
rect 8362 4352 8402 4386
rect 8436 4352 8476 4386
rect 8510 4352 8550 4386
rect 8669 4379 8674 4411
rect 8777 4443 8811 4477
rect 9734 4658 9738 4711
rect 9908 4658 9912 4711
rect 9734 4571 9738 4624
rect 9908 4571 9912 4624
rect 10498 4678 10532 4712
rect 13496 4713 13530 4730
rect 10498 4610 10532 4644
rect 10498 4542 10532 4576
rect 9551 4509 9585 4537
rect 9551 4441 9585 4475
rect 8777 4393 8811 4409
rect 8901 4382 8948 4416
rect 8982 4382 9029 4416
rect 9063 4382 9110 4416
rect 9144 4382 9191 4416
rect 9225 4382 9271 4416
rect 9305 4382 9351 4416
rect 10498 4474 10532 4508
rect 7913 4298 7947 4314
rect 8669 4324 8703 4379
rect 9551 4373 9585 4407
rect 8669 4290 8811 4324
rect 8063 4242 8104 4276
rect 8138 4242 8179 4276
rect 8213 4242 8254 4276
rect 8288 4242 8328 4276
rect 8362 4242 8402 4276
rect 8436 4242 8476 4276
rect 8510 4242 8550 4276
rect 8777 4245 8811 4290
rect 8901 4272 8948 4306
rect 8982 4272 9029 4306
rect 9063 4272 9110 4306
rect 9144 4272 9191 4306
rect 9225 4272 9271 4306
rect 9305 4272 9351 4306
rect 9551 4305 9585 4339
rect 7913 4230 7947 4242
rect 7913 4162 7947 4169
rect 8669 4212 8703 4228
rect 8669 4144 8703 4178
rect 6705 4010 6739 4048
rect 7403 4066 7437 4096
rect 7403 3998 7437 4032
rect 6561 3889 6595 3909
rect 6561 3815 6595 3840
rect 7403 3930 7437 3964
rect 7403 3862 7437 3890
rect 7590 4079 7760 4096
rect 7624 4078 7760 4079
rect 7624 4045 7658 4078
rect 7590 4044 7658 4045
rect 7692 4076 7760 4078
rect 7692 4044 7726 4076
rect 7590 4042 7726 4044
rect 7590 4010 7760 4042
rect 7624 4009 7760 4010
rect 7624 3976 7658 4009
rect 7590 3975 7658 3976
rect 7692 4008 7760 4009
rect 7692 3975 7726 4008
rect 7590 3974 7726 3975
rect 7590 3941 7760 3974
rect 7624 3940 7760 3941
rect 7624 3907 7658 3940
rect 7590 3872 7658 3907
rect 7913 4094 7947 4096
rect 8631 4093 8669 4127
rect 7913 4026 7947 4060
rect 7913 3958 7947 3992
rect 8669 4076 8703 4093
rect 8669 4008 8703 4042
rect 8777 4177 8811 4211
rect 8777 4109 8811 4143
rect 9551 4237 9585 4271
rect 9551 4169 9585 4203
rect 9551 4130 9585 4135
rect 8952 4096 8991 4130
rect 9025 4096 9063 4130
rect 9097 4096 9135 4130
rect 9169 4096 9207 4130
rect 9241 4096 9279 4130
rect 9313 4096 9351 4130
rect 9397 4101 9585 4130
rect 9397 4096 9551 4101
rect 8777 4041 8811 4075
rect 8777 3991 8811 4007
rect 9734 4317 9738 4377
rect 9908 4317 9912 4377
rect 9734 4223 9738 4283
rect 9908 4223 9912 4283
rect 9734 4130 9738 4189
rect 9908 4130 9912 4189
rect 10498 4406 10532 4440
rect 10498 4338 10532 4372
rect 10614 4633 10648 4671
rect 10614 4560 10648 4599
rect 10926 4633 10960 4671
rect 10926 4560 10960 4599
rect 10614 4487 10648 4526
rect 10614 4414 10648 4453
rect 10614 4341 10648 4380
rect 10770 4475 10804 4513
rect 10770 4402 10804 4441
rect 10770 4329 10804 4368
rect 10498 4270 10532 4304
rect 10498 4202 10532 4236
rect 10498 4134 10532 4168
rect 11238 4633 11272 4671
rect 11238 4560 11272 4599
rect 10926 4487 10960 4526
rect 10926 4414 10960 4453
rect 10926 4341 10960 4380
rect 11082 4475 11116 4513
rect 11082 4402 11116 4441
rect 11082 4329 11116 4368
rect 10770 4256 10804 4295
rect 10770 4183 10804 4222
rect 11550 4633 11584 4671
rect 11550 4560 11584 4599
rect 11238 4487 11272 4526
rect 11238 4414 11272 4453
rect 11238 4341 11272 4380
rect 11394 4475 11428 4513
rect 11394 4402 11428 4441
rect 11394 4329 11428 4368
rect 11082 4256 11116 4295
rect 11082 4183 11116 4222
rect 11862 4633 11896 4671
rect 11862 4560 11896 4599
rect 11550 4487 11584 4526
rect 11550 4414 11584 4453
rect 11550 4341 11584 4380
rect 11706 4475 11740 4513
rect 11706 4402 11740 4441
rect 11706 4329 11740 4368
rect 11394 4256 11428 4295
rect 11394 4183 11428 4222
rect 12174 4633 12208 4671
rect 12174 4560 12208 4599
rect 11862 4487 11896 4526
rect 11862 4414 11896 4453
rect 11862 4341 11896 4380
rect 12018 4475 12052 4513
rect 12018 4402 12052 4441
rect 12018 4329 12052 4368
rect 11706 4256 11740 4295
rect 11706 4183 11740 4222
rect 12486 4633 12520 4671
rect 12486 4560 12520 4599
rect 12174 4487 12208 4526
rect 12174 4414 12208 4453
rect 12174 4341 12208 4380
rect 12330 4475 12364 4513
rect 12330 4402 12364 4441
rect 12330 4329 12364 4368
rect 12018 4256 12052 4295
rect 12018 4183 12052 4222
rect 12798 4633 12832 4671
rect 12798 4560 12832 4599
rect 12486 4487 12520 4526
rect 12486 4414 12520 4453
rect 12486 4341 12520 4380
rect 12642 4475 12676 4513
rect 12642 4402 12676 4441
rect 12642 4329 12676 4368
rect 12330 4256 12364 4295
rect 12330 4183 12364 4222
rect 13110 4631 13144 4671
rect 13110 4557 13144 4597
rect 12798 4487 12832 4526
rect 12798 4414 12832 4453
rect 12798 4341 12832 4380
rect 12954 4475 12988 4513
rect 12954 4402 12988 4441
rect 12954 4329 12988 4368
rect 12642 4256 12676 4295
rect 12642 4183 12676 4222
rect 12954 4256 12988 4295
rect 12954 4183 12988 4222
rect 13110 4483 13144 4523
rect 13110 4408 13144 4449
rect 13110 4333 13144 4374
rect 13110 4258 13144 4299
rect 13110 4183 13144 4224
rect 13496 4645 13530 4657
rect 13496 4577 13530 4584
rect 13496 4509 13530 4511
rect 13496 4472 13530 4475
rect 13496 4399 13530 4407
rect 13496 4326 13530 4339
rect 13496 4253 13530 4271
rect 13496 4180 13530 4203
rect 9551 4033 9585 4067
rect 8669 3958 8703 3974
rect 9551 3965 9585 3999
rect 7947 3890 8029 3924
rect 8063 3890 8104 3924
rect 8138 3890 8179 3924
rect 8213 3890 8254 3924
rect 8288 3890 8328 3924
rect 8362 3890 8402 3924
rect 8436 3890 8476 3924
rect 8510 3890 8550 3924
rect 8584 3890 8614 3924
rect 8703 3890 8741 3924
rect 8901 3920 8948 3954
rect 8982 3920 9029 3954
rect 9063 3920 9110 3954
rect 9144 3920 9191 3954
rect 9225 3920 9271 3954
rect 9305 3920 9351 3954
rect 10498 3995 10532 4100
rect 13496 4107 13530 4135
rect 10697 4037 10735 4071
rect 10769 4037 10807 4071
rect 10841 4037 10879 4071
rect 10913 4037 10951 4071
rect 10985 4037 11023 4071
rect 11057 4037 11095 4071
rect 11129 4037 11167 4071
rect 11201 4037 11239 4071
rect 11273 4037 11311 4071
rect 11345 4037 11383 4071
rect 11417 4037 11455 4071
rect 11489 4037 11527 4071
rect 11561 4037 11599 4071
rect 11633 4037 11672 4071
rect 11706 4037 11745 4071
rect 11779 4037 11818 4071
rect 11852 4037 11891 4071
rect 11925 4037 11964 4071
rect 11998 4037 12037 4071
rect 12071 4037 12110 4071
rect 12144 4037 12183 4071
rect 12217 4037 12256 4071
rect 12290 4037 12329 4071
rect 12363 4037 12402 4071
rect 12436 4037 12475 4071
rect 12509 4037 12548 4071
rect 12582 4037 12621 4071
rect 12655 4037 12694 4071
rect 12728 4037 12767 4071
rect 12801 4037 12840 4071
rect 12874 4037 12913 4071
rect 12947 4037 12986 4071
rect 13020 4037 13059 4071
rect 13496 4033 13530 4067
rect 10566 3995 10600 3999
rect 10634 3995 10668 3999
rect 10702 3995 10736 3999
rect 10770 3995 10804 3999
rect 10498 3965 10510 3995
rect 10566 3965 10583 3995
rect 10634 3965 10656 3995
rect 10702 3965 10729 3995
rect 10770 3965 10802 3995
rect 10838 3965 10872 3999
rect 10906 3995 10940 3999
rect 10974 3995 11008 3999
rect 11042 3995 11076 3999
rect 11110 3995 11144 3999
rect 11178 3995 11212 3999
rect 11246 3995 11280 3999
rect 11314 3995 11348 3999
rect 10909 3965 10940 3995
rect 10982 3965 11008 3995
rect 11055 3965 11076 3995
rect 11128 3965 11144 3995
rect 11201 3965 11212 3995
rect 11274 3965 11280 3995
rect 11347 3965 11348 3995
rect 11382 3995 11416 3999
rect 11450 3995 11484 3999
rect 11518 3995 11552 3999
rect 11586 3995 11620 3999
rect 11654 3995 11688 3999
rect 11382 3965 11386 3995
rect 11450 3965 11460 3995
rect 11518 3965 11534 3995
rect 11586 3965 11608 3995
rect 11654 3965 11682 3995
rect 11722 3965 11756 3999
rect 11790 3965 11824 3999
rect 11858 3995 11892 3999
rect 11926 3995 11960 3999
rect 11994 3995 12028 3999
rect 12062 3995 12096 3999
rect 12130 3995 12164 3999
rect 11864 3965 11892 3995
rect 11938 3965 11960 3995
rect 12012 3965 12028 3995
rect 12086 3965 12096 3995
rect 12160 3965 12164 3995
rect 12198 3995 12232 3999
rect 12266 3995 12300 3999
rect 12334 3995 12368 3999
rect 12402 3995 12436 3999
rect 12470 3995 12504 3999
rect 12538 3995 12572 3999
rect 12198 3965 12200 3995
rect 12266 3965 12274 3995
rect 12334 3965 12348 3995
rect 12402 3965 12422 3995
rect 12470 3965 12496 3995
rect 12538 3965 12570 3995
rect 12606 3965 12640 3999
rect 12674 3995 12708 3999
rect 12742 3995 12776 3999
rect 12810 3995 12844 3999
rect 12878 3995 12912 3999
rect 12946 3995 12980 3999
rect 12678 3965 12708 3995
rect 12752 3965 12776 3995
rect 12826 3965 12844 3995
rect 12900 3965 12912 3995
rect 12974 3965 12980 3995
rect 13014 3995 13048 3999
rect 10544 3961 10583 3965
rect 10617 3961 10656 3965
rect 10690 3961 10729 3965
rect 10763 3961 10802 3965
rect 10836 3961 10875 3965
rect 10909 3961 10948 3965
rect 10982 3961 11021 3965
rect 11055 3961 11094 3965
rect 11128 3961 11167 3965
rect 11201 3961 11240 3965
rect 11274 3961 11313 3965
rect 11347 3961 11386 3965
rect 11420 3961 11460 3965
rect 11494 3961 11534 3965
rect 11568 3961 11608 3965
rect 11642 3961 11682 3965
rect 11716 3961 11756 3965
rect 11790 3961 11830 3965
rect 11864 3961 11904 3965
rect 11938 3961 11978 3965
rect 12012 3961 12052 3965
rect 12086 3961 12126 3965
rect 12160 3961 12200 3965
rect 12234 3961 12274 3965
rect 12308 3961 12348 3965
rect 12382 3961 12422 3965
rect 12456 3961 12496 3965
rect 12530 3961 12570 3965
rect 12604 3961 12644 3965
rect 12678 3961 12718 3965
rect 12752 3961 12792 3965
rect 12826 3961 12866 3965
rect 12900 3961 12940 3965
rect 12974 3961 13014 3965
rect 13082 3995 13116 3999
rect 13150 3995 13184 3999
rect 13218 3995 13252 3999
rect 13286 3995 13320 3999
rect 13354 3995 13388 3999
rect 13422 3995 13530 3999
rect 13082 3965 13088 3995
rect 13150 3965 13162 3995
rect 13218 3965 13236 3995
rect 13286 3965 13310 3995
rect 13354 3965 13384 3995
rect 13422 3965 13458 3995
rect 13048 3961 13088 3965
rect 13122 3961 13162 3965
rect 13196 3961 13236 3965
rect 13270 3961 13310 3965
rect 13344 3961 13384 3965
rect 13418 3961 13458 3965
rect 13492 3961 13530 3995
rect 9551 3897 9585 3931
rect 6814 3786 6852 3820
rect 6886 3786 6924 3820
rect 6958 3786 6996 3820
rect 7030 3786 7068 3820
rect 7102 3786 7140 3820
rect 7174 3786 7212 3820
rect 7403 3815 7437 3828
rect 6561 3736 6595 3771
rect 6561 3667 6595 3702
rect 6561 3598 6595 3633
rect 6561 3488 6595 3564
rect 7589 3781 7590 3816
rect 7403 3726 7437 3760
rect 7403 3658 7437 3692
rect 7403 3590 7437 3624
rect 7403 3522 7437 3556
rect 4793 3454 4949 3460
rect 4983 3454 4987 3488
rect 5051 3454 5061 3488
rect 5119 3454 5134 3488
rect 5187 3454 5207 3488
rect 5255 3454 5280 3488
rect 5323 3454 5353 3488
rect 5391 3454 5425 3488
rect 5460 3454 5493 3488
rect 5533 3454 5561 3488
rect 5606 3454 5629 3488
rect 5679 3454 5697 3488
rect 5752 3454 5765 3488
rect 5825 3454 5833 3488
rect 5898 3454 5901 3488
rect 5935 3454 5937 3488
rect 6003 3454 6010 3488
rect 6071 3454 6083 3488
rect 6139 3454 6156 3488
rect 6207 3454 6229 3488
rect 6275 3454 6302 3488
rect 6343 3454 6375 3488
rect 6411 3454 6445 3488
rect 6482 3454 6513 3488
rect 6555 3454 6581 3488
rect 6628 3454 6649 3488
rect 6701 3454 6717 3488
rect 6774 3454 6785 3488
rect 6847 3454 6853 3488
rect 6920 3454 6921 3488
rect 6955 3454 6959 3488
rect 7023 3454 7032 3488
rect 7091 3454 7105 3488
rect 7159 3454 7178 3488
rect 7227 3454 7251 3488
rect 7295 3454 7324 3488
rect 7363 3454 7397 3488
rect 7431 3454 7437 3488
rect 7760 3781 7767 3816
rect 7913 3842 7947 3856
rect 0 3242 68 3295
rect 102 3242 170 3261
rect 0 3204 170 3242
rect 7590 3204 7760 3498
rect 0 3170 7760 3204
rect 7664 64 7760 3170
rect 7913 3760 7947 3788
rect 8669 3863 8703 3890
rect 8669 3795 8703 3829
rect 9551 3829 9585 3863
rect 7913 3686 7947 3720
rect 8063 3714 8104 3748
rect 8138 3714 8179 3748
rect 8213 3714 8254 3748
rect 8288 3714 8328 3748
rect 8362 3714 8402 3748
rect 8436 3714 8476 3748
rect 8510 3714 8550 3748
rect 8669 3745 8703 3761
rect 8777 3799 8821 3815
rect 8811 3765 8821 3799
rect 8777 3731 8821 3765
rect 8901 3744 8948 3778
rect 8982 3744 9029 3778
rect 9063 3744 9110 3778
rect 9144 3744 9191 3778
rect 9225 3744 9271 3778
rect 9305 3744 9351 3778
rect 9551 3761 9585 3795
rect 7913 3618 7947 3645
rect 8811 3697 8821 3731
rect 8777 3663 8821 3697
rect 8063 3604 8101 3638
rect 8135 3604 8173 3638
rect 8811 3629 8821 3663
rect 7913 3550 7947 3564
rect 7913 3482 7947 3483
rect 7913 3414 7947 3448
rect 7913 3346 7947 3380
rect 7913 3278 7947 3312
rect 7913 3210 7947 3244
rect 7913 3142 7947 3176
rect 8269 3577 8303 3593
rect 8269 3509 8303 3543
rect 8777 3514 8821 3629
rect 9551 3693 9585 3727
rect 9551 3625 9585 3659
rect 8901 3568 8942 3602
rect 8976 3568 9017 3602
rect 9051 3568 9092 3602
rect 9126 3568 9166 3602
rect 9200 3568 9240 3602
rect 9274 3568 9314 3602
rect 9348 3568 9388 3602
rect 9551 3557 9585 3591
rect 7913 3074 7947 3108
rect 8017 3117 8219 3148
rect 8017 3083 8029 3117
rect 8063 3083 8101 3117
rect 8135 3083 8173 3117
rect 8207 3083 8219 3117
rect 8269 3043 8303 3475
rect 8411 3477 8459 3511
rect 8493 3477 8541 3511
rect 8575 3477 8622 3511
rect 8656 3477 8703 3511
rect 8777 3480 8789 3514
rect 8823 3480 8861 3514
rect 9551 3489 9585 3523
rect 8377 3343 8737 3477
rect 8411 3309 8737 3343
rect 8377 3304 8737 3309
rect 9551 3421 9585 3455
rect 9551 3353 9585 3387
rect 8377 3275 8411 3304
rect 8377 3225 8411 3241
rect 9551 3285 9585 3319
rect 9551 3217 9585 3251
rect 9908 3431 11286 3443
rect 9934 3397 9975 3431
rect 10009 3397 10050 3431
rect 10084 3397 10125 3431
rect 10159 3397 10200 3431
rect 10234 3397 10275 3431
rect 10309 3397 10350 3431
rect 10384 3397 10425 3431
rect 10459 3397 10500 3431
rect 10534 3397 10574 3431
rect 10608 3397 10648 3431
rect 10682 3397 10722 3431
rect 10756 3397 10796 3431
rect 10830 3397 10870 3431
rect 10904 3397 10944 3431
rect 10978 3397 11018 3431
rect 11052 3397 11092 3431
rect 11126 3397 11166 3431
rect 11200 3397 11240 3431
rect 11274 3397 11286 3431
rect 9908 3370 11286 3397
rect 11132 3336 11166 3370
rect 11200 3336 11286 3370
rect 11132 3302 11252 3336
rect 9840 3261 9942 3295
rect 11132 3268 11184 3302
rect 9738 3200 9942 3261
rect 11064 3234 11184 3268
rect 11064 3200 11116 3234
rect 9551 3149 9585 3183
rect 8455 3117 9405 3148
rect 8455 3083 8467 3117
rect 8501 3083 8542 3117
rect 8576 3083 8617 3117
rect 8651 3083 8692 3117
rect 8726 3083 8767 3117
rect 8801 3083 8841 3117
rect 8875 3083 8915 3117
rect 8949 3083 8989 3117
rect 9023 3083 9063 3117
rect 9097 3083 9137 3117
rect 9171 3083 9211 3117
rect 9245 3083 9285 3117
rect 9319 3083 9359 3117
rect 9393 3083 9405 3117
rect 7913 3006 7947 3040
rect 8231 3009 8269 3043
rect 9551 3081 9585 3115
rect 9551 3013 9619 3047
rect 9653 3013 9687 3047
rect 9721 3013 9755 3047
rect 9789 3013 9823 3047
rect 9857 3013 9891 3047
rect 9925 3013 9959 3047
rect 9993 3013 10027 3047
rect 10061 3013 10095 3047
rect 10129 3013 10163 3047
rect 10197 3013 10231 3047
rect 10265 3013 10299 3047
rect 10333 3013 10367 3047
rect 10401 3013 10435 3047
rect 10469 3013 10503 3047
rect 10537 3013 10571 3047
rect 10605 3013 10639 3047
rect 10673 3013 10707 3047
rect 10741 3013 10775 3047
rect 10809 3013 10843 3047
rect 10877 3013 10963 3047
rect 7913 2938 7947 2972
rect 10929 2945 10963 2979
rect 7913 2871 7947 2904
rect 8106 2877 8148 2911
rect 8182 2877 8224 2911
rect 8258 2877 8300 2911
rect 8334 2877 8376 2911
rect 8410 2877 8452 2911
rect 8486 2877 8528 2911
rect 8562 2877 8604 2911
rect 8638 2877 8680 2911
rect 8714 2877 8756 2911
rect 8790 2877 8832 2911
rect 8866 2877 8908 2911
rect 8942 2877 8984 2911
rect 9018 2877 9061 2911
rect 9095 2877 9138 2911
rect 9172 2877 9215 2911
rect 10929 2877 10963 2911
rect 7913 2802 7947 2836
rect 10929 2817 10963 2843
rect 7913 2734 7947 2764
rect 7913 2666 7947 2691
rect 7913 2598 7947 2618
rect 7913 2530 7947 2545
rect 7913 2462 7947 2472
rect 7913 2394 7947 2399
rect 7913 2287 7947 2292
rect 7913 2214 7947 2224
rect 7913 2141 7947 2156
rect 7913 2068 7947 2088
rect 7913 1995 7947 2020
rect 7913 1922 7947 1952
rect 7913 1850 7947 1884
rect 7913 1782 7947 1815
rect 7913 1714 7947 1742
rect 7913 1646 7947 1669
rect 7913 1578 7947 1596
rect 7913 1510 7947 1523
rect 7913 1442 7947 1450
rect 7913 1374 7947 1377
rect 7913 1338 7947 1340
rect 7913 1265 7947 1272
rect 7913 1192 7947 1204
rect 7913 1119 7947 1136
rect 7913 1046 7947 1068
rect 7913 973 7947 1000
rect 7913 900 7947 932
rect 7913 830 7947 864
rect 8053 2745 8087 2783
rect 8053 2673 8087 2711
rect 8965 2745 8999 2783
rect 8965 2673 8999 2711
rect 8053 2601 8087 2639
rect 8053 2529 8087 2567
rect 8053 2457 8087 2495
rect 8053 2385 8087 2423
rect 8053 2313 8087 2351
rect 8053 2241 8087 2279
rect 8053 2169 8087 2207
rect 8053 2097 8087 2135
rect 8053 2025 8087 2063
rect 8053 1953 8087 1991
rect 8053 1881 8087 1919
rect 8053 1809 8087 1847
rect 8053 1737 8087 1775
rect 8053 1665 8087 1703
rect 8053 1593 8087 1631
rect 8053 1521 8087 1559
rect 8053 1449 8087 1487
rect 8053 1377 8087 1415
rect 8053 1305 8087 1343
rect 8053 1233 8087 1271
rect 8053 1161 8087 1199
rect 8053 1089 8087 1127
rect 8053 1017 8087 1055
rect 8053 944 8087 983
rect 8053 871 8087 910
rect 8509 2585 8543 2625
rect 8509 2511 8543 2551
rect 8509 2437 8543 2477
rect 8509 2363 8543 2403
rect 8509 2289 8543 2329
rect 8509 2215 8543 2255
rect 8509 2141 8543 2181
rect 8509 2067 8543 2107
rect 8509 1993 8543 2033
rect 8509 1919 8543 1959
rect 8509 1845 8543 1885
rect 8509 1771 8543 1811
rect 8509 1696 8543 1737
rect 8509 1621 8543 1662
rect 8509 1546 8543 1587
rect 8509 1471 8543 1512
rect 8509 1396 8543 1437
rect 8509 1321 8543 1362
rect 8509 1246 8543 1287
rect 8509 1171 8543 1212
rect 8509 1096 8543 1137
rect 8509 1021 8543 1062
rect 8509 946 8543 987
rect 8509 871 8543 912
rect 9877 2745 9911 2783
rect 9877 2673 9911 2711
rect 8965 2601 8999 2639
rect 8965 2529 8999 2567
rect 8965 2457 8999 2495
rect 8965 2385 8999 2423
rect 8965 2313 8999 2351
rect 8965 2241 8999 2279
rect 8965 2169 8999 2207
rect 8965 2097 8999 2135
rect 8965 2025 8999 2063
rect 8965 1953 8999 1991
rect 8965 1881 8999 1919
rect 8965 1809 8999 1847
rect 8965 1737 8999 1775
rect 8965 1665 8999 1703
rect 8965 1593 8999 1631
rect 8965 1521 8999 1559
rect 8965 1449 8999 1487
rect 8965 1377 8999 1415
rect 8965 1305 8999 1343
rect 8965 1233 8999 1271
rect 8965 1161 8999 1199
rect 8965 1089 8999 1127
rect 8965 1017 8999 1055
rect 8965 944 8999 983
rect 8965 871 8999 910
rect 9421 2585 9455 2625
rect 9421 2511 9455 2551
rect 9421 2437 9455 2477
rect 9421 2363 9455 2403
rect 9421 2289 9455 2329
rect 9421 2215 9455 2255
rect 9421 2141 9455 2181
rect 9421 2067 9455 2107
rect 9421 1993 9455 2033
rect 9421 1919 9455 1959
rect 9421 1845 9455 1885
rect 9421 1771 9455 1811
rect 9421 1696 9455 1737
rect 9421 1621 9455 1662
rect 9421 1546 9455 1587
rect 9421 1471 9455 1512
rect 9421 1396 9455 1437
rect 9421 1321 9455 1362
rect 9421 1246 9455 1287
rect 9421 1171 9455 1212
rect 9421 1096 9455 1137
rect 9421 1021 9455 1062
rect 9421 946 9455 987
rect 9421 871 9455 912
rect 10789 2745 10823 2783
rect 10789 2673 10823 2711
rect 9877 2601 9911 2639
rect 9877 2529 9911 2567
rect 9877 2457 9911 2495
rect 9877 2385 9911 2423
rect 9877 2313 9911 2351
rect 9877 2241 9911 2279
rect 9877 2169 9911 2207
rect 9877 2097 9911 2135
rect 9877 2025 9911 2063
rect 9877 1953 9911 1991
rect 9877 1881 9911 1919
rect 9877 1809 9911 1847
rect 9877 1737 9911 1775
rect 9877 1665 9911 1703
rect 9877 1593 9911 1631
rect 9877 1521 9911 1559
rect 9877 1449 9911 1487
rect 9877 1377 9911 1415
rect 9877 1305 9911 1343
rect 9877 1233 9911 1271
rect 9877 1161 9911 1199
rect 9877 1089 9911 1127
rect 9877 1017 9911 1055
rect 9877 944 9911 983
rect 9877 871 9911 910
rect 10333 2585 10367 2625
rect 10333 2511 10367 2551
rect 10333 2437 10367 2477
rect 10333 2363 10367 2403
rect 10333 2289 10367 2329
rect 10333 2215 10367 2255
rect 10333 2141 10367 2181
rect 10333 2067 10367 2107
rect 10333 1993 10367 2033
rect 10333 1919 10367 1959
rect 10333 1845 10367 1885
rect 10333 1771 10367 1811
rect 10333 1696 10367 1737
rect 10333 1621 10367 1662
rect 10333 1546 10367 1587
rect 10333 1471 10367 1512
rect 10333 1396 10367 1437
rect 10333 1321 10367 1362
rect 10333 1246 10367 1287
rect 10333 1171 10367 1212
rect 10333 1096 10367 1137
rect 10333 1021 10367 1062
rect 10333 946 10367 987
rect 10333 871 10367 912
rect 10789 2601 10823 2639
rect 10789 2529 10823 2567
rect 10789 2457 10823 2495
rect 10789 2385 10823 2423
rect 10789 2313 10823 2351
rect 10789 2241 10823 2279
rect 10789 2169 10823 2207
rect 10789 2097 10823 2135
rect 10789 2025 10823 2063
rect 10789 1953 10823 1991
rect 10789 1881 10823 1919
rect 10789 1809 10823 1847
rect 10789 1737 10823 1775
rect 10789 1665 10823 1703
rect 10789 1593 10823 1631
rect 10789 1521 10823 1559
rect 10789 1449 10823 1487
rect 10789 1377 10823 1415
rect 10789 1305 10823 1343
rect 10789 1233 10823 1271
rect 10789 1161 10823 1199
rect 10789 1089 10823 1127
rect 10789 1017 10823 1055
rect 10789 944 10823 983
rect 10789 871 10823 910
rect 10929 2744 10963 2775
rect 10929 2673 10963 2707
rect 10929 2605 10963 2637
rect 10929 2537 10963 2564
rect 10929 2469 10963 2491
rect 10929 2401 10963 2418
rect 10929 2333 10963 2345
rect 10929 2265 10963 2272
rect 10929 2197 10963 2199
rect 10929 2159 10963 2163
rect 10929 2085 10963 2095
rect 10929 2011 10963 2027
rect 10929 1937 10963 1959
rect 10929 1863 10963 1891
rect 10929 1789 10963 1823
rect 10929 1721 10963 1755
rect 10929 1653 10963 1681
rect 10929 1585 10963 1607
rect 10929 1517 10963 1533
rect 10929 1449 10963 1459
rect 10929 1381 10963 1385
rect 10929 1345 10963 1347
rect 10929 1271 10963 1279
rect 10929 1197 10963 1211
rect 10929 1123 10963 1143
rect 10929 1049 10963 1075
rect 10929 975 10963 1007
rect 10929 905 10963 939
rect 10929 837 10963 867
rect 7913 755 7947 793
rect 10929 755 10963 793
rect 7913 721 7919 755
rect 7971 721 7992 755
rect 8039 721 8065 755
rect 8107 721 8138 755
rect 8175 721 8209 755
rect 8245 721 8277 755
rect 8318 721 8345 755
rect 8391 721 8413 755
rect 8464 721 8481 755
rect 8537 721 8549 755
rect 8610 721 8617 755
rect 8683 721 8685 755
rect 8719 721 8722 755
rect 8787 721 8795 755
rect 8856 721 8868 755
rect 8925 721 8941 755
rect 8994 721 9014 755
rect 9063 721 9087 755
rect 9132 721 9160 755
rect 9201 721 9233 755
rect 9270 721 9305 755
rect 9340 721 9374 755
rect 9413 721 9443 755
rect 9486 721 9512 755
rect 9559 721 9581 755
rect 9632 721 9650 755
rect 9705 721 9719 755
rect 9778 721 9788 755
rect 9851 721 9857 755
rect 9924 721 9926 755
rect 9960 721 9963 755
rect 10029 721 10036 755
rect 10070 721 10109 755
rect 10143 721 10183 755
rect 10217 721 10257 755
rect 10291 721 10331 755
rect 10365 721 10405 755
rect 10439 721 10479 755
rect 10513 721 10553 755
rect 10587 721 10627 755
rect 10661 721 10701 755
rect 10735 721 10775 755
rect 10809 721 10849 755
rect 10883 721 10923 755
rect 10957 721 10963 755
rect 7913 687 7947 721
rect 7913 619 7947 649
rect 7913 551 7947 567
rect 7913 483 7947 485
rect 7913 436 7947 449
rect 7913 353 7947 381
rect 10929 687 10963 721
rect 10929 619 10963 653
rect 10929 551 10963 585
rect 10929 483 10963 517
rect 10929 415 10963 449
rect 10929 347 10963 381
rect 7913 313 7937 319
rect 7971 313 7985 347
rect 8040 313 8058 347
rect 8109 313 8131 347
rect 8178 313 8204 347
rect 8247 313 8277 347
rect 8316 313 8350 347
rect 8385 313 8420 347
rect 8457 313 8489 347
rect 8530 313 8558 347
rect 8603 313 8627 347
rect 8676 313 8696 347
rect 8749 313 8765 347
rect 8822 313 8834 347
rect 8895 313 8903 347
rect 8968 313 8972 347
rect 9006 313 9007 347
rect 9075 313 9081 347
rect 9144 313 9155 347
rect 9213 313 9229 347
rect 9282 313 9303 347
rect 9351 313 9377 347
rect 9420 313 9451 347
rect 9489 313 9524 347
rect 9559 313 9593 347
rect 9633 313 9662 347
rect 9707 313 9731 347
rect 9781 313 9800 347
rect 9855 313 9869 347
rect 9929 313 9938 347
rect 10003 313 10007 347
rect 10041 313 10043 347
rect 10110 313 10117 347
rect 10179 313 10191 347
rect 10248 313 10265 347
rect 10317 313 10339 347
rect 10386 313 10413 347
rect 10455 313 10487 347
rect 10524 313 10559 347
rect 10595 313 10628 347
rect 10669 313 10697 347
rect 10743 313 10766 347
rect 10817 313 10835 347
rect 10891 313 10905 347
rect 10939 313 10963 347
rect 12540 3339 12552 3373
rect 12608 3339 12629 3373
rect 12663 3339 12706 3373
rect 12774 3339 12783 3373
rect 12842 3339 12860 3373
rect 12910 3339 12938 3373
rect 12978 3339 13012 3373
rect 13050 3339 13080 3373
rect 13128 3339 13148 3373
rect 13206 3339 13216 3373
rect 13318 3339 13328 3373
rect 13362 3339 13400 3373
rect 12540 3247 12574 3339
rect 13366 3271 13400 3305
rect 12540 3179 12574 3213
rect 12540 3111 12574 3145
rect 12624 3234 12658 3250
rect 12624 3166 12658 3200
rect 13366 3203 13400 3229
rect 12814 3157 12852 3191
rect 12886 3157 12924 3191
rect 12958 3157 12996 3191
rect 13030 3157 13068 3191
rect 13102 3157 13140 3191
rect 12624 3111 12658 3132
rect 13366 3135 13400 3157
rect 12658 3077 12696 3111
rect 12540 3043 12574 3077
rect 13366 3047 13400 3085
rect 12540 2975 12552 3009
rect 12586 2975 12630 3009
rect 12686 2975 12707 3009
rect 12754 2975 12784 3009
rect 12822 2975 12856 3009
rect 12895 2975 12924 3009
rect 12972 2975 12992 3009
rect 13049 2975 13060 3009
rect 13126 2975 13128 3009
rect 13162 2975 13169 3009
rect 13230 2975 13246 3009
rect 13298 2975 13332 3009
rect 13366 2975 13400 3013
rect 13693 3032 13709 6602
rect 14083 3032 14099 6602
rect 13693 2997 14099 3032
rect 13693 2963 13709 2997
rect 13743 2963 13777 2997
rect 13811 2963 13845 2997
rect 13879 2963 13913 2997
rect 13947 2963 13981 2997
rect 14015 2963 14049 2997
rect 14083 2963 14099 2997
rect 13693 2928 14099 2963
rect 13693 2894 13709 2928
rect 13743 2894 13777 2928
rect 13811 2894 13845 2928
rect 13879 2894 13913 2928
rect 13947 2894 13981 2928
rect 14015 2894 14049 2928
rect 14083 2894 14099 2928
rect 13693 2859 14099 2894
rect 13693 2825 13709 2859
rect 13743 2825 13777 2859
rect 13811 2825 13845 2859
rect 13879 2825 13913 2859
rect 13947 2825 13981 2859
rect 14015 2825 14049 2859
rect 14083 2825 14099 2859
rect 13693 2790 14099 2825
rect 13693 2756 13709 2790
rect 13743 2756 13777 2790
rect 13811 2756 13845 2790
rect 13879 2756 13913 2790
rect 13947 2756 13981 2790
rect 14015 2756 14049 2790
rect 14083 2756 14099 2790
rect 13693 2732 14099 2756
rect 11439 2714 14099 2732
rect 11439 2680 11448 2714
rect 11482 2695 11522 2714
rect 11556 2695 11596 2714
rect 11630 2695 11670 2714
rect 11704 2695 11744 2714
rect 11778 2695 11818 2714
rect 11852 2695 11892 2714
rect 11926 2695 11966 2714
rect 12000 2695 12040 2714
rect 12074 2695 12114 2714
rect 12148 2695 12188 2714
rect 12222 2695 12262 2714
rect 12296 2695 12336 2714
rect 12370 2695 12410 2714
rect 12444 2695 12484 2714
rect 12518 2695 12558 2714
rect 11510 2680 11522 2695
rect 11580 2680 11596 2695
rect 11650 2680 11670 2695
rect 11720 2680 11744 2695
rect 11790 2680 11818 2695
rect 11860 2680 11892 2695
rect 11439 2661 11476 2680
rect 11510 2661 11546 2680
rect 11580 2661 11616 2680
rect 11650 2661 11686 2680
rect 11720 2661 11756 2680
rect 11790 2661 11826 2680
rect 11860 2661 11896 2680
rect 11930 2661 11966 2695
rect 12000 2661 12036 2695
rect 12074 2680 12106 2695
rect 12148 2680 12176 2695
rect 12222 2680 12246 2695
rect 12296 2680 12316 2695
rect 12370 2680 12385 2695
rect 12444 2680 12454 2695
rect 12518 2680 12523 2695
rect 12070 2661 12106 2680
rect 12140 2661 12176 2680
rect 12210 2661 12246 2680
rect 12280 2661 12316 2680
rect 12350 2661 12385 2680
rect 12419 2661 12454 2680
rect 12488 2661 12523 2680
rect 12557 2680 12558 2695
rect 12592 2695 12632 2714
rect 12666 2695 12706 2714
rect 12740 2695 12780 2714
rect 12814 2695 12854 2714
rect 12888 2695 12928 2714
rect 12962 2695 13002 2714
rect 13036 2695 13076 2714
rect 13110 2695 13150 2714
rect 13184 2695 13224 2714
rect 13258 2695 13298 2714
rect 13332 2695 13372 2714
rect 13406 2695 13446 2714
rect 13480 2695 13520 2714
rect 13554 2695 13594 2714
rect 13628 2695 13668 2714
rect 13702 2695 13741 2714
rect 13775 2695 13814 2714
rect 13848 2695 13887 2714
rect 13921 2695 13960 2714
rect 13994 2695 14033 2714
rect 14067 2695 14099 2714
rect 12557 2661 12592 2680
rect 12626 2680 12632 2695
rect 12695 2680 12706 2695
rect 12764 2680 12780 2695
rect 12833 2680 12854 2695
rect 12902 2680 12928 2695
rect 12971 2680 13002 2695
rect 12626 2661 12661 2680
rect 12695 2661 12730 2680
rect 12764 2661 12799 2680
rect 12833 2661 12868 2680
rect 12902 2661 12937 2680
rect 12971 2661 13006 2680
rect 13040 2661 13075 2695
rect 13110 2680 13144 2695
rect 13184 2680 13213 2695
rect 13258 2680 13282 2695
rect 13332 2680 13351 2695
rect 13406 2680 13420 2695
rect 13480 2680 13489 2695
rect 13554 2680 13558 2695
rect 13109 2661 13144 2680
rect 13178 2661 13213 2680
rect 13247 2661 13282 2680
rect 13316 2661 13351 2680
rect 13385 2661 13420 2680
rect 13454 2661 13489 2680
rect 13523 2661 13558 2680
rect 13592 2680 13594 2695
rect 13661 2680 13668 2695
rect 13730 2680 13741 2695
rect 13799 2680 13814 2695
rect 13868 2680 13887 2695
rect 13937 2680 13960 2695
rect 14006 2680 14033 2695
rect 13592 2661 13627 2680
rect 13661 2661 13696 2680
rect 13730 2661 13765 2680
rect 13799 2661 13834 2680
rect 13868 2661 13903 2680
rect 13937 2661 13972 2680
rect 14006 2661 14041 2680
rect 14075 2661 14099 2695
rect 11439 2642 14099 2661
rect 11439 2608 11448 2642
rect 11482 2627 11522 2642
rect 11556 2627 11596 2642
rect 11630 2627 11670 2642
rect 11704 2627 11744 2642
rect 11778 2627 11818 2642
rect 11852 2627 11892 2642
rect 11926 2627 11966 2642
rect 12000 2627 12040 2642
rect 12074 2627 12114 2642
rect 12148 2627 12188 2642
rect 12222 2627 12262 2642
rect 12296 2627 12336 2642
rect 12370 2627 12410 2642
rect 12444 2627 12484 2642
rect 12518 2627 12558 2642
rect 11510 2608 11522 2627
rect 11580 2608 11596 2627
rect 11650 2608 11670 2627
rect 11720 2608 11744 2627
rect 11790 2608 11818 2627
rect 11860 2608 11892 2627
rect 11439 2593 11476 2608
rect 11510 2593 11546 2608
rect 11580 2593 11616 2608
rect 11650 2593 11686 2608
rect 11720 2593 11756 2608
rect 11790 2593 11826 2608
rect 11860 2593 11896 2608
rect 11930 2593 11966 2627
rect 12000 2593 12036 2627
rect 12074 2608 12106 2627
rect 12148 2608 12176 2627
rect 12222 2608 12246 2627
rect 12296 2608 12316 2627
rect 12370 2608 12385 2627
rect 12444 2608 12454 2627
rect 12518 2608 12523 2627
rect 12070 2593 12106 2608
rect 12140 2593 12176 2608
rect 12210 2593 12246 2608
rect 12280 2593 12316 2608
rect 12350 2593 12385 2608
rect 12419 2593 12454 2608
rect 12488 2593 12523 2608
rect 12557 2608 12558 2627
rect 12592 2627 12632 2642
rect 12666 2627 12706 2642
rect 12740 2627 12780 2642
rect 12814 2627 12854 2642
rect 12888 2627 12928 2642
rect 12962 2627 13002 2642
rect 13036 2627 13076 2642
rect 13110 2627 13150 2642
rect 13184 2627 13224 2642
rect 13258 2627 13298 2642
rect 13332 2627 13372 2642
rect 13406 2627 13446 2642
rect 13480 2627 13520 2642
rect 13554 2627 13594 2642
rect 13628 2627 13668 2642
rect 13702 2627 13741 2642
rect 13775 2627 13814 2642
rect 13848 2627 13887 2642
rect 13921 2627 13960 2642
rect 13994 2627 14033 2642
rect 14067 2627 14099 2642
rect 12557 2593 12592 2608
rect 12626 2608 12632 2627
rect 12695 2608 12706 2627
rect 12764 2608 12780 2627
rect 12833 2608 12854 2627
rect 12902 2608 12928 2627
rect 12971 2608 13002 2627
rect 12626 2593 12661 2608
rect 12695 2593 12730 2608
rect 12764 2593 12799 2608
rect 12833 2593 12868 2608
rect 12902 2593 12937 2608
rect 12971 2593 13006 2608
rect 13040 2593 13075 2627
rect 13110 2608 13144 2627
rect 13184 2608 13213 2627
rect 13258 2608 13282 2627
rect 13332 2608 13351 2627
rect 13406 2608 13420 2627
rect 13480 2608 13489 2627
rect 13554 2608 13558 2627
rect 13109 2593 13144 2608
rect 13178 2593 13213 2608
rect 13247 2593 13282 2608
rect 13316 2593 13351 2608
rect 13385 2593 13420 2608
rect 13454 2593 13489 2608
rect 13523 2593 13558 2608
rect 13592 2608 13594 2627
rect 13661 2608 13668 2627
rect 13730 2608 13741 2627
rect 13799 2608 13814 2627
rect 13868 2608 13887 2627
rect 13937 2608 13960 2627
rect 14006 2608 14033 2627
rect 13592 2593 13627 2608
rect 13661 2593 13696 2608
rect 13730 2593 13765 2608
rect 13799 2593 13834 2608
rect 13868 2593 13903 2608
rect 13937 2593 13972 2608
rect 14006 2593 14041 2608
rect 14075 2593 14099 2627
rect 11439 2570 14099 2593
rect 11439 2536 11448 2570
rect 11482 2559 11522 2570
rect 11556 2559 11596 2570
rect 11630 2559 11670 2570
rect 11704 2559 11744 2570
rect 11778 2559 11818 2570
rect 11852 2559 11892 2570
rect 11926 2559 11966 2570
rect 12000 2559 12040 2570
rect 12074 2559 12114 2570
rect 12148 2559 12188 2570
rect 12222 2559 12262 2570
rect 12296 2559 12336 2570
rect 12370 2559 12410 2570
rect 12444 2559 12484 2570
rect 12518 2559 12558 2570
rect 11510 2536 11522 2559
rect 11580 2536 11596 2559
rect 11650 2536 11670 2559
rect 11720 2536 11744 2559
rect 11790 2536 11818 2559
rect 11860 2536 11892 2559
rect 11439 2525 11476 2536
rect 11510 2525 11546 2536
rect 11580 2525 11616 2536
rect 11650 2525 11686 2536
rect 11720 2525 11756 2536
rect 11790 2525 11826 2536
rect 11860 2525 11896 2536
rect 11930 2525 11966 2559
rect 12000 2525 12036 2559
rect 12074 2536 12106 2559
rect 12148 2536 12176 2559
rect 12222 2536 12246 2559
rect 12296 2536 12316 2559
rect 12370 2536 12385 2559
rect 12444 2536 12454 2559
rect 12518 2536 12523 2559
rect 12070 2525 12106 2536
rect 12140 2525 12176 2536
rect 12210 2525 12246 2536
rect 12280 2525 12316 2536
rect 12350 2525 12385 2536
rect 12419 2525 12454 2536
rect 12488 2525 12523 2536
rect 12557 2536 12558 2559
rect 12592 2559 12632 2570
rect 12666 2559 12706 2570
rect 12740 2559 12780 2570
rect 12814 2559 12854 2570
rect 12888 2559 12928 2570
rect 12962 2559 13002 2570
rect 13036 2559 13076 2570
rect 13110 2559 13150 2570
rect 13184 2559 13224 2570
rect 13258 2559 13298 2570
rect 13332 2559 13372 2570
rect 13406 2559 13446 2570
rect 13480 2559 13520 2570
rect 13554 2559 13594 2570
rect 13628 2559 13668 2570
rect 13702 2559 13741 2570
rect 13775 2559 13814 2570
rect 13848 2559 13887 2570
rect 13921 2559 13960 2570
rect 13994 2559 14033 2570
rect 14067 2559 14099 2570
rect 12557 2525 12592 2536
rect 12626 2536 12632 2559
rect 12695 2536 12706 2559
rect 12764 2536 12780 2559
rect 12833 2536 12854 2559
rect 12902 2536 12928 2559
rect 12971 2536 13002 2559
rect 12626 2525 12661 2536
rect 12695 2525 12730 2536
rect 12764 2525 12799 2536
rect 12833 2525 12868 2536
rect 12902 2525 12937 2536
rect 12971 2525 13006 2536
rect 13040 2525 13075 2559
rect 13110 2536 13144 2559
rect 13184 2536 13213 2559
rect 13258 2536 13282 2559
rect 13332 2536 13351 2559
rect 13406 2536 13420 2559
rect 13480 2536 13489 2559
rect 13554 2536 13558 2559
rect 13109 2525 13144 2536
rect 13178 2525 13213 2536
rect 13247 2525 13282 2536
rect 13316 2525 13351 2536
rect 13385 2525 13420 2536
rect 13454 2525 13489 2536
rect 13523 2525 13558 2536
rect 13592 2536 13594 2559
rect 13661 2536 13668 2559
rect 13730 2536 13741 2559
rect 13799 2536 13814 2559
rect 13868 2536 13887 2559
rect 13937 2536 13960 2559
rect 14006 2536 14033 2559
rect 13592 2525 13627 2536
rect 13661 2525 13696 2536
rect 13730 2525 13765 2536
rect 13799 2525 13834 2536
rect 13868 2525 13903 2536
rect 13937 2525 13972 2536
rect 14006 2525 14041 2536
rect 14075 2525 14099 2559
rect 11439 2498 14099 2525
rect 11439 2464 11448 2498
rect 11482 2491 11522 2498
rect 11556 2491 11596 2498
rect 11630 2491 11670 2498
rect 11704 2491 11744 2498
rect 11778 2491 11818 2498
rect 11852 2491 11892 2498
rect 11926 2491 11966 2498
rect 12000 2491 12040 2498
rect 12074 2491 12114 2498
rect 12148 2491 12188 2498
rect 12222 2491 12262 2498
rect 12296 2491 12336 2498
rect 12370 2491 12410 2498
rect 12444 2491 12484 2498
rect 12518 2491 12558 2498
rect 11510 2464 11522 2491
rect 11580 2464 11596 2491
rect 11650 2464 11670 2491
rect 11720 2464 11744 2491
rect 11790 2464 11818 2491
rect 11860 2464 11892 2491
rect 11439 2457 11476 2464
rect 11510 2457 11546 2464
rect 11580 2457 11616 2464
rect 11650 2457 11686 2464
rect 11720 2457 11756 2464
rect 11790 2457 11826 2464
rect 11860 2457 11896 2464
rect 11930 2457 11966 2491
rect 12000 2457 12036 2491
rect 12074 2464 12106 2491
rect 12148 2464 12176 2491
rect 12222 2464 12246 2491
rect 12296 2464 12316 2491
rect 12370 2464 12385 2491
rect 12444 2464 12454 2491
rect 12518 2464 12523 2491
rect 12070 2457 12106 2464
rect 12140 2457 12176 2464
rect 12210 2457 12246 2464
rect 12280 2457 12316 2464
rect 12350 2457 12385 2464
rect 12419 2457 12454 2464
rect 12488 2457 12523 2464
rect 12557 2464 12558 2491
rect 12592 2491 12632 2498
rect 12666 2491 12706 2498
rect 12740 2491 12780 2498
rect 12814 2491 12854 2498
rect 12888 2491 12928 2498
rect 12962 2491 13002 2498
rect 13036 2491 13076 2498
rect 13110 2491 13150 2498
rect 13184 2491 13224 2498
rect 13258 2491 13298 2498
rect 13332 2491 13372 2498
rect 13406 2491 13446 2498
rect 13480 2491 13520 2498
rect 13554 2491 13594 2498
rect 13628 2491 13668 2498
rect 13702 2491 13741 2498
rect 13775 2491 13814 2498
rect 13848 2491 13887 2498
rect 13921 2491 13960 2498
rect 13994 2491 14033 2498
rect 14067 2491 14099 2498
rect 12557 2457 12592 2464
rect 12626 2464 12632 2491
rect 12695 2464 12706 2491
rect 12764 2464 12780 2491
rect 12833 2464 12854 2491
rect 12902 2464 12928 2491
rect 12971 2464 13002 2491
rect 12626 2457 12661 2464
rect 12695 2457 12730 2464
rect 12764 2457 12799 2464
rect 12833 2457 12868 2464
rect 12902 2457 12937 2464
rect 12971 2457 13006 2464
rect 13040 2457 13075 2491
rect 13110 2464 13144 2491
rect 13184 2464 13213 2491
rect 13258 2464 13282 2491
rect 13332 2464 13351 2491
rect 13406 2464 13420 2491
rect 13480 2464 13489 2491
rect 13554 2464 13558 2491
rect 13109 2457 13144 2464
rect 13178 2457 13213 2464
rect 13247 2457 13282 2464
rect 13316 2457 13351 2464
rect 13385 2457 13420 2464
rect 13454 2457 13489 2464
rect 13523 2457 13558 2464
rect 13592 2464 13594 2491
rect 13661 2464 13668 2491
rect 13730 2464 13741 2491
rect 13799 2464 13814 2491
rect 13868 2464 13887 2491
rect 13937 2464 13960 2491
rect 14006 2464 14033 2491
rect 13592 2457 13627 2464
rect 13661 2457 13696 2464
rect 13730 2457 13765 2464
rect 13799 2457 13834 2464
rect 13868 2457 13903 2464
rect 13937 2457 13972 2464
rect 14006 2457 14041 2464
rect 14075 2457 14099 2491
rect 11439 2426 14099 2457
rect 11439 2392 11448 2426
rect 11482 2423 11522 2426
rect 11556 2423 11596 2426
rect 11630 2423 11670 2426
rect 11704 2423 11744 2426
rect 11778 2423 11818 2426
rect 11852 2423 11892 2426
rect 11926 2423 11966 2426
rect 12000 2423 12040 2426
rect 12074 2423 12114 2426
rect 12148 2423 12188 2426
rect 12222 2423 12262 2426
rect 12296 2423 12336 2426
rect 12370 2423 12410 2426
rect 12444 2423 12484 2426
rect 12518 2423 12558 2426
rect 11510 2392 11522 2423
rect 11580 2392 11596 2423
rect 11650 2392 11670 2423
rect 11720 2392 11744 2423
rect 11790 2392 11818 2423
rect 11860 2392 11892 2423
rect 11439 2389 11476 2392
rect 11510 2389 11546 2392
rect 11580 2389 11616 2392
rect 11650 2389 11686 2392
rect 11720 2389 11756 2392
rect 11790 2389 11826 2392
rect 11860 2389 11896 2392
rect 11930 2389 11966 2423
rect 12000 2389 12036 2423
rect 12074 2392 12106 2423
rect 12148 2392 12176 2423
rect 12222 2392 12246 2423
rect 12296 2392 12316 2423
rect 12370 2392 12385 2423
rect 12444 2392 12454 2423
rect 12518 2392 12523 2423
rect 12070 2389 12106 2392
rect 12140 2389 12176 2392
rect 12210 2389 12246 2392
rect 12280 2389 12316 2392
rect 12350 2389 12385 2392
rect 12419 2389 12454 2392
rect 12488 2389 12523 2392
rect 12557 2392 12558 2423
rect 12592 2423 12632 2426
rect 12666 2423 12706 2426
rect 12740 2423 12780 2426
rect 12814 2423 12854 2426
rect 12888 2423 12928 2426
rect 12962 2423 13002 2426
rect 13036 2423 13076 2426
rect 13110 2423 13150 2426
rect 13184 2423 13224 2426
rect 13258 2423 13298 2426
rect 13332 2423 13372 2426
rect 13406 2423 13446 2426
rect 13480 2423 13520 2426
rect 13554 2423 13594 2426
rect 13628 2423 13668 2426
rect 13702 2423 13741 2426
rect 13775 2423 13814 2426
rect 13848 2423 13887 2426
rect 13921 2423 13960 2426
rect 13994 2423 14033 2426
rect 14067 2423 14099 2426
rect 12557 2389 12592 2392
rect 12626 2392 12632 2423
rect 12695 2392 12706 2423
rect 12764 2392 12780 2423
rect 12833 2392 12854 2423
rect 12902 2392 12928 2423
rect 12971 2392 13002 2423
rect 12626 2389 12661 2392
rect 12695 2389 12730 2392
rect 12764 2389 12799 2392
rect 12833 2389 12868 2392
rect 12902 2389 12937 2392
rect 12971 2389 13006 2392
rect 13040 2389 13075 2423
rect 13110 2392 13144 2423
rect 13184 2392 13213 2423
rect 13258 2392 13282 2423
rect 13332 2392 13351 2423
rect 13406 2392 13420 2423
rect 13480 2392 13489 2423
rect 13554 2392 13558 2423
rect 13109 2389 13144 2392
rect 13178 2389 13213 2392
rect 13247 2389 13282 2392
rect 13316 2389 13351 2392
rect 13385 2389 13420 2392
rect 13454 2389 13489 2392
rect 13523 2389 13558 2392
rect 13592 2392 13594 2423
rect 13661 2392 13668 2423
rect 13730 2392 13741 2423
rect 13799 2392 13814 2423
rect 13868 2392 13887 2423
rect 13937 2392 13960 2423
rect 14006 2392 14033 2423
rect 13592 2389 13627 2392
rect 13661 2389 13696 2392
rect 13730 2389 13765 2392
rect 13799 2389 13834 2392
rect 13868 2389 13903 2392
rect 13937 2389 13972 2392
rect 14006 2389 14041 2392
rect 14075 2389 14099 2423
rect 11439 2355 14099 2389
rect 11439 2354 11476 2355
rect 11510 2354 11546 2355
rect 11580 2354 11616 2355
rect 11650 2354 11686 2355
rect 11720 2354 11756 2355
rect 11790 2354 11826 2355
rect 11860 2354 11896 2355
rect 11439 2320 11448 2354
rect 11510 2321 11522 2354
rect 11580 2321 11596 2354
rect 11650 2321 11670 2354
rect 11720 2321 11744 2354
rect 11790 2321 11818 2354
rect 11860 2321 11892 2354
rect 11930 2321 11966 2355
rect 12000 2321 12036 2355
rect 12070 2354 12106 2355
rect 12140 2354 12176 2355
rect 12210 2354 12246 2355
rect 12280 2354 12316 2355
rect 12350 2354 12385 2355
rect 12419 2354 12454 2355
rect 12488 2354 12523 2355
rect 12074 2321 12106 2354
rect 12148 2321 12176 2354
rect 12222 2321 12246 2354
rect 12296 2321 12316 2354
rect 12370 2321 12385 2354
rect 12444 2321 12454 2354
rect 12518 2321 12523 2354
rect 12557 2354 12592 2355
rect 12557 2321 12558 2354
rect 11482 2320 11522 2321
rect 11556 2320 11596 2321
rect 11630 2320 11670 2321
rect 11704 2320 11744 2321
rect 11778 2320 11818 2321
rect 11852 2320 11892 2321
rect 11926 2320 11966 2321
rect 12000 2320 12040 2321
rect 12074 2320 12114 2321
rect 12148 2320 12188 2321
rect 12222 2320 12262 2321
rect 12296 2320 12336 2321
rect 12370 2320 12410 2321
rect 12444 2320 12484 2321
rect 12518 2320 12558 2321
rect 12626 2354 12661 2355
rect 12695 2354 12730 2355
rect 12764 2354 12799 2355
rect 12833 2354 12868 2355
rect 12902 2354 12937 2355
rect 12971 2354 13006 2355
rect 12626 2321 12632 2354
rect 12695 2321 12706 2354
rect 12764 2321 12780 2354
rect 12833 2321 12854 2354
rect 12902 2321 12928 2354
rect 12971 2321 13002 2354
rect 13040 2321 13075 2355
rect 13109 2354 13144 2355
rect 13178 2354 13213 2355
rect 13247 2354 13282 2355
rect 13316 2354 13351 2355
rect 13385 2354 13420 2355
rect 13454 2354 13489 2355
rect 13523 2354 13558 2355
rect 13110 2321 13144 2354
rect 13184 2321 13213 2354
rect 13258 2321 13282 2354
rect 13332 2321 13351 2354
rect 13406 2321 13420 2354
rect 13480 2321 13489 2354
rect 13554 2321 13558 2354
rect 13592 2354 13627 2355
rect 13661 2354 13696 2355
rect 13730 2354 13765 2355
rect 13799 2354 13834 2355
rect 13868 2354 13903 2355
rect 13937 2354 13972 2355
rect 14006 2354 14041 2355
rect 13592 2321 13594 2354
rect 13661 2321 13668 2354
rect 13730 2321 13741 2354
rect 13799 2321 13814 2354
rect 13868 2321 13887 2354
rect 13937 2321 13960 2354
rect 14006 2321 14033 2354
rect 14075 2321 14099 2355
rect 12592 2320 12632 2321
rect 12666 2320 12706 2321
rect 12740 2320 12780 2321
rect 12814 2320 12854 2321
rect 12888 2320 12928 2321
rect 12962 2320 13002 2321
rect 13036 2320 13076 2321
rect 13110 2320 13150 2321
rect 13184 2320 13224 2321
rect 13258 2320 13298 2321
rect 13332 2320 13372 2321
rect 13406 2320 13446 2321
rect 13480 2320 13520 2321
rect 13554 2320 13594 2321
rect 13628 2320 13668 2321
rect 13702 2320 13741 2321
rect 13775 2320 13814 2321
rect 13848 2320 13887 2321
rect 13921 2320 13960 2321
rect 13994 2320 14033 2321
rect 14067 2320 14099 2321
rect 11439 2287 14099 2320
rect 11439 2282 11476 2287
rect 11510 2282 11546 2287
rect 11580 2282 11616 2287
rect 11650 2282 11686 2287
rect 11720 2282 11756 2287
rect 11790 2282 11826 2287
rect 11860 2282 11896 2287
rect 11439 2248 11448 2282
rect 11510 2253 11522 2282
rect 11580 2253 11596 2282
rect 11650 2253 11670 2282
rect 11720 2253 11744 2282
rect 11790 2253 11818 2282
rect 11860 2253 11892 2282
rect 11930 2253 11966 2287
rect 12000 2253 12036 2287
rect 12070 2282 12106 2287
rect 12140 2282 12176 2287
rect 12210 2282 12246 2287
rect 12280 2282 12316 2287
rect 12350 2282 12385 2287
rect 12419 2282 12454 2287
rect 12488 2282 12523 2287
rect 12074 2253 12106 2282
rect 12148 2253 12176 2282
rect 12222 2253 12246 2282
rect 12296 2253 12316 2282
rect 12370 2253 12385 2282
rect 12444 2253 12454 2282
rect 12518 2253 12523 2282
rect 12557 2282 12592 2287
rect 12557 2253 12558 2282
rect 11482 2248 11522 2253
rect 11556 2248 11596 2253
rect 11630 2248 11670 2253
rect 11704 2248 11744 2253
rect 11778 2248 11818 2253
rect 11852 2248 11892 2253
rect 11926 2248 11966 2253
rect 12000 2248 12040 2253
rect 12074 2248 12114 2253
rect 12148 2248 12188 2253
rect 12222 2248 12262 2253
rect 12296 2248 12336 2253
rect 12370 2248 12410 2253
rect 12444 2248 12484 2253
rect 12518 2248 12558 2253
rect 12626 2282 12661 2287
rect 12695 2282 12730 2287
rect 12764 2282 12799 2287
rect 12833 2282 12868 2287
rect 12902 2282 12937 2287
rect 12971 2282 13006 2287
rect 12626 2253 12632 2282
rect 12695 2253 12706 2282
rect 12764 2253 12780 2282
rect 12833 2253 12854 2282
rect 12902 2253 12928 2282
rect 12971 2253 13002 2282
rect 13040 2253 13075 2287
rect 13109 2282 13144 2287
rect 13178 2282 13213 2287
rect 13247 2282 13282 2287
rect 13316 2282 13351 2287
rect 13385 2282 13420 2287
rect 13454 2282 13489 2287
rect 13523 2282 13558 2287
rect 13110 2253 13144 2282
rect 13184 2253 13213 2282
rect 13258 2253 13282 2282
rect 13332 2253 13351 2282
rect 13406 2253 13420 2282
rect 13480 2253 13489 2282
rect 13554 2253 13558 2282
rect 13592 2282 13627 2287
rect 13661 2282 13696 2287
rect 13730 2282 13765 2287
rect 13799 2282 13834 2287
rect 13868 2282 13903 2287
rect 13937 2282 13972 2287
rect 14006 2282 14041 2287
rect 13592 2253 13594 2282
rect 13661 2253 13668 2282
rect 13730 2253 13741 2282
rect 13799 2253 13814 2282
rect 13868 2253 13887 2282
rect 13937 2253 13960 2282
rect 14006 2253 14033 2282
rect 14075 2253 14099 2287
rect 12592 2248 12632 2253
rect 12666 2248 12706 2253
rect 12740 2248 12780 2253
rect 12814 2248 12854 2253
rect 12888 2248 12928 2253
rect 12962 2248 13002 2253
rect 13036 2248 13076 2253
rect 13110 2248 13150 2253
rect 13184 2248 13224 2253
rect 13258 2248 13298 2253
rect 13332 2248 13372 2253
rect 13406 2248 13446 2253
rect 13480 2248 13520 2253
rect 13554 2248 13594 2253
rect 13628 2248 13668 2253
rect 13702 2248 13741 2253
rect 13775 2248 13814 2253
rect 13848 2248 13887 2253
rect 13921 2248 13960 2253
rect 13994 2248 14033 2253
rect 14067 2248 14099 2253
rect 11439 2219 14099 2248
rect 11439 2210 11476 2219
rect 11510 2210 11546 2219
rect 11580 2210 11616 2219
rect 11650 2210 11686 2219
rect 11720 2210 11756 2219
rect 11790 2210 11826 2219
rect 11860 2210 11896 2219
rect 11439 2176 11448 2210
rect 11510 2185 11522 2210
rect 11580 2185 11596 2210
rect 11650 2185 11670 2210
rect 11720 2185 11744 2210
rect 11790 2185 11818 2210
rect 11860 2185 11892 2210
rect 11930 2185 11966 2219
rect 12000 2185 12036 2219
rect 12070 2210 12106 2219
rect 12140 2210 12176 2219
rect 12210 2210 12246 2219
rect 12280 2210 12316 2219
rect 12350 2210 12385 2219
rect 12419 2210 12454 2219
rect 12488 2210 12523 2219
rect 12074 2185 12106 2210
rect 12148 2185 12176 2210
rect 12222 2185 12246 2210
rect 12296 2185 12316 2210
rect 12370 2185 12385 2210
rect 12444 2185 12454 2210
rect 12518 2185 12523 2210
rect 12557 2210 12592 2219
rect 12557 2185 12558 2210
rect 11482 2176 11522 2185
rect 11556 2176 11596 2185
rect 11630 2176 11670 2185
rect 11704 2176 11744 2185
rect 11778 2176 11818 2185
rect 11852 2176 11892 2185
rect 11926 2176 11966 2185
rect 12000 2176 12040 2185
rect 12074 2176 12114 2185
rect 12148 2176 12188 2185
rect 12222 2176 12262 2185
rect 12296 2176 12336 2185
rect 12370 2176 12410 2185
rect 12444 2176 12484 2185
rect 12518 2176 12558 2185
rect 12626 2210 12661 2219
rect 12695 2210 12730 2219
rect 12764 2210 12799 2219
rect 12833 2210 12868 2219
rect 12902 2210 12937 2219
rect 12971 2210 13006 2219
rect 12626 2185 12632 2210
rect 12695 2185 12706 2210
rect 12764 2185 12780 2210
rect 12833 2185 12854 2210
rect 12902 2185 12928 2210
rect 12971 2185 13002 2210
rect 13040 2185 13075 2219
rect 13109 2210 13144 2219
rect 13178 2210 13213 2219
rect 13247 2210 13282 2219
rect 13316 2210 13351 2219
rect 13385 2210 13420 2219
rect 13454 2210 13489 2219
rect 13523 2210 13558 2219
rect 13110 2185 13144 2210
rect 13184 2185 13213 2210
rect 13258 2185 13282 2210
rect 13332 2185 13351 2210
rect 13406 2185 13420 2210
rect 13480 2185 13489 2210
rect 13554 2185 13558 2210
rect 13592 2210 13627 2219
rect 13661 2210 13696 2219
rect 13730 2210 13765 2219
rect 13799 2210 13834 2219
rect 13868 2210 13903 2219
rect 13937 2210 13972 2219
rect 14006 2210 14041 2219
rect 13592 2185 13594 2210
rect 13661 2185 13668 2210
rect 13730 2185 13741 2210
rect 13799 2185 13814 2210
rect 13868 2185 13887 2210
rect 13937 2185 13960 2210
rect 14006 2185 14033 2210
rect 14075 2185 14099 2219
rect 12592 2176 12632 2185
rect 12666 2176 12706 2185
rect 12740 2176 12780 2185
rect 12814 2176 12854 2185
rect 12888 2176 12928 2185
rect 12962 2176 13002 2185
rect 13036 2176 13076 2185
rect 13110 2176 13150 2185
rect 13184 2176 13224 2185
rect 13258 2176 13298 2185
rect 13332 2176 13372 2185
rect 13406 2176 13446 2185
rect 13480 2176 13520 2185
rect 13554 2176 13594 2185
rect 13628 2176 13668 2185
rect 13702 2176 13741 2185
rect 13775 2176 13814 2185
rect 13848 2176 13887 2185
rect 13921 2176 13960 2185
rect 13994 2176 14033 2185
rect 14067 2176 14099 2185
rect 11439 2151 14099 2176
rect 11439 2138 11476 2151
rect 11510 2138 11546 2151
rect 11580 2138 11616 2151
rect 11650 2138 11686 2151
rect 11720 2138 11756 2151
rect 11790 2138 11826 2151
rect 11860 2138 11896 2151
rect 11439 2104 11448 2138
rect 11510 2117 11522 2138
rect 11580 2117 11596 2138
rect 11650 2117 11670 2138
rect 11720 2117 11744 2138
rect 11790 2117 11818 2138
rect 11860 2117 11892 2138
rect 11930 2117 11966 2151
rect 12000 2117 12036 2151
rect 12070 2138 12106 2151
rect 12140 2138 12176 2151
rect 12210 2138 12246 2151
rect 12280 2138 12316 2151
rect 12350 2138 12385 2151
rect 12419 2138 12454 2151
rect 12488 2138 12523 2151
rect 12074 2117 12106 2138
rect 12148 2117 12176 2138
rect 12222 2117 12246 2138
rect 12296 2117 12316 2138
rect 12370 2117 12385 2138
rect 12444 2117 12454 2138
rect 12518 2117 12523 2138
rect 12557 2138 12592 2151
rect 12557 2117 12558 2138
rect 11482 2104 11522 2117
rect 11556 2104 11596 2117
rect 11630 2104 11670 2117
rect 11704 2104 11744 2117
rect 11778 2104 11818 2117
rect 11852 2104 11892 2117
rect 11926 2104 11966 2117
rect 12000 2104 12040 2117
rect 12074 2104 12114 2117
rect 12148 2104 12188 2117
rect 12222 2104 12262 2117
rect 12296 2104 12336 2117
rect 12370 2104 12410 2117
rect 12444 2104 12484 2117
rect 12518 2104 12558 2117
rect 12626 2138 12661 2151
rect 12695 2138 12730 2151
rect 12764 2138 12799 2151
rect 12833 2138 12868 2151
rect 12902 2138 12937 2151
rect 12971 2138 13006 2151
rect 12626 2117 12632 2138
rect 12695 2117 12706 2138
rect 12764 2117 12780 2138
rect 12833 2117 12854 2138
rect 12902 2117 12928 2138
rect 12971 2117 13002 2138
rect 13040 2117 13075 2151
rect 13109 2138 13144 2151
rect 13178 2138 13213 2151
rect 13247 2138 13282 2151
rect 13316 2138 13351 2151
rect 13385 2138 13420 2151
rect 13454 2138 13489 2151
rect 13523 2138 13558 2151
rect 13110 2117 13144 2138
rect 13184 2117 13213 2138
rect 13258 2117 13282 2138
rect 13332 2117 13351 2138
rect 13406 2117 13420 2138
rect 13480 2117 13489 2138
rect 13554 2117 13558 2138
rect 13592 2138 13627 2151
rect 13661 2138 13696 2151
rect 13730 2138 13765 2151
rect 13799 2138 13834 2151
rect 13868 2138 13903 2151
rect 13937 2138 13972 2151
rect 14006 2138 14041 2151
rect 13592 2117 13594 2138
rect 13661 2117 13668 2138
rect 13730 2117 13741 2138
rect 13799 2117 13814 2138
rect 13868 2117 13887 2138
rect 13937 2117 13960 2138
rect 14006 2117 14033 2138
rect 14075 2117 14099 2151
rect 12592 2104 12632 2117
rect 12666 2104 12706 2117
rect 12740 2104 12780 2117
rect 12814 2104 12854 2117
rect 12888 2104 12928 2117
rect 12962 2104 13002 2117
rect 13036 2104 13076 2117
rect 13110 2104 13150 2117
rect 13184 2104 13224 2117
rect 13258 2104 13298 2117
rect 13332 2104 13372 2117
rect 13406 2104 13446 2117
rect 13480 2104 13520 2117
rect 13554 2104 13594 2117
rect 13628 2104 13668 2117
rect 13702 2104 13741 2117
rect 13775 2104 13814 2117
rect 13848 2104 13887 2117
rect 13921 2104 13960 2117
rect 13994 2104 14033 2117
rect 14067 2104 14099 2117
rect 11439 2083 14099 2104
rect 11439 2066 11476 2083
rect 11510 2066 11546 2083
rect 11580 2066 11616 2083
rect 11650 2066 11686 2083
rect 11720 2066 11756 2083
rect 11790 2066 11826 2083
rect 11860 2066 11896 2083
rect 11439 2032 11448 2066
rect 11510 2049 11522 2066
rect 11580 2049 11596 2066
rect 11650 2049 11670 2066
rect 11720 2049 11744 2066
rect 11790 2049 11818 2066
rect 11860 2049 11892 2066
rect 11930 2049 11966 2083
rect 12000 2049 12036 2083
rect 12070 2066 12106 2083
rect 12140 2066 12176 2083
rect 12210 2066 12246 2083
rect 12280 2066 12316 2083
rect 12350 2066 12385 2083
rect 12419 2066 12454 2083
rect 12488 2066 12523 2083
rect 12074 2049 12106 2066
rect 12148 2049 12176 2066
rect 12222 2049 12246 2066
rect 12296 2049 12316 2066
rect 12370 2049 12385 2066
rect 12444 2049 12454 2066
rect 12518 2049 12523 2066
rect 12557 2066 12592 2083
rect 12557 2049 12558 2066
rect 11482 2032 11522 2049
rect 11556 2032 11596 2049
rect 11630 2032 11670 2049
rect 11704 2032 11744 2049
rect 11778 2032 11818 2049
rect 11852 2032 11892 2049
rect 11926 2032 11966 2049
rect 12000 2032 12040 2049
rect 12074 2032 12114 2049
rect 12148 2032 12188 2049
rect 12222 2032 12262 2049
rect 12296 2032 12336 2049
rect 12370 2032 12410 2049
rect 12444 2032 12484 2049
rect 12518 2032 12558 2049
rect 12626 2066 12661 2083
rect 12695 2066 12730 2083
rect 12764 2066 12799 2083
rect 12833 2066 12868 2083
rect 12902 2066 12937 2083
rect 12971 2066 13006 2083
rect 12626 2049 12632 2066
rect 12695 2049 12706 2066
rect 12764 2049 12780 2066
rect 12833 2049 12854 2066
rect 12902 2049 12928 2066
rect 12971 2049 13002 2066
rect 13040 2049 13075 2083
rect 13109 2066 13144 2083
rect 13178 2066 13213 2083
rect 13247 2066 13282 2083
rect 13316 2066 13351 2083
rect 13385 2066 13420 2083
rect 13454 2066 13489 2083
rect 13523 2066 13558 2083
rect 13110 2049 13144 2066
rect 13184 2049 13213 2066
rect 13258 2049 13282 2066
rect 13332 2049 13351 2066
rect 13406 2049 13420 2066
rect 13480 2049 13489 2066
rect 13554 2049 13558 2066
rect 13592 2066 13627 2083
rect 13661 2066 13696 2083
rect 13730 2066 13765 2083
rect 13799 2066 13834 2083
rect 13868 2066 13903 2083
rect 13937 2066 13972 2083
rect 14006 2066 14041 2083
rect 13592 2049 13594 2066
rect 13661 2049 13668 2066
rect 13730 2049 13741 2066
rect 13799 2049 13814 2066
rect 13868 2049 13887 2066
rect 13937 2049 13960 2066
rect 14006 2049 14033 2066
rect 14075 2049 14099 2083
rect 12592 2032 12632 2049
rect 12666 2032 12706 2049
rect 12740 2032 12780 2049
rect 12814 2032 12854 2049
rect 12888 2032 12928 2049
rect 12962 2032 13002 2049
rect 13036 2032 13076 2049
rect 13110 2032 13150 2049
rect 13184 2032 13224 2049
rect 13258 2032 13298 2049
rect 13332 2032 13372 2049
rect 13406 2032 13446 2049
rect 13480 2032 13520 2049
rect 13554 2032 13594 2049
rect 13628 2032 13668 2049
rect 13702 2032 13741 2049
rect 13775 2032 13814 2049
rect 13848 2032 13887 2049
rect 13921 2032 13960 2049
rect 13994 2032 14033 2049
rect 14067 2032 14099 2049
rect 11439 2015 14099 2032
rect 11439 1994 11476 2015
rect 11510 1994 11546 2015
rect 11580 1994 11616 2015
rect 11650 1994 11686 2015
rect 11720 1994 11756 2015
rect 11790 1994 11826 2015
rect 11860 1994 11896 2015
rect 11439 1960 11448 1994
rect 11510 1981 11522 1994
rect 11580 1981 11596 1994
rect 11650 1981 11670 1994
rect 11720 1981 11744 1994
rect 11790 1981 11818 1994
rect 11860 1981 11892 1994
rect 11930 1981 11966 2015
rect 12000 1981 12036 2015
rect 12070 1994 12106 2015
rect 12140 1994 12176 2015
rect 12210 1994 12246 2015
rect 12280 1994 12316 2015
rect 12350 1994 12385 2015
rect 12419 1994 12454 2015
rect 12488 1994 12523 2015
rect 12074 1981 12106 1994
rect 12148 1981 12176 1994
rect 12222 1981 12246 1994
rect 12296 1981 12316 1994
rect 12370 1981 12385 1994
rect 12444 1981 12454 1994
rect 12518 1981 12523 1994
rect 12557 1994 12592 2015
rect 12557 1981 12558 1994
rect 11482 1960 11522 1981
rect 11556 1960 11596 1981
rect 11630 1960 11670 1981
rect 11704 1960 11744 1981
rect 11778 1960 11818 1981
rect 11852 1960 11892 1981
rect 11926 1960 11966 1981
rect 12000 1960 12040 1981
rect 12074 1960 12114 1981
rect 12148 1960 12188 1981
rect 12222 1960 12262 1981
rect 12296 1960 12336 1981
rect 12370 1960 12410 1981
rect 12444 1960 12484 1981
rect 12518 1960 12558 1981
rect 12626 1994 12661 2015
rect 12695 1994 12730 2015
rect 12764 1994 12799 2015
rect 12833 1994 12868 2015
rect 12902 1994 12937 2015
rect 12971 1994 13006 2015
rect 12626 1981 12632 1994
rect 12695 1981 12706 1994
rect 12764 1981 12780 1994
rect 12833 1981 12854 1994
rect 12902 1981 12928 1994
rect 12971 1981 13002 1994
rect 13040 1981 13075 2015
rect 13109 1994 13144 2015
rect 13178 1994 13213 2015
rect 13247 1994 13282 2015
rect 13316 1994 13351 2015
rect 13385 1994 13420 2015
rect 13454 1994 13489 2015
rect 13523 1994 13558 2015
rect 13110 1981 13144 1994
rect 13184 1981 13213 1994
rect 13258 1981 13282 1994
rect 13332 1981 13351 1994
rect 13406 1981 13420 1994
rect 13480 1981 13489 1994
rect 13554 1981 13558 1994
rect 13592 1994 13627 2015
rect 13661 1994 13696 2015
rect 13730 1994 13765 2015
rect 13799 1994 13834 2015
rect 13868 1994 13903 2015
rect 13937 1994 13972 2015
rect 14006 1994 14041 2015
rect 13592 1981 13594 1994
rect 13661 1981 13668 1994
rect 13730 1981 13741 1994
rect 13799 1981 13814 1994
rect 13868 1981 13887 1994
rect 13937 1981 13960 1994
rect 14006 1981 14033 1994
rect 14075 1981 14099 2015
rect 12592 1960 12632 1981
rect 12666 1960 12706 1981
rect 12740 1960 12780 1981
rect 12814 1960 12854 1981
rect 12888 1960 12928 1981
rect 12962 1960 13002 1981
rect 13036 1960 13076 1981
rect 13110 1960 13150 1981
rect 13184 1960 13224 1981
rect 13258 1960 13298 1981
rect 13332 1960 13372 1981
rect 13406 1960 13446 1981
rect 13480 1960 13520 1981
rect 13554 1960 13594 1981
rect 13628 1960 13668 1981
rect 13702 1960 13741 1981
rect 13775 1960 13814 1981
rect 13848 1960 13887 1981
rect 13921 1960 13960 1981
rect 13994 1960 14033 1981
rect 14067 1960 14099 1981
rect 11439 1947 14099 1960
rect 11439 1922 11476 1947
rect 11510 1922 11546 1947
rect 11580 1922 11616 1947
rect 11650 1922 11686 1947
rect 11720 1922 11756 1947
rect 11790 1922 11826 1947
rect 11860 1922 11896 1947
rect 11439 1888 11448 1922
rect 11510 1913 11522 1922
rect 11580 1913 11596 1922
rect 11650 1913 11670 1922
rect 11720 1913 11744 1922
rect 11790 1913 11818 1922
rect 11860 1913 11892 1922
rect 11930 1913 11966 1947
rect 12000 1913 12036 1947
rect 12070 1922 12106 1947
rect 12140 1922 12176 1947
rect 12210 1922 12246 1947
rect 12280 1922 12316 1947
rect 12350 1922 12385 1947
rect 12419 1922 12454 1947
rect 12488 1922 12523 1947
rect 12074 1913 12106 1922
rect 12148 1913 12176 1922
rect 12222 1913 12246 1922
rect 12296 1913 12316 1922
rect 12370 1913 12385 1922
rect 12444 1913 12454 1922
rect 12518 1913 12523 1922
rect 12557 1922 12592 1947
rect 12557 1913 12558 1922
rect 11482 1888 11522 1913
rect 11556 1888 11596 1913
rect 11630 1888 11670 1913
rect 11704 1888 11744 1913
rect 11778 1888 11818 1913
rect 11852 1888 11892 1913
rect 11926 1888 11966 1913
rect 12000 1888 12040 1913
rect 12074 1888 12114 1913
rect 12148 1888 12188 1913
rect 12222 1888 12262 1913
rect 12296 1888 12336 1913
rect 12370 1888 12410 1913
rect 12444 1888 12484 1913
rect 12518 1888 12558 1913
rect 12626 1922 12661 1947
rect 12695 1922 12730 1947
rect 12764 1922 12799 1947
rect 12833 1922 12868 1947
rect 12902 1922 12937 1947
rect 12971 1922 13006 1947
rect 12626 1913 12632 1922
rect 12695 1913 12706 1922
rect 12764 1913 12780 1922
rect 12833 1913 12854 1922
rect 12902 1913 12928 1922
rect 12971 1913 13002 1922
rect 13040 1913 13075 1947
rect 13109 1922 13144 1947
rect 13178 1922 13213 1947
rect 13247 1922 13282 1947
rect 13316 1922 13351 1947
rect 13385 1922 13420 1947
rect 13454 1922 13489 1947
rect 13523 1922 13558 1947
rect 13110 1913 13144 1922
rect 13184 1913 13213 1922
rect 13258 1913 13282 1922
rect 13332 1913 13351 1922
rect 13406 1913 13420 1922
rect 13480 1913 13489 1922
rect 13554 1913 13558 1922
rect 13592 1922 13627 1947
rect 13661 1922 13696 1947
rect 13730 1922 13765 1947
rect 13799 1922 13834 1947
rect 13868 1922 13903 1947
rect 13937 1922 13972 1947
rect 14006 1922 14041 1947
rect 13592 1913 13594 1922
rect 13661 1913 13668 1922
rect 13730 1913 13741 1922
rect 13799 1913 13814 1922
rect 13868 1913 13887 1922
rect 13937 1913 13960 1922
rect 14006 1913 14033 1922
rect 14075 1913 14099 1947
rect 12592 1888 12632 1913
rect 12666 1888 12706 1913
rect 12740 1888 12780 1913
rect 12814 1888 12854 1913
rect 12888 1888 12928 1913
rect 12962 1888 13002 1913
rect 13036 1888 13076 1913
rect 13110 1888 13150 1913
rect 13184 1888 13224 1913
rect 13258 1888 13298 1913
rect 13332 1888 13372 1913
rect 13406 1888 13446 1913
rect 13480 1888 13520 1913
rect 13554 1888 13594 1913
rect 13628 1888 13668 1913
rect 13702 1888 13741 1913
rect 13775 1888 13814 1913
rect 13848 1888 13887 1913
rect 13921 1888 13960 1913
rect 13994 1888 14033 1913
rect 14067 1888 14099 1913
rect 11439 1879 14099 1888
rect 11439 1850 11476 1879
rect 11510 1850 11546 1879
rect 11580 1850 11616 1879
rect 11650 1850 11686 1879
rect 11720 1850 11756 1879
rect 11790 1850 11826 1879
rect 11860 1850 11896 1879
rect 11439 1816 11448 1850
rect 11510 1845 11522 1850
rect 11580 1845 11596 1850
rect 11650 1845 11670 1850
rect 11720 1845 11744 1850
rect 11790 1845 11818 1850
rect 11860 1845 11892 1850
rect 11930 1845 11966 1879
rect 12000 1845 12036 1879
rect 12070 1850 12106 1879
rect 12140 1850 12176 1879
rect 12210 1850 12246 1879
rect 12280 1850 12316 1879
rect 12350 1850 12385 1879
rect 12419 1850 12454 1879
rect 12488 1850 12523 1879
rect 12074 1845 12106 1850
rect 12148 1845 12176 1850
rect 12222 1845 12246 1850
rect 12296 1845 12316 1850
rect 12370 1845 12385 1850
rect 12444 1845 12454 1850
rect 12518 1845 12523 1850
rect 12557 1850 12592 1879
rect 12557 1845 12558 1850
rect 11482 1816 11522 1845
rect 11556 1816 11596 1845
rect 11630 1816 11670 1845
rect 11704 1816 11744 1845
rect 11778 1816 11818 1845
rect 11852 1816 11892 1845
rect 11926 1816 11966 1845
rect 12000 1816 12040 1845
rect 12074 1816 12114 1845
rect 12148 1816 12188 1845
rect 12222 1816 12262 1845
rect 12296 1816 12336 1845
rect 12370 1816 12410 1845
rect 12444 1816 12484 1845
rect 12518 1816 12558 1845
rect 12626 1850 12661 1879
rect 12695 1850 12730 1879
rect 12764 1850 12799 1879
rect 12833 1850 12868 1879
rect 12902 1850 12937 1879
rect 12971 1850 13006 1879
rect 12626 1845 12632 1850
rect 12695 1845 12706 1850
rect 12764 1845 12780 1850
rect 12833 1845 12854 1850
rect 12902 1845 12928 1850
rect 12971 1845 13002 1850
rect 13040 1845 13075 1879
rect 13109 1850 13144 1879
rect 13178 1850 13213 1879
rect 13247 1850 13282 1879
rect 13316 1850 13351 1879
rect 13385 1850 13420 1879
rect 13454 1850 13489 1879
rect 13523 1850 13558 1879
rect 13110 1845 13144 1850
rect 13184 1845 13213 1850
rect 13258 1845 13282 1850
rect 13332 1845 13351 1850
rect 13406 1845 13420 1850
rect 13480 1845 13489 1850
rect 13554 1845 13558 1850
rect 13592 1850 13627 1879
rect 13661 1850 13696 1879
rect 13730 1850 13765 1879
rect 13799 1850 13834 1879
rect 13868 1850 13903 1879
rect 13937 1850 13972 1879
rect 14006 1850 14041 1879
rect 13592 1845 13594 1850
rect 13661 1845 13668 1850
rect 13730 1845 13741 1850
rect 13799 1845 13814 1850
rect 13868 1845 13887 1850
rect 13937 1845 13960 1850
rect 14006 1845 14033 1850
rect 14075 1845 14099 1879
rect 12592 1816 12632 1845
rect 12666 1816 12706 1845
rect 12740 1816 12780 1845
rect 12814 1816 12854 1845
rect 12888 1816 12928 1845
rect 12962 1816 13002 1845
rect 13036 1816 13076 1845
rect 13110 1816 13150 1845
rect 13184 1816 13224 1845
rect 13258 1816 13298 1845
rect 13332 1816 13372 1845
rect 13406 1816 13446 1845
rect 13480 1816 13520 1845
rect 13554 1816 13594 1845
rect 13628 1816 13668 1845
rect 13702 1816 13741 1845
rect 13775 1816 13814 1845
rect 13848 1816 13887 1845
rect 13921 1816 13960 1845
rect 13994 1816 14033 1845
rect 14067 1816 14099 1845
rect 11439 1811 14099 1816
rect 11439 1778 11476 1811
rect 11510 1778 11546 1811
rect 11580 1778 11616 1811
rect 11650 1778 11686 1811
rect 11720 1778 11756 1811
rect 11790 1778 11826 1811
rect 11860 1778 11896 1811
rect 11439 1744 11448 1778
rect 11510 1777 11522 1778
rect 11580 1777 11596 1778
rect 11650 1777 11670 1778
rect 11720 1777 11744 1778
rect 11790 1777 11818 1778
rect 11860 1777 11892 1778
rect 11930 1777 11966 1811
rect 12000 1777 12036 1811
rect 12070 1778 12106 1811
rect 12140 1778 12176 1811
rect 12210 1778 12246 1811
rect 12280 1778 12316 1811
rect 12350 1778 12385 1811
rect 12419 1778 12454 1811
rect 12488 1778 12523 1811
rect 12074 1777 12106 1778
rect 12148 1777 12176 1778
rect 12222 1777 12246 1778
rect 12296 1777 12316 1778
rect 12370 1777 12385 1778
rect 12444 1777 12454 1778
rect 12518 1777 12523 1778
rect 12557 1778 12592 1811
rect 12557 1777 12558 1778
rect 11482 1744 11522 1777
rect 11556 1744 11596 1777
rect 11630 1744 11670 1777
rect 11704 1744 11744 1777
rect 11778 1744 11818 1777
rect 11852 1744 11892 1777
rect 11926 1744 11966 1777
rect 12000 1744 12040 1777
rect 12074 1744 12114 1777
rect 12148 1744 12188 1777
rect 12222 1744 12262 1777
rect 12296 1744 12336 1777
rect 12370 1744 12410 1777
rect 12444 1744 12484 1777
rect 12518 1744 12558 1777
rect 12626 1778 12661 1811
rect 12695 1778 12730 1811
rect 12764 1778 12799 1811
rect 12833 1778 12868 1811
rect 12902 1778 12937 1811
rect 12971 1778 13006 1811
rect 12626 1777 12632 1778
rect 12695 1777 12706 1778
rect 12764 1777 12780 1778
rect 12833 1777 12854 1778
rect 12902 1777 12928 1778
rect 12971 1777 13002 1778
rect 13040 1777 13075 1811
rect 13109 1778 13144 1811
rect 13178 1778 13213 1811
rect 13247 1778 13282 1811
rect 13316 1778 13351 1811
rect 13385 1778 13420 1811
rect 13454 1778 13489 1811
rect 13523 1778 13558 1811
rect 13110 1777 13144 1778
rect 13184 1777 13213 1778
rect 13258 1777 13282 1778
rect 13332 1777 13351 1778
rect 13406 1777 13420 1778
rect 13480 1777 13489 1778
rect 13554 1777 13558 1778
rect 13592 1778 13627 1811
rect 13661 1778 13696 1811
rect 13730 1778 13765 1811
rect 13799 1778 13834 1811
rect 13868 1778 13903 1811
rect 13937 1778 13972 1811
rect 14006 1778 14041 1811
rect 13592 1777 13594 1778
rect 13661 1777 13668 1778
rect 13730 1777 13741 1778
rect 13799 1777 13814 1778
rect 13868 1777 13887 1778
rect 13937 1777 13960 1778
rect 14006 1777 14033 1778
rect 14075 1777 14099 1811
rect 12592 1744 12632 1777
rect 12666 1744 12706 1777
rect 12740 1744 12780 1777
rect 12814 1744 12854 1777
rect 12888 1744 12928 1777
rect 12962 1744 13002 1777
rect 13036 1744 13076 1777
rect 13110 1744 13150 1777
rect 13184 1744 13224 1777
rect 13258 1744 13298 1777
rect 13332 1744 13372 1777
rect 13406 1744 13446 1777
rect 13480 1744 13520 1777
rect 13554 1744 13594 1777
rect 13628 1744 13668 1777
rect 13702 1744 13741 1777
rect 13775 1744 13814 1777
rect 13848 1744 13887 1777
rect 13921 1744 13960 1777
rect 13994 1744 14033 1777
rect 14067 1744 14099 1777
rect 11439 1743 14099 1744
rect 11439 1709 11476 1743
rect 11510 1709 11546 1743
rect 11580 1709 11616 1743
rect 11650 1709 11686 1743
rect 11720 1709 11756 1743
rect 11790 1709 11826 1743
rect 11860 1709 11896 1743
rect 11930 1709 11966 1743
rect 12000 1709 12036 1743
rect 12070 1709 12106 1743
rect 12140 1709 12176 1743
rect 12210 1709 12246 1743
rect 12280 1709 12316 1743
rect 12350 1709 12385 1743
rect 12419 1709 12454 1743
rect 12488 1709 12523 1743
rect 12557 1709 12592 1743
rect 12626 1709 12661 1743
rect 12695 1709 12730 1743
rect 12764 1709 12799 1743
rect 12833 1709 12868 1743
rect 12902 1709 12937 1743
rect 12971 1709 13006 1743
rect 13040 1709 13075 1743
rect 13109 1709 13144 1743
rect 13178 1709 13213 1743
rect 13247 1709 13282 1743
rect 13316 1709 13351 1743
rect 13385 1709 13420 1743
rect 13454 1709 13489 1743
rect 13523 1709 13558 1743
rect 13592 1709 13627 1743
rect 13661 1709 13696 1743
rect 13730 1709 13765 1743
rect 13799 1709 13834 1743
rect 13868 1709 13903 1743
rect 13937 1709 13972 1743
rect 14006 1709 14041 1743
rect 14075 1709 14099 1743
rect 11439 1675 14099 1709
rect 11439 1641 11476 1675
rect 11510 1641 11546 1675
rect 11580 1641 11616 1675
rect 11650 1641 11686 1675
rect 11720 1641 11756 1675
rect 11790 1641 11826 1675
rect 11860 1641 11896 1675
rect 11930 1641 11966 1675
rect 12000 1641 12036 1675
rect 12070 1641 12106 1675
rect 12140 1641 12176 1675
rect 12210 1641 12246 1675
rect 12280 1641 12316 1675
rect 12350 1641 12385 1675
rect 12419 1641 12454 1675
rect 12488 1641 12523 1675
rect 12557 1641 12592 1675
rect 12626 1641 12661 1675
rect 12695 1641 12730 1675
rect 12764 1641 12799 1675
rect 12833 1641 12868 1675
rect 12902 1641 12937 1675
rect 12971 1641 13006 1675
rect 13040 1641 13075 1675
rect 13109 1641 13144 1675
rect 13178 1641 13213 1675
rect 13247 1641 13282 1675
rect 13316 1641 13351 1675
rect 13385 1641 13420 1675
rect 13454 1641 13489 1675
rect 13523 1641 13558 1675
rect 13592 1641 13627 1675
rect 13661 1641 13696 1675
rect 13730 1641 13765 1675
rect 13799 1641 13834 1675
rect 13868 1641 13903 1675
rect 13937 1641 13972 1675
rect 14006 1641 14041 1675
rect 14075 1641 14099 1675
rect 11439 1566 14099 1641
rect 11439 1532 12957 1566
rect 12991 1532 13030 1566
rect 13064 1532 13103 1566
rect 13137 1532 13176 1566
rect 13210 1532 13249 1566
rect 13283 1532 13321 1566
rect 13355 1532 13393 1566
rect 13427 1532 13465 1566
rect 13499 1532 13537 1566
rect 13571 1532 13609 1566
rect 13643 1532 13681 1566
rect 13715 1532 13753 1566
rect 13787 1532 13825 1566
rect 13859 1532 13897 1566
rect 13931 1532 13969 1566
rect 14003 1532 14041 1566
rect 14075 1532 14099 1566
rect 11439 1498 14099 1532
rect 11439 1464 12957 1498
rect 12991 1464 13030 1498
rect 13064 1464 13103 1498
rect 13137 1464 13176 1498
rect 13210 1464 13249 1498
rect 13283 1464 13321 1498
rect 13355 1464 13393 1498
rect 13427 1464 13465 1498
rect 13499 1464 13537 1498
rect 13571 1464 13609 1498
rect 13643 1464 13681 1498
rect 13715 1464 13753 1498
rect 13787 1464 13825 1498
rect 13859 1464 13897 1498
rect 13931 1464 13969 1498
rect 14003 1464 14041 1498
rect 14075 1464 14099 1498
rect 11439 1430 14099 1464
rect 11439 1396 12957 1430
rect 12991 1396 13030 1430
rect 13064 1396 13103 1430
rect 13137 1396 13176 1430
rect 13210 1396 13249 1430
rect 13283 1396 13321 1430
rect 13355 1396 13393 1430
rect 13427 1396 13465 1430
rect 13499 1396 13537 1430
rect 13571 1396 13609 1430
rect 13643 1396 13681 1430
rect 13715 1396 13753 1430
rect 13787 1396 13825 1430
rect 13859 1396 13897 1430
rect 13931 1396 13969 1430
rect 14003 1396 14041 1430
rect 14075 1396 14099 1430
rect 11116 106 11252 140
rect 11116 64 11286 106
rect 7664 0 11286 64
<< viali >>
rect 74 6433 108 6467
rect 146 6433 180 6467
rect 218 6433 252 6467
rect 290 6433 324 6467
rect 362 6433 396 6467
rect 434 6433 468 6467
rect 506 6433 540 6467
rect 578 6433 612 6467
rect 650 6433 684 6467
rect 722 6433 756 6467
rect 794 6433 828 6467
rect 866 6433 900 6467
rect 938 6433 972 6467
rect 1010 6433 1044 6467
rect 1082 6433 1116 6467
rect 1154 6433 1188 6467
rect 1226 6433 1260 6467
rect 1298 6433 1332 6467
rect 1370 6433 1404 6467
rect 1442 6433 1476 6467
rect 1514 6433 1548 6467
rect 1586 6433 1620 6467
rect 1658 6433 1692 6467
rect 1730 6433 1764 6467
rect 1802 6433 1836 6467
rect 1874 6433 1908 6467
rect 1946 6433 1980 6467
rect 2018 6433 2052 6467
rect 2090 6433 2124 6467
rect 2162 6433 2196 6467
rect 2234 6433 2268 6467
rect 2306 6433 2340 6467
rect 2378 6433 2412 6467
rect 2450 6433 2484 6467
rect 2522 6433 2556 6467
rect 2594 6433 2628 6467
rect 2666 6433 2700 6467
rect 2738 6433 2772 6467
rect 2810 6433 2844 6467
rect 2882 6433 2916 6467
rect 2954 6433 2988 6467
rect 3026 6433 3060 6467
rect 3098 6433 3132 6467
rect 3170 6433 3204 6467
rect 3242 6433 3276 6467
rect 3314 6433 3348 6467
rect 3386 6433 3420 6467
rect 3458 6433 3492 6467
rect 3530 6433 3564 6467
rect 3602 6433 3636 6467
rect 3674 6433 3708 6467
rect 3746 6433 3780 6467
rect 3818 6433 3852 6467
rect 3890 6433 3924 6467
rect 3962 6433 3996 6467
rect 4034 6433 4068 6467
rect 4106 6433 4140 6467
rect 4178 6433 4212 6467
rect 4250 6433 4284 6467
rect 4322 6433 4356 6467
rect 4394 6433 4428 6467
rect 4466 6433 4500 6467
rect 4538 6433 4572 6467
rect 4610 6433 4644 6467
rect 4682 6433 4716 6467
rect 4754 6433 4788 6467
rect 4826 6433 4860 6467
rect 4898 6433 4932 6467
rect 4971 6433 5005 6467
rect 5044 6433 5078 6467
rect 5117 6433 5151 6467
rect 5190 6433 5224 6467
rect 5263 6433 5297 6467
rect 5336 6433 5370 6467
rect 5409 6433 5443 6467
rect 5482 6433 5516 6467
rect 5555 6433 5589 6467
rect 5628 6433 5662 6467
rect 5701 6433 5735 6467
rect 5774 6433 5808 6467
rect 5847 6433 5881 6467
rect 5920 6433 5954 6467
rect 5993 6433 6027 6467
rect 6066 6433 6100 6467
rect 6139 6433 6173 6467
rect 6212 6433 6246 6467
rect 6285 6433 6319 6467
rect 6358 6433 6392 6467
rect 6431 6433 6465 6467
rect 6504 6433 6538 6467
rect 6577 6433 6611 6467
rect 6650 6433 6684 6467
rect 6723 6433 6757 6467
rect 6796 6433 6830 6467
rect 6869 6433 6903 6467
rect 6942 6433 6976 6467
rect 7015 6433 7049 6467
rect 7088 6433 7122 6467
rect 7161 6433 7195 6467
rect 7234 6433 7268 6467
rect 7307 6433 7341 6467
rect 7380 6433 7414 6467
rect 7453 6433 7487 6467
rect 7526 6433 7560 6467
rect 7599 6433 7633 6467
rect 7672 6433 7706 6467
rect 7745 6433 7779 6467
rect 7818 6433 7852 6467
rect 7891 6433 7925 6467
rect 7964 6433 7998 6467
rect 8037 6433 8071 6467
rect 8110 6433 8144 6467
rect 8183 6433 8217 6467
rect 8256 6433 8290 6467
rect 8329 6433 8363 6467
rect 8402 6433 8436 6467
rect 8475 6433 8509 6467
rect 8548 6433 8582 6467
rect 8621 6433 8655 6467
rect 8694 6433 8728 6467
rect 8767 6433 8801 6467
rect 8840 6433 8874 6467
rect 8913 6433 8947 6467
rect 8986 6433 9020 6467
rect 9059 6433 9093 6467
rect 9132 6433 9166 6467
rect 9205 6433 9239 6467
rect 9278 6433 9312 6467
rect 9351 6433 9385 6467
rect 9424 6433 9458 6467
rect 9497 6433 9531 6467
rect 9570 6433 9604 6467
rect 9643 6433 9677 6467
rect 9716 6433 9750 6467
rect 9789 6433 9823 6467
rect 9862 6433 9896 6467
rect 68 6361 102 6395
rect 68 6289 102 6323
rect 68 6217 102 6251
rect 68 6145 102 6179
rect 68 6073 102 6107
rect 68 6001 102 6035
rect 68 5929 102 5963
rect 68 5857 102 5891
rect 68 5785 102 5819
rect 68 5713 102 5747
rect 68 5641 102 5675
rect 68 5569 102 5603
rect 68 5497 102 5531
rect 68 5425 102 5459
rect 68 5353 102 5387
rect 68 5281 102 5315
rect 68 5209 102 5243
rect 68 5137 102 5171
rect 68 5065 102 5099
rect 68 4993 102 5027
rect 68 4921 102 4955
rect 68 4848 102 4882
rect 68 4775 102 4809
rect 68 4702 102 4736
rect 68 4629 102 4663
rect 68 4556 102 4590
rect 68 4483 102 4517
rect 68 4410 102 4444
rect 68 4337 102 4371
rect 68 4264 102 4298
rect 68 4191 102 4225
rect 68 4118 102 4152
rect 68 4045 102 4079
rect 68 3972 102 4006
rect 68 3899 102 3933
rect 68 3826 102 3860
rect 68 3753 102 3787
rect 68 3680 102 3714
rect 68 3607 102 3641
rect 68 3534 102 3568
rect 68 3461 102 3495
rect 323 6066 357 6094
rect 395 6066 429 6100
rect 473 6066 483 6100
rect 483 6066 507 6100
rect 551 6066 585 6100
rect 629 6066 653 6100
rect 653 6066 663 6100
rect 707 6066 721 6100
rect 721 6066 741 6100
rect 784 6066 789 6100
rect 789 6066 818 6100
rect 950 6066 959 6100
rect 959 6066 984 6100
rect 1027 6066 1061 6100
rect 1104 6066 1129 6100
rect 1129 6066 1138 6100
rect 1181 6066 1197 6100
rect 1197 6066 1215 6100
rect 1258 6066 1265 6100
rect 1265 6066 1292 6100
rect 1335 6066 1367 6100
rect 1367 6066 1369 6100
rect 1412 6066 1435 6100
rect 1435 6066 1446 6100
rect 1488 6066 1503 6100
rect 1503 6066 1522 6100
rect 1564 6066 1571 6100
rect 1571 6066 1598 6100
rect 1640 6066 1673 6100
rect 1673 6066 1674 6100
rect 1806 6066 1809 6100
rect 1809 6066 1840 6100
rect 1883 6066 1911 6100
rect 1911 6066 1917 6100
rect 1960 6066 1979 6100
rect 1979 6066 1994 6100
rect 2037 6066 2047 6100
rect 2047 6066 2071 6100
rect 2114 6066 2115 6100
rect 2115 6066 2148 6100
rect 2191 6066 2217 6100
rect 2217 6066 2225 6100
rect 2268 6066 2285 6100
rect 2285 6066 2302 6100
rect 2344 6066 2353 6100
rect 2353 6066 2378 6100
rect 2420 6066 2421 6100
rect 2421 6066 2454 6100
rect 2496 6066 2523 6100
rect 2523 6066 2530 6100
rect 2662 6066 2693 6100
rect 2693 6066 2696 6100
rect 2739 6066 2761 6100
rect 2761 6066 2773 6100
rect 2816 6066 2829 6100
rect 2829 6066 2850 6100
rect 2893 6066 2897 6100
rect 2897 6066 2927 6100
rect 2970 6066 2999 6100
rect 2999 6066 3004 6100
rect 3047 6066 3067 6100
rect 3067 6066 3081 6100
rect 3124 6066 3135 6100
rect 3135 6066 3158 6100
rect 3200 6066 3203 6100
rect 3203 6066 3234 6100
rect 3276 6066 3305 6100
rect 3305 6066 3310 6100
rect 3352 6066 3373 6100
rect 3373 6066 3386 6100
rect 3518 6066 3543 6100
rect 3543 6066 3552 6100
rect 3595 6066 3611 6100
rect 3611 6066 3629 6100
rect 3671 6066 3679 6100
rect 3679 6066 3705 6100
rect 3747 6066 3781 6100
rect 3823 6066 3849 6100
rect 3849 6066 3857 6100
rect 3899 6066 3917 6100
rect 3917 6066 3933 6100
rect 3975 6066 3985 6100
rect 3985 6066 4009 6100
rect 4051 6066 4053 6100
rect 4053 6066 4085 6100
rect 4127 6066 4155 6100
rect 4155 6066 4161 6100
rect 4203 6066 4223 6100
rect 4223 6066 4237 6100
rect 4379 6066 4393 6100
rect 4393 6066 4413 6100
rect 4455 6066 4461 6100
rect 4461 6066 4489 6100
rect 4531 6066 4563 6100
rect 4563 6066 4565 6100
rect 4607 6066 4631 6100
rect 4631 6066 4641 6100
rect 4683 6066 4699 6100
rect 4699 6066 4717 6100
rect 4759 6066 4767 6100
rect 4767 6066 4793 6100
rect 4831 6066 4835 6094
rect 4835 6066 4937 6094
rect 4987 6066 4989 6100
rect 4989 6066 5021 6100
rect 5061 6066 5091 6100
rect 5091 6066 5095 6100
rect 5135 6066 5159 6100
rect 5159 6066 5169 6100
rect 5209 6066 5227 6100
rect 5227 6066 5243 6100
rect 5283 6066 5295 6100
rect 5295 6066 5317 6100
rect 5357 6066 5363 6100
rect 5363 6066 5391 6100
rect 5431 6066 5465 6100
rect 5505 6066 5533 6100
rect 5533 6066 5539 6100
rect 5579 6066 5601 6100
rect 5601 6066 5613 6100
rect 5652 6066 5669 6100
rect 5669 6066 5686 6100
rect 5725 6066 5737 6100
rect 5737 6066 5759 6100
rect 5798 6066 5805 6100
rect 5805 6066 5832 6100
rect 5871 6066 5873 6100
rect 5873 6066 5905 6100
rect 5944 6066 5975 6100
rect 5975 6066 5978 6100
rect 6017 6066 6043 6100
rect 6043 6066 6051 6100
rect 6090 6066 6111 6100
rect 6111 6066 6124 6100
rect 6163 6066 6179 6100
rect 6179 6066 6197 6100
rect 6236 6066 6247 6100
rect 6247 6066 6270 6100
rect 6309 6066 6315 6100
rect 6315 6066 6343 6100
rect 6382 6066 6383 6100
rect 6383 6066 6416 6100
rect 6455 6066 6485 6100
rect 6485 6066 6489 6100
rect 6528 6066 6553 6100
rect 6553 6066 6562 6100
rect 6601 6066 6621 6100
rect 6621 6066 6635 6100
rect 6674 6066 6689 6100
rect 6689 6066 6708 6100
rect 6747 6066 6757 6100
rect 6757 6066 6781 6100
rect 6820 6066 6825 6100
rect 6825 6066 6854 6100
rect 6893 6066 6927 6100
rect 6966 6066 6995 6100
rect 6995 6066 7000 6100
rect 7039 6066 7063 6100
rect 7063 6066 7073 6100
rect 7112 6066 7131 6100
rect 7131 6066 7146 6100
rect 7185 6066 7199 6100
rect 7199 6066 7219 6100
rect 7258 6066 7267 6100
rect 7267 6066 7292 6100
rect 7331 6066 7335 6100
rect 7335 6066 7365 6100
rect 323 6060 357 6066
rect 323 5998 357 6022
rect 323 5988 357 5998
rect 323 5930 357 5950
rect 323 5916 357 5930
rect 323 5862 357 5878
rect 323 5844 357 5862
rect 4831 6032 4915 6066
rect 4915 6032 4937 6066
rect 4831 5998 4937 6032
rect 4831 5970 4915 5998
rect 4831 5936 4835 5970
rect 4835 5936 4869 5970
rect 4869 5964 4915 5970
rect 4915 5964 4937 5998
rect 4869 5936 4937 5964
rect 4831 5930 4937 5936
rect 4831 5902 4915 5930
rect 4831 5868 4835 5902
rect 4835 5868 4869 5902
rect 4869 5896 4915 5902
rect 4915 5896 4937 5930
rect 4869 5868 4937 5896
rect 4831 5862 4937 5868
rect 696 5825 730 5859
rect 781 5825 815 5859
rect 866 5825 900 5859
rect 952 5825 986 5859
rect 1038 5825 1072 5859
rect 1552 5825 1586 5859
rect 1637 5825 1671 5859
rect 1722 5825 1756 5859
rect 1808 5825 1842 5859
rect 1894 5825 1928 5859
rect 2408 5825 2434 5859
rect 2434 5825 2442 5859
rect 2493 5825 2508 5859
rect 2508 5825 2527 5859
rect 2578 5825 2581 5859
rect 2581 5825 2612 5859
rect 2664 5825 2688 5859
rect 2688 5825 2698 5859
rect 2750 5825 2761 5859
rect 2761 5825 2784 5859
rect 3264 5825 3278 5859
rect 3278 5825 3298 5859
rect 3349 5825 3381 5859
rect 3381 5825 3383 5859
rect 3434 5825 3450 5859
rect 3450 5825 3468 5859
rect 3520 5825 3554 5859
rect 3606 5825 3623 5859
rect 3623 5825 3640 5859
rect 4120 5825 4140 5859
rect 4140 5825 4154 5859
rect 4205 5825 4209 5859
rect 4209 5825 4239 5859
rect 4290 5825 4313 5859
rect 4313 5825 4324 5859
rect 4376 5825 4382 5859
rect 4382 5825 4410 5859
rect 4462 5825 4485 5859
rect 4485 5825 4496 5859
rect 4831 5834 4915 5862
rect 323 5794 357 5806
rect 323 5772 357 5794
rect 323 5726 357 5734
rect 4831 5800 4835 5834
rect 4835 5800 4869 5834
rect 4869 5828 4915 5834
rect 4915 5828 4937 5862
rect 4869 5800 4937 5828
rect 4831 5794 4937 5800
rect 4831 5766 4915 5794
rect 4831 5732 4835 5766
rect 4835 5732 4869 5766
rect 4869 5760 4915 5766
rect 4915 5760 4937 5794
rect 4869 5732 4937 5760
rect 323 5700 357 5726
rect 323 5658 357 5662
rect 323 5628 357 5658
rect 323 5556 357 5590
rect 323 5488 357 5518
rect 323 5484 357 5488
rect 323 5420 357 5446
rect 323 5412 357 5420
rect 323 5352 357 5374
rect 323 5340 357 5352
rect 323 5284 357 5302
rect 323 5268 357 5284
rect 323 5216 357 5230
rect 323 5196 357 5216
rect 323 5148 357 5158
rect 323 5124 357 5148
rect 323 5080 357 5086
rect 323 5052 357 5080
rect 323 5012 357 5014
rect 323 4980 357 5012
rect 323 4910 357 4942
rect 323 4908 357 4910
rect 323 4842 357 4870
rect 323 4836 357 4842
rect 323 4774 357 4798
rect 323 4764 357 4774
rect 323 4706 357 4726
rect 323 4692 357 4706
rect 323 4638 357 4654
rect 323 4620 357 4638
rect 323 4570 357 4582
rect 323 4548 357 4570
rect 323 4502 357 4510
rect 323 4476 357 4502
rect 323 4434 357 4438
rect 323 4404 357 4434
rect 323 4332 357 4366
rect 323 4264 357 4294
rect 323 4260 357 4264
rect 323 4196 357 4222
rect 323 4188 357 4196
rect 323 4128 357 4150
rect 323 4116 357 4128
rect 323 4060 357 4078
rect 323 4044 357 4060
rect 323 3992 357 4005
rect 323 3971 357 3992
rect 323 3924 357 3932
rect 323 3898 357 3924
rect 323 3856 357 3859
rect 323 3825 357 3856
rect 323 3754 357 3786
rect 439 5697 473 5731
rect 439 5624 473 5658
rect 439 5551 473 5585
rect 439 5478 473 5512
rect 439 5405 473 5439
rect 439 5332 473 5366
rect 439 5259 473 5293
rect 439 5186 473 5220
rect 439 5113 473 5147
rect 439 5040 473 5074
rect 439 4967 473 5001
rect 439 4894 473 4928
rect 439 4821 473 4855
rect 439 4747 473 4781
rect 439 4673 473 4707
rect 439 4599 473 4633
rect 439 4525 473 4559
rect 439 4451 473 4485
rect 439 4377 473 4411
rect 439 4303 473 4337
rect 439 4229 473 4263
rect 439 4155 473 4189
rect 439 4081 473 4115
rect 439 4007 473 4041
rect 439 3933 473 3967
rect 439 3859 473 3893
rect 439 3785 473 3819
rect 1295 5697 1329 5731
rect 1295 5624 1329 5658
rect 1295 5551 1329 5585
rect 1295 5478 1329 5512
rect 1295 5405 1329 5439
rect 1295 5332 1329 5366
rect 1295 5259 1329 5293
rect 1295 5186 1329 5220
rect 1295 5113 1329 5147
rect 1295 5040 1329 5074
rect 1295 4967 1329 5001
rect 1295 4894 1329 4928
rect 1295 4821 1329 4855
rect 1295 4747 1329 4781
rect 1295 4673 1329 4707
rect 1295 4599 1329 4633
rect 1295 4525 1329 4559
rect 1295 4451 1329 4485
rect 1295 4377 1329 4411
rect 1295 4303 1329 4337
rect 1295 4229 1329 4263
rect 1295 4155 1329 4189
rect 1295 4081 1329 4115
rect 1295 4007 1329 4041
rect 1295 3933 1329 3967
rect 1295 3859 1329 3893
rect 1295 3785 1329 3819
rect 2151 5697 2185 5731
rect 2151 5624 2185 5658
rect 2151 5551 2185 5585
rect 2151 5478 2185 5512
rect 2151 5405 2185 5439
rect 2151 5332 2185 5366
rect 2151 5259 2185 5293
rect 2151 5186 2185 5220
rect 2151 5113 2185 5147
rect 2151 5040 2185 5074
rect 2151 4967 2185 5001
rect 2151 4894 2185 4928
rect 2151 4821 2185 4855
rect 2151 4747 2185 4781
rect 2151 4673 2185 4707
rect 2151 4599 2185 4633
rect 2151 4525 2185 4559
rect 2151 4451 2185 4485
rect 2151 4377 2185 4411
rect 2151 4303 2185 4337
rect 2151 4229 2185 4263
rect 2151 4155 2185 4189
rect 2151 4081 2185 4115
rect 2151 4007 2185 4041
rect 2151 3933 2185 3967
rect 2151 3859 2185 3893
rect 2151 3785 2185 3819
rect 3007 5697 3041 5731
rect 3007 5624 3041 5658
rect 3007 5551 3041 5585
rect 3007 5478 3041 5512
rect 3007 5405 3041 5439
rect 3007 5332 3041 5366
rect 3007 5259 3041 5293
rect 3007 5186 3041 5220
rect 3007 5113 3041 5147
rect 3007 5040 3041 5074
rect 3007 4967 3041 5001
rect 3007 4894 3041 4928
rect 3007 4821 3041 4855
rect 3007 4747 3041 4781
rect 3007 4673 3041 4707
rect 3007 4599 3041 4633
rect 3007 4525 3041 4559
rect 3007 4451 3041 4485
rect 3007 4377 3041 4411
rect 3007 4303 3041 4337
rect 3007 4229 3041 4263
rect 3007 4155 3041 4189
rect 3007 4081 3041 4115
rect 3007 4007 3041 4041
rect 3007 3933 3041 3967
rect 3007 3859 3041 3893
rect 3007 3785 3041 3819
rect 3863 5697 3897 5731
rect 3863 5624 3897 5658
rect 3863 5551 3897 5585
rect 3863 5478 3897 5512
rect 3863 5405 3897 5439
rect 3863 5332 3897 5366
rect 3863 5259 3897 5293
rect 3863 5186 3897 5220
rect 3863 5113 3897 5147
rect 3863 5040 3897 5074
rect 3863 4967 3897 5001
rect 3863 4894 3897 4928
rect 3863 4821 3897 4855
rect 3863 4747 3897 4781
rect 3863 4673 3897 4707
rect 3863 4599 3897 4633
rect 3863 4525 3897 4559
rect 3863 4451 3897 4485
rect 3863 4377 3897 4411
rect 3863 4303 3897 4337
rect 3863 4229 3897 4263
rect 3863 4155 3897 4189
rect 3863 4081 3897 4115
rect 3863 4007 3897 4041
rect 3863 3933 3897 3967
rect 3863 3859 3897 3893
rect 3863 3785 3897 3819
rect 4719 5697 4753 5731
rect 4719 5624 4753 5658
rect 4719 5551 4753 5585
rect 4719 5478 4753 5512
rect 4719 5405 4753 5439
rect 4719 5332 4753 5366
rect 4719 5259 4753 5293
rect 4719 5186 4753 5220
rect 4719 5113 4753 5147
rect 4719 5040 4753 5074
rect 4719 4967 4753 5001
rect 4719 4894 4753 4928
rect 4719 4821 4753 4855
rect 4719 4747 4753 4781
rect 4719 4673 4753 4707
rect 4719 4599 4753 4633
rect 4719 4525 4753 4559
rect 4719 4451 4753 4485
rect 4719 4377 4753 4411
rect 4719 4303 4753 4337
rect 4719 4229 4753 4263
rect 4719 4155 4753 4189
rect 4719 4081 4753 4115
rect 4719 4007 4753 4041
rect 4719 3933 4753 3967
rect 4719 3859 4753 3893
rect 4719 3785 4753 3819
rect 4831 5726 4937 5732
rect 4831 5698 4915 5726
rect 4831 5664 4835 5698
rect 4835 5664 4869 5698
rect 4869 5692 4915 5698
rect 4915 5692 4937 5726
rect 4869 5664 4937 5692
rect 4831 5658 4937 5664
rect 4831 5630 4915 5658
rect 4831 5596 4835 5630
rect 4835 5596 4869 5630
rect 4869 5624 4915 5630
rect 4915 5624 4937 5658
rect 4869 5596 4937 5624
rect 4831 5590 4937 5596
rect 4831 5562 4915 5590
rect 4831 5528 4835 5562
rect 4835 5528 4869 5562
rect 4869 5556 4915 5562
rect 4915 5556 4937 5590
rect 4869 5528 4937 5556
rect 4831 5522 4937 5528
rect 4831 5494 4915 5522
rect 4831 5460 4835 5494
rect 4835 5460 4869 5494
rect 4869 5488 4915 5494
rect 4915 5488 4937 5522
rect 4869 5460 4937 5488
rect 4831 5454 4937 5460
rect 4831 5426 4915 5454
rect 4831 5392 4835 5426
rect 4835 5392 4869 5426
rect 4869 5420 4915 5426
rect 4915 5420 4937 5454
rect 4869 5392 4937 5420
rect 4831 5386 4937 5392
rect 4831 5358 4915 5386
rect 4831 5324 4835 5358
rect 4835 5324 4869 5358
rect 4869 5352 4915 5358
rect 4915 5352 4937 5386
rect 4869 5324 4937 5352
rect 4831 5318 4937 5324
rect 4831 5290 4915 5318
rect 4831 5256 4835 5290
rect 4835 5256 4869 5290
rect 4869 5284 4915 5290
rect 4915 5284 4937 5318
rect 4869 5256 4937 5284
rect 4831 5250 4937 5256
rect 4831 5222 4915 5250
rect 4831 5188 4835 5222
rect 4835 5188 4869 5222
rect 4869 5216 4915 5222
rect 4915 5216 4937 5250
rect 4869 5188 4937 5216
rect 4831 5182 4937 5188
rect 4831 5154 4915 5182
rect 4831 5120 4835 5154
rect 4835 5120 4869 5154
rect 4869 5148 4915 5154
rect 4915 5148 4937 5182
rect 4869 5120 4937 5148
rect 4831 5114 4937 5120
rect 4831 5086 4915 5114
rect 4831 5052 4835 5086
rect 4835 5052 4869 5086
rect 4869 5080 4915 5086
rect 4915 5080 4937 5114
rect 4869 5052 4937 5080
rect 4831 5046 4937 5052
rect 4831 5018 4915 5046
rect 4831 4984 4835 5018
rect 4835 4984 4869 5018
rect 4869 5012 4915 5018
rect 4915 5012 4937 5046
rect 4869 4984 4937 5012
rect 4831 4978 4937 4984
rect 4831 4950 4915 4978
rect 4831 4916 4835 4950
rect 4835 4916 4869 4950
rect 4869 4944 4915 4950
rect 4915 4944 4937 4978
rect 4869 4916 4937 4944
rect 4831 4910 4937 4916
rect 4831 4882 4915 4910
rect 4831 4848 4835 4882
rect 4835 4848 4869 4882
rect 4869 4876 4915 4882
rect 4915 4876 4937 4910
rect 4869 4848 4937 4876
rect 4831 4842 4937 4848
rect 4831 4814 4915 4842
rect 4831 4780 4835 4814
rect 4835 4780 4869 4814
rect 4869 4808 4915 4814
rect 4915 4808 4937 4842
rect 4869 4780 4937 4808
rect 4831 4774 4937 4780
rect 4831 4746 4915 4774
rect 4831 4712 4835 4746
rect 4835 4712 4869 4746
rect 4869 4740 4915 4746
rect 4915 4740 4937 4774
rect 4869 4712 4937 4740
rect 4831 4706 4937 4712
rect 4831 4678 4915 4706
rect 4831 4644 4835 4678
rect 4835 4644 4869 4678
rect 4869 4672 4915 4678
rect 4915 4672 4937 4706
rect 4869 4644 4937 4672
rect 4831 4638 4937 4644
rect 4831 4610 4915 4638
rect 4831 4576 4835 4610
rect 4835 4576 4869 4610
rect 4869 4604 4915 4610
rect 4915 4604 4937 4638
rect 4869 4576 4937 4604
rect 4831 4570 4937 4576
rect 4831 4542 4915 4570
rect 4831 4508 4835 4542
rect 4835 4508 4869 4542
rect 4869 4536 4915 4542
rect 4915 4536 4937 4570
rect 4869 4508 4937 4536
rect 4831 4502 4937 4508
rect 4831 4474 4915 4502
rect 4831 4440 4835 4474
rect 4835 4440 4869 4474
rect 4869 4468 4915 4474
rect 4915 4468 4937 4502
rect 4869 4440 4937 4468
rect 4831 4434 4937 4440
rect 4831 4406 4915 4434
rect 4831 4372 4835 4406
rect 4835 4372 4869 4406
rect 4869 4400 4915 4406
rect 4915 4400 4937 4434
rect 4869 4372 4937 4400
rect 4831 4366 4937 4372
rect 4831 4338 4915 4366
rect 4831 4304 4835 4338
rect 4835 4304 4869 4338
rect 4869 4332 4915 4338
rect 4915 4332 4937 4366
rect 4869 4304 4937 4332
rect 4831 4298 4937 4304
rect 4831 4270 4915 4298
rect 4831 4236 4835 4270
rect 4835 4236 4869 4270
rect 4869 4264 4915 4270
rect 4915 4264 4937 4298
rect 4869 4236 4937 4264
rect 4831 4230 4937 4236
rect 4831 4202 4915 4230
rect 4831 4168 4835 4202
rect 4835 4168 4869 4202
rect 4869 4196 4915 4202
rect 4915 4196 4937 4230
rect 4869 4168 4937 4196
rect 4831 4162 4937 4168
rect 4831 4134 4915 4162
rect 4831 4100 4835 4134
rect 4835 4100 4869 4134
rect 4869 4128 4915 4134
rect 4915 4128 4937 4162
rect 4869 4100 4937 4128
rect 4831 4094 4937 4100
rect 4831 4066 4915 4094
rect 4831 4044 4835 4066
rect 4835 4044 4869 4066
rect 4869 4060 4915 4066
rect 4915 4060 4937 4094
rect 4869 4044 4937 4060
rect 4831 3998 4865 4005
rect 4831 3971 4835 3998
rect 4835 3971 4865 3998
rect 4903 3992 4915 4005
rect 4915 3992 4937 4005
rect 4903 3971 4937 3992
rect 4831 3930 4865 3932
rect 4831 3898 4835 3930
rect 4835 3898 4865 3930
rect 4903 3924 4915 3932
rect 4915 3924 4937 3932
rect 4903 3898 4937 3924
rect 4831 3828 4835 3859
rect 4835 3828 4865 3859
rect 4903 3856 4915 3859
rect 4915 3856 4937 3859
rect 4831 3825 4865 3828
rect 4903 3825 4937 3856
rect 323 3752 357 3754
rect 4831 3760 4835 3786
rect 4835 3760 4865 3786
rect 4831 3752 4865 3760
rect 4903 3754 4937 3786
rect 4903 3752 4915 3754
rect 4915 3752 4937 3754
rect 323 3686 357 3713
rect 696 3695 730 3729
rect 781 3695 799 3729
rect 799 3695 815 3729
rect 866 3695 868 3729
rect 868 3695 900 3729
rect 952 3695 971 3729
rect 971 3695 986 3729
rect 1038 3695 1040 3729
rect 1040 3695 1072 3729
rect 1552 3695 1586 3729
rect 1637 3695 1656 3729
rect 1656 3695 1671 3729
rect 1722 3695 1725 3729
rect 1725 3695 1756 3729
rect 1808 3695 1828 3729
rect 1828 3695 1842 3729
rect 1894 3695 1897 3729
rect 1897 3695 1928 3729
rect 2408 3695 2442 3729
rect 2493 3695 2527 3729
rect 2578 3695 2612 3729
rect 2664 3695 2698 3729
rect 2750 3695 2784 3729
rect 3264 3695 3298 3729
rect 3349 3695 3367 3729
rect 3367 3695 3383 3729
rect 3434 3695 3436 3729
rect 3436 3695 3468 3729
rect 3520 3695 3539 3729
rect 3539 3695 3554 3729
rect 3606 3695 3608 3729
rect 3608 3695 3640 3729
rect 4120 3695 4154 3729
rect 4205 3695 4223 3729
rect 4223 3695 4239 3729
rect 4290 3695 4292 3729
rect 4292 3695 4324 3729
rect 4376 3695 4395 3729
rect 4395 3695 4410 3729
rect 4462 3695 4464 3729
rect 4464 3695 4496 3729
rect 323 3679 357 3686
rect 323 3618 357 3640
rect 323 3606 357 3618
rect 323 3533 357 3567
rect 323 3460 357 3494
rect 4831 3692 4835 3713
rect 4835 3692 4865 3713
rect 4831 3679 4865 3692
rect 4903 3686 4937 3713
rect 4903 3679 4915 3686
rect 4915 3679 4937 3686
rect 4831 3624 4835 3640
rect 4835 3624 4865 3640
rect 4831 3606 4865 3624
rect 4903 3618 4937 3640
rect 4903 3606 4915 3618
rect 4915 3606 4937 3618
rect 4831 3556 4835 3567
rect 4835 3556 4865 3567
rect 4831 3533 4865 3556
rect 4903 3533 4937 3567
rect 4831 3488 4835 3494
rect 4835 3488 4865 3494
rect 395 3454 425 3488
rect 425 3454 429 3488
rect 468 3454 493 3488
rect 493 3454 502 3488
rect 541 3454 561 3488
rect 561 3454 575 3488
rect 614 3454 629 3488
rect 629 3454 648 3488
rect 687 3454 697 3488
rect 697 3454 721 3488
rect 760 3454 765 3488
rect 765 3454 794 3488
rect 833 3454 867 3488
rect 906 3454 935 3488
rect 935 3454 940 3488
rect 979 3454 1003 3488
rect 1003 3454 1013 3488
rect 1052 3454 1071 3488
rect 1071 3454 1086 3488
rect 1125 3454 1139 3488
rect 1139 3454 1159 3488
rect 1198 3454 1207 3488
rect 1207 3454 1232 3488
rect 1271 3454 1275 3488
rect 1275 3454 1305 3488
rect 1344 3454 1377 3488
rect 1377 3454 1378 3488
rect 1417 3454 1445 3488
rect 1445 3454 1451 3488
rect 1490 3454 1513 3488
rect 1513 3454 1524 3488
rect 1563 3454 1581 3488
rect 1581 3454 1597 3488
rect 1636 3454 1649 3488
rect 1649 3454 1670 3488
rect 1709 3454 1717 3488
rect 1717 3454 1743 3488
rect 1782 3454 1785 3488
rect 1785 3454 1816 3488
rect 1855 3454 1887 3488
rect 1887 3454 1889 3488
rect 1928 3454 1955 3488
rect 1955 3454 1962 3488
rect 2001 3454 2023 3488
rect 2023 3454 2035 3488
rect 2074 3454 2091 3488
rect 2091 3454 2108 3488
rect 2147 3454 2159 3488
rect 2159 3454 2181 3488
rect 2220 3454 2227 3488
rect 2227 3454 2254 3488
rect 2293 3454 2295 3488
rect 2295 3454 2327 3488
rect 2366 3454 2397 3488
rect 2397 3454 2400 3488
rect 2439 3454 2465 3488
rect 2465 3454 2473 3488
rect 2512 3454 2533 3488
rect 2533 3454 2546 3488
rect 2585 3454 2601 3488
rect 2601 3454 2619 3488
rect 2658 3454 2669 3488
rect 2669 3454 2692 3488
rect 2731 3454 2737 3488
rect 2737 3454 2765 3488
rect 2804 3454 2805 3488
rect 2805 3454 2838 3488
rect 2877 3454 2907 3488
rect 2907 3454 2911 3488
rect 2950 3454 2975 3488
rect 2975 3454 2984 3488
rect 3023 3454 3043 3488
rect 3043 3454 3057 3488
rect 3096 3454 3111 3488
rect 3111 3454 3130 3488
rect 3169 3454 3179 3488
rect 3179 3454 3203 3488
rect 3242 3454 3247 3488
rect 3247 3454 3276 3488
rect 3315 3454 3349 3488
rect 3388 3454 3417 3488
rect 3417 3454 3422 3488
rect 3461 3454 3485 3488
rect 3485 3454 3495 3488
rect 3534 3454 3553 3488
rect 3553 3454 3568 3488
rect 3607 3454 3621 3488
rect 3621 3454 3641 3488
rect 3679 3454 3689 3488
rect 3689 3454 3713 3488
rect 3751 3454 3757 3488
rect 3757 3454 3785 3488
rect 3823 3454 3825 3488
rect 3825 3454 3857 3488
rect 3895 3454 3927 3488
rect 3927 3454 3929 3488
rect 3967 3454 3995 3488
rect 3995 3454 4001 3488
rect 4039 3454 4063 3488
rect 4063 3454 4073 3488
rect 4111 3454 4131 3488
rect 4131 3454 4145 3488
rect 4183 3454 4199 3488
rect 4199 3454 4217 3488
rect 4255 3454 4267 3488
rect 4267 3454 4289 3488
rect 4327 3454 4335 3488
rect 4335 3454 4361 3488
rect 4399 3454 4403 3488
rect 4403 3454 4433 3488
rect 4471 3454 4505 3488
rect 4543 3454 4573 3488
rect 4573 3454 4577 3488
rect 4615 3454 4641 3488
rect 4641 3454 4649 3488
rect 4687 3454 4709 3488
rect 4709 3454 4721 3488
rect 4759 3454 4793 3488
rect 4831 3460 4865 3488
rect 4903 3460 4937 3494
rect 6561 5994 6595 6028
rect 6561 5922 6595 5955
rect 6561 5921 6595 5922
rect 7403 6060 7437 6094
rect 7403 5984 7437 6018
rect 7403 5936 7437 5942
rect 7403 5908 7437 5936
rect 6561 5854 6595 5882
rect 6561 5848 6595 5854
rect 6561 5786 6595 5809
rect 6561 5775 6595 5786
rect 6561 5718 6595 5736
rect 6561 5702 6595 5718
rect 6561 5650 6595 5663
rect 6561 5629 6595 5650
rect 6561 5582 6595 5590
rect 6561 5556 6595 5582
rect 6561 5514 6595 5517
rect 6561 5483 6595 5514
rect 6561 5412 6595 5443
rect 6561 5409 6595 5412
rect 6561 5344 6595 5369
rect 6561 5335 6595 5344
rect 6561 5276 6595 5295
rect 6561 5261 6595 5276
rect 6561 5208 6595 5221
rect 6561 5187 6595 5208
rect 6561 5140 6595 5147
rect 6561 5113 6595 5140
rect 6561 5072 6595 5073
rect 6561 5039 6595 5072
rect 6561 4970 6595 4999
rect 6561 4965 6595 4970
rect 6561 4902 6595 4925
rect 6561 4891 6595 4902
rect 6561 4834 6595 4851
rect 6561 4817 6595 4834
rect 6561 4766 6595 4777
rect 6561 4743 6595 4766
rect 6561 4698 6595 4703
rect 6561 4669 6595 4698
rect 6561 4596 6595 4629
rect 6561 4595 6595 4596
rect 6561 4528 6595 4555
rect 6561 4521 6595 4528
rect 6561 4460 6595 4481
rect 6561 4447 6595 4460
rect 6561 4392 6595 4407
rect 6561 4373 6595 4392
rect 6561 4323 6595 4333
rect 6561 4299 6595 4323
rect 6561 4254 6595 4259
rect 6561 4225 6595 4254
rect 6561 4151 6595 4185
rect 6561 4081 6595 4111
rect 6561 4077 6595 4081
rect 6561 4012 6595 4037
rect 6561 4003 6595 4012
rect 6705 5848 6739 5882
rect 6705 5776 6739 5810
rect 6705 5704 6739 5738
rect 6705 5632 6739 5666
rect 6705 5560 6739 5594
rect 6705 5488 6739 5522
rect 6705 5416 6739 5450
rect 6705 5344 6739 5378
rect 6705 5272 6739 5306
rect 6705 5200 6739 5234
rect 6705 5128 6739 5162
rect 6705 5056 6739 5090
rect 6705 4984 6739 5018
rect 6705 4912 6739 4946
rect 6705 4840 6739 4874
rect 6705 4768 6739 4802
rect 6705 4696 6739 4730
rect 6705 4624 6739 4658
rect 6705 4552 6739 4586
rect 6705 4480 6739 4514
rect 6705 4408 6739 4442
rect 6705 4336 6739 4370
rect 6705 4264 6739 4298
rect 6705 4192 6739 4226
rect 6705 4120 6739 4154
rect 6941 5848 6975 5882
rect 6941 5775 6975 5809
rect 6941 5702 6975 5736
rect 6941 5629 6975 5663
rect 6941 5556 6975 5590
rect 6941 5483 6975 5517
rect 6941 5410 6975 5444
rect 6941 5337 6975 5371
rect 6941 5264 6975 5298
rect 6941 5191 6975 5225
rect 6941 5118 6975 5152
rect 6941 5045 6975 5079
rect 6941 4972 6975 5006
rect 6941 4899 6975 4933
rect 6941 4826 6975 4860
rect 6941 4753 6975 4787
rect 6941 4680 6975 4714
rect 6941 4607 6975 4641
rect 6941 4534 6975 4568
rect 6941 4461 6975 4495
rect 6941 4388 6975 4422
rect 6941 4315 6975 4349
rect 6941 4242 6975 4276
rect 6941 4169 6975 4203
rect 6941 4096 6975 4130
rect 7051 5848 7085 5882
rect 7051 5775 7085 5809
rect 7051 5702 7085 5736
rect 7051 5629 7085 5663
rect 7051 5556 7085 5590
rect 7051 5483 7085 5517
rect 7051 5410 7085 5444
rect 7051 5337 7085 5371
rect 7051 5264 7085 5298
rect 7051 5191 7085 5225
rect 7051 5118 7085 5152
rect 7051 5045 7085 5079
rect 7051 4972 7085 5006
rect 7051 4899 7085 4933
rect 7051 4826 7085 4860
rect 7051 4753 7085 4787
rect 7051 4680 7085 4714
rect 7051 4607 7085 4641
rect 7051 4534 7085 4568
rect 7051 4461 7085 4495
rect 7051 4388 7085 4422
rect 7051 4315 7085 4349
rect 7051 4242 7085 4276
rect 7051 4169 7085 4203
rect 7051 4096 7085 4130
rect 7287 5848 7321 5882
rect 7287 5775 7321 5809
rect 7287 5702 7321 5736
rect 7287 5629 7321 5663
rect 7287 5556 7321 5590
rect 7287 5483 7321 5517
rect 7287 5410 7321 5444
rect 7287 5337 7321 5371
rect 7287 5264 7321 5298
rect 7287 5191 7321 5225
rect 7287 5118 7321 5152
rect 7287 5045 7321 5079
rect 7287 4972 7321 5006
rect 7287 4899 7321 4933
rect 7287 4826 7321 4860
rect 7287 4753 7321 4787
rect 7287 4680 7321 4714
rect 7287 4607 7321 4641
rect 7287 4534 7321 4568
rect 7287 4461 7321 4495
rect 7287 4388 7321 4422
rect 7287 4315 7321 4349
rect 7287 4242 7321 4276
rect 7287 4169 7321 4203
rect 7287 4096 7321 4130
rect 7403 5834 7437 5866
rect 7403 5832 7437 5834
rect 7403 5766 7437 5790
rect 7403 5756 7437 5766
rect 7403 5698 7437 5714
rect 7403 5680 7437 5698
rect 7403 5630 7437 5638
rect 7403 5604 7437 5630
rect 7403 5528 7437 5562
rect 7403 5460 7437 5486
rect 7403 5452 7437 5460
rect 7403 5392 7437 5410
rect 7403 5376 7437 5392
rect 7403 5324 7437 5334
rect 7403 5300 7437 5324
rect 7403 5256 7437 5258
rect 7403 5224 7437 5256
rect 7403 5154 7437 5182
rect 7403 5148 7437 5154
rect 7403 5086 7437 5106
rect 7403 5072 7437 5086
rect 7403 5018 7437 5029
rect 7403 4995 7437 5018
rect 7403 4950 7437 4952
rect 7403 4918 7437 4950
rect 7589 5977 7590 6008
rect 7590 5977 7623 6008
rect 7925 6107 7959 6141
rect 7998 6107 8032 6141
rect 8071 6107 8105 6141
rect 8144 6107 8178 6141
rect 8217 6107 8251 6141
rect 8290 6107 8324 6141
rect 8363 6107 8397 6141
rect 8436 6107 8470 6141
rect 8509 6107 8543 6141
rect 8582 6107 8616 6141
rect 8655 6107 8689 6141
rect 8728 6107 8762 6141
rect 8801 6107 8835 6141
rect 8874 6107 8908 6141
rect 8947 6107 8981 6141
rect 9021 6107 9055 6141
rect 9095 6107 9129 6141
rect 9169 6107 9203 6141
rect 9243 6107 9277 6141
rect 9317 6107 9351 6141
rect 9391 6107 9425 6141
rect 9465 6107 9499 6141
rect 9539 6107 9573 6141
rect 7913 6066 7947 6069
rect 7913 6035 7947 6066
rect 7589 5974 7623 5977
rect 7661 5976 7692 6008
rect 7692 5976 7695 6008
rect 7733 5980 7767 6008
rect 7661 5974 7695 5976
rect 7733 5974 7760 5980
rect 7760 5974 7767 5980
rect 7589 5908 7590 5932
rect 7590 5908 7623 5932
rect 7589 5898 7623 5908
rect 7661 5907 7692 5932
rect 7692 5907 7695 5932
rect 7733 5912 7767 5932
rect 7661 5898 7695 5907
rect 7733 5898 7760 5912
rect 7760 5898 7767 5912
rect 7589 5839 7590 5856
rect 7590 5839 7623 5856
rect 7589 5822 7623 5839
rect 7661 5838 7692 5856
rect 7692 5838 7695 5856
rect 7733 5844 7767 5856
rect 7661 5822 7695 5838
rect 7733 5822 7760 5844
rect 7760 5822 7767 5844
rect 7589 5770 7590 5780
rect 7590 5770 7623 5780
rect 7589 5746 7623 5770
rect 7661 5769 7692 5780
rect 7692 5769 7695 5780
rect 7733 5776 7767 5780
rect 7661 5746 7695 5769
rect 7733 5746 7760 5776
rect 7760 5746 7767 5776
rect 7589 5701 7590 5704
rect 7590 5701 7623 5704
rect 7589 5670 7623 5701
rect 7661 5700 7692 5704
rect 7692 5700 7695 5704
rect 7661 5670 7695 5700
rect 7733 5674 7760 5704
rect 7760 5674 7767 5704
rect 7733 5670 7767 5674
rect 7589 5597 7623 5628
rect 7589 5594 7590 5597
rect 7590 5594 7623 5597
rect 7661 5596 7695 5628
rect 7733 5606 7760 5628
rect 7760 5606 7767 5628
rect 7661 5594 7692 5596
rect 7692 5594 7695 5596
rect 7733 5594 7767 5606
rect 7589 5528 7623 5552
rect 7589 5518 7590 5528
rect 7590 5518 7623 5528
rect 7661 5527 7695 5552
rect 7733 5538 7760 5552
rect 7760 5538 7767 5552
rect 7661 5518 7692 5527
rect 7692 5518 7695 5527
rect 7733 5518 7767 5538
rect 7589 5459 7623 5477
rect 7589 5443 7590 5459
rect 7590 5443 7623 5459
rect 7661 5458 7695 5477
rect 7733 5470 7760 5477
rect 7760 5470 7767 5477
rect 7661 5443 7692 5458
rect 7692 5443 7695 5458
rect 7733 5443 7767 5470
rect 7589 5390 7623 5402
rect 7589 5368 7590 5390
rect 7590 5368 7623 5390
rect 7661 5389 7695 5402
rect 7661 5368 7692 5389
rect 7692 5368 7695 5389
rect 7733 5368 7767 5402
rect 7589 5321 7623 5327
rect 7589 5293 7590 5321
rect 7590 5293 7623 5321
rect 7661 5320 7695 5327
rect 7661 5293 7692 5320
rect 7692 5293 7695 5320
rect 7733 5300 7767 5327
rect 7733 5293 7760 5300
rect 7760 5293 7767 5300
rect 7589 5218 7590 5252
rect 7590 5218 7623 5252
rect 7661 5251 7695 5252
rect 7661 5218 7692 5251
rect 7692 5218 7695 5251
rect 7733 5232 7767 5252
rect 7733 5218 7760 5232
rect 7760 5218 7767 5232
rect 7589 5149 7590 5177
rect 7590 5149 7623 5177
rect 7589 5143 7623 5149
rect 7661 5148 7692 5177
rect 7692 5148 7695 5177
rect 7733 5164 7767 5177
rect 7661 5143 7695 5148
rect 7733 5143 7760 5164
rect 7760 5143 7767 5164
rect 7589 5080 7590 5102
rect 7590 5080 7623 5102
rect 7589 5068 7623 5080
rect 7661 5079 7692 5102
rect 7692 5079 7695 5102
rect 7733 5096 7767 5102
rect 7661 5068 7695 5079
rect 7733 5068 7760 5096
rect 7760 5068 7767 5096
rect 7589 5011 7590 5027
rect 7590 5011 7623 5027
rect 7589 4993 7623 5011
rect 7661 5010 7692 5027
rect 7692 5010 7695 5027
rect 7661 4993 7695 5010
rect 7733 4994 7760 5027
rect 7760 4994 7767 5027
rect 7733 4993 7767 4994
rect 7589 4942 7590 4952
rect 7590 4942 7623 4952
rect 7589 4918 7623 4942
rect 7661 4941 7692 4952
rect 7692 4941 7695 4952
rect 7661 4918 7695 4941
rect 7733 4926 7760 4952
rect 7760 4926 7767 4952
rect 7733 4918 7767 4926
rect 7913 5964 7947 5993
rect 7913 5959 7947 5964
rect 7913 5896 7947 5917
rect 7913 5883 7947 5896
rect 7913 5828 7947 5841
rect 7913 5807 7947 5828
rect 7913 5760 7947 5765
rect 7913 5731 7947 5760
rect 7913 5658 7947 5689
rect 7913 5655 7947 5658
rect 7913 5590 7947 5613
rect 7913 5579 7947 5590
rect 7913 5522 7947 5536
rect 7913 5502 7947 5522
rect 7913 5454 7947 5459
rect 7913 5425 7947 5454
rect 7913 5352 7947 5382
rect 7913 5348 7947 5352
rect 8027 5950 8061 5984
rect 8104 5950 8138 5984
rect 8181 5950 8215 5984
rect 8259 5950 8293 5984
rect 8933 5950 8967 5984
rect 9013 5950 9047 5984
rect 9093 5950 9127 5984
rect 9174 5950 9208 5984
rect 9255 5950 9289 5984
rect 9336 5950 9370 5984
rect 9417 5950 9451 5984
rect 8777 5903 8811 5907
rect 8777 5873 8811 5903
rect 8849 5873 8883 5907
rect 8095 5794 8129 5828
rect 8175 5794 8209 5828
rect 8255 5794 8289 5828
rect 8336 5794 8370 5828
rect 8417 5794 8451 5828
rect 8498 5794 8532 5828
rect 8579 5794 8613 5828
rect 8933 5794 8967 5828
rect 9014 5794 9048 5828
rect 9095 5794 9129 5828
rect 9177 5794 9211 5828
rect 9259 5794 9293 5828
rect 9341 5794 9375 5828
rect 9423 5794 9457 5828
rect 8027 5638 8061 5672
rect 8107 5638 8141 5672
rect 8187 5638 8221 5672
rect 8268 5638 8302 5672
rect 8349 5638 8383 5672
rect 8864 5638 8898 5672
rect 8943 5638 8977 5672
rect 9023 5638 9057 5672
rect 9103 5638 9137 5672
rect 9183 5638 9217 5672
rect 9263 5638 9297 5672
rect 9343 5638 9377 5672
rect 9423 5638 9457 5672
rect 8095 5482 8129 5516
rect 8175 5482 8209 5516
rect 8255 5482 8289 5516
rect 8336 5482 8370 5516
rect 8417 5482 8451 5516
rect 8498 5482 8532 5516
rect 8579 5482 8613 5516
rect 8867 5528 8901 5562
rect 8946 5528 8980 5562
rect 9025 5528 9059 5562
rect 9104 5528 9138 5562
rect 9183 5528 9217 5562
rect 9263 5528 9297 5562
rect 9343 5528 9377 5562
rect 9423 5528 9457 5562
rect 8681 5450 8715 5484
rect 8753 5481 8777 5484
rect 8777 5481 8787 5484
rect 8753 5450 8787 5481
rect 8027 5326 8061 5360
rect 8105 5326 8139 5360
rect 8184 5326 8218 5360
rect 8263 5326 8297 5360
rect 8342 5326 8376 5360
rect 8421 5326 8455 5360
rect 8500 5326 8534 5360
rect 8579 5326 8613 5360
rect 8862 5352 8896 5386
rect 8937 5352 8971 5386
rect 9012 5352 9046 5386
rect 9087 5352 9121 5386
rect 9162 5352 9196 5386
rect 9237 5352 9271 5386
rect 9312 5352 9346 5386
rect 9387 5352 9421 5386
rect 9463 5352 9497 5386
rect 9539 5359 9551 5386
rect 9551 5359 9573 5386
rect 9539 5352 9573 5359
rect 7913 5284 7947 5305
rect 7913 5271 7947 5284
rect 7913 5216 7947 5228
rect 8029 5216 8063 5250
rect 8104 5216 8138 5250
rect 8179 5216 8213 5250
rect 8254 5216 8288 5250
rect 8330 5216 8364 5250
rect 8406 5216 8440 5250
rect 8482 5216 8516 5250
rect 9764 5982 9870 6088
rect 10510 6378 10544 6412
rect 10584 6378 10617 6412
rect 10617 6378 10618 6412
rect 10658 6378 10685 6412
rect 10685 6378 10692 6412
rect 10732 6378 10753 6412
rect 10753 6378 10766 6412
rect 10806 6378 10821 6412
rect 10821 6378 10840 6412
rect 10880 6378 10889 6412
rect 10889 6378 10914 6412
rect 10954 6378 10957 6412
rect 10957 6378 10988 6412
rect 11028 6378 11059 6412
rect 11059 6378 11062 6412
rect 11102 6378 11127 6412
rect 11127 6378 11136 6412
rect 11176 6378 11195 6412
rect 11195 6378 11210 6412
rect 11250 6378 11263 6412
rect 11263 6378 11284 6412
rect 11324 6378 11331 6412
rect 11331 6378 11358 6412
rect 11398 6378 11399 6412
rect 11399 6378 11432 6412
rect 11472 6378 11480 6412
rect 11480 6378 11506 6412
rect 11546 6378 11548 6412
rect 11548 6378 11580 6412
rect 11620 6378 11650 6412
rect 11650 6378 11654 6412
rect 11694 6378 11718 6412
rect 11718 6378 11728 6412
rect 11768 6378 11786 6412
rect 11786 6378 11802 6412
rect 11842 6378 11854 6412
rect 11854 6378 11876 6412
rect 11916 6378 11922 6412
rect 11922 6378 11950 6412
rect 11990 6378 12024 6412
rect 12064 6378 12092 6412
rect 12092 6378 12098 6412
rect 12138 6378 12160 6412
rect 12160 6378 12172 6412
rect 12212 6378 12228 6412
rect 12228 6378 12246 6412
rect 12286 6378 12296 6412
rect 12296 6378 12320 6412
rect 12360 6378 12364 6412
rect 12364 6378 12394 6412
rect 12434 6378 12466 6412
rect 12466 6378 12468 6412
rect 12508 6378 12534 6412
rect 12534 6378 12542 6412
rect 12581 6378 12602 6412
rect 12602 6378 12615 6412
rect 12654 6378 12670 6412
rect 12670 6378 12688 6412
rect 12727 6378 12738 6412
rect 12738 6378 12761 6412
rect 12800 6378 12806 6412
rect 12806 6378 12834 6412
rect 12873 6378 12874 6412
rect 12874 6378 12907 6412
rect 12946 6378 12976 6412
rect 12976 6378 12980 6412
rect 13019 6378 13044 6412
rect 13044 6378 13053 6412
rect 13092 6378 13112 6412
rect 13112 6378 13126 6412
rect 13165 6378 13199 6412
rect 13238 6378 13258 6412
rect 13258 6378 13272 6412
rect 13311 6378 13326 6412
rect 13326 6378 13345 6412
rect 13384 6378 13394 6412
rect 13394 6378 13418 6412
rect 13496 6340 13530 6374
rect 10707 6243 10709 6277
rect 10709 6243 10741 6277
rect 10779 6243 10811 6277
rect 10811 6243 10813 6277
rect 11046 6232 11152 6338
rect 13496 6294 13530 6300
rect 13100 6277 13134 6280
rect 13172 6277 13206 6280
rect 11979 6243 12013 6277
rect 12051 6243 12085 6277
rect 12580 6243 12584 6277
rect 12584 6243 12614 6277
rect 12652 6243 12686 6277
rect 11290 6158 11324 6192
rect 11362 6158 11396 6192
rect 10870 6062 10904 6096
rect 10870 5990 10904 6024
rect 10870 5918 10904 5952
rect 11222 6062 11256 6096
rect 11222 5990 11256 6024
rect 11222 5918 11256 5952
rect 10614 5692 10720 5798
rect 11406 5714 11512 5820
rect 11588 5758 11622 5792
rect 11588 5686 11622 5720
rect 11940 5758 11974 5792
rect 11764 5684 11798 5718
rect 11940 5686 11974 5720
rect 11764 5612 11798 5646
rect 12897 6171 13003 6277
rect 13100 6246 13130 6277
rect 13130 6246 13134 6277
rect 13172 6246 13198 6277
rect 13198 6246 13206 6277
rect 13496 6266 13530 6294
rect 13496 6192 13530 6226
rect 13496 6124 13530 6152
rect 13496 6118 13530 6124
rect 13496 6056 13530 6078
rect 12713 6021 12747 6055
rect 12713 5949 12747 5983
rect 12713 5877 12747 5911
rect 12713 5805 12747 5839
rect 12292 5758 12326 5792
rect 12116 5684 12150 5718
rect 12292 5686 12326 5720
rect 12378 5758 12412 5792
rect 12713 5733 12747 5767
rect 13225 6021 13259 6055
rect 13225 5949 13259 5983
rect 13225 5877 13259 5911
rect 13225 5805 13259 5839
rect 13225 5733 13259 5767
rect 13496 6044 13530 6056
rect 13496 5988 13530 6005
rect 13496 5971 13530 5988
rect 13496 5920 13530 5932
rect 13496 5898 13530 5920
rect 13496 5852 13530 5859
rect 13496 5825 13530 5852
rect 13496 5784 13530 5786
rect 13496 5752 13530 5784
rect 12378 5686 12412 5720
rect 12116 5612 12150 5646
rect 13496 5682 13530 5713
rect 13496 5679 13530 5682
rect 13496 5606 13530 5640
rect 13496 5563 13530 5567
rect 13496 5533 13530 5563
rect 12381 5477 12385 5478
rect 12385 5477 12415 5478
rect 12453 5477 12487 5478
rect 12381 5444 12415 5477
rect 12453 5444 12487 5477
rect 13496 5461 13530 5494
rect 13496 5460 13530 5461
rect 9551 5223 9585 5226
rect 7913 5194 7947 5216
rect 8600 5176 8634 5210
rect 8672 5189 8706 5210
rect 8672 5176 8703 5189
rect 8703 5176 8706 5189
rect 8893 5176 8927 5210
rect 8974 5176 9008 5210
rect 9055 5176 9089 5210
rect 9136 5176 9170 5210
rect 9217 5176 9251 5210
rect 9297 5176 9331 5210
rect 9377 5176 9411 5210
rect 9551 5192 9585 5223
rect 7913 5148 7947 5151
rect 7913 5117 7947 5148
rect 7913 5046 7947 5074
rect 9551 5121 9585 5150
rect 9551 5116 9585 5121
rect 8862 5066 8896 5100
rect 8941 5066 8975 5100
rect 9021 5066 9055 5100
rect 9101 5066 9135 5100
rect 9181 5066 9215 5100
rect 9261 5066 9295 5100
rect 9341 5066 9375 5100
rect 9421 5066 9455 5100
rect 7913 5040 7947 5046
rect 7913 4978 7947 4997
rect 9551 5053 9585 5073
rect 9551 5039 9585 5053
rect 7913 4963 7947 4978
rect 8029 4960 8063 4994
rect 8111 4960 8145 4994
rect 8192 4960 8226 4994
rect 8273 4960 8307 4994
rect 8354 4960 8388 4994
rect 8435 4960 8469 4994
rect 9551 4985 9585 4996
rect 9551 4962 9585 4985
rect 7403 4678 7437 4708
rect 7403 4674 7437 4678
rect 7403 4610 7437 4636
rect 8585 4887 8619 4921
rect 8657 4899 8669 4921
rect 8669 4899 8691 4921
rect 8657 4887 8691 4899
rect 8867 4890 8901 4924
rect 8942 4890 8976 4924
rect 9017 4890 9051 4924
rect 9092 4890 9126 4924
rect 9167 4890 9201 4924
rect 9242 4890 9276 4924
rect 9317 4890 9351 4924
rect 9391 4890 9425 4924
rect 9465 4890 9499 4924
rect 9539 4917 9573 4924
rect 9539 4890 9551 4917
rect 9551 4890 9573 4917
rect 9734 5192 9738 5226
rect 9738 5192 9768 5226
rect 9806 5192 9840 5226
rect 9878 5192 9908 5226
rect 9908 5192 9912 5226
rect 9734 5117 9738 5151
rect 9738 5117 9768 5151
rect 9806 5117 9840 5151
rect 9878 5117 9908 5151
rect 9908 5117 9912 5151
rect 9734 5042 9738 5076
rect 9738 5042 9768 5076
rect 9806 5042 9840 5076
rect 9878 5042 9908 5076
rect 9908 5042 9912 5076
rect 9734 4967 9738 5001
rect 9738 4967 9768 5001
rect 9806 4967 9840 5001
rect 9878 4967 9908 5001
rect 9908 4967 9912 5001
rect 9734 4893 9738 4927
rect 9738 4893 9768 4927
rect 9806 4893 9840 4927
rect 9878 4893 9908 4927
rect 9908 4893 9912 4927
rect 10770 5336 10804 5370
rect 10770 5253 10804 5287
rect 8029 4784 8063 4818
rect 8111 4784 8145 4818
rect 8192 4784 8226 4818
rect 8273 4784 8307 4818
rect 8354 4784 8388 4818
rect 8435 4784 8469 4818
rect 8715 4714 8749 4748
rect 8787 4714 8821 4748
rect 8918 4714 8952 4748
rect 8991 4714 9025 4748
rect 9063 4714 9097 4748
rect 9135 4714 9169 4748
rect 9207 4714 9241 4748
rect 9279 4714 9313 4748
rect 9351 4714 9385 4748
rect 10614 5178 10648 5212
rect 10614 5095 10648 5129
rect 10614 5011 10648 5045
rect 11082 5336 11116 5370
rect 11082 5253 11116 5287
rect 10770 5169 10804 5203
rect 10770 5085 10804 5119
rect 10770 5001 10804 5035
rect 10926 5178 10960 5212
rect 10926 5095 10960 5129
rect 10926 5011 10960 5045
rect 10614 4927 10648 4961
rect 10614 4843 10648 4877
rect 11394 5336 11428 5370
rect 11394 5253 11428 5287
rect 11082 5169 11116 5203
rect 11082 5085 11116 5119
rect 11082 5001 11116 5035
rect 11238 5178 11272 5212
rect 11238 5095 11272 5129
rect 11238 5011 11272 5045
rect 10926 4927 10960 4961
rect 10926 4843 10960 4877
rect 11706 5336 11740 5370
rect 11706 5253 11740 5287
rect 11394 5169 11428 5203
rect 11394 5085 11428 5119
rect 11394 5001 11428 5035
rect 11550 5178 11584 5212
rect 11550 5095 11584 5129
rect 11550 5011 11584 5045
rect 11238 4927 11272 4961
rect 11238 4843 11272 4877
rect 11706 5169 11740 5203
rect 11706 5085 11740 5119
rect 11706 5001 11740 5035
rect 11862 5336 11896 5370
rect 12500 5362 12534 5396
rect 11862 5254 11896 5288
rect 11862 5172 11896 5206
rect 11862 5090 11896 5124
rect 11862 5008 11896 5042
rect 11550 4927 11584 4961
rect 11550 4843 11584 4877
rect 11862 4926 11896 4960
rect 11862 4843 11896 4877
rect 11972 5321 12006 5355
rect 11972 5241 12006 5275
rect 11972 5161 12006 5195
rect 11972 5080 12006 5114
rect 11972 4999 12006 5033
rect 11972 4918 12006 4952
rect 11972 4837 12006 4871
rect 12324 5321 12358 5355
rect 12324 5242 12358 5276
rect 12324 5163 12358 5197
rect 12324 5083 12358 5117
rect 12324 5003 12358 5037
rect 12852 5392 12886 5426
rect 12500 5290 12534 5324
rect 12500 5218 12534 5252
rect 12500 5146 12534 5180
rect 12500 5074 12534 5108
rect 12500 5001 12534 5035
rect 12676 5321 12710 5355
rect 12676 5242 12710 5276
rect 12676 5163 12710 5197
rect 12676 5083 12710 5117
rect 12676 5003 12710 5037
rect 12324 4923 12358 4957
rect 12324 4843 12358 4877
rect 13205 5392 13239 5426
rect 12852 5314 12886 5348
rect 12852 5236 12886 5270
rect 12852 5158 12886 5192
rect 12852 5080 12886 5114
rect 12852 5001 12886 5035
rect 13028 5321 13062 5355
rect 13028 5242 13062 5276
rect 13028 5163 13062 5197
rect 13028 5083 13062 5117
rect 13028 5003 13062 5037
rect 12676 4923 12710 4957
rect 12676 4843 12710 4877
rect 13496 5393 13530 5421
rect 13496 5387 13530 5393
rect 13205 5314 13239 5348
rect 13205 5236 13239 5270
rect 13205 5158 13239 5192
rect 13205 5080 13239 5114
rect 13205 5001 13239 5035
rect 13380 5321 13414 5355
rect 13380 5242 13414 5276
rect 13380 5163 13414 5197
rect 13380 5083 13414 5117
rect 13380 5003 13414 5037
rect 13028 4923 13062 4957
rect 13028 4843 13062 4877
rect 13380 4923 13414 4957
rect 13380 4843 13414 4877
rect 13496 5325 13530 5348
rect 13496 5314 13530 5325
rect 13496 5257 13530 5275
rect 13496 5241 13530 5257
rect 13496 5189 13530 5202
rect 13496 5168 13530 5189
rect 13496 5121 13530 5129
rect 13496 5095 13530 5121
rect 13496 5053 13530 5056
rect 13496 5022 13530 5053
rect 13496 4951 13530 4983
rect 13496 4949 13530 4951
rect 13496 4883 13530 4910
rect 13496 4876 13530 4883
rect 13496 4815 13530 4837
rect 13496 4803 13530 4815
rect 7913 4706 7947 4708
rect 7913 4674 7947 4706
rect 9551 4713 9585 4745
rect 9551 4711 9585 4713
rect 9551 4645 9585 4658
rect 7403 4602 7437 4610
rect 7403 4542 7437 4564
rect 7403 4530 7437 4542
rect 7403 4474 7437 4492
rect 7403 4458 7437 4474
rect 7403 4406 7437 4420
rect 7403 4386 7437 4406
rect 7403 4338 7437 4348
rect 7403 4314 7437 4338
rect 7403 4270 7437 4276
rect 7403 4242 7437 4270
rect 7403 4202 7437 4203
rect 7403 4169 7437 4202
rect 7403 4100 7437 4130
rect 7403 4096 7437 4100
rect 7589 4631 7767 4634
rect 7589 4597 7590 4631
rect 7590 4597 7624 4631
rect 7624 4630 7767 4631
rect 7624 4597 7658 4630
rect 7589 4596 7658 4597
rect 7658 4596 7692 4630
rect 7692 4620 7767 4630
rect 7692 4596 7726 4620
rect 7589 4586 7726 4596
rect 7726 4586 7760 4620
rect 7760 4586 7767 4620
rect 7589 4562 7767 4586
rect 7589 4528 7590 4562
rect 7590 4528 7624 4562
rect 7624 4561 7767 4562
rect 7624 4528 7658 4561
rect 7589 4527 7658 4528
rect 7658 4527 7692 4561
rect 7692 4552 7767 4561
rect 7692 4527 7726 4552
rect 7589 4518 7726 4527
rect 7726 4518 7760 4552
rect 7760 4518 7767 4552
rect 7589 4493 7767 4518
rect 7589 4459 7590 4493
rect 7590 4459 7624 4493
rect 7624 4492 7767 4493
rect 7624 4459 7658 4492
rect 7589 4458 7658 4459
rect 7658 4458 7692 4492
rect 7692 4484 7767 4492
rect 7692 4458 7726 4484
rect 7589 4450 7726 4458
rect 7726 4450 7760 4484
rect 7760 4450 7767 4484
rect 7589 4424 7767 4450
rect 7589 4390 7590 4424
rect 7590 4390 7624 4424
rect 7624 4423 7767 4424
rect 7624 4390 7658 4423
rect 7589 4389 7658 4390
rect 7658 4389 7692 4423
rect 7692 4416 7767 4423
rect 7692 4389 7726 4416
rect 7589 4382 7726 4389
rect 7726 4382 7760 4416
rect 7760 4382 7767 4416
rect 7589 4355 7767 4382
rect 7589 4321 7590 4355
rect 7590 4321 7624 4355
rect 7624 4354 7767 4355
rect 7624 4321 7658 4354
rect 7589 4320 7658 4321
rect 7658 4320 7692 4354
rect 7692 4348 7767 4354
rect 7692 4320 7726 4348
rect 7589 4314 7726 4320
rect 7726 4314 7760 4348
rect 7760 4314 7767 4348
rect 7589 4286 7767 4314
rect 7589 4252 7590 4286
rect 7590 4252 7624 4286
rect 7624 4285 7767 4286
rect 7624 4252 7658 4285
rect 7589 4251 7658 4252
rect 7658 4251 7692 4285
rect 7692 4280 7767 4285
rect 7692 4251 7726 4280
rect 7589 4246 7726 4251
rect 7726 4246 7760 4280
rect 7760 4246 7767 4280
rect 7589 4217 7767 4246
rect 7589 4183 7590 4217
rect 7590 4183 7624 4217
rect 7624 4216 7767 4217
rect 7624 4183 7658 4216
rect 7589 4182 7658 4183
rect 7658 4182 7692 4216
rect 7692 4212 7767 4216
rect 7692 4182 7726 4212
rect 7589 4178 7726 4182
rect 7726 4178 7760 4212
rect 7760 4178 7767 4212
rect 7589 4148 7767 4178
rect 7589 4114 7590 4148
rect 7590 4114 7624 4148
rect 7624 4147 7767 4148
rect 7624 4114 7658 4147
rect 7589 4113 7658 4114
rect 7658 4113 7692 4147
rect 7692 4144 7767 4147
rect 7692 4113 7726 4144
rect 7589 4110 7726 4113
rect 7726 4110 7760 4144
rect 7760 4110 7767 4144
rect 7589 4096 7767 4110
rect 7913 4604 7947 4636
rect 8029 4608 8063 4642
rect 8110 4608 8144 4642
rect 8191 4608 8225 4642
rect 8272 4608 8306 4642
rect 8353 4608 8387 4642
rect 8433 4608 8467 4642
rect 8513 4608 8547 4642
rect 9551 4624 9585 4645
rect 7913 4602 7947 4604
rect 7913 4536 7947 4564
rect 7913 4530 7947 4536
rect 7913 4468 7947 4492
rect 7913 4458 7947 4468
rect 7913 4400 7947 4420
rect 7913 4386 7947 4400
rect 8867 4538 8901 4572
rect 8948 4538 8982 4572
rect 9029 4538 9063 4572
rect 9110 4538 9144 4572
rect 9191 4538 9225 4572
rect 9271 4538 9305 4572
rect 9351 4538 9385 4572
rect 9551 4543 9585 4571
rect 8674 4479 8703 4485
rect 8703 4479 8708 4485
rect 8674 4451 8708 4479
rect 8674 4411 8703 4413
rect 8703 4411 8708 4413
rect 8029 4352 8063 4386
rect 8104 4352 8138 4386
rect 8179 4352 8213 4386
rect 8254 4352 8288 4386
rect 8328 4352 8362 4386
rect 8402 4352 8436 4386
rect 8476 4352 8510 4386
rect 8550 4352 8584 4386
rect 8674 4379 8708 4411
rect 9551 4537 9585 4543
rect 9734 4711 9738 4745
rect 9738 4711 9768 4745
rect 9806 4711 9840 4745
rect 9878 4711 9908 4745
rect 9908 4711 9912 4745
rect 9734 4624 9738 4658
rect 9738 4624 9768 4658
rect 9806 4624 9840 4658
rect 9878 4624 9908 4658
rect 9908 4624 9912 4658
rect 9734 4537 9738 4571
rect 9738 4537 9768 4571
rect 9806 4537 9840 4571
rect 9878 4537 9908 4571
rect 9908 4537 9912 4571
rect 13496 4747 13530 4764
rect 13496 4730 13530 4747
rect 8867 4382 8901 4416
rect 8948 4382 8982 4416
rect 9029 4382 9063 4416
rect 9110 4382 9144 4416
rect 9191 4382 9225 4416
rect 9271 4382 9305 4416
rect 9351 4382 9385 4416
rect 7913 4332 7947 4348
rect 7913 4314 7947 4332
rect 7913 4264 7947 4276
rect 7913 4242 7947 4264
rect 8029 4242 8063 4276
rect 8104 4242 8138 4276
rect 8179 4242 8213 4276
rect 8254 4242 8288 4276
rect 8328 4242 8362 4276
rect 8402 4242 8436 4276
rect 8476 4242 8510 4276
rect 8550 4242 8584 4276
rect 8867 4272 8901 4306
rect 8948 4272 8982 4306
rect 9029 4272 9063 4306
rect 9110 4272 9144 4306
rect 9191 4272 9225 4306
rect 9271 4272 9305 4306
rect 9351 4272 9385 4306
rect 7913 4196 7947 4203
rect 7913 4169 7947 4196
rect 7913 4128 7947 4130
rect 7913 4096 7947 4128
rect 6705 4048 6739 4082
rect 6705 3976 6739 4010
rect 6561 3943 6595 3963
rect 6561 3929 6595 3943
rect 6561 3874 6595 3889
rect 6561 3855 6595 3874
rect 7403 3896 7437 3924
rect 7403 3890 7437 3896
rect 8597 4093 8631 4127
rect 8669 4110 8703 4127
rect 8669 4093 8703 4110
rect 8918 4096 8952 4130
rect 8991 4096 9025 4130
rect 9063 4096 9097 4130
rect 9135 4096 9169 4130
rect 9207 4096 9241 4130
rect 9279 4096 9313 4130
rect 9351 4096 9385 4130
rect 9734 4377 9738 4411
rect 9738 4377 9768 4411
rect 9806 4377 9840 4411
rect 9878 4377 9908 4411
rect 9908 4377 9912 4411
rect 9734 4283 9738 4317
rect 9738 4283 9768 4317
rect 9806 4283 9840 4317
rect 9878 4283 9908 4317
rect 9908 4283 9912 4317
rect 9734 4189 9738 4223
rect 9738 4189 9768 4223
rect 9806 4189 9840 4223
rect 9878 4189 9908 4223
rect 9908 4189 9912 4223
rect 9734 4096 9738 4130
rect 9738 4096 9768 4130
rect 9806 4096 9840 4130
rect 9878 4096 9908 4130
rect 9908 4096 9912 4130
rect 10614 4671 10648 4705
rect 10614 4599 10648 4633
rect 10614 4526 10648 4560
rect 10926 4671 10960 4705
rect 10926 4599 10960 4633
rect 10614 4453 10648 4487
rect 10614 4380 10648 4414
rect 10614 4307 10648 4341
rect 10770 4513 10804 4547
rect 10770 4441 10804 4475
rect 10770 4368 10804 4402
rect 10770 4295 10804 4329
rect 10926 4526 10960 4560
rect 11238 4671 11272 4705
rect 11238 4599 11272 4633
rect 10926 4453 10960 4487
rect 10926 4380 10960 4414
rect 10926 4307 10960 4341
rect 11082 4513 11116 4547
rect 11082 4441 11116 4475
rect 11082 4368 11116 4402
rect 10770 4222 10804 4256
rect 10770 4149 10804 4183
rect 11082 4295 11116 4329
rect 11238 4526 11272 4560
rect 11550 4671 11584 4705
rect 11550 4599 11584 4633
rect 11238 4453 11272 4487
rect 11238 4380 11272 4414
rect 11238 4307 11272 4341
rect 11394 4513 11428 4547
rect 11394 4441 11428 4475
rect 11394 4368 11428 4402
rect 11082 4222 11116 4256
rect 11082 4149 11116 4183
rect 11394 4295 11428 4329
rect 11550 4526 11584 4560
rect 11862 4671 11896 4705
rect 11862 4599 11896 4633
rect 11550 4453 11584 4487
rect 11550 4380 11584 4414
rect 11550 4307 11584 4341
rect 11706 4513 11740 4547
rect 11706 4441 11740 4475
rect 11706 4368 11740 4402
rect 11394 4222 11428 4256
rect 11394 4149 11428 4183
rect 11706 4295 11740 4329
rect 11862 4526 11896 4560
rect 12174 4671 12208 4705
rect 12174 4599 12208 4633
rect 11862 4453 11896 4487
rect 11862 4380 11896 4414
rect 11862 4307 11896 4341
rect 12018 4513 12052 4547
rect 12018 4441 12052 4475
rect 12018 4368 12052 4402
rect 11706 4222 11740 4256
rect 11706 4149 11740 4183
rect 12018 4295 12052 4329
rect 12174 4526 12208 4560
rect 12486 4671 12520 4705
rect 12486 4599 12520 4633
rect 12174 4453 12208 4487
rect 12174 4380 12208 4414
rect 12174 4307 12208 4341
rect 12330 4513 12364 4547
rect 12330 4441 12364 4475
rect 12330 4368 12364 4402
rect 12018 4222 12052 4256
rect 12018 4149 12052 4183
rect 12330 4295 12364 4329
rect 12486 4526 12520 4560
rect 12798 4671 12832 4705
rect 12798 4599 12832 4633
rect 12486 4453 12520 4487
rect 12486 4380 12520 4414
rect 12486 4307 12520 4341
rect 12642 4513 12676 4547
rect 12642 4441 12676 4475
rect 12642 4368 12676 4402
rect 12330 4222 12364 4256
rect 12330 4149 12364 4183
rect 12642 4295 12676 4329
rect 12798 4526 12832 4560
rect 13110 4671 13144 4705
rect 13110 4597 13144 4631
rect 12798 4453 12832 4487
rect 12798 4380 12832 4414
rect 12798 4307 12832 4341
rect 12954 4513 12988 4547
rect 12954 4441 12988 4475
rect 12954 4368 12988 4402
rect 12642 4222 12676 4256
rect 12642 4149 12676 4183
rect 12954 4295 12988 4329
rect 12954 4222 12988 4256
rect 12954 4149 12988 4183
rect 13110 4523 13144 4557
rect 13110 4449 13144 4483
rect 13110 4374 13144 4408
rect 13110 4299 13144 4333
rect 13110 4224 13144 4258
rect 13110 4149 13144 4183
rect 13496 4679 13530 4691
rect 13496 4657 13530 4679
rect 13496 4611 13530 4618
rect 13496 4584 13530 4611
rect 13496 4543 13530 4545
rect 13496 4511 13530 4543
rect 13496 4441 13530 4472
rect 13496 4438 13530 4441
rect 13496 4373 13530 4399
rect 13496 4365 13530 4373
rect 13496 4305 13530 4326
rect 13496 4292 13530 4305
rect 13496 4237 13530 4253
rect 13496 4219 13530 4237
rect 13496 4169 13530 4180
rect 7913 3890 7947 3924
rect 8029 3890 8063 3924
rect 8104 3890 8138 3924
rect 8179 3890 8213 3924
rect 8254 3890 8288 3924
rect 8328 3890 8362 3924
rect 8402 3890 8436 3924
rect 8476 3890 8510 3924
rect 8550 3890 8584 3924
rect 8669 3890 8703 3924
rect 8741 3890 8775 3924
rect 8867 3920 8901 3954
rect 8948 3920 8982 3954
rect 9029 3920 9063 3954
rect 9110 3920 9144 3954
rect 9191 3920 9225 3954
rect 9271 3920 9305 3954
rect 9351 3920 9385 3954
rect 13496 4146 13530 4169
rect 13496 4101 13530 4107
rect 13496 4073 13530 4101
rect 10663 4037 10697 4071
rect 10735 4037 10769 4071
rect 10807 4037 10841 4071
rect 10879 4037 10913 4071
rect 10951 4037 10985 4071
rect 11023 4037 11057 4071
rect 11095 4037 11129 4071
rect 11167 4037 11201 4071
rect 11239 4037 11273 4071
rect 11311 4037 11345 4071
rect 11383 4037 11417 4071
rect 11455 4037 11489 4071
rect 11527 4037 11561 4071
rect 11599 4037 11633 4071
rect 11672 4037 11706 4071
rect 11745 4037 11779 4071
rect 11818 4037 11852 4071
rect 11891 4037 11925 4071
rect 11964 4037 11998 4071
rect 12037 4037 12071 4071
rect 12110 4037 12144 4071
rect 12183 4037 12217 4071
rect 12256 4037 12290 4071
rect 12329 4037 12363 4071
rect 12402 4037 12436 4071
rect 12475 4037 12509 4071
rect 12548 4037 12582 4071
rect 12621 4037 12655 4071
rect 12694 4037 12728 4071
rect 12767 4037 12801 4071
rect 12840 4037 12874 4071
rect 12913 4037 12947 4071
rect 12986 4037 13020 4071
rect 13059 4037 13093 4071
rect 10510 3965 10532 3995
rect 10532 3965 10544 3995
rect 10583 3965 10600 3995
rect 10600 3965 10617 3995
rect 10656 3965 10668 3995
rect 10668 3965 10690 3995
rect 10729 3965 10736 3995
rect 10736 3965 10763 3995
rect 10802 3965 10804 3995
rect 10804 3965 10836 3995
rect 10875 3965 10906 3995
rect 10906 3965 10909 3995
rect 10948 3965 10974 3995
rect 10974 3965 10982 3995
rect 11021 3965 11042 3995
rect 11042 3965 11055 3995
rect 11094 3965 11110 3995
rect 11110 3965 11128 3995
rect 11167 3965 11178 3995
rect 11178 3965 11201 3995
rect 11240 3965 11246 3995
rect 11246 3965 11274 3995
rect 11313 3965 11314 3995
rect 11314 3965 11347 3995
rect 11386 3965 11416 3995
rect 11416 3965 11420 3995
rect 11460 3965 11484 3995
rect 11484 3965 11494 3995
rect 11534 3965 11552 3995
rect 11552 3965 11568 3995
rect 11608 3965 11620 3995
rect 11620 3965 11642 3995
rect 11682 3965 11688 3995
rect 11688 3965 11716 3995
rect 11756 3965 11790 3995
rect 11830 3965 11858 3995
rect 11858 3965 11864 3995
rect 11904 3965 11926 3995
rect 11926 3965 11938 3995
rect 11978 3965 11994 3995
rect 11994 3965 12012 3995
rect 12052 3965 12062 3995
rect 12062 3965 12086 3995
rect 12126 3965 12130 3995
rect 12130 3965 12160 3995
rect 12200 3965 12232 3995
rect 12232 3965 12234 3995
rect 12274 3965 12300 3995
rect 12300 3965 12308 3995
rect 12348 3965 12368 3995
rect 12368 3965 12382 3995
rect 12422 3965 12436 3995
rect 12436 3965 12456 3995
rect 12496 3965 12504 3995
rect 12504 3965 12530 3995
rect 12570 3965 12572 3995
rect 12572 3965 12604 3995
rect 12644 3965 12674 3995
rect 12674 3965 12678 3995
rect 12718 3965 12742 3995
rect 12742 3965 12752 3995
rect 12792 3965 12810 3995
rect 12810 3965 12826 3995
rect 12866 3965 12878 3995
rect 12878 3965 12900 3995
rect 12940 3965 12946 3995
rect 12946 3965 12974 3995
rect 10510 3961 10544 3965
rect 10583 3961 10617 3965
rect 10656 3961 10690 3965
rect 10729 3961 10763 3965
rect 10802 3961 10836 3965
rect 10875 3961 10909 3965
rect 10948 3961 10982 3965
rect 11021 3961 11055 3965
rect 11094 3961 11128 3965
rect 11167 3961 11201 3965
rect 11240 3961 11274 3965
rect 11313 3961 11347 3965
rect 11386 3961 11420 3965
rect 11460 3961 11494 3965
rect 11534 3961 11568 3965
rect 11608 3961 11642 3965
rect 11682 3961 11716 3965
rect 11756 3961 11790 3965
rect 11830 3961 11864 3965
rect 11904 3961 11938 3965
rect 11978 3961 12012 3965
rect 12052 3961 12086 3965
rect 12126 3961 12160 3965
rect 12200 3961 12234 3965
rect 12274 3961 12308 3965
rect 12348 3961 12382 3965
rect 12422 3961 12456 3965
rect 12496 3961 12530 3965
rect 12570 3961 12604 3965
rect 12644 3961 12678 3965
rect 12718 3961 12752 3965
rect 12792 3961 12826 3965
rect 12866 3961 12900 3965
rect 12940 3961 12974 3965
rect 13014 3961 13048 3995
rect 13088 3965 13116 3995
rect 13116 3965 13122 3995
rect 13162 3965 13184 3995
rect 13184 3965 13196 3995
rect 13236 3965 13252 3995
rect 13252 3965 13270 3995
rect 13310 3965 13320 3995
rect 13320 3965 13344 3995
rect 13384 3965 13388 3995
rect 13388 3965 13418 3995
rect 13088 3961 13122 3965
rect 13162 3961 13196 3965
rect 13236 3961 13270 3965
rect 13310 3961 13344 3965
rect 13384 3961 13418 3965
rect 13458 3961 13492 3995
rect 6561 3805 6595 3815
rect 6561 3781 6595 3805
rect 6780 3786 6814 3820
rect 6852 3786 6886 3820
rect 6924 3786 6958 3820
rect 6996 3786 7030 3820
rect 7068 3786 7102 3820
rect 7140 3786 7174 3820
rect 7212 3786 7246 3820
rect 7403 3794 7437 3815
rect 7403 3781 7437 3794
rect 7589 3816 7590 3850
rect 7590 3816 7623 3850
rect 7661 3816 7695 3850
rect 7733 3816 7760 3850
rect 7760 3816 7767 3850
rect 4987 3454 5017 3488
rect 5017 3454 5021 3488
rect 5061 3454 5085 3488
rect 5085 3454 5095 3488
rect 5134 3454 5153 3488
rect 5153 3454 5168 3488
rect 5207 3454 5221 3488
rect 5221 3454 5241 3488
rect 5280 3454 5289 3488
rect 5289 3454 5314 3488
rect 5353 3454 5357 3488
rect 5357 3454 5387 3488
rect 5426 3454 5459 3488
rect 5459 3454 5460 3488
rect 5499 3454 5527 3488
rect 5527 3454 5533 3488
rect 5572 3454 5595 3488
rect 5595 3454 5606 3488
rect 5645 3454 5663 3488
rect 5663 3454 5679 3488
rect 5718 3454 5731 3488
rect 5731 3454 5752 3488
rect 5791 3454 5799 3488
rect 5799 3454 5825 3488
rect 5864 3454 5867 3488
rect 5867 3454 5898 3488
rect 5937 3454 5969 3488
rect 5969 3454 5971 3488
rect 6010 3454 6037 3488
rect 6037 3454 6044 3488
rect 6083 3454 6105 3488
rect 6105 3454 6117 3488
rect 6156 3454 6173 3488
rect 6173 3454 6190 3488
rect 6229 3454 6241 3488
rect 6241 3454 6263 3488
rect 6302 3454 6309 3488
rect 6309 3454 6336 3488
rect 6375 3454 6377 3488
rect 6377 3454 6409 3488
rect 6448 3454 6479 3488
rect 6479 3454 6482 3488
rect 6521 3454 6547 3488
rect 6547 3454 6555 3488
rect 6594 3454 6615 3488
rect 6615 3454 6628 3488
rect 6667 3454 6683 3488
rect 6683 3454 6701 3488
rect 6740 3454 6751 3488
rect 6751 3454 6774 3488
rect 6813 3454 6819 3488
rect 6819 3454 6847 3488
rect 6886 3454 6887 3488
rect 6887 3454 6920 3488
rect 6959 3454 6989 3488
rect 6989 3454 6993 3488
rect 7032 3454 7057 3488
rect 7057 3454 7066 3488
rect 7105 3454 7125 3488
rect 7125 3454 7139 3488
rect 7178 3454 7193 3488
rect 7193 3454 7212 3488
rect 7251 3454 7261 3488
rect 7261 3454 7285 3488
rect 7324 3454 7329 3488
rect 7329 3454 7358 3488
rect 7397 3454 7431 3488
rect 7913 3822 7947 3842
rect 7913 3808 7947 3822
rect 68 3388 102 3422
rect 68 3315 102 3349
rect 68 3261 102 3276
rect 68 3242 102 3261
rect 7913 3754 7947 3760
rect 7913 3726 7947 3754
rect 9734 3837 9738 3943
rect 9738 3837 9908 3943
rect 9908 3837 9912 3943
rect 8029 3714 8063 3748
rect 8104 3714 8138 3748
rect 8179 3714 8213 3748
rect 8254 3714 8288 3748
rect 8328 3714 8362 3748
rect 8402 3714 8436 3748
rect 8476 3714 8510 3748
rect 8550 3714 8584 3748
rect 8867 3744 8901 3778
rect 8948 3744 8982 3778
rect 9029 3744 9063 3778
rect 9110 3744 9144 3778
rect 9191 3744 9225 3778
rect 9271 3744 9305 3778
rect 9351 3744 9385 3778
rect 7913 3652 7947 3679
rect 7913 3645 7947 3652
rect 8029 3604 8063 3638
rect 8101 3604 8135 3638
rect 8173 3604 8207 3638
rect 7913 3584 7947 3598
rect 7913 3564 7947 3584
rect 7913 3516 7947 3517
rect 7913 3483 7947 3516
rect 8867 3568 8901 3602
rect 8942 3568 8976 3602
rect 9017 3568 9051 3602
rect 9092 3568 9126 3602
rect 9166 3568 9200 3602
rect 9240 3568 9274 3602
rect 9314 3568 9348 3602
rect 9388 3568 9422 3602
rect 8029 3083 8063 3117
rect 8101 3083 8135 3117
rect 8173 3083 8207 3117
rect 8377 3477 8411 3511
rect 8459 3477 8493 3511
rect 8541 3477 8575 3511
rect 8622 3477 8656 3511
rect 8703 3477 8737 3511
rect 8789 3480 8823 3514
rect 8861 3480 8895 3514
rect 9750 3397 9784 3431
rect 9825 3397 9859 3431
rect 9900 3397 9908 3431
rect 9908 3397 9934 3431
rect 9975 3397 10009 3431
rect 10050 3397 10084 3431
rect 10125 3397 10159 3431
rect 10200 3397 10234 3431
rect 10275 3397 10309 3431
rect 10350 3397 10384 3431
rect 10425 3397 10459 3431
rect 10500 3397 10534 3431
rect 10574 3397 10608 3431
rect 10648 3397 10682 3431
rect 10722 3397 10756 3431
rect 10796 3397 10830 3431
rect 10870 3397 10904 3431
rect 10944 3397 10978 3431
rect 11018 3397 11052 3431
rect 11092 3397 11126 3431
rect 11166 3397 11200 3431
rect 11240 3397 11274 3431
rect 8467 3083 8501 3117
rect 8542 3083 8576 3117
rect 8617 3083 8651 3117
rect 8692 3083 8726 3117
rect 8767 3083 8801 3117
rect 8841 3083 8875 3117
rect 8915 3083 8949 3117
rect 8989 3083 9023 3117
rect 9063 3083 9097 3117
rect 9137 3083 9171 3117
rect 9211 3083 9245 3117
rect 9285 3083 9319 3117
rect 9359 3083 9393 3117
rect 8197 3009 8231 3043
rect 8269 3009 8303 3043
rect 8072 2877 8106 2911
rect 8148 2877 8182 2911
rect 8224 2877 8258 2911
rect 8300 2877 8334 2911
rect 8376 2877 8410 2911
rect 8452 2877 8486 2911
rect 8528 2877 8562 2911
rect 8604 2877 8638 2911
rect 8680 2877 8714 2911
rect 8756 2877 8790 2911
rect 8832 2877 8866 2911
rect 8908 2877 8942 2911
rect 8984 2877 9018 2911
rect 9061 2877 9095 2911
rect 9138 2877 9172 2911
rect 9215 2877 9249 2911
rect 7913 2870 7947 2871
rect 7913 2837 7947 2870
rect 7913 2768 7947 2798
rect 7913 2764 7947 2768
rect 7913 2700 7947 2725
rect 7913 2691 7947 2700
rect 7913 2632 7947 2652
rect 7913 2618 7947 2632
rect 7913 2564 7947 2579
rect 7913 2545 7947 2564
rect 7913 2496 7947 2506
rect 7913 2472 7947 2496
rect 7913 2428 7947 2433
rect 7913 2399 7947 2428
rect 7913 2326 7947 2360
rect 7913 2258 7947 2287
rect 7913 2253 7947 2258
rect 7913 2190 7947 2214
rect 7913 2180 7947 2190
rect 7913 2122 7947 2141
rect 7913 2107 7947 2122
rect 7913 2054 7947 2068
rect 7913 2034 7947 2054
rect 7913 1986 7947 1995
rect 7913 1961 7947 1986
rect 7913 1918 7947 1922
rect 7913 1888 7947 1918
rect 7913 1816 7947 1849
rect 7913 1815 7947 1816
rect 7913 1748 7947 1776
rect 7913 1742 7947 1748
rect 7913 1680 7947 1703
rect 7913 1669 7947 1680
rect 7913 1612 7947 1630
rect 7913 1596 7947 1612
rect 7913 1544 7947 1557
rect 7913 1523 7947 1544
rect 7913 1476 7947 1484
rect 7913 1450 7947 1476
rect 7913 1408 7947 1411
rect 7913 1377 7947 1408
rect 7913 1306 7947 1338
rect 7913 1304 7947 1306
rect 7913 1238 7947 1265
rect 7913 1231 7947 1238
rect 7913 1170 7947 1192
rect 7913 1158 7947 1170
rect 7913 1102 7947 1119
rect 7913 1085 7947 1102
rect 7913 1034 7947 1046
rect 7913 1012 7947 1034
rect 7913 966 7947 973
rect 7913 939 7947 966
rect 7913 898 7947 900
rect 7913 866 7947 898
rect 8053 2783 8087 2817
rect 8053 2711 8087 2745
rect 8053 2639 8087 2673
rect 8965 2783 8999 2817
rect 8965 2711 8999 2745
rect 8053 2567 8087 2601
rect 8053 2495 8087 2529
rect 8053 2423 8087 2457
rect 8053 2351 8087 2385
rect 8053 2279 8087 2313
rect 8053 2207 8087 2241
rect 8053 2135 8087 2169
rect 8053 2063 8087 2097
rect 8053 1991 8087 2025
rect 8053 1919 8087 1953
rect 8053 1847 8087 1881
rect 8053 1775 8087 1809
rect 8053 1703 8087 1737
rect 8053 1631 8087 1665
rect 8053 1559 8087 1593
rect 8053 1487 8087 1521
rect 8053 1415 8087 1449
rect 8053 1343 8087 1377
rect 8053 1271 8087 1305
rect 8053 1199 8087 1233
rect 8053 1127 8087 1161
rect 8053 1055 8087 1089
rect 8053 983 8087 1017
rect 8053 910 8087 944
rect 8053 837 8087 871
rect 8509 2625 8543 2659
rect 8509 2551 8543 2585
rect 8509 2477 8543 2511
rect 8509 2403 8543 2437
rect 8509 2329 8543 2363
rect 8509 2255 8543 2289
rect 8509 2181 8543 2215
rect 8509 2107 8543 2141
rect 8509 2033 8543 2067
rect 8509 1959 8543 1993
rect 8509 1885 8543 1919
rect 8509 1811 8543 1845
rect 8509 1737 8543 1771
rect 8509 1662 8543 1696
rect 8509 1587 8543 1621
rect 8509 1512 8543 1546
rect 8509 1437 8543 1471
rect 8509 1362 8543 1396
rect 8509 1287 8543 1321
rect 8509 1212 8543 1246
rect 8509 1137 8543 1171
rect 8509 1062 8543 1096
rect 8509 987 8543 1021
rect 8509 912 8543 946
rect 8509 837 8543 871
rect 8965 2639 8999 2673
rect 9877 2783 9911 2817
rect 9877 2711 9911 2745
rect 8965 2567 8999 2601
rect 8965 2495 8999 2529
rect 8965 2423 8999 2457
rect 8965 2351 8999 2385
rect 8965 2279 8999 2313
rect 8965 2207 8999 2241
rect 8965 2135 8999 2169
rect 8965 2063 8999 2097
rect 8965 1991 8999 2025
rect 8965 1919 8999 1953
rect 8965 1847 8999 1881
rect 8965 1775 8999 1809
rect 8965 1703 8999 1737
rect 8965 1631 8999 1665
rect 8965 1559 8999 1593
rect 8965 1487 8999 1521
rect 8965 1415 8999 1449
rect 8965 1343 8999 1377
rect 8965 1271 8999 1305
rect 8965 1199 8999 1233
rect 8965 1127 8999 1161
rect 8965 1055 8999 1089
rect 8965 983 8999 1017
rect 8965 910 8999 944
rect 8965 837 8999 871
rect 9421 2625 9455 2659
rect 9421 2551 9455 2585
rect 9421 2477 9455 2511
rect 9421 2403 9455 2437
rect 9421 2329 9455 2363
rect 9421 2255 9455 2289
rect 9421 2181 9455 2215
rect 9421 2107 9455 2141
rect 9421 2033 9455 2067
rect 9421 1959 9455 1993
rect 9421 1885 9455 1919
rect 9421 1811 9455 1845
rect 9421 1737 9455 1771
rect 9421 1662 9455 1696
rect 9421 1587 9455 1621
rect 9421 1512 9455 1546
rect 9421 1437 9455 1471
rect 9421 1362 9455 1396
rect 9421 1287 9455 1321
rect 9421 1212 9455 1246
rect 9421 1137 9455 1171
rect 9421 1062 9455 1096
rect 9421 987 9455 1021
rect 9421 912 9455 946
rect 9421 837 9455 871
rect 9877 2639 9911 2673
rect 10789 2783 10823 2817
rect 10789 2711 10823 2745
rect 9877 2567 9911 2601
rect 9877 2495 9911 2529
rect 9877 2423 9911 2457
rect 9877 2351 9911 2385
rect 9877 2279 9911 2313
rect 9877 2207 9911 2241
rect 9877 2135 9911 2169
rect 9877 2063 9911 2097
rect 9877 1991 9911 2025
rect 9877 1919 9911 1953
rect 9877 1847 9911 1881
rect 9877 1775 9911 1809
rect 9877 1703 9911 1737
rect 9877 1631 9911 1665
rect 9877 1559 9911 1593
rect 9877 1487 9911 1521
rect 9877 1415 9911 1449
rect 9877 1343 9911 1377
rect 9877 1271 9911 1305
rect 9877 1199 9911 1233
rect 9877 1127 9911 1161
rect 9877 1055 9911 1089
rect 9877 983 9911 1017
rect 9877 910 9911 944
rect 9877 837 9911 871
rect 10333 2625 10367 2659
rect 10333 2551 10367 2585
rect 10333 2477 10367 2511
rect 10333 2403 10367 2437
rect 10333 2329 10367 2363
rect 10333 2255 10367 2289
rect 10333 2181 10367 2215
rect 10333 2107 10367 2141
rect 10333 2033 10367 2067
rect 10333 1959 10367 1993
rect 10333 1885 10367 1919
rect 10333 1811 10367 1845
rect 10333 1737 10367 1771
rect 10333 1662 10367 1696
rect 10333 1587 10367 1621
rect 10333 1512 10367 1546
rect 10333 1437 10367 1471
rect 10333 1362 10367 1396
rect 10333 1287 10367 1321
rect 10333 1212 10367 1246
rect 10333 1137 10367 1171
rect 10333 1062 10367 1096
rect 10333 987 10367 1021
rect 10333 912 10367 946
rect 10333 837 10367 871
rect 10789 2639 10823 2673
rect 10789 2567 10823 2601
rect 10789 2495 10823 2529
rect 10789 2423 10823 2457
rect 10789 2351 10823 2385
rect 10789 2279 10823 2313
rect 10789 2207 10823 2241
rect 10789 2135 10823 2169
rect 10789 2063 10823 2097
rect 10789 1991 10823 2025
rect 10789 1919 10823 1953
rect 10789 1847 10823 1881
rect 10789 1775 10823 1809
rect 10789 1703 10823 1737
rect 10789 1631 10823 1665
rect 10789 1559 10823 1593
rect 10789 1487 10823 1521
rect 10789 1415 10823 1449
rect 10789 1343 10823 1377
rect 10789 1271 10823 1305
rect 10789 1199 10823 1233
rect 10789 1127 10823 1161
rect 10789 1055 10823 1089
rect 10789 983 10823 1017
rect 10789 910 10823 944
rect 10789 837 10823 871
rect 10929 2809 10963 2817
rect 10929 2783 10963 2809
rect 10929 2741 10963 2744
rect 10929 2710 10963 2741
rect 10929 2639 10963 2671
rect 10929 2637 10963 2639
rect 10929 2571 10963 2598
rect 10929 2564 10963 2571
rect 10929 2503 10963 2525
rect 10929 2491 10963 2503
rect 10929 2435 10963 2452
rect 10929 2418 10963 2435
rect 10929 2367 10963 2379
rect 10929 2345 10963 2367
rect 10929 2299 10963 2306
rect 10929 2272 10963 2299
rect 10929 2231 10963 2233
rect 10929 2199 10963 2231
rect 10929 2129 10963 2159
rect 10929 2125 10963 2129
rect 10929 2061 10963 2085
rect 10929 2051 10963 2061
rect 10929 1993 10963 2011
rect 10929 1977 10963 1993
rect 10929 1925 10963 1937
rect 10929 1903 10963 1925
rect 10929 1857 10963 1863
rect 10929 1829 10963 1857
rect 10929 1755 10963 1789
rect 10929 1687 10963 1715
rect 10929 1681 10963 1687
rect 10929 1619 10963 1641
rect 10929 1607 10963 1619
rect 10929 1551 10963 1567
rect 10929 1533 10963 1551
rect 10929 1483 10963 1493
rect 10929 1459 10963 1483
rect 10929 1415 10963 1419
rect 10929 1385 10963 1415
rect 10929 1313 10963 1345
rect 10929 1311 10963 1313
rect 10929 1245 10963 1271
rect 10929 1237 10963 1245
rect 10929 1177 10963 1197
rect 10929 1163 10963 1177
rect 10929 1109 10963 1123
rect 10929 1089 10963 1109
rect 10929 1041 10963 1049
rect 10929 1015 10963 1041
rect 10929 973 10963 975
rect 10929 941 10963 973
rect 10929 871 10963 901
rect 10929 867 10963 871
rect 7913 796 7947 827
rect 7913 793 7947 796
rect 10929 803 10963 827
rect 10929 793 10963 803
rect 7919 721 7937 755
rect 7937 721 7953 755
rect 7992 721 8005 755
rect 8005 721 8026 755
rect 8065 721 8073 755
rect 8073 721 8099 755
rect 8138 721 8141 755
rect 8141 721 8172 755
rect 8211 721 8243 755
rect 8243 721 8245 755
rect 8284 721 8311 755
rect 8311 721 8318 755
rect 8357 721 8379 755
rect 8379 721 8391 755
rect 8430 721 8447 755
rect 8447 721 8464 755
rect 8503 721 8515 755
rect 8515 721 8537 755
rect 8576 721 8583 755
rect 8583 721 8610 755
rect 8649 721 8651 755
rect 8651 721 8683 755
rect 8722 721 8753 755
rect 8753 721 8756 755
rect 8795 721 8822 755
rect 8822 721 8829 755
rect 8868 721 8891 755
rect 8891 721 8902 755
rect 8941 721 8960 755
rect 8960 721 8975 755
rect 9014 721 9029 755
rect 9029 721 9048 755
rect 9087 721 9098 755
rect 9098 721 9121 755
rect 9160 721 9167 755
rect 9167 721 9194 755
rect 9233 721 9236 755
rect 9236 721 9267 755
rect 9306 721 9339 755
rect 9339 721 9340 755
rect 9379 721 9408 755
rect 9408 721 9413 755
rect 9452 721 9477 755
rect 9477 721 9486 755
rect 9525 721 9546 755
rect 9546 721 9559 755
rect 9598 721 9615 755
rect 9615 721 9632 755
rect 9671 721 9684 755
rect 9684 721 9705 755
rect 9744 721 9753 755
rect 9753 721 9778 755
rect 9817 721 9822 755
rect 9822 721 9851 755
rect 9890 721 9891 755
rect 9891 721 9924 755
rect 9963 721 9995 755
rect 9995 721 9997 755
rect 10036 721 10070 755
rect 10109 721 10143 755
rect 10183 721 10217 755
rect 10257 721 10291 755
rect 10331 721 10365 755
rect 10405 721 10439 755
rect 10479 721 10513 755
rect 10553 721 10587 755
rect 10627 721 10661 755
rect 10701 721 10735 755
rect 10775 721 10809 755
rect 10849 721 10883 755
rect 10923 721 10957 755
rect 7913 653 7947 683
rect 7913 649 7947 653
rect 7913 585 7947 601
rect 7913 567 7947 585
rect 7913 517 7947 519
rect 7913 485 7947 517
rect 7913 415 7947 436
rect 7913 402 7947 415
rect 7913 347 7947 353
rect 7913 319 7937 347
rect 7937 319 7947 347
rect 7985 313 8006 347
rect 8006 313 8019 347
rect 8058 313 8075 347
rect 8075 313 8092 347
rect 8131 313 8144 347
rect 8144 313 8165 347
rect 8204 313 8213 347
rect 8213 313 8238 347
rect 8277 313 8282 347
rect 8282 313 8311 347
rect 8350 313 8351 347
rect 8351 313 8384 347
rect 8423 313 8454 347
rect 8454 313 8457 347
rect 8496 313 8523 347
rect 8523 313 8530 347
rect 8569 313 8592 347
rect 8592 313 8603 347
rect 8642 313 8661 347
rect 8661 313 8676 347
rect 8715 313 8730 347
rect 8730 313 8749 347
rect 8788 313 8799 347
rect 8799 313 8822 347
rect 8861 313 8868 347
rect 8868 313 8895 347
rect 8934 313 8937 347
rect 8937 313 8968 347
rect 9007 313 9041 347
rect 9081 313 9110 347
rect 9110 313 9115 347
rect 9155 313 9179 347
rect 9179 313 9189 347
rect 9229 313 9248 347
rect 9248 313 9263 347
rect 9303 313 9317 347
rect 9317 313 9337 347
rect 9377 313 9386 347
rect 9386 313 9411 347
rect 9451 313 9455 347
rect 9455 313 9485 347
rect 9525 313 9558 347
rect 9558 313 9559 347
rect 9599 313 9627 347
rect 9627 313 9633 347
rect 9673 313 9696 347
rect 9696 313 9707 347
rect 9747 313 9765 347
rect 9765 313 9781 347
rect 9821 313 9834 347
rect 9834 313 9855 347
rect 9895 313 9903 347
rect 9903 313 9929 347
rect 9969 313 9972 347
rect 9972 313 10003 347
rect 10043 313 10076 347
rect 10076 313 10077 347
rect 10117 313 10145 347
rect 10145 313 10151 347
rect 10191 313 10214 347
rect 10214 313 10225 347
rect 10265 313 10283 347
rect 10283 313 10299 347
rect 10339 313 10352 347
rect 10352 313 10373 347
rect 10413 313 10421 347
rect 10421 313 10447 347
rect 10487 313 10490 347
rect 10490 313 10521 347
rect 10561 313 10593 347
rect 10593 313 10595 347
rect 10635 313 10662 347
rect 10662 313 10669 347
rect 10709 313 10731 347
rect 10731 313 10743 347
rect 10783 313 10800 347
rect 10800 313 10817 347
rect 10857 313 10869 347
rect 10869 313 10891 347
rect 12552 3339 12574 3373
rect 12574 3339 12586 3373
rect 12629 3339 12663 3373
rect 12706 3339 12740 3373
rect 12783 3339 12808 3373
rect 12808 3339 12817 3373
rect 12860 3339 12876 3373
rect 12876 3339 12894 3373
rect 12938 3339 12944 3373
rect 12944 3339 12972 3373
rect 13016 3339 13046 3373
rect 13046 3339 13050 3373
rect 13094 3339 13114 3373
rect 13114 3339 13128 3373
rect 13172 3339 13182 3373
rect 13182 3339 13206 3373
rect 13250 3339 13284 3373
rect 13328 3339 13362 3373
rect 13366 3237 13400 3263
rect 13366 3229 13400 3237
rect 12780 3157 12814 3191
rect 12852 3157 12886 3191
rect 12924 3157 12958 3191
rect 12996 3157 13030 3191
rect 13068 3157 13102 3191
rect 13140 3157 13174 3191
rect 13366 3169 13400 3191
rect 13366 3157 13400 3169
rect 12624 3077 12658 3111
rect 12696 3077 12730 3111
rect 13366 3101 13400 3119
rect 13366 3085 13400 3101
rect 13366 3013 13400 3047
rect 12552 2975 12586 3009
rect 12630 2975 12652 3009
rect 12652 2975 12664 3009
rect 12707 2975 12720 3009
rect 12720 2975 12741 3009
rect 12784 2975 12788 3009
rect 12788 2975 12818 3009
rect 12861 2975 12890 3009
rect 12890 2975 12895 3009
rect 12938 2975 12958 3009
rect 12958 2975 12972 3009
rect 13015 2975 13026 3009
rect 13026 2975 13049 3009
rect 13092 2975 13094 3009
rect 13094 2975 13126 3009
rect 13169 2975 13196 3009
rect 13196 2975 13203 3009
rect 13246 2975 13264 3009
rect 13264 2975 13280 3009
rect 11448 2695 11482 2714
rect 11522 2695 11556 2714
rect 11596 2695 11630 2714
rect 11670 2695 11704 2714
rect 11744 2695 11778 2714
rect 11818 2695 11852 2714
rect 11892 2695 11926 2714
rect 11966 2695 12000 2714
rect 12040 2695 12074 2714
rect 12114 2695 12148 2714
rect 12188 2695 12222 2714
rect 12262 2695 12296 2714
rect 12336 2695 12370 2714
rect 12410 2695 12444 2714
rect 12484 2695 12518 2714
rect 11448 2680 11476 2695
rect 11476 2680 11482 2695
rect 11522 2680 11546 2695
rect 11546 2680 11556 2695
rect 11596 2680 11616 2695
rect 11616 2680 11630 2695
rect 11670 2680 11686 2695
rect 11686 2680 11704 2695
rect 11744 2680 11756 2695
rect 11756 2680 11778 2695
rect 11818 2680 11826 2695
rect 11826 2680 11852 2695
rect 11892 2680 11896 2695
rect 11896 2680 11926 2695
rect 11966 2680 12000 2695
rect 12040 2680 12070 2695
rect 12070 2680 12074 2695
rect 12114 2680 12140 2695
rect 12140 2680 12148 2695
rect 12188 2680 12210 2695
rect 12210 2680 12222 2695
rect 12262 2680 12280 2695
rect 12280 2680 12296 2695
rect 12336 2680 12350 2695
rect 12350 2680 12370 2695
rect 12410 2680 12419 2695
rect 12419 2680 12444 2695
rect 12484 2680 12488 2695
rect 12488 2680 12518 2695
rect 12558 2680 12592 2714
rect 12632 2695 12666 2714
rect 12706 2695 12740 2714
rect 12780 2695 12814 2714
rect 12854 2695 12888 2714
rect 12928 2695 12962 2714
rect 13002 2695 13036 2714
rect 13076 2695 13110 2714
rect 13150 2695 13184 2714
rect 13224 2695 13258 2714
rect 13298 2695 13332 2714
rect 13372 2695 13406 2714
rect 13446 2695 13480 2714
rect 13520 2695 13554 2714
rect 13594 2695 13628 2714
rect 13668 2695 13702 2714
rect 13741 2695 13775 2714
rect 13814 2695 13848 2714
rect 13887 2695 13921 2714
rect 13960 2695 13994 2714
rect 14033 2695 14067 2714
rect 12632 2680 12661 2695
rect 12661 2680 12666 2695
rect 12706 2680 12730 2695
rect 12730 2680 12740 2695
rect 12780 2680 12799 2695
rect 12799 2680 12814 2695
rect 12854 2680 12868 2695
rect 12868 2680 12888 2695
rect 12928 2680 12937 2695
rect 12937 2680 12962 2695
rect 13002 2680 13006 2695
rect 13006 2680 13036 2695
rect 13076 2680 13109 2695
rect 13109 2680 13110 2695
rect 13150 2680 13178 2695
rect 13178 2680 13184 2695
rect 13224 2680 13247 2695
rect 13247 2680 13258 2695
rect 13298 2680 13316 2695
rect 13316 2680 13332 2695
rect 13372 2680 13385 2695
rect 13385 2680 13406 2695
rect 13446 2680 13454 2695
rect 13454 2680 13480 2695
rect 13520 2680 13523 2695
rect 13523 2680 13554 2695
rect 13594 2680 13627 2695
rect 13627 2680 13628 2695
rect 13668 2680 13696 2695
rect 13696 2680 13702 2695
rect 13741 2680 13765 2695
rect 13765 2680 13775 2695
rect 13814 2680 13834 2695
rect 13834 2680 13848 2695
rect 13887 2680 13903 2695
rect 13903 2680 13921 2695
rect 13960 2680 13972 2695
rect 13972 2680 13994 2695
rect 14033 2680 14041 2695
rect 14041 2680 14067 2695
rect 11448 2627 11482 2642
rect 11522 2627 11556 2642
rect 11596 2627 11630 2642
rect 11670 2627 11704 2642
rect 11744 2627 11778 2642
rect 11818 2627 11852 2642
rect 11892 2627 11926 2642
rect 11966 2627 12000 2642
rect 12040 2627 12074 2642
rect 12114 2627 12148 2642
rect 12188 2627 12222 2642
rect 12262 2627 12296 2642
rect 12336 2627 12370 2642
rect 12410 2627 12444 2642
rect 12484 2627 12518 2642
rect 11448 2608 11476 2627
rect 11476 2608 11482 2627
rect 11522 2608 11546 2627
rect 11546 2608 11556 2627
rect 11596 2608 11616 2627
rect 11616 2608 11630 2627
rect 11670 2608 11686 2627
rect 11686 2608 11704 2627
rect 11744 2608 11756 2627
rect 11756 2608 11778 2627
rect 11818 2608 11826 2627
rect 11826 2608 11852 2627
rect 11892 2608 11896 2627
rect 11896 2608 11926 2627
rect 11966 2608 12000 2627
rect 12040 2608 12070 2627
rect 12070 2608 12074 2627
rect 12114 2608 12140 2627
rect 12140 2608 12148 2627
rect 12188 2608 12210 2627
rect 12210 2608 12222 2627
rect 12262 2608 12280 2627
rect 12280 2608 12296 2627
rect 12336 2608 12350 2627
rect 12350 2608 12370 2627
rect 12410 2608 12419 2627
rect 12419 2608 12444 2627
rect 12484 2608 12488 2627
rect 12488 2608 12518 2627
rect 12558 2608 12592 2642
rect 12632 2627 12666 2642
rect 12706 2627 12740 2642
rect 12780 2627 12814 2642
rect 12854 2627 12888 2642
rect 12928 2627 12962 2642
rect 13002 2627 13036 2642
rect 13076 2627 13110 2642
rect 13150 2627 13184 2642
rect 13224 2627 13258 2642
rect 13298 2627 13332 2642
rect 13372 2627 13406 2642
rect 13446 2627 13480 2642
rect 13520 2627 13554 2642
rect 13594 2627 13628 2642
rect 13668 2627 13702 2642
rect 13741 2627 13775 2642
rect 13814 2627 13848 2642
rect 13887 2627 13921 2642
rect 13960 2627 13994 2642
rect 14033 2627 14067 2642
rect 12632 2608 12661 2627
rect 12661 2608 12666 2627
rect 12706 2608 12730 2627
rect 12730 2608 12740 2627
rect 12780 2608 12799 2627
rect 12799 2608 12814 2627
rect 12854 2608 12868 2627
rect 12868 2608 12888 2627
rect 12928 2608 12937 2627
rect 12937 2608 12962 2627
rect 13002 2608 13006 2627
rect 13006 2608 13036 2627
rect 13076 2608 13109 2627
rect 13109 2608 13110 2627
rect 13150 2608 13178 2627
rect 13178 2608 13184 2627
rect 13224 2608 13247 2627
rect 13247 2608 13258 2627
rect 13298 2608 13316 2627
rect 13316 2608 13332 2627
rect 13372 2608 13385 2627
rect 13385 2608 13406 2627
rect 13446 2608 13454 2627
rect 13454 2608 13480 2627
rect 13520 2608 13523 2627
rect 13523 2608 13554 2627
rect 13594 2608 13627 2627
rect 13627 2608 13628 2627
rect 13668 2608 13696 2627
rect 13696 2608 13702 2627
rect 13741 2608 13765 2627
rect 13765 2608 13775 2627
rect 13814 2608 13834 2627
rect 13834 2608 13848 2627
rect 13887 2608 13903 2627
rect 13903 2608 13921 2627
rect 13960 2608 13972 2627
rect 13972 2608 13994 2627
rect 14033 2608 14041 2627
rect 14041 2608 14067 2627
rect 11448 2559 11482 2570
rect 11522 2559 11556 2570
rect 11596 2559 11630 2570
rect 11670 2559 11704 2570
rect 11744 2559 11778 2570
rect 11818 2559 11852 2570
rect 11892 2559 11926 2570
rect 11966 2559 12000 2570
rect 12040 2559 12074 2570
rect 12114 2559 12148 2570
rect 12188 2559 12222 2570
rect 12262 2559 12296 2570
rect 12336 2559 12370 2570
rect 12410 2559 12444 2570
rect 12484 2559 12518 2570
rect 11448 2536 11476 2559
rect 11476 2536 11482 2559
rect 11522 2536 11546 2559
rect 11546 2536 11556 2559
rect 11596 2536 11616 2559
rect 11616 2536 11630 2559
rect 11670 2536 11686 2559
rect 11686 2536 11704 2559
rect 11744 2536 11756 2559
rect 11756 2536 11778 2559
rect 11818 2536 11826 2559
rect 11826 2536 11852 2559
rect 11892 2536 11896 2559
rect 11896 2536 11926 2559
rect 11966 2536 12000 2559
rect 12040 2536 12070 2559
rect 12070 2536 12074 2559
rect 12114 2536 12140 2559
rect 12140 2536 12148 2559
rect 12188 2536 12210 2559
rect 12210 2536 12222 2559
rect 12262 2536 12280 2559
rect 12280 2536 12296 2559
rect 12336 2536 12350 2559
rect 12350 2536 12370 2559
rect 12410 2536 12419 2559
rect 12419 2536 12444 2559
rect 12484 2536 12488 2559
rect 12488 2536 12518 2559
rect 12558 2536 12592 2570
rect 12632 2559 12666 2570
rect 12706 2559 12740 2570
rect 12780 2559 12814 2570
rect 12854 2559 12888 2570
rect 12928 2559 12962 2570
rect 13002 2559 13036 2570
rect 13076 2559 13110 2570
rect 13150 2559 13184 2570
rect 13224 2559 13258 2570
rect 13298 2559 13332 2570
rect 13372 2559 13406 2570
rect 13446 2559 13480 2570
rect 13520 2559 13554 2570
rect 13594 2559 13628 2570
rect 13668 2559 13702 2570
rect 13741 2559 13775 2570
rect 13814 2559 13848 2570
rect 13887 2559 13921 2570
rect 13960 2559 13994 2570
rect 14033 2559 14067 2570
rect 12632 2536 12661 2559
rect 12661 2536 12666 2559
rect 12706 2536 12730 2559
rect 12730 2536 12740 2559
rect 12780 2536 12799 2559
rect 12799 2536 12814 2559
rect 12854 2536 12868 2559
rect 12868 2536 12888 2559
rect 12928 2536 12937 2559
rect 12937 2536 12962 2559
rect 13002 2536 13006 2559
rect 13006 2536 13036 2559
rect 13076 2536 13109 2559
rect 13109 2536 13110 2559
rect 13150 2536 13178 2559
rect 13178 2536 13184 2559
rect 13224 2536 13247 2559
rect 13247 2536 13258 2559
rect 13298 2536 13316 2559
rect 13316 2536 13332 2559
rect 13372 2536 13385 2559
rect 13385 2536 13406 2559
rect 13446 2536 13454 2559
rect 13454 2536 13480 2559
rect 13520 2536 13523 2559
rect 13523 2536 13554 2559
rect 13594 2536 13627 2559
rect 13627 2536 13628 2559
rect 13668 2536 13696 2559
rect 13696 2536 13702 2559
rect 13741 2536 13765 2559
rect 13765 2536 13775 2559
rect 13814 2536 13834 2559
rect 13834 2536 13848 2559
rect 13887 2536 13903 2559
rect 13903 2536 13921 2559
rect 13960 2536 13972 2559
rect 13972 2536 13994 2559
rect 14033 2536 14041 2559
rect 14041 2536 14067 2559
rect 11448 2491 11482 2498
rect 11522 2491 11556 2498
rect 11596 2491 11630 2498
rect 11670 2491 11704 2498
rect 11744 2491 11778 2498
rect 11818 2491 11852 2498
rect 11892 2491 11926 2498
rect 11966 2491 12000 2498
rect 12040 2491 12074 2498
rect 12114 2491 12148 2498
rect 12188 2491 12222 2498
rect 12262 2491 12296 2498
rect 12336 2491 12370 2498
rect 12410 2491 12444 2498
rect 12484 2491 12518 2498
rect 11448 2464 11476 2491
rect 11476 2464 11482 2491
rect 11522 2464 11546 2491
rect 11546 2464 11556 2491
rect 11596 2464 11616 2491
rect 11616 2464 11630 2491
rect 11670 2464 11686 2491
rect 11686 2464 11704 2491
rect 11744 2464 11756 2491
rect 11756 2464 11778 2491
rect 11818 2464 11826 2491
rect 11826 2464 11852 2491
rect 11892 2464 11896 2491
rect 11896 2464 11926 2491
rect 11966 2464 12000 2491
rect 12040 2464 12070 2491
rect 12070 2464 12074 2491
rect 12114 2464 12140 2491
rect 12140 2464 12148 2491
rect 12188 2464 12210 2491
rect 12210 2464 12222 2491
rect 12262 2464 12280 2491
rect 12280 2464 12296 2491
rect 12336 2464 12350 2491
rect 12350 2464 12370 2491
rect 12410 2464 12419 2491
rect 12419 2464 12444 2491
rect 12484 2464 12488 2491
rect 12488 2464 12518 2491
rect 12558 2464 12592 2498
rect 12632 2491 12666 2498
rect 12706 2491 12740 2498
rect 12780 2491 12814 2498
rect 12854 2491 12888 2498
rect 12928 2491 12962 2498
rect 13002 2491 13036 2498
rect 13076 2491 13110 2498
rect 13150 2491 13184 2498
rect 13224 2491 13258 2498
rect 13298 2491 13332 2498
rect 13372 2491 13406 2498
rect 13446 2491 13480 2498
rect 13520 2491 13554 2498
rect 13594 2491 13628 2498
rect 13668 2491 13702 2498
rect 13741 2491 13775 2498
rect 13814 2491 13848 2498
rect 13887 2491 13921 2498
rect 13960 2491 13994 2498
rect 14033 2491 14067 2498
rect 12632 2464 12661 2491
rect 12661 2464 12666 2491
rect 12706 2464 12730 2491
rect 12730 2464 12740 2491
rect 12780 2464 12799 2491
rect 12799 2464 12814 2491
rect 12854 2464 12868 2491
rect 12868 2464 12888 2491
rect 12928 2464 12937 2491
rect 12937 2464 12962 2491
rect 13002 2464 13006 2491
rect 13006 2464 13036 2491
rect 13076 2464 13109 2491
rect 13109 2464 13110 2491
rect 13150 2464 13178 2491
rect 13178 2464 13184 2491
rect 13224 2464 13247 2491
rect 13247 2464 13258 2491
rect 13298 2464 13316 2491
rect 13316 2464 13332 2491
rect 13372 2464 13385 2491
rect 13385 2464 13406 2491
rect 13446 2464 13454 2491
rect 13454 2464 13480 2491
rect 13520 2464 13523 2491
rect 13523 2464 13554 2491
rect 13594 2464 13627 2491
rect 13627 2464 13628 2491
rect 13668 2464 13696 2491
rect 13696 2464 13702 2491
rect 13741 2464 13765 2491
rect 13765 2464 13775 2491
rect 13814 2464 13834 2491
rect 13834 2464 13848 2491
rect 13887 2464 13903 2491
rect 13903 2464 13921 2491
rect 13960 2464 13972 2491
rect 13972 2464 13994 2491
rect 14033 2464 14041 2491
rect 14041 2464 14067 2491
rect 11448 2423 11482 2426
rect 11522 2423 11556 2426
rect 11596 2423 11630 2426
rect 11670 2423 11704 2426
rect 11744 2423 11778 2426
rect 11818 2423 11852 2426
rect 11892 2423 11926 2426
rect 11966 2423 12000 2426
rect 12040 2423 12074 2426
rect 12114 2423 12148 2426
rect 12188 2423 12222 2426
rect 12262 2423 12296 2426
rect 12336 2423 12370 2426
rect 12410 2423 12444 2426
rect 12484 2423 12518 2426
rect 11448 2392 11476 2423
rect 11476 2392 11482 2423
rect 11522 2392 11546 2423
rect 11546 2392 11556 2423
rect 11596 2392 11616 2423
rect 11616 2392 11630 2423
rect 11670 2392 11686 2423
rect 11686 2392 11704 2423
rect 11744 2392 11756 2423
rect 11756 2392 11778 2423
rect 11818 2392 11826 2423
rect 11826 2392 11852 2423
rect 11892 2392 11896 2423
rect 11896 2392 11926 2423
rect 11966 2392 12000 2423
rect 12040 2392 12070 2423
rect 12070 2392 12074 2423
rect 12114 2392 12140 2423
rect 12140 2392 12148 2423
rect 12188 2392 12210 2423
rect 12210 2392 12222 2423
rect 12262 2392 12280 2423
rect 12280 2392 12296 2423
rect 12336 2392 12350 2423
rect 12350 2392 12370 2423
rect 12410 2392 12419 2423
rect 12419 2392 12444 2423
rect 12484 2392 12488 2423
rect 12488 2392 12518 2423
rect 12558 2392 12592 2426
rect 12632 2423 12666 2426
rect 12706 2423 12740 2426
rect 12780 2423 12814 2426
rect 12854 2423 12888 2426
rect 12928 2423 12962 2426
rect 13002 2423 13036 2426
rect 13076 2423 13110 2426
rect 13150 2423 13184 2426
rect 13224 2423 13258 2426
rect 13298 2423 13332 2426
rect 13372 2423 13406 2426
rect 13446 2423 13480 2426
rect 13520 2423 13554 2426
rect 13594 2423 13628 2426
rect 13668 2423 13702 2426
rect 13741 2423 13775 2426
rect 13814 2423 13848 2426
rect 13887 2423 13921 2426
rect 13960 2423 13994 2426
rect 14033 2423 14067 2426
rect 12632 2392 12661 2423
rect 12661 2392 12666 2423
rect 12706 2392 12730 2423
rect 12730 2392 12740 2423
rect 12780 2392 12799 2423
rect 12799 2392 12814 2423
rect 12854 2392 12868 2423
rect 12868 2392 12888 2423
rect 12928 2392 12937 2423
rect 12937 2392 12962 2423
rect 13002 2392 13006 2423
rect 13006 2392 13036 2423
rect 13076 2392 13109 2423
rect 13109 2392 13110 2423
rect 13150 2392 13178 2423
rect 13178 2392 13184 2423
rect 13224 2392 13247 2423
rect 13247 2392 13258 2423
rect 13298 2392 13316 2423
rect 13316 2392 13332 2423
rect 13372 2392 13385 2423
rect 13385 2392 13406 2423
rect 13446 2392 13454 2423
rect 13454 2392 13480 2423
rect 13520 2392 13523 2423
rect 13523 2392 13554 2423
rect 13594 2392 13627 2423
rect 13627 2392 13628 2423
rect 13668 2392 13696 2423
rect 13696 2392 13702 2423
rect 13741 2392 13765 2423
rect 13765 2392 13775 2423
rect 13814 2392 13834 2423
rect 13834 2392 13848 2423
rect 13887 2392 13903 2423
rect 13903 2392 13921 2423
rect 13960 2392 13972 2423
rect 13972 2392 13994 2423
rect 14033 2392 14041 2423
rect 14041 2392 14067 2423
rect 11448 2321 11476 2354
rect 11476 2321 11482 2354
rect 11522 2321 11546 2354
rect 11546 2321 11556 2354
rect 11596 2321 11616 2354
rect 11616 2321 11630 2354
rect 11670 2321 11686 2354
rect 11686 2321 11704 2354
rect 11744 2321 11756 2354
rect 11756 2321 11778 2354
rect 11818 2321 11826 2354
rect 11826 2321 11852 2354
rect 11892 2321 11896 2354
rect 11896 2321 11926 2354
rect 11966 2321 12000 2354
rect 12040 2321 12070 2354
rect 12070 2321 12074 2354
rect 12114 2321 12140 2354
rect 12140 2321 12148 2354
rect 12188 2321 12210 2354
rect 12210 2321 12222 2354
rect 12262 2321 12280 2354
rect 12280 2321 12296 2354
rect 12336 2321 12350 2354
rect 12350 2321 12370 2354
rect 12410 2321 12419 2354
rect 12419 2321 12444 2354
rect 12484 2321 12488 2354
rect 12488 2321 12518 2354
rect 11448 2320 11482 2321
rect 11522 2320 11556 2321
rect 11596 2320 11630 2321
rect 11670 2320 11704 2321
rect 11744 2320 11778 2321
rect 11818 2320 11852 2321
rect 11892 2320 11926 2321
rect 11966 2320 12000 2321
rect 12040 2320 12074 2321
rect 12114 2320 12148 2321
rect 12188 2320 12222 2321
rect 12262 2320 12296 2321
rect 12336 2320 12370 2321
rect 12410 2320 12444 2321
rect 12484 2320 12518 2321
rect 12558 2320 12592 2354
rect 12632 2321 12661 2354
rect 12661 2321 12666 2354
rect 12706 2321 12730 2354
rect 12730 2321 12740 2354
rect 12780 2321 12799 2354
rect 12799 2321 12814 2354
rect 12854 2321 12868 2354
rect 12868 2321 12888 2354
rect 12928 2321 12937 2354
rect 12937 2321 12962 2354
rect 13002 2321 13006 2354
rect 13006 2321 13036 2354
rect 13076 2321 13109 2354
rect 13109 2321 13110 2354
rect 13150 2321 13178 2354
rect 13178 2321 13184 2354
rect 13224 2321 13247 2354
rect 13247 2321 13258 2354
rect 13298 2321 13316 2354
rect 13316 2321 13332 2354
rect 13372 2321 13385 2354
rect 13385 2321 13406 2354
rect 13446 2321 13454 2354
rect 13454 2321 13480 2354
rect 13520 2321 13523 2354
rect 13523 2321 13554 2354
rect 13594 2321 13627 2354
rect 13627 2321 13628 2354
rect 13668 2321 13696 2354
rect 13696 2321 13702 2354
rect 13741 2321 13765 2354
rect 13765 2321 13775 2354
rect 13814 2321 13834 2354
rect 13834 2321 13848 2354
rect 13887 2321 13903 2354
rect 13903 2321 13921 2354
rect 13960 2321 13972 2354
rect 13972 2321 13994 2354
rect 14033 2321 14041 2354
rect 14041 2321 14067 2354
rect 12632 2320 12666 2321
rect 12706 2320 12740 2321
rect 12780 2320 12814 2321
rect 12854 2320 12888 2321
rect 12928 2320 12962 2321
rect 13002 2320 13036 2321
rect 13076 2320 13110 2321
rect 13150 2320 13184 2321
rect 13224 2320 13258 2321
rect 13298 2320 13332 2321
rect 13372 2320 13406 2321
rect 13446 2320 13480 2321
rect 13520 2320 13554 2321
rect 13594 2320 13628 2321
rect 13668 2320 13702 2321
rect 13741 2320 13775 2321
rect 13814 2320 13848 2321
rect 13887 2320 13921 2321
rect 13960 2320 13994 2321
rect 14033 2320 14067 2321
rect 11448 2253 11476 2282
rect 11476 2253 11482 2282
rect 11522 2253 11546 2282
rect 11546 2253 11556 2282
rect 11596 2253 11616 2282
rect 11616 2253 11630 2282
rect 11670 2253 11686 2282
rect 11686 2253 11704 2282
rect 11744 2253 11756 2282
rect 11756 2253 11778 2282
rect 11818 2253 11826 2282
rect 11826 2253 11852 2282
rect 11892 2253 11896 2282
rect 11896 2253 11926 2282
rect 11966 2253 12000 2282
rect 12040 2253 12070 2282
rect 12070 2253 12074 2282
rect 12114 2253 12140 2282
rect 12140 2253 12148 2282
rect 12188 2253 12210 2282
rect 12210 2253 12222 2282
rect 12262 2253 12280 2282
rect 12280 2253 12296 2282
rect 12336 2253 12350 2282
rect 12350 2253 12370 2282
rect 12410 2253 12419 2282
rect 12419 2253 12444 2282
rect 12484 2253 12488 2282
rect 12488 2253 12518 2282
rect 11448 2248 11482 2253
rect 11522 2248 11556 2253
rect 11596 2248 11630 2253
rect 11670 2248 11704 2253
rect 11744 2248 11778 2253
rect 11818 2248 11852 2253
rect 11892 2248 11926 2253
rect 11966 2248 12000 2253
rect 12040 2248 12074 2253
rect 12114 2248 12148 2253
rect 12188 2248 12222 2253
rect 12262 2248 12296 2253
rect 12336 2248 12370 2253
rect 12410 2248 12444 2253
rect 12484 2248 12518 2253
rect 12558 2248 12592 2282
rect 12632 2253 12661 2282
rect 12661 2253 12666 2282
rect 12706 2253 12730 2282
rect 12730 2253 12740 2282
rect 12780 2253 12799 2282
rect 12799 2253 12814 2282
rect 12854 2253 12868 2282
rect 12868 2253 12888 2282
rect 12928 2253 12937 2282
rect 12937 2253 12962 2282
rect 13002 2253 13006 2282
rect 13006 2253 13036 2282
rect 13076 2253 13109 2282
rect 13109 2253 13110 2282
rect 13150 2253 13178 2282
rect 13178 2253 13184 2282
rect 13224 2253 13247 2282
rect 13247 2253 13258 2282
rect 13298 2253 13316 2282
rect 13316 2253 13332 2282
rect 13372 2253 13385 2282
rect 13385 2253 13406 2282
rect 13446 2253 13454 2282
rect 13454 2253 13480 2282
rect 13520 2253 13523 2282
rect 13523 2253 13554 2282
rect 13594 2253 13627 2282
rect 13627 2253 13628 2282
rect 13668 2253 13696 2282
rect 13696 2253 13702 2282
rect 13741 2253 13765 2282
rect 13765 2253 13775 2282
rect 13814 2253 13834 2282
rect 13834 2253 13848 2282
rect 13887 2253 13903 2282
rect 13903 2253 13921 2282
rect 13960 2253 13972 2282
rect 13972 2253 13994 2282
rect 14033 2253 14041 2282
rect 14041 2253 14067 2282
rect 12632 2248 12666 2253
rect 12706 2248 12740 2253
rect 12780 2248 12814 2253
rect 12854 2248 12888 2253
rect 12928 2248 12962 2253
rect 13002 2248 13036 2253
rect 13076 2248 13110 2253
rect 13150 2248 13184 2253
rect 13224 2248 13258 2253
rect 13298 2248 13332 2253
rect 13372 2248 13406 2253
rect 13446 2248 13480 2253
rect 13520 2248 13554 2253
rect 13594 2248 13628 2253
rect 13668 2248 13702 2253
rect 13741 2248 13775 2253
rect 13814 2248 13848 2253
rect 13887 2248 13921 2253
rect 13960 2248 13994 2253
rect 14033 2248 14067 2253
rect 11448 2185 11476 2210
rect 11476 2185 11482 2210
rect 11522 2185 11546 2210
rect 11546 2185 11556 2210
rect 11596 2185 11616 2210
rect 11616 2185 11630 2210
rect 11670 2185 11686 2210
rect 11686 2185 11704 2210
rect 11744 2185 11756 2210
rect 11756 2185 11778 2210
rect 11818 2185 11826 2210
rect 11826 2185 11852 2210
rect 11892 2185 11896 2210
rect 11896 2185 11926 2210
rect 11966 2185 12000 2210
rect 12040 2185 12070 2210
rect 12070 2185 12074 2210
rect 12114 2185 12140 2210
rect 12140 2185 12148 2210
rect 12188 2185 12210 2210
rect 12210 2185 12222 2210
rect 12262 2185 12280 2210
rect 12280 2185 12296 2210
rect 12336 2185 12350 2210
rect 12350 2185 12370 2210
rect 12410 2185 12419 2210
rect 12419 2185 12444 2210
rect 12484 2185 12488 2210
rect 12488 2185 12518 2210
rect 11448 2176 11482 2185
rect 11522 2176 11556 2185
rect 11596 2176 11630 2185
rect 11670 2176 11704 2185
rect 11744 2176 11778 2185
rect 11818 2176 11852 2185
rect 11892 2176 11926 2185
rect 11966 2176 12000 2185
rect 12040 2176 12074 2185
rect 12114 2176 12148 2185
rect 12188 2176 12222 2185
rect 12262 2176 12296 2185
rect 12336 2176 12370 2185
rect 12410 2176 12444 2185
rect 12484 2176 12518 2185
rect 12558 2176 12592 2210
rect 12632 2185 12661 2210
rect 12661 2185 12666 2210
rect 12706 2185 12730 2210
rect 12730 2185 12740 2210
rect 12780 2185 12799 2210
rect 12799 2185 12814 2210
rect 12854 2185 12868 2210
rect 12868 2185 12888 2210
rect 12928 2185 12937 2210
rect 12937 2185 12962 2210
rect 13002 2185 13006 2210
rect 13006 2185 13036 2210
rect 13076 2185 13109 2210
rect 13109 2185 13110 2210
rect 13150 2185 13178 2210
rect 13178 2185 13184 2210
rect 13224 2185 13247 2210
rect 13247 2185 13258 2210
rect 13298 2185 13316 2210
rect 13316 2185 13332 2210
rect 13372 2185 13385 2210
rect 13385 2185 13406 2210
rect 13446 2185 13454 2210
rect 13454 2185 13480 2210
rect 13520 2185 13523 2210
rect 13523 2185 13554 2210
rect 13594 2185 13627 2210
rect 13627 2185 13628 2210
rect 13668 2185 13696 2210
rect 13696 2185 13702 2210
rect 13741 2185 13765 2210
rect 13765 2185 13775 2210
rect 13814 2185 13834 2210
rect 13834 2185 13848 2210
rect 13887 2185 13903 2210
rect 13903 2185 13921 2210
rect 13960 2185 13972 2210
rect 13972 2185 13994 2210
rect 14033 2185 14041 2210
rect 14041 2185 14067 2210
rect 12632 2176 12666 2185
rect 12706 2176 12740 2185
rect 12780 2176 12814 2185
rect 12854 2176 12888 2185
rect 12928 2176 12962 2185
rect 13002 2176 13036 2185
rect 13076 2176 13110 2185
rect 13150 2176 13184 2185
rect 13224 2176 13258 2185
rect 13298 2176 13332 2185
rect 13372 2176 13406 2185
rect 13446 2176 13480 2185
rect 13520 2176 13554 2185
rect 13594 2176 13628 2185
rect 13668 2176 13702 2185
rect 13741 2176 13775 2185
rect 13814 2176 13848 2185
rect 13887 2176 13921 2185
rect 13960 2176 13994 2185
rect 14033 2176 14067 2185
rect 11448 2117 11476 2138
rect 11476 2117 11482 2138
rect 11522 2117 11546 2138
rect 11546 2117 11556 2138
rect 11596 2117 11616 2138
rect 11616 2117 11630 2138
rect 11670 2117 11686 2138
rect 11686 2117 11704 2138
rect 11744 2117 11756 2138
rect 11756 2117 11778 2138
rect 11818 2117 11826 2138
rect 11826 2117 11852 2138
rect 11892 2117 11896 2138
rect 11896 2117 11926 2138
rect 11966 2117 12000 2138
rect 12040 2117 12070 2138
rect 12070 2117 12074 2138
rect 12114 2117 12140 2138
rect 12140 2117 12148 2138
rect 12188 2117 12210 2138
rect 12210 2117 12222 2138
rect 12262 2117 12280 2138
rect 12280 2117 12296 2138
rect 12336 2117 12350 2138
rect 12350 2117 12370 2138
rect 12410 2117 12419 2138
rect 12419 2117 12444 2138
rect 12484 2117 12488 2138
rect 12488 2117 12518 2138
rect 11448 2104 11482 2117
rect 11522 2104 11556 2117
rect 11596 2104 11630 2117
rect 11670 2104 11704 2117
rect 11744 2104 11778 2117
rect 11818 2104 11852 2117
rect 11892 2104 11926 2117
rect 11966 2104 12000 2117
rect 12040 2104 12074 2117
rect 12114 2104 12148 2117
rect 12188 2104 12222 2117
rect 12262 2104 12296 2117
rect 12336 2104 12370 2117
rect 12410 2104 12444 2117
rect 12484 2104 12518 2117
rect 12558 2104 12592 2138
rect 12632 2117 12661 2138
rect 12661 2117 12666 2138
rect 12706 2117 12730 2138
rect 12730 2117 12740 2138
rect 12780 2117 12799 2138
rect 12799 2117 12814 2138
rect 12854 2117 12868 2138
rect 12868 2117 12888 2138
rect 12928 2117 12937 2138
rect 12937 2117 12962 2138
rect 13002 2117 13006 2138
rect 13006 2117 13036 2138
rect 13076 2117 13109 2138
rect 13109 2117 13110 2138
rect 13150 2117 13178 2138
rect 13178 2117 13184 2138
rect 13224 2117 13247 2138
rect 13247 2117 13258 2138
rect 13298 2117 13316 2138
rect 13316 2117 13332 2138
rect 13372 2117 13385 2138
rect 13385 2117 13406 2138
rect 13446 2117 13454 2138
rect 13454 2117 13480 2138
rect 13520 2117 13523 2138
rect 13523 2117 13554 2138
rect 13594 2117 13627 2138
rect 13627 2117 13628 2138
rect 13668 2117 13696 2138
rect 13696 2117 13702 2138
rect 13741 2117 13765 2138
rect 13765 2117 13775 2138
rect 13814 2117 13834 2138
rect 13834 2117 13848 2138
rect 13887 2117 13903 2138
rect 13903 2117 13921 2138
rect 13960 2117 13972 2138
rect 13972 2117 13994 2138
rect 14033 2117 14041 2138
rect 14041 2117 14067 2138
rect 12632 2104 12666 2117
rect 12706 2104 12740 2117
rect 12780 2104 12814 2117
rect 12854 2104 12888 2117
rect 12928 2104 12962 2117
rect 13002 2104 13036 2117
rect 13076 2104 13110 2117
rect 13150 2104 13184 2117
rect 13224 2104 13258 2117
rect 13298 2104 13332 2117
rect 13372 2104 13406 2117
rect 13446 2104 13480 2117
rect 13520 2104 13554 2117
rect 13594 2104 13628 2117
rect 13668 2104 13702 2117
rect 13741 2104 13775 2117
rect 13814 2104 13848 2117
rect 13887 2104 13921 2117
rect 13960 2104 13994 2117
rect 14033 2104 14067 2117
rect 11448 2049 11476 2066
rect 11476 2049 11482 2066
rect 11522 2049 11546 2066
rect 11546 2049 11556 2066
rect 11596 2049 11616 2066
rect 11616 2049 11630 2066
rect 11670 2049 11686 2066
rect 11686 2049 11704 2066
rect 11744 2049 11756 2066
rect 11756 2049 11778 2066
rect 11818 2049 11826 2066
rect 11826 2049 11852 2066
rect 11892 2049 11896 2066
rect 11896 2049 11926 2066
rect 11966 2049 12000 2066
rect 12040 2049 12070 2066
rect 12070 2049 12074 2066
rect 12114 2049 12140 2066
rect 12140 2049 12148 2066
rect 12188 2049 12210 2066
rect 12210 2049 12222 2066
rect 12262 2049 12280 2066
rect 12280 2049 12296 2066
rect 12336 2049 12350 2066
rect 12350 2049 12370 2066
rect 12410 2049 12419 2066
rect 12419 2049 12444 2066
rect 12484 2049 12488 2066
rect 12488 2049 12518 2066
rect 11448 2032 11482 2049
rect 11522 2032 11556 2049
rect 11596 2032 11630 2049
rect 11670 2032 11704 2049
rect 11744 2032 11778 2049
rect 11818 2032 11852 2049
rect 11892 2032 11926 2049
rect 11966 2032 12000 2049
rect 12040 2032 12074 2049
rect 12114 2032 12148 2049
rect 12188 2032 12222 2049
rect 12262 2032 12296 2049
rect 12336 2032 12370 2049
rect 12410 2032 12444 2049
rect 12484 2032 12518 2049
rect 12558 2032 12592 2066
rect 12632 2049 12661 2066
rect 12661 2049 12666 2066
rect 12706 2049 12730 2066
rect 12730 2049 12740 2066
rect 12780 2049 12799 2066
rect 12799 2049 12814 2066
rect 12854 2049 12868 2066
rect 12868 2049 12888 2066
rect 12928 2049 12937 2066
rect 12937 2049 12962 2066
rect 13002 2049 13006 2066
rect 13006 2049 13036 2066
rect 13076 2049 13109 2066
rect 13109 2049 13110 2066
rect 13150 2049 13178 2066
rect 13178 2049 13184 2066
rect 13224 2049 13247 2066
rect 13247 2049 13258 2066
rect 13298 2049 13316 2066
rect 13316 2049 13332 2066
rect 13372 2049 13385 2066
rect 13385 2049 13406 2066
rect 13446 2049 13454 2066
rect 13454 2049 13480 2066
rect 13520 2049 13523 2066
rect 13523 2049 13554 2066
rect 13594 2049 13627 2066
rect 13627 2049 13628 2066
rect 13668 2049 13696 2066
rect 13696 2049 13702 2066
rect 13741 2049 13765 2066
rect 13765 2049 13775 2066
rect 13814 2049 13834 2066
rect 13834 2049 13848 2066
rect 13887 2049 13903 2066
rect 13903 2049 13921 2066
rect 13960 2049 13972 2066
rect 13972 2049 13994 2066
rect 14033 2049 14041 2066
rect 14041 2049 14067 2066
rect 12632 2032 12666 2049
rect 12706 2032 12740 2049
rect 12780 2032 12814 2049
rect 12854 2032 12888 2049
rect 12928 2032 12962 2049
rect 13002 2032 13036 2049
rect 13076 2032 13110 2049
rect 13150 2032 13184 2049
rect 13224 2032 13258 2049
rect 13298 2032 13332 2049
rect 13372 2032 13406 2049
rect 13446 2032 13480 2049
rect 13520 2032 13554 2049
rect 13594 2032 13628 2049
rect 13668 2032 13702 2049
rect 13741 2032 13775 2049
rect 13814 2032 13848 2049
rect 13887 2032 13921 2049
rect 13960 2032 13994 2049
rect 14033 2032 14067 2049
rect 11448 1981 11476 1994
rect 11476 1981 11482 1994
rect 11522 1981 11546 1994
rect 11546 1981 11556 1994
rect 11596 1981 11616 1994
rect 11616 1981 11630 1994
rect 11670 1981 11686 1994
rect 11686 1981 11704 1994
rect 11744 1981 11756 1994
rect 11756 1981 11778 1994
rect 11818 1981 11826 1994
rect 11826 1981 11852 1994
rect 11892 1981 11896 1994
rect 11896 1981 11926 1994
rect 11966 1981 12000 1994
rect 12040 1981 12070 1994
rect 12070 1981 12074 1994
rect 12114 1981 12140 1994
rect 12140 1981 12148 1994
rect 12188 1981 12210 1994
rect 12210 1981 12222 1994
rect 12262 1981 12280 1994
rect 12280 1981 12296 1994
rect 12336 1981 12350 1994
rect 12350 1981 12370 1994
rect 12410 1981 12419 1994
rect 12419 1981 12444 1994
rect 12484 1981 12488 1994
rect 12488 1981 12518 1994
rect 11448 1960 11482 1981
rect 11522 1960 11556 1981
rect 11596 1960 11630 1981
rect 11670 1960 11704 1981
rect 11744 1960 11778 1981
rect 11818 1960 11852 1981
rect 11892 1960 11926 1981
rect 11966 1960 12000 1981
rect 12040 1960 12074 1981
rect 12114 1960 12148 1981
rect 12188 1960 12222 1981
rect 12262 1960 12296 1981
rect 12336 1960 12370 1981
rect 12410 1960 12444 1981
rect 12484 1960 12518 1981
rect 12558 1960 12592 1994
rect 12632 1981 12661 1994
rect 12661 1981 12666 1994
rect 12706 1981 12730 1994
rect 12730 1981 12740 1994
rect 12780 1981 12799 1994
rect 12799 1981 12814 1994
rect 12854 1981 12868 1994
rect 12868 1981 12888 1994
rect 12928 1981 12937 1994
rect 12937 1981 12962 1994
rect 13002 1981 13006 1994
rect 13006 1981 13036 1994
rect 13076 1981 13109 1994
rect 13109 1981 13110 1994
rect 13150 1981 13178 1994
rect 13178 1981 13184 1994
rect 13224 1981 13247 1994
rect 13247 1981 13258 1994
rect 13298 1981 13316 1994
rect 13316 1981 13332 1994
rect 13372 1981 13385 1994
rect 13385 1981 13406 1994
rect 13446 1981 13454 1994
rect 13454 1981 13480 1994
rect 13520 1981 13523 1994
rect 13523 1981 13554 1994
rect 13594 1981 13627 1994
rect 13627 1981 13628 1994
rect 13668 1981 13696 1994
rect 13696 1981 13702 1994
rect 13741 1981 13765 1994
rect 13765 1981 13775 1994
rect 13814 1981 13834 1994
rect 13834 1981 13848 1994
rect 13887 1981 13903 1994
rect 13903 1981 13921 1994
rect 13960 1981 13972 1994
rect 13972 1981 13994 1994
rect 14033 1981 14041 1994
rect 14041 1981 14067 1994
rect 12632 1960 12666 1981
rect 12706 1960 12740 1981
rect 12780 1960 12814 1981
rect 12854 1960 12888 1981
rect 12928 1960 12962 1981
rect 13002 1960 13036 1981
rect 13076 1960 13110 1981
rect 13150 1960 13184 1981
rect 13224 1960 13258 1981
rect 13298 1960 13332 1981
rect 13372 1960 13406 1981
rect 13446 1960 13480 1981
rect 13520 1960 13554 1981
rect 13594 1960 13628 1981
rect 13668 1960 13702 1981
rect 13741 1960 13775 1981
rect 13814 1960 13848 1981
rect 13887 1960 13921 1981
rect 13960 1960 13994 1981
rect 14033 1960 14067 1981
rect 11448 1913 11476 1922
rect 11476 1913 11482 1922
rect 11522 1913 11546 1922
rect 11546 1913 11556 1922
rect 11596 1913 11616 1922
rect 11616 1913 11630 1922
rect 11670 1913 11686 1922
rect 11686 1913 11704 1922
rect 11744 1913 11756 1922
rect 11756 1913 11778 1922
rect 11818 1913 11826 1922
rect 11826 1913 11852 1922
rect 11892 1913 11896 1922
rect 11896 1913 11926 1922
rect 11966 1913 12000 1922
rect 12040 1913 12070 1922
rect 12070 1913 12074 1922
rect 12114 1913 12140 1922
rect 12140 1913 12148 1922
rect 12188 1913 12210 1922
rect 12210 1913 12222 1922
rect 12262 1913 12280 1922
rect 12280 1913 12296 1922
rect 12336 1913 12350 1922
rect 12350 1913 12370 1922
rect 12410 1913 12419 1922
rect 12419 1913 12444 1922
rect 12484 1913 12488 1922
rect 12488 1913 12518 1922
rect 11448 1888 11482 1913
rect 11522 1888 11556 1913
rect 11596 1888 11630 1913
rect 11670 1888 11704 1913
rect 11744 1888 11778 1913
rect 11818 1888 11852 1913
rect 11892 1888 11926 1913
rect 11966 1888 12000 1913
rect 12040 1888 12074 1913
rect 12114 1888 12148 1913
rect 12188 1888 12222 1913
rect 12262 1888 12296 1913
rect 12336 1888 12370 1913
rect 12410 1888 12444 1913
rect 12484 1888 12518 1913
rect 12558 1888 12592 1922
rect 12632 1913 12661 1922
rect 12661 1913 12666 1922
rect 12706 1913 12730 1922
rect 12730 1913 12740 1922
rect 12780 1913 12799 1922
rect 12799 1913 12814 1922
rect 12854 1913 12868 1922
rect 12868 1913 12888 1922
rect 12928 1913 12937 1922
rect 12937 1913 12962 1922
rect 13002 1913 13006 1922
rect 13006 1913 13036 1922
rect 13076 1913 13109 1922
rect 13109 1913 13110 1922
rect 13150 1913 13178 1922
rect 13178 1913 13184 1922
rect 13224 1913 13247 1922
rect 13247 1913 13258 1922
rect 13298 1913 13316 1922
rect 13316 1913 13332 1922
rect 13372 1913 13385 1922
rect 13385 1913 13406 1922
rect 13446 1913 13454 1922
rect 13454 1913 13480 1922
rect 13520 1913 13523 1922
rect 13523 1913 13554 1922
rect 13594 1913 13627 1922
rect 13627 1913 13628 1922
rect 13668 1913 13696 1922
rect 13696 1913 13702 1922
rect 13741 1913 13765 1922
rect 13765 1913 13775 1922
rect 13814 1913 13834 1922
rect 13834 1913 13848 1922
rect 13887 1913 13903 1922
rect 13903 1913 13921 1922
rect 13960 1913 13972 1922
rect 13972 1913 13994 1922
rect 14033 1913 14041 1922
rect 14041 1913 14067 1922
rect 12632 1888 12666 1913
rect 12706 1888 12740 1913
rect 12780 1888 12814 1913
rect 12854 1888 12888 1913
rect 12928 1888 12962 1913
rect 13002 1888 13036 1913
rect 13076 1888 13110 1913
rect 13150 1888 13184 1913
rect 13224 1888 13258 1913
rect 13298 1888 13332 1913
rect 13372 1888 13406 1913
rect 13446 1888 13480 1913
rect 13520 1888 13554 1913
rect 13594 1888 13628 1913
rect 13668 1888 13702 1913
rect 13741 1888 13775 1913
rect 13814 1888 13848 1913
rect 13887 1888 13921 1913
rect 13960 1888 13994 1913
rect 14033 1888 14067 1913
rect 11448 1845 11476 1850
rect 11476 1845 11482 1850
rect 11522 1845 11546 1850
rect 11546 1845 11556 1850
rect 11596 1845 11616 1850
rect 11616 1845 11630 1850
rect 11670 1845 11686 1850
rect 11686 1845 11704 1850
rect 11744 1845 11756 1850
rect 11756 1845 11778 1850
rect 11818 1845 11826 1850
rect 11826 1845 11852 1850
rect 11892 1845 11896 1850
rect 11896 1845 11926 1850
rect 11966 1845 12000 1850
rect 12040 1845 12070 1850
rect 12070 1845 12074 1850
rect 12114 1845 12140 1850
rect 12140 1845 12148 1850
rect 12188 1845 12210 1850
rect 12210 1845 12222 1850
rect 12262 1845 12280 1850
rect 12280 1845 12296 1850
rect 12336 1845 12350 1850
rect 12350 1845 12370 1850
rect 12410 1845 12419 1850
rect 12419 1845 12444 1850
rect 12484 1845 12488 1850
rect 12488 1845 12518 1850
rect 11448 1816 11482 1845
rect 11522 1816 11556 1845
rect 11596 1816 11630 1845
rect 11670 1816 11704 1845
rect 11744 1816 11778 1845
rect 11818 1816 11852 1845
rect 11892 1816 11926 1845
rect 11966 1816 12000 1845
rect 12040 1816 12074 1845
rect 12114 1816 12148 1845
rect 12188 1816 12222 1845
rect 12262 1816 12296 1845
rect 12336 1816 12370 1845
rect 12410 1816 12444 1845
rect 12484 1816 12518 1845
rect 12558 1816 12592 1850
rect 12632 1845 12661 1850
rect 12661 1845 12666 1850
rect 12706 1845 12730 1850
rect 12730 1845 12740 1850
rect 12780 1845 12799 1850
rect 12799 1845 12814 1850
rect 12854 1845 12868 1850
rect 12868 1845 12888 1850
rect 12928 1845 12937 1850
rect 12937 1845 12962 1850
rect 13002 1845 13006 1850
rect 13006 1845 13036 1850
rect 13076 1845 13109 1850
rect 13109 1845 13110 1850
rect 13150 1845 13178 1850
rect 13178 1845 13184 1850
rect 13224 1845 13247 1850
rect 13247 1845 13258 1850
rect 13298 1845 13316 1850
rect 13316 1845 13332 1850
rect 13372 1845 13385 1850
rect 13385 1845 13406 1850
rect 13446 1845 13454 1850
rect 13454 1845 13480 1850
rect 13520 1845 13523 1850
rect 13523 1845 13554 1850
rect 13594 1845 13627 1850
rect 13627 1845 13628 1850
rect 13668 1845 13696 1850
rect 13696 1845 13702 1850
rect 13741 1845 13765 1850
rect 13765 1845 13775 1850
rect 13814 1845 13834 1850
rect 13834 1845 13848 1850
rect 13887 1845 13903 1850
rect 13903 1845 13921 1850
rect 13960 1845 13972 1850
rect 13972 1845 13994 1850
rect 14033 1845 14041 1850
rect 14041 1845 14067 1850
rect 12632 1816 12666 1845
rect 12706 1816 12740 1845
rect 12780 1816 12814 1845
rect 12854 1816 12888 1845
rect 12928 1816 12962 1845
rect 13002 1816 13036 1845
rect 13076 1816 13110 1845
rect 13150 1816 13184 1845
rect 13224 1816 13258 1845
rect 13298 1816 13332 1845
rect 13372 1816 13406 1845
rect 13446 1816 13480 1845
rect 13520 1816 13554 1845
rect 13594 1816 13628 1845
rect 13668 1816 13702 1845
rect 13741 1816 13775 1845
rect 13814 1816 13848 1845
rect 13887 1816 13921 1845
rect 13960 1816 13994 1845
rect 14033 1816 14067 1845
rect 11448 1777 11476 1778
rect 11476 1777 11482 1778
rect 11522 1777 11546 1778
rect 11546 1777 11556 1778
rect 11596 1777 11616 1778
rect 11616 1777 11630 1778
rect 11670 1777 11686 1778
rect 11686 1777 11704 1778
rect 11744 1777 11756 1778
rect 11756 1777 11778 1778
rect 11818 1777 11826 1778
rect 11826 1777 11852 1778
rect 11892 1777 11896 1778
rect 11896 1777 11926 1778
rect 11966 1777 12000 1778
rect 12040 1777 12070 1778
rect 12070 1777 12074 1778
rect 12114 1777 12140 1778
rect 12140 1777 12148 1778
rect 12188 1777 12210 1778
rect 12210 1777 12222 1778
rect 12262 1777 12280 1778
rect 12280 1777 12296 1778
rect 12336 1777 12350 1778
rect 12350 1777 12370 1778
rect 12410 1777 12419 1778
rect 12419 1777 12444 1778
rect 12484 1777 12488 1778
rect 12488 1777 12518 1778
rect 11448 1744 11482 1777
rect 11522 1744 11556 1777
rect 11596 1744 11630 1777
rect 11670 1744 11704 1777
rect 11744 1744 11778 1777
rect 11818 1744 11852 1777
rect 11892 1744 11926 1777
rect 11966 1744 12000 1777
rect 12040 1744 12074 1777
rect 12114 1744 12148 1777
rect 12188 1744 12222 1777
rect 12262 1744 12296 1777
rect 12336 1744 12370 1777
rect 12410 1744 12444 1777
rect 12484 1744 12518 1777
rect 12558 1744 12592 1778
rect 12632 1777 12661 1778
rect 12661 1777 12666 1778
rect 12706 1777 12730 1778
rect 12730 1777 12740 1778
rect 12780 1777 12799 1778
rect 12799 1777 12814 1778
rect 12854 1777 12868 1778
rect 12868 1777 12888 1778
rect 12928 1777 12937 1778
rect 12937 1777 12962 1778
rect 13002 1777 13006 1778
rect 13006 1777 13036 1778
rect 13076 1777 13109 1778
rect 13109 1777 13110 1778
rect 13150 1777 13178 1778
rect 13178 1777 13184 1778
rect 13224 1777 13247 1778
rect 13247 1777 13258 1778
rect 13298 1777 13316 1778
rect 13316 1777 13332 1778
rect 13372 1777 13385 1778
rect 13385 1777 13406 1778
rect 13446 1777 13454 1778
rect 13454 1777 13480 1778
rect 13520 1777 13523 1778
rect 13523 1777 13554 1778
rect 13594 1777 13627 1778
rect 13627 1777 13628 1778
rect 13668 1777 13696 1778
rect 13696 1777 13702 1778
rect 13741 1777 13765 1778
rect 13765 1777 13775 1778
rect 13814 1777 13834 1778
rect 13834 1777 13848 1778
rect 13887 1777 13903 1778
rect 13903 1777 13921 1778
rect 13960 1777 13972 1778
rect 13972 1777 13994 1778
rect 14033 1777 14041 1778
rect 14041 1777 14067 1778
rect 12632 1744 12666 1777
rect 12706 1744 12740 1777
rect 12780 1744 12814 1777
rect 12854 1744 12888 1777
rect 12928 1744 12962 1777
rect 13002 1744 13036 1777
rect 13076 1744 13110 1777
rect 13150 1744 13184 1777
rect 13224 1744 13258 1777
rect 13298 1744 13332 1777
rect 13372 1744 13406 1777
rect 13446 1744 13480 1777
rect 13520 1744 13554 1777
rect 13594 1744 13628 1777
rect 13668 1744 13702 1777
rect 13741 1744 13775 1777
rect 13814 1744 13848 1777
rect 13887 1744 13921 1777
rect 13960 1744 13994 1777
rect 14033 1744 14067 1777
<< metal1 >>
rect 62 6467 4320 6473
rect 62 6433 74 6467
rect 108 6433 146 6467
rect 180 6433 218 6467
rect 252 6433 290 6467
rect 324 6433 362 6467
rect 396 6433 434 6467
rect 468 6433 506 6467
rect 540 6433 578 6467
rect 612 6433 650 6467
rect 684 6433 722 6467
rect 756 6433 794 6467
rect 828 6433 866 6467
rect 900 6433 938 6467
rect 972 6433 1010 6467
rect 1044 6433 1082 6467
rect 1116 6433 1154 6467
rect 1188 6433 1226 6467
rect 1260 6433 1298 6467
rect 1332 6433 1370 6467
rect 1404 6433 1442 6467
rect 1476 6433 1514 6467
rect 1548 6433 1586 6467
rect 1620 6433 1658 6467
rect 1692 6433 1730 6467
rect 1764 6433 1802 6467
rect 1836 6433 1874 6467
rect 1908 6433 1946 6467
rect 1980 6433 2018 6467
rect 2052 6433 2090 6467
rect 2124 6433 2162 6467
rect 2196 6433 2234 6467
rect 2268 6433 2306 6467
rect 2340 6433 2378 6467
rect 2412 6433 2450 6467
rect 2484 6433 2522 6467
rect 2556 6433 2594 6467
rect 2628 6433 2666 6467
rect 2700 6433 2738 6467
rect 2772 6433 2810 6467
rect 2844 6433 2882 6467
rect 2916 6433 2954 6467
rect 2988 6433 3026 6467
rect 3060 6433 3098 6467
rect 3132 6433 3170 6467
rect 3204 6433 3242 6467
rect 3276 6433 3314 6467
rect 3348 6433 3386 6467
rect 3420 6433 3458 6467
rect 3492 6433 3530 6467
rect 3564 6433 3602 6467
rect 3636 6433 3674 6467
rect 3708 6433 3746 6467
rect 3780 6433 3818 6467
rect 3852 6433 3890 6467
rect 3924 6433 3962 6467
rect 3996 6433 4034 6467
rect 4068 6433 4106 6467
rect 4140 6433 4178 6467
rect 4212 6433 4250 6467
rect 4284 6433 4320 6467
rect 62 6427 4320 6433
rect 62 6412 118 6427
tri 118 6412 133 6427 nw
tri 4308 6421 4314 6427 ne
rect 4314 6421 4320 6427
rect 4372 6421 4385 6473
rect 4437 6421 4450 6473
rect 4502 6421 4516 6473
rect 4568 6467 7589 6473
rect 4572 6433 4610 6467
rect 4644 6433 4682 6467
rect 4716 6433 4754 6467
rect 4788 6433 4826 6467
rect 4860 6433 4898 6467
rect 4932 6433 4971 6467
rect 5005 6433 5044 6467
rect 5078 6433 5117 6467
rect 5151 6433 5190 6467
rect 5224 6433 5263 6467
rect 5297 6433 5336 6467
rect 5370 6433 5409 6467
rect 5443 6433 5482 6467
rect 5516 6433 5555 6467
rect 5589 6433 5628 6467
rect 5662 6433 5701 6467
rect 5735 6433 5774 6467
rect 5808 6433 5847 6467
rect 5881 6433 5920 6467
rect 5954 6433 5993 6467
rect 6027 6433 6066 6467
rect 6100 6433 6139 6467
rect 6173 6433 6212 6467
rect 6246 6433 6285 6467
rect 6319 6433 6358 6467
rect 6392 6433 6431 6467
rect 6465 6433 6504 6467
rect 6538 6433 6577 6467
rect 6611 6433 6650 6467
rect 6684 6433 6723 6467
rect 6757 6433 6796 6467
rect 6830 6433 6869 6467
rect 6903 6433 6942 6467
rect 6976 6433 7015 6467
rect 7049 6433 7088 6467
rect 7122 6433 7161 6467
rect 7195 6433 7234 6467
rect 7268 6433 7307 6467
rect 7341 6433 7380 6467
rect 7414 6433 7453 6467
rect 7487 6433 7526 6467
rect 7560 6433 7589 6467
rect 4568 6427 7589 6433
rect 4568 6421 4574 6427
tri 4574 6421 4580 6427 nw
tri 7577 6421 7583 6427 ne
rect 7583 6421 7589 6427
rect 7641 6421 7653 6473
rect 7705 6467 7717 6473
rect 7769 6467 13536 6473
rect 7706 6433 7717 6467
rect 7779 6433 7818 6467
rect 7852 6433 7891 6467
rect 7925 6433 7964 6467
rect 7998 6433 8037 6467
rect 8071 6433 8110 6467
rect 8144 6433 8183 6467
rect 8217 6433 8256 6467
rect 8290 6433 8329 6467
rect 8363 6433 8402 6467
rect 8436 6433 8475 6467
rect 8509 6433 8548 6467
rect 8582 6433 8621 6467
rect 8655 6433 8694 6467
rect 8728 6433 8767 6467
rect 8801 6433 8840 6467
rect 8874 6433 8913 6467
rect 8947 6433 8986 6467
rect 9020 6433 9059 6467
rect 9093 6433 9132 6467
rect 9166 6433 9205 6467
rect 9239 6433 9278 6467
rect 9312 6433 9351 6467
rect 9385 6433 9424 6467
rect 9458 6433 9497 6467
rect 9531 6433 9570 6467
rect 9604 6433 9643 6467
rect 9677 6433 9693 6467
rect 9750 6433 9757 6467
rect 9896 6433 13536 6467
rect 7705 6421 7717 6433
rect 7769 6427 9693 6433
rect 7769 6421 7775 6427
tri 7775 6421 7781 6427 nw
tri 9418 6421 9424 6427 ne
rect 9424 6421 9693 6427
tri 9424 6412 9433 6421 ne
rect 9433 6415 9693 6421
rect 9745 6415 9757 6433
rect 9809 6415 9821 6433
rect 9873 6415 13536 6433
rect 9433 6412 13536 6415
rect 62 6395 108 6412
tri 108 6402 118 6412 nw
tri 9433 6402 9443 6412 ne
rect 9443 6402 10510 6412
rect 62 6361 68 6395
rect 102 6361 108 6395
tri 9443 6387 9458 6402 ne
rect 9458 6401 10510 6402
rect 9458 6387 9693 6401
tri 905 6378 914 6387 se
rect 914 6378 9401 6387
tri 9401 6378 9410 6387 sw
tri 9458 6378 9467 6387 ne
rect 9467 6378 9693 6387
tri 901 6374 905 6378 se
rect 905 6374 9410 6378
tri 9410 6374 9414 6378 sw
tri 9467 6374 9471 6378 ne
rect 9471 6374 9693 6378
rect 62 6323 108 6361
tri 867 6340 901 6374 se
rect 901 6357 9414 6374
tri 9414 6357 9431 6374 sw
tri 9471 6357 9488 6374 ne
rect 9488 6357 9693 6374
rect 901 6340 9431 6357
tri 9431 6340 9448 6357 sw
tri 9488 6340 9505 6357 ne
rect 9505 6349 9693 6357
rect 9745 6349 9757 6401
rect 9809 6349 9821 6401
rect 9873 6378 10510 6401
rect 10544 6378 10584 6412
rect 10618 6378 10658 6412
rect 10692 6378 10732 6412
rect 10766 6378 10806 6412
rect 10840 6378 10880 6412
rect 10914 6378 10954 6412
rect 10988 6378 11028 6412
rect 11062 6378 11102 6412
rect 11136 6378 11176 6412
rect 11210 6378 11250 6412
rect 11284 6378 11324 6412
rect 11358 6378 11398 6412
rect 11432 6378 11472 6412
rect 11506 6378 11546 6412
rect 11580 6378 11620 6412
rect 11654 6378 11694 6412
rect 11728 6378 11768 6412
rect 11802 6378 11842 6412
rect 11876 6378 11916 6412
rect 11950 6378 11990 6412
rect 12024 6378 12064 6412
rect 12098 6378 12138 6412
rect 12172 6378 12212 6412
rect 12246 6378 12286 6412
rect 12320 6378 12360 6412
rect 12394 6378 12434 6412
rect 12468 6378 12508 6412
rect 12542 6378 12581 6412
rect 12615 6378 12654 6412
rect 12688 6378 12727 6412
rect 12761 6378 12800 6412
rect 12834 6378 12873 6412
rect 12907 6378 12946 6412
rect 12980 6378 13019 6412
rect 13053 6378 13092 6412
rect 13126 6378 13165 6412
rect 13199 6378 13238 6412
rect 13272 6378 13311 6412
rect 13345 6378 13384 6412
rect 13418 6378 13536 6412
rect 9873 6374 13536 6378
rect 9873 6372 13496 6374
rect 9873 6349 9971 6372
rect 9505 6340 9971 6349
tri 9971 6340 10003 6372 nw
tri 13401 6344 13429 6372 ne
rect 13429 6344 13496 6372
tri 865 6338 867 6340 se
rect 867 6338 9448 6340
tri 9448 6338 9450 6340 sw
tri 9505 6338 9507 6340 ne
rect 9507 6338 9969 6340
tri 9969 6338 9971 6340 nw
rect 11034 6338 11164 6344
tri 13429 6340 13433 6344 ne
rect 13433 6340 13496 6344
rect 13530 6340 13536 6374
rect 62 6289 68 6323
rect 102 6289 108 6323
rect 62 6251 108 6289
rect 62 6217 68 6251
rect 102 6217 108 6251
rect 62 6179 108 6217
rect 62 6145 68 6179
rect 102 6145 108 6179
rect 62 6107 108 6145
rect 62 6073 68 6107
rect 102 6073 108 6107
tri 858 6331 865 6338 se
rect 865 6335 9450 6338
rect 865 6331 931 6335
tri 931 6331 935 6335 nw
tri 1689 6331 1693 6335 ne
rect 1693 6331 1766 6335
rect 62 6035 108 6073
rect 62 6001 68 6035
rect 102 6001 108 6035
rect 62 5963 108 6001
rect 62 5929 68 5963
rect 102 5929 108 5963
rect 62 5891 108 5929
rect 62 5857 68 5891
rect 102 5857 108 5891
rect 62 5819 108 5857
rect 62 5785 68 5819
rect 102 5785 108 5819
rect 62 5747 108 5785
rect 62 5713 68 5747
rect 102 5713 108 5747
rect 62 5675 108 5713
rect 62 5641 68 5675
rect 102 5641 108 5675
rect 62 5603 108 5641
rect 62 5569 68 5603
rect 102 5569 108 5603
rect 62 5531 108 5569
rect 62 5497 68 5531
rect 102 5497 108 5531
rect 62 5459 108 5497
rect 62 5425 68 5459
rect 102 5425 108 5459
rect 62 5387 108 5425
rect 62 5353 68 5387
rect 102 5353 108 5387
rect 62 5315 108 5353
rect 62 5281 68 5315
rect 102 5281 108 5315
rect 62 5243 108 5281
rect 62 5209 68 5243
rect 102 5209 108 5243
rect 62 5171 108 5209
rect 62 5137 68 5171
rect 102 5137 108 5171
rect 62 5099 108 5137
rect 62 5065 68 5099
rect 102 5065 108 5099
rect 62 5027 108 5065
rect 62 4993 68 5027
rect 102 4993 108 5027
rect 62 4955 108 4993
rect 62 4921 68 4955
rect 102 4921 108 4955
rect 62 4882 108 4921
rect 62 4848 68 4882
rect 102 4848 108 4882
rect 62 4809 108 4848
rect 62 4775 68 4809
rect 102 4775 108 4809
rect 62 4736 108 4775
rect 62 4702 68 4736
rect 102 4702 108 4736
rect 62 4663 108 4702
rect 62 4629 68 4663
rect 102 4629 108 4663
rect 62 4590 108 4629
rect 62 4556 68 4590
rect 102 4556 108 4590
rect 62 4517 108 4556
rect 62 4483 68 4517
rect 102 4483 108 4517
rect 62 4444 108 4483
rect 62 4410 68 4444
rect 102 4410 108 4444
rect 62 4371 108 4410
rect 62 4337 68 4371
rect 102 4337 108 4371
rect 62 4298 108 4337
rect 62 4264 68 4298
rect 102 4264 108 4298
rect 62 4225 108 4264
rect 62 4191 68 4225
rect 102 4191 108 4225
rect 62 4152 108 4191
rect 62 4118 68 4152
rect 102 4118 108 4152
rect 62 4079 108 4118
rect 62 4045 68 4079
rect 102 4045 108 4079
rect 62 4006 108 4045
rect 62 3972 68 4006
rect 102 3972 108 4006
rect 62 3933 108 3972
rect 62 3899 68 3933
rect 102 3899 108 3933
rect 62 3860 108 3899
rect 62 3826 68 3860
rect 102 3826 108 3860
rect 62 3787 108 3826
rect 62 3753 68 3787
rect 102 3753 108 3787
rect 62 3714 108 3753
rect 62 3680 68 3714
rect 102 3680 108 3714
rect 62 3641 108 3680
rect 62 3607 68 3641
rect 102 3607 108 3641
rect 62 3568 108 3607
rect 62 3534 68 3568
rect 102 3534 108 3568
rect 62 3495 108 3534
tri 42 3461 62 3481 se
rect 62 3461 68 3495
rect 102 3461 108 3495
rect 317 6100 830 6106
rect 317 6094 395 6100
rect 317 6060 323 6094
rect 357 6066 395 6094
rect 429 6066 473 6100
rect 507 6066 551 6100
rect 585 6066 629 6100
rect 663 6066 707 6100
rect 741 6066 784 6100
rect 818 6066 830 6100
rect 357 6060 830 6066
rect 317 6039 809 6060
tri 809 6039 830 6060 nw
rect 317 6022 760 6039
rect 317 5988 323 6022
rect 357 5990 760 6022
tri 760 5990 809 6039 nw
tri 809 5990 858 6039 se
rect 858 5990 910 6331
tri 910 6310 931 6331 nw
tri 1693 6310 1714 6331 ne
rect 938 6100 1376 6106
rect 1428 6100 1458 6106
rect 1510 6100 1540 6106
rect 1592 6100 1622 6106
rect 938 6066 950 6100
rect 984 6066 1027 6100
rect 1061 6066 1104 6100
rect 1138 6066 1181 6100
rect 1215 6066 1258 6100
rect 1292 6066 1335 6100
rect 1369 6066 1376 6100
rect 1446 6066 1458 6100
rect 1522 6066 1540 6100
rect 1598 6066 1622 6100
rect 938 6060 1376 6066
tri 938 6039 959 6060 ne
rect 959 6054 1376 6060
rect 1428 6054 1458 6066
rect 1510 6054 1540 6066
rect 1592 6054 1622 6066
rect 1674 6060 1686 6106
rect 1674 6054 1680 6060
tri 1680 6054 1686 6060 nw
rect 959 6039 1665 6054
tri 1665 6039 1680 6054 nw
tri 910 5990 959 6039 sw
tri 959 5990 1008 6039 ne
rect 1008 5990 1616 6039
tri 1616 5990 1665 6039 nw
tri 1665 5990 1714 6039 se
rect 1714 5990 1766 6331
tri 1766 6310 1791 6335 nw
tri 9323 6310 9348 6335 ne
rect 9348 6310 9450 6335
tri 9348 6307 9351 6310 ne
rect 9351 6307 9450 6310
tri 2600 6277 2630 6307 se
rect 2630 6277 8878 6307
tri 8878 6277 8908 6307 sw
tri 9351 6277 9381 6307 ne
rect 9381 6300 9450 6307
tri 9450 6300 9488 6338 sw
tri 9507 6300 9545 6338 ne
rect 9545 6335 9908 6338
rect 9545 6300 9693 6335
rect 9381 6277 9488 6300
tri 9488 6277 9511 6300 sw
tri 9545 6277 9568 6300 ne
rect 9568 6283 9693 6300
rect 9745 6283 9757 6335
rect 9809 6283 9821 6335
rect 9873 6283 9908 6335
rect 9568 6277 9908 6283
tri 9908 6277 9969 6338 nw
tri 11009 6283 11034 6308 se
rect 11034 6283 11046 6338
rect 11152 6300 11164 6338
tri 13433 6308 13465 6340 ne
rect 13465 6308 13536 6340
tri 11164 6300 11172 6308 sw
tri 13465 6300 13473 6308 ne
rect 13473 6300 13536 6308
rect 11152 6283 11172 6300
tri 11172 6283 11189 6300 sw
tri 13473 6288 13485 6300 ne
rect 13485 6288 13496 6300
tri 2570 6247 2600 6277 se
rect 2600 6255 8908 6277
rect 2600 6247 2644 6255
tri 2644 6247 2652 6255 nw
tri 8802 6247 8810 6255 ne
rect 8810 6247 8908 6255
rect 2570 6243 2640 6247
tri 2640 6243 2644 6247 nw
tri 8810 6243 8814 6247 ne
rect 8814 6243 8908 6247
tri 8908 6243 8942 6277 sw
tri 9381 6243 9415 6277 ne
rect 9415 6243 9511 6277
tri 9511 6243 9545 6277 sw
rect 2570 6232 2629 6243
tri 2629 6232 2640 6243 nw
tri 8814 6232 8825 6243 ne
rect 8825 6232 8942 6243
tri 8942 6232 8953 6243 sw
tri 9415 6232 9426 6243 ne
rect 9426 6232 9545 6243
tri 9545 6232 9556 6243 sw
rect 1794 6100 2542 6106
rect 1794 6066 1806 6100
rect 1840 6066 1883 6100
rect 1917 6066 1960 6100
rect 1994 6066 2037 6100
rect 2071 6066 2114 6100
rect 2148 6066 2191 6100
rect 2225 6066 2268 6100
rect 2302 6066 2344 6100
rect 2378 6066 2420 6100
rect 2454 6066 2496 6100
rect 2530 6066 2542 6100
rect 1794 6060 2542 6066
tri 1794 6039 1815 6060 ne
rect 1815 6039 2521 6060
tri 2521 6039 2542 6060 nw
tri 1766 5990 1815 6039 sw
tri 1815 5990 1864 6039 ne
rect 1864 5990 2472 6039
tri 2472 5990 2521 6039 nw
tri 2521 5990 2570 6039 se
rect 2570 5990 2622 6232
tri 2622 6225 2629 6232 nw
tri 8825 6227 8830 6232 ne
rect 8830 6227 8953 6232
tri 8953 6227 8958 6232 sw
tri 9426 6227 9431 6232 ne
rect 9431 6227 9556 6232
tri 9556 6227 9561 6232 sw
rect 10220 6231 10226 6283
rect 10278 6231 10290 6283
rect 10342 6277 10825 6283
rect 10342 6243 10707 6277
rect 10741 6243 10779 6277
rect 10813 6243 10825 6277
rect 10342 6231 10825 6243
rect 10962 6231 10968 6283
rect 11020 6231 11032 6283
rect 11152 6277 13015 6283
rect 11152 6243 11979 6277
rect 12013 6243 12051 6277
rect 12085 6243 12580 6277
rect 12614 6243 12652 6277
rect 12686 6243 12897 6277
rect 11152 6232 12897 6243
rect 11084 6231 12897 6232
tri 3480 6225 3482 6227 se
rect 3482 6225 8668 6227
tri 3447 6192 3480 6225 se
rect 3480 6192 8668 6225
tri 3426 6171 3447 6192 se
rect 3447 6175 8668 6192
rect 8720 6175 8732 6227
rect 8784 6175 8790 6227
rect 8830 6175 8836 6227
rect 8888 6175 8900 6227
rect 8952 6175 8958 6227
rect 9431 6175 9437 6227
rect 9489 6175 9503 6227
rect 9555 6175 9561 6227
tri 11029 6226 11034 6231 ne
rect 11034 6226 12897 6231
tri 12824 6198 12852 6226 ne
rect 12852 6198 12897 6226
tri 9717 6192 9723 6198 se
rect 9723 6192 11408 6198
tri 9700 6175 9717 6192 se
rect 9717 6175 11290 6192
rect 3447 6171 3499 6175
tri 3499 6171 3503 6175 nw
tri 4257 6171 4261 6175 ne
rect 4261 6171 4342 6175
rect 3426 6158 3486 6171
tri 3486 6158 3499 6171 nw
tri 4261 6158 4274 6171 ne
rect 4274 6158 4342 6171
tri 4342 6158 4359 6175 nw
tri 9683 6158 9700 6175 se
rect 9700 6158 11290 6175
rect 11324 6158 11362 6192
rect 11396 6158 11408 6192
tri 12852 6171 12879 6198 ne
rect 12879 6171 12897 6198
rect 13003 6171 13015 6277
rect 13088 6280 13112 6288
rect 13164 6280 13180 6288
rect 13088 6246 13100 6280
rect 13164 6246 13172 6280
rect 13088 6236 13112 6246
rect 13164 6236 13180 6246
rect 13232 6236 13238 6288
tri 13485 6283 13490 6288 ne
rect 13490 6266 13496 6288
rect 13530 6266 13536 6300
rect 13490 6226 13536 6266
tri 13485 6192 13490 6197 se
rect 13490 6192 13496 6226
rect 13530 6192 13536 6226
tri 12879 6165 12885 6171 ne
rect 12885 6165 13015 6171
tri 13458 6165 13485 6192 se
rect 13485 6165 13536 6192
rect 3426 6152 3480 6158
tri 3480 6152 3486 6158 nw
tri 4274 6152 4280 6158 ne
rect 4280 6152 4336 6158
tri 4336 6152 4342 6158 nw
tri 9678 6153 9683 6158 se
rect 9683 6153 11408 6158
tri 8985 6152 8986 6153 se
rect 8986 6152 8992 6153
rect 2650 6100 3398 6106
rect 2650 6066 2662 6100
rect 2696 6066 2739 6100
rect 2773 6066 2816 6100
rect 2850 6066 2893 6100
rect 2927 6066 2970 6100
rect 3004 6066 3047 6100
rect 3081 6066 3124 6100
rect 3158 6066 3200 6100
rect 3234 6066 3276 6100
rect 3310 6066 3352 6100
rect 3386 6066 3398 6100
rect 2650 6060 3398 6066
tri 2650 6039 2671 6060 ne
rect 2671 6039 3377 6060
tri 3377 6039 3398 6060 nw
tri 2622 5990 2671 6039 sw
tri 2671 5990 2720 6039 ne
rect 2720 5990 3328 6039
tri 3328 5990 3377 6039 nw
tri 3377 5990 3426 6039 se
rect 3426 5990 3478 6152
tri 3478 6150 3480 6152 nw
tri 4280 6150 4282 6152 ne
rect 3506 6100 4249 6106
rect 3506 6066 3518 6100
rect 3552 6066 3595 6100
rect 3629 6066 3671 6100
rect 3705 6066 3747 6100
rect 3781 6066 3823 6100
rect 3857 6066 3899 6100
rect 3933 6066 3975 6100
rect 4009 6066 4051 6100
rect 4085 6066 4127 6100
rect 4161 6066 4203 6100
rect 4237 6066 4249 6100
rect 3506 6060 4249 6066
tri 3506 6039 3527 6060 ne
rect 3527 6039 4228 6060
tri 4228 6039 4249 6060 nw
tri 3478 5990 3527 6039 sw
tri 3527 5990 3576 6039 ne
rect 3576 5990 4174 6039
rect 357 5988 733 5990
rect 317 5963 733 5988
tri 733 5963 760 5990 nw
tri 782 5963 809 5990 se
rect 809 5963 959 5990
tri 959 5963 986 5990 sw
tri 1008 5963 1035 5990 ne
rect 1035 5963 1589 5990
tri 1589 5963 1616 5990 nw
tri 1638 5963 1665 5990 se
rect 1665 5963 1815 5990
tri 1815 5963 1842 5990 sw
tri 1864 5963 1891 5990 ne
rect 1891 5963 2445 5990
tri 2445 5963 2472 5990 nw
tri 2494 5963 2521 5990 se
rect 2521 5963 2671 5990
tri 2671 5963 2698 5990 sw
tri 2720 5963 2747 5990 ne
rect 2747 5963 3301 5990
tri 3301 5963 3328 5990 nw
tri 3350 5963 3377 5990 se
rect 3377 5963 3527 5990
tri 3527 5963 3554 5990 sw
tri 3576 5963 3603 5990 ne
rect 3603 5985 4174 5990
tri 4174 5985 4228 6039 nw
tri 4228 5985 4282 6039 se
rect 4282 5985 4334 6152
tri 4334 6150 4336 6152 nw
tri 8983 6150 8985 6152 se
rect 8985 6150 8992 6152
tri 8980 6147 8983 6150 se
rect 8983 6147 8992 6150
tri 7901 6141 7907 6147 se
rect 7907 6141 7913 6147
tri 7867 6107 7901 6141 se
rect 7901 6107 7913 6141
tri 7866 6106 7867 6107 se
rect 7867 6106 7913 6107
rect 4367 6100 7913 6106
rect 4367 6066 4379 6100
rect 4413 6066 4455 6100
rect 4489 6066 4531 6100
rect 4565 6066 4607 6100
rect 4641 6066 4683 6100
rect 4717 6066 4757 6100
rect 4367 6060 4757 6066
tri 4367 6039 4388 6060 ne
rect 4388 6048 4757 6060
rect 4809 6048 4821 6100
rect 4873 6094 4885 6100
rect 4937 6066 4987 6100
rect 5021 6066 5061 6100
rect 5095 6066 5135 6100
rect 5169 6066 5209 6100
rect 5243 6066 5283 6100
rect 5317 6066 5357 6100
rect 5391 6066 5431 6100
rect 5465 6066 5505 6100
rect 5539 6066 5579 6100
rect 5613 6066 5652 6100
rect 5686 6066 5725 6100
rect 5759 6066 5798 6100
rect 5832 6066 5871 6100
rect 5905 6066 5944 6100
rect 5978 6066 6017 6100
rect 6051 6066 6090 6100
rect 6124 6066 6163 6100
rect 6197 6066 6236 6100
rect 6270 6066 6309 6100
rect 6343 6066 6382 6100
rect 6416 6066 6455 6100
rect 6489 6066 6528 6100
rect 6562 6066 6601 6100
rect 6635 6066 6674 6100
rect 6708 6066 6747 6100
rect 6781 6066 6820 6100
rect 6854 6066 6893 6100
rect 6927 6066 6966 6100
rect 7000 6066 7039 6100
rect 7073 6066 7112 6100
rect 7146 6066 7185 6100
rect 7219 6066 7258 6100
rect 7292 6066 7331 6100
rect 7365 6095 7913 6100
rect 7965 6095 7979 6147
rect 8031 6141 8045 6147
rect 8097 6141 8111 6147
rect 8163 6141 8992 6147
rect 9044 6141 9056 6153
rect 9108 6141 9121 6153
rect 9173 6141 9186 6153
rect 9238 6152 9244 6153
tri 9244 6152 9245 6153 sw
tri 9677 6152 9678 6153 se
rect 9678 6152 11408 6153
tri 13445 6152 13458 6165 se
rect 13458 6152 13536 6165
rect 9238 6147 9245 6152
tri 9245 6147 9250 6152 sw
tri 9672 6147 9677 6152 se
rect 9677 6147 9723 6152
rect 9238 6141 9585 6147
rect 8032 6107 8045 6141
rect 8105 6107 8111 6141
rect 8178 6107 8217 6141
rect 8251 6107 8290 6141
rect 8324 6107 8363 6141
rect 8397 6107 8436 6141
rect 8470 6107 8509 6141
rect 8543 6107 8582 6141
rect 8616 6107 8655 6141
rect 8689 6107 8728 6141
rect 8762 6107 8801 6141
rect 8835 6107 8874 6141
rect 8908 6107 8947 6141
rect 8981 6107 8992 6141
rect 9055 6107 9056 6141
rect 9238 6107 9243 6141
rect 9277 6107 9317 6141
rect 9351 6107 9391 6141
rect 9425 6107 9465 6141
rect 9499 6107 9539 6141
rect 9573 6107 9585 6141
tri 9657 6132 9672 6147 se
rect 9672 6132 9723 6147
tri 9723 6132 9743 6152 nw
tri 13425 6132 13445 6152 se
rect 13445 6132 13496 6152
tri 9643 6118 9657 6132 se
rect 9657 6118 9709 6132
tri 9709 6118 9723 6132 nw
tri 13411 6118 13425 6132 se
rect 13425 6118 13496 6132
rect 13530 6118 13536 6152
rect 8031 6095 8045 6107
rect 8097 6095 8111 6107
rect 8163 6101 8992 6107
rect 9044 6101 9056 6107
rect 9108 6101 9121 6107
rect 9173 6101 9186 6107
rect 9238 6101 9585 6107
tri 9626 6101 9643 6118 se
rect 9643 6101 9687 6118
rect 8163 6096 8170 6101
tri 8170 6096 8175 6101 nw
tri 9621 6096 9626 6101 se
rect 9626 6096 9687 6101
tri 9687 6096 9709 6118 nw
tri 13401 6108 13411 6118 se
rect 13411 6108 13536 6118
rect 9757 6096 13536 6108
rect 8163 6095 8169 6096
tri 8169 6095 8170 6096 nw
tri 9620 6095 9621 6096 se
rect 9621 6095 9679 6096
rect 7365 6094 7977 6095
rect 7365 6066 7403 6094
rect 4937 6060 7403 6066
rect 7437 6088 7977 6094
tri 7977 6088 7984 6095 nw
tri 9613 6088 9620 6095 se
rect 9620 6088 9679 6095
tri 9679 6088 9687 6096 nw
rect 9757 6088 10870 6096
rect 7437 6075 7959 6088
rect 7437 6060 7907 6075
tri 7959 6070 7977 6088 nw
tri 9598 6073 9613 6088 se
rect 9613 6073 9658 6088
rect 4388 6039 4831 6048
tri 4334 5985 4388 6039 sw
tri 4388 5985 4442 6039 ne
rect 4442 6035 4831 6039
rect 4442 5985 4757 6035
rect 3603 5973 4162 5985
tri 4162 5973 4174 5985 nw
tri 4216 5973 4228 5985 se
rect 4228 5973 4388 5985
tri 4388 5973 4400 5985 sw
tri 4442 5973 4454 5985 ne
rect 4454 5983 4757 5985
rect 4809 5983 4821 6035
rect 4454 5973 4831 5983
rect 3603 5963 4108 5973
rect 317 5950 684 5963
rect 317 5916 323 5950
rect 357 5916 684 5950
rect 317 5914 684 5916
tri 684 5914 733 5963 nw
tri 733 5914 782 5963 se
rect 782 5914 986 5963
tri 986 5914 1035 5963 sw
tri 1035 5914 1084 5963 ne
rect 1084 5914 1540 5963
tri 1540 5914 1589 5963 nw
tri 1589 5914 1638 5963 se
rect 1638 5914 1842 5963
tri 1842 5914 1891 5963 sw
tri 1891 5914 1940 5963 ne
rect 1940 5914 2396 5963
tri 2396 5914 2445 5963 nw
tri 2445 5914 2494 5963 se
rect 2494 5914 2698 5963
tri 2698 5914 2747 5963 sw
tri 2747 5914 2796 5963 ne
rect 2796 5914 3252 5963
tri 3252 5914 3301 5963 nw
tri 3301 5914 3350 5963 se
rect 3350 5914 3554 5963
tri 3554 5914 3603 5963 sw
tri 3603 5914 3652 5963 ne
rect 3652 5919 4108 5963
tri 4108 5919 4162 5973 nw
tri 4162 5919 4216 5973 se
rect 4216 5919 4400 5973
tri 4400 5919 4454 5973 sw
tri 4454 5919 4508 5973 ne
rect 4508 5970 4831 5973
rect 4508 5919 4757 5970
rect 3652 5914 4080 5919
rect 317 5878 656 5914
tri 656 5886 684 5914 nw
tri 705 5886 733 5914 se
rect 733 5886 1035 5914
rect 317 5844 323 5878
rect 357 5844 656 5878
rect 317 5806 656 5844
rect 317 5772 323 5806
rect 357 5772 656 5806
rect 317 5734 656 5772
rect 317 5700 323 5734
rect 357 5731 656 5734
rect 357 5700 439 5731
rect 317 5697 439 5700
rect 473 5697 656 5731
rect 317 5662 656 5697
rect 317 5628 323 5662
rect 357 5658 656 5662
rect 357 5628 439 5658
rect 317 5624 439 5628
rect 473 5624 656 5658
rect 317 5590 656 5624
rect 317 5556 323 5590
rect 357 5585 656 5590
rect 357 5556 439 5585
rect 317 5551 439 5556
rect 473 5551 656 5585
rect 317 5518 656 5551
rect 317 5484 323 5518
rect 357 5512 656 5518
rect 357 5484 439 5512
rect 317 5478 439 5484
rect 473 5478 656 5512
rect 317 5446 656 5478
rect 317 5412 323 5446
rect 357 5439 656 5446
rect 357 5412 439 5439
rect 317 5405 439 5412
rect 473 5405 656 5439
rect 317 5374 656 5405
rect 317 5340 323 5374
rect 357 5366 656 5374
rect 357 5340 439 5366
rect 317 5332 439 5340
rect 473 5332 656 5366
rect 317 5302 656 5332
rect 317 5268 323 5302
rect 357 5293 656 5302
rect 357 5268 439 5293
rect 317 5259 439 5268
rect 473 5259 656 5293
rect 317 5230 656 5259
rect 317 5196 323 5230
rect 357 5220 656 5230
rect 357 5196 439 5220
rect 317 5186 439 5196
rect 473 5186 656 5220
rect 317 5158 656 5186
rect 317 5124 323 5158
rect 357 5147 656 5158
rect 357 5124 439 5147
rect 317 5113 439 5124
rect 473 5113 656 5147
rect 317 5086 656 5113
rect 317 5052 323 5086
rect 357 5074 656 5086
rect 357 5052 439 5074
rect 317 5040 439 5052
rect 473 5040 656 5074
rect 317 5014 656 5040
rect 317 4980 323 5014
rect 357 5001 656 5014
rect 357 4980 439 5001
rect 317 4967 439 4980
rect 473 4967 656 5001
rect 317 4942 656 4967
rect 317 4908 323 4942
rect 357 4928 656 4942
rect 357 4908 439 4928
rect 317 4894 439 4908
rect 473 4894 656 4928
rect 317 4870 656 4894
rect 317 4836 323 4870
rect 357 4855 656 4870
rect 357 4836 439 4855
rect 317 4821 439 4836
rect 473 4821 656 4855
rect 317 4798 656 4821
rect 317 4764 323 4798
rect 357 4781 656 4798
rect 357 4764 439 4781
rect 317 4747 439 4764
rect 473 4747 656 4781
rect 317 4726 656 4747
rect 317 4692 323 4726
rect 357 4707 656 4726
rect 357 4692 439 4707
rect 317 4673 439 4692
rect 473 4673 656 4707
rect 317 4654 656 4673
rect 317 4620 323 4654
rect 357 4633 656 4654
rect 357 4620 439 4633
rect 317 4599 439 4620
rect 473 4599 656 4633
rect 317 4582 656 4599
rect 317 4548 323 4582
rect 357 4559 656 4582
rect 357 4548 439 4559
rect 317 4525 439 4548
rect 473 4525 656 4559
rect 317 4510 656 4525
rect 317 4476 323 4510
rect 357 4485 656 4510
rect 357 4476 439 4485
rect 317 4451 439 4476
rect 473 4451 656 4485
rect 317 4438 656 4451
rect 317 4404 323 4438
rect 357 4411 656 4438
rect 357 4404 439 4411
rect 317 4377 439 4404
rect 473 4377 656 4411
rect 317 4366 656 4377
rect 317 4332 323 4366
rect 357 4337 656 4366
rect 357 4332 439 4337
rect 317 4303 439 4332
rect 473 4303 656 4337
rect 317 4294 656 4303
rect 317 4260 323 4294
rect 357 4263 656 4294
rect 357 4260 439 4263
rect 317 4229 439 4260
rect 473 4229 656 4263
rect 317 4222 656 4229
rect 317 4188 323 4222
rect 357 4189 656 4222
rect 357 4188 439 4189
rect 317 4155 439 4188
rect 473 4155 656 4189
rect 317 4150 656 4155
rect 317 4116 323 4150
rect 357 4116 656 4150
rect 317 4115 656 4116
rect 317 4081 439 4115
rect 473 4081 656 4115
rect 317 4078 656 4081
rect 317 4044 323 4078
rect 357 4044 656 4078
rect 317 4041 656 4044
rect 317 4007 439 4041
rect 473 4007 656 4041
rect 317 4005 656 4007
rect 317 3971 323 4005
rect 357 3971 656 4005
rect 317 3967 656 3971
rect 317 3933 439 3967
rect 473 3933 656 3967
rect 317 3932 656 3933
rect 317 3898 323 3932
rect 357 3898 656 3932
rect 317 3893 656 3898
rect 317 3859 439 3893
rect 473 3859 656 3893
rect 317 3825 323 3859
rect 357 3825 656 3859
rect 317 3819 656 3825
rect 317 3786 439 3819
rect 317 3752 323 3786
rect 357 3785 439 3786
rect 473 3785 656 3819
rect 357 3752 656 3785
rect 317 3713 656 3752
rect 317 3679 323 3713
rect 357 3679 656 3713
tri 684 5865 705 5886 se
rect 705 5865 1035 5886
tri 1035 5865 1084 5914 sw
tri 1084 5886 1112 5914 ne
rect 684 5859 1084 5865
rect 684 5825 696 5859
rect 730 5825 781 5859
rect 815 5825 866 5859
rect 900 5825 952 5859
rect 986 5825 1038 5859
rect 1072 5825 1084 5859
rect 684 3729 1084 5825
rect 684 3695 696 3729
rect 730 3695 781 3729
rect 815 3695 866 3729
rect 900 3695 952 3729
rect 986 3695 1038 3729
rect 1072 3695 1084 3729
rect 684 3689 1084 3695
rect 1112 5731 1512 5914
tri 1512 5886 1540 5914 nw
tri 1561 5886 1589 5914 se
rect 1589 5886 1891 5914
rect 1112 5697 1295 5731
rect 1329 5697 1512 5731
rect 1112 5658 1512 5697
rect 1112 5624 1295 5658
rect 1329 5624 1512 5658
rect 1112 5585 1512 5624
rect 1112 5551 1295 5585
rect 1329 5551 1512 5585
rect 1112 5512 1512 5551
rect 1112 5478 1295 5512
rect 1329 5478 1512 5512
rect 1112 5439 1512 5478
rect 1112 5405 1295 5439
rect 1329 5405 1512 5439
rect 1112 5366 1512 5405
rect 1112 5332 1295 5366
rect 1329 5332 1512 5366
rect 1112 5293 1512 5332
rect 1112 5259 1295 5293
rect 1329 5259 1512 5293
rect 1112 5220 1512 5259
rect 1112 5186 1295 5220
rect 1329 5186 1512 5220
rect 1112 5147 1512 5186
rect 1112 5113 1295 5147
rect 1329 5113 1512 5147
rect 1112 5074 1512 5113
rect 1112 5040 1295 5074
rect 1329 5040 1512 5074
rect 1112 5001 1512 5040
rect 1112 4967 1295 5001
rect 1329 4967 1512 5001
rect 1112 4928 1512 4967
rect 1112 4894 1295 4928
rect 1329 4894 1512 4928
rect 1112 4855 1512 4894
rect 1112 4821 1295 4855
rect 1329 4821 1512 4855
rect 1112 4781 1512 4821
rect 1112 4747 1295 4781
rect 1329 4747 1512 4781
rect 1112 4707 1512 4747
rect 1112 4673 1295 4707
rect 1329 4673 1512 4707
rect 1112 4633 1512 4673
rect 1112 4599 1295 4633
rect 1329 4599 1512 4633
rect 1112 4559 1512 4599
rect 1112 4525 1295 4559
rect 1329 4525 1512 4559
rect 1112 4485 1512 4525
rect 1112 4451 1295 4485
rect 1329 4451 1512 4485
rect 1112 4411 1512 4451
rect 1112 4377 1295 4411
rect 1329 4377 1512 4411
rect 1112 4337 1512 4377
rect 1112 4303 1295 4337
rect 1329 4303 1512 4337
rect 1112 4263 1512 4303
rect 1112 4229 1295 4263
rect 1329 4229 1512 4263
rect 1112 4189 1512 4229
rect 1112 4155 1295 4189
rect 1329 4155 1512 4189
rect 1112 4115 1512 4155
rect 1112 4081 1295 4115
rect 1329 4081 1512 4115
rect 1112 4041 1512 4081
rect 1112 4007 1295 4041
rect 1329 4007 1512 4041
rect 1112 3967 1512 4007
rect 1112 3933 1295 3967
rect 1329 3933 1512 3967
rect 1112 3893 1512 3933
rect 1112 3859 1295 3893
rect 1329 3859 1512 3893
rect 1112 3819 1512 3859
rect 1112 3785 1295 3819
rect 1329 3785 1512 3819
rect 317 3645 656 3679
tri 656 3645 671 3660 sw
tri 1097 3645 1112 3660 se
rect 1112 3645 1512 3785
tri 1540 5865 1561 5886 se
rect 1561 5865 1891 5886
tri 1891 5865 1940 5914 sw
tri 1940 5886 1968 5914 ne
rect 1540 5859 1940 5865
rect 1540 5825 1552 5859
rect 1586 5825 1637 5859
rect 1671 5825 1722 5859
rect 1756 5825 1808 5859
rect 1842 5825 1894 5859
rect 1928 5825 1940 5859
rect 1540 3729 1940 5825
rect 1540 3695 1552 3729
rect 1586 3695 1637 3729
rect 1671 3695 1722 3729
rect 1756 3695 1808 3729
rect 1842 3695 1894 3729
rect 1928 3695 1940 3729
rect 1540 3689 1940 3695
rect 1968 5731 2368 5914
tri 2368 5886 2396 5914 nw
tri 2417 5886 2445 5914 se
rect 2445 5886 2747 5914
rect 1968 5697 2151 5731
rect 2185 5697 2368 5731
rect 1968 5658 2368 5697
rect 1968 5624 2151 5658
rect 2185 5624 2368 5658
rect 1968 5585 2368 5624
rect 1968 5551 2151 5585
rect 2185 5551 2368 5585
rect 1968 5512 2368 5551
rect 1968 5478 2151 5512
rect 2185 5478 2368 5512
rect 1968 5439 2368 5478
rect 1968 5405 2151 5439
rect 2185 5405 2368 5439
rect 1968 5366 2368 5405
rect 1968 5332 2151 5366
rect 2185 5332 2368 5366
rect 1968 5293 2368 5332
rect 1968 5259 2151 5293
rect 2185 5259 2368 5293
rect 1968 5220 2368 5259
rect 1968 5186 2151 5220
rect 2185 5186 2368 5220
rect 1968 5147 2368 5186
rect 1968 5113 2151 5147
rect 2185 5113 2368 5147
rect 1968 5074 2368 5113
rect 1968 5040 2151 5074
rect 2185 5040 2368 5074
rect 1968 5001 2368 5040
rect 1968 4967 2151 5001
rect 2185 4967 2368 5001
rect 1968 4928 2368 4967
rect 1968 4894 2151 4928
rect 2185 4894 2368 4928
rect 1968 4855 2368 4894
rect 1968 4821 2151 4855
rect 2185 4821 2368 4855
rect 1968 4781 2368 4821
rect 1968 4747 2151 4781
rect 2185 4747 2368 4781
rect 1968 4707 2368 4747
rect 1968 4673 2151 4707
rect 2185 4673 2368 4707
rect 1968 4633 2368 4673
rect 1968 4599 2151 4633
rect 2185 4599 2368 4633
rect 1968 4559 2368 4599
rect 1968 4525 2151 4559
rect 2185 4525 2368 4559
rect 1968 4485 2368 4525
rect 1968 4451 2151 4485
rect 2185 4451 2368 4485
rect 1968 4411 2368 4451
rect 1968 4377 2151 4411
rect 2185 4377 2368 4411
rect 1968 4337 2368 4377
rect 1968 4303 2151 4337
rect 2185 4303 2368 4337
rect 1968 4263 2368 4303
rect 1968 4229 2151 4263
rect 2185 4229 2368 4263
rect 1968 4189 2368 4229
rect 1968 4155 2151 4189
rect 2185 4155 2368 4189
rect 1968 4115 2368 4155
rect 1968 4081 2151 4115
rect 2185 4081 2368 4115
rect 1968 4041 2368 4081
rect 1968 4007 2151 4041
rect 2185 4007 2368 4041
rect 1968 3967 2368 4007
rect 1968 3933 2151 3967
rect 2185 3933 2368 3967
rect 1968 3893 2368 3933
rect 1968 3859 2151 3893
rect 2185 3859 2368 3893
rect 1968 3819 2368 3859
rect 1968 3785 2151 3819
rect 2185 3785 2368 3819
tri 1512 3645 1527 3660 sw
tri 1953 3645 1968 3660 se
rect 1968 3645 2368 3785
tri 2396 5865 2417 5886 se
rect 2417 5865 2747 5886
tri 2747 5865 2796 5914 sw
tri 2796 5886 2824 5914 ne
rect 2396 5859 2796 5865
rect 2396 5825 2408 5859
rect 2442 5825 2493 5859
rect 2527 5825 2578 5859
rect 2612 5825 2664 5859
rect 2698 5825 2750 5859
rect 2784 5825 2796 5859
rect 2396 3729 2796 5825
rect 2396 3695 2408 3729
rect 2442 3695 2493 3729
rect 2527 3695 2578 3729
rect 2612 3695 2664 3729
rect 2698 3695 2750 3729
rect 2784 3695 2796 3729
rect 2396 3689 2796 3695
rect 2824 5731 3224 5914
tri 3224 5886 3252 5914 nw
tri 3273 5886 3301 5914 se
rect 3301 5886 3603 5914
rect 2824 5697 3007 5731
rect 3041 5697 3224 5731
rect 2824 5658 3224 5697
rect 2824 5624 3007 5658
rect 3041 5624 3224 5658
rect 2824 5585 3224 5624
rect 2824 5551 3007 5585
rect 3041 5551 3224 5585
rect 2824 5512 3224 5551
rect 2824 5478 3007 5512
rect 3041 5478 3224 5512
rect 2824 5439 3224 5478
rect 2824 5405 3007 5439
rect 3041 5405 3224 5439
rect 2824 5366 3224 5405
rect 2824 5332 3007 5366
rect 3041 5332 3224 5366
rect 2824 5293 3224 5332
rect 2824 5259 3007 5293
rect 3041 5259 3224 5293
rect 2824 5220 3224 5259
rect 2824 5186 3007 5220
rect 3041 5186 3224 5220
rect 2824 5147 3224 5186
rect 2824 5113 3007 5147
rect 3041 5113 3224 5147
rect 2824 5074 3224 5113
rect 2824 5040 3007 5074
rect 3041 5040 3224 5074
rect 2824 5001 3224 5040
rect 2824 4967 3007 5001
rect 3041 4967 3224 5001
rect 2824 4928 3224 4967
rect 2824 4894 3007 4928
rect 3041 4894 3224 4928
rect 2824 4855 3224 4894
rect 2824 4821 3007 4855
rect 3041 4821 3224 4855
rect 2824 4781 3224 4821
rect 2824 4747 3007 4781
rect 3041 4747 3224 4781
rect 2824 4707 3224 4747
rect 2824 4673 3007 4707
rect 3041 4673 3224 4707
rect 2824 4633 3224 4673
rect 2824 4599 3007 4633
rect 3041 4599 3224 4633
rect 2824 4559 3224 4599
rect 2824 4525 3007 4559
rect 3041 4525 3224 4559
rect 2824 4485 3224 4525
rect 2824 4451 3007 4485
rect 3041 4451 3224 4485
rect 2824 4411 3224 4451
rect 2824 4377 3007 4411
rect 3041 4377 3224 4411
rect 2824 4337 3224 4377
rect 2824 4303 3007 4337
rect 3041 4303 3224 4337
rect 2824 4263 3224 4303
rect 2824 4229 3007 4263
rect 3041 4229 3224 4263
rect 2824 4189 3224 4229
rect 2824 4155 3007 4189
rect 3041 4155 3224 4189
rect 2824 4115 3224 4155
rect 2824 4081 3007 4115
rect 3041 4081 3224 4115
rect 2824 4041 3224 4081
rect 2824 4007 3007 4041
rect 3041 4007 3224 4041
rect 2824 3967 3224 4007
rect 2824 3933 3007 3967
rect 3041 3933 3224 3967
rect 2824 3893 3224 3933
rect 2824 3859 3007 3893
rect 3041 3859 3224 3893
rect 2824 3819 3224 3859
rect 2824 3785 3007 3819
rect 3041 3785 3224 3819
tri 2368 3645 2383 3660 sw
tri 2809 3645 2824 3660 se
rect 2824 3645 3224 3785
tri 3252 5865 3273 5886 se
rect 3273 5865 3603 5886
tri 3603 5865 3652 5914 sw
tri 3652 5886 3680 5914 ne
rect 3252 5859 3652 5865
rect 3252 5825 3264 5859
rect 3298 5825 3349 5859
rect 3383 5825 3434 5859
rect 3468 5825 3520 5859
rect 3554 5825 3606 5859
rect 3640 5825 3652 5859
rect 3252 3729 3652 5825
rect 3252 3695 3264 3729
rect 3298 3695 3349 3729
rect 3383 3695 3434 3729
rect 3468 3695 3520 3729
rect 3554 3695 3606 3729
rect 3640 3695 3652 3729
rect 3252 3689 3652 3695
rect 3680 5731 4080 5914
tri 4080 5891 4108 5919 nw
tri 4134 5891 4162 5919 se
rect 4162 5891 4454 5919
rect 3680 5697 3863 5731
rect 3897 5697 4080 5731
rect 3680 5658 4080 5697
rect 3680 5624 3863 5658
rect 3897 5624 4080 5658
rect 3680 5585 4080 5624
rect 3680 5551 3863 5585
rect 3897 5551 4080 5585
rect 3680 5512 4080 5551
rect 3680 5478 3863 5512
rect 3897 5478 4080 5512
rect 3680 5439 4080 5478
rect 3680 5405 3863 5439
rect 3897 5405 4080 5439
rect 3680 5366 4080 5405
rect 3680 5332 3863 5366
rect 3897 5332 4080 5366
rect 3680 5293 4080 5332
rect 3680 5259 3863 5293
rect 3897 5259 4080 5293
rect 3680 5220 4080 5259
rect 3680 5186 3863 5220
rect 3897 5186 4080 5220
rect 3680 5147 4080 5186
rect 3680 5113 3863 5147
rect 3897 5113 4080 5147
rect 3680 5074 4080 5113
rect 3680 5040 3863 5074
rect 3897 5040 4080 5074
rect 3680 5001 4080 5040
rect 3680 4967 3863 5001
rect 3897 4967 4080 5001
rect 3680 4928 4080 4967
rect 3680 4894 3863 4928
rect 3897 4894 4080 4928
rect 3680 4855 4080 4894
rect 3680 4821 3863 4855
rect 3897 4821 4080 4855
rect 3680 4781 4080 4821
rect 3680 4747 3863 4781
rect 3897 4747 4080 4781
rect 3680 4707 4080 4747
rect 3680 4673 3863 4707
rect 3897 4673 4080 4707
rect 3680 4633 4080 4673
rect 3680 4599 3863 4633
rect 3897 4599 4080 4633
rect 3680 4559 4080 4599
rect 3680 4525 3863 4559
rect 3897 4525 4080 4559
rect 3680 4485 4080 4525
rect 3680 4451 3863 4485
rect 3897 4451 4080 4485
rect 3680 4411 4080 4451
rect 3680 4377 3863 4411
rect 3897 4377 4080 4411
rect 3680 4337 4080 4377
rect 3680 4303 3863 4337
rect 3897 4303 4080 4337
rect 3680 4263 4080 4303
rect 3680 4229 3863 4263
rect 3897 4229 4080 4263
rect 3680 4189 4080 4229
rect 3680 4155 3863 4189
rect 3897 4155 4080 4189
rect 3680 4115 4080 4155
rect 3680 4081 3863 4115
rect 3897 4081 4080 4115
rect 3680 4041 4080 4081
rect 3680 4007 3863 4041
rect 3897 4007 4080 4041
rect 3680 3967 4080 4007
rect 3680 3933 3863 3967
rect 3897 3933 4080 3967
rect 3680 3893 4080 3933
rect 3680 3859 3863 3893
rect 3897 3859 4080 3893
rect 3680 3819 4080 3859
rect 3680 3785 3863 3819
rect 3897 3785 4080 3819
tri 3224 3645 3239 3660 sw
tri 3665 3645 3680 3660 se
rect 3680 3645 4080 3785
tri 4108 5865 4134 5891 se
rect 4134 5865 4454 5891
tri 4454 5865 4508 5919 sw
tri 4508 5891 4536 5919 ne
rect 4536 5918 4757 5919
rect 4809 5918 4821 5970
rect 4536 5905 4831 5918
rect 4108 5859 4508 5865
rect 4108 5825 4120 5859
rect 4154 5825 4205 5859
rect 4239 5825 4290 5859
rect 4324 5825 4376 5859
rect 4410 5825 4462 5859
rect 4496 5825 4508 5859
rect 4108 3729 4508 5825
rect 4108 3695 4120 3729
rect 4154 3695 4205 3729
rect 4239 3695 4290 3729
rect 4324 3695 4376 3729
rect 4410 3695 4462 3729
rect 4496 3695 4508 3729
rect 4108 3689 4508 3695
rect 4536 5853 4757 5905
rect 4809 5853 4821 5905
rect 4536 5840 4831 5853
rect 4536 5788 4757 5840
rect 4809 5788 4821 5840
rect 4536 5775 4831 5788
rect 4536 5731 4757 5775
rect 4536 5697 4719 5731
rect 4753 5723 4757 5731
rect 4809 5723 4821 5775
rect 4753 5710 4831 5723
rect 4753 5697 4757 5710
rect 4536 5658 4757 5697
rect 4809 5658 4821 5710
rect 4536 5624 4719 5658
rect 4753 5645 4831 5658
rect 4753 5624 4757 5645
rect 4536 5593 4757 5624
rect 4809 5593 4821 5645
rect 4536 5585 4831 5593
rect 4536 5551 4719 5585
rect 4753 5580 4831 5585
rect 4753 5551 4757 5580
rect 4536 5528 4757 5551
rect 4809 5528 4821 5580
rect 4536 5515 4831 5528
rect 4536 5512 4757 5515
rect 4536 5478 4719 5512
rect 4753 5478 4757 5512
rect 4536 5463 4757 5478
rect 4809 5463 4821 5515
rect 4536 5450 4831 5463
rect 4536 5439 4757 5450
rect 4536 5405 4719 5439
rect 4753 5405 4757 5439
rect 4536 5398 4757 5405
rect 4809 5398 4821 5450
rect 4536 5385 4831 5398
rect 4536 5366 4757 5385
rect 4536 5332 4719 5366
rect 4753 5333 4757 5366
rect 4809 5333 4821 5385
rect 4753 5332 4831 5333
rect 4536 5320 4831 5332
rect 4536 5293 4757 5320
rect 4536 5259 4719 5293
rect 4753 5268 4757 5293
rect 4809 5268 4821 5320
rect 4753 5259 4831 5268
rect 4536 5255 4831 5259
rect 4536 5220 4757 5255
rect 4536 5186 4719 5220
rect 4753 5203 4757 5220
rect 4809 5203 4821 5255
rect 4753 5190 4831 5203
rect 4753 5186 4757 5190
rect 4536 5147 4757 5186
rect 4536 5113 4719 5147
rect 4753 5138 4757 5147
rect 4809 5138 4821 5190
rect 4753 5125 4831 5138
rect 4753 5113 4757 5125
rect 4536 5074 4757 5113
rect 4536 5040 4719 5074
rect 4753 5073 4757 5074
rect 4809 5073 4821 5125
rect 4753 5060 4831 5073
rect 4753 5040 4757 5060
rect 4536 5008 4757 5040
rect 4809 5008 4821 5060
rect 4536 5001 4831 5008
rect 4536 4967 4719 5001
rect 4753 4995 4831 5001
rect 4753 4967 4757 4995
rect 4536 4943 4757 4967
rect 4809 4943 4821 4995
rect 4536 4930 4831 4943
rect 4536 4928 4757 4930
rect 4536 4894 4719 4928
rect 4753 4894 4757 4928
rect 4536 4878 4757 4894
rect 4809 4878 4821 4930
rect 4536 4865 4831 4878
rect 4536 4855 4757 4865
rect 4536 4821 4719 4855
rect 4753 4821 4757 4855
rect 4536 4813 4757 4821
rect 4809 4813 4821 4865
rect 4536 4800 4831 4813
rect 4536 4781 4757 4800
rect 4536 4747 4719 4781
rect 4753 4748 4757 4781
rect 4809 4748 4821 4800
rect 4753 4747 4831 4748
rect 4536 4735 4831 4747
rect 4536 4707 4757 4735
rect 4536 4673 4719 4707
rect 4753 4683 4757 4707
rect 4809 4683 4821 4735
rect 4753 4673 4831 4683
rect 4536 4670 4831 4673
rect 4536 4633 4757 4670
rect 4536 4599 4719 4633
rect 4753 4618 4757 4633
rect 4809 4618 4821 4670
rect 4753 4605 4831 4618
rect 4753 4599 4757 4605
rect 4536 4559 4757 4599
rect 4536 4525 4719 4559
rect 4753 4553 4757 4559
rect 4809 4553 4821 4605
rect 4753 4540 4831 4553
rect 4753 4525 4757 4540
rect 4536 4488 4757 4525
rect 4809 4488 4821 4540
rect 4536 4485 4831 4488
rect 4536 4451 4719 4485
rect 4753 4475 4831 4485
rect 4753 4451 4757 4475
rect 4536 4423 4757 4451
rect 4809 4423 4821 4475
rect 4536 4411 4831 4423
rect 4536 4377 4719 4411
rect 4753 4410 4831 4411
rect 4753 4377 4757 4410
rect 4536 4358 4757 4377
rect 4809 4358 4821 4410
rect 4536 4345 4831 4358
rect 4536 4337 4757 4345
rect 4536 4303 4719 4337
rect 4753 4303 4757 4337
rect 4536 4293 4757 4303
rect 4809 4293 4821 4345
rect 4536 4280 4831 4293
rect 4536 4263 4757 4280
rect 4536 4229 4719 4263
rect 4753 4229 4757 4263
rect 4536 4228 4757 4229
rect 4809 4228 4821 4280
rect 4536 4215 4831 4228
rect 4536 4189 4757 4215
rect 4536 4155 4719 4189
rect 4753 4163 4757 4189
rect 4809 4163 4821 4215
rect 4753 4155 4831 4163
rect 4536 4150 4831 4155
rect 4536 4115 4757 4150
rect 4536 4081 4719 4115
rect 4753 4098 4757 4115
rect 4809 4098 4821 4150
rect 4753 4085 4831 4098
rect 4753 4081 4757 4085
rect 4536 4041 4757 4081
rect 4536 4007 4719 4041
rect 4753 4033 4757 4041
rect 4809 4033 4821 4085
rect 4873 4033 4885 4044
rect 4937 4033 4943 6060
tri 4943 6035 4968 6060 nw
tri 6530 6035 6555 6060 ne
rect 4753 4020 4943 4033
rect 4753 4007 4757 4020
rect 4536 3968 4757 4007
rect 4809 3968 4821 4020
rect 4873 3968 4885 4020
rect 4937 3968 4943 4020
rect 4536 3967 4943 3968
rect 4536 3933 4719 3967
rect 4753 3955 4943 3967
rect 4753 3933 4757 3955
rect 4536 3903 4757 3933
rect 4809 3903 4821 3955
rect 4873 3903 4885 3955
rect 4536 3898 4831 3903
rect 4865 3898 4903 3903
rect 4937 3898 4943 3955
rect 4536 3893 4943 3898
rect 4536 3859 4719 3893
rect 4753 3890 4943 3893
rect 4753 3859 4757 3890
rect 4536 3819 4757 3859
rect 4536 3785 4719 3819
rect 4753 3785 4757 3819
tri 4080 3645 4095 3660 sw
tri 4521 3645 4536 3660 se
rect 4536 3645 4757 3785
rect 317 3640 671 3645
tri 671 3640 676 3645 sw
tri 1092 3640 1097 3645 se
rect 1097 3640 1527 3645
tri 1527 3640 1532 3645 sw
tri 1948 3640 1953 3645 se
rect 1953 3640 2383 3645
tri 2383 3640 2388 3645 sw
tri 2804 3640 2809 3645 se
rect 2809 3640 3239 3645
tri 3239 3640 3244 3645 sw
tri 3660 3640 3665 3645 se
rect 3665 3640 4095 3645
tri 4095 3640 4100 3645 sw
tri 4516 3640 4521 3645 se
rect 4521 3640 4757 3645
rect 317 3606 323 3640
rect 357 3614 676 3640
tri 676 3614 702 3640 sw
tri 1066 3614 1092 3640 se
rect 1092 3614 1532 3640
tri 1532 3614 1558 3640 sw
tri 1922 3614 1948 3640 se
rect 1948 3614 2388 3640
tri 2388 3614 2414 3640 sw
tri 2778 3614 2804 3640 se
rect 2804 3614 3244 3640
tri 3244 3614 3270 3640 sw
tri 3634 3614 3660 3640 se
rect 3660 3614 4100 3640
tri 4100 3614 4126 3640 sw
tri 4490 3614 4516 3640 se
rect 4516 3614 4757 3640
rect 357 3606 4757 3614
rect 317 3596 4757 3606
rect 317 3567 1376 3596
rect 317 3533 323 3567
rect 357 3544 1376 3567
rect 1428 3544 1441 3596
rect 1493 3544 1506 3596
rect 1558 3544 1572 3596
rect 1624 3544 1638 3596
rect 1690 3544 4757 3596
rect 357 3533 4757 3544
rect 317 3532 4757 3533
rect 317 3494 1376 3532
tri 41 3460 42 3461 se
rect 42 3460 108 3461
tri 108 3460 129 3481 sw
rect 317 3460 323 3494
rect 357 3488 1376 3494
rect 1428 3488 1441 3532
rect 1493 3488 1506 3532
rect 1558 3488 1572 3532
rect 1624 3488 1638 3532
rect 1690 3488 4757 3532
rect 4937 3517 4943 3890
rect 6555 6028 6601 6060
tri 6601 6035 6626 6060 nw
tri 7372 6035 7397 6060 ne
rect 6555 5994 6561 6028
rect 6595 5994 6601 6028
rect 6555 5955 6601 5994
rect 6555 5921 6561 5955
rect 6595 5921 6601 5955
rect 6555 5882 6601 5921
rect 7397 6018 7443 6060
tri 7443 6035 7468 6060 nw
tri 7866 6035 7891 6060 ne
rect 7891 6035 7907 6060
tri 7891 6020 7906 6035 ne
rect 7906 6023 7907 6035
rect 7906 6020 7959 6023
rect 8592 6021 8598 6073
rect 8650 6021 8662 6073
rect 8714 6067 8720 6073
tri 8720 6067 8726 6073 sw
tri 9592 6067 9598 6073 se
rect 9598 6067 9658 6073
tri 9658 6067 9679 6088 nw
rect 9757 6080 9764 6088
rect 9870 6080 10870 6088
rect 8714 6021 9612 6067
tri 9612 6021 9658 6067 nw
rect 7397 5984 7403 6018
rect 7437 5984 7443 6018
rect 7397 5942 7443 5984
rect 7397 5908 7403 5942
rect 7437 5908 7443 5942
rect 6555 5848 6561 5882
rect 6595 5848 6601 5882
rect 6555 5809 6601 5848
rect 6555 5775 6561 5809
rect 6595 5775 6601 5809
rect 6555 5736 6601 5775
rect 6555 5702 6561 5736
rect 6595 5702 6601 5736
rect 6555 5663 6601 5702
rect 6555 5629 6561 5663
rect 6595 5629 6601 5663
rect 6555 5590 6601 5629
rect 6555 5556 6561 5590
rect 6595 5556 6601 5590
rect 6555 5517 6601 5556
rect 6555 5483 6561 5517
rect 6595 5483 6601 5517
rect 6555 5443 6601 5483
rect 6555 5409 6561 5443
rect 6595 5409 6601 5443
rect 6555 5369 6601 5409
rect 6555 5335 6561 5369
rect 6595 5335 6601 5369
rect 6555 5295 6601 5335
rect 6555 5261 6561 5295
rect 6595 5261 6601 5295
rect 6555 5221 6601 5261
rect 6555 5187 6561 5221
rect 6595 5187 6601 5221
rect 6555 5147 6601 5187
rect 6555 5113 6561 5147
rect 6595 5113 6601 5147
rect 6555 5073 6601 5113
rect 6555 5039 6561 5073
rect 6595 5039 6601 5073
rect 6555 4999 6601 5039
rect 6555 4965 6561 4999
rect 6595 4965 6601 4999
rect 6555 4925 6601 4965
rect 6555 4891 6561 4925
rect 6595 4891 6601 4925
rect 6555 4851 6601 4891
rect 6555 4817 6561 4851
rect 6595 4817 6601 4851
rect 6555 4777 6601 4817
rect 6555 4743 6561 4777
rect 6595 4743 6601 4777
rect 6555 4703 6601 4743
rect 6555 4669 6561 4703
rect 6595 4669 6601 4703
rect 6555 4629 6601 4669
rect 6555 4595 6561 4629
rect 6595 4595 6601 4629
rect 6555 4555 6601 4595
rect 6555 4521 6561 4555
rect 6595 4521 6601 4555
rect 6555 4481 6601 4521
rect 6555 4447 6561 4481
rect 6595 4447 6601 4481
rect 6555 4407 6601 4447
rect 6555 4373 6561 4407
rect 6595 4373 6601 4407
rect 6555 4333 6601 4373
rect 6555 4299 6561 4333
rect 6595 4299 6601 4333
rect 6555 4259 6601 4299
rect 6555 4225 6561 4259
rect 6595 4225 6601 4259
rect 6555 4185 6601 4225
rect 6555 4151 6561 4185
rect 6595 4151 6601 4185
rect 6555 4111 6601 4151
rect 6555 4077 6561 4111
rect 6595 4077 6601 4111
rect 6555 4037 6601 4077
rect 6555 4003 6561 4037
rect 6595 4003 6601 4037
rect 6555 3963 6601 4003
rect 6699 5882 6745 5894
rect 6699 5848 6705 5882
rect 6739 5848 6745 5882
rect 6699 5810 6745 5848
rect 6699 5776 6705 5810
rect 6739 5776 6745 5810
rect 6699 5738 6745 5776
rect 6699 5704 6705 5738
rect 6739 5704 6745 5738
rect 6699 5666 6745 5704
rect 6699 5632 6705 5666
rect 6739 5632 6745 5666
rect 6699 5594 6745 5632
rect 6699 5560 6705 5594
rect 6739 5560 6745 5594
rect 6699 5522 6745 5560
rect 6699 5488 6705 5522
rect 6739 5488 6745 5522
rect 6699 5450 6745 5488
rect 6699 5416 6705 5450
rect 6739 5416 6745 5450
rect 6699 5378 6745 5416
rect 6699 5344 6705 5378
rect 6739 5344 6745 5378
rect 6699 5306 6745 5344
rect 6699 5272 6705 5306
rect 6739 5272 6745 5306
rect 6699 5234 6745 5272
rect 6699 5200 6705 5234
rect 6739 5200 6745 5234
rect 6699 5162 6745 5200
rect 6699 5128 6705 5162
rect 6739 5128 6745 5162
rect 6699 5090 6745 5128
rect 6699 5056 6705 5090
rect 6739 5056 6745 5090
rect 6699 5018 6745 5056
rect 6699 4984 6705 5018
rect 6739 4984 6745 5018
rect 6699 4946 6745 4984
rect 6699 4912 6705 4946
rect 6739 4912 6745 4946
rect 6699 4874 6745 4912
rect 6699 4840 6705 4874
rect 6739 4840 6745 4874
rect 6699 4802 6745 4840
rect 6699 4768 6705 4802
rect 6739 4768 6745 4802
rect 6699 4730 6745 4768
rect 6699 4696 6705 4730
rect 6739 4696 6745 4730
rect 6699 4658 6745 4696
rect 6699 4624 6705 4658
rect 6739 4624 6745 4658
rect 6699 4586 6745 4624
rect 6699 4552 6705 4586
rect 6739 4552 6745 4586
rect 6699 4514 6745 4552
rect 6699 4480 6705 4514
rect 6739 4480 6745 4514
rect 6699 4442 6745 4480
rect 6699 4408 6705 4442
rect 6739 4408 6745 4442
rect 6699 4370 6745 4408
rect 6699 4336 6705 4370
rect 6739 4336 6745 4370
rect 6699 4298 6745 4336
rect 6699 4264 6705 4298
rect 6739 4264 6745 4298
rect 6699 4226 6745 4264
rect 6699 4192 6705 4226
rect 6739 4192 6745 4226
rect 6935 5882 6981 5894
rect 6935 5848 6941 5882
rect 6975 5848 6981 5882
rect 6935 5809 6981 5848
rect 6935 5775 6941 5809
rect 6975 5775 6981 5809
rect 6935 5736 6981 5775
rect 6935 5702 6941 5736
rect 6975 5702 6981 5736
rect 6935 5663 6981 5702
rect 6935 5629 6941 5663
rect 6975 5629 6981 5663
rect 6935 5590 6981 5629
rect 6935 5556 6941 5590
rect 6975 5556 6981 5590
rect 6935 5517 6981 5556
rect 6935 5483 6941 5517
rect 6975 5483 6981 5517
rect 6935 5444 6981 5483
rect 6935 5410 6941 5444
rect 6975 5410 6981 5444
rect 6935 5371 6981 5410
rect 6935 5337 6941 5371
rect 6975 5337 6981 5371
rect 6935 5298 6981 5337
rect 6935 5264 6941 5298
rect 6975 5264 6981 5298
rect 6935 5225 6981 5264
rect 6935 5191 6941 5225
rect 6975 5191 6981 5225
rect 6935 5152 6981 5191
rect 6935 5118 6941 5152
rect 6975 5118 6981 5152
rect 6935 5079 6981 5118
rect 6935 5045 6941 5079
rect 6975 5045 6981 5079
rect 6935 5006 6981 5045
rect 6935 4972 6941 5006
rect 6975 4972 6981 5006
rect 6935 4933 6981 4972
rect 6935 4899 6941 4933
rect 6975 4899 6981 4933
rect 6935 4860 6981 4899
rect 6935 4826 6941 4860
rect 6975 4826 6981 4860
rect 6935 4787 6981 4826
rect 6935 4753 6941 4787
rect 6975 4753 6981 4787
rect 6935 4714 6981 4753
rect 6935 4680 6941 4714
rect 6975 4680 6981 4714
rect 6935 4641 6981 4680
rect 6935 4607 6941 4641
rect 6975 4607 6981 4641
rect 6935 4568 6981 4607
rect 6935 4534 6941 4568
rect 6975 4534 6981 4568
rect 6935 4495 6981 4534
rect 6935 4461 6941 4495
rect 6975 4461 6981 4495
rect 6935 4422 6981 4461
rect 6935 4388 6941 4422
rect 6975 4388 6981 4422
rect 6935 4349 6981 4388
rect 6935 4315 6941 4349
rect 6975 4315 6981 4349
rect 6935 4276 6981 4315
rect 6935 4242 6941 4276
rect 6975 4242 6981 4276
rect 6699 4154 6745 4192
rect 6699 4120 6705 4154
rect 6739 4120 6745 4154
rect 6699 4082 6745 4120
tri 6932 4214 6935 4217 se
rect 6935 4214 6981 4242
rect 7045 5882 7091 5894
rect 7045 5848 7051 5882
rect 7085 5848 7091 5882
rect 7045 5809 7091 5848
rect 7045 5775 7051 5809
rect 7085 5775 7091 5809
rect 7045 5736 7091 5775
rect 7045 5702 7051 5736
rect 7085 5702 7091 5736
rect 7045 5663 7091 5702
rect 7045 5629 7051 5663
rect 7085 5629 7091 5663
rect 7045 5590 7091 5629
rect 7045 5556 7051 5590
rect 7085 5556 7091 5590
rect 7045 5517 7091 5556
rect 7045 5483 7051 5517
rect 7085 5483 7091 5517
rect 7045 5444 7091 5483
rect 7045 5410 7051 5444
rect 7085 5410 7091 5444
rect 7045 5371 7091 5410
rect 7045 5337 7051 5371
rect 7085 5337 7091 5371
rect 7045 5298 7091 5337
rect 7045 5264 7051 5298
rect 7085 5264 7091 5298
rect 7045 5225 7091 5264
rect 7045 5191 7051 5225
rect 7085 5191 7091 5225
rect 7045 5152 7091 5191
rect 7045 5118 7051 5152
rect 7085 5118 7091 5152
rect 7045 5079 7091 5118
rect 7045 5045 7051 5079
rect 7085 5045 7091 5079
rect 7045 5006 7091 5045
rect 7045 4972 7051 5006
rect 7085 4972 7091 5006
rect 7045 4933 7091 4972
rect 7045 4899 7051 4933
rect 7085 4899 7091 4933
rect 7045 4860 7091 4899
rect 7045 4826 7051 4860
rect 7085 4826 7091 4860
rect 7045 4787 7091 4826
rect 7045 4753 7051 4787
rect 7085 4753 7091 4787
rect 7045 4714 7091 4753
rect 7045 4680 7051 4714
rect 7085 4680 7091 4714
rect 7045 4641 7091 4680
rect 7045 4607 7051 4641
rect 7085 4607 7091 4641
rect 7045 4568 7091 4607
rect 7045 4534 7051 4568
rect 7085 4534 7091 4568
rect 7045 4495 7091 4534
rect 7045 4461 7051 4495
rect 7085 4461 7091 4495
rect 7045 4422 7091 4461
rect 7045 4388 7051 4422
rect 7085 4388 7091 4422
rect 7045 4349 7091 4388
rect 7045 4315 7051 4349
rect 7085 4315 7091 4349
rect 7045 4276 7091 4315
rect 7045 4242 7051 4276
rect 7085 4242 7091 4276
tri 6981 4214 6984 4217 sw
rect 6932 4208 6984 4214
rect 6932 4142 6984 4156
rect 6932 4084 6984 4090
tri 7042 4214 7045 4217 se
rect 7045 4214 7091 4242
rect 7281 5882 7327 5894
rect 7281 5848 7287 5882
rect 7321 5848 7327 5882
rect 7281 5809 7327 5848
rect 7281 5775 7287 5809
rect 7321 5775 7327 5809
rect 7281 5736 7327 5775
rect 7281 5702 7287 5736
rect 7321 5702 7327 5736
rect 7281 5663 7327 5702
rect 7281 5629 7287 5663
rect 7321 5629 7327 5663
rect 7281 5590 7327 5629
rect 7281 5556 7287 5590
rect 7321 5556 7327 5590
rect 7281 5517 7327 5556
rect 7281 5483 7287 5517
rect 7321 5483 7327 5517
rect 7281 5444 7327 5483
rect 7281 5410 7287 5444
rect 7321 5410 7327 5444
rect 7281 5371 7327 5410
rect 7281 5337 7287 5371
rect 7321 5337 7327 5371
rect 7281 5298 7327 5337
rect 7281 5264 7287 5298
rect 7321 5264 7327 5298
rect 7281 5225 7327 5264
rect 7281 5191 7287 5225
rect 7321 5191 7327 5225
rect 7281 5152 7327 5191
rect 7281 5118 7287 5152
rect 7321 5118 7327 5152
rect 7281 5079 7327 5118
rect 7281 5045 7287 5079
rect 7321 5045 7327 5079
rect 7281 5006 7327 5045
rect 7281 4972 7287 5006
rect 7321 4972 7327 5006
rect 7281 4933 7327 4972
rect 7281 4899 7287 4933
rect 7321 4899 7327 4933
rect 7397 5866 7443 5908
rect 7397 5832 7403 5866
rect 7437 5832 7443 5866
rect 7397 5790 7443 5832
rect 7397 5756 7403 5790
rect 7437 5756 7443 5790
rect 7397 5714 7443 5756
rect 7397 5680 7403 5714
rect 7437 5680 7443 5714
rect 7397 5638 7443 5680
rect 7397 5604 7403 5638
rect 7437 5604 7443 5638
rect 7397 5562 7443 5604
rect 7397 5528 7403 5562
rect 7437 5528 7443 5562
rect 7397 5486 7443 5528
rect 7397 5452 7403 5486
rect 7437 5452 7443 5486
rect 7397 5410 7443 5452
rect 7397 5376 7403 5410
rect 7437 5376 7443 5410
rect 7397 5334 7443 5376
rect 7397 5300 7403 5334
rect 7437 5300 7443 5334
rect 7397 5258 7443 5300
rect 7397 5224 7403 5258
rect 7437 5224 7443 5258
rect 7397 5182 7443 5224
rect 7397 5148 7403 5182
rect 7437 5148 7443 5182
rect 7397 5106 7443 5148
rect 7397 5072 7403 5106
rect 7437 5072 7443 5106
rect 7397 5029 7443 5072
rect 7397 4995 7403 5029
rect 7437 4995 7443 5029
rect 7397 4952 7443 4995
rect 7397 4918 7403 4952
rect 7437 4918 7443 4952
rect 7397 4906 7443 4918
rect 7583 6014 7773 6020
tri 7906 6019 7907 6020 ne
rect 7583 6008 7592 6014
rect 7583 5974 7589 6008
rect 7583 5962 7592 5974
rect 7644 5962 7656 6014
rect 7708 5962 7720 6014
rect 7772 5962 7773 6014
rect 7583 5949 7773 5962
rect 7583 5932 7592 5949
rect 7583 5898 7589 5932
rect 7583 5897 7592 5898
rect 7644 5897 7656 5949
rect 7708 5897 7720 5949
rect 7772 5897 7773 5949
rect 7583 5884 7773 5897
rect 7583 5856 7592 5884
rect 7583 5822 7589 5856
rect 7644 5832 7656 5884
rect 7708 5832 7720 5884
rect 7772 5832 7773 5884
rect 7623 5822 7661 5832
rect 7695 5822 7733 5832
rect 7767 5822 7773 5832
rect 7583 5819 7773 5822
rect 7583 5780 7592 5819
rect 7583 5746 7589 5780
rect 7644 5767 7656 5819
rect 7708 5767 7720 5819
rect 7772 5767 7773 5819
rect 7623 5754 7661 5767
rect 7695 5754 7733 5767
rect 7767 5754 7773 5767
rect 7583 5704 7592 5746
rect 7583 5670 7589 5704
rect 7644 5702 7656 5754
rect 7708 5702 7720 5754
rect 7772 5702 7773 5754
rect 7623 5689 7661 5702
rect 7695 5689 7733 5702
rect 7767 5689 7773 5702
rect 7583 5637 7592 5670
rect 7644 5637 7656 5689
rect 7708 5637 7720 5689
rect 7772 5637 7773 5689
rect 7583 5628 7773 5637
rect 7583 5594 7589 5628
rect 7623 5624 7661 5628
rect 7695 5624 7733 5628
rect 7767 5624 7773 5628
rect 7583 5572 7592 5594
rect 7644 5572 7656 5624
rect 7708 5572 7720 5624
rect 7772 5572 7773 5624
rect 7583 5558 7773 5572
rect 7583 5552 7592 5558
rect 7583 5518 7589 5552
rect 7583 5506 7592 5518
rect 7644 5506 7656 5558
rect 7708 5506 7720 5558
rect 7772 5506 7773 5558
rect 7583 5492 7773 5506
rect 7583 5477 7592 5492
rect 7583 5443 7589 5477
rect 7583 5440 7592 5443
rect 7644 5440 7656 5492
rect 7708 5440 7720 5492
rect 7772 5440 7773 5492
rect 7583 5426 7773 5440
rect 7583 5402 7592 5426
rect 7583 5368 7589 5402
rect 7644 5374 7656 5426
rect 7708 5374 7720 5426
rect 7772 5374 7773 5426
rect 7623 5368 7661 5374
rect 7695 5368 7733 5374
rect 7767 5368 7773 5374
rect 7583 5360 7773 5368
rect 7583 5327 7592 5360
rect 7583 5293 7589 5327
rect 7644 5308 7656 5360
rect 7708 5308 7720 5360
rect 7772 5308 7773 5360
rect 7623 5294 7661 5308
rect 7695 5294 7733 5308
rect 7767 5294 7773 5308
rect 7583 5252 7592 5293
rect 7583 5218 7589 5252
rect 7644 5242 7656 5294
rect 7708 5242 7720 5294
rect 7772 5242 7773 5294
rect 7623 5228 7661 5242
rect 7695 5228 7733 5242
rect 7767 5228 7773 5242
rect 7583 5177 7592 5218
rect 7583 5143 7589 5177
rect 7644 5176 7656 5228
rect 7708 5176 7720 5228
rect 7772 5176 7773 5228
rect 7623 5162 7661 5176
rect 7695 5162 7733 5176
rect 7767 5162 7773 5176
rect 7583 5110 7592 5143
rect 7644 5110 7656 5162
rect 7708 5110 7720 5162
rect 7772 5110 7773 5162
rect 7583 5102 7773 5110
rect 7583 5068 7589 5102
rect 7623 5096 7661 5102
rect 7695 5096 7733 5102
rect 7767 5096 7773 5102
rect 7583 5044 7592 5068
rect 7644 5044 7656 5096
rect 7708 5044 7720 5096
rect 7772 5044 7773 5096
rect 7583 5030 7773 5044
rect 7583 5027 7592 5030
rect 7583 4993 7589 5027
rect 7583 4978 7592 4993
rect 7644 4978 7656 5030
rect 7708 4978 7720 5030
rect 7772 4978 7773 5030
rect 7583 4964 7773 4978
rect 7583 4952 7592 4964
rect 7583 4918 7589 4952
rect 7583 4912 7592 4918
rect 7644 4912 7656 4964
rect 7708 4912 7720 4964
rect 7772 4912 7773 4964
rect 7907 6010 7959 6020
rect 7907 5945 7959 5958
rect 8015 5984 8203 5993
rect 8255 5984 8269 5993
rect 8015 5950 8027 5984
rect 8061 5950 8104 5984
rect 8138 5950 8181 5984
rect 8255 5950 8259 5984
rect 8015 5941 8203 5950
rect 8255 5941 8269 5950
rect 8321 5941 8327 5993
rect 8830 5941 8836 5993
rect 8888 5941 8900 5993
rect 8952 5990 8958 5993
tri 8958 5990 8961 5993 sw
rect 8952 5984 9463 5990
rect 8967 5950 9013 5984
rect 9047 5950 9093 5984
rect 9127 5950 9174 5984
rect 9208 5950 9255 5984
rect 9289 5950 9336 5984
rect 9370 5950 9417 5984
rect 9451 5950 9463 5984
rect 9873 6062 10870 6080
rect 10904 6062 11222 6096
rect 11256 6078 13536 6096
rect 11256 6062 13496 6078
rect 9873 6055 13496 6062
rect 9873 6024 12713 6055
rect 9873 5990 10870 6024
rect 10904 5990 11222 6024
rect 11256 6021 12713 6024
rect 12747 6021 13225 6055
rect 13259 6044 13496 6055
rect 13530 6044 13536 6078
rect 13259 6021 13536 6044
rect 11256 6005 13536 6021
rect 11256 5990 13496 6005
rect 9873 5983 13496 5990
rect 9873 5964 12713 5983
rect 9757 5958 12713 5964
tri 10812 5952 10818 5958 ne
rect 10818 5952 12713 5958
rect 8952 5944 9463 5950
tri 10818 5944 10826 5952 ne
rect 10826 5944 10870 5952
rect 8952 5941 8958 5944
tri 8958 5941 8961 5944 nw
tri 10826 5941 10829 5944 ne
rect 10829 5941 10870 5944
tri 10829 5919 10851 5941 ne
rect 10851 5919 10870 5941
rect 7907 5883 7913 5893
rect 7947 5883 7959 5893
rect 7907 5880 7959 5883
rect 8454 5867 8460 5919
rect 8512 5867 8527 5919
rect 8579 5918 8585 5919
tri 8585 5918 8586 5919 sw
tri 10851 5918 10852 5919 ne
rect 10852 5918 10870 5919
rect 10904 5918 11222 5952
rect 11256 5949 12713 5952
rect 12747 5949 13225 5983
rect 13259 5971 13496 5983
rect 13530 5971 13536 6005
rect 13259 5949 13536 5971
rect 11256 5932 13536 5949
rect 11256 5918 13496 5932
rect 8579 5913 8586 5918
tri 8586 5913 8591 5918 sw
tri 10852 5913 10857 5918 ne
rect 10857 5913 13496 5918
rect 8579 5911 10767 5913
tri 10767 5911 10769 5913 sw
tri 10857 5911 10859 5913 ne
rect 10859 5911 13496 5913
rect 8579 5907 10769 5911
rect 8579 5873 8777 5907
rect 8811 5873 8849 5907
rect 8883 5878 10769 5907
tri 10769 5878 10802 5911 sw
tri 10859 5906 10864 5911 ne
rect 10864 5906 12713 5911
tri 12506 5878 12534 5906 ne
rect 12534 5878 12713 5906
rect 8883 5873 12418 5878
tri 12534 5877 12535 5878 ne
rect 12535 5877 12713 5878
rect 12747 5877 13225 5911
rect 13259 5898 13496 5911
rect 13530 5898 13536 5932
rect 13259 5877 13536 5898
rect 8579 5867 12418 5873
tri 10747 5859 10755 5867 ne
rect 10755 5859 12418 5867
tri 12535 5859 12553 5877 ne
rect 12553 5859 13536 5877
tri 10755 5839 10775 5859 ne
rect 10775 5839 12418 5859
tri 12553 5839 12573 5859 ne
rect 12573 5839 13496 5859
tri 8661 5834 8666 5839 se
rect 8666 5834 8718 5839
rect 7907 5815 7913 5828
rect 7947 5815 7959 5828
rect 8083 5828 8277 5834
rect 8329 5828 8343 5834
rect 8395 5828 8718 5834
rect 8083 5794 8095 5828
rect 8129 5794 8175 5828
rect 8209 5794 8255 5828
rect 8329 5794 8336 5828
rect 8395 5794 8417 5828
rect 8451 5794 8498 5828
rect 8532 5794 8579 5828
rect 8613 5794 8718 5828
rect 8083 5782 8277 5794
rect 8329 5782 8343 5794
rect 8395 5787 8718 5794
rect 8719 5788 8720 5838
rect 8756 5788 8757 5838
rect 8758 5828 10386 5839
rect 8758 5794 8933 5828
rect 8967 5794 9014 5828
rect 9048 5794 9095 5828
rect 9129 5794 9177 5828
rect 9211 5794 9259 5828
rect 9293 5794 9341 5828
rect 9375 5794 9423 5828
rect 9457 5794 10386 5828
rect 8758 5787 10386 5794
rect 10438 5787 10450 5839
rect 10502 5787 10508 5839
tri 10775 5832 10782 5839 ne
rect 10782 5832 12418 5839
tri 11375 5820 11387 5832 ne
rect 11387 5820 11518 5832
tri 11387 5810 11397 5820 ne
rect 11397 5810 11406 5820
tri 10596 5798 10608 5810 se
rect 10608 5798 10726 5810
tri 11397 5807 11400 5810 ne
tri 10585 5787 10596 5798 se
rect 10596 5787 10614 5798
rect 8395 5782 8484 5787
tri 8484 5782 8489 5787 nw
tri 10580 5782 10585 5787 se
rect 10585 5782 10614 5787
rect 7907 5750 7913 5763
rect 7947 5750 7959 5763
tri 10557 5759 10580 5782 se
rect 10580 5759 10614 5782
rect 8512 5707 8518 5759
rect 8570 5707 8582 5759
rect 8634 5709 10614 5759
rect 8634 5707 8640 5709
tri 8640 5707 8642 5709 nw
tri 10579 5707 10581 5709 ne
rect 10581 5707 10614 5709
rect 7907 5689 7959 5698
tri 10581 5692 10596 5707 ne
rect 10596 5692 10614 5707
rect 10720 5692 10726 5798
rect 11400 5714 11406 5810
rect 11512 5714 11518 5820
tri 11518 5807 11543 5832 nw
tri 12347 5807 12372 5832 ne
rect 11578 5752 11584 5804
rect 11636 5752 11648 5804
rect 11700 5792 12332 5804
rect 11700 5758 11940 5792
rect 11974 5758 12292 5792
rect 12326 5758 12332 5792
rect 11700 5752 11706 5758
tri 11706 5752 11712 5758 nw
tri 11909 5752 11915 5758 ne
rect 11915 5752 11980 5758
tri 11578 5748 11582 5752 ne
rect 11400 5702 11518 5714
rect 11582 5733 11634 5752
tri 11634 5733 11653 5752 nw
tri 11915 5733 11934 5752 ne
rect 11582 5720 11628 5733
tri 11628 5727 11634 5733 nw
rect 7907 5685 7913 5689
rect 7947 5685 7959 5689
tri 10596 5686 10602 5692 ne
rect 10602 5686 10726 5692
tri 10602 5684 10604 5686 ne
rect 10604 5684 10726 5686
tri 10604 5681 10607 5684 ne
rect 10607 5681 10726 5684
rect 7907 5620 7959 5633
rect 8015 5672 8203 5681
rect 8255 5672 8269 5681
rect 8321 5679 8392 5681
tri 8392 5679 8394 5681 sw
rect 8321 5678 8394 5679
tri 8394 5678 8395 5679 sw
rect 8321 5672 8395 5678
rect 8015 5638 8027 5672
rect 8061 5638 8107 5672
rect 8141 5638 8187 5672
rect 8255 5638 8268 5672
rect 8321 5638 8349 5672
rect 8383 5638 8395 5672
rect 8015 5629 8203 5638
rect 8255 5629 8269 5638
rect 8321 5632 8395 5638
rect 8321 5629 8392 5632
tri 8392 5629 8395 5632 nw
rect 8750 5629 8756 5681
rect 8808 5629 8820 5681
rect 8872 5679 8878 5681
tri 8878 5679 8880 5681 sw
tri 10607 5680 10608 5681 ne
rect 10608 5680 10726 5681
rect 11582 5686 11588 5720
rect 11622 5686 11628 5720
rect 8872 5678 8880 5679
tri 8880 5678 8881 5679 sw
rect 8872 5672 9469 5678
rect 11582 5674 11628 5686
rect 11758 5718 11804 5730
rect 11758 5684 11764 5718
rect 11798 5684 11804 5718
rect 8898 5638 8943 5672
rect 8977 5638 9023 5672
rect 9057 5638 9103 5672
rect 9137 5638 9183 5672
rect 9217 5638 9263 5672
rect 9297 5638 9343 5672
rect 9377 5638 9423 5672
rect 9457 5638 9469 5672
tri 11739 5652 11758 5671 se
rect 11758 5652 11804 5684
rect 11934 5720 11980 5752
tri 11980 5733 12005 5758 nw
tri 12261 5733 12286 5758 ne
rect 11934 5686 11940 5720
rect 11974 5686 11980 5720
rect 11934 5674 11980 5686
rect 12110 5718 12156 5730
rect 12110 5684 12116 5718
rect 12150 5684 12156 5718
rect 8872 5632 9469 5638
rect 8872 5629 8878 5632
tri 8878 5629 8881 5632 nw
rect 9522 5600 9528 5652
rect 9580 5600 9594 5652
rect 9646 5646 9652 5652
tri 9652 5646 9658 5652 sw
tri 11733 5646 11739 5652 se
rect 11739 5646 11804 5652
tri 11804 5646 11829 5671 sw
tri 12085 5646 12110 5671 se
rect 12110 5646 12156 5684
rect 12286 5720 12332 5758
rect 12286 5686 12292 5720
rect 12326 5686 12332 5720
rect 12286 5674 12332 5686
rect 12372 5792 12418 5832
tri 12573 5805 12607 5839 ne
rect 12607 5805 12713 5839
rect 12747 5805 13225 5839
rect 13259 5825 13496 5839
rect 13530 5825 13536 5859
rect 13259 5805 13536 5825
rect 12372 5758 12378 5792
rect 12412 5758 12418 5792
tri 12607 5786 12626 5805 ne
rect 12626 5786 13536 5805
tri 12626 5767 12645 5786 ne
rect 12645 5767 13496 5786
rect 12372 5720 12418 5758
tri 12645 5733 12679 5767 ne
rect 12679 5733 12713 5767
rect 12747 5733 13225 5767
rect 13259 5752 13496 5767
rect 13530 5752 13536 5786
rect 13259 5733 13536 5752
rect 12372 5686 12378 5720
rect 12412 5686 12418 5720
tri 12679 5713 12699 5733 ne
rect 12699 5713 13536 5733
tri 12699 5705 12707 5713 ne
rect 12707 5705 13496 5713
rect 12372 5674 12418 5686
tri 13335 5680 13360 5705 ne
rect 13360 5679 13496 5705
rect 13530 5679 13536 5713
tri 12156 5646 12181 5671 sw
rect 9646 5612 11764 5646
rect 11798 5612 12116 5646
rect 12150 5612 13250 5646
rect 9646 5606 13250 5612
rect 9646 5600 12898 5606
tri 12815 5575 12840 5600 ne
rect 7907 5555 7959 5568
rect 8855 5562 10466 5572
rect 8855 5528 8867 5562
rect 8901 5528 8946 5562
rect 8980 5528 9025 5562
rect 9059 5528 9104 5562
rect 9138 5528 9183 5562
rect 9217 5528 9263 5562
rect 9297 5528 9343 5562
rect 9377 5528 9423 5562
rect 9457 5528 10466 5562
rect 7907 5502 7913 5503
rect 7947 5502 7959 5503
rect 7907 5489 7959 5502
rect 8083 5516 8277 5526
rect 8329 5516 8343 5526
rect 8395 5516 8625 5526
rect 8855 5520 10466 5528
rect 10518 5520 10530 5572
rect 10582 5520 12586 5572
rect 8083 5482 8095 5516
rect 8129 5482 8175 5516
rect 8209 5482 8255 5516
rect 8329 5482 8336 5516
rect 8395 5482 8417 5516
rect 8451 5482 8498 5516
rect 8532 5482 8579 5516
rect 8613 5482 8625 5516
tri 12509 5495 12534 5520 ne
rect 8083 5474 8277 5482
rect 8329 5474 8343 5482
rect 8395 5474 8625 5482
rect 8669 5484 9278 5490
rect 8669 5450 8681 5484
rect 8715 5450 8753 5484
rect 8787 5450 9278 5484
rect 8669 5438 9278 5450
rect 9330 5438 9344 5490
rect 9396 5478 12499 5490
rect 9396 5444 12381 5478
rect 12415 5444 12453 5478
rect 12487 5444 12499 5478
rect 9396 5438 12499 5444
rect 7907 5425 7913 5437
rect 7947 5425 7959 5437
tri 12527 5426 12534 5433 se
rect 12534 5426 12586 5520
rect 7907 5423 7959 5425
tri 12509 5408 12527 5426 se
rect 12527 5408 12586 5426
tri 8984 5396 8986 5398 se
rect 8986 5396 8992 5398
tri 8980 5392 8984 5396 se
rect 8984 5392 8992 5396
rect 8850 5386 8992 5392
rect 9044 5386 9056 5398
rect 9108 5386 9121 5398
rect 9173 5386 9186 5398
rect 9238 5396 9244 5398
tri 9244 5396 9246 5398 sw
rect 12494 5396 12586 5408
rect 9238 5392 9246 5396
tri 9246 5392 9250 5396 sw
rect 9238 5386 9585 5392
rect 7907 5357 7913 5371
rect 7947 5357 7959 5371
tri 8191 5366 8197 5372 se
rect 8197 5366 8203 5372
rect 8015 5360 8203 5366
rect 8255 5360 8269 5372
rect 8321 5366 8327 5372
tri 8327 5366 8333 5372 sw
rect 8321 5360 8625 5366
rect 8015 5326 8027 5360
rect 8061 5326 8105 5360
rect 8139 5326 8184 5360
rect 8255 5326 8263 5360
rect 8321 5326 8342 5360
rect 8376 5326 8421 5360
rect 8455 5326 8500 5360
rect 8534 5326 8579 5360
rect 8613 5352 8625 5360
tri 8625 5352 8639 5366 sw
rect 8850 5352 8862 5386
rect 8896 5352 8937 5386
rect 8971 5352 8992 5386
rect 9046 5352 9056 5386
rect 9271 5352 9312 5386
rect 9346 5352 9387 5386
rect 9421 5352 9463 5386
rect 9497 5352 9539 5386
rect 9573 5352 9585 5386
rect 8613 5336 8639 5352
tri 8639 5336 8655 5352 sw
rect 8850 5346 8992 5352
rect 9044 5346 9056 5352
rect 9108 5346 9121 5352
rect 9173 5346 9186 5352
rect 9238 5346 9585 5352
rect 10300 5375 10672 5382
rect 10674 5381 10710 5382
tri 10293 5336 10300 5343 se
rect 8613 5326 8655 5336
rect 8015 5320 8203 5326
rect 8255 5320 8269 5326
rect 8321 5321 8655 5326
tri 8655 5321 8670 5336 sw
tri 10278 5321 10293 5336 se
rect 10293 5323 10300 5336
rect 10352 5323 10672 5375
rect 10293 5321 10672 5323
rect 8321 5320 8670 5321
rect 7907 5291 7913 5305
rect 7947 5291 7959 5305
tri 8607 5302 8625 5320 ne
rect 8625 5318 8670 5320
tri 8670 5318 8673 5321 sw
tri 10275 5318 10278 5321 se
rect 10278 5318 10672 5321
rect 8625 5302 10208 5318
tri 8625 5290 8637 5302 ne
rect 8637 5290 10208 5302
tri 8637 5288 8639 5290 ne
rect 8639 5288 10208 5290
tri 8639 5287 8640 5288 ne
rect 8640 5287 10208 5288
tri 8640 5266 8661 5287 ne
rect 8661 5266 10208 5287
rect 10209 5267 10210 5317
rect 10246 5267 10247 5317
rect 10248 5310 10672 5318
rect 10248 5266 10300 5310
tri 10286 5259 10293 5266 ne
rect 10293 5259 10300 5266
tri 8426 5256 8429 5259 se
rect 8429 5256 8435 5259
rect 7907 5228 7959 5239
rect 7907 5225 7913 5228
rect 7947 5225 7959 5228
rect 8017 5250 8435 5256
rect 8487 5250 8502 5259
rect 8017 5216 8029 5250
rect 8063 5216 8104 5250
rect 8138 5216 8179 5250
rect 8213 5216 8254 5250
rect 8288 5216 8330 5250
rect 8364 5216 8406 5250
rect 8017 5210 8435 5216
tri 8426 5207 8429 5210 ne
rect 8429 5207 8435 5210
rect 8487 5207 8502 5216
rect 8554 5207 8560 5259
tri 10293 5253 10299 5259 ne
rect 10299 5258 10300 5259
rect 10352 5258 10672 5310
rect 10299 5253 10672 5258
rect 10673 5253 10711 5381
rect 10712 5370 11746 5382
rect 10712 5336 10770 5370
rect 10804 5336 11082 5370
rect 11116 5336 11394 5370
rect 11428 5336 11706 5370
rect 11740 5336 11746 5370
rect 10712 5287 11746 5336
rect 10712 5253 10770 5287
rect 10804 5253 11082 5287
rect 11116 5253 11394 5287
rect 11428 5253 11706 5287
rect 11740 5253 11746 5287
tri 10299 5252 10300 5253 ne
rect 10300 5252 10672 5253
rect 10674 5252 10710 5253
rect 10712 5252 11746 5253
tri 10739 5241 10750 5252 ne
rect 10750 5241 10824 5252
tri 10824 5241 10835 5252 nw
tri 11051 5241 11062 5252 ne
rect 11062 5241 11136 5252
tri 11136 5241 11147 5252 nw
tri 11363 5241 11374 5252 ne
rect 11374 5241 11448 5252
tri 11448 5241 11459 5252 nw
tri 11675 5241 11686 5252 ne
rect 11686 5241 11746 5252
tri 10750 5238 10753 5241 ne
rect 10753 5238 10810 5241
rect 9545 5226 9591 5238
rect 8588 5210 8674 5219
rect 7907 5167 7959 5173
rect 8588 5176 8600 5210
rect 8634 5176 8672 5210
rect 8588 5167 8674 5176
rect 8726 5167 8740 5219
rect 8792 5167 8798 5219
rect 8881 5210 9278 5221
rect 9330 5210 9344 5221
rect 9396 5210 9423 5221
rect 8881 5176 8893 5210
rect 8927 5176 8974 5210
rect 9008 5176 9055 5210
rect 9089 5176 9136 5210
rect 9170 5176 9217 5210
rect 9251 5176 9278 5210
rect 9331 5176 9344 5210
rect 9411 5176 9423 5210
rect 8881 5170 9278 5176
tri 9271 5169 9272 5170 ne
rect 9272 5169 9278 5170
rect 9330 5169 9344 5176
rect 9396 5169 9423 5176
rect 9545 5192 9551 5226
rect 9585 5192 9591 5226
rect 7907 5151 7953 5167
tri 7953 5161 7959 5167 nw
rect 7907 5117 7913 5151
rect 7947 5117 7953 5151
rect 7907 5074 7953 5117
rect 9545 5150 9591 5192
rect 9545 5116 9551 5150
rect 9585 5116 9591 5150
rect 7907 5040 7913 5074
rect 7947 5040 7953 5074
rect 8748 5060 8754 5112
rect 8806 5060 8820 5112
rect 8872 5100 9467 5112
rect 8896 5066 8941 5100
rect 8975 5066 9021 5100
rect 9055 5066 9101 5100
rect 9135 5066 9181 5100
rect 9215 5066 9261 5100
rect 9295 5066 9341 5100
rect 9375 5066 9421 5100
rect 9455 5066 9467 5100
rect 8872 5060 9467 5066
rect 9545 5073 9591 5116
rect 7907 5011 7953 5040
rect 9545 5039 9551 5073
rect 9585 5039 9591 5073
tri 7953 5011 7970 5028 sw
rect 7907 5003 7970 5011
tri 7970 5003 7978 5011 sw
rect 7907 4951 7913 5003
rect 7965 4951 7979 5003
rect 8031 4994 8045 5003
rect 8031 4951 8045 4960
rect 8097 4951 8111 5003
rect 8163 5001 8169 5003
tri 8169 5001 8171 5003 sw
rect 8163 5000 8171 5001
tri 8171 5000 8172 5001 sw
rect 8163 4994 8481 5000
rect 8163 4960 8192 4994
rect 8226 4960 8273 4994
rect 8307 4960 8354 4994
rect 8388 4960 8435 4994
rect 8469 4960 8481 4994
rect 8163 4954 8481 4960
rect 8163 4951 8169 4954
tri 8169 4951 8172 4954 nw
rect 8509 4951 8515 5003
rect 8567 4951 8582 5003
rect 8634 4951 8640 5003
rect 9545 4996 9591 5039
rect 9545 4962 9551 4996
rect 9585 4962 9591 4996
tri 9542 4952 9545 4955 se
rect 9545 4952 9591 4962
tri 8548 4927 8572 4951 ne
rect 8572 4927 8640 4951
tri 8640 4927 8665 4952 sw
tri 9526 4936 9542 4952 se
rect 9542 4936 9591 4952
tri 8980 4930 8986 4936 se
rect 8986 4930 8992 4936
tri 8572 4926 8573 4927 ne
rect 7583 4906 7773 4912
rect 8573 4921 8703 4927
rect 7281 4887 7327 4899
tri 7327 4887 7343 4903 sw
rect 8573 4887 8585 4921
rect 8619 4887 8657 4921
rect 8691 4887 8703 4921
rect 7281 4878 7343 4887
tri 7343 4878 7352 4887 sw
rect 8573 4881 8703 4887
rect 8855 4924 8992 4930
rect 9044 4924 9056 4936
rect 9108 4924 9121 4936
rect 9173 4924 9186 4936
rect 9238 4930 9244 4936
tri 9244 4930 9250 4936 sw
tri 9520 4930 9526 4936 se
rect 9526 4930 9591 4936
rect 9238 4924 9591 4930
rect 8855 4890 8867 4924
rect 8901 4890 8942 4924
rect 8976 4890 8992 4924
rect 9051 4890 9056 4924
rect 9238 4890 9242 4924
rect 9276 4890 9317 4924
rect 9351 4890 9391 4924
rect 9425 4890 9465 4924
rect 9499 4890 9539 4924
rect 9573 4890 9591 4924
rect 8855 4884 8992 4890
rect 9044 4884 9056 4890
rect 9108 4884 9121 4890
rect 9173 4884 9186 4890
rect 9238 4884 9591 4890
rect 9693 5232 9918 5238
rect 9745 5226 9757 5232
rect 9809 5226 9821 5232
rect 9873 5226 9918 5232
tri 10753 5227 10764 5238 ne
rect 9873 5192 9878 5226
rect 9912 5192 9918 5226
rect 9745 5180 9757 5192
rect 9809 5180 9821 5192
rect 9873 5180 9918 5192
rect 9693 5159 9918 5180
rect 9745 5151 9757 5159
rect 9809 5151 9821 5159
rect 9873 5151 9918 5159
rect 9873 5117 9878 5151
rect 9912 5117 9918 5151
rect 9745 5107 9757 5117
rect 9809 5107 9821 5117
rect 9873 5107 9918 5117
rect 9693 5086 9918 5107
rect 9745 5076 9757 5086
rect 9809 5076 9821 5086
rect 9873 5076 9918 5086
rect 9873 5042 9878 5076
rect 9912 5042 9918 5076
rect 9745 5034 9757 5042
rect 9809 5034 9821 5042
rect 9873 5034 9918 5042
rect 9693 5013 9918 5034
rect 9745 5001 9757 5013
rect 9809 5001 9821 5013
rect 9873 5001 9918 5013
rect 9873 4967 9878 5001
rect 9912 4967 9918 5001
rect 10608 5212 10654 5224
rect 10608 5178 10614 5212
rect 10648 5178 10654 5212
rect 10608 5129 10654 5178
rect 10608 5095 10614 5129
rect 10648 5095 10654 5129
rect 10608 5045 10654 5095
rect 10608 5011 10614 5045
rect 10648 5011 10654 5045
tri 10605 4983 10608 4986 se
rect 10608 4983 10654 5011
rect 10764 5203 10810 5238
tri 10810 5227 10824 5241 nw
tri 11062 5227 11076 5241 ne
rect 10764 5169 10770 5203
rect 10804 5169 10810 5203
rect 10764 5119 10810 5169
rect 10764 5085 10770 5119
rect 10804 5085 10810 5119
rect 10764 5035 10810 5085
rect 10764 5001 10770 5035
rect 10804 5001 10810 5035
rect 10764 4989 10810 5001
rect 10920 5212 10966 5224
rect 10920 5178 10926 5212
rect 10960 5178 10966 5212
rect 10920 5129 10966 5178
rect 10920 5095 10926 5129
rect 10960 5095 10966 5129
rect 10920 5045 10966 5095
rect 10920 5011 10926 5045
rect 10960 5011 10966 5045
tri 10654 4983 10657 4986 sw
tri 10917 4983 10920 4986 se
rect 10920 4983 10966 5011
rect 11076 5203 11122 5241
tri 11122 5227 11136 5241 nw
tri 11374 5227 11388 5241 ne
rect 11076 5169 11082 5203
rect 11116 5169 11122 5203
rect 11076 5119 11122 5169
rect 11076 5085 11082 5119
rect 11116 5085 11122 5119
rect 11076 5035 11122 5085
rect 11076 5001 11082 5035
rect 11116 5001 11122 5035
rect 11076 4989 11122 5001
rect 11232 5212 11278 5224
rect 11232 5178 11238 5212
rect 11272 5178 11278 5212
rect 11232 5129 11278 5178
rect 11232 5095 11238 5129
rect 11272 5095 11278 5129
rect 11232 5045 11278 5095
rect 11232 5011 11238 5045
rect 11272 5011 11278 5045
tri 10966 4983 10969 4986 sw
tri 11229 4983 11232 4986 se
rect 11232 4983 11278 5011
rect 11388 5203 11434 5241
tri 11434 5227 11448 5241 nw
tri 11686 5227 11700 5241 ne
rect 11388 5169 11394 5203
rect 11428 5169 11434 5203
rect 11388 5119 11434 5169
rect 11388 5085 11394 5119
rect 11428 5085 11434 5119
rect 11388 5035 11434 5085
rect 11388 5001 11394 5035
rect 11428 5001 11434 5035
rect 11388 4989 11434 5001
rect 11544 5212 11590 5224
rect 11544 5178 11550 5212
rect 11584 5178 11590 5212
rect 11544 5129 11590 5178
rect 11544 5095 11550 5129
rect 11584 5095 11590 5129
rect 11544 5045 11590 5095
rect 11544 5011 11550 5045
rect 11584 5011 11590 5045
tri 11278 4983 11281 4986 sw
tri 11541 4983 11544 4986 se
rect 11544 4983 11590 5011
rect 11700 5203 11746 5241
rect 11700 5169 11706 5203
rect 11740 5169 11746 5203
rect 11700 5119 11746 5169
rect 11700 5085 11706 5119
rect 11740 5085 11746 5119
rect 11700 5035 11746 5085
rect 11700 5001 11706 5035
rect 11740 5001 11746 5035
rect 11700 4989 11746 5001
rect 11856 5370 11902 5382
rect 11856 5336 11862 5370
rect 11896 5336 11902 5370
rect 11856 5288 11902 5336
rect 11856 5254 11862 5288
rect 11896 5254 11902 5288
rect 11856 5206 11902 5254
rect 11856 5172 11862 5206
rect 11896 5172 11902 5206
rect 11856 5124 11902 5172
rect 11856 5090 11862 5124
rect 11896 5090 11902 5124
rect 11856 5042 11902 5090
rect 11856 5008 11862 5042
rect 11896 5008 11902 5042
tri 11590 4983 11593 4986 sw
tri 11853 4983 11856 4986 se
rect 11856 4983 11902 5008
rect 9745 4961 9757 4967
rect 9809 4961 9821 4967
rect 9873 4961 9918 4967
tri 10583 4961 10605 4983 se
rect 10605 4961 10657 4983
tri 10657 4961 10679 4983 sw
tri 10895 4961 10917 4983 se
rect 10917 4961 10969 4983
tri 10969 4961 10991 4983 sw
tri 11207 4961 11229 4983 se
rect 11229 4961 11281 4983
tri 11281 4961 11303 4983 sw
tri 11519 4961 11541 4983 se
rect 11541 4961 11593 4983
tri 11593 4961 11615 4983 sw
tri 11831 4961 11853 4983 se
rect 11853 4961 11902 4983
rect 9693 4939 9918 4961
rect 9745 4927 9757 4939
rect 9809 4927 9821 4939
rect 9873 4927 9918 4939
tri 10266 4927 10300 4961 se
rect 10300 4934 10523 4961
rect 10525 4960 10561 4961
rect 10300 4927 10380 4934
rect 9873 4893 9878 4927
rect 9912 4893 9918 4927
tri 10265 4926 10266 4927 se
rect 10266 4926 10380 4927
tri 10257 4918 10265 4926 se
rect 10265 4918 10380 4926
tri 10249 4910 10257 4918 se
rect 10257 4910 10380 4918
rect 9745 4887 9757 4893
rect 9809 4887 9821 4893
rect 9873 4887 9918 4893
rect 9693 4881 9918 4887
tri 10220 4881 10249 4910 se
rect 10249 4882 10380 4910
rect 10432 4882 10523 4934
rect 10249 4881 10523 4882
tri 10217 4878 10220 4881 se
rect 10220 4878 10523 4881
rect 7281 4877 8534 4878
tri 8534 4877 8535 4878 sw
tri 10216 4877 10217 4878 se
rect 10217 4877 10523 4878
rect 7281 4872 8535 4877
rect 7281 4860 7347 4872
rect 7281 4826 7287 4860
rect 7321 4826 7347 4860
rect 7281 4820 7347 4826
rect 7399 4820 7411 4872
rect 7463 4820 7475 4872
rect 7527 4820 8225 4872
rect 8277 4820 8289 4872
rect 8341 4820 8353 4872
rect 8405 4853 8535 4872
tri 8535 4853 8559 4877 sw
tri 10192 4853 10216 4877 se
rect 10216 4868 10523 4877
rect 10216 4853 10380 4868
rect 8405 4820 10380 4853
rect 7281 4818 10380 4820
rect 7281 4806 8029 4818
rect 7281 4787 7347 4806
rect 7281 4753 7287 4787
rect 7321 4754 7347 4787
rect 7399 4754 7411 4806
rect 7463 4754 7475 4806
rect 7527 4784 8029 4806
rect 8063 4784 8111 4818
rect 8145 4784 8192 4818
rect 8226 4806 8273 4818
rect 8307 4806 8354 4818
rect 8388 4806 8435 4818
rect 7527 4754 8225 4784
rect 8277 4754 8289 4784
rect 8341 4754 8353 4806
rect 8405 4784 8435 4806
rect 8469 4816 10380 4818
rect 10432 4831 10523 4868
rect 10524 4832 10562 4960
rect 10563 4927 10614 4961
rect 10648 4927 10926 4961
rect 10960 4927 11238 4961
rect 11272 4927 11550 4961
rect 11584 4960 11902 4961
rect 11584 4927 11862 4960
rect 10563 4926 11862 4927
rect 11896 4926 11902 4960
rect 10563 4877 11902 4926
rect 10563 4843 10614 4877
rect 10648 4843 10926 4877
rect 10960 4843 11238 4877
rect 11272 4843 11550 4877
rect 11584 4843 11862 4877
rect 11896 4843 11902 4877
rect 10525 4831 10561 4832
rect 10563 4831 11902 4843
rect 11966 5355 12012 5367
rect 11966 5321 11972 5355
rect 12006 5321 12012 5355
rect 11966 5275 12012 5321
rect 11966 5241 11972 5275
rect 12006 5241 12012 5275
rect 11966 5195 12012 5241
rect 11966 5161 11972 5195
rect 12006 5161 12012 5195
rect 11966 5114 12012 5161
rect 11966 5080 11972 5114
rect 12006 5080 12012 5114
rect 11966 5033 12012 5080
rect 11966 4999 11972 5033
rect 12006 4999 12012 5033
rect 11966 4952 12012 4999
rect 11966 4918 11972 4952
rect 12006 4918 12012 4952
rect 11966 4871 12012 4918
rect 11966 4837 11972 4871
rect 12006 4837 12012 4871
rect 8469 4785 10432 4816
tri 10432 4806 10457 4831 nw
tri 11947 4806 11966 4825 se
rect 11966 4806 12012 4837
rect 12318 5355 12364 5367
rect 12318 5321 12324 5355
rect 12358 5321 12364 5355
rect 12318 5276 12364 5321
rect 12318 5242 12324 5276
rect 12358 5242 12364 5276
rect 12318 5197 12364 5242
rect 12318 5163 12324 5197
rect 12358 5163 12364 5197
rect 12318 5117 12364 5163
rect 12318 5083 12324 5117
rect 12358 5083 12364 5117
rect 12318 5037 12364 5083
rect 12318 5003 12324 5037
rect 12358 5003 12364 5037
rect 12318 4983 12364 5003
rect 12494 5362 12500 5396
rect 12534 5362 12586 5396
rect 12840 5426 12898 5600
tri 12898 5581 12923 5606 nw
tri 13167 5581 13192 5606 ne
rect 12840 5392 12852 5426
rect 12886 5392 12898 5426
rect 12494 5324 12586 5362
rect 12494 5290 12500 5324
rect 12534 5290 12586 5324
rect 12494 5252 12586 5290
rect 12494 5218 12500 5252
rect 12534 5218 12586 5252
rect 12494 5180 12586 5218
rect 12494 5146 12500 5180
rect 12534 5146 12586 5180
rect 12494 5108 12586 5146
rect 12494 5074 12500 5108
rect 12534 5074 12586 5108
rect 12494 5035 12586 5074
rect 12494 5001 12500 5035
rect 12534 5001 12586 5035
rect 12494 4989 12586 5001
rect 12670 5355 12716 5367
rect 12670 5321 12676 5355
rect 12710 5321 12716 5355
rect 12670 5276 12716 5321
rect 12670 5242 12676 5276
rect 12710 5242 12716 5276
rect 12670 5197 12716 5242
rect 12670 5163 12676 5197
rect 12710 5163 12716 5197
rect 12670 5117 12716 5163
rect 12670 5083 12676 5117
rect 12710 5083 12716 5117
rect 12670 5037 12716 5083
rect 12670 5003 12676 5037
rect 12710 5003 12716 5037
tri 12364 4983 12367 4986 sw
tri 12667 4983 12670 4986 se
rect 12670 4983 12716 5003
rect 12840 5348 12898 5392
rect 13192 5426 13250 5606
rect 13192 5392 13205 5426
rect 13239 5392 13250 5426
rect 12840 5314 12852 5348
rect 12886 5314 12898 5348
rect 12840 5270 12898 5314
rect 12840 5236 12852 5270
rect 12886 5236 12898 5270
rect 12840 5192 12898 5236
rect 12840 5158 12852 5192
rect 12886 5158 12898 5192
rect 12840 5114 12898 5158
rect 12840 5080 12852 5114
rect 12886 5080 12898 5114
rect 12840 5035 12898 5080
rect 12840 5001 12852 5035
rect 12886 5001 12898 5035
rect 12840 4989 12898 5001
rect 13022 5355 13068 5367
rect 13022 5321 13028 5355
rect 13062 5321 13068 5355
rect 13022 5276 13068 5321
rect 13022 5242 13028 5276
rect 13062 5242 13068 5276
rect 13022 5197 13068 5242
rect 13022 5163 13028 5197
rect 13062 5163 13068 5197
rect 13022 5117 13068 5163
rect 13022 5083 13028 5117
rect 13062 5083 13068 5117
rect 13022 5037 13068 5083
rect 13022 5003 13028 5037
rect 13062 5003 13068 5037
tri 12716 4983 12719 4986 sw
tri 13019 4983 13022 4986 se
rect 13022 4983 13068 5003
rect 13192 5348 13250 5392
rect 13192 5314 13205 5348
rect 13239 5314 13250 5348
rect 13192 5270 13250 5314
rect 13192 5236 13205 5270
rect 13239 5236 13250 5270
rect 13192 5192 13250 5236
rect 13192 5158 13205 5192
rect 13239 5158 13250 5192
rect 13192 5114 13250 5158
rect 13192 5080 13205 5114
rect 13239 5080 13250 5114
rect 13192 5035 13250 5080
rect 13192 5001 13205 5035
rect 13239 5001 13250 5035
rect 13192 4989 13250 5001
rect 13360 5640 13536 5679
rect 13360 5606 13496 5640
rect 13530 5606 13536 5640
rect 13360 5567 13536 5606
rect 13360 5533 13496 5567
rect 13530 5533 13536 5567
rect 13360 5494 13536 5533
rect 13360 5460 13496 5494
rect 13530 5460 13536 5494
rect 13360 5421 13536 5460
rect 13360 5387 13496 5421
rect 13530 5387 13536 5421
rect 13360 5355 13536 5387
rect 13360 5321 13380 5355
rect 13414 5348 13536 5355
rect 13414 5321 13496 5348
rect 13360 5314 13496 5321
rect 13530 5314 13536 5348
rect 13360 5276 13536 5314
rect 13360 5242 13380 5276
rect 13414 5275 13536 5276
rect 13414 5242 13496 5275
rect 13360 5241 13496 5242
rect 13530 5241 13536 5275
rect 13360 5202 13536 5241
rect 13360 5197 13496 5202
rect 13360 5163 13380 5197
rect 13414 5168 13496 5197
rect 13530 5168 13536 5202
rect 13414 5163 13536 5168
rect 13360 5129 13536 5163
rect 13360 5117 13496 5129
rect 13360 5083 13380 5117
rect 13414 5095 13496 5117
rect 13530 5095 13536 5129
rect 13414 5083 13536 5095
rect 13360 5056 13536 5083
rect 13360 5037 13496 5056
rect 13360 5003 13380 5037
rect 13414 5022 13496 5037
rect 13530 5022 13536 5056
rect 13414 5003 13536 5022
tri 13068 4983 13071 4986 sw
tri 13357 4983 13360 4986 se
rect 13360 4983 13536 5003
rect 12318 4961 12367 4983
tri 12367 4961 12389 4983 sw
tri 12645 4961 12667 4983 se
rect 12667 4961 12719 4983
tri 12719 4961 12741 4983 sw
tri 12997 4961 13019 4983 se
rect 13019 4961 13071 4983
tri 13071 4961 13093 4983 sw
tri 13335 4961 13357 4983 se
rect 13357 4961 13496 4983
rect 12318 4957 13496 4961
rect 12318 4923 12324 4957
rect 12358 4923 12676 4957
rect 12710 4923 13028 4957
rect 13062 4923 13380 4957
rect 13414 4949 13496 4957
rect 13530 4949 13536 4983
rect 13414 4923 13536 4949
rect 12318 4910 13536 4923
rect 12318 4877 13496 4910
rect 12318 4843 12324 4877
rect 12358 4843 12676 4877
rect 12710 4843 13028 4877
rect 13062 4843 13380 4877
rect 13414 4876 13496 4877
rect 13530 4876 13536 4910
rect 13414 4843 13536 4876
rect 12318 4837 13536 4843
rect 12318 4831 13496 4837
tri 13335 4806 13360 4831 ne
tri 11944 4803 11947 4806 se
rect 11947 4803 12012 4806
tri 11941 4800 11944 4803 se
rect 11944 4800 12012 4803
rect 8469 4784 8543 4785
rect 8405 4764 8543 4784
tri 8543 4764 8564 4785 nw
tri 10192 4764 10213 4785 ne
rect 10213 4764 10432 4785
rect 8405 4754 8527 4764
rect 7321 4753 8527 4754
rect 7281 4748 8527 4753
tri 8527 4748 8543 4764 nw
tri 10213 4757 10220 4764 ne
rect 10220 4757 10432 4764
rect 8703 4748 8754 4757
rect 8806 4748 8820 4757
rect 7281 4714 7327 4748
tri 7327 4723 7352 4748 nw
rect 7281 4680 7287 4714
rect 7321 4680 7327 4714
rect 7281 4641 7327 4680
rect 7281 4607 7287 4641
rect 7321 4607 7327 4641
rect 7281 4568 7327 4607
rect 7281 4534 7287 4568
rect 7321 4534 7327 4568
rect 7281 4495 7327 4534
rect 7281 4461 7287 4495
rect 7321 4461 7327 4495
rect 7281 4422 7327 4461
rect 7281 4388 7287 4422
rect 7321 4388 7327 4422
rect 7281 4349 7327 4388
rect 7281 4315 7287 4349
rect 7321 4315 7327 4349
rect 7281 4276 7327 4315
rect 7281 4242 7287 4276
rect 7321 4242 7327 4276
tri 7091 4214 7094 4217 sw
rect 7042 4208 7094 4214
rect 7042 4142 7094 4156
rect 7042 4084 7094 4090
rect 7281 4203 7327 4242
rect 7281 4169 7287 4203
rect 7321 4169 7327 4203
rect 7281 4130 7327 4169
rect 7281 4096 7287 4130
rect 7321 4096 7327 4130
rect 7281 4084 7327 4096
rect 7397 4708 7953 4720
rect 7397 4674 7403 4708
rect 7437 4674 7913 4708
rect 7947 4674 7953 4708
rect 8703 4714 8715 4748
rect 8749 4714 8754 4748
rect 8703 4705 8754 4714
rect 8806 4705 8820 4714
rect 8872 4705 8878 4757
rect 8906 4748 9361 4754
rect 8906 4714 8918 4748
rect 8952 4714 8991 4748
rect 9025 4714 9063 4748
rect 9097 4714 9135 4748
rect 9169 4714 9207 4748
rect 9241 4714 9279 4748
rect 9313 4714 9351 4748
rect 8906 4708 9361 4714
tri 9349 4705 9352 4708 ne
rect 9352 4705 9361 4708
tri 9352 4702 9355 4705 ne
rect 9355 4702 9361 4705
rect 9413 4702 9427 4754
rect 9479 4702 9485 4754
rect 9545 4745 9591 4757
rect 9545 4711 9551 4745
rect 9585 4711 9591 4745
tri 9524 4676 9545 4697 se
rect 9545 4676 9591 4711
rect 7397 4671 7465 4674
tri 7465 4671 7468 4674 nw
tri 7866 4671 7869 4674 ne
rect 7869 4671 7953 4674
tri 7953 4671 7958 4676 sw
tri 9520 4672 9524 4676 se
rect 9524 4672 9591 4676
rect 7397 4658 7452 4671
tri 7452 4658 7465 4671 nw
tri 7869 4658 7882 4671 ne
rect 7882 4658 7958 4671
tri 7958 4658 7971 4671 sw
rect 7397 4636 7443 4658
tri 7443 4649 7452 4658 nw
tri 7882 4649 7891 4658 ne
rect 7891 4651 7971 4658
tri 7971 4651 7978 4658 sw
rect 7891 4649 7913 4651
tri 7891 4646 7894 4649 ne
rect 7894 4646 7913 4649
rect 7397 4602 7403 4636
rect 7437 4602 7443 4636
rect 7397 4564 7443 4602
rect 7397 4530 7403 4564
rect 7437 4530 7443 4564
rect 7397 4492 7443 4530
rect 7397 4458 7403 4492
rect 7437 4458 7443 4492
rect 7397 4420 7443 4458
rect 7397 4386 7403 4420
rect 7437 4386 7443 4420
rect 7397 4348 7443 4386
rect 7397 4314 7403 4348
rect 7437 4314 7443 4348
rect 7397 4276 7443 4314
rect 7397 4242 7403 4276
rect 7437 4242 7443 4276
rect 7397 4203 7443 4242
rect 7397 4169 7403 4203
rect 7437 4169 7443 4203
rect 7397 4130 7443 4169
rect 7397 4096 7403 4130
rect 7437 4096 7443 4130
rect 7397 4084 7443 4096
rect 7583 4640 7773 4646
tri 7894 4642 7898 4646 ne
rect 7898 4642 7913 4646
rect 7583 4634 7592 4640
rect 7644 4634 7656 4640
rect 7708 4634 7720 4640
rect 7583 4096 7589 4634
rect 7772 4588 7773 4640
tri 7898 4636 7904 4642 ne
rect 7904 4636 7913 4642
tri 7904 4633 7907 4636 ne
rect 7767 4569 7773 4588
rect 7772 4517 7773 4569
rect 7767 4498 7773 4517
rect 7772 4446 7773 4498
rect 7767 4427 7773 4446
rect 7772 4375 7773 4427
rect 7767 4356 7773 4375
rect 7772 4304 7773 4356
rect 7767 4285 7773 4304
rect 7772 4233 7773 4285
rect 7767 4214 7773 4233
rect 7772 4162 7773 4214
rect 7767 4142 7773 4162
rect 7583 4090 7592 4096
rect 7644 4090 7656 4096
rect 7708 4090 7720 4096
rect 7772 4090 7773 4142
rect 7583 4084 7773 4090
rect 7907 4599 7913 4636
rect 7965 4599 7979 4651
rect 8031 4642 8045 4651
rect 8097 4642 8111 4651
rect 8163 4648 8169 4651
tri 8169 4648 8172 4651 sw
rect 8163 4642 8559 4648
rect 8097 4608 8110 4642
rect 8163 4608 8191 4642
rect 8225 4608 8272 4642
rect 8306 4608 8353 4642
rect 8387 4608 8433 4642
rect 8467 4608 8513 4642
rect 8547 4608 8559 4642
rect 8986 4620 8992 4672
rect 9044 4620 9056 4672
rect 9108 4620 9121 4672
rect 9173 4620 9186 4672
rect 9238 4658 9591 4672
rect 9238 4624 9551 4658
rect 9585 4624 9591 4658
rect 9238 4620 9591 4624
rect 8031 4599 8045 4608
rect 8097 4599 8111 4608
rect 8163 4602 8559 4608
tri 9520 4602 9538 4620 ne
rect 9538 4602 9591 4620
rect 8163 4599 8169 4602
tri 8169 4599 8172 4602 nw
tri 9538 4599 9541 4602 ne
rect 9541 4599 9591 4602
rect 7907 4597 7976 4599
tri 7976 4597 7978 4599 nw
tri 9541 4597 9543 4599 ne
rect 9543 4597 9591 4599
rect 7907 4584 7963 4597
tri 7963 4584 7976 4597 nw
tri 9543 4595 9545 4597 ne
rect 7907 4564 7953 4584
tri 7953 4574 7963 4584 nw
rect 7907 4530 7913 4564
rect 7947 4530 7953 4564
rect 7907 4492 7953 4530
rect 8828 4526 8834 4578
rect 8886 4572 8900 4578
rect 8952 4572 9397 4578
rect 8982 4538 9029 4572
rect 9063 4538 9110 4572
rect 9144 4538 9191 4572
rect 9225 4538 9271 4572
rect 9305 4538 9351 4572
rect 9385 4538 9397 4572
rect 8886 4526 8900 4538
rect 8952 4532 9397 4538
rect 9545 4571 9591 4597
rect 9545 4537 9551 4571
rect 9585 4537 9591 4571
rect 8952 4526 8958 4532
tri 8958 4526 8964 4532 nw
rect 9545 4525 9591 4537
rect 9693 4751 9918 4757
rect 9745 4745 9757 4751
rect 9809 4745 9821 4751
rect 9873 4745 9918 4751
rect 9873 4711 9878 4745
rect 9912 4711 9918 4745
tri 10220 4742 10235 4757 ne
rect 10235 4742 10432 4757
rect 11686 4748 11692 4800
rect 11744 4748 11756 4800
rect 11808 4788 12012 4800
rect 11808 4764 11988 4788
tri 11988 4764 12012 4788 nw
rect 13360 4803 13496 4831
rect 13530 4803 13536 4837
rect 13360 4764 13536 4803
rect 11808 4748 11972 4764
tri 11972 4748 11988 4764 nw
tri 10235 4730 10247 4742 ne
rect 10247 4736 10432 4742
rect 10247 4730 10380 4736
rect 9745 4699 9757 4711
rect 9809 4699 9821 4711
rect 9873 4699 9918 4711
tri 10247 4705 10272 4730 ne
rect 10272 4705 10380 4730
rect 9693 4667 9918 4699
tri 10272 4671 10306 4705 ne
rect 10306 4684 10380 4705
tri 10432 4730 10444 4742 sw
rect 13360 4730 13496 4764
rect 13530 4730 13536 4764
rect 10432 4717 10444 4730
tri 10444 4717 10457 4730 sw
rect 10432 4684 10523 4717
rect 10525 4716 10561 4717
rect 10306 4671 10523 4684
rect 9745 4658 9757 4667
rect 9809 4658 9821 4667
rect 9873 4658 9918 4667
rect 9873 4624 9878 4658
rect 9912 4624 9918 4658
tri 10306 4657 10320 4671 ne
rect 10320 4670 10523 4671
rect 10320 4657 10380 4670
tri 10320 4633 10344 4657 ne
rect 10344 4633 10380 4657
rect 9745 4615 9757 4624
rect 9809 4615 9821 4624
rect 9873 4615 9918 4624
rect 9693 4583 9918 4615
tri 10344 4612 10365 4633 ne
rect 10365 4618 10380 4633
rect 10432 4618 10523 4670
rect 10365 4612 10523 4618
tri 10365 4599 10378 4612 ne
rect 10378 4599 10523 4612
tri 10378 4597 10380 4599 ne
rect 10380 4597 10523 4599
tri 10380 4587 10390 4597 ne
rect 10390 4587 10523 4597
rect 10524 4588 10562 4716
rect 10563 4705 13150 4717
rect 10563 4671 10614 4705
rect 10648 4671 10926 4705
rect 10960 4671 11238 4705
rect 11272 4671 11550 4705
rect 11584 4671 11862 4705
rect 11896 4671 12174 4705
rect 12208 4671 12486 4705
rect 12520 4671 12798 4705
rect 12832 4671 13110 4705
rect 13144 4671 13150 4705
rect 10563 4633 13150 4671
rect 10563 4599 10614 4633
rect 10648 4599 10926 4633
rect 10960 4599 11238 4633
rect 11272 4599 11550 4633
rect 11584 4599 11862 4633
rect 11896 4599 12174 4633
rect 12208 4599 12486 4633
rect 12520 4599 12798 4633
rect 12832 4631 13150 4633
rect 12832 4599 13110 4631
rect 10563 4597 13110 4599
rect 13144 4597 13150 4631
rect 10525 4587 10561 4588
rect 10563 4587 13150 4597
tri 10583 4584 10586 4587 ne
rect 10586 4584 10676 4587
tri 10676 4584 10679 4587 nw
tri 10895 4584 10898 4587 ne
rect 10898 4584 10988 4587
tri 10988 4584 10991 4587 nw
tri 11207 4584 11210 4587 ne
rect 11210 4584 11300 4587
tri 11300 4584 11303 4587 nw
tri 11519 4584 11522 4587 ne
rect 11522 4584 11612 4587
tri 11612 4584 11615 4587 nw
tri 11831 4584 11834 4587 ne
rect 11834 4584 11924 4587
tri 11924 4584 11927 4587 nw
tri 12143 4584 12146 4587 ne
rect 12146 4584 12236 4587
tri 12236 4584 12239 4587 nw
tri 12455 4584 12458 4587 ne
rect 12458 4584 12548 4587
tri 12548 4584 12551 4587 nw
tri 12767 4584 12770 4587 ne
rect 12770 4584 12860 4587
tri 12860 4584 12863 4587 nw
tri 13079 4584 13082 4587 ne
rect 13082 4584 13150 4587
rect 9745 4571 9757 4583
rect 9809 4571 9821 4583
rect 9873 4571 9918 4583
tri 10586 4581 10589 4584 ne
rect 10589 4581 10654 4584
rect 9873 4537 9878 4571
rect 9912 4537 9918 4571
rect 9745 4531 9757 4537
rect 9809 4531 9821 4537
rect 9873 4531 9918 4537
rect 9693 4525 9918 4531
rect 10220 4575 10272 4581
tri 10589 4562 10608 4581 ne
tri 10211 4513 10220 4522 se
rect 10220 4513 10272 4523
tri 10209 4511 10211 4513 se
rect 10211 4511 10272 4513
tri 10195 4497 10209 4511 se
rect 10209 4509 10272 4511
rect 10209 4497 10220 4509
rect 7907 4458 7913 4492
rect 7947 4458 7953 4492
rect 7907 4420 7953 4458
rect 7907 4386 7913 4420
rect 7947 4386 7953 4420
rect 8668 4485 10220 4497
rect 8668 4451 8674 4485
rect 8708 4457 10220 4485
rect 8708 4451 10272 4457
rect 10608 4560 10654 4581
tri 10654 4562 10676 4584 nw
tri 10898 4562 10920 4584 ne
rect 10608 4526 10614 4560
rect 10648 4526 10654 4560
rect 10920 4560 10966 4584
tri 10966 4562 10988 4584 nw
tri 11210 4562 11232 4584 ne
rect 10608 4487 10654 4526
rect 10608 4453 10614 4487
rect 10648 4453 10654 4487
rect 8668 4441 8729 4451
tri 8729 4441 8739 4451 nw
rect 8668 4438 8726 4441
tri 8726 4438 8729 4441 nw
rect 8668 4413 8714 4438
tri 8714 4426 8726 4438 nw
tri 8506 4392 8509 4395 se
rect 8509 4392 8515 4395
rect 7907 4348 7953 4386
rect 7907 4314 7913 4348
rect 7947 4314 7953 4348
rect 8017 4386 8515 4392
rect 8567 4386 8582 4395
rect 8017 4352 8029 4386
rect 8063 4352 8104 4386
rect 8138 4352 8179 4386
rect 8213 4352 8254 4386
rect 8288 4352 8328 4386
rect 8362 4352 8402 4386
rect 8436 4352 8476 4386
rect 8510 4352 8515 4386
rect 8017 4346 8515 4352
tri 8506 4343 8509 4346 ne
rect 8509 4343 8515 4346
rect 8567 4343 8582 4352
rect 8634 4343 8640 4395
rect 8668 4379 8674 4413
rect 8708 4379 8714 4413
rect 8668 4367 8714 4379
rect 8855 4416 9361 4422
rect 8855 4382 8867 4416
rect 8901 4382 8948 4416
rect 8982 4382 9029 4416
rect 9063 4382 9110 4416
rect 9144 4382 9191 4416
rect 9225 4382 9271 4416
rect 9305 4382 9351 4416
rect 8855 4376 9361 4382
tri 9349 4370 9355 4376 ne
rect 9355 4370 9361 4376
rect 9413 4370 9427 4422
rect 9479 4370 9485 4422
rect 9693 4417 9918 4423
rect 9745 4411 9757 4417
rect 9809 4411 9821 4417
rect 9873 4411 9918 4417
rect 9873 4377 9878 4411
rect 9912 4377 9918 4411
rect 9745 4365 9757 4377
rect 9809 4365 9821 4377
rect 9873 4365 9918 4377
rect 9693 4349 9918 4365
rect 9745 4317 9757 4349
rect 9809 4317 9821 4349
rect 9873 4317 9918 4349
rect 7907 4276 7953 4314
rect 8855 4306 9361 4312
rect 7907 4242 7913 4276
rect 7947 4242 7953 4276
rect 7907 4203 7953 4242
rect 8017 4276 8623 4282
rect 8017 4242 8029 4276
rect 8063 4242 8104 4276
rect 8138 4242 8179 4276
rect 8213 4242 8254 4276
rect 8288 4242 8328 4276
rect 8362 4242 8402 4276
rect 8436 4242 8476 4276
rect 8510 4242 8550 4276
rect 8584 4272 8623 4276
tri 8623 4272 8633 4282 sw
rect 8855 4272 8867 4306
rect 8901 4272 8948 4306
rect 8982 4272 9029 4306
rect 9063 4272 9110 4306
rect 9144 4272 9191 4306
rect 9225 4272 9271 4306
rect 9305 4272 9351 4306
rect 8584 4258 8633 4272
tri 8633 4258 8647 4272 sw
rect 8855 4266 9361 4272
tri 9349 4260 9355 4266 ne
rect 9355 4260 9361 4266
rect 9413 4260 9427 4312
rect 9479 4260 9485 4312
rect 9522 4310 9574 4316
rect 8584 4256 8647 4258
tri 8647 4256 8649 4258 sw
tri 9521 4256 9522 4257 se
rect 9522 4256 9574 4258
rect 8584 4242 8649 4256
rect 8017 4236 8649 4242
tri 8603 4223 8616 4236 ne
rect 8616 4232 8649 4236
tri 8649 4232 8673 4256 sw
tri 9497 4232 9521 4256 se
rect 9521 4244 9574 4256
rect 9521 4232 9522 4244
rect 8616 4223 9522 4232
tri 8616 4216 8623 4223 ne
rect 8623 4216 9522 4223
rect 7907 4169 7913 4203
rect 7947 4169 7953 4203
tri 8623 4189 8650 4216 ne
rect 8650 4192 9522 4216
rect 8650 4189 9574 4192
tri 8650 4186 8653 4189 ne
rect 8653 4186 9574 4189
rect 9873 4297 9878 4317
rect 9693 4283 9734 4297
rect 9768 4283 9806 4297
rect 9840 4283 9878 4297
rect 9912 4283 9918 4317
rect 10608 4414 10654 4453
rect 10608 4380 10614 4414
rect 10648 4380 10654 4414
rect 10608 4341 10654 4380
rect 10608 4307 10614 4341
rect 10648 4307 10654 4341
rect 10608 4295 10654 4307
rect 10764 4547 10810 4559
rect 10764 4513 10770 4547
rect 10804 4513 10810 4547
rect 10764 4475 10810 4513
rect 10764 4441 10770 4475
rect 10804 4441 10810 4475
rect 10764 4402 10810 4441
rect 10764 4368 10770 4402
rect 10804 4368 10810 4402
rect 10764 4329 10810 4368
rect 10764 4295 10770 4329
rect 10804 4295 10810 4329
rect 10920 4526 10926 4560
rect 10960 4526 10966 4560
rect 11232 4560 11278 4584
tri 11278 4562 11300 4584 nw
tri 11522 4562 11544 4584 ne
rect 10920 4487 10966 4526
rect 10920 4453 10926 4487
rect 10960 4453 10966 4487
rect 10920 4414 10966 4453
rect 10920 4380 10926 4414
rect 10960 4380 10966 4414
rect 10920 4341 10966 4380
rect 10920 4307 10926 4341
rect 10960 4307 10966 4341
rect 10920 4295 10966 4307
rect 11076 4547 11122 4559
rect 11076 4513 11082 4547
rect 11116 4513 11122 4547
rect 11076 4475 11122 4513
rect 11076 4441 11082 4475
rect 11116 4441 11122 4475
rect 11076 4402 11122 4441
rect 11076 4368 11082 4402
rect 11116 4368 11122 4402
rect 11076 4329 11122 4368
rect 11076 4295 11082 4329
rect 11116 4295 11122 4329
rect 11232 4526 11238 4560
rect 11272 4526 11278 4560
rect 11544 4560 11590 4584
tri 11590 4562 11612 4584 nw
tri 11834 4562 11856 4584 ne
rect 11232 4487 11278 4526
rect 11232 4453 11238 4487
rect 11272 4453 11278 4487
rect 11232 4414 11278 4453
rect 11232 4380 11238 4414
rect 11272 4380 11278 4414
rect 11232 4341 11278 4380
rect 11232 4307 11238 4341
rect 11272 4307 11278 4341
rect 11232 4295 11278 4307
rect 11388 4547 11434 4559
rect 11388 4513 11394 4547
rect 11428 4513 11434 4547
rect 11388 4475 11434 4513
rect 11388 4441 11394 4475
rect 11428 4441 11434 4475
rect 11388 4402 11434 4441
rect 11388 4368 11394 4402
rect 11428 4368 11434 4402
rect 11388 4329 11434 4368
rect 11388 4295 11394 4329
rect 11428 4295 11434 4329
rect 11544 4526 11550 4560
rect 11584 4526 11590 4560
rect 11856 4560 11902 4584
tri 11902 4562 11924 4584 nw
tri 12146 4562 12168 4584 ne
rect 11544 4487 11590 4526
rect 11544 4453 11550 4487
rect 11584 4453 11590 4487
rect 11544 4414 11590 4453
rect 11544 4380 11550 4414
rect 11584 4380 11590 4414
rect 11544 4341 11590 4380
rect 11544 4307 11550 4341
rect 11584 4307 11590 4341
rect 11544 4295 11590 4307
rect 11700 4547 11746 4559
rect 11700 4513 11706 4547
rect 11740 4513 11746 4547
rect 11700 4475 11746 4513
rect 11700 4441 11706 4475
rect 11740 4441 11746 4475
rect 11700 4402 11746 4441
rect 11700 4368 11706 4402
rect 11740 4368 11746 4402
rect 11700 4329 11746 4368
rect 11700 4295 11706 4329
rect 11740 4295 11746 4329
rect 11856 4526 11862 4560
rect 11896 4526 11902 4560
rect 12168 4560 12214 4584
tri 12214 4562 12236 4584 nw
tri 12458 4562 12480 4584 ne
rect 11856 4487 11902 4526
rect 11856 4453 11862 4487
rect 11896 4453 11902 4487
rect 11856 4414 11902 4453
rect 11856 4380 11862 4414
rect 11896 4380 11902 4414
rect 11856 4341 11902 4380
rect 11856 4307 11862 4341
rect 11896 4307 11902 4341
rect 11856 4295 11902 4307
rect 12012 4547 12058 4559
rect 12012 4513 12018 4547
rect 12052 4513 12058 4547
rect 12012 4475 12058 4513
rect 12012 4441 12018 4475
rect 12052 4441 12058 4475
rect 12012 4402 12058 4441
rect 12012 4368 12018 4402
rect 12052 4368 12058 4402
rect 12012 4329 12058 4368
rect 12012 4295 12018 4329
rect 12052 4295 12058 4329
rect 12168 4526 12174 4560
rect 12208 4526 12214 4560
rect 12480 4560 12526 4584
tri 12526 4562 12548 4584 nw
tri 12770 4562 12792 4584 ne
rect 12168 4487 12214 4526
rect 12168 4453 12174 4487
rect 12208 4453 12214 4487
rect 12168 4414 12214 4453
rect 12168 4380 12174 4414
rect 12208 4380 12214 4414
rect 12168 4341 12214 4380
rect 12168 4307 12174 4341
rect 12208 4307 12214 4341
rect 12168 4295 12214 4307
rect 12324 4547 12370 4559
rect 12324 4513 12330 4547
rect 12364 4513 12370 4547
rect 12324 4475 12370 4513
rect 12324 4441 12330 4475
rect 12364 4441 12370 4475
rect 12324 4402 12370 4441
rect 12324 4368 12330 4402
rect 12364 4368 12370 4402
rect 12324 4329 12370 4368
rect 12324 4295 12330 4329
rect 12364 4295 12370 4329
rect 12480 4526 12486 4560
rect 12520 4526 12526 4560
rect 12792 4560 12838 4584
tri 12838 4562 12860 4584 nw
tri 13082 4562 13104 4584 ne
rect 12480 4487 12526 4526
rect 12480 4453 12486 4487
rect 12520 4453 12526 4487
rect 12480 4414 12526 4453
rect 12480 4380 12486 4414
rect 12520 4380 12526 4414
rect 12480 4341 12526 4380
rect 12480 4307 12486 4341
rect 12520 4307 12526 4341
rect 12480 4295 12526 4307
rect 12636 4547 12682 4559
rect 12636 4513 12642 4547
rect 12676 4513 12682 4547
rect 12636 4475 12682 4513
rect 12636 4441 12642 4475
rect 12676 4441 12682 4475
rect 12636 4402 12682 4441
rect 12636 4368 12642 4402
rect 12676 4368 12682 4402
rect 12636 4329 12682 4368
rect 12636 4295 12642 4329
rect 12676 4295 12682 4329
rect 12792 4526 12798 4560
rect 12832 4526 12838 4560
rect 12792 4487 12838 4526
rect 12792 4453 12798 4487
rect 12832 4453 12838 4487
rect 12792 4414 12838 4453
rect 12792 4380 12798 4414
rect 12832 4380 12838 4414
rect 12792 4341 12838 4380
rect 12792 4307 12798 4341
rect 12832 4307 12838 4341
rect 12792 4295 12838 4307
rect 12948 4547 12994 4559
rect 12948 4513 12954 4547
rect 12988 4513 12994 4547
rect 12948 4475 12994 4513
rect 12948 4441 12954 4475
rect 12988 4441 12994 4475
rect 12948 4402 12994 4441
rect 12948 4368 12954 4402
rect 12988 4368 12994 4402
rect 12948 4329 12994 4368
rect 12948 4295 12954 4329
rect 12988 4295 12994 4329
rect 9693 4280 9918 4283
rect 9745 4228 9757 4280
rect 9809 4228 9821 4280
rect 9873 4228 9918 4280
tri 10739 4267 10764 4292 se
rect 10764 4267 10810 4295
tri 10810 4267 10835 4292 sw
tri 11051 4267 11076 4292 se
rect 11076 4267 11122 4295
tri 11122 4267 11147 4292 sw
tri 11363 4267 11388 4292 se
rect 11388 4267 11434 4295
tri 11434 4267 11459 4292 sw
tri 11675 4267 11700 4292 se
rect 11700 4267 11746 4295
tri 11746 4267 11771 4292 sw
tri 11987 4267 12012 4292 se
rect 12012 4267 12058 4295
tri 12058 4267 12083 4292 sw
tri 12299 4267 12324 4292 se
rect 12324 4267 12370 4295
tri 12370 4267 12395 4292 sw
tri 12611 4267 12636 4292 se
rect 12636 4267 12682 4295
tri 12682 4267 12707 4292 sw
tri 12923 4267 12948 4292 se
rect 12948 4267 12994 4295
tri 10177 4258 10186 4267 se
rect 10186 4261 10679 4267
rect 10681 4266 10717 4267
rect 10186 4258 10300 4261
tri 10175 4256 10177 4258 se
rect 10177 4256 10300 4258
rect 9693 4223 9918 4228
rect 9693 4211 9734 4223
rect 9768 4211 9806 4223
rect 9840 4211 9878 4223
rect 9873 4189 9878 4211
rect 9912 4189 9918 4223
tri 10141 4222 10175 4256 se
rect 10175 4222 10300 4256
tri 10138 4219 10141 4222 se
rect 10141 4219 10300 4222
rect 7907 4130 7953 4169
rect 9745 4159 9757 4189
rect 9809 4159 9821 4189
rect 9873 4159 9918 4189
tri 10102 4183 10138 4219 se
rect 10138 4209 10300 4219
rect 10352 4209 10679 4261
rect 10138 4195 10679 4209
rect 10138 4183 10300 4195
rect 9693 4142 9918 4159
tri 10068 4149 10102 4183 se
rect 10102 4149 10300 4183
tri 10065 4146 10068 4149 se
rect 10068 4146 10300 4149
rect 7907 4096 7913 4130
rect 7947 4096 7953 4130
rect 7907 4084 7953 4096
rect 8585 4127 8754 4136
rect 8585 4093 8597 4127
rect 8631 4093 8669 4127
rect 8703 4093 8754 4127
rect 8585 4084 8754 4093
rect 8806 4084 8820 4136
rect 8872 4084 8878 4136
rect 8906 4130 8992 4136
rect 8906 4096 8918 4130
rect 8952 4096 8991 4130
rect 8906 4084 8992 4096
rect 9044 4084 9056 4136
rect 9108 4084 9121 4136
rect 9173 4084 9186 4136
rect 9238 4130 9397 4136
rect 9241 4096 9279 4130
rect 9313 4096 9351 4130
rect 9385 4096 9397 4130
rect 9238 4084 9397 4096
rect 9745 4130 9757 4142
rect 9809 4130 9821 4142
rect 9873 4130 9918 4142
tri 10056 4137 10065 4146 se
rect 10065 4143 10300 4146
rect 10352 4143 10679 4195
rect 10065 4137 10679 4143
rect 10680 4138 10718 4266
rect 10719 4256 12994 4267
rect 10719 4222 10770 4256
rect 10804 4222 11082 4256
rect 11116 4222 11394 4256
rect 11428 4222 11706 4256
rect 11740 4222 12018 4256
rect 12052 4222 12330 4256
rect 12364 4222 12642 4256
rect 12676 4222 12954 4256
rect 12988 4222 12994 4256
rect 10719 4183 12994 4222
rect 10719 4149 10770 4183
rect 10804 4149 11082 4183
rect 11116 4149 11394 4183
rect 11428 4149 11706 4183
rect 11740 4149 12018 4183
rect 12052 4149 12330 4183
rect 12364 4149 12642 4183
rect 12676 4149 12954 4183
rect 12988 4149 12994 4183
rect 10681 4137 10717 4138
rect 10719 4137 12994 4149
rect 13104 4557 13150 4584
rect 13104 4523 13110 4557
rect 13144 4523 13150 4557
rect 13104 4483 13150 4523
rect 13104 4449 13110 4483
rect 13144 4449 13150 4483
rect 13104 4408 13150 4449
rect 13104 4374 13110 4408
rect 13144 4374 13150 4408
rect 13104 4333 13150 4374
rect 13104 4299 13110 4333
rect 13144 4299 13150 4333
rect 13104 4258 13150 4299
rect 13104 4224 13110 4258
rect 13144 4224 13150 4258
rect 13104 4183 13150 4224
rect 13104 4149 13110 4183
rect 13144 4149 13150 4183
rect 13104 4137 13150 4149
rect 13360 4691 13536 4730
rect 13360 4657 13496 4691
rect 13530 4657 13536 4691
rect 13360 4618 13536 4657
rect 13360 4584 13496 4618
rect 13530 4584 13536 4618
rect 13360 4545 13536 4584
rect 13360 4511 13496 4545
rect 13530 4511 13536 4545
rect 13360 4472 13536 4511
rect 13360 4438 13496 4472
rect 13530 4438 13536 4472
rect 13360 4399 13536 4438
rect 13360 4365 13496 4399
rect 13530 4365 13536 4399
rect 13360 4326 13536 4365
rect 13360 4292 13496 4326
rect 13530 4292 13536 4326
rect 13360 4253 13536 4292
rect 13360 4219 13496 4253
rect 13530 4219 13536 4253
rect 13360 4180 13536 4219
rect 13360 4146 13496 4180
rect 13530 4146 13536 4180
rect 9873 4096 9878 4130
rect 9912 4096 9918 4130
tri 10026 4107 10056 4137 se
rect 10056 4107 10123 4137
tri 10123 4107 10153 4137 nw
rect 13360 4107 13536 4146
rect 9745 4090 9757 4096
rect 9809 4090 9821 4096
rect 9873 4090 9918 4096
rect 9693 4084 9918 4090
tri 10003 4084 10026 4107 se
rect 10026 4084 10089 4107
rect 6699 4048 6705 4082
rect 6739 4073 6745 4082
tri 10000 4081 10003 4084 se
rect 10003 4081 10089 4084
tri 6745 4073 6753 4081 sw
tri 9992 4073 10000 4081 se
rect 10000 4073 10089 4081
tri 10089 4073 10123 4107 nw
rect 6739 4071 6753 4073
tri 6753 4071 6755 4073 sw
tri 9990 4071 9992 4073 se
rect 9992 4071 10087 4073
tri 10087 4071 10089 4073 nw
rect 6739 4056 6755 4071
tri 6755 4056 6770 4071 sw
tri 9975 4056 9990 4071 se
rect 9990 4056 10072 4071
tri 10072 4056 10087 4071 nw
rect 6739 4048 7167 4056
rect 6699 4010 7167 4048
rect 6699 3976 6705 4010
rect 6739 4004 7167 4010
rect 7219 4004 7233 4056
rect 7285 4004 7299 4056
rect 7351 4037 10053 4056
tri 10053 4037 10072 4056 nw
rect 7351 4016 10011 4037
rect 7351 4004 8508 4016
rect 6739 3992 8508 4004
rect 6739 3976 7167 3992
rect 6699 3964 7167 3976
rect 6555 3929 6561 3963
rect 6595 3929 6601 3963
tri 7137 3961 7140 3964 ne
rect 7140 3961 7167 3964
tri 7140 3954 7147 3961 ne
rect 7147 3954 7167 3961
tri 7147 3940 7161 3954 ne
rect 7161 3940 7167 3954
rect 7219 3940 7233 3992
rect 7285 3940 7299 3992
rect 7351 3964 8508 3992
rect 8560 3964 8574 4016
rect 8626 3995 10011 4016
tri 10011 3995 10053 4037 nw
rect 10548 4029 10554 4081
rect 10606 4029 10618 4081
rect 10670 4071 13105 4081
rect 10697 4037 10735 4071
rect 10769 4037 10807 4071
rect 10841 4037 10879 4071
rect 10913 4037 10951 4071
rect 10985 4037 11023 4071
rect 11057 4037 11095 4071
rect 11129 4037 11167 4071
rect 11201 4037 11239 4071
rect 11273 4037 11311 4071
rect 11345 4037 11383 4071
rect 11417 4037 11455 4071
rect 11489 4037 11527 4071
rect 11561 4037 11599 4071
rect 11633 4037 11672 4071
rect 11706 4037 11745 4071
rect 11779 4037 11818 4071
rect 11852 4037 11891 4071
rect 11925 4037 11964 4071
rect 11998 4037 12037 4071
rect 12071 4037 12110 4071
rect 12144 4037 12183 4071
rect 12217 4037 12256 4071
rect 12290 4037 12329 4071
rect 12363 4037 12402 4071
rect 12436 4037 12475 4071
rect 12509 4037 12548 4071
rect 12582 4037 12621 4071
rect 12655 4037 12694 4071
rect 12728 4037 12767 4071
rect 12801 4037 12840 4071
rect 12874 4037 12913 4071
rect 12947 4037 12986 4071
rect 13020 4037 13059 4071
rect 13093 4037 13105 4071
rect 10670 4029 13105 4037
rect 13360 4073 13496 4107
rect 13530 4073 13536 4107
tri 13335 4001 13360 4026 se
rect 13360 4001 13536 4073
tri 10092 3995 10098 4001 se
rect 10098 3995 13536 4001
rect 8626 3988 10004 3995
tri 10004 3988 10011 3995 nw
tri 10085 3988 10092 3995 se
rect 10092 3988 10510 3995
rect 8626 3964 8813 3988
tri 8813 3964 8837 3988 nw
tri 10061 3964 10085 3988 se
rect 10085 3964 10510 3988
rect 7351 3961 7378 3964
tri 7378 3961 7381 3964 nw
tri 10058 3961 10061 3964 se
rect 10061 3961 10510 3964
rect 10544 3961 10583 3995
rect 10617 3961 10656 3995
rect 10690 3961 10729 3995
rect 10763 3961 10802 3995
rect 10836 3961 10875 3995
rect 10909 3961 10948 3995
rect 10982 3961 11021 3995
rect 11055 3961 11094 3995
rect 11128 3961 11167 3995
rect 11201 3961 11240 3995
rect 11274 3961 11313 3995
rect 11347 3961 11386 3995
rect 11420 3961 11460 3995
rect 11494 3961 11534 3995
rect 11568 3961 11608 3995
rect 11642 3961 11682 3995
rect 11716 3961 11756 3995
rect 11790 3961 11830 3995
rect 11864 3961 11904 3995
rect 11938 3961 11978 3995
rect 12012 3961 12052 3995
rect 12086 3961 12126 3995
rect 12160 3961 12200 3995
rect 12234 3961 12274 3995
rect 12308 3961 12348 3995
rect 12382 3961 12422 3995
rect 12456 3961 12496 3995
rect 12530 3961 12570 3995
rect 12604 3961 12644 3995
rect 12678 3961 12718 3995
rect 12752 3961 12792 3995
rect 12826 3961 12866 3995
rect 12900 3961 12940 3995
rect 12974 3961 13014 3995
rect 13048 3961 13088 3995
rect 13122 3961 13162 3995
rect 13196 3961 13236 3995
rect 13270 3961 13310 3995
rect 13344 3961 13384 3995
rect 13418 3961 13458 3995
rect 13492 3961 13536 3995
rect 7351 3954 7371 3961
tri 7371 3954 7378 3961 nw
tri 10057 3960 10058 3961 se
rect 10058 3960 13536 3961
rect 8855 3954 9359 3960
rect 7351 3940 7357 3954
tri 7357 3940 7371 3954 nw
rect 6555 3889 6601 3929
rect 7397 3924 7913 3936
rect 6555 3855 6561 3889
rect 6595 3855 6601 3889
rect 6555 3815 6601 3855
rect 6852 3904 6904 3910
tri 6851 3850 6852 3851 se
rect 6852 3850 6904 3852
rect 7397 3890 7403 3924
rect 7437 3890 7913 3924
tri 6904 3850 6905 3851 sw
tri 6827 3826 6851 3850 se
rect 6851 3838 6905 3850
rect 6851 3826 6852 3838
rect 6555 3781 6561 3815
rect 6595 3781 6601 3815
rect 6555 3769 6601 3781
rect 6768 3820 6852 3826
rect 6904 3826 6905 3838
tri 6905 3826 6929 3850 sw
rect 6904 3820 7258 3826
rect 6768 3786 6780 3820
rect 6814 3786 6852 3820
rect 6904 3786 6924 3820
rect 6958 3786 6996 3820
rect 7030 3786 7068 3820
rect 7102 3786 7140 3820
rect 7174 3786 7212 3820
rect 7246 3786 7258 3820
rect 6768 3780 7258 3786
rect 7397 3815 7443 3890
tri 7443 3865 7468 3890 nw
tri 7866 3865 7891 3890 ne
rect 7891 3884 7913 3890
rect 7965 3884 7979 3936
rect 8031 3924 8045 3936
rect 8097 3924 8111 3936
rect 8163 3930 8169 3936
tri 8169 3930 8175 3936 sw
rect 8163 3924 8596 3930
rect 8097 3890 8104 3924
rect 8163 3890 8179 3924
rect 8213 3890 8254 3924
rect 8288 3890 8328 3924
rect 8362 3890 8402 3924
rect 8436 3890 8476 3924
rect 8510 3890 8550 3924
rect 8584 3890 8596 3924
rect 8031 3884 8045 3890
rect 8097 3884 8111 3890
rect 8163 3884 8596 3890
rect 8657 3924 8787 3930
rect 8657 3890 8669 3924
rect 8703 3890 8741 3924
rect 8775 3920 8787 3924
tri 8787 3920 8790 3923 sw
rect 8855 3920 8867 3954
rect 8901 3920 8948 3954
rect 8982 3920 9029 3954
rect 9063 3920 9110 3954
rect 9144 3920 9191 3954
rect 9225 3920 9271 3954
rect 9305 3920 9351 3954
rect 8775 3890 8790 3920
rect 8657 3884 8790 3890
rect 7891 3865 7953 3884
tri 7891 3862 7894 3865 ne
rect 7894 3862 7953 3865
rect 7397 3781 7403 3815
rect 7437 3781 7443 3815
rect 7397 3769 7443 3781
rect 7583 3850 7773 3862
rect 7583 3816 7589 3850
rect 7623 3827 7661 3850
rect 7695 3827 7733 3850
rect 7767 3827 7773 3850
tri 7894 3849 7907 3862 ne
rect 7583 3775 7592 3816
rect 7644 3775 7656 3827
rect 7708 3775 7720 3827
rect 7772 3775 7773 3827
rect 7583 3769 7773 3775
rect 7907 3842 7953 3862
tri 7953 3859 7978 3884 nw
tri 8766 3863 8787 3884 ne
rect 8787 3872 8790 3884
tri 8790 3872 8838 3920 sw
rect 8855 3914 9359 3920
tri 9347 3908 9353 3914 ne
rect 9353 3908 9359 3914
rect 9411 3908 9425 3960
rect 9477 3908 9483 3960
tri 10052 3955 10057 3960 se
rect 10057 3955 13536 3960
rect 9680 3949 13536 3955
rect 9732 3943 9744 3949
rect 9796 3943 9808 3949
rect 9860 3943 13536 3949
rect 9732 3897 9734 3943
rect 9680 3883 9734 3897
rect 9912 3887 13536 3943
rect 8787 3863 9278 3872
tri 8787 3859 8791 3863 ne
rect 8791 3859 9278 3863
rect 7907 3808 7913 3842
rect 7947 3808 7953 3842
tri 8791 3837 8813 3859 ne
rect 8813 3837 9278 3859
tri 8813 3831 8819 3837 ne
rect 8819 3831 9278 3837
tri 9261 3820 9272 3831 ne
rect 9272 3820 9278 3831
rect 9330 3820 9344 3872
rect 9396 3820 9402 3872
rect 9732 3837 9734 3883
rect 9912 3837 11647 3887
rect 9732 3831 9744 3837
rect 9796 3831 9808 3837
rect 9860 3831 11647 3837
rect 9680 3825 11647 3831
tri 11647 3825 11709 3887 nw
tri 11727 3825 11733 3831 se
rect 11733 3825 12450 3831
tri 11722 3820 11727 3825 se
rect 11727 3820 12450 3825
rect 7907 3760 7953 3808
tri 11689 3787 11722 3820 se
rect 11722 3787 12450 3820
tri 10959 3784 10962 3787 se
rect 10962 3784 10968 3787
rect 6527 3739 7578 3741
tri 7578 3739 7580 3741 sw
rect 6527 3726 7580 3739
tri 7580 3726 7593 3739 sw
rect 7907 3726 7913 3760
rect 7947 3726 7953 3760
rect 6527 3714 7593 3726
tri 7593 3714 7605 3726 sw
rect 6527 3695 7605 3714
rect 4971 3679 5032 3695
tri 5032 3679 5048 3695 nw
tri 7550 3679 7566 3695 ne
rect 7566 3679 7605 3695
tri 7605 3679 7640 3714 sw
rect 7907 3679 7953 3726
rect 4971 3604 5023 3679
tri 5023 3670 5032 3679 nw
tri 7566 3670 7575 3679 ne
rect 7575 3670 7640 3679
tri 7575 3665 7580 3670 ne
rect 7580 3665 7640 3670
tri 7640 3665 7654 3679 sw
tri 7580 3645 7600 3665 ne
rect 7600 3645 7654 3665
tri 7654 3645 7674 3665 sw
rect 7907 3645 7913 3679
rect 7947 3645 7953 3679
tri 7600 3638 7607 3645 ne
rect 7607 3638 7674 3645
tri 7674 3638 7681 3645 sw
tri 7607 3624 7621 3638 ne
rect 7621 3624 7681 3638
tri 5023 3604 5043 3624 sw
tri 7621 3604 7641 3624 ne
rect 7641 3604 7681 3624
tri 7681 3604 7715 3638 sw
rect 4971 3602 5043 3604
tri 5043 3602 5045 3604 sw
tri 7641 3602 7643 3604 ne
rect 7643 3602 7715 3604
tri 7715 3602 7717 3604 sw
rect 4971 3599 5045 3602
tri 5045 3599 5048 3602 sw
tri 7643 3599 7646 3602 ne
rect 7646 3599 7717 3602
rect 4971 3598 7600 3599
tri 7600 3598 7601 3599 sw
tri 7646 3598 7647 3599 ne
rect 7647 3598 7717 3599
tri 7717 3598 7721 3602 sw
rect 7907 3598 7953 3645
rect 8017 3748 8596 3754
rect 8017 3714 8029 3748
rect 8063 3714 8104 3748
rect 8138 3714 8179 3748
rect 8213 3714 8254 3748
rect 8288 3714 8328 3748
rect 8362 3714 8402 3748
rect 8436 3714 8476 3748
rect 8510 3714 8550 3748
rect 8584 3714 8596 3748
rect 8748 3732 8754 3784
rect 8806 3732 8820 3784
rect 8872 3778 10968 3784
rect 8901 3744 8948 3778
rect 8982 3744 9029 3778
rect 9063 3744 9110 3778
rect 9144 3744 9191 3778
rect 9225 3744 9271 3778
rect 9305 3744 9351 3778
rect 9385 3744 10968 3778
rect 8872 3738 10968 3744
rect 8872 3732 8878 3738
tri 8878 3732 8884 3738 nw
tri 10959 3735 10962 3738 ne
rect 10962 3735 10968 3738
rect 11020 3735 11032 3787
rect 11084 3735 11090 3787
tri 11658 3756 11689 3787 se
rect 11689 3779 12450 3787
rect 12502 3779 12516 3831
rect 12568 3779 13034 3831
rect 13086 3779 13100 3831
rect 13152 3779 13158 3831
rect 11689 3756 11733 3779
tri 11733 3756 11756 3779 nw
tri 11637 3735 11658 3756 se
tri 11634 3732 11637 3735 se
rect 11637 3732 11658 3735
tri 11631 3729 11634 3732 se
rect 11634 3729 11658 3732
rect 8017 3704 8596 3714
tri 8596 3704 8621 3729 sw
tri 11611 3709 11631 3729 se
rect 11631 3709 11658 3729
tri 10543 3704 10548 3709 se
rect 10548 3704 10554 3709
rect 8017 3657 10554 3704
rect 10606 3657 10618 3709
rect 10670 3657 10676 3709
tri 11583 3681 11611 3709 se
rect 11611 3681 11658 3709
tri 11658 3681 11733 3756 nw
tri 11559 3657 11583 3681 se
rect 8017 3638 8223 3657
rect 8017 3604 8029 3638
rect 8063 3604 8101 3638
rect 8135 3604 8173 3638
rect 8207 3604 8223 3638
rect 8017 3602 8223 3604
tri 8223 3602 8278 3657 nw
tri 11510 3608 11559 3657 se
rect 11559 3608 11583 3657
rect 8855 3602 9361 3608
rect 9413 3602 9427 3608
rect 8017 3598 8219 3602
tri 8219 3598 8223 3602 nw
rect 4971 3585 7601 3598
tri 7601 3585 7614 3598 sw
tri 7647 3591 7654 3598 ne
rect 7654 3591 7721 3598
tri 7721 3591 7728 3598 sw
tri 7654 3585 7660 3591 ne
rect 7660 3585 7728 3591
rect 4971 3564 7614 3585
tri 7614 3564 7635 3585 sw
tri 7660 3564 7681 3585 ne
rect 7681 3564 7728 3585
tri 7728 3564 7755 3591 sw
rect 7907 3564 7913 3598
rect 7947 3570 7953 3598
tri 7953 3570 7978 3595 sw
rect 7947 3564 8749 3570
rect 4971 3547 7635 3564
tri 7578 3519 7606 3547 ne
rect 7606 3545 7635 3547
tri 7635 3545 7654 3564 sw
tri 7681 3545 7700 3564 ne
rect 7700 3545 7755 3564
rect 7606 3519 7654 3545
tri 4943 3517 4945 3519 sw
tri 7606 3517 7608 3519 ne
rect 7608 3517 7654 3519
tri 7654 3517 7682 3545 sw
tri 7700 3517 7728 3545 ne
rect 7728 3517 7755 3545
tri 7755 3517 7802 3564 sw
rect 7907 3523 8749 3564
rect 8855 3568 8867 3602
rect 8901 3568 8942 3602
rect 8976 3568 9017 3602
rect 9051 3568 9092 3602
rect 9126 3568 9166 3602
rect 9200 3568 9240 3602
rect 9274 3568 9314 3602
rect 9348 3568 9361 3602
rect 9422 3568 9427 3602
rect 8855 3562 9361 3568
tri 9349 3556 9355 3562 ne
rect 9355 3556 9361 3562
rect 9413 3556 9427 3568
rect 9479 3556 9485 3608
tri 11508 3606 11510 3608 se
rect 11510 3606 11583 3608
tri 11583 3606 11658 3681 nw
rect 11794 3671 11800 3723
rect 11852 3671 11866 3723
rect 11918 3671 13843 3723
rect 11794 3659 13843 3671
rect 11794 3607 11800 3659
rect 11852 3607 11866 3659
rect 11918 3607 13843 3659
rect 13959 3607 13965 3723
tri 11458 3556 11508 3606 se
tri 11433 3531 11458 3556 se
rect 11458 3531 11508 3556
tri 11508 3531 11583 3606 nw
tri 11425 3523 11433 3531 se
rect 11433 3523 11448 3531
rect 4937 3494 4945 3517
tri 4945 3494 4968 3517 sw
tri 7608 3511 7614 3517 ne
rect 7614 3511 7682 3517
tri 7682 3511 7688 3517 sw
tri 7728 3511 7734 3517 ne
rect 7734 3511 7802 3517
tri 7614 3494 7631 3511 ne
rect 7631 3494 7688 3511
rect 357 3460 395 3488
tri 35 3454 41 3460 se
rect 41 3454 129 3460
tri 129 3454 135 3460 sw
rect 317 3454 395 3460
rect 429 3454 468 3488
rect 502 3454 541 3488
rect 575 3454 614 3488
rect 648 3454 687 3488
rect 721 3454 760 3488
rect 794 3454 833 3488
rect 867 3454 906 3488
rect 940 3454 979 3488
rect 1013 3454 1052 3488
rect 1086 3454 1125 3488
rect 1159 3454 1198 3488
rect 1232 3454 1271 3488
rect 1305 3454 1344 3488
rect 1558 3480 1563 3488
rect 1624 3480 1636 3488
rect 1690 3480 1709 3488
rect 1378 3454 1417 3480
rect 1451 3454 1490 3480
rect 1524 3454 1563 3480
rect 1597 3454 1636 3480
rect 1670 3454 1709 3480
rect 1743 3454 1782 3488
rect 1816 3454 1855 3488
rect 1889 3454 1928 3488
rect 1962 3454 2001 3488
rect 2035 3454 2074 3488
rect 2108 3454 2147 3488
rect 2181 3454 2220 3488
rect 2254 3454 2293 3488
rect 2327 3454 2366 3488
rect 2400 3454 2439 3488
rect 2473 3454 2512 3488
rect 2546 3454 2585 3488
rect 2619 3454 2658 3488
rect 2692 3454 2731 3488
rect 2765 3454 2804 3488
rect 2838 3454 2877 3488
rect 2911 3454 2950 3488
rect 2984 3454 3023 3488
rect 3057 3454 3096 3488
rect 3130 3454 3169 3488
rect 3203 3454 3242 3488
rect 3276 3454 3315 3488
rect 3349 3454 3388 3488
rect 3422 3454 3461 3488
rect 3495 3454 3534 3488
rect 3568 3454 3607 3488
rect 3641 3454 3679 3488
rect 3713 3454 3751 3488
rect 3785 3454 3823 3488
rect 3857 3454 3895 3488
rect 3929 3454 3967 3488
rect 4001 3454 4039 3488
rect 4073 3454 4111 3488
rect 4145 3454 4183 3488
rect 4217 3454 4255 3488
rect 4289 3454 4327 3488
rect 4361 3454 4399 3488
rect 4433 3454 4471 3488
rect 4505 3454 4543 3488
rect 4577 3454 4615 3488
rect 4649 3454 4687 3488
rect 4721 3454 4757 3488
rect 4937 3488 7443 3494
rect 4937 3454 4987 3488
rect 5021 3454 5061 3488
rect 5095 3454 5134 3488
rect 5168 3454 5207 3488
rect 5241 3454 5280 3488
rect 5314 3454 5353 3488
rect 5387 3454 5426 3488
rect 5460 3454 5499 3488
rect 5533 3454 5572 3488
rect 5606 3454 5645 3488
rect 5679 3454 5718 3488
rect 5752 3454 5791 3488
rect 5825 3454 5864 3488
rect 5898 3454 5937 3488
rect 5971 3454 6010 3488
rect 6044 3454 6083 3488
rect 6117 3454 6156 3488
rect 6190 3454 6229 3488
rect 6263 3454 6302 3488
rect 6336 3454 6375 3488
rect 6409 3454 6448 3488
rect 6482 3454 6521 3488
rect 6555 3454 6594 3488
rect 6628 3454 6667 3488
rect 6701 3454 6740 3488
rect 6774 3454 6813 3488
rect 6847 3454 6886 3488
rect 6920 3454 6959 3488
rect 6993 3454 7032 3488
rect 7066 3454 7105 3488
rect 7139 3454 7178 3488
rect 7212 3454 7251 3488
rect 7285 3454 7324 3488
rect 7358 3454 7397 3488
rect 7431 3454 7443 3488
tri 7631 3483 7642 3494 ne
rect 7642 3483 7688 3494
tri 7688 3483 7716 3511 sw
tri 7734 3483 7762 3511 ne
rect 7762 3483 7802 3511
tri 7802 3483 7836 3517 sw
tri 7642 3477 7648 3483 ne
rect 7648 3477 7716 3483
tri 7716 3477 7722 3483 sw
tri 7762 3477 7768 3483 ne
rect 7768 3477 7836 3483
tri 7836 3477 7842 3483 sw
tri 12 3431 35 3454 se
rect 35 3431 135 3454
tri 135 3431 158 3454 sw
rect 317 3448 7443 3454
tri 7648 3448 7677 3477 ne
rect 7677 3471 7722 3477
tri 7722 3471 7728 3477 sw
tri 7768 3471 7774 3477 ne
rect 7774 3471 7842 3477
rect 7677 3448 7728 3471
tri 7677 3437 7688 3448 ne
rect 7688 3437 7728 3448
tri 7728 3437 7762 3471 sw
tri 7774 3443 7802 3471 ne
rect 7802 3443 7842 3471
tri 7842 3443 7876 3477 sw
rect 7907 3471 7913 3523
rect 7965 3471 7979 3523
rect 8031 3471 8045 3523
rect 8097 3471 8111 3523
rect 8163 3511 8749 3523
rect 8163 3477 8377 3511
rect 8411 3477 8459 3511
rect 8493 3477 8541 3511
rect 8575 3477 8622 3511
rect 8656 3477 8703 3511
rect 8737 3477 8749 3511
rect 8163 3471 8749 3477
rect 8777 3514 11448 3523
rect 8777 3480 8789 3514
rect 8823 3480 8861 3514
rect 8895 3480 11448 3514
rect 8777 3471 11448 3480
tri 11448 3471 11508 3531 nw
rect 11980 3499 11986 3551
rect 12038 3499 12052 3551
rect 12104 3499 14029 3551
rect 11980 3487 14029 3499
tri 7802 3437 7808 3443 ne
rect 7808 3437 9450 3443
tri 7688 3431 7694 3437 ne
rect 7694 3431 7762 3437
tri 7762 3431 7768 3437 sw
tri 7808 3431 7814 3437 ne
rect 7814 3431 9450 3437
tri 3 3422 12 3431 se
rect 12 3422 158 3431
tri -31 3388 3 3422 se
rect 3 3388 68 3422
rect 102 3408 158 3422
tri 158 3408 181 3431 sw
tri 7694 3420 7705 3431 ne
rect 7705 3420 7768 3431
rect 102 3388 4320 3408
tri -46 3373 -31 3388 se
rect -31 3373 4320 3388
tri -70 3349 -46 3373 se
rect -46 3356 4320 3373
rect 4372 3356 4385 3408
rect 4437 3356 4450 3408
rect 4502 3356 4516 3408
rect 4568 3397 6598 3408
tri 6598 3397 6609 3408 sw
rect 4568 3373 6609 3397
tri 6609 3373 6633 3397 sw
rect 4568 3356 6633 3373
rect -46 3349 6633 3356
tri -104 3315 -70 3349 se
rect -70 3315 68 3349
rect 102 3344 6633 3349
rect 102 3315 4320 3344
tri -143 3276 -104 3315 se
rect -104 3292 4320 3315
rect 4372 3292 4385 3344
rect 4437 3292 4450 3344
rect 4502 3292 4516 3344
rect 4568 3339 6633 3344
tri 6633 3339 6667 3373 sw
rect 7042 3368 7048 3420
rect 7100 3368 7114 3420
rect 7166 3397 7659 3420
tri 7659 3397 7682 3420 sw
tri 7705 3397 7728 3420 ne
rect 7728 3397 7768 3420
tri 7768 3397 7802 3431 sw
tri 7814 3397 7848 3431 ne
rect 7848 3397 9450 3431
rect 7166 3391 7682 3397
tri 7682 3391 7688 3397 sw
tri 7728 3391 7734 3397 ne
rect 7734 3391 7802 3397
rect 7166 3373 7688 3391
tri 7688 3373 7706 3391 sw
tri 7734 3373 7752 3391 ne
rect 7752 3373 7802 3391
tri 7802 3373 7826 3397 sw
tri 7848 3391 7854 3397 ne
rect 7854 3391 9450 3397
rect 9502 3391 9516 3443
rect 9568 3391 9574 3443
rect 9680 3391 9686 3443
rect 9738 3391 9750 3443
rect 9802 3391 9815 3443
rect 9867 3431 11286 3443
rect 11980 3435 11986 3487
rect 12038 3435 12052 3487
rect 12104 3435 14029 3487
rect 14145 3435 14151 3551
rect 9867 3397 9900 3431
rect 9934 3397 9975 3431
rect 10009 3397 10050 3431
rect 10084 3397 10125 3431
rect 10159 3397 10200 3431
rect 10234 3397 10275 3431
rect 10309 3397 10350 3431
rect 10384 3397 10425 3431
rect 10459 3397 10500 3431
rect 10534 3397 10574 3431
rect 10608 3397 10648 3431
rect 10682 3397 10722 3431
rect 10756 3397 10796 3431
rect 10830 3397 10870 3431
rect 10904 3397 10944 3431
rect 10978 3397 11018 3431
rect 11052 3397 11092 3431
rect 11126 3397 11166 3431
rect 11200 3397 11240 3431
rect 11274 3397 11286 3431
rect 9867 3391 11286 3397
rect 12540 3373 13406 3379
rect 7166 3368 7706 3373
tri 7637 3346 7659 3368 ne
rect 7659 3357 7706 3368
tri 7706 3357 7722 3373 sw
tri 7752 3363 7762 3373 ne
rect 7762 3363 7826 3373
tri 7826 3363 7836 3373 sw
tri 7762 3357 7768 3363 ne
rect 7768 3357 8507 3363
rect 7659 3346 7722 3357
tri 7659 3340 7665 3346 ne
rect 7665 3340 7722 3346
rect 4568 3292 6667 3339
rect -104 3280 6667 3292
rect -104 3276 4320 3280
tri -177 3242 -143 3276 se
rect -143 3242 68 3276
rect 102 3242 4320 3276
tri -190 3229 -177 3242 se
rect -177 3229 4320 3242
tri -209 3210 -190 3229 se
rect -190 3228 4320 3229
rect 4372 3228 4385 3280
rect 4437 3228 4450 3280
rect 4502 3228 4516 3280
rect 4568 3263 6667 3280
tri 6667 3263 6743 3339 sw
rect 6943 3288 6949 3340
rect 7001 3288 7015 3340
rect 7067 3339 7619 3340
tri 7619 3339 7620 3340 sw
tri 7665 3339 7666 3340 ne
rect 7666 3339 7722 3340
tri 7722 3339 7740 3357 sw
tri 7768 3339 7786 3357 ne
rect 7786 3339 8507 3357
rect 7067 3323 7620 3339
tri 7620 3323 7636 3339 sw
tri 7666 3323 7682 3339 ne
rect 7682 3323 7740 3339
rect 7067 3288 7636 3323
tri 7597 3266 7619 3288 ne
rect 7619 3277 7636 3288
tri 7636 3277 7682 3323 sw
tri 7682 3283 7722 3323 ne
rect 7722 3317 7740 3323
tri 7740 3317 7762 3339 sw
tri 7786 3317 7808 3339 ne
rect 7808 3317 8507 3339
rect 7722 3283 7762 3317
tri 7762 3283 7796 3317 sw
tri 7808 3311 7814 3317 ne
rect 7814 3311 8507 3317
rect 8559 3311 8571 3363
rect 8623 3311 11508 3363
rect 11560 3311 11572 3363
rect 11624 3311 11630 3363
rect 12540 3339 12552 3373
rect 12586 3339 12629 3373
rect 12663 3339 12706 3373
rect 12740 3339 12783 3373
rect 12817 3339 12860 3373
rect 12894 3339 12938 3373
rect 12972 3339 13016 3373
rect 13050 3339 13094 3373
rect 13128 3339 13172 3373
rect 13206 3339 13250 3373
rect 13284 3339 13328 3373
rect 13362 3339 13406 3373
rect 12540 3333 13406 3339
tri 13335 3311 13357 3333 ne
rect 13357 3311 13406 3333
tri 13357 3308 13360 3311 ne
tri 7722 3277 7728 3283 ne
rect 7728 3277 13330 3283
rect 7619 3266 7682 3277
tri 7619 3263 7622 3266 ne
rect 7622 3263 7682 3266
tri 7682 3263 7696 3277 sw
tri 7728 3263 7742 3277 ne
rect 7742 3263 13330 3277
rect 4568 3229 6743 3263
tri 6743 3229 6777 3263 sw
tri 7622 3260 7625 3263 ne
rect 7625 3260 7696 3263
rect 4568 3228 6777 3229
rect -190 3210 6777 3228
tri 6777 3210 6796 3229 sw
rect -209 3164 6796 3210
rect 6852 3208 6858 3260
rect 6910 3208 6924 3260
rect 6976 3229 7539 3260
tri 7539 3229 7570 3260 sw
tri 7625 3229 7656 3260 ne
rect 7656 3249 7696 3260
tri 7696 3249 7710 3263 sw
tri 7742 3249 7756 3263 ne
rect 7756 3249 13330 3263
rect 7656 3229 7710 3249
tri 7710 3229 7730 3249 sw
tri 7756 3231 7774 3249 ne
rect 7774 3231 13330 3249
tri 13204 3229 13206 3231 ne
rect 13206 3229 13330 3231
rect 6976 3208 7570 3229
tri 7517 3191 7534 3208 ne
rect 7534 3197 7570 3208
tri 7570 3197 7602 3229 sw
tri 7656 3203 7682 3229 ne
rect 7682 3203 7730 3229
tri 7730 3203 7756 3229 sw
tri 13206 3206 13229 3229 ne
tri 7682 3197 7688 3203 ne
rect 7688 3197 13186 3203
rect 7534 3191 7602 3197
tri 7602 3191 7608 3197 sw
tri 7688 3191 7694 3197 ne
rect 7694 3191 13186 3197
tri 7534 3186 7539 3191 ne
rect 7539 3186 7608 3191
tri 7539 3164 7561 3186 ne
rect 7561 3164 7608 3186
tri 7561 3157 7568 3164 ne
rect 7568 3157 7608 3164
tri 7608 3157 7642 3191 sw
tri 7694 3157 7728 3191 ne
rect 7728 3157 12780 3191
rect 12814 3157 12852 3191
rect 12886 3157 12924 3191
rect 12958 3157 12996 3191
rect 13030 3157 13068 3191
rect 13102 3157 13140 3191
rect 13174 3157 13186 3191
tri 7568 3123 7602 3157 ne
rect 7602 3123 7642 3157
tri 7642 3123 7676 3157 sw
tri 7728 3151 7734 3157 ne
rect 7734 3151 13186 3157
tri 13216 3123 13229 3136 se
rect 13229 3123 13330 3229
tri 7602 3119 7606 3123 ne
rect 7606 3119 7676 3123
tri 7676 3119 7680 3123 sw
tri 7606 3117 7608 3119 ne
rect 7608 3117 7680 3119
tri 7680 3117 7682 3119 sw
rect 8017 3117 12736 3123
tri 13212 3119 13216 3123 se
rect 13216 3119 13330 3123
tri 7608 3083 7642 3117 ne
rect 7642 3083 7682 3117
tri 7682 3083 7716 3117 sw
rect 8017 3083 8029 3117
rect 8063 3083 8101 3117
rect 8135 3083 8173 3117
rect 8207 3083 8467 3117
rect 8501 3083 8542 3117
rect 8576 3083 8617 3117
rect 8651 3083 8692 3117
rect 8726 3083 8767 3117
rect 8801 3083 8841 3117
rect 8875 3083 8915 3117
rect 8949 3083 8989 3117
rect 9023 3083 9063 3117
rect 9097 3083 9137 3117
rect 9171 3083 9211 3117
rect 9245 3083 9285 3117
rect 9319 3083 9359 3117
rect 9393 3111 12736 3117
tri 13204 3111 13212 3119 se
rect 13212 3111 13330 3119
rect 13360 3263 13406 3311
rect 13360 3229 13366 3263
rect 13400 3229 13406 3263
rect 13360 3191 13406 3229
rect 13360 3157 13366 3191
rect 13400 3157 13406 3191
rect 13360 3119 13406 3157
rect 9393 3083 12624 3111
tri 7642 3077 7648 3083 ne
rect 7648 3077 7716 3083
tri 7716 3077 7722 3083 sw
rect 8017 3077 12624 3083
rect 12658 3077 12696 3111
rect 12730 3077 12736 3111
tri 7648 3049 7676 3077 ne
rect 7676 3049 7722 3077
tri 7722 3049 7750 3077 sw
tri 12606 3065 12618 3077 ne
rect 12618 3065 12736 3077
rect 13360 3085 13366 3119
rect 13400 3085 13406 3119
tri 7676 3047 7678 3049 ne
rect 7678 3047 9319 3049
tri 9319 3047 9321 3049 sw
tri 7678 3043 7682 3047 ne
rect 7682 3043 9321 3047
tri 7682 3009 7716 3043 ne
rect 7716 3009 8197 3043
rect 8231 3009 8269 3043
rect 8303 3013 9321 3043
tri 9321 3013 9355 3047 sw
rect 8303 3009 9355 3013
tri 9355 3009 9359 3013 sw
tri 7716 2975 7750 3009 ne
rect 7750 2975 9359 3009
tri 9359 2975 9393 3009 sw
rect 9412 2997 9418 3049
rect 9470 2997 9482 3049
rect 9534 2997 10330 3049
rect 10382 2997 10394 3049
rect 10446 2997 11616 3049
rect 11668 2997 11680 3049
rect 11732 2997 11738 3049
rect 13360 3047 13406 3085
tri 13335 3015 13360 3040 se
rect 13360 3015 13366 3047
tri 12538 3013 12540 3015 se
rect 12540 3013 13366 3015
rect 13400 3013 13406 3047
tri 12534 3009 12538 3013 se
rect 12538 3009 13406 3013
tri 12522 2997 12534 3009 se
rect 12534 2997 12552 3009
tri 12500 2975 12522 2997 se
rect 12522 2975 12552 2997
rect 12586 2975 12630 3009
rect 12664 2975 12707 3009
rect 12741 2975 12784 3009
rect 12818 2975 12861 3009
rect 12895 2975 12938 3009
rect 12972 2975 13015 3009
rect 13049 2975 13092 3009
rect 13126 2975 13169 3009
rect 13203 2975 13246 3009
rect 13280 2975 13406 3009
tri 7750 2945 7780 2975 ne
rect 7780 2969 9393 2975
tri 9393 2969 9399 2975 sw
tri 12494 2969 12500 2975 se
rect 12500 2973 13406 2975
tri 13406 2973 13431 2998 sw
rect 12500 2969 13619 2973
rect 7780 2945 13619 2969
tri 9275 2917 9303 2945 ne
rect 9303 2921 13619 2945
rect 13671 2921 13685 2973
rect 13737 2921 13751 2973
rect 13803 2921 13817 2973
rect 13869 2921 13883 2973
rect 13935 2921 13949 2973
rect 14001 2921 14015 2973
rect 14067 2921 14073 2973
rect 9303 2917 14073 2921
rect 8060 2911 8587 2917
rect 7907 2871 7953 2883
rect 8060 2877 8072 2911
rect 8106 2877 8148 2911
rect 8182 2877 8224 2911
rect 8258 2877 8300 2911
rect 8334 2877 8376 2911
rect 8410 2877 8452 2911
rect 8486 2877 8528 2911
rect 8562 2877 8587 2911
rect 8060 2871 8587 2877
rect 7907 2837 7913 2871
rect 7947 2837 7953 2871
tri 8575 2865 8581 2871 ne
rect 8581 2865 8587 2871
rect 8639 2865 8653 2917
rect 8705 2911 9261 2917
rect 8714 2877 8756 2911
rect 8790 2877 8832 2911
rect 8866 2877 8908 2911
rect 8942 2877 8984 2911
rect 9018 2877 9061 2911
rect 9095 2877 9138 2911
rect 9172 2877 9215 2911
rect 9249 2877 9261 2911
rect 8705 2871 9261 2877
tri 9303 2871 9349 2917 ne
rect 9349 2909 14073 2917
rect 9349 2871 13619 2909
rect 8705 2865 8711 2871
tri 8711 2865 8717 2871 nw
tri 9349 2865 9355 2871 ne
rect 9355 2865 13619 2871
tri 9355 2857 9363 2865 ne
rect 9363 2857 13619 2865
rect 13671 2857 13685 2909
rect 13737 2857 13751 2909
rect 13803 2857 13817 2909
rect 13869 2857 13883 2909
rect 13935 2857 13949 2909
rect 14001 2857 14015 2909
rect 14067 2857 14073 2909
tri 7904 2831 7907 2834 se
rect 7907 2831 7953 2837
tri 7953 2831 7956 2834 sw
rect 7904 2825 7956 2831
rect 7904 2764 7913 2773
rect 7947 2764 7956 2773
rect 7904 2760 7956 2764
rect 7904 2695 7913 2708
rect 7947 2695 7956 2708
rect 7904 2630 7913 2643
rect 7947 2630 7956 2643
rect 7904 2565 7913 2578
rect 7947 2565 7956 2578
rect 7904 2506 7956 2513
rect 7904 2500 7913 2506
rect 7947 2500 7956 2506
rect 7904 2435 7956 2448
rect 7904 2370 7956 2383
rect 7904 2305 7956 2318
rect 7904 2240 7956 2253
rect 7904 2180 7913 2188
rect 7947 2180 7956 2188
rect 7904 2175 7956 2180
rect 7904 2110 7913 2123
rect 7947 2110 7956 2123
rect 7904 2045 7913 2058
rect 7947 2045 7956 2058
rect 7904 1980 7913 1993
rect 7947 1980 7956 1993
rect 7904 1922 7956 1928
rect 7904 1915 7913 1922
rect 7947 1915 7956 1922
rect 7904 1850 7956 1863
rect 7904 1785 7956 1798
rect 7904 1720 7956 1733
rect 7904 1655 7956 1668
rect 7904 1596 7913 1603
rect 7947 1596 7956 1603
rect 7904 1590 7956 1596
rect 7904 1525 7913 1538
rect 7947 1525 7956 1538
rect 7904 1460 7913 1473
rect 7947 1460 7956 1473
rect 7904 1395 7913 1408
rect 7947 1395 7956 1408
rect 7904 1338 7956 1343
rect 7904 1330 7913 1338
rect 7947 1330 7956 1338
rect 7904 1265 7956 1278
rect 7904 1200 7956 1213
rect 7904 1135 7956 1148
rect 7904 1070 7956 1083
rect 7904 1012 7913 1018
rect 7947 1012 7956 1018
rect 7904 1005 7956 1012
rect 7904 941 7913 953
rect 7947 941 7956 953
rect 7904 877 7913 889
rect 7947 877 7956 889
rect 8047 2823 10829 2829
rect 8047 2817 8225 2823
rect 8047 2783 8053 2817
rect 8087 2783 8225 2817
rect 8047 2771 8225 2783
rect 8277 2771 8289 2823
rect 8341 2771 8353 2823
rect 8405 2817 10829 2823
rect 8405 2783 8965 2817
rect 8999 2783 9877 2817
rect 9911 2783 10789 2817
rect 10823 2783 10829 2817
rect 8405 2771 10829 2783
rect 8047 2757 10829 2771
rect 8047 2745 8225 2757
rect 8047 2711 8053 2745
rect 8087 2711 8225 2745
rect 8047 2705 8225 2711
rect 8277 2705 8289 2757
rect 8341 2705 8353 2757
rect 8405 2745 10829 2757
rect 8405 2711 8965 2745
rect 8999 2711 9877 2745
rect 9911 2711 10789 2745
rect 10823 2711 10829 2745
rect 8405 2705 10829 2711
rect 8047 2699 10829 2705
rect 8047 2680 8099 2699
tri 8099 2680 8118 2699 nw
tri 8934 2680 8953 2699 ne
rect 8953 2680 9011 2699
tri 9011 2680 9030 2699 nw
tri 9846 2680 9865 2699 ne
rect 9865 2680 9923 2699
tri 9923 2680 9942 2699 nw
tri 10758 2680 10777 2699 ne
rect 10777 2680 10829 2699
rect 8047 2673 8093 2680
tri 8093 2674 8099 2680 nw
tri 8953 2674 8959 2680 ne
rect 8047 2639 8053 2673
rect 8087 2639 8093 2673
rect 8959 2673 9005 2680
tri 9005 2674 9011 2680 nw
tri 9865 2674 9871 2680 ne
rect 8047 2601 8093 2639
rect 8047 2567 8053 2601
rect 8087 2567 8093 2601
rect 8047 2529 8093 2567
rect 8047 2495 8053 2529
rect 8087 2495 8093 2529
rect 8047 2457 8093 2495
rect 8047 2423 8053 2457
rect 8087 2423 8093 2457
rect 8047 2385 8093 2423
rect 8047 2351 8053 2385
rect 8087 2351 8093 2385
rect 8047 2313 8093 2351
rect 8047 2279 8053 2313
rect 8087 2279 8093 2313
rect 8047 2241 8093 2279
rect 8047 2207 8053 2241
rect 8087 2207 8093 2241
rect 8047 2169 8093 2207
rect 8047 2135 8053 2169
rect 8087 2135 8093 2169
rect 8503 2659 8549 2671
rect 8503 2625 8509 2659
rect 8543 2625 8549 2659
rect 8503 2585 8549 2625
rect 8503 2551 8509 2585
rect 8543 2551 8549 2585
rect 8503 2511 8549 2551
rect 8503 2477 8509 2511
rect 8543 2477 8549 2511
rect 8503 2437 8549 2477
rect 8503 2403 8509 2437
rect 8543 2403 8549 2437
rect 8503 2363 8549 2403
rect 8503 2329 8509 2363
rect 8543 2329 8549 2363
rect 8503 2289 8549 2329
rect 8503 2255 8509 2289
rect 8543 2255 8549 2289
rect 8503 2215 8549 2255
rect 8503 2181 8509 2215
rect 8543 2181 8549 2215
tri 8501 2157 8503 2159 ne
rect 8047 2097 8093 2135
rect 8047 2063 8053 2097
rect 8087 2063 8093 2097
rect 8047 2025 8093 2063
rect 8047 1991 8053 2025
rect 8087 1991 8093 2025
rect 8047 1953 8093 1991
rect 8047 1919 8053 1953
rect 8087 1919 8093 1953
rect 8047 1881 8093 1919
rect 8047 1847 8053 1881
rect 8087 1847 8093 1881
rect 8047 1809 8093 1847
rect 8047 1775 8053 1809
rect 8087 1775 8093 1809
rect 8047 1737 8093 1775
rect 8047 1703 8053 1737
rect 8087 1703 8093 1737
rect 8047 1665 8093 1703
rect 8047 1631 8053 1665
rect 8087 1631 8093 1665
rect 8047 1593 8093 1631
rect 8047 1559 8053 1593
rect 8087 1559 8093 1593
rect 8047 1521 8093 1559
rect 8047 1487 8053 1521
rect 8087 1487 8093 1521
rect 8047 1449 8093 1487
rect 8047 1415 8053 1449
rect 8087 1415 8093 1449
rect 8047 1377 8093 1415
rect 8047 1343 8053 1377
rect 8087 1343 8093 1377
rect 8047 1305 8093 1343
rect 8047 1271 8053 1305
rect 8087 1271 8093 1305
rect 8047 1233 8093 1271
rect 8047 1199 8053 1233
rect 8087 1199 8093 1233
rect 8047 1161 8093 1199
rect 8047 1127 8053 1161
rect 8087 1127 8093 1161
rect 8047 1089 8093 1127
rect 8047 1055 8053 1089
rect 8087 1055 8093 1089
rect 8047 1017 8093 1055
rect 8047 983 8053 1017
rect 8087 983 8093 1017
rect 8047 944 8093 983
rect 8047 910 8053 944
rect 8087 910 8093 944
rect 8047 871 8093 910
rect 8047 837 8053 871
rect 8087 837 8093 871
rect 8047 825 8093 837
rect 8503 2141 8549 2181
rect 8959 2639 8965 2673
rect 8999 2639 9005 2673
rect 9871 2673 9917 2680
tri 9917 2674 9923 2680 nw
tri 10777 2674 10783 2680 ne
rect 8959 2601 9005 2639
rect 8959 2567 8965 2601
rect 8999 2567 9005 2601
rect 8959 2529 9005 2567
rect 8959 2495 8965 2529
rect 8999 2495 9005 2529
rect 8959 2457 9005 2495
rect 8959 2423 8965 2457
rect 8999 2423 9005 2457
rect 8959 2385 9005 2423
rect 8959 2351 8965 2385
rect 8999 2351 9005 2385
rect 8959 2313 9005 2351
rect 8959 2279 8965 2313
rect 8999 2279 9005 2313
rect 8959 2241 9005 2279
rect 8959 2207 8965 2241
rect 8999 2207 9005 2241
rect 8959 2169 9005 2207
tri 8549 2155 8553 2159 nw
rect 8503 2107 8509 2141
rect 8543 2107 8549 2141
rect 8503 2067 8549 2107
rect 8503 2033 8509 2067
rect 8543 2033 8549 2067
rect 8503 1993 8549 2033
rect 8503 1959 8509 1993
rect 8543 1959 8549 1993
rect 8503 1919 8549 1959
rect 8503 1885 8509 1919
rect 8543 1885 8549 1919
rect 8503 1845 8549 1885
rect 8503 1811 8509 1845
rect 8543 1811 8549 1845
rect 8503 1771 8549 1811
rect 8503 1737 8509 1771
rect 8543 1737 8549 1771
rect 8503 1696 8549 1737
rect 8503 1662 8509 1696
rect 8543 1662 8549 1696
rect 8503 1621 8549 1662
rect 8503 1587 8509 1621
rect 8543 1587 8549 1621
rect 8503 1546 8549 1587
rect 8503 1512 8509 1546
rect 8543 1512 8549 1546
rect 8503 1471 8549 1512
rect 8503 1437 8509 1471
rect 8543 1437 8549 1471
rect 8503 1396 8549 1437
rect 8503 1362 8509 1396
rect 8543 1362 8549 1396
rect 8503 1321 8549 1362
rect 8503 1287 8509 1321
rect 8543 1287 8549 1321
rect 8503 1246 8549 1287
rect 8503 1212 8509 1246
rect 8543 1212 8549 1246
rect 8503 1171 8549 1212
rect 8503 1137 8509 1171
rect 8543 1137 8549 1171
rect 8503 1096 8549 1137
rect 8503 1062 8509 1096
rect 8543 1062 8549 1096
rect 8503 1021 8549 1062
rect 8503 987 8509 1021
rect 8543 987 8549 1021
rect 8503 946 8549 987
rect 8503 912 8509 946
rect 8543 912 8549 946
rect 8503 871 8549 912
rect 8503 837 8509 871
rect 8543 837 8549 871
rect 8503 825 8549 837
rect 8959 2135 8965 2169
rect 8999 2135 9005 2169
rect 9415 2659 9461 2671
rect 9415 2625 9421 2659
rect 9455 2625 9461 2659
rect 9415 2585 9461 2625
rect 9415 2551 9421 2585
rect 9455 2551 9461 2585
rect 9415 2511 9461 2551
rect 9415 2477 9421 2511
rect 9455 2477 9461 2511
rect 9415 2437 9461 2477
rect 9415 2403 9421 2437
rect 9455 2403 9461 2437
rect 9415 2363 9461 2403
rect 9415 2329 9421 2363
rect 9455 2329 9461 2363
rect 9415 2289 9461 2329
rect 9415 2255 9421 2289
rect 9455 2255 9461 2289
rect 9415 2215 9461 2255
rect 9415 2181 9421 2215
rect 9455 2181 9461 2215
tri 9412 2156 9415 2159 ne
rect 8959 2097 9005 2135
rect 8959 2063 8965 2097
rect 8999 2063 9005 2097
rect 8959 2025 9005 2063
rect 8959 1991 8965 2025
rect 8999 1991 9005 2025
rect 8959 1953 9005 1991
rect 8959 1919 8965 1953
rect 8999 1919 9005 1953
rect 8959 1881 9005 1919
rect 8959 1847 8965 1881
rect 8999 1847 9005 1881
rect 8959 1809 9005 1847
rect 8959 1775 8965 1809
rect 8999 1775 9005 1809
rect 8959 1737 9005 1775
rect 8959 1703 8965 1737
rect 8999 1703 9005 1737
rect 8959 1665 9005 1703
rect 8959 1631 8965 1665
rect 8999 1631 9005 1665
rect 8959 1593 9005 1631
rect 8959 1559 8965 1593
rect 8999 1559 9005 1593
rect 8959 1521 9005 1559
rect 8959 1487 8965 1521
rect 8999 1487 9005 1521
rect 8959 1449 9005 1487
rect 8959 1415 8965 1449
rect 8999 1415 9005 1449
rect 8959 1377 9005 1415
rect 8959 1343 8965 1377
rect 8999 1343 9005 1377
rect 8959 1305 9005 1343
rect 8959 1271 8965 1305
rect 8999 1271 9005 1305
rect 8959 1233 9005 1271
rect 8959 1199 8965 1233
rect 8999 1199 9005 1233
rect 8959 1161 9005 1199
rect 8959 1127 8965 1161
rect 8999 1127 9005 1161
rect 8959 1089 9005 1127
rect 8959 1055 8965 1089
rect 8999 1055 9005 1089
rect 8959 1017 9005 1055
rect 8959 983 8965 1017
rect 8999 983 9005 1017
rect 8959 944 9005 983
rect 8959 910 8965 944
rect 8999 910 9005 944
rect 8959 871 9005 910
rect 8959 837 8965 871
rect 8999 837 9005 871
rect 8959 825 9005 837
rect 9415 2141 9461 2181
rect 9871 2639 9877 2673
rect 9911 2639 9917 2673
rect 10783 2673 10829 2680
rect 9871 2601 9917 2639
rect 9871 2567 9877 2601
rect 9911 2567 9917 2601
rect 9871 2529 9917 2567
rect 9871 2495 9877 2529
rect 9911 2495 9917 2529
rect 9871 2457 9917 2495
rect 9871 2423 9877 2457
rect 9911 2423 9917 2457
rect 9871 2385 9917 2423
rect 9871 2351 9877 2385
rect 9911 2351 9917 2385
rect 9871 2313 9917 2351
rect 9871 2279 9877 2313
rect 9911 2279 9917 2313
rect 9871 2241 9917 2279
rect 9871 2207 9877 2241
rect 9911 2207 9917 2241
rect 9871 2169 9917 2207
tri 9461 2156 9464 2159 nw
rect 9415 2107 9421 2141
rect 9455 2107 9461 2141
rect 9415 2067 9461 2107
rect 9415 2033 9421 2067
rect 9455 2033 9461 2067
rect 9415 1993 9461 2033
rect 9415 1959 9421 1993
rect 9455 1959 9461 1993
rect 9415 1919 9461 1959
rect 9415 1885 9421 1919
rect 9455 1885 9461 1919
rect 9415 1845 9461 1885
rect 9415 1811 9421 1845
rect 9455 1811 9461 1845
rect 9415 1771 9461 1811
rect 9415 1737 9421 1771
rect 9455 1737 9461 1771
rect 9415 1696 9461 1737
rect 9415 1662 9421 1696
rect 9455 1662 9461 1696
rect 9415 1621 9461 1662
rect 9415 1587 9421 1621
rect 9455 1587 9461 1621
rect 9415 1546 9461 1587
rect 9415 1512 9421 1546
rect 9455 1512 9461 1546
rect 9415 1471 9461 1512
rect 9415 1437 9421 1471
rect 9455 1437 9461 1471
rect 9415 1396 9461 1437
rect 9415 1362 9421 1396
rect 9455 1362 9461 1396
rect 9415 1321 9461 1362
rect 9415 1287 9421 1321
rect 9455 1287 9461 1321
rect 9415 1246 9461 1287
rect 9415 1212 9421 1246
rect 9455 1212 9461 1246
rect 9415 1171 9461 1212
rect 9415 1137 9421 1171
rect 9455 1137 9461 1171
rect 9415 1096 9461 1137
rect 9415 1062 9421 1096
rect 9455 1062 9461 1096
rect 9415 1021 9461 1062
rect 9415 987 9421 1021
rect 9455 987 9461 1021
rect 9415 946 9461 987
rect 9415 912 9421 946
rect 9455 912 9461 946
rect 9415 871 9461 912
rect 9415 837 9421 871
rect 9455 837 9461 871
rect 9415 825 9461 837
rect 9871 2135 9877 2169
rect 9911 2135 9917 2169
rect 10327 2659 10373 2671
rect 10327 2625 10333 2659
rect 10367 2625 10373 2659
rect 10327 2585 10373 2625
rect 10327 2551 10333 2585
rect 10367 2551 10373 2585
rect 10327 2511 10373 2551
rect 10327 2477 10333 2511
rect 10367 2477 10373 2511
rect 10327 2437 10373 2477
rect 10327 2403 10333 2437
rect 10367 2403 10373 2437
rect 10327 2363 10373 2403
rect 10327 2329 10333 2363
rect 10367 2329 10373 2363
rect 10327 2289 10373 2329
rect 10327 2255 10333 2289
rect 10367 2255 10373 2289
rect 10327 2215 10373 2255
rect 10327 2181 10333 2215
rect 10367 2181 10373 2215
tri 10324 2156 10327 2159 ne
rect 9871 2097 9917 2135
rect 9871 2063 9877 2097
rect 9911 2063 9917 2097
rect 9871 2025 9917 2063
rect 9871 1991 9877 2025
rect 9911 1991 9917 2025
rect 9871 1953 9917 1991
rect 9871 1919 9877 1953
rect 9911 1919 9917 1953
rect 9871 1881 9917 1919
rect 9871 1847 9877 1881
rect 9911 1847 9917 1881
rect 9871 1809 9917 1847
rect 9871 1775 9877 1809
rect 9911 1775 9917 1809
rect 9871 1737 9917 1775
rect 9871 1703 9877 1737
rect 9911 1703 9917 1737
rect 9871 1665 9917 1703
rect 9871 1631 9877 1665
rect 9911 1631 9917 1665
rect 9871 1593 9917 1631
rect 9871 1559 9877 1593
rect 9911 1559 9917 1593
rect 9871 1521 9917 1559
rect 9871 1487 9877 1521
rect 9911 1487 9917 1521
rect 9871 1449 9917 1487
rect 9871 1415 9877 1449
rect 9911 1415 9917 1449
rect 9871 1377 9917 1415
rect 9871 1343 9877 1377
rect 9911 1343 9917 1377
rect 9871 1305 9917 1343
rect 9871 1271 9877 1305
rect 9911 1271 9917 1305
rect 9871 1233 9917 1271
rect 9871 1199 9877 1233
rect 9911 1199 9917 1233
rect 9871 1161 9917 1199
rect 9871 1127 9877 1161
rect 9911 1127 9917 1161
rect 9871 1089 9917 1127
rect 9871 1055 9877 1089
rect 9911 1055 9917 1089
rect 9871 1017 9917 1055
rect 9871 983 9877 1017
rect 9911 983 9917 1017
rect 9871 944 9917 983
rect 9871 910 9877 944
rect 9911 910 9917 944
rect 9871 871 9917 910
rect 9871 837 9877 871
rect 9911 837 9917 871
rect 9871 825 9917 837
rect 10327 2141 10373 2181
rect 10783 2639 10789 2673
rect 10823 2639 10829 2673
rect 10783 2601 10829 2639
rect 10783 2567 10789 2601
rect 10823 2567 10829 2601
rect 10783 2529 10829 2567
rect 10783 2495 10789 2529
rect 10823 2495 10829 2529
rect 10783 2457 10829 2495
rect 10783 2423 10789 2457
rect 10823 2423 10829 2457
rect 10783 2385 10829 2423
rect 10783 2351 10789 2385
rect 10823 2351 10829 2385
rect 10783 2313 10829 2351
rect 10783 2279 10789 2313
rect 10823 2279 10829 2313
rect 10783 2241 10829 2279
rect 10783 2207 10789 2241
rect 10823 2207 10829 2241
rect 10783 2169 10829 2207
tri 10373 2156 10376 2159 nw
rect 10327 2107 10333 2141
rect 10367 2107 10373 2141
rect 10327 2067 10373 2107
rect 10327 2033 10333 2067
rect 10367 2033 10373 2067
rect 10327 1993 10373 2033
rect 10327 1959 10333 1993
rect 10367 1959 10373 1993
rect 10327 1919 10373 1959
rect 10327 1885 10333 1919
rect 10367 1885 10373 1919
rect 10327 1845 10373 1885
rect 10327 1811 10333 1845
rect 10367 1811 10373 1845
rect 10327 1771 10373 1811
rect 10327 1737 10333 1771
rect 10367 1737 10373 1771
rect 10327 1696 10373 1737
rect 10327 1662 10333 1696
rect 10367 1662 10373 1696
rect 10327 1621 10373 1662
rect 10327 1587 10333 1621
rect 10367 1587 10373 1621
rect 10327 1546 10373 1587
rect 10327 1512 10333 1546
rect 10367 1512 10373 1546
rect 10327 1471 10373 1512
rect 10327 1437 10333 1471
rect 10367 1437 10373 1471
rect 10327 1396 10373 1437
rect 10327 1362 10333 1396
rect 10367 1362 10373 1396
rect 10327 1321 10373 1362
rect 10327 1287 10333 1321
rect 10367 1287 10373 1321
rect 10327 1246 10373 1287
rect 10327 1212 10333 1246
rect 10367 1212 10373 1246
rect 10327 1171 10373 1212
rect 10327 1137 10333 1171
rect 10367 1137 10373 1171
rect 10327 1096 10373 1137
rect 10327 1062 10333 1096
rect 10367 1062 10373 1096
rect 10327 1021 10373 1062
rect 10327 987 10333 1021
rect 10367 987 10373 1021
rect 10327 946 10373 987
rect 10327 912 10333 946
rect 10367 912 10373 946
rect 10327 871 10373 912
rect 10327 837 10333 871
rect 10367 837 10373 871
rect 10327 825 10373 837
rect 10783 2135 10789 2169
rect 10823 2135 10829 2169
rect 10783 2097 10829 2135
rect 10783 2063 10789 2097
rect 10823 2063 10829 2097
rect 10783 2025 10829 2063
rect 10783 1991 10789 2025
rect 10823 1991 10829 2025
rect 10783 1953 10829 1991
rect 10783 1919 10789 1953
rect 10823 1919 10829 1953
rect 10783 1881 10829 1919
rect 10783 1847 10789 1881
rect 10823 1847 10829 1881
rect 10783 1809 10829 1847
rect 10783 1775 10789 1809
rect 10823 1775 10829 1809
rect 10783 1737 10829 1775
rect 10783 1703 10789 1737
rect 10823 1703 10829 1737
rect 10783 1665 10829 1703
rect 10783 1631 10789 1665
rect 10823 1631 10829 1665
rect 10783 1593 10829 1631
rect 10783 1559 10789 1593
rect 10823 1559 10829 1593
rect 10783 1521 10829 1559
rect 10783 1487 10789 1521
rect 10823 1487 10829 1521
rect 10783 1449 10829 1487
rect 10783 1415 10789 1449
rect 10823 1415 10829 1449
rect 10783 1377 10829 1415
rect 10783 1343 10789 1377
rect 10823 1343 10829 1377
rect 10783 1305 10829 1343
rect 10783 1271 10789 1305
rect 10823 1271 10829 1305
rect 10783 1233 10829 1271
rect 10783 1199 10789 1233
rect 10823 1199 10829 1233
rect 10783 1161 10829 1199
rect 10783 1127 10789 1161
rect 10823 1127 10829 1161
rect 10783 1089 10829 1127
rect 10783 1055 10789 1089
rect 10823 1055 10829 1089
rect 10783 1017 10829 1055
rect 10783 983 10789 1017
rect 10823 983 10829 1017
rect 10783 944 10829 983
rect 10783 910 10789 944
rect 10823 910 10829 944
rect 10783 871 10829 910
rect 10783 837 10789 871
rect 10823 837 10829 871
rect 10783 825 10829 837
rect 10923 2817 10969 2829
rect 10923 2783 10929 2817
rect 10963 2783 10969 2817
rect 10923 2744 10969 2783
rect 10923 2710 10929 2744
rect 10963 2710 10969 2744
rect 10923 2671 10969 2710
rect 10923 2637 10929 2671
rect 10963 2637 10969 2671
rect 10923 2598 10969 2637
rect 10923 2564 10929 2598
rect 10963 2564 10969 2598
rect 10923 2525 10969 2564
rect 10923 2491 10929 2525
rect 10963 2491 10969 2525
rect 10923 2452 10969 2491
rect 10923 2418 10929 2452
rect 10963 2418 10969 2452
rect 10923 2379 10969 2418
rect 10923 2345 10929 2379
rect 10963 2345 10969 2379
rect 10923 2306 10969 2345
rect 10923 2272 10929 2306
rect 10963 2272 10969 2306
rect 10923 2233 10969 2272
rect 10923 2199 10929 2233
rect 10963 2199 10969 2233
rect 10923 2159 10969 2199
rect 10923 2125 10929 2159
rect 10963 2125 10969 2159
rect 10923 2085 10969 2125
rect 10923 2051 10929 2085
rect 10963 2051 10969 2085
rect 10923 2011 10969 2051
rect 10923 1977 10929 2011
rect 10963 1977 10969 2011
rect 10923 1937 10969 1977
rect 10923 1903 10929 1937
rect 10963 1903 10969 1937
rect 10923 1863 10969 1903
rect 10923 1829 10929 1863
rect 10963 1829 10969 1863
rect 10923 1789 10969 1829
rect 10923 1755 10929 1789
rect 10963 1755 10969 1789
rect 10923 1715 10969 1755
rect 11436 2714 14079 2729
rect 11436 2680 11448 2714
rect 11482 2680 11522 2714
rect 11556 2680 11596 2714
rect 11630 2680 11670 2714
rect 11704 2680 11744 2714
rect 11778 2680 11818 2714
rect 11852 2680 11892 2714
rect 11926 2680 11966 2714
rect 12000 2680 12040 2714
rect 12074 2680 12114 2714
rect 12148 2680 12188 2714
rect 12222 2680 12262 2714
rect 12296 2680 12336 2714
rect 12370 2680 12410 2714
rect 12444 2680 12484 2714
rect 12518 2680 12558 2714
rect 12592 2680 12632 2714
rect 12666 2680 12706 2714
rect 12740 2680 12780 2714
rect 12814 2680 12854 2714
rect 12888 2680 12928 2714
rect 12962 2680 13002 2714
rect 13036 2680 13076 2714
rect 13110 2680 13150 2714
rect 13184 2680 13224 2714
rect 13258 2680 13298 2714
rect 13332 2680 13372 2714
rect 13406 2680 13446 2714
rect 13480 2680 13520 2714
rect 13554 2680 13594 2714
rect 13628 2680 13668 2714
rect 13702 2680 13741 2714
rect 13775 2680 13814 2714
rect 13848 2680 13887 2714
rect 13921 2680 13960 2714
rect 13994 2680 14033 2714
rect 14067 2680 14079 2714
rect 11436 2642 14079 2680
rect 11436 2608 11448 2642
rect 11482 2608 11522 2642
rect 11556 2608 11596 2642
rect 11630 2608 11670 2642
rect 11704 2608 11744 2642
rect 11778 2608 11818 2642
rect 11852 2608 11892 2642
rect 11926 2608 11966 2642
rect 12000 2608 12040 2642
rect 12074 2608 12114 2642
rect 12148 2608 12188 2642
rect 12222 2608 12262 2642
rect 12296 2608 12336 2642
rect 12370 2608 12410 2642
rect 12444 2608 12484 2642
rect 12518 2608 12558 2642
rect 12592 2608 12632 2642
rect 12666 2608 12706 2642
rect 12740 2608 12780 2642
rect 12814 2608 12854 2642
rect 12888 2608 12928 2642
rect 12962 2608 13002 2642
rect 13036 2608 13076 2642
rect 13110 2608 13150 2642
rect 13184 2608 13224 2642
rect 13258 2608 13298 2642
rect 13332 2608 13372 2642
rect 13406 2608 13446 2642
rect 13480 2608 13520 2642
rect 13554 2608 13594 2642
rect 13628 2608 13668 2642
rect 13702 2608 13741 2642
rect 13775 2608 13814 2642
rect 13848 2608 13887 2642
rect 13921 2608 13960 2642
rect 13994 2608 14033 2642
rect 14067 2608 14079 2642
rect 11436 2570 14079 2608
rect 11436 2536 11448 2570
rect 11482 2536 11522 2570
rect 11556 2536 11596 2570
rect 11630 2536 11670 2570
rect 11704 2536 11744 2570
rect 11778 2536 11818 2570
rect 11852 2536 11892 2570
rect 11926 2536 11966 2570
rect 12000 2536 12040 2570
rect 12074 2536 12114 2570
rect 12148 2536 12188 2570
rect 12222 2536 12262 2570
rect 12296 2536 12336 2570
rect 12370 2536 12410 2570
rect 12444 2536 12484 2570
rect 12518 2536 12558 2570
rect 12592 2536 12632 2570
rect 12666 2536 12706 2570
rect 12740 2536 12780 2570
rect 12814 2536 12854 2570
rect 12888 2536 12928 2570
rect 12962 2536 13002 2570
rect 13036 2536 13076 2570
rect 13110 2536 13150 2570
rect 13184 2536 13224 2570
rect 13258 2536 13298 2570
rect 13332 2536 13372 2570
rect 13406 2536 13446 2570
rect 13480 2536 13520 2570
rect 13554 2536 13594 2570
rect 13628 2536 13668 2570
rect 13702 2536 13741 2570
rect 13775 2536 13814 2570
rect 13848 2536 13887 2570
rect 13921 2536 13960 2570
rect 13994 2536 14033 2570
rect 14067 2536 14079 2570
rect 11436 2498 14079 2536
rect 11436 2464 11448 2498
rect 11482 2464 11522 2498
rect 11556 2464 11596 2498
rect 11630 2464 11670 2498
rect 11704 2464 11744 2498
rect 11778 2464 11818 2498
rect 11852 2464 11892 2498
rect 11926 2464 11966 2498
rect 12000 2464 12040 2498
rect 12074 2464 12114 2498
rect 12148 2464 12188 2498
rect 12222 2464 12262 2498
rect 12296 2464 12336 2498
rect 12370 2464 12410 2498
rect 12444 2464 12484 2498
rect 12518 2464 12558 2498
rect 12592 2464 12632 2498
rect 12666 2464 12706 2498
rect 12740 2464 12780 2498
rect 12814 2464 12854 2498
rect 12888 2464 12928 2498
rect 12962 2464 13002 2498
rect 13036 2464 13076 2498
rect 13110 2464 13150 2498
rect 13184 2464 13224 2498
rect 13258 2464 13298 2498
rect 13332 2464 13372 2498
rect 13406 2464 13446 2498
rect 13480 2464 13520 2498
rect 13554 2464 13594 2498
rect 13628 2464 13668 2498
rect 13702 2464 13741 2498
rect 13775 2464 13814 2498
rect 13848 2464 13887 2498
rect 13921 2464 13960 2498
rect 13994 2464 14033 2498
rect 14067 2464 14079 2498
rect 11436 2454 14079 2464
rect 11436 2426 12145 2454
rect 12197 2426 14079 2454
rect 11436 2392 11448 2426
rect 11482 2392 11522 2426
rect 11556 2392 11596 2426
rect 11630 2392 11670 2426
rect 11704 2392 11744 2426
rect 11778 2392 11818 2426
rect 11852 2392 11892 2426
rect 11926 2392 11966 2426
rect 12000 2392 12040 2426
rect 12074 2400 12114 2426
rect 12074 2392 12090 2400
rect 12148 2392 12188 2402
rect 12222 2392 12262 2426
rect 12296 2411 12336 2426
rect 12335 2392 12336 2411
rect 12370 2392 12410 2426
rect 12444 2392 12484 2426
rect 12518 2392 12558 2426
rect 12592 2392 12632 2426
rect 12666 2392 12706 2426
rect 12740 2392 12780 2426
rect 12814 2392 12854 2426
rect 12888 2392 12928 2426
rect 12962 2392 13002 2426
rect 13036 2392 13076 2426
rect 13110 2392 13150 2426
rect 13184 2392 13224 2426
rect 13258 2392 13298 2426
rect 13332 2392 13372 2426
rect 13406 2392 13446 2426
rect 13480 2392 13520 2426
rect 13554 2392 13594 2426
rect 13628 2392 13668 2426
rect 13702 2392 13741 2426
rect 13775 2392 13814 2426
rect 13848 2392 13887 2426
rect 13921 2392 13960 2426
rect 13994 2392 14033 2426
rect 14067 2392 14079 2426
rect 11436 2354 12090 2392
rect 12142 2359 12283 2392
rect 12335 2359 14079 2392
rect 12142 2357 14079 2359
rect 12142 2354 12228 2357
rect 12280 2354 14079 2357
rect 11436 2320 11448 2354
rect 11482 2320 11522 2354
rect 11556 2320 11596 2354
rect 11630 2320 11670 2354
rect 11704 2320 11744 2354
rect 11778 2320 11818 2354
rect 11852 2320 11892 2354
rect 11926 2320 11966 2354
rect 12000 2346 12040 2354
rect 12074 2348 12090 2354
rect 12074 2346 12114 2348
rect 12000 2320 12035 2346
rect 12087 2320 12114 2346
rect 12148 2320 12188 2354
rect 12222 2320 12228 2354
rect 12296 2320 12336 2354
rect 12370 2320 12410 2354
rect 12444 2320 12484 2354
rect 12518 2320 12558 2354
rect 12592 2320 12632 2354
rect 12666 2320 12706 2354
rect 12740 2320 12780 2354
rect 12814 2320 12854 2354
rect 12888 2320 12928 2354
rect 12962 2320 13002 2354
rect 13036 2320 13076 2354
rect 13110 2320 13150 2354
rect 13184 2320 13224 2354
rect 13258 2320 13298 2354
rect 13332 2320 13372 2354
rect 13406 2320 13446 2354
rect 13480 2320 13520 2354
rect 13554 2320 13594 2354
rect 13628 2320 13668 2354
rect 13702 2320 13741 2354
rect 13775 2320 13814 2354
rect 13848 2320 13887 2354
rect 13921 2320 13960 2354
rect 13994 2320 14033 2354
rect 14067 2320 14079 2354
rect 11436 2294 12035 2320
rect 12087 2305 12228 2320
rect 12280 2305 14079 2320
rect 12087 2303 14079 2305
rect 12087 2294 12173 2303
rect 11436 2292 12173 2294
rect 11436 2282 11980 2292
rect 12032 2282 12173 2292
rect 12225 2282 14079 2303
rect 11436 2248 11448 2282
rect 11482 2248 11522 2282
rect 11556 2248 11596 2282
rect 11630 2248 11670 2282
rect 11704 2248 11744 2282
rect 11778 2248 11818 2282
rect 11852 2248 11892 2282
rect 11926 2248 11966 2282
rect 12032 2248 12040 2282
rect 12074 2248 12114 2282
rect 12148 2251 12173 2282
rect 12225 2251 12262 2282
rect 12148 2249 12188 2251
rect 12170 2248 12188 2249
rect 12222 2248 12262 2251
rect 12296 2248 12336 2282
rect 12370 2248 12410 2282
rect 12444 2248 12484 2282
rect 12518 2248 12558 2282
rect 12592 2248 12632 2282
rect 12666 2248 12706 2282
rect 12740 2248 12780 2282
rect 12814 2248 12854 2282
rect 12888 2248 12928 2282
rect 12962 2248 13002 2282
rect 13036 2248 13076 2282
rect 13110 2248 13150 2282
rect 13184 2248 13224 2282
rect 13258 2248 13298 2282
rect 13332 2248 13372 2282
rect 13406 2248 13446 2282
rect 13480 2248 13520 2282
rect 13554 2248 13594 2282
rect 13628 2248 13668 2282
rect 13702 2248 13741 2282
rect 13775 2248 13814 2282
rect 13848 2248 13887 2282
rect 13921 2248 13960 2282
rect 13994 2248 14033 2282
rect 14067 2248 14079 2282
rect 11436 2240 11980 2248
rect 12032 2240 12118 2248
rect 11436 2238 12118 2240
rect 11436 2210 11925 2238
rect 11977 2210 12118 2238
rect 12170 2210 14079 2248
rect 11436 2176 11448 2210
rect 11482 2176 11522 2210
rect 11556 2176 11596 2210
rect 11630 2176 11670 2210
rect 11704 2176 11744 2210
rect 11778 2176 11818 2210
rect 11852 2184 11892 2210
rect 11852 2176 11870 2184
rect 11926 2176 11966 2186
rect 12000 2176 12040 2210
rect 12074 2195 12114 2210
rect 12170 2197 12188 2210
rect 12148 2176 12188 2197
rect 12222 2176 12262 2210
rect 12296 2176 12336 2210
rect 12370 2176 12410 2210
rect 12444 2176 12484 2210
rect 12518 2176 12558 2210
rect 12592 2176 12632 2210
rect 12666 2176 12706 2210
rect 12740 2176 12780 2210
rect 12814 2176 12854 2210
rect 12888 2176 12928 2210
rect 12962 2176 13002 2210
rect 13036 2176 13076 2210
rect 13110 2176 13150 2210
rect 13184 2176 13224 2210
rect 13258 2176 13298 2210
rect 13332 2176 13372 2210
rect 13406 2176 13446 2210
rect 13480 2176 13520 2210
rect 13554 2176 13594 2210
rect 13628 2176 13668 2210
rect 13702 2176 13741 2210
rect 13775 2176 13814 2210
rect 13848 2176 13887 2210
rect 13921 2176 13960 2210
rect 13994 2176 14033 2210
rect 14067 2176 14079 2210
rect 11436 2138 11870 2176
rect 11922 2143 12063 2176
rect 12115 2143 14079 2176
rect 11922 2141 14079 2143
rect 11922 2138 12008 2141
rect 12060 2138 14079 2141
rect 11436 2104 11448 2138
rect 11482 2104 11522 2138
rect 11556 2104 11596 2138
rect 11630 2104 11670 2138
rect 11704 2104 11744 2138
rect 11778 2130 11818 2138
rect 11852 2132 11870 2138
rect 11852 2130 11892 2132
rect 11778 2104 11815 2130
rect 11867 2104 11892 2130
rect 11926 2104 11966 2138
rect 12000 2104 12008 2138
rect 12074 2104 12114 2138
rect 12148 2104 12188 2138
rect 12222 2104 12262 2138
rect 12296 2104 12336 2138
rect 12370 2104 12410 2138
rect 12444 2104 12484 2138
rect 12518 2104 12558 2138
rect 12592 2104 12632 2138
rect 12666 2104 12706 2138
rect 12740 2104 12780 2138
rect 12814 2104 12854 2138
rect 12888 2104 12928 2138
rect 12962 2104 13002 2138
rect 13036 2104 13076 2138
rect 13110 2104 13150 2138
rect 13184 2104 13224 2138
rect 13258 2104 13298 2138
rect 13332 2104 13372 2138
rect 13406 2104 13446 2138
rect 13480 2104 13520 2138
rect 13554 2104 13594 2138
rect 13628 2104 13668 2138
rect 13702 2104 13741 2138
rect 13775 2104 13814 2138
rect 13848 2104 13887 2138
rect 13921 2104 13960 2138
rect 13994 2104 14033 2138
rect 14067 2104 14079 2138
rect 11436 2078 11815 2104
rect 11867 2089 12008 2104
rect 12060 2089 14079 2104
rect 11867 2087 14079 2089
rect 11867 2078 11953 2087
rect 11436 2076 11953 2078
rect 11436 2066 11760 2076
rect 11812 2066 11953 2076
rect 12005 2066 14079 2087
rect 11436 2032 11448 2066
rect 11482 2032 11522 2066
rect 11556 2032 11596 2066
rect 11630 2032 11670 2066
rect 11704 2032 11744 2066
rect 11812 2032 11818 2066
rect 11852 2032 11892 2066
rect 11926 2035 11953 2066
rect 12005 2035 12040 2066
rect 11926 2033 11966 2035
rect 11950 2032 11966 2033
rect 12000 2032 12040 2035
rect 12074 2032 12114 2066
rect 12148 2032 12188 2066
rect 12222 2032 12262 2066
rect 12296 2032 12336 2066
rect 12370 2032 12410 2066
rect 12444 2032 12484 2066
rect 12518 2032 12558 2066
rect 12592 2032 12632 2066
rect 12666 2032 12706 2066
rect 12740 2032 12780 2066
rect 12814 2032 12854 2066
rect 12888 2032 12928 2066
rect 12962 2032 13002 2066
rect 13036 2032 13076 2066
rect 13110 2032 13150 2066
rect 13184 2032 13224 2066
rect 13258 2032 13298 2066
rect 13332 2032 13372 2066
rect 13406 2032 13446 2066
rect 13480 2032 13520 2066
rect 13554 2032 13594 2066
rect 13628 2032 13668 2066
rect 13702 2032 13741 2066
rect 13775 2032 13814 2066
rect 13848 2032 13887 2066
rect 13921 2032 13960 2066
rect 13994 2032 14033 2066
rect 14067 2032 14079 2066
rect 11436 2024 11760 2032
rect 11812 2024 11898 2032
rect 11436 2022 11898 2024
rect 11436 1994 11705 2022
rect 11757 1994 11898 2022
rect 11950 1994 14079 2032
rect 11436 1960 11448 1994
rect 11482 1960 11522 1994
rect 11556 1960 11596 1994
rect 11630 1960 11670 1994
rect 11704 1970 11705 1994
rect 11704 1960 11744 1970
rect 11778 1960 11818 1994
rect 11852 1979 11892 1994
rect 11950 1981 11966 1994
rect 11926 1960 11966 1981
rect 12000 1960 12040 1994
rect 12074 1960 12114 1994
rect 12148 1960 12188 1994
rect 12222 1960 12262 1994
rect 12296 1960 12336 1994
rect 12370 1960 12410 1994
rect 12444 1960 12484 1994
rect 12518 1960 12558 1994
rect 12592 1960 12632 1994
rect 12666 1960 12706 1994
rect 12740 1960 12780 1994
rect 12814 1960 12854 1994
rect 12888 1960 12928 1994
rect 12962 1960 13002 1994
rect 13036 1960 13076 1994
rect 13110 1960 13150 1994
rect 13184 1960 13224 1994
rect 13258 1960 13298 1994
rect 13332 1960 13372 1994
rect 13406 1960 13446 1994
rect 13480 1960 13520 1994
rect 13554 1960 13594 1994
rect 13628 1960 13668 1994
rect 13702 1960 13741 1994
rect 13775 1960 13814 1994
rect 13848 1960 13887 1994
rect 13921 1960 13960 1994
rect 13994 1960 14033 1994
rect 14067 1960 14079 1994
rect 11436 1927 11843 1960
rect 11895 1927 14079 1960
rect 11436 1922 14079 1927
rect 11436 1888 11448 1922
rect 11482 1888 11522 1922
rect 11556 1888 11596 1922
rect 11630 1888 11670 1922
rect 11704 1888 11744 1922
rect 11778 1888 11818 1922
rect 11852 1888 11892 1922
rect 11926 1888 11966 1922
rect 12000 1888 12040 1922
rect 12074 1888 12114 1922
rect 12148 1888 12188 1922
rect 12222 1888 12262 1922
rect 12296 1888 12336 1922
rect 12370 1888 12410 1922
rect 12444 1888 12484 1922
rect 12518 1888 12558 1922
rect 12592 1888 12632 1922
rect 12666 1888 12706 1922
rect 12740 1888 12780 1922
rect 12814 1888 12854 1922
rect 12888 1888 12928 1922
rect 12962 1888 13002 1922
rect 13036 1888 13076 1922
rect 13110 1888 13150 1922
rect 13184 1888 13224 1922
rect 13258 1888 13298 1922
rect 13332 1888 13372 1922
rect 13406 1888 13446 1922
rect 13480 1888 13520 1922
rect 13554 1888 13594 1922
rect 13628 1888 13668 1922
rect 13702 1888 13741 1922
rect 13775 1888 13814 1922
rect 13848 1888 13887 1922
rect 13921 1888 13960 1922
rect 13994 1888 14033 1922
rect 14067 1888 14079 1922
rect 11436 1850 14079 1888
rect 11436 1816 11448 1850
rect 11482 1816 11522 1850
rect 11556 1816 11596 1850
rect 11630 1816 11670 1850
rect 11704 1816 11744 1850
rect 11778 1816 11818 1850
rect 11852 1816 11892 1850
rect 11926 1816 11966 1850
rect 12000 1816 12040 1850
rect 12074 1816 12114 1850
rect 12148 1816 12188 1850
rect 12222 1816 12262 1850
rect 12296 1816 12336 1850
rect 12370 1816 12410 1850
rect 12444 1816 12484 1850
rect 12518 1816 12558 1850
rect 12592 1816 12632 1850
rect 12666 1816 12706 1850
rect 12740 1816 12780 1850
rect 12814 1816 12854 1850
rect 12888 1816 12928 1850
rect 12962 1816 13002 1850
rect 13036 1816 13076 1850
rect 13110 1816 13150 1850
rect 13184 1816 13224 1850
rect 13258 1816 13298 1850
rect 13332 1816 13372 1850
rect 13406 1816 13446 1850
rect 13480 1816 13520 1850
rect 13554 1816 13594 1850
rect 13628 1816 13668 1850
rect 13702 1816 13741 1850
rect 13775 1816 13814 1850
rect 13848 1816 13887 1850
rect 13921 1816 13960 1850
rect 13994 1816 14033 1850
rect 14067 1816 14079 1850
rect 11436 1778 14079 1816
rect 11436 1744 11448 1778
rect 11482 1744 11522 1778
rect 11556 1744 11596 1778
rect 11630 1744 11670 1778
rect 11704 1744 11744 1778
rect 11778 1744 11818 1778
rect 11852 1744 11892 1778
rect 11926 1744 11966 1778
rect 12000 1744 12040 1778
rect 12074 1744 12114 1778
rect 12148 1744 12188 1778
rect 12222 1744 12262 1778
rect 12296 1744 12336 1778
rect 12370 1744 12410 1778
rect 12444 1744 12484 1778
rect 12518 1744 12558 1778
rect 12592 1744 12632 1778
rect 12666 1744 12706 1778
rect 12740 1744 12780 1778
rect 12814 1744 12854 1778
rect 12888 1744 12928 1778
rect 12962 1744 13002 1778
rect 13036 1744 13076 1778
rect 13110 1744 13150 1778
rect 13184 1744 13224 1778
rect 13258 1744 13298 1778
rect 13332 1744 13372 1778
rect 13406 1744 13446 1778
rect 13480 1744 13520 1778
rect 13554 1744 13594 1778
rect 13628 1744 13668 1778
rect 13702 1744 13741 1778
rect 13775 1744 13814 1778
rect 13848 1744 13887 1778
rect 13921 1744 13960 1778
rect 13994 1744 14033 1778
rect 14067 1744 14079 1778
rect 11436 1729 14079 1744
rect 10923 1681 10929 1715
rect 10963 1681 10969 1715
rect 10923 1641 10969 1681
rect 10923 1607 10929 1641
rect 10963 1607 10969 1641
rect 10923 1567 10969 1607
rect 10923 1533 10929 1567
rect 10963 1533 10969 1567
rect 10923 1493 10969 1533
rect 10923 1459 10929 1493
rect 10963 1459 10969 1493
rect 10923 1419 10969 1459
rect 10923 1385 10929 1419
rect 10963 1385 10969 1419
rect 10923 1345 10969 1385
rect 10923 1311 10929 1345
rect 10963 1311 10969 1345
rect 10923 1271 10969 1311
rect 10923 1237 10929 1271
rect 10963 1237 10969 1271
rect 10923 1197 10969 1237
rect 10923 1163 10929 1197
rect 10963 1163 10969 1197
rect 10923 1123 10969 1163
rect 10923 1089 10929 1123
rect 10963 1089 10969 1123
rect 10923 1049 10969 1089
rect 10923 1015 10929 1049
rect 10963 1015 10969 1049
rect 10923 975 10969 1015
rect 10923 941 10929 975
rect 10963 941 10969 975
rect 10923 901 10969 941
rect 10923 867 10929 901
rect 10963 867 10969 901
rect 10923 827 10969 867
rect 7904 813 7913 825
rect 7947 813 7956 825
rect 10923 793 10929 827
rect 10963 793 10969 827
tri 7956 761 7981 786 sw
tri 10898 761 10923 786 se
rect 10923 761 10969 793
rect 7904 755 8992 761
rect 9044 755 9056 761
rect 9108 755 9121 761
rect 9173 755 9186 761
rect 9238 755 10969 761
rect 7904 749 7919 755
rect 7953 749 7992 755
rect 7956 721 7992 749
rect 8026 721 8065 755
rect 8099 721 8138 755
rect 8172 721 8211 755
rect 8245 721 8284 755
rect 8318 721 8357 755
rect 8391 721 8430 755
rect 8464 721 8503 755
rect 8537 721 8576 755
rect 8610 721 8649 755
rect 8683 721 8722 755
rect 8756 721 8795 755
rect 8829 721 8868 755
rect 8902 721 8941 755
rect 8975 721 8992 755
rect 9048 721 9056 755
rect 9267 721 9306 755
rect 9340 721 9379 755
rect 9413 721 9452 755
rect 9486 721 9525 755
rect 9559 721 9598 755
rect 9632 721 9671 755
rect 9705 721 9744 755
rect 9778 721 9817 755
rect 9851 721 9890 755
rect 9924 721 9963 755
rect 9997 721 10036 755
rect 10070 721 10109 755
rect 10143 721 10183 755
rect 10217 721 10257 755
rect 10291 721 10331 755
rect 10365 721 10405 755
rect 10439 721 10479 755
rect 10513 721 10553 755
rect 10587 721 10627 755
rect 10661 721 10701 755
rect 10735 721 10775 755
rect 10809 721 10849 755
rect 10883 721 10923 755
rect 10957 721 10969 755
rect 7956 715 8992 721
rect 7904 685 7956 697
tri 7956 690 7981 715 nw
tri 8980 709 8986 715 ne
rect 8986 709 8992 715
rect 9044 709 9056 721
rect 9108 709 9121 721
rect 9173 709 9186 721
rect 9238 715 10969 721
rect 9238 709 9244 715
tri 9244 709 9250 715 nw
tri 10898 709 10904 715 ne
rect 10904 709 10969 715
tri 10904 690 10923 709 ne
rect 10923 690 10969 709
rect 7904 621 7956 633
rect 7904 567 7913 569
rect 7947 567 7956 569
rect 7904 557 7956 567
rect 7904 493 7913 505
rect 7947 493 7956 505
rect 7904 436 7956 441
rect 7904 429 7913 436
rect 7947 429 7956 436
rect 7904 365 7956 377
tri 7956 353 7981 378 sw
tri 8980 353 8986 359 se
rect 8986 353 8992 359
rect 7956 347 8992 353
rect 7956 313 7985 347
rect 8019 313 8058 347
rect 8092 313 8131 347
rect 8165 313 8204 347
rect 8238 313 8277 347
rect 8311 313 8350 347
rect 8384 313 8423 347
rect 8457 313 8496 347
rect 8530 313 8569 347
rect 8603 313 8642 347
rect 8676 313 8715 347
rect 8749 313 8788 347
rect 8822 313 8861 347
rect 8895 313 8934 347
rect 8968 313 8992 347
rect 7904 307 8992 313
rect 9044 307 9056 359
rect 9108 347 9121 359
rect 9173 347 9186 359
rect 9238 353 9244 359
tri 9244 353 9250 359 sw
rect 9238 347 10923 353
rect 9115 313 9121 347
rect 9263 313 9303 347
rect 9337 313 9377 347
rect 9411 313 9451 347
rect 9485 313 9525 347
rect 9559 313 9599 347
rect 9633 313 9673 347
rect 9707 313 9747 347
rect 9781 313 9821 347
rect 9855 313 9895 347
rect 9929 313 9969 347
rect 10003 313 10043 347
rect 10077 313 10117 347
rect 10151 313 10191 347
rect 10225 313 10265 347
rect 10299 313 10339 347
rect 10373 313 10413 347
rect 10447 313 10487 347
rect 10521 313 10561 347
rect 10595 313 10635 347
rect 10669 313 10709 347
rect 10743 313 10783 347
rect 10817 313 10857 347
rect 10891 313 10923 347
rect 9108 307 9121 313
rect 9173 307 9186 313
rect 9238 307 10923 313
<< rmetal1 >>
rect 8718 5838 8720 5839
rect 8718 5788 8719 5838
rect 8718 5787 8720 5788
rect 8756 5838 8758 5839
rect 8757 5788 8758 5838
rect 8756 5787 8758 5788
rect 10672 5381 10674 5382
rect 10710 5381 10712 5382
rect 10208 5317 10210 5318
rect 10208 5267 10209 5317
rect 10208 5266 10210 5267
rect 10246 5317 10248 5318
rect 10247 5267 10248 5317
rect 10246 5266 10248 5267
rect 10672 5253 10673 5381
rect 10711 5253 10712 5381
rect 10672 5252 10674 5253
rect 10710 5252 10712 5253
rect 10523 4960 10525 4961
rect 10561 4960 10563 4961
rect 10523 4832 10524 4960
rect 10562 4832 10563 4960
rect 10523 4831 10525 4832
rect 10561 4831 10563 4832
rect 10523 4716 10525 4717
rect 10561 4716 10563 4717
rect 10523 4588 10524 4716
rect 10562 4588 10563 4716
rect 10523 4587 10525 4588
rect 10561 4587 10563 4588
rect 10679 4266 10681 4267
rect 10717 4266 10719 4267
rect 10679 4138 10680 4266
rect 10718 4138 10719 4266
rect 10679 4137 10681 4138
rect 10717 4137 10719 4138
<< via1 >>
rect 4320 6467 4372 6473
rect 4320 6433 4322 6467
rect 4322 6433 4356 6467
rect 4356 6433 4372 6467
rect 4320 6421 4372 6433
rect 4385 6467 4437 6473
rect 4385 6433 4394 6467
rect 4394 6433 4428 6467
rect 4428 6433 4437 6467
rect 4385 6421 4437 6433
rect 4450 6467 4502 6473
rect 4450 6433 4466 6467
rect 4466 6433 4500 6467
rect 4500 6433 4502 6467
rect 4450 6421 4502 6433
rect 4516 6467 4568 6473
rect 7589 6467 7641 6473
rect 4516 6433 4538 6467
rect 4538 6433 4568 6467
rect 7589 6433 7599 6467
rect 7599 6433 7633 6467
rect 7633 6433 7641 6467
rect 4516 6421 4568 6433
rect 7589 6421 7641 6433
rect 7653 6467 7705 6473
rect 7717 6467 7769 6473
rect 7653 6433 7672 6467
rect 7672 6433 7705 6467
rect 7717 6433 7745 6467
rect 7745 6433 7769 6467
rect 9693 6433 9716 6467
rect 9716 6433 9745 6467
rect 9757 6433 9789 6467
rect 9789 6433 9809 6467
rect 9821 6433 9823 6467
rect 9823 6433 9862 6467
rect 9862 6433 9873 6467
rect 7653 6421 7705 6433
rect 7717 6421 7769 6433
rect 9693 6415 9745 6433
rect 9757 6415 9809 6433
rect 9821 6415 9873 6433
rect 9693 6349 9745 6401
rect 9757 6349 9809 6401
rect 9821 6349 9873 6401
rect 1376 6100 1428 6106
rect 1458 6100 1510 6106
rect 1540 6100 1592 6106
rect 1622 6100 1674 6106
rect 1376 6066 1412 6100
rect 1412 6066 1428 6100
rect 1458 6066 1488 6100
rect 1488 6066 1510 6100
rect 1540 6066 1564 6100
rect 1564 6066 1592 6100
rect 1622 6066 1640 6100
rect 1640 6066 1674 6100
rect 1376 6054 1428 6066
rect 1458 6054 1510 6066
rect 1540 6054 1592 6066
rect 1622 6054 1674 6066
rect 9693 6283 9745 6335
rect 9757 6283 9809 6335
rect 9821 6283 9873 6335
rect 10226 6231 10278 6283
rect 10290 6231 10342 6283
rect 10968 6231 11020 6283
rect 11032 6232 11046 6283
rect 11046 6232 11084 6283
rect 11032 6231 11084 6232
rect 8668 6175 8720 6227
rect 8732 6175 8784 6227
rect 8836 6175 8888 6227
rect 8900 6175 8952 6227
rect 9437 6175 9489 6227
rect 9503 6175 9555 6227
rect 13112 6280 13164 6288
rect 13180 6280 13232 6288
rect 13112 6246 13134 6280
rect 13134 6246 13164 6280
rect 13180 6246 13206 6280
rect 13206 6246 13232 6280
rect 13112 6236 13164 6246
rect 13180 6236 13232 6246
rect 7913 6141 7965 6147
rect 7913 6107 7925 6141
rect 7925 6107 7959 6141
rect 7959 6107 7965 6141
rect 4757 6066 4759 6100
rect 4759 6066 4793 6100
rect 4793 6066 4809 6100
rect 4757 6048 4809 6066
rect 4821 6094 4873 6100
rect 4885 6094 4937 6100
rect 4821 6048 4831 6094
rect 4831 6048 4873 6094
rect 4885 6048 4937 6094
rect 7913 6095 7965 6107
rect 7979 6141 8031 6147
rect 8045 6141 8097 6147
rect 8111 6141 8163 6147
rect 8992 6141 9044 6153
rect 9056 6141 9108 6153
rect 9121 6141 9173 6153
rect 9186 6141 9238 6153
rect 7979 6107 7998 6141
rect 7998 6107 8031 6141
rect 8045 6107 8071 6141
rect 8071 6107 8097 6141
rect 8111 6107 8144 6141
rect 8144 6107 8163 6141
rect 8992 6107 9021 6141
rect 9021 6107 9044 6141
rect 9056 6107 9095 6141
rect 9095 6107 9108 6141
rect 9121 6107 9129 6141
rect 9129 6107 9169 6141
rect 9169 6107 9173 6141
rect 9186 6107 9203 6141
rect 9203 6107 9238 6141
rect 7979 6095 8031 6107
rect 8045 6095 8097 6107
rect 8111 6095 8163 6107
rect 8992 6101 9044 6107
rect 9056 6101 9108 6107
rect 9121 6101 9173 6107
rect 9186 6101 9238 6107
rect 7907 6069 7959 6075
rect 4757 5983 4809 6035
rect 4821 5983 4831 6035
rect 4831 5983 4873 6035
rect 4885 5983 4937 6035
rect 4757 5918 4809 5970
rect 4821 5918 4831 5970
rect 4831 5918 4873 5970
rect 4885 5918 4937 5970
rect 4757 5853 4809 5905
rect 4821 5853 4831 5905
rect 4831 5853 4873 5905
rect 4885 5853 4937 5905
rect 4757 5788 4809 5840
rect 4821 5788 4831 5840
rect 4831 5788 4873 5840
rect 4885 5788 4937 5840
rect 4757 5723 4809 5775
rect 4821 5723 4831 5775
rect 4831 5723 4873 5775
rect 4885 5723 4937 5775
rect 4757 5658 4809 5710
rect 4821 5658 4831 5710
rect 4831 5658 4873 5710
rect 4885 5658 4937 5710
rect 4757 5593 4809 5645
rect 4821 5593 4831 5645
rect 4831 5593 4873 5645
rect 4885 5593 4937 5645
rect 4757 5528 4809 5580
rect 4821 5528 4831 5580
rect 4831 5528 4873 5580
rect 4885 5528 4937 5580
rect 4757 5463 4809 5515
rect 4821 5463 4831 5515
rect 4831 5463 4873 5515
rect 4885 5463 4937 5515
rect 4757 5398 4809 5450
rect 4821 5398 4831 5450
rect 4831 5398 4873 5450
rect 4885 5398 4937 5450
rect 4757 5333 4809 5385
rect 4821 5333 4831 5385
rect 4831 5333 4873 5385
rect 4885 5333 4937 5385
rect 4757 5268 4809 5320
rect 4821 5268 4831 5320
rect 4831 5268 4873 5320
rect 4885 5268 4937 5320
rect 4757 5203 4809 5255
rect 4821 5203 4831 5255
rect 4831 5203 4873 5255
rect 4885 5203 4937 5255
rect 4757 5138 4809 5190
rect 4821 5138 4831 5190
rect 4831 5138 4873 5190
rect 4885 5138 4937 5190
rect 4757 5073 4809 5125
rect 4821 5073 4831 5125
rect 4831 5073 4873 5125
rect 4885 5073 4937 5125
rect 4757 5008 4809 5060
rect 4821 5008 4831 5060
rect 4831 5008 4873 5060
rect 4885 5008 4937 5060
rect 4757 4943 4809 4995
rect 4821 4943 4831 4995
rect 4831 4943 4873 4995
rect 4885 4943 4937 4995
rect 4757 4878 4809 4930
rect 4821 4878 4831 4930
rect 4831 4878 4873 4930
rect 4885 4878 4937 4930
rect 4757 4813 4809 4865
rect 4821 4813 4831 4865
rect 4831 4813 4873 4865
rect 4885 4813 4937 4865
rect 4757 4748 4809 4800
rect 4821 4748 4831 4800
rect 4831 4748 4873 4800
rect 4885 4748 4937 4800
rect 4757 4683 4809 4735
rect 4821 4683 4831 4735
rect 4831 4683 4873 4735
rect 4885 4683 4937 4735
rect 4757 4618 4809 4670
rect 4821 4618 4831 4670
rect 4831 4618 4873 4670
rect 4885 4618 4937 4670
rect 4757 4553 4809 4605
rect 4821 4553 4831 4605
rect 4831 4553 4873 4605
rect 4885 4553 4937 4605
rect 4757 4488 4809 4540
rect 4821 4488 4831 4540
rect 4831 4488 4873 4540
rect 4885 4488 4937 4540
rect 4757 4423 4809 4475
rect 4821 4423 4831 4475
rect 4831 4423 4873 4475
rect 4885 4423 4937 4475
rect 4757 4358 4809 4410
rect 4821 4358 4831 4410
rect 4831 4358 4873 4410
rect 4885 4358 4937 4410
rect 4757 4293 4809 4345
rect 4821 4293 4831 4345
rect 4831 4293 4873 4345
rect 4885 4293 4937 4345
rect 4757 4228 4809 4280
rect 4821 4228 4831 4280
rect 4831 4228 4873 4280
rect 4885 4228 4937 4280
rect 4757 4163 4809 4215
rect 4821 4163 4831 4215
rect 4831 4163 4873 4215
rect 4885 4163 4937 4215
rect 4757 4098 4809 4150
rect 4821 4098 4831 4150
rect 4831 4098 4873 4150
rect 4885 4098 4937 4150
rect 4757 4033 4809 4085
rect 4821 4044 4831 4085
rect 4831 4044 4873 4085
rect 4885 4044 4937 4085
rect 4821 4033 4873 4044
rect 4885 4033 4937 4044
rect 4757 3968 4809 4020
rect 4821 4005 4873 4020
rect 4821 3971 4831 4005
rect 4831 3971 4865 4005
rect 4865 3971 4873 4005
rect 4821 3968 4873 3971
rect 4885 4005 4937 4020
rect 4885 3971 4903 4005
rect 4903 3971 4937 4005
rect 4885 3968 4937 3971
rect 4757 3903 4809 3955
rect 4821 3932 4873 3955
rect 4821 3903 4831 3932
rect 4831 3903 4865 3932
rect 4865 3903 4873 3932
rect 4885 3932 4937 3955
rect 4885 3903 4903 3932
rect 4903 3903 4937 3932
rect 4757 3859 4937 3890
rect 4757 3825 4831 3859
rect 4831 3825 4865 3859
rect 4865 3825 4903 3859
rect 4903 3825 4937 3859
rect 4757 3786 4937 3825
rect 4757 3752 4831 3786
rect 4831 3752 4865 3786
rect 4865 3752 4903 3786
rect 4903 3752 4937 3786
rect 4757 3713 4937 3752
rect 4757 3679 4831 3713
rect 4831 3679 4865 3713
rect 4865 3679 4903 3713
rect 4903 3679 4937 3713
rect 4757 3640 4937 3679
rect 4757 3606 4831 3640
rect 4831 3606 4865 3640
rect 4865 3606 4903 3640
rect 4903 3606 4937 3640
rect 1376 3544 1428 3596
rect 1441 3544 1493 3596
rect 1506 3544 1558 3596
rect 1572 3544 1624 3596
rect 1638 3544 1690 3596
rect 4757 3567 4937 3606
rect 4757 3533 4831 3567
rect 4831 3533 4865 3567
rect 4865 3533 4903 3567
rect 4903 3533 4937 3567
rect 1376 3488 1428 3532
rect 1441 3488 1493 3532
rect 1506 3488 1558 3532
rect 1572 3488 1624 3532
rect 1638 3488 1690 3532
rect 4757 3494 4937 3533
rect 7907 6035 7913 6069
rect 7913 6035 7947 6069
rect 7947 6035 7959 6069
rect 7907 6023 7959 6035
rect 8598 6021 8650 6073
rect 8662 6021 8714 6073
rect 6932 4203 6984 4208
rect 6932 4169 6941 4203
rect 6941 4169 6975 4203
rect 6975 4169 6984 4203
rect 6932 4156 6984 4169
rect 6932 4130 6984 4142
rect 6932 4096 6941 4130
rect 6941 4096 6975 4130
rect 6975 4096 6984 4130
rect 6932 4090 6984 4096
rect 7592 6008 7644 6014
rect 7592 5974 7623 6008
rect 7623 5974 7644 6008
rect 7592 5962 7644 5974
rect 7656 6008 7708 6014
rect 7656 5974 7661 6008
rect 7661 5974 7695 6008
rect 7695 5974 7708 6008
rect 7656 5962 7708 5974
rect 7720 6008 7772 6014
rect 7720 5974 7733 6008
rect 7733 5974 7767 6008
rect 7767 5974 7772 6008
rect 7720 5962 7772 5974
rect 7592 5932 7644 5949
rect 7592 5898 7623 5932
rect 7623 5898 7644 5932
rect 7592 5897 7644 5898
rect 7656 5932 7708 5949
rect 7656 5898 7661 5932
rect 7661 5898 7695 5932
rect 7695 5898 7708 5932
rect 7656 5897 7708 5898
rect 7720 5932 7772 5949
rect 7720 5898 7733 5932
rect 7733 5898 7767 5932
rect 7767 5898 7772 5932
rect 7720 5897 7772 5898
rect 7592 5856 7644 5884
rect 7592 5832 7623 5856
rect 7623 5832 7644 5856
rect 7656 5856 7708 5884
rect 7656 5832 7661 5856
rect 7661 5832 7695 5856
rect 7695 5832 7708 5856
rect 7720 5856 7772 5884
rect 7720 5832 7733 5856
rect 7733 5832 7767 5856
rect 7767 5832 7772 5856
rect 7592 5780 7644 5819
rect 7592 5767 7623 5780
rect 7623 5767 7644 5780
rect 7656 5780 7708 5819
rect 7656 5767 7661 5780
rect 7661 5767 7695 5780
rect 7695 5767 7708 5780
rect 7720 5780 7772 5819
rect 7720 5767 7733 5780
rect 7733 5767 7767 5780
rect 7767 5767 7772 5780
rect 7592 5746 7623 5754
rect 7623 5746 7644 5754
rect 7592 5704 7644 5746
rect 7592 5702 7623 5704
rect 7623 5702 7644 5704
rect 7656 5746 7661 5754
rect 7661 5746 7695 5754
rect 7695 5746 7708 5754
rect 7656 5704 7708 5746
rect 7656 5702 7661 5704
rect 7661 5702 7695 5704
rect 7695 5702 7708 5704
rect 7720 5746 7733 5754
rect 7733 5746 7767 5754
rect 7767 5746 7772 5754
rect 7720 5704 7772 5746
rect 7720 5702 7733 5704
rect 7733 5702 7767 5704
rect 7767 5702 7772 5704
rect 7592 5670 7623 5689
rect 7623 5670 7644 5689
rect 7592 5637 7644 5670
rect 7656 5670 7661 5689
rect 7661 5670 7695 5689
rect 7695 5670 7708 5689
rect 7656 5637 7708 5670
rect 7720 5670 7733 5689
rect 7733 5670 7767 5689
rect 7767 5670 7772 5689
rect 7720 5637 7772 5670
rect 7592 5594 7623 5624
rect 7623 5594 7644 5624
rect 7592 5572 7644 5594
rect 7656 5594 7661 5624
rect 7661 5594 7695 5624
rect 7695 5594 7708 5624
rect 7656 5572 7708 5594
rect 7720 5594 7733 5624
rect 7733 5594 7767 5624
rect 7767 5594 7772 5624
rect 7720 5572 7772 5594
rect 7592 5552 7644 5558
rect 7592 5518 7623 5552
rect 7623 5518 7644 5552
rect 7592 5506 7644 5518
rect 7656 5552 7708 5558
rect 7656 5518 7661 5552
rect 7661 5518 7695 5552
rect 7695 5518 7708 5552
rect 7656 5506 7708 5518
rect 7720 5552 7772 5558
rect 7720 5518 7733 5552
rect 7733 5518 7767 5552
rect 7767 5518 7772 5552
rect 7720 5506 7772 5518
rect 7592 5477 7644 5492
rect 7592 5443 7623 5477
rect 7623 5443 7644 5477
rect 7592 5440 7644 5443
rect 7656 5477 7708 5492
rect 7656 5443 7661 5477
rect 7661 5443 7695 5477
rect 7695 5443 7708 5477
rect 7656 5440 7708 5443
rect 7720 5477 7772 5492
rect 7720 5443 7733 5477
rect 7733 5443 7767 5477
rect 7767 5443 7772 5477
rect 7720 5440 7772 5443
rect 7592 5402 7644 5426
rect 7592 5374 7623 5402
rect 7623 5374 7644 5402
rect 7656 5402 7708 5426
rect 7656 5374 7661 5402
rect 7661 5374 7695 5402
rect 7695 5374 7708 5402
rect 7720 5402 7772 5426
rect 7720 5374 7733 5402
rect 7733 5374 7767 5402
rect 7767 5374 7772 5402
rect 7592 5327 7644 5360
rect 7592 5308 7623 5327
rect 7623 5308 7644 5327
rect 7656 5327 7708 5360
rect 7656 5308 7661 5327
rect 7661 5308 7695 5327
rect 7695 5308 7708 5327
rect 7720 5327 7772 5360
rect 7720 5308 7733 5327
rect 7733 5308 7767 5327
rect 7767 5308 7772 5327
rect 7592 5293 7623 5294
rect 7623 5293 7644 5294
rect 7592 5252 7644 5293
rect 7592 5242 7623 5252
rect 7623 5242 7644 5252
rect 7656 5293 7661 5294
rect 7661 5293 7695 5294
rect 7695 5293 7708 5294
rect 7656 5252 7708 5293
rect 7656 5242 7661 5252
rect 7661 5242 7695 5252
rect 7695 5242 7708 5252
rect 7720 5293 7733 5294
rect 7733 5293 7767 5294
rect 7767 5293 7772 5294
rect 7720 5252 7772 5293
rect 7720 5242 7733 5252
rect 7733 5242 7767 5252
rect 7767 5242 7772 5252
rect 7592 5218 7623 5228
rect 7623 5218 7644 5228
rect 7592 5177 7644 5218
rect 7592 5176 7623 5177
rect 7623 5176 7644 5177
rect 7656 5218 7661 5228
rect 7661 5218 7695 5228
rect 7695 5218 7708 5228
rect 7656 5177 7708 5218
rect 7656 5176 7661 5177
rect 7661 5176 7695 5177
rect 7695 5176 7708 5177
rect 7720 5218 7733 5228
rect 7733 5218 7767 5228
rect 7767 5218 7772 5228
rect 7720 5177 7772 5218
rect 7720 5176 7733 5177
rect 7733 5176 7767 5177
rect 7767 5176 7772 5177
rect 7592 5143 7623 5162
rect 7623 5143 7644 5162
rect 7592 5110 7644 5143
rect 7656 5143 7661 5162
rect 7661 5143 7695 5162
rect 7695 5143 7708 5162
rect 7656 5110 7708 5143
rect 7720 5143 7733 5162
rect 7733 5143 7767 5162
rect 7767 5143 7772 5162
rect 7720 5110 7772 5143
rect 7592 5068 7623 5096
rect 7623 5068 7644 5096
rect 7592 5044 7644 5068
rect 7656 5068 7661 5096
rect 7661 5068 7695 5096
rect 7695 5068 7708 5096
rect 7656 5044 7708 5068
rect 7720 5068 7733 5096
rect 7733 5068 7767 5096
rect 7767 5068 7772 5096
rect 7720 5044 7772 5068
rect 7592 5027 7644 5030
rect 7592 4993 7623 5027
rect 7623 4993 7644 5027
rect 7592 4978 7644 4993
rect 7656 5027 7708 5030
rect 7656 4993 7661 5027
rect 7661 4993 7695 5027
rect 7695 4993 7708 5027
rect 7656 4978 7708 4993
rect 7720 5027 7772 5030
rect 7720 4993 7733 5027
rect 7733 4993 7767 5027
rect 7767 4993 7772 5027
rect 7720 4978 7772 4993
rect 7592 4952 7644 4964
rect 7592 4918 7623 4952
rect 7623 4918 7644 4952
rect 7592 4912 7644 4918
rect 7656 4952 7708 4964
rect 7656 4918 7661 4952
rect 7661 4918 7695 4952
rect 7695 4918 7708 4952
rect 7656 4912 7708 4918
rect 7720 4952 7772 4964
rect 7720 4918 7733 4952
rect 7733 4918 7767 4952
rect 7767 4918 7772 4952
rect 7720 4912 7772 4918
rect 7907 5993 7959 6010
rect 7907 5959 7913 5993
rect 7913 5959 7947 5993
rect 7947 5959 7959 5993
rect 7907 5958 7959 5959
rect 7907 5917 7959 5945
rect 8203 5984 8255 5993
rect 8269 5984 8321 5993
rect 8203 5950 8215 5984
rect 8215 5950 8255 5984
rect 8269 5950 8293 5984
rect 8293 5950 8321 5984
rect 8203 5941 8255 5950
rect 8269 5941 8321 5950
rect 8836 5941 8888 5993
rect 8900 5984 8952 5993
rect 8900 5950 8933 5984
rect 8933 5950 8952 5984
rect 9757 5982 9764 6080
rect 9764 5982 9870 6080
rect 9870 5982 9873 6080
rect 9757 5964 9873 5982
rect 8900 5941 8952 5950
rect 7907 5893 7913 5917
rect 7913 5893 7947 5917
rect 7947 5893 7959 5917
rect 7907 5841 7959 5880
rect 8460 5867 8512 5919
rect 8527 5867 8579 5919
rect 7907 5828 7913 5841
rect 7913 5828 7947 5841
rect 7947 5828 7959 5841
rect 7907 5807 7913 5815
rect 7913 5807 7947 5815
rect 7947 5807 7959 5815
rect 7907 5765 7959 5807
rect 8277 5828 8329 5834
rect 8343 5828 8395 5834
rect 8277 5794 8289 5828
rect 8289 5794 8329 5828
rect 8343 5794 8370 5828
rect 8370 5794 8395 5828
rect 8277 5782 8329 5794
rect 8343 5782 8395 5794
rect 10386 5787 10438 5839
rect 10450 5787 10502 5839
rect 7907 5763 7913 5765
rect 7913 5763 7947 5765
rect 7947 5763 7959 5765
rect 7907 5731 7913 5750
rect 7913 5731 7947 5750
rect 7947 5731 7959 5750
rect 7907 5698 7959 5731
rect 8518 5707 8570 5759
rect 8582 5707 8634 5759
rect 11584 5792 11636 5804
rect 11584 5758 11588 5792
rect 11588 5758 11622 5792
rect 11622 5758 11636 5792
rect 11584 5752 11636 5758
rect 11648 5752 11700 5804
rect 7907 5655 7913 5685
rect 7913 5655 7947 5685
rect 7947 5655 7959 5685
rect 7907 5633 7959 5655
rect 8203 5672 8255 5681
rect 8269 5672 8321 5681
rect 8203 5638 8221 5672
rect 8221 5638 8255 5672
rect 8269 5638 8302 5672
rect 8302 5638 8321 5672
rect 8203 5629 8255 5638
rect 8269 5629 8321 5638
rect 8756 5629 8808 5681
rect 8820 5672 8872 5681
rect 8820 5638 8864 5672
rect 8864 5638 8872 5672
rect 8820 5629 8872 5638
rect 7907 5613 7959 5620
rect 7907 5579 7913 5613
rect 7913 5579 7947 5613
rect 7947 5579 7959 5613
rect 9528 5600 9580 5652
rect 9594 5600 9646 5652
rect 7907 5568 7959 5579
rect 7907 5536 7959 5555
rect 7907 5503 7913 5536
rect 7913 5503 7947 5536
rect 7947 5503 7959 5536
rect 7907 5459 7959 5489
rect 8277 5516 8329 5526
rect 8343 5516 8395 5526
rect 10466 5520 10518 5572
rect 10530 5520 10582 5572
rect 8277 5482 8289 5516
rect 8289 5482 8329 5516
rect 8343 5482 8370 5516
rect 8370 5482 8395 5516
rect 8277 5474 8329 5482
rect 8343 5474 8395 5482
rect 7907 5437 7913 5459
rect 7913 5437 7947 5459
rect 7947 5437 7959 5459
rect 9278 5438 9330 5490
rect 9344 5438 9396 5490
rect 7907 5382 7959 5423
rect 7907 5371 7913 5382
rect 7913 5371 7947 5382
rect 7947 5371 7959 5382
rect 8992 5386 9044 5398
rect 9056 5386 9108 5398
rect 9121 5386 9173 5398
rect 9186 5386 9238 5398
rect 7907 5348 7913 5357
rect 7913 5348 7947 5357
rect 7947 5348 7959 5357
rect 7907 5305 7959 5348
rect 8203 5360 8255 5372
rect 8269 5360 8321 5372
rect 8203 5326 8218 5360
rect 8218 5326 8255 5360
rect 8269 5326 8297 5360
rect 8297 5326 8321 5360
rect 8992 5352 9012 5386
rect 9012 5352 9044 5386
rect 9056 5352 9087 5386
rect 9087 5352 9108 5386
rect 9121 5352 9162 5386
rect 9162 5352 9173 5386
rect 9186 5352 9196 5386
rect 9196 5352 9237 5386
rect 9237 5352 9238 5386
rect 8992 5346 9044 5352
rect 9056 5346 9108 5352
rect 9121 5346 9173 5352
rect 9186 5346 9238 5352
rect 8203 5320 8255 5326
rect 8269 5320 8321 5326
rect 10300 5323 10352 5375
rect 7907 5271 7913 5291
rect 7913 5271 7947 5291
rect 7947 5271 7959 5291
rect 7907 5239 7959 5271
rect 7907 5194 7913 5225
rect 7913 5194 7947 5225
rect 7947 5194 7959 5225
rect 8435 5250 8487 5259
rect 8502 5250 8554 5259
rect 8435 5216 8440 5250
rect 8440 5216 8482 5250
rect 8482 5216 8487 5250
rect 8502 5216 8516 5250
rect 8516 5216 8554 5250
rect 8435 5207 8487 5216
rect 8502 5207 8554 5216
rect 10300 5258 10352 5310
rect 8674 5210 8726 5219
rect 7907 5173 7959 5194
rect 8674 5176 8706 5210
rect 8706 5176 8726 5210
rect 8674 5167 8726 5176
rect 8740 5167 8792 5219
rect 9278 5210 9330 5221
rect 9344 5210 9396 5221
rect 9278 5176 9297 5210
rect 9297 5176 9330 5210
rect 9344 5176 9377 5210
rect 9377 5176 9396 5210
rect 9278 5169 9330 5176
rect 9344 5169 9396 5176
rect 8754 5060 8806 5112
rect 8820 5100 8872 5112
rect 8820 5066 8862 5100
rect 8862 5066 8872 5100
rect 8820 5060 8872 5066
rect 7913 4997 7965 5003
rect 7913 4963 7947 4997
rect 7947 4963 7965 4997
rect 7913 4951 7965 4963
rect 7979 4994 8031 5003
rect 8045 4994 8097 5003
rect 7979 4960 8029 4994
rect 8029 4960 8031 4994
rect 8045 4960 8063 4994
rect 8063 4960 8097 4994
rect 7979 4951 8031 4960
rect 8045 4951 8097 4960
rect 8111 4994 8163 5003
rect 8111 4960 8145 4994
rect 8145 4960 8163 4994
rect 8111 4951 8163 4960
rect 8515 4951 8567 5003
rect 8582 4951 8634 5003
rect 8992 4924 9044 4936
rect 9056 4924 9108 4936
rect 9121 4924 9173 4936
rect 9186 4924 9238 4936
rect 8992 4890 9017 4924
rect 9017 4890 9044 4924
rect 9056 4890 9092 4924
rect 9092 4890 9108 4924
rect 9121 4890 9126 4924
rect 9126 4890 9167 4924
rect 9167 4890 9173 4924
rect 9186 4890 9201 4924
rect 9201 4890 9238 4924
rect 8992 4884 9044 4890
rect 9056 4884 9108 4890
rect 9121 4884 9173 4890
rect 9186 4884 9238 4890
rect 9693 5226 9745 5232
rect 9757 5226 9809 5232
rect 9821 5226 9873 5232
rect 9693 5192 9734 5226
rect 9734 5192 9745 5226
rect 9757 5192 9768 5226
rect 9768 5192 9806 5226
rect 9806 5192 9809 5226
rect 9821 5192 9840 5226
rect 9840 5192 9873 5226
rect 9693 5180 9745 5192
rect 9757 5180 9809 5192
rect 9821 5180 9873 5192
rect 9693 5151 9745 5159
rect 9757 5151 9809 5159
rect 9821 5151 9873 5159
rect 9693 5117 9734 5151
rect 9734 5117 9745 5151
rect 9757 5117 9768 5151
rect 9768 5117 9806 5151
rect 9806 5117 9809 5151
rect 9821 5117 9840 5151
rect 9840 5117 9873 5151
rect 9693 5107 9745 5117
rect 9757 5107 9809 5117
rect 9821 5107 9873 5117
rect 9693 5076 9745 5086
rect 9757 5076 9809 5086
rect 9821 5076 9873 5086
rect 9693 5042 9734 5076
rect 9734 5042 9745 5076
rect 9757 5042 9768 5076
rect 9768 5042 9806 5076
rect 9806 5042 9809 5076
rect 9821 5042 9840 5076
rect 9840 5042 9873 5076
rect 9693 5034 9745 5042
rect 9757 5034 9809 5042
rect 9821 5034 9873 5042
rect 9693 5001 9745 5013
rect 9757 5001 9809 5013
rect 9821 5001 9873 5013
rect 9693 4967 9734 5001
rect 9734 4967 9745 5001
rect 9757 4967 9768 5001
rect 9768 4967 9806 5001
rect 9806 4967 9809 5001
rect 9821 4967 9840 5001
rect 9840 4967 9873 5001
rect 9693 4961 9745 4967
rect 9757 4961 9809 4967
rect 9821 4961 9873 4967
rect 9693 4927 9745 4939
rect 9757 4927 9809 4939
rect 9821 4927 9873 4939
rect 9693 4893 9734 4927
rect 9734 4893 9745 4927
rect 9757 4893 9768 4927
rect 9768 4893 9806 4927
rect 9806 4893 9809 4927
rect 9821 4893 9840 4927
rect 9840 4893 9873 4927
rect 9693 4887 9745 4893
rect 9757 4887 9809 4893
rect 9821 4887 9873 4893
rect 10380 4882 10432 4934
rect 7347 4820 7399 4872
rect 7411 4820 7463 4872
rect 7475 4820 7527 4872
rect 8225 4820 8277 4872
rect 8289 4820 8341 4872
rect 8353 4820 8405 4872
rect 7347 4754 7399 4806
rect 7411 4754 7463 4806
rect 7475 4754 7527 4806
rect 8225 4784 8226 4806
rect 8226 4784 8273 4806
rect 8273 4784 8277 4806
rect 8289 4784 8307 4806
rect 8307 4784 8341 4806
rect 8225 4754 8277 4784
rect 8289 4754 8341 4784
rect 8353 4784 8354 4806
rect 8354 4784 8388 4806
rect 8388 4784 8405 4806
rect 10380 4816 10432 4868
rect 8353 4754 8405 4784
rect 8754 4748 8806 4757
rect 8820 4748 8872 4757
rect 7042 4203 7094 4208
rect 7042 4169 7051 4203
rect 7051 4169 7085 4203
rect 7085 4169 7094 4203
rect 7042 4156 7094 4169
rect 7042 4130 7094 4142
rect 7042 4096 7051 4130
rect 7051 4096 7085 4130
rect 7085 4096 7094 4130
rect 7042 4090 7094 4096
rect 8754 4714 8787 4748
rect 8787 4714 8806 4748
rect 8820 4714 8821 4748
rect 8821 4714 8872 4748
rect 8754 4705 8806 4714
rect 8820 4705 8872 4714
rect 9361 4748 9413 4754
rect 9361 4714 9385 4748
rect 9385 4714 9413 4748
rect 9361 4702 9413 4714
rect 9427 4702 9479 4754
rect 7592 4634 7644 4640
rect 7656 4634 7708 4640
rect 7720 4634 7772 4640
rect 7592 4588 7644 4634
rect 7656 4588 7708 4634
rect 7720 4588 7767 4634
rect 7767 4588 7772 4634
rect 7913 4636 7965 4651
rect 7592 4517 7644 4569
rect 7656 4517 7708 4569
rect 7720 4517 7767 4569
rect 7767 4517 7772 4569
rect 7592 4446 7644 4498
rect 7656 4446 7708 4498
rect 7720 4446 7767 4498
rect 7767 4446 7772 4498
rect 7592 4375 7644 4427
rect 7656 4375 7708 4427
rect 7720 4375 7767 4427
rect 7767 4375 7772 4427
rect 7592 4304 7644 4356
rect 7656 4304 7708 4356
rect 7720 4304 7767 4356
rect 7767 4304 7772 4356
rect 7592 4233 7644 4285
rect 7656 4233 7708 4285
rect 7720 4233 7767 4285
rect 7767 4233 7772 4285
rect 7592 4162 7644 4214
rect 7656 4162 7708 4214
rect 7720 4162 7767 4214
rect 7767 4162 7772 4214
rect 7592 4096 7644 4142
rect 7656 4096 7708 4142
rect 7720 4096 7767 4142
rect 7767 4096 7772 4142
rect 7592 4090 7644 4096
rect 7656 4090 7708 4096
rect 7720 4090 7772 4096
rect 7913 4602 7947 4636
rect 7947 4602 7965 4636
rect 7913 4599 7965 4602
rect 7979 4642 8031 4651
rect 8045 4642 8097 4651
rect 8111 4642 8163 4651
rect 7979 4608 8029 4642
rect 8029 4608 8031 4642
rect 8045 4608 8063 4642
rect 8063 4608 8097 4642
rect 8111 4608 8144 4642
rect 8144 4608 8163 4642
rect 8992 4620 9044 4672
rect 9056 4620 9108 4672
rect 9121 4620 9173 4672
rect 9186 4620 9238 4672
rect 7979 4599 8031 4608
rect 8045 4599 8097 4608
rect 8111 4599 8163 4608
rect 8834 4572 8886 4578
rect 8900 4572 8952 4578
rect 8834 4538 8867 4572
rect 8867 4538 8886 4572
rect 8900 4538 8901 4572
rect 8901 4538 8948 4572
rect 8948 4538 8952 4572
rect 8834 4526 8886 4538
rect 8900 4526 8952 4538
rect 9693 4745 9745 4751
rect 9757 4745 9809 4751
rect 9821 4745 9873 4751
rect 9693 4711 9734 4745
rect 9734 4711 9745 4745
rect 9757 4711 9768 4745
rect 9768 4711 9806 4745
rect 9806 4711 9809 4745
rect 9821 4711 9840 4745
rect 9840 4711 9873 4745
rect 11692 4748 11744 4800
rect 11756 4748 11808 4800
rect 9693 4699 9745 4711
rect 9757 4699 9809 4711
rect 9821 4699 9873 4711
rect 10380 4684 10432 4736
rect 9693 4658 9745 4667
rect 9757 4658 9809 4667
rect 9821 4658 9873 4667
rect 9693 4624 9734 4658
rect 9734 4624 9745 4658
rect 9757 4624 9768 4658
rect 9768 4624 9806 4658
rect 9806 4624 9809 4658
rect 9821 4624 9840 4658
rect 9840 4624 9873 4658
rect 9693 4615 9745 4624
rect 9757 4615 9809 4624
rect 9821 4615 9873 4624
rect 10380 4618 10432 4670
rect 9693 4571 9745 4583
rect 9757 4571 9809 4583
rect 9821 4571 9873 4583
rect 9693 4537 9734 4571
rect 9734 4537 9745 4571
rect 9757 4537 9768 4571
rect 9768 4537 9806 4571
rect 9806 4537 9809 4571
rect 9821 4537 9840 4571
rect 9840 4537 9873 4571
rect 9693 4531 9745 4537
rect 9757 4531 9809 4537
rect 9821 4531 9873 4537
rect 10220 4523 10272 4575
rect 10220 4457 10272 4509
rect 8515 4386 8567 4395
rect 8582 4386 8634 4395
rect 8515 4352 8550 4386
rect 8550 4352 8567 4386
rect 8582 4352 8584 4386
rect 8584 4352 8634 4386
rect 8515 4343 8567 4352
rect 8582 4343 8634 4352
rect 9361 4416 9413 4422
rect 9361 4382 9385 4416
rect 9385 4382 9413 4416
rect 9361 4370 9413 4382
rect 9427 4370 9479 4422
rect 9693 4411 9745 4417
rect 9757 4411 9809 4417
rect 9821 4411 9873 4417
rect 9693 4377 9734 4411
rect 9734 4377 9745 4411
rect 9757 4377 9768 4411
rect 9768 4377 9806 4411
rect 9806 4377 9809 4411
rect 9821 4377 9840 4411
rect 9840 4377 9873 4411
rect 9693 4365 9745 4377
rect 9757 4365 9809 4377
rect 9821 4365 9873 4377
rect 9693 4317 9745 4349
rect 9757 4317 9809 4349
rect 9821 4317 9873 4349
rect 9361 4306 9413 4312
rect 9361 4272 9385 4306
rect 9385 4272 9413 4306
rect 9361 4260 9413 4272
rect 9427 4260 9479 4312
rect 9522 4258 9574 4310
rect 9522 4192 9574 4244
rect 9693 4297 9734 4317
rect 9734 4297 9745 4317
rect 9757 4297 9768 4317
rect 9768 4297 9806 4317
rect 9806 4297 9809 4317
rect 9821 4297 9840 4317
rect 9840 4297 9873 4317
rect 9693 4228 9745 4280
rect 9757 4228 9809 4280
rect 9821 4228 9873 4280
rect 9693 4189 9734 4211
rect 9734 4189 9745 4211
rect 9757 4189 9768 4211
rect 9768 4189 9806 4211
rect 9806 4189 9809 4211
rect 9821 4189 9840 4211
rect 9840 4189 9873 4211
rect 9693 4159 9745 4189
rect 9757 4159 9809 4189
rect 9821 4159 9873 4189
rect 10300 4209 10352 4261
rect 8754 4084 8806 4136
rect 8820 4084 8872 4136
rect 8992 4130 9044 4136
rect 8992 4096 9025 4130
rect 9025 4096 9044 4130
rect 8992 4084 9044 4096
rect 9056 4130 9108 4136
rect 9056 4096 9063 4130
rect 9063 4096 9097 4130
rect 9097 4096 9108 4130
rect 9056 4084 9108 4096
rect 9121 4130 9173 4136
rect 9121 4096 9135 4130
rect 9135 4096 9169 4130
rect 9169 4096 9173 4130
rect 9121 4084 9173 4096
rect 9186 4130 9238 4136
rect 9186 4096 9207 4130
rect 9207 4096 9238 4130
rect 9186 4084 9238 4096
rect 9693 4130 9745 4142
rect 9757 4130 9809 4142
rect 9821 4130 9873 4142
rect 10300 4143 10352 4195
rect 9693 4096 9734 4130
rect 9734 4096 9745 4130
rect 9757 4096 9768 4130
rect 9768 4096 9806 4130
rect 9806 4096 9809 4130
rect 9821 4096 9840 4130
rect 9840 4096 9873 4130
rect 9693 4090 9745 4096
rect 9757 4090 9809 4096
rect 9821 4090 9873 4096
rect 7167 4004 7219 4056
rect 7233 4004 7285 4056
rect 7299 4004 7351 4056
rect 7167 3940 7219 3992
rect 7233 3940 7285 3992
rect 7299 3940 7351 3992
rect 8508 3964 8560 4016
rect 8574 3964 8626 4016
rect 10554 4029 10606 4081
rect 10618 4071 10670 4081
rect 10618 4037 10663 4071
rect 10663 4037 10670 4071
rect 10618 4029 10670 4037
rect 9359 3954 9411 3960
rect 7913 3924 7965 3936
rect 6852 3852 6904 3904
rect 7913 3890 7947 3924
rect 7947 3890 7965 3924
rect 6852 3820 6904 3838
rect 6852 3786 6886 3820
rect 6886 3786 6904 3820
rect 7913 3884 7965 3890
rect 7979 3924 8031 3936
rect 8045 3924 8097 3936
rect 8111 3924 8163 3936
rect 7979 3890 8029 3924
rect 8029 3890 8031 3924
rect 8045 3890 8063 3924
rect 8063 3890 8097 3924
rect 8111 3890 8138 3924
rect 8138 3890 8163 3924
rect 7979 3884 8031 3890
rect 8045 3884 8097 3890
rect 8111 3884 8163 3890
rect 9359 3920 9385 3954
rect 9385 3920 9411 3954
rect 7592 3816 7623 3827
rect 7623 3816 7644 3827
rect 7592 3775 7644 3816
rect 7656 3816 7661 3827
rect 7661 3816 7695 3827
rect 7695 3816 7708 3827
rect 7656 3775 7708 3816
rect 7720 3816 7733 3827
rect 7733 3816 7767 3827
rect 7767 3816 7772 3827
rect 7720 3775 7772 3816
rect 9359 3908 9411 3920
rect 9425 3908 9477 3960
rect 9680 3897 9732 3949
rect 9744 3943 9796 3949
rect 9808 3943 9860 3949
rect 9744 3897 9796 3943
rect 9808 3897 9860 3943
rect 9278 3820 9330 3872
rect 9344 3820 9396 3872
rect 9680 3831 9732 3883
rect 9744 3837 9796 3883
rect 9808 3837 9860 3883
rect 9744 3831 9796 3837
rect 9808 3831 9860 3837
rect 8754 3732 8806 3784
rect 8820 3778 8872 3784
rect 8820 3744 8867 3778
rect 8867 3744 8872 3778
rect 8820 3732 8872 3744
rect 10968 3735 11020 3787
rect 11032 3735 11084 3787
rect 12450 3779 12502 3831
rect 12516 3779 12568 3831
rect 13034 3779 13086 3831
rect 13100 3779 13152 3831
rect 10554 3657 10606 3709
rect 10618 3657 10670 3709
rect 9361 3602 9413 3608
rect 9361 3568 9388 3602
rect 9388 3568 9413 3602
rect 9361 3556 9413 3568
rect 9427 3556 9479 3608
rect 11800 3671 11852 3723
rect 11866 3671 11918 3723
rect 11800 3607 11852 3659
rect 11866 3607 11918 3659
rect 13843 3607 13959 3723
rect 4757 3488 4831 3494
rect 1376 3480 1378 3488
rect 1378 3480 1417 3488
rect 1417 3480 1428 3488
rect 1441 3480 1451 3488
rect 1451 3480 1490 3488
rect 1490 3480 1493 3488
rect 1506 3480 1524 3488
rect 1524 3480 1558 3488
rect 1572 3480 1597 3488
rect 1597 3480 1624 3488
rect 1638 3480 1670 3488
rect 1670 3480 1690 3488
rect 4757 3454 4759 3488
rect 4759 3454 4793 3488
rect 4793 3460 4831 3488
rect 4831 3460 4865 3494
rect 4865 3460 4903 3494
rect 4903 3460 4937 3494
rect 4793 3454 4937 3460
rect 7913 3517 7965 3523
rect 7913 3483 7947 3517
rect 7947 3483 7965 3517
rect 7913 3471 7965 3483
rect 7979 3471 8031 3523
rect 8045 3471 8097 3523
rect 8111 3471 8163 3523
rect 11986 3499 12038 3551
rect 12052 3499 12104 3551
rect 4320 3356 4372 3408
rect 4385 3356 4437 3408
rect 4450 3356 4502 3408
rect 4516 3356 4568 3408
rect 4320 3292 4372 3344
rect 4385 3292 4437 3344
rect 4450 3292 4502 3344
rect 4516 3292 4568 3344
rect 7048 3368 7100 3420
rect 7114 3368 7166 3420
rect 9450 3391 9502 3443
rect 9516 3391 9568 3443
rect 9686 3391 9738 3443
rect 9750 3431 9802 3443
rect 9750 3397 9784 3431
rect 9784 3397 9802 3431
rect 9750 3391 9802 3397
rect 9815 3431 9867 3443
rect 11986 3435 12038 3487
rect 12052 3435 12104 3487
rect 14029 3435 14145 3551
rect 9815 3397 9825 3431
rect 9825 3397 9859 3431
rect 9859 3397 9867 3431
rect 9815 3391 9867 3397
rect 4320 3228 4372 3280
rect 4385 3228 4437 3280
rect 4450 3228 4502 3280
rect 4516 3228 4568 3280
rect 6949 3288 7001 3340
rect 7015 3288 7067 3340
rect 8507 3311 8559 3363
rect 8571 3311 8623 3363
rect 11508 3311 11560 3363
rect 11572 3311 11624 3363
rect 6858 3208 6910 3260
rect 6924 3208 6976 3260
rect 9418 2997 9470 3049
rect 9482 2997 9534 3049
rect 10330 2997 10382 3049
rect 10394 2997 10446 3049
rect 11616 2997 11668 3049
rect 11680 2997 11732 3049
rect 13619 2921 13671 2973
rect 13685 2921 13737 2973
rect 13751 2921 13803 2973
rect 13817 2921 13869 2973
rect 13883 2921 13935 2973
rect 13949 2921 14001 2973
rect 14015 2921 14067 2973
rect 8587 2911 8639 2917
rect 8587 2877 8604 2911
rect 8604 2877 8638 2911
rect 8638 2877 8639 2911
rect 8587 2865 8639 2877
rect 8653 2911 8705 2917
rect 8653 2877 8680 2911
rect 8680 2877 8705 2911
rect 8653 2865 8705 2877
rect 13619 2857 13671 2909
rect 13685 2857 13737 2909
rect 13751 2857 13803 2909
rect 13817 2857 13869 2909
rect 13883 2857 13935 2909
rect 13949 2857 14001 2909
rect 14015 2857 14067 2909
rect 7904 2798 7956 2825
rect 7904 2773 7913 2798
rect 7913 2773 7947 2798
rect 7947 2773 7956 2798
rect 7904 2725 7956 2760
rect 7904 2708 7913 2725
rect 7913 2708 7947 2725
rect 7947 2708 7956 2725
rect 7904 2691 7913 2695
rect 7913 2691 7947 2695
rect 7947 2691 7956 2695
rect 7904 2652 7956 2691
rect 7904 2643 7913 2652
rect 7913 2643 7947 2652
rect 7947 2643 7956 2652
rect 7904 2618 7913 2630
rect 7913 2618 7947 2630
rect 7947 2618 7956 2630
rect 7904 2579 7956 2618
rect 7904 2578 7913 2579
rect 7913 2578 7947 2579
rect 7947 2578 7956 2579
rect 7904 2545 7913 2565
rect 7913 2545 7947 2565
rect 7947 2545 7956 2565
rect 7904 2513 7956 2545
rect 7904 2472 7913 2500
rect 7913 2472 7947 2500
rect 7947 2472 7956 2500
rect 7904 2448 7956 2472
rect 7904 2433 7956 2435
rect 7904 2399 7913 2433
rect 7913 2399 7947 2433
rect 7947 2399 7956 2433
rect 7904 2383 7956 2399
rect 7904 2360 7956 2370
rect 7904 2326 7913 2360
rect 7913 2326 7947 2360
rect 7947 2326 7956 2360
rect 7904 2318 7956 2326
rect 7904 2287 7956 2305
rect 7904 2253 7913 2287
rect 7913 2253 7947 2287
rect 7947 2253 7956 2287
rect 7904 2214 7956 2240
rect 7904 2188 7913 2214
rect 7913 2188 7947 2214
rect 7947 2188 7956 2214
rect 7904 2141 7956 2175
rect 7904 2123 7913 2141
rect 7913 2123 7947 2141
rect 7947 2123 7956 2141
rect 7904 2107 7913 2110
rect 7913 2107 7947 2110
rect 7947 2107 7956 2110
rect 7904 2068 7956 2107
rect 7904 2058 7913 2068
rect 7913 2058 7947 2068
rect 7947 2058 7956 2068
rect 7904 2034 7913 2045
rect 7913 2034 7947 2045
rect 7947 2034 7956 2045
rect 7904 1995 7956 2034
rect 7904 1993 7913 1995
rect 7913 1993 7947 1995
rect 7947 1993 7956 1995
rect 7904 1961 7913 1980
rect 7913 1961 7947 1980
rect 7947 1961 7956 1980
rect 7904 1928 7956 1961
rect 7904 1888 7913 1915
rect 7913 1888 7947 1915
rect 7947 1888 7956 1915
rect 7904 1863 7956 1888
rect 7904 1849 7956 1850
rect 7904 1815 7913 1849
rect 7913 1815 7947 1849
rect 7947 1815 7956 1849
rect 7904 1798 7956 1815
rect 7904 1776 7956 1785
rect 7904 1742 7913 1776
rect 7913 1742 7947 1776
rect 7947 1742 7956 1776
rect 7904 1733 7956 1742
rect 7904 1703 7956 1720
rect 7904 1669 7913 1703
rect 7913 1669 7947 1703
rect 7947 1669 7956 1703
rect 7904 1668 7956 1669
rect 7904 1630 7956 1655
rect 7904 1603 7913 1630
rect 7913 1603 7947 1630
rect 7947 1603 7956 1630
rect 7904 1557 7956 1590
rect 7904 1538 7913 1557
rect 7913 1538 7947 1557
rect 7947 1538 7956 1557
rect 7904 1523 7913 1525
rect 7913 1523 7947 1525
rect 7947 1523 7956 1525
rect 7904 1484 7956 1523
rect 7904 1473 7913 1484
rect 7913 1473 7947 1484
rect 7947 1473 7956 1484
rect 7904 1450 7913 1460
rect 7913 1450 7947 1460
rect 7947 1450 7956 1460
rect 7904 1411 7956 1450
rect 7904 1408 7913 1411
rect 7913 1408 7947 1411
rect 7947 1408 7956 1411
rect 7904 1377 7913 1395
rect 7913 1377 7947 1395
rect 7947 1377 7956 1395
rect 7904 1343 7956 1377
rect 7904 1304 7913 1330
rect 7913 1304 7947 1330
rect 7947 1304 7956 1330
rect 7904 1278 7956 1304
rect 7904 1231 7913 1265
rect 7913 1231 7947 1265
rect 7947 1231 7956 1265
rect 7904 1213 7956 1231
rect 7904 1192 7956 1200
rect 7904 1158 7913 1192
rect 7913 1158 7947 1192
rect 7947 1158 7956 1192
rect 7904 1148 7956 1158
rect 7904 1119 7956 1135
rect 7904 1085 7913 1119
rect 7913 1085 7947 1119
rect 7947 1085 7956 1119
rect 7904 1083 7956 1085
rect 7904 1046 7956 1070
rect 7904 1018 7913 1046
rect 7913 1018 7947 1046
rect 7947 1018 7956 1046
rect 7904 973 7956 1005
rect 7904 953 7913 973
rect 7913 953 7947 973
rect 7947 953 7956 973
rect 7904 939 7913 941
rect 7913 939 7947 941
rect 7947 939 7956 941
rect 7904 900 7956 939
rect 7904 889 7913 900
rect 7913 889 7947 900
rect 7947 889 7956 900
rect 7904 866 7913 877
rect 7913 866 7947 877
rect 7947 866 7956 877
rect 7904 827 7956 866
rect 7904 825 7913 827
rect 7913 825 7947 827
rect 7947 825 7956 827
rect 8225 2771 8277 2823
rect 8289 2771 8341 2823
rect 8353 2771 8405 2823
rect 8225 2705 8277 2757
rect 8289 2705 8341 2757
rect 8353 2705 8405 2757
rect 12145 2426 12197 2454
rect 12145 2402 12148 2426
rect 12148 2402 12188 2426
rect 12188 2402 12197 2426
rect 12090 2392 12114 2400
rect 12114 2392 12142 2400
rect 12283 2392 12296 2411
rect 12296 2392 12335 2411
rect 12090 2354 12142 2392
rect 12283 2359 12335 2392
rect 12228 2354 12280 2357
rect 12090 2348 12114 2354
rect 12114 2348 12142 2354
rect 12035 2320 12040 2346
rect 12040 2320 12074 2346
rect 12074 2320 12087 2346
rect 12228 2320 12262 2354
rect 12262 2320 12280 2354
rect 12035 2294 12087 2320
rect 12228 2305 12280 2320
rect 11980 2282 12032 2292
rect 12173 2282 12225 2303
rect 11980 2248 12000 2282
rect 12000 2248 12032 2282
rect 12173 2251 12188 2282
rect 12188 2251 12222 2282
rect 12222 2251 12225 2282
rect 12118 2248 12148 2249
rect 12148 2248 12170 2249
rect 11980 2240 12032 2248
rect 11925 2210 11977 2238
rect 12118 2210 12170 2248
rect 11925 2186 11926 2210
rect 11926 2186 11966 2210
rect 11966 2186 11977 2210
rect 11870 2176 11892 2184
rect 11892 2176 11922 2184
rect 12118 2197 12148 2210
rect 12148 2197 12170 2210
rect 12063 2176 12074 2195
rect 12074 2176 12114 2195
rect 12114 2176 12115 2195
rect 11870 2138 11922 2176
rect 12063 2143 12115 2176
rect 12008 2138 12060 2141
rect 11870 2132 11892 2138
rect 11892 2132 11922 2138
rect 11815 2104 11818 2130
rect 11818 2104 11852 2130
rect 11852 2104 11867 2130
rect 12008 2104 12040 2138
rect 12040 2104 12060 2138
rect 11815 2078 11867 2104
rect 12008 2089 12060 2104
rect 11760 2066 11812 2076
rect 11953 2066 12005 2087
rect 11760 2032 11778 2066
rect 11778 2032 11812 2066
rect 11953 2035 11966 2066
rect 11966 2035 12000 2066
rect 12000 2035 12005 2066
rect 11898 2032 11926 2033
rect 11926 2032 11950 2033
rect 11760 2024 11812 2032
rect 11705 1994 11757 2022
rect 11898 1994 11950 2032
rect 11705 1970 11744 1994
rect 11744 1970 11757 1994
rect 11898 1981 11926 1994
rect 11926 1981 11950 1994
rect 11843 1960 11852 1979
rect 11852 1960 11892 1979
rect 11892 1960 11895 1979
rect 11843 1927 11895 1960
rect 7904 793 7913 813
rect 7913 793 7947 813
rect 7947 793 7956 813
rect 7904 761 7956 793
rect 8992 755 9044 761
rect 9056 755 9108 761
rect 9121 755 9173 761
rect 9186 755 9238 761
rect 7904 721 7919 749
rect 7919 721 7953 749
rect 7953 721 7956 749
rect 8992 721 9014 755
rect 9014 721 9044 755
rect 9056 721 9087 755
rect 9087 721 9108 755
rect 9121 721 9160 755
rect 9160 721 9173 755
rect 9186 721 9194 755
rect 9194 721 9233 755
rect 9233 721 9238 755
rect 7904 697 7956 721
rect 8992 709 9044 721
rect 9056 709 9108 721
rect 9121 709 9173 721
rect 9186 709 9238 721
rect 7904 683 7956 685
rect 7904 649 7913 683
rect 7913 649 7947 683
rect 7947 649 7956 683
rect 7904 633 7956 649
rect 7904 601 7956 621
rect 7904 569 7913 601
rect 7913 569 7947 601
rect 7947 569 7956 601
rect 7904 519 7956 557
rect 7904 505 7913 519
rect 7913 505 7947 519
rect 7947 505 7956 519
rect 7904 485 7913 493
rect 7913 485 7947 493
rect 7947 485 7956 493
rect 7904 441 7956 485
rect 7904 402 7913 429
rect 7913 402 7947 429
rect 7947 402 7956 429
rect 7904 377 7956 402
rect 7904 353 7956 365
rect 7904 319 7913 353
rect 7913 319 7947 353
rect 7947 319 7956 353
rect 8992 347 9044 359
rect 7904 313 7956 319
rect 8992 313 9007 347
rect 9007 313 9041 347
rect 9041 313 9044 347
rect 8992 307 9044 313
rect 9056 347 9108 359
rect 9121 347 9173 359
rect 9186 347 9238 359
rect 9056 313 9081 347
rect 9081 313 9108 347
rect 9121 313 9155 347
rect 9155 313 9173 347
rect 9186 313 9189 347
rect 9189 313 9229 347
rect 9229 313 9238 347
rect 9056 307 9108 313
rect 9121 307 9173 313
rect 9186 307 9238 313
<< metal2 >>
rect -132 3108 -80 6473
rect -40 3108 12 6473
rect 1370 6106 1696 6473
tri 2474 6421 2526 6473 se
rect 2526 6421 3100 6473
tri 2468 6415 2474 6421 se
rect 2474 6415 3100 6421
tri 2454 6401 2468 6415 se
rect 2468 6401 3100 6415
tri 2402 6349 2454 6401 se
rect 2454 6349 3100 6401
tri 2388 6335 2402 6349 se
rect 2402 6335 3100 6349
tri 2336 6283 2388 6335 se
rect 2388 6283 3100 6335
rect 1370 6054 1376 6106
rect 1428 6054 1458 6106
rect 1510 6054 1540 6106
rect 1592 6054 1622 6106
rect 1674 6054 1696 6106
rect 1370 3596 1696 6054
rect 1370 3544 1376 3596
rect 1428 3544 1441 3596
rect 1493 3544 1506 3596
rect 1558 3544 1572 3596
rect 1624 3544 1638 3596
rect 1690 3544 1696 3596
rect 1370 3532 1696 3544
rect 1370 3480 1376 3532
rect 1428 3480 1441 3532
rect 1493 3480 1506 3532
rect 1558 3480 1572 3532
rect 1624 3480 1638 3532
rect 1690 3480 1696 3532
rect 1370 3108 1696 3480
tri 2290 6237 2336 6283 se
rect 2336 6237 3100 6283
rect 2290 3108 3100 6237
rect 4314 6421 4320 6473
rect 4372 6421 4385 6473
rect 4437 6421 4450 6473
rect 4502 6421 4516 6473
rect 4568 6421 4574 6473
rect 4314 3408 4574 6421
rect 4314 3356 4320 3408
rect 4372 3356 4385 3408
rect 4437 3356 4450 3408
rect 4502 3356 4516 3408
rect 4568 3356 4574 3408
rect 4314 3344 4574 3356
rect 4314 3292 4320 3344
rect 4372 3292 4385 3344
rect 4437 3292 4450 3344
rect 4502 3292 4516 3344
rect 4568 3292 4574 3344
rect 4314 3280 4574 3292
rect 4314 3228 4320 3280
rect 4372 3228 4385 3280
rect 4437 3228 4450 3280
rect 4502 3228 4516 3280
rect 4568 3228 4574 3280
rect 4757 6100 5017 6473
rect 4809 6048 4821 6100
rect 4873 6048 4885 6100
rect 4937 6048 5017 6100
rect 4757 6035 5017 6048
rect 4809 5983 4821 6035
rect 4873 5983 4885 6035
rect 4937 5983 5017 6035
rect 4757 5970 5017 5983
rect 4809 5918 4821 5970
rect 4873 5918 4885 5970
rect 4937 5918 5017 5970
rect 4757 5905 5017 5918
rect 4809 5853 4821 5905
rect 4873 5853 4885 5905
rect 4937 5853 5017 5905
rect 4757 5840 5017 5853
rect 4809 5788 4821 5840
rect 4873 5788 4885 5840
rect 4937 5788 5017 5840
rect 4757 5775 5017 5788
rect 4809 5723 4821 5775
rect 4873 5723 4885 5775
rect 4937 5723 5017 5775
rect 4757 5710 5017 5723
rect 4809 5658 4821 5710
rect 4873 5658 4885 5710
rect 4937 5658 5017 5710
rect 4757 5645 5017 5658
rect 4809 5593 4821 5645
rect 4873 5593 4885 5645
rect 4937 5593 5017 5645
rect 4757 5580 5017 5593
rect 4809 5528 4821 5580
rect 4873 5528 4885 5580
rect 4937 5528 5017 5580
rect 4757 5515 5017 5528
rect 4809 5463 4821 5515
rect 4873 5463 4885 5515
rect 4937 5463 5017 5515
rect 4757 5450 5017 5463
rect 4809 5398 4821 5450
rect 4873 5398 4885 5450
rect 4937 5398 5017 5450
rect 4757 5385 5017 5398
rect 4809 5333 4821 5385
rect 4873 5333 4885 5385
rect 4937 5333 5017 5385
rect 4757 5320 5017 5333
rect 4809 5268 4821 5320
rect 4873 5268 4885 5320
rect 4937 5268 5017 5320
rect 4757 5255 5017 5268
rect 4809 5203 4821 5255
rect 4873 5203 4885 5255
rect 4937 5203 5017 5255
rect 4757 5190 5017 5203
rect 4809 5138 4821 5190
rect 4873 5138 4885 5190
rect 4937 5138 5017 5190
rect 4757 5125 5017 5138
rect 4809 5073 4821 5125
rect 4873 5073 4885 5125
rect 4937 5073 5017 5125
rect 4757 5060 5017 5073
rect 4809 5008 4821 5060
rect 4873 5008 4885 5060
rect 4937 5008 5017 5060
rect 4757 4995 5017 5008
rect 4809 4943 4821 4995
rect 4873 4943 4885 4995
rect 4937 4943 5017 4995
rect 4757 4930 5017 4943
rect 4809 4878 4821 4930
rect 4873 4878 4885 4930
rect 4937 4878 5017 4930
rect 4757 4865 5017 4878
rect 4809 4813 4821 4865
rect 4873 4813 4885 4865
rect 4937 4813 5017 4865
rect 4757 4800 5017 4813
rect 4809 4748 4821 4800
rect 4873 4748 4885 4800
rect 4937 4748 5017 4800
rect 4757 4735 5017 4748
rect 4809 4683 4821 4735
rect 4873 4683 4885 4735
rect 4937 4683 5017 4735
rect 4757 4670 5017 4683
rect 4809 4618 4821 4670
rect 4873 4618 4885 4670
rect 4937 4618 5017 4670
rect 4757 4605 5017 4618
rect 4809 4553 4821 4605
rect 4873 4553 4885 4605
rect 4937 4553 5017 4605
rect 4757 4540 5017 4553
rect 4809 4488 4821 4540
rect 4873 4488 4885 4540
rect 4937 4488 5017 4540
rect 4757 4475 5017 4488
rect 4809 4423 4821 4475
rect 4873 4423 4885 4475
rect 4937 4423 5017 4475
rect 4757 4410 5017 4423
rect 4809 4358 4821 4410
rect 4873 4358 4885 4410
rect 4937 4358 5017 4410
rect 4757 4345 5017 4358
rect 4809 4293 4821 4345
rect 4873 4293 4885 4345
rect 4937 4293 5017 4345
rect 4757 4280 5017 4293
rect 4809 4228 4821 4280
rect 4873 4228 4885 4280
rect 4937 4228 5017 4280
rect 4757 4215 5017 4228
rect 4809 4163 4821 4215
rect 4873 4163 4885 4215
rect 4937 4163 5017 4215
rect 4757 4150 5017 4163
rect 4809 4098 4821 4150
rect 4873 4098 4885 4150
rect 4937 4098 5017 4150
rect 4757 4085 5017 4098
rect 4809 4033 4821 4085
rect 4873 4033 4885 4085
rect 4937 4033 5017 4085
rect 4757 4020 5017 4033
rect 4809 3968 4821 4020
rect 4873 3968 4885 4020
rect 4937 3968 5017 4020
rect 4757 3955 5017 3968
rect 4809 3903 4821 3955
rect 4873 3903 4885 3955
rect 4937 3903 5017 3955
rect 4757 3890 5017 3903
rect 4937 3454 5017 3890
rect 4757 3228 5017 3454
tri 4314 3208 4334 3228 ne
rect 4334 3208 4554 3228
tri 4554 3208 4574 3228 nw
tri 4334 3162 4380 3208 ne
rect 4380 3162 4508 3208
tri 4508 3162 4554 3208 nw
rect 5564 3108 5616 6473
rect 5656 3108 5708 6473
rect 6932 4208 6984 4214
rect 6932 4142 6984 4156
rect 6852 3904 6904 3910
rect 6852 3838 6904 3852
rect 6852 3260 6904 3786
rect 6932 3363 6984 4090
rect 7042 4208 7094 4214
rect 7042 4142 7094 4156
rect 7042 3443 7094 4090
rect 7161 4143 7291 6473
rect 7347 4872 7527 6473
rect 7399 4820 7411 4872
rect 7463 4820 7475 4872
rect 7347 4806 7527 4820
rect 7399 4754 7411 4806
rect 7463 4754 7475 4806
rect 7347 4748 7527 4754
rect 7583 6421 7589 6473
rect 7641 6421 7653 6473
rect 7705 6421 7717 6473
rect 7769 6421 7776 6473
rect 7583 6014 7776 6421
rect 7583 5962 7592 6014
rect 7644 5962 7656 6014
rect 7708 5962 7720 6014
rect 7772 5962 7776 6014
rect 7583 5949 7776 5962
rect 7583 5897 7592 5949
rect 7644 5897 7656 5949
rect 7708 5897 7720 5949
rect 7772 5897 7776 5949
rect 7583 5884 7776 5897
rect 7583 5832 7592 5884
rect 7644 5832 7656 5884
rect 7708 5832 7720 5884
rect 7772 5832 7776 5884
rect 7583 5819 7776 5832
rect 7583 5767 7592 5819
rect 7644 5767 7656 5819
rect 7708 5767 7720 5819
rect 7772 5767 7776 5819
rect 7583 5754 7776 5767
rect 7583 5702 7592 5754
rect 7644 5702 7656 5754
rect 7708 5702 7720 5754
rect 7772 5702 7776 5754
rect 7583 5689 7776 5702
rect 7583 5637 7592 5689
rect 7644 5637 7656 5689
rect 7708 5637 7720 5689
rect 7772 5637 7776 5689
rect 7583 5624 7776 5637
rect 7583 5572 7592 5624
rect 7644 5572 7656 5624
rect 7708 5572 7720 5624
rect 7772 5572 7776 5624
rect 7583 5558 7776 5572
rect 7583 5506 7592 5558
rect 7644 5506 7656 5558
rect 7708 5506 7720 5558
rect 7772 5506 7776 5558
rect 7583 5492 7776 5506
rect 7583 5440 7592 5492
rect 7644 5440 7656 5492
rect 7708 5440 7720 5492
rect 7772 5440 7776 5492
rect 7583 5426 7776 5440
rect 7583 5374 7592 5426
rect 7644 5374 7656 5426
rect 7708 5374 7720 5426
rect 7772 5374 7776 5426
rect 7583 5360 7776 5374
rect 7583 5308 7592 5360
rect 7644 5308 7656 5360
rect 7708 5308 7720 5360
rect 7772 5308 7776 5360
rect 7583 5294 7776 5308
rect 7583 5242 7592 5294
rect 7644 5242 7656 5294
rect 7708 5242 7720 5294
rect 7772 5242 7776 5294
rect 7583 5228 7776 5242
rect 7583 5176 7592 5228
rect 7644 5176 7656 5228
rect 7708 5176 7720 5228
rect 7772 5176 7776 5228
rect 7583 5162 7776 5176
rect 7583 5110 7592 5162
rect 7644 5110 7656 5162
rect 7708 5110 7720 5162
rect 7772 5110 7776 5162
rect 7583 5096 7776 5110
rect 7583 5044 7592 5096
rect 7644 5044 7656 5096
rect 7708 5044 7720 5096
rect 7772 5044 7776 5096
rect 7583 5030 7776 5044
rect 7583 4978 7592 5030
rect 7644 4978 7656 5030
rect 7708 4978 7720 5030
rect 7772 4978 7776 5030
rect 7583 4964 7776 4978
rect 7583 4912 7592 4964
rect 7644 4912 7656 4964
rect 7708 4912 7720 4964
rect 7772 4912 7776 4964
rect 7583 4640 7776 4912
rect 7583 4588 7592 4640
rect 7644 4588 7656 4640
rect 7708 4588 7720 4640
rect 7772 4588 7776 4640
rect 7583 4569 7776 4588
rect 7583 4517 7592 4569
rect 7644 4517 7656 4569
rect 7708 4517 7720 4569
rect 7772 4517 7776 4569
rect 7583 4498 7776 4517
rect 7583 4446 7592 4498
rect 7644 4446 7656 4498
rect 7708 4446 7720 4498
rect 7772 4446 7776 4498
rect 7583 4427 7776 4446
rect 7583 4375 7592 4427
rect 7644 4375 7656 4427
rect 7708 4375 7720 4427
rect 7772 4375 7776 4427
rect 7583 4356 7776 4375
rect 7583 4304 7592 4356
rect 7644 4304 7656 4356
rect 7708 4304 7720 4356
rect 7772 4304 7776 4356
rect 7583 4285 7776 4304
rect 7583 4233 7592 4285
rect 7644 4233 7656 4285
rect 7708 4233 7720 4285
rect 7772 4233 7776 4285
rect 7583 4214 7776 4233
rect 7583 4162 7592 4214
rect 7644 4162 7656 4214
rect 7708 4162 7720 4214
rect 7772 4162 7776 4214
tri 7291 4143 7307 4159 sw
rect 7161 4142 7307 4143
tri 7307 4142 7308 4143 sw
rect 7583 4142 7776 4162
rect 7161 4090 7308 4142
tri 7308 4090 7360 4142 sw
rect 7583 4090 7592 4142
rect 7644 4090 7656 4142
rect 7708 4090 7720 4142
rect 7772 4090 7776 4142
rect 7161 4084 7360 4090
tri 7360 4084 7366 4090 sw
rect 7161 4081 7366 4084
tri 7366 4081 7369 4084 sw
rect 7161 4056 7369 4081
tri 7369 4056 7394 4081 sw
rect 7161 4004 7167 4056
rect 7219 4004 7233 4056
rect 7285 4004 7299 4056
rect 7351 4004 7394 4056
rect 7161 3992 7394 4004
rect 7161 3940 7167 3992
rect 7219 3940 7233 3992
rect 7285 3940 7299 3992
rect 7351 3940 7394 3992
tri 7161 3936 7165 3940 ne
rect 7165 3936 7394 3940
tri 7165 3884 7217 3936 ne
rect 7217 3884 7394 3936
tri 7217 3883 7218 3884 ne
rect 7218 3883 7394 3884
tri 7218 3872 7229 3883 ne
rect 7229 3872 7394 3883
tri 7229 3837 7264 3872 ne
tri 7094 3443 7096 3445 sw
rect 7042 3420 7096 3443
tri 7096 3420 7119 3443 sw
rect 7042 3368 7048 3420
rect 7100 3368 7114 3420
rect 7166 3368 7172 3420
tri 6984 3363 6986 3365 sw
rect 6932 3340 6986 3363
tri 6986 3340 7009 3363 sw
rect 6932 3299 6949 3340
tri 6932 3288 6943 3299 ne
rect 6943 3288 6949 3299
rect 7001 3288 7015 3340
rect 7067 3288 7073 3340
tri 6904 3260 6929 3285 sw
rect 6852 3208 6858 3260
rect 6910 3208 6924 3260
rect 6976 3208 6982 3260
rect 7264 2969 7394 3872
rect 7583 3827 7776 4090
rect 7583 3775 7592 3827
rect 7644 3775 7656 3827
rect 7708 3775 7720 3827
rect 7772 3775 7776 3827
rect 7583 2969 7776 3775
rect 7904 6147 8169 6473
rect 8662 6175 8668 6227
rect 8720 6175 8732 6227
rect 8784 6175 8802 6227
rect 8830 6175 8836 6227
rect 8888 6175 8900 6227
rect 8952 6175 8958 6227
tri 8725 6153 8747 6175 ne
rect 8747 6153 8802 6175
tri 8881 6153 8903 6175 ne
rect 8903 6153 8958 6175
tri 8747 6150 8750 6153 ne
rect 7904 6095 7913 6147
rect 7965 6095 7979 6147
rect 8031 6095 8045 6147
rect 8097 6095 8111 6147
rect 8163 6095 8169 6147
rect 7904 6075 8169 6095
rect 7904 6023 7907 6075
rect 7959 6023 8169 6075
rect 7904 6010 8169 6023
rect 8592 6021 8598 6073
rect 8650 6021 8662 6073
rect 8714 6021 8720 6073
rect 7904 5958 7907 6010
rect 7959 5958 8169 6010
tri 8643 5996 8668 6021 ne
rect 7904 5945 8169 5958
rect 7904 5893 7907 5945
rect 7959 5893 8169 5945
rect 7904 5880 8169 5893
rect 7904 5828 7907 5880
rect 7959 5828 8169 5880
rect 7904 5815 8169 5828
rect 7904 5763 7907 5815
rect 7959 5763 8169 5815
rect 7904 5750 8169 5763
rect 7904 5698 7907 5750
rect 7959 5698 8169 5750
rect 7904 5685 8169 5698
rect 7904 5633 7907 5685
rect 7959 5633 8169 5685
rect 7904 5620 8169 5633
rect 7904 5568 7907 5620
rect 7959 5568 8169 5620
rect 7904 5555 8169 5568
rect 7904 5503 7907 5555
rect 7959 5503 8169 5555
rect 7904 5489 8169 5503
rect 7904 5437 7907 5489
rect 7959 5437 8169 5489
rect 7904 5423 8169 5437
rect 7904 5371 7907 5423
rect 7959 5371 8169 5423
rect 7904 5357 8169 5371
rect 7904 5305 7907 5357
rect 7959 5305 8169 5357
rect 8197 5941 8203 5993
rect 8255 5941 8269 5993
rect 8321 5941 8327 5993
rect 8197 5919 8246 5941
tri 8246 5919 8268 5941 nw
rect 8197 5681 8243 5919
tri 8243 5916 8246 5919 nw
rect 8429 5867 8460 5919
rect 8512 5867 8527 5919
rect 8579 5867 8585 5919
rect 8429 5839 8484 5867
tri 8484 5839 8512 5867 nw
rect 8271 5782 8277 5834
rect 8329 5782 8343 5834
rect 8395 5782 8401 5834
tri 8330 5759 8353 5782 ne
rect 8353 5759 8401 5782
tri 8353 5757 8355 5759 ne
tri 8243 5681 8268 5706 sw
rect 8197 5629 8203 5681
rect 8255 5629 8269 5681
rect 8321 5629 8327 5681
rect 8197 5398 8243 5629
tri 8243 5604 8268 5629 nw
tri 8329 5526 8355 5552 se
rect 8355 5526 8401 5759
rect 8271 5474 8277 5526
rect 8329 5474 8343 5526
rect 8395 5474 8401 5526
tri 8243 5398 8254 5409 sw
rect 8197 5372 8254 5398
tri 8254 5372 8280 5398 sw
rect 8197 5320 8203 5372
rect 8255 5320 8269 5372
rect 8321 5320 8327 5372
rect 7904 5291 8169 5305
rect 7904 5239 7907 5291
rect 7959 5239 8169 5291
rect 7904 5225 8169 5239
rect 7904 5173 7907 5225
rect 7959 5173 8169 5225
rect 8429 5259 8481 5839
tri 8481 5836 8484 5839 nw
rect 8512 5707 8518 5759
rect 8570 5707 8582 5759
rect 8634 5707 8640 5759
tri 8563 5682 8588 5707 ne
tri 8481 5259 8506 5284 sw
rect 8429 5207 8435 5259
rect 8487 5207 8502 5259
rect 8554 5207 8560 5259
rect 7904 5003 8169 5173
tri 8573 5013 8588 5028 se
rect 8588 5013 8640 5707
tri 8563 5003 8573 5013 se
rect 8573 5003 8640 5013
rect 7904 4951 7913 5003
rect 7965 4951 7979 5003
rect 8031 4951 8045 5003
rect 8097 4951 8111 5003
rect 8163 4951 8169 5003
rect 8509 4951 8515 5003
rect 8567 4951 8582 5003
rect 8634 4951 8640 5003
rect 7904 4651 8169 4951
tri 8563 4939 8575 4951 ne
rect 8575 4939 8640 4951
tri 8575 4936 8578 4939 ne
rect 8578 4936 8640 4939
tri 8578 4926 8588 4936 ne
rect 7904 4599 7913 4651
rect 7965 4599 7979 4651
rect 8031 4599 8045 4651
rect 8097 4599 8111 4651
rect 8163 4599 8169 4651
rect 7904 3936 8169 4599
rect 7904 3884 7913 3936
rect 7965 3884 7979 3936
rect 8031 3884 8045 3936
rect 8097 3884 8111 3936
rect 8163 3884 8169 3936
rect 7904 3523 8169 3884
rect 7904 3471 7913 3523
rect 7965 3471 7979 3523
rect 8031 3471 8045 3523
rect 8097 3471 8111 3523
rect 8163 3471 8169 3523
rect 7904 2825 8169 3471
rect 7956 2773 8169 2825
rect 7904 2760 8169 2773
rect 7956 2708 8169 2760
rect 7904 2695 8169 2708
rect 8225 4872 8405 4878
rect 8277 4820 8289 4872
rect 8341 4820 8353 4872
rect 8225 4806 8405 4820
rect 8277 4754 8289 4806
rect 8341 4754 8353 4806
rect 8225 2823 8405 4754
tri 8563 4395 8588 4420 se
rect 8588 4395 8640 4936
rect 8509 4343 8515 4395
rect 8567 4343 8582 4395
rect 8634 4343 8640 4395
rect 8668 5232 8720 6021
rect 8750 5681 8802 6153
tri 8903 6150 8906 6153 ne
tri 8881 5993 8906 6018 se
rect 8906 5993 8958 6153
rect 8830 5941 8836 5993
rect 8888 5941 8900 5993
rect 8952 5941 8958 5993
tri 8881 5916 8906 5941 ne
tri 8802 5681 8827 5706 sw
rect 8750 5629 8756 5681
rect 8808 5629 8820 5681
rect 8872 5629 8878 5681
tri 8801 5604 8826 5629 ne
tri 8720 5232 8732 5244 sw
rect 8668 5221 8732 5232
tri 8732 5221 8743 5232 sw
rect 8668 5219 8743 5221
tri 8743 5219 8745 5221 sw
rect 8668 5167 8674 5219
rect 8726 5167 8740 5219
rect 8792 5167 8798 5219
rect 8668 5159 8737 5167
tri 8737 5159 8745 5167 nw
rect 8502 3964 8508 4016
rect 8560 3964 8574 4016
rect 8626 3964 8632 4016
tri 8555 3960 8559 3964 ne
rect 8559 3960 8632 3964
tri 8559 3939 8580 3960 ne
rect 8580 3662 8632 3960
rect 8668 3698 8720 5159
tri 8720 5142 8737 5159 nw
tri 8801 5112 8826 5137 se
rect 8826 5112 8878 5629
rect 8748 5060 8754 5112
rect 8806 5060 8820 5112
rect 8872 5060 8878 5112
rect 8748 4705 8754 4757
rect 8806 4705 8820 4757
rect 8872 4705 8878 4757
rect 8748 4702 8822 4705
tri 8822 4702 8825 4705 nw
rect 8748 4699 8819 4702
tri 8819 4699 8822 4702 nw
rect 8748 4684 8804 4699
tri 8804 4684 8819 4699 nw
rect 8748 4159 8800 4684
tri 8800 4680 8804 4684 nw
tri 8886 4583 8906 4603 se
rect 8906 4583 8958 5941
tri 8881 4578 8886 4583 se
rect 8886 4578 8958 4583
rect 8828 4526 8834 4578
rect 8886 4526 8900 4578
rect 8952 4526 8958 4578
rect 8986 6153 9244 6473
rect 9680 6467 9873 6473
rect 9680 6415 9693 6467
rect 9745 6415 9757 6467
rect 9809 6415 9821 6467
rect 9680 6401 9873 6415
rect 9680 6349 9693 6401
rect 9745 6349 9757 6401
rect 9809 6349 9821 6401
rect 9680 6335 9873 6349
rect 9680 6283 9693 6335
rect 9745 6283 9757 6335
rect 9809 6283 9821 6335
rect 8986 6101 8992 6153
rect 9044 6101 9056 6153
rect 9108 6101 9121 6153
rect 9173 6101 9186 6153
rect 9238 6101 9244 6153
rect 8986 5398 9244 6101
rect 9431 6175 9437 6227
rect 9489 6175 9503 6227
rect 9555 6175 9561 6227
rect 8986 5346 8992 5398
rect 9044 5346 9056 5398
rect 9108 5346 9121 5398
rect 9173 5346 9186 5398
rect 9238 5346 9244 5398
rect 8986 4936 9244 5346
rect 8986 4884 8992 4936
rect 9044 4884 9056 4936
rect 9108 4884 9121 4936
rect 9173 4884 9186 4936
rect 9238 4884 9244 4936
rect 8986 4672 9244 4884
rect 8986 4620 8992 4672
rect 9044 4620 9056 4672
rect 9108 4620 9121 4672
rect 9173 4620 9186 4672
rect 9238 4620 9244 4672
tri 8800 4159 8802 4161 sw
rect 8748 4143 8802 4159
tri 8802 4143 8818 4159 sw
rect 8748 4142 8818 4143
tri 8818 4142 8819 4143 sw
rect 8748 4136 8819 4142
tri 8819 4136 8825 4142 sw
rect 8986 4136 9244 4620
rect 8748 4084 8754 4136
rect 8806 4084 8820 4136
rect 8872 4084 8878 4136
rect 8986 4084 8992 4136
rect 9044 4084 9056 4136
rect 9108 4084 9121 4136
rect 9173 4084 9186 4136
rect 9238 4084 9244 4136
rect 8748 4081 8822 4084
tri 8822 4081 8825 4084 nw
rect 8748 3787 8800 4081
tri 8800 4059 8822 4081 nw
tri 8800 3787 8822 3809 sw
rect 8748 3784 8822 3787
tri 8822 3784 8825 3787 sw
rect 8748 3732 8754 3784
rect 8806 3732 8820 3784
rect 8872 3732 8878 3784
tri 8720 3698 8726 3704 sw
rect 8668 3682 8726 3698
tri 8668 3667 8683 3682 ne
rect 8683 3667 8726 3682
tri 8632 3662 8637 3667 sw
tri 8683 3662 8688 3667 ne
rect 8688 3662 8726 3667
rect 8580 3657 8637 3662
tri 8637 3657 8642 3662 sw
tri 8688 3657 8693 3662 ne
rect 8693 3657 8726 3662
tri 8726 3657 8767 3698 sw
rect 8580 3645 8642 3657
tri 8580 3608 8617 3645 ne
rect 8617 3639 8642 3645
tri 8642 3639 8660 3657 sw
tri 8693 3639 8711 3657 ne
rect 8711 3639 8767 3657
rect 8617 3608 8660 3639
tri 8660 3608 8691 3639 sw
tri 8711 3624 8726 3639 ne
rect 8726 3624 8767 3639
tri 8767 3624 8800 3657 sw
tri 8726 3608 8742 3624 ne
rect 8742 3608 8800 3624
tri 8617 3588 8637 3608 ne
rect 8637 3588 8691 3608
tri 8691 3588 8711 3608 sw
tri 8742 3602 8748 3608 ne
tri 8637 3566 8659 3588 ne
rect 8277 2771 8289 2823
rect 8341 2771 8353 2823
rect 8225 2757 8405 2771
rect 8277 2705 8289 2757
rect 8341 2705 8353 2757
rect 8225 2699 8405 2705
rect 8501 3311 8507 3363
rect 8559 3311 8571 3363
rect 8623 3311 8629 3363
rect 7956 2643 8169 2695
rect 8501 2671 8553 3311
tri 8553 3286 8578 3311 nw
tri 8637 2973 8659 2995 se
rect 8659 2973 8711 3588
tri 8585 2921 8637 2973 se
rect 8637 2921 8711 2973
tri 8581 2917 8585 2921 se
rect 8585 2917 8711 2921
rect 8581 2865 8587 2917
rect 8639 2865 8653 2917
rect 8705 2865 8711 2917
rect 7904 2630 8169 2643
rect 7956 2578 8169 2630
rect 7904 2565 8169 2578
rect 7956 2513 8169 2565
rect 7904 2500 8169 2513
rect 7956 2448 8169 2500
rect 7904 2435 8169 2448
rect 7956 2383 8169 2435
rect 7904 2370 8169 2383
rect 7956 2318 8169 2370
rect 7904 2305 8169 2318
rect 7956 2253 8169 2305
rect 7904 2240 8169 2253
rect 7956 2188 8169 2240
rect 7904 2175 8169 2188
rect 7956 2123 8169 2175
rect 7904 2110 8169 2123
rect 7956 2058 8169 2110
rect 7904 2045 8169 2058
rect 7956 1993 8169 2045
rect 7904 1980 8169 1993
rect 7956 1928 8169 1980
rect 7904 1915 8169 1928
rect 7956 1863 8169 1915
rect 7904 1850 8169 1863
rect 7956 1798 8169 1850
rect 7904 1785 8169 1798
rect 7956 1733 8169 1785
rect 7904 1720 8169 1733
rect 7956 1668 8169 1720
rect 7904 1655 8169 1668
rect 7956 1603 8169 1655
rect 7904 1590 8169 1603
rect 7956 1538 8169 1590
rect 7904 1525 8169 1538
rect 7956 1473 8169 1525
rect 7904 1460 8169 1473
rect 7956 1408 8169 1460
rect 7904 1395 8169 1408
rect 7956 1343 8169 1395
rect 7904 1330 8169 1343
rect 7956 1278 8169 1330
rect 7904 1265 8169 1278
rect 7956 1213 8169 1265
rect 7904 1200 8169 1213
rect 7956 1148 8169 1200
rect 7904 1135 8169 1148
rect 7956 1083 8169 1135
rect 7904 1070 8169 1083
rect 7956 1018 8169 1070
rect 7904 1005 8169 1018
rect 7956 953 8169 1005
rect 7904 941 8169 953
rect 7956 889 8169 941
rect 7904 877 8169 889
rect 7956 825 8169 877
rect 7904 813 8169 825
rect 7956 761 8169 813
tri 8169 761 8170 762 sw
rect 7904 749 8170 761
rect 7956 697 8170 749
rect 7904 685 8170 697
rect 7956 633 8170 685
rect 7904 621 8170 633
rect 7956 569 8170 621
rect 7904 557 8170 569
rect 7956 505 8170 557
rect 7904 493 8170 505
rect 7956 441 8170 493
rect 7904 429 8170 441
rect 7956 377 8170 429
rect 7904 365 8170 377
rect 7956 313 8170 365
rect 7904 307 8170 313
rect 8748 -53 8800 3608
rect 8986 761 9244 4084
rect 9272 5438 9278 5490
rect 9330 5438 9344 5490
rect 9396 5438 9402 5490
rect 9272 5232 9318 5438
tri 9318 5413 9343 5438 nw
tri 9318 5232 9332 5246 sw
rect 9272 5221 9332 5232
tri 9332 5221 9343 5232 sw
rect 9272 5169 9278 5221
rect 9330 5169 9344 5221
rect 9396 5169 9402 5221
rect 9272 5159 9333 5169
tri 9333 5159 9343 5169 nw
rect 9272 3883 9318 5159
tri 9318 5144 9333 5159 nw
tri 9406 4754 9431 4779 se
rect 9431 4754 9485 6175
tri 9485 6150 9510 6175 nw
rect 9680 6080 9873 6283
rect 9680 5964 9757 6080
rect 9355 4702 9361 4754
rect 9413 4702 9427 4754
rect 9479 4702 9485 4754
tri 9406 4699 9409 4702 ne
rect 9409 4699 9485 4702
tri 9409 4684 9424 4699 ne
rect 9424 4684 9485 4699
tri 9424 4677 9431 4684 ne
tri 9403 4422 9431 4450 se
rect 9431 4422 9485 4684
rect 9355 4370 9361 4422
rect 9413 4370 9427 4422
rect 9479 4370 9485 4422
rect 9522 5600 9528 5652
rect 9580 5600 9594 5652
rect 9646 5600 9652 5652
rect 9522 5572 9624 5600
tri 9624 5572 9652 5600 nw
rect 9355 4260 9361 4312
rect 9413 4260 9427 4312
rect 9479 4260 9485 4312
tri 9406 4258 9408 4260 ne
rect 9408 4258 9485 4260
tri 9408 4244 9422 4258 ne
rect 9422 4244 9485 4258
tri 9422 4235 9431 4244 ne
tri 9406 3960 9431 3985 se
rect 9431 3960 9485 4244
rect 9353 3908 9359 3960
rect 9411 3908 9425 3960
rect 9477 3908 9485 3960
tri 9406 3897 9417 3908 ne
rect 9417 3897 9485 3908
tri 9318 3883 9332 3897 sw
tri 9417 3883 9431 3897 ne
rect 9272 3872 9332 3883
tri 9332 3872 9343 3883 sw
rect 9272 3820 9278 3872
rect 9330 3820 9344 3872
rect 9396 3820 9402 3872
tri 9406 3608 9431 3633 se
rect 9431 3608 9485 3897
rect 9355 3556 9361 3608
rect 9413 3556 9427 3608
rect 9479 3556 9485 3608
rect 9522 4310 9574 5572
tri 9574 5522 9624 5572 nw
rect 9522 4244 9574 4258
tri 9497 3443 9522 3468 se
rect 9522 3443 9574 4192
rect 9444 3391 9450 3443
rect 9502 3391 9516 3443
rect 9568 3391 9574 3443
rect 9680 5232 9873 5964
rect 9680 5180 9693 5232
rect 9745 5180 9757 5232
rect 9809 5180 9821 5232
rect 9680 5159 9873 5180
rect 9680 5107 9693 5159
rect 9745 5107 9757 5159
rect 9809 5107 9821 5159
rect 9680 5086 9873 5107
rect 9680 5034 9693 5086
rect 9745 5034 9757 5086
rect 9809 5034 9821 5086
rect 9680 5013 9873 5034
rect 9680 4961 9693 5013
rect 9745 4961 9757 5013
rect 9809 4961 9821 5013
rect 9680 4939 9873 4961
rect 9680 4887 9693 4939
rect 9745 4887 9757 4939
rect 9809 4887 9821 4939
rect 9680 4751 9873 4887
rect 9680 4699 9693 4751
rect 9745 4699 9757 4751
rect 9809 4699 9821 4751
rect 9680 4667 9873 4699
rect 9680 4615 9693 4667
rect 9745 4615 9757 4667
rect 9809 4615 9821 4667
rect 9680 4583 9873 4615
rect 9680 4531 9693 4583
rect 9745 4531 9757 4583
rect 9809 4531 9821 4583
rect 9680 4417 9873 4531
rect 9680 4365 9693 4417
rect 9745 4365 9757 4417
rect 9809 4365 9821 4417
rect 9680 4349 9873 4365
rect 9680 4297 9693 4349
rect 9745 4297 9757 4349
rect 9809 4297 9821 4349
rect 9680 4280 9873 4297
rect 9680 4228 9693 4280
rect 9745 4228 9757 4280
rect 9809 4228 9821 4280
rect 9680 4211 9873 4228
rect 9680 4159 9693 4211
rect 9745 4159 9757 4211
rect 9809 4159 9821 4211
rect 9680 4142 9873 4159
rect 9680 4090 9693 4142
rect 9745 4090 9757 4142
rect 9809 4090 9821 4142
rect 9680 3949 9873 4090
rect 9732 3897 9744 3949
rect 9796 3897 9808 3949
rect 9860 3897 9873 3949
rect 9680 3883 9873 3897
rect 9732 3831 9744 3883
rect 9796 3831 9808 3883
rect 9860 3831 9873 3883
rect 9680 3443 9873 3831
rect 9680 3391 9686 3443
rect 9738 3391 9750 3443
rect 9802 3391 9815 3443
rect 9867 3391 9873 3443
rect 9412 2997 9418 3049
rect 9470 2997 9482 3049
rect 9534 2997 9540 3049
rect 9412 2973 9465 2997
tri 9465 2973 9489 2997 nw
rect 9412 2671 9464 2973
tri 9464 2972 9465 2973 nw
rect 9680 2969 9873 3391
rect 10220 6231 10226 6283
rect 10278 6231 10290 6283
rect 10342 6231 10348 6283
rect 10220 4575 10272 6231
tri 10272 6155 10348 6231 nw
rect 10962 6231 10968 6283
rect 11020 6231 11032 6283
rect 11084 6231 11090 6283
rect 10380 5787 10386 5839
rect 10438 5787 10450 5839
rect 10502 5787 10508 5839
rect 10220 4509 10272 4523
rect 8986 709 8992 761
rect 9044 709 9056 761
rect 9108 709 9121 761
rect 9173 709 9186 761
rect 9238 709 9244 761
rect 8986 359 9244 709
rect 8986 307 8992 359
rect 9044 307 9056 359
rect 9108 307 9121 359
rect 9173 307 9186 359
rect 9238 307 9244 359
rect 10220 -53 10272 4457
rect 10300 5375 10352 5381
rect 10300 5310 10352 5323
rect 10300 4261 10352 5258
rect 10380 4934 10432 5787
tri 10432 5754 10465 5787 nw
rect 10460 5520 10466 5572
rect 10518 5520 10530 5572
rect 10582 5520 10588 5572
tri 10515 5487 10548 5520 ne
rect 10380 4868 10432 4882
rect 10380 4736 10432 4816
rect 10380 4670 10432 4684
rect 10380 4612 10432 4618
rect 10300 4195 10352 4209
rect 10300 4137 10352 4143
rect 10548 4081 10588 5520
tri 10588 4081 10621 4114 sw
rect 10548 4029 10554 4081
rect 10606 4029 10618 4081
rect 10670 4029 10676 4081
rect 10548 3735 10588 4029
tri 10588 3996 10621 4029 nw
rect 10962 3787 11002 6231
tri 11002 6206 11027 6231 nw
rect 11578 5752 11584 5804
rect 11636 5752 11648 5804
rect 11700 5752 11706 5804
tri 11002 3787 11027 3812 sw
tri 10588 3735 10595 3742 sw
rect 10962 3735 10968 3787
rect 11020 3735 11032 3787
rect 11084 3735 11090 3787
rect 10548 3723 10595 3735
tri 10595 3723 10607 3735 sw
rect 10548 3709 10607 3723
tri 10607 3709 10621 3723 sw
rect 10548 3657 10554 3709
rect 10606 3657 10618 3709
rect 10670 3657 10676 3709
rect 10548 3611 10588 3657
tri 10588 3624 10621 3657 nw
tri 11553 3363 11578 3388 se
rect 11578 3363 11630 5752
tri 11630 5727 11655 5752 nw
rect 11502 3311 11508 3363
rect 11560 3311 11572 3363
rect 11624 3311 11630 3363
rect 11686 4748 11692 4800
rect 11744 4748 11756 4800
rect 11808 4748 11814 4800
tri 11661 3049 11686 3074 se
rect 11686 3049 11738 4748
tri 11738 4723 11763 4748 nw
rect 11794 3671 11800 3723
rect 11852 3671 11866 3723
rect 11918 3671 11924 3723
rect 11794 3659 11924 3671
rect 11794 3607 11800 3659
rect 11852 3607 11866 3659
rect 11918 3607 11924 3659
rect 11794 3367 11924 3607
rect 11980 3499 11986 3551
rect 12038 3499 12052 3551
rect 12104 3499 12110 3551
rect 11980 3487 12110 3499
rect 11980 3435 11986 3487
rect 12038 3435 12052 3487
rect 12104 3435 12110 3487
rect 11980 3367 12110 3435
rect 12166 3367 12388 6473
rect 13106 6288 13158 6473
tri 13158 6288 13183 6313 sw
rect 13106 6236 13112 6288
rect 13164 6236 13180 6288
rect 13232 6236 13238 6288
tri 13081 3831 13106 3856 se
rect 13106 3831 13158 6236
tri 13158 6211 13183 6236 nw
rect 12444 3779 12450 3831
rect 12502 3779 12516 3831
rect 12568 3779 12574 3831
rect 13028 3779 13034 3831
rect 13086 3779 13100 3831
rect 13152 3779 13158 3831
rect 10324 2997 10330 3049
rect 10382 2997 10394 3049
rect 10446 2997 10452 3049
rect 11610 2997 11616 3049
rect 11668 2997 11680 3049
rect 11732 2997 11738 3049
rect 10324 2973 10377 2997
tri 10377 2973 10401 2997 nw
rect 10324 2671 10376 2973
tri 10376 2972 10377 2973 nw
rect 12139 2402 12145 2454
rect 12197 2402 12203 2454
rect 12084 2348 12090 2400
rect 12142 2348 12148 2400
rect 12277 2359 12283 2411
rect 12335 2359 12341 2411
rect 12029 2294 12035 2346
rect 12087 2294 12093 2346
rect 12222 2305 12228 2357
rect 12280 2305 12286 2357
rect 11974 2240 11980 2292
rect 12032 2240 12038 2292
rect 12167 2251 12173 2303
rect 12225 2251 12231 2303
rect 11919 2186 11925 2238
rect 11977 2186 11983 2238
rect 12112 2197 12118 2249
rect 12170 2197 12176 2249
rect 11864 2132 11870 2184
rect 11922 2132 11928 2184
rect 12057 2143 12063 2195
rect 12115 2143 12121 2195
rect 11809 2078 11815 2130
rect 11867 2078 11873 2130
rect 12002 2089 12008 2141
rect 12060 2089 12066 2141
rect 11754 2024 11760 2076
rect 11812 2024 11818 2076
rect 11947 2035 11953 2087
rect 12005 2035 12011 2087
rect 11699 1970 11705 2022
rect 11757 1970 11763 2022
rect 11892 1981 11898 2033
rect 11950 1981 11956 2033
rect 11837 1927 11843 1979
rect 11895 1927 11901 1979
rect 12444 1279 12496 3779
tri 12496 3753 12522 3779 nw
rect 13613 2973 13757 6473
rect 13837 3723 13965 6473
rect 13837 3607 13843 3723
rect 13959 3607 13965 3723
rect 14023 3551 14151 6473
rect 14023 3435 14029 3551
rect 14145 3435 14151 3551
tri 13757 2973 14151 3367 sw
rect 13613 2921 13619 2973
rect 13671 2921 13685 2973
rect 13737 2921 13751 2973
rect 13803 2921 13817 2973
rect 13869 2921 13883 2973
rect 13935 2921 13949 2973
rect 14001 2921 14015 2973
rect 14067 2921 14151 2973
rect 13613 2909 14151 2921
rect 13613 2857 13619 2909
rect 13671 2857 13685 2909
rect 13737 2857 13751 2909
rect 13803 2857 13817 2909
rect 13869 2857 13883 2909
rect 13935 2857 13949 2909
rect 14001 2857 14015 2909
rect 14067 2857 14151 2909
rect 13613 1279 14151 2857
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 1 12624 1 0 3077
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform -1 0 8883 0 1 5873
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform -1 0 13206 0 1 6246
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform -1 0 8895 0 1 3480
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform -1 0 8303 0 1 3009
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform -1 0 8821 0 -1 4748
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform -1 0 8703 0 -1 4127
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1704896540
transform -1 0 8706 0 -1 5210
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1704896540
transform -1 0 12686 0 -1 6277
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1704896540
transform -1 0 8775 0 -1 3924
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1704896540
transform -1 0 8691 0 -1 4921
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1704896540
transform 0 -1 12150 1 0 5612
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1704896540
transform 0 -1 11798 1 0 5612
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1704896540
transform 0 -1 12412 1 0 5686
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1704896540
transform 0 -1 12326 1 0 5686
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1704896540
transform 0 -1 11974 1 0 5686
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1704896540
transform 0 -1 11622 1 0 5686
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1704896540
transform 0 -1 8708 1 0 4379
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1704896540
transform 1 0 10707 0 -1 6277
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1704896540
transform 1 0 11979 0 -1 6277
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1704896540
transform 1 0 11290 0 1 6158
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1704896540
transform 1 0 8681 0 1 5450
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1704896540
transform 1 0 12381 0 1 5444
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1704896540
transform 0 1 9764 -1 0 6088
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_1
timestamp 1704896540
transform -1 0 13003 0 -1 6277
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_2
timestamp 1704896540
transform 0 1 10614 1 0 5692
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_3
timestamp 1704896540
transform 0 -1 11512 1 0 5714
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_4
timestamp 1704896540
transform 1 0 11046 0 1 6232
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 11256 1 0 5918
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 10904 1 0 5918
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform 0 -1 13259 -1 0 6055
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_1
timestamp 1704896540
transform 0 -1 12747 -1 0 6055
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1704896540
transform 1 0 12780 0 1 3243
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1704896540
transform 1 0 12780 0 1 3071
box -12 -6 550 40
use L1M1_CDNS_52468879185285  L1M1_CDNS_52468879185285_0
timestamp 1704896540
transform 0 -1 9896 -1 0 6395
box -12 -6 118 328
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1704896540
transform 1 0 12780 0 1 3157
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1704896540
transform 1 0 6780 0 -1 3820
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform -1 0 11814 0 1 4748
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform -1 0 10588 0 1 5520
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform -1 0 10676 0 1 4029
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform -1 0 8720 0 -1 6073
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform 1 0 10380 0 -1 5839
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform 1 0 8662 0 -1 6227
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform 1 0 8750 0 -1 5681
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform 1 0 8512 0 -1 5759
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1704896540
transform 1 0 10220 0 -1 6283
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1704896540
transform 1 0 8830 0 -1 6227
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1704896540
transform 1 0 8830 0 -1 5993
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1704896540
transform 1 0 11578 0 1 5752
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1704896540
transform 1 0 11502 0 1 3311
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1704896540
transform 1 0 10548 0 1 3657
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1704896540
transform 1 0 8501 0 1 3311
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1704896540
transform 1 0 10962 0 1 6231
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1704896540
transform 1 0 10962 0 1 3735
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1704896540
transform 1 0 11610 0 1 2997
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1704896540
transform 1 0 9412 0 1 2997
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1704896540
transform 1 0 10324 0 1 2997
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1704896540
transform 1 0 12192 0 1 2466
box 0 0 192 244
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1704896540
transform 1 0 11699 0 1 1970
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_1
timestamp 1704896540
transform 1 0 11754 0 1 2024
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_2
timestamp 1704896540
transform 1 0 11809 0 1 2078
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_3
timestamp 1704896540
transform 1 0 11864 0 1 2132
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_4
timestamp 1704896540
transform 1 0 11919 0 1 2186
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_5
timestamp 1704896540
transform 1 0 11974 0 1 2240
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_6
timestamp 1704896540
transform 1 0 12029 0 1 2294
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_7
timestamp 1704896540
transform 1 0 12084 0 1 2348
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_8
timestamp 1704896540
transform 1 0 12139 0 1 2402
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_9
timestamp 1704896540
transform 1 0 12277 0 1 2359
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_10
timestamp 1704896540
transform 1 0 12222 0 1 2305
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_11
timestamp 1704896540
transform 1 0 12167 0 1 2251
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_12
timestamp 1704896540
transform 1 0 12112 0 1 2197
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_13
timestamp 1704896540
transform 1 0 12057 0 1 2143
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_14
timestamp 1704896540
transform 1 0 12002 0 1 2089
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_15
timestamp 1704896540
transform 1 0 11947 0 1 2035
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_16
timestamp 1704896540
transform 1 0 11837 0 1 1927
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_17
timestamp 1704896540
transform 1 0 11892 0 1 1981
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1704896540
transform 1 0 11617 0 -1 1917
box 0 0 192 180
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_0
timestamp 1704896540
transform 0 1 8501 -1 0 2671
box 0 0 512 52
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_1
timestamp 1704896540
transform 0 1 10324 -1 0 2671
box 0 0 512 52
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_2
timestamp 1704896540
transform 0 1 9412 -1 0 2671
box 0 0 512 52
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1704896540
transform 0 1 8859 -1 0 4879
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_1
timestamp 1704896540
transform 0 1 8859 -1 0 5341
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_2
timestamp 1704896540
transform 0 1 8859 -1 0 4703
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_3
timestamp 1704896540
transform 0 1 8021 -1 0 4231
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_4
timestamp 1704896540
transform 0 1 8021 -1 0 3879
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_5
timestamp 1704896540
transform 0 1 8859 1 0 4935
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_6
timestamp 1704896540
transform 0 1 8021 1 0 3935
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_7
timestamp 1704896540
transform 0 1 8859 1 0 5397
box -79 -26 199 626
use nfet_CDNS_52468879185319  nfet_CDNS_52468879185319_0
timestamp 1704896540
transform 0 1 8859 -1 0 4261
box -79 -26 375 626
use nfet_CDNS_52468879185319  nfet_CDNS_52468879185319_1
timestamp 1704896540
transform 0 1 8859 -1 0 3909
box -79 -26 375 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_0
timestamp 1704896540
transform 0 1 8859 -1 0 4527
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_1
timestamp 1704896540
transform 0 -1 9459 1 0 5683
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_2
timestamp 1704896540
transform 0 -1 9459 1 0 5839
box -79 -26 179 626
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_0
timestamp 1704896540
transform 0 1 8021 1 0 4653
box -79 -26 375 626
use nfet_CDNS_52468879185392  nfet_CDNS_52468879185392_0
timestamp 1704896540
transform 0 -1 8621 1 0 5371
box -79 -26 647 626
use nfet_CDNS_524688791851173  nfet_CDNS_524688791851173_0
timestamp 1704896540
transform 0 1 8021 -1 0 4597
box -79 -26 279 626
use nfet_CDNS_524688791851173  nfet_CDNS_524688791851173_1
timestamp 1704896540
transform 0 1 8021 1 0 5005
box -79 -26 279 626
use nfet_CDNS_524688791851651  nfet_CDNS_524688791851651_0
timestamp 1704896540
transform -1 0 4708 0 1 3777
box -79 -26 1735 2026
use nfet_CDNS_524688791851651  nfet_CDNS_524688791851651_1
timestamp 1704896540
transform -1 0 2140 0 1 3777
box -79 -26 1735 2026
use nfet_CDNS_524688791851652  nfet_CDNS_524688791851652_0
timestamp 1704896540
transform -1 0 2996 0 1 3777
box -79 -26 879 2026
use nfet_CDNS_524688791851653  nfet_CDNS_524688791851653_0
timestamp 1704896540
transform 0 1 8021 -1 0 3593
box -79 -26 479 226
use nfet_CDNS_524688791851654  nfet_CDNS_524688791851654_0
timestamp 1704896540
transform -1 0 8954 0 1 829
box -79 -26 935 2026
use nfet_CDNS_524688791851655  nfet_CDNS_524688791851655_0
timestamp 1704896540
transform 1 0 9010 0 1 829
box -79 -26 1847 2026
use nfet_CDNS_524688791851656  nfet_CDNS_524688791851656_0
timestamp 1704896540
transform -1 0 7276 0 -1 5890
box -79 -26 259 2026
use nfet_CDNS_524688791851656  nfet_CDNS_524688791851656_1
timestamp 1704896540
transform -1 0 6930 0 -1 5890
box -79 -26 259 2026
use nfet_CDNS_524688791851657  nfet_CDNS_524688791851657_0
timestamp 1704896540
transform 0 1 8459 -1 0 3293
box -79 -26 179 1026
use pfet_CDNS_52468879185134  pfet_CDNS_52468879185134_0
timestamp 1704896540
transform -1 0 12137 0 1 4829
box -119 -66 239 666
use pfet_CDNS_52468879185134  pfet_CDNS_52468879185134_1
timestamp 1704896540
transform -1 0 12313 0 1 4829
box -119 -66 239 666
use pfet_CDNS_52468879185134  pfet_CDNS_52468879185134_2
timestamp 1704896540
transform -1 0 12702 0 -1 6195
box -119 -66 239 666
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_0
timestamp 1704896540
transform -1 0 11467 0 -1 6195
box -119 -66 319 666
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_1
timestamp 1704896540
transform -1 0 10859 0 -1 6195
box -119 -66 319 666
use pfet_CDNS_524688791851658  pfet_CDNS_524688791851658_0
timestamp 1704896540
transform 0 -1 13306 -1 0 3232
box -89 -36 205 636
use pfet_CDNS_524688791851659  pfet_CDNS_524688791851659_0
timestamp 1704896540
transform -1 0 13369 0 1 4829
box -119 -66 767 666
use pfet_CDNS_524688791851660  pfet_CDNS_524688791851660_0
timestamp 1704896540
transform -1 0 11851 0 1 4829
box -119 -66 1311 666
use pfet_CDNS_524688791851661  pfet_CDNS_524688791851661_0
timestamp 1704896540
transform -1 0 12665 0 1 4829
box -119 -66 415 666
use pfet_CDNS_524688791851661  pfet_CDNS_524688791851661_1
timestamp 1704896540
transform -1 0 11211 0 -1 6195
box -119 -66 415 666
use pfet_CDNS_524688791851662  pfet_CDNS_524688791851662_0
timestamp 1704896540
transform 1 0 12758 0 -1 6195
box -119 -66 575 666
use pfet_CDNS_524688791851663  pfet_CDNS_524688791851663_0
timestamp 1704896540
transform -1 0 12281 0 -1 6195
box -119 -66 767 666
use pfet_CDNS_524688791851664  pfet_CDNS_524688791851664_0
timestamp 1704896540
transform 1 0 10659 0 -1 4719
box -119 -66 2559 666
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform -1 0 8319 0 -1 3593
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform -1 0 8827 0 -1 4527
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform -1 0 8827 0 -1 5531
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1704896540
transform -1 0 8427 0 -1 3359
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1704896540
transform 0 -1 13214 1 0 6227
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1704896540
transform 0 -1 12702 1 0 6227
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1704896540
transform 0 -1 12320 1 0 5461
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1704896540
transform 0 -1 12137 1 0 5461
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1704896540
transform 1 0 8653 0 -1 4949
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1704896540
transform 1 0 8653 0 -1 5205
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1704896540
transform 1 0 12608 0 1 3116
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_11
timestamp 1704896540
transform 1 0 8653 0 1 3745
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1704896540
transform -1 0 8827 0 1 3613
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1704896540
transform 0 1 12369 1 0 5461
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1704896540
transform 1 0 8653 0 1 4395
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1704896540
transform 0 1 10659 1 0 6227
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1704896540
transform -1 0 8827 0 1 3991
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1704896540
transform -1 0 8827 0 -1 5953
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_2
timestamp 1704896540
transform 1 0 8653 0 1 3958
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1704896540
transform 0 1 2219 -1 0 3745
box 0 0 66 746
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1704896540
transform 1 0 8653 0 -1 5939
box 0 0 66 542
use PYL1_CDNS_52468879185370  PYL1_CDNS_52468879185370_0
timestamp 1704896540
transform -1 0 8827 0 -1 5341
box 0 0 66 678
use PYL1_CDNS_52468879185370  PYL1_CDNS_52468879185370_1
timestamp 1704896540
transform 0 1 11267 1 0 6227
box 0 0 66 678
use PYL1_CDNS_52468879185370  PYL1_CDNS_52468879185370_2
timestamp 1704896540
transform 0 -1 13399 1 0 5461
box 0 0 66 678
use PYL1_CDNS_524688791851203  PYL1_CDNS_524688791851203_0
timestamp 1704896540
transform 0 1 6776 -1 0 3836
box 0 0 66 474
use PYL1_CDNS_524688791851646  PYL1_CDNS_524688791851646_0
timestamp 1704896540
transform 0 -1 2114 1 0 5809
box 0 0 66 1630
use PYL1_CDNS_524688791851647  PYL1_CDNS_524688791851647_0
timestamp 1704896540
transform 0 -1 10778 1 0 2861
box 0 0 66 2718
use PYL1_CDNS_524688791851648  PYL1_CDNS_524688791851648_0
timestamp 1704896540
transform 0 1 10658 -1 0 4087
box 0 0 66 2446
use PYL1_CDNS_524688791851649  PYL1_CDNS_524688791851649_0
timestamp 1704896540
transform 0 1 10629 -1 0 5527
box 0 0 66 1222
use sky130_fd_io__sio_pudrvr_reg_csw_res  sky130_fd_io__sio_pudrvr_reg_csw_res_0
timestamp 1704896540
transform 1 0 4997 0 -1 6012
box -26 0 1530 2317
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1704896540
transform -1 0 8810 0 1 5787
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1704896540
transform 1 0 10156 0 -1 5318
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_5246887918565  sky130_fd_io__tk_em1s_CDNS_5246887918565_0
timestamp 1704896540
transform -1 0 10771 0 1 4137
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_5246887918565  sky130_fd_io__tk_em1s_CDNS_5246887918565_1
timestamp 1704896540
transform -1 0 10764 0 1 5252
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_5246887918565  sky130_fd_io__tk_em1s_CDNS_5246887918565_2
timestamp 1704896540
transform 1 0 10471 0 1 4587
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_5246887918565  sky130_fd_io__tk_em1s_CDNS_5246887918565_3
timestamp 1704896540
transform 1 0 10471 0 1 4831
box 0 0 1 1
<< labels >>
flabel locali 8671 5155 8671 5155 0 FreeSans 300 90 0 0 slow_h_n
flabel locali 8670 4078 8670 4078 0 FreeSans 300 90 0 0 drvhi_h_n_s
flabel locali 8782 3752 8782 3752 0 FreeSans 300 270 0 0 drvhi_h
flabel locali s 8806 5123 8806 5123 0 FreeSans 300 270 0 0 drvhi_h_n_s
flabel locali 12036 5517 12036 5517 0 FreeSans 300 0 0 0 drvhi_h_n_s
flabel comment s 2674 6149 2674 6149 0 FreeSans 1000 0 0 0 condiode
flabel comment s 5784 6151 5784 6151 0 FreeSans 1000 0 0 0 condiode
flabel comment s 8810 6148 8810 6148 0 FreeSans 1000 0 0 0 condiode
flabel comment s 12270 6459 12270 6459 3 FreeSans 200 270 0 0 vnb
flabel comment s 4743 4503 4743 4503 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 3892 4503 3892 4503 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 3036 4503 3036 4503 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 2182 4503 2182 4503 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 7561 4412 7561 4412 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 3603 6106 3603 6106 0 FreeSans 300 180 0 0 vgnd_io
flabel comment s 7862 6106 7862 6106 0 FreeSans 300 180 0 0 vgnd_io
flabel comment s 9466 5815 9466 5815 0 FreeSans 300 180 0 0 vref_nng
flabel comment s 9401 5894 9401 5894 0 FreeSans 300 180 0 0 ncap_s3
flabel comment s 9446 4736 9446 4736 0 FreeSans 300 0 0 0 ncap_s2
flabel comment s 9445 4915 9445 4915 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 9406 5699 9406 5699 0 FreeSans 300 0 0 0 ncap_s1
flabel comment s 9463 5096 9463 5096 0 FreeSans 300 180 0 0 ncap_s1
flabel comment s 9460 4117 9460 4117 0 FreeSans 300 180 0 0 vgnd_io
flabel comment s 9440 3938 9440 3938 0 FreeSans 300 180 0 0 int_2
flabel comment s 9454 5360 9454 5360 0 FreeSans 300 180 0 0 vgnd_io
flabel comment s 9452 4594 9452 4594 0 FreeSans 300 0 0 0 ncap_s3
flabel comment s 9478 4376 9478 4376 0 FreeSans 300 180 0 0 ncap_s2
flabel comment s 7030 3773 7030 3773 0 FreeSans 300 0 0 0 m1_vpwr
flabel comment s 8049 4041 8049 4041 0 FreeSans 300 180 0 0 int_4
flabel comment s 8036 3941 8036 3941 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 8051 4219 8051 4219 0 FreeSans 300 180 0 0 nng_sd
flabel comment s 8060 4662 8060 4662 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 8067 5010 8067 5010 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 8047 4814 8047 4814 0 FreeSans 300 180 0 0 vref_nng
flabel comment s 8044 4392 8044 4392 0 FreeSans 300 180 0 0 puen_reg_h_n
flabel comment s 9431 5545 9431 5545 0 FreeSans 300 180 0 0 hvpsw_s
flabel comment s 9389 5208 9389 5208 0 FreeSans 300 180 0 0 hvnsw_s
flabel comment s 8646 3667 8646 3667 0 FreeSans 300 180 0 0 hvpsw_s
flabel comment s 10329 2985 10329 2985 0 FreeSans 300 270 0 0 lvpsw_s
flabel comment s 8713 3818 8713 3818 0 FreeSans 300 270 0 0 hvnsw_s
flabel comment s 8776 4098 8776 4098 0 FreeSans 300 90 0 0 puen_reg_h
flabel comment s 7866 5907 7866 5907 0 FreeSans 300 0 0 0 m2_ncap_s3
flabel comment s 8772 5829 8772 5829 0 FreeSans 300 270 0 0 slow_h
flabel comment s 11074 5841 11074 5841 0 FreeSans 300 270 0 0 drvhi_h_n_s
flabel comment s 12900 6120 12900 6120 0 FreeSans 300 0 0 0 drvhi_h_n_s
flabel comment s 12643 6296 12643 6296 0 FreeSans 300 0 0 0 drvhi_h_n_s
flabel comment s 13230 5737 13230 5737 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 11466 5861 11466 5861 0 FreeSans 300 0 0 0 slow_h
flabel comment s 10608 5836 10608 5836 0 FreeSans 300 270 0 0 puen_reg_h_n
flabel comment s 12955 6292 12955 6292 0 FreeSans 300 0 0 0 drvhi_h
flabel comment s 12571 5842 12571 5842 0 FreeSans 300 90 0 0 hvnsw_s
flabel comment s 12682 5361 12682 5361 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 12325 5212 12325 5212 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 12165 5219 12165 5219 0 FreeSans 300 90 0 0 int_1
flabel comment s 11989 5214 11989 5214 0 FreeSans 300 90 0 0 int_3
flabel comment s 11915 5783 11915 5783 0 FreeSans 300 0 0 0 int_5
flabel comment s 13026 5341 13026 5341 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 13400 5481 13400 5481 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 13202 5369 13202 5369 0 FreeSans 300 90 0 0 nng_sd
flabel comment s 12849 5365 12849 5365 0 FreeSans 300 90 0 0 nng_sd
flabel comment s 12491 5343 12491 5343 0 FreeSans 300 270 0 0 hvpsw_s
flabel comment s 7983 5228 7983 5228 0 FreeSans 300 180 0 0 slow_h
flabel comment s 9440 3586 9440 3586 0 FreeSans 300 180 0 0 int_2
flabel comment s 9440 4286 9440 4286 0 FreeSans 300 180 0 0 int_2
flabel comment s 9083 3786 9083 3786 0 FreeSans 300 0 0 0 li_drvhi_h_n_s
flabel comment s 11855 3486 11855 3486 0 FreeSans 300 270 0 0 voutref
flabel comment s 12044 3486 12044 3486 0 FreeSans 300 270 0 0 refleak_bias
flabel comment s 14092 6311 14092 6311 0 FreeSans 300 270 0 0 refleak_bias
flabel comment s 6728 3868 6728 3868 0 FreeSans 300 0 0 0 vrefin
flabel comment s 13903 6311 13903 6311 0 FreeSans 300 270 0 0 voutref
flabel comment s 10178 6197 10178 6197 0 FreeSans 300 180 0 0 int_3
flabel comment s 1638 4847 1638 4847 0 FreeSans 300 0 0 0 vref_nng
flabel comment s 4101 4847 4101 4847 0 FreeSans 300 0 0 0 vref_nng
flabel comment s 6740 4003 6740 4003 0 FreeSans 300 0 0 0 m1_vrefin
flabel comment s 4098 4094 4098 4094 0 FreeSans 300 0 0 0 vrefin
flabel comment s 1723 4508 1723 4508 0 FreeSans 300 90 0 0 m2_int_3
flabel comment s 1635 4094 1635 4094 0 FreeSans 300 0 0 0 vrefin
flabel comment s 1324 4503 1324 4503 0 FreeSans 300 270 0 0 vgnd_io
flabel comment s 3751 5861 3751 5861 0 FreeSans 300 0 0 0 ncap_s1
flabel comment s 1176 5873 1176 5873 0 FreeSans 300 0 0 0 ncap_s2
flabel comment s 2724 5877 2724 5877 0 FreeSans 300 0 0 0 ncap_s3
flabel comment s 5036 5892 5036 5892 0 FreeSans 300 0 0 0 int_5
flabel comment s 13675 3257 13675 3257 0 FreeSans 300 270 0 0 vpwr_ka
flabel comment s 10227 6451 10227 6451 0 FreeSans 300 180 0 0 lvpsw_s
flabel comment s -107 6386 -107 6386 3 FreeSans 200 270 0 0 pu_h_n<0>
flabel comment s 13076 3186 13076 3186 0 FreeSans 300 90 0 0 psh_int_1
flabel comment s 6500 5910 6500 5910 0 FreeSans 300 0 0 0 nng_sd
flabel comment s 1599 5558 1599 5558 0 FreeSans 300 0 0 0 m1_vpwr
flabel comment s 4068 5558 4068 5558 0 FreeSans 300 0 0 0 m1_vpwr
flabel comment s 4852 5987 4852 5987 0 FreeSans 300 0 0 0 ncap_s2
flabel comment s 7471 5901 7471 5901 0 FreeSans 300 0 0 0 m1_ncap_s1
flabel comment s 8719 5661 8719 5661 0 FreeSans 300 90 0 0 hvnsw_s
flabel comment s 8715 4822 8715 4822 0 FreeSans 300 270 0 0 puen_reg_h_n
flabel comment s 8714 4494 8714 4494 0 FreeSans 300 270 0 0 puen_reg_h
flabel comment s 10230 5474 10230 5474 0 FreeSans 300 0 0 0 hvnsw_s
flabel comment s 8766 4462 8766 4462 0 FreeSans 300 90 0 0 ncap_s3
flabel comment s 3191 5907 3191 5907 0 FreeSans 300 0 0 0 m1_ncap_s3
flabel comment s -16 6386 -16 6386 3 FreeSans 200 270 0 0 pu_h_n<1>
flabel comment s 11191 4747 11191 4747 0 FreeSans 300 180 0 0 hvpsw_s
flabel comment s 10216 5110 10216 5110 0 FreeSans 300 180 0 0 vpwr
flabel comment s 10557 3526 10557 3526 0 FreeSans 300 90 0 0 hvpsw_s
flabel comment s 10221 5540 10221 5540 0 FreeSans 300 180 0 0 hvpsw_s
flabel comment s -107 3143 -107 3143 3 FreeSans 200 90 0 0 pu_h_n<0>
flabel comment s -16 3143 -16 3143 3 FreeSans 200 90 0 0 pu_h_n<1>
flabel comment s 3595 6058 3595 6058 0 FreeSans 300 0 0 0 int_5
flabel comment s 12899 6351 12899 6351 0 FreeSans 300 0 0 0 nng_sd
flabel comment s 12038 6302 12038 6302 0 FreeSans 300 0 0 0 slow_h_n
flabel comment s 5588 3136 5588 3136 3 FreeSans 200 90 0 0 od_h
flabel comment s 12429 5463 12429 5463 0 FreeSans 300 0 0 0 hvnsw_s
flabel comment s 5678 3136 5678 3136 3 FreeSans 200 90 0 0 oe_hs_h
flabel comment s 12720 5737 12720 5737 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 5588 6417 5588 6417 3 FreeSans 200 270 0 0 od_h
flabel comment s 5678 6417 5678 6417 3 FreeSans 200 270 0 0 oe_hs_h
flabel comment s 10948 6293 10948 6293 0 FreeSans 300 180 0 0 puen_reg_h
flabel comment s 7862 6188 7862 6188 0 FreeSans 300 180 0 0 int_3
flabel comment s 10638 6184 10638 6184 0 FreeSans 300 180 0 0 int_3
flabel comment s 11073 5598 11073 5598 0 FreeSans 300 0 0 0 vcc_io
flabel comment s 2694 6352 2694 6352 0 FreeSans 300 180 0 0 nng_sd
flabel comment s 790 5265 790 5265 0 FreeSans 300 270 0 0 m2_nng_sd
flabel comment s 13674 6417 13674 6417 3 FreeSans 200 270 0 0 vpwr_ka
flabel comment s 13674 3400 13674 3400 3 FreeSans 200 90 0 0 vpwr_ka
flabel comment s 7856 6370 7856 6370 0 FreeSans 300 0 0 0 nng_sd
flabel comment s 9421 5480 9421 5480 0 FreeSans 300 180 0 0 hvnsw_s
flabel comment s 11042 4062 11042 4062 0 FreeSans 300 180 0 0 hvpsw_s
flabel comment s 10179 5893 10179 5893 0 FreeSans 300 0 0 0 slow_h
flabel comment s 8583 4494 8583 4494 0 FreeSans 300 270 0 0 nng_sd
flabel comment s 2567 6417 2567 6417 3 FreeSans 200 270 0 0 vgnd_io
flabel comment s 2567 3115 2567 3115 3 FreeSans 200 90 0 0 vgnd_io
flabel comment s 10233 5630 10233 5630 0 FreeSans 300 0 0 0 puen_reg_h_n
flabel comment s 8501 4519 8501 4519 0 FreeSans 300 90 0 0 ncap_s2
flabel comment s 9375 4021 9375 4021 0 FreeSans 300 270 0 0 hvnsw_s
flabel comment s 9071 3892 9071 3892 0 FreeSans 300 0 0 0 m1_hvnsw_s
flabel comment s 8630 3573 8630 3573 0 FreeSans 300 0 0 0 hvnsw_s
flabel comment s 10051 5803 10051 5803 0 FreeSans 300 180 0 0 vref_nng
flabel comment s 10313 4342 10313 4342 0 FreeSans 300 90 0 0 vrefin
flabel comment s 10323 4735 10323 4735 0 FreeSans 300 90 0 0 vrefin
flabel comment s 10415 4742 10415 4742 0 FreeSans 300 270 0 0 vref_nng
flabel comment s 11769 5791 11769 5791 0 FreeSans 300 270 0 0 nng_sd
flabel comment s 12298 6046 12298 6046 0 FreeSans 300 0 0 0 int_5
flabel comment s 11603 6046 11603 6046 0 FreeSans 300 0 0 0 int_5
flabel comment s 12105 5791 12105 5791 0 FreeSans 300 270 0 0 nng_sd
flabel comment s 10084 5294 10084 5294 0 FreeSans 300 180 0 0 vrefin
flabel metal1 s 10078 3471 10239 3523 0 FreeSans 200 0 0 0 drvhi_h
port 2 nsew
flabel metal1 s 10057 6152 10132 6198 0 FreeSans 200 0 0 0 slow_h_n
port 3 nsew
flabel metal1 s 10072 4785 10192 4853 0 FreeSans 200 0 0 0 vref_nng
port 5 nsew
flabel metal1 s 10091 4451 10220 4497 0 FreeSans 200 0 0 0 puen_reg_h
port 4 nsew
flabel metal1 s 10186 4137 10300 4267 0 FreeSans 200 0 0 0 vrefin
port 6 nsew
flabel metal2 s 4757 3228 5017 3277 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 4757 6427 5017 6473 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 1370 6427 1696 6473 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 1370 3108 1696 3164 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 9680 6427 9873 6473 0 FreeSans 200 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 7583 6421 7776 6473 0 FreeSans 200 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 7904 6427 8169 6473 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 8986 6427 9244 6473 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 7264 2969 7394 3049 0 FreeSans 200 0 0 0 vrefin
port 6 nsew
flabel metal2 s 7161 6427 7291 6473 0 FreeSans 200 0 0 0 vrefin
port 6 nsew
flabel metal2 s 7347 6427 7527 6473 0 FreeSans 200 0 0 0 vref_nng
port 5 nsew
flabel metal2 s 13106 6434 13158 6473 0 FreeSans 200 0 0 0 drvhi_h
port 2 nsew
flabel metal2 s 10220 -53 10272 -5 0 FreeSans 200 0 0 0 puen_reg_h
port 4 nsew
flabel metal2 s 8748 -53 8800 -6 0 FreeSans 200 0 0 0 slow_h_n
port 3 nsew
flabel metal2 s 8986 307 9244 373 0 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal2 s 7583 2969 7776 3049 0 FreeSans 200 0 0 0 vcc_io
port 8 nsew
flabel metal2 s 9680 2969 9873 3049 0 FreeSans 200 0 0 0 vcc_io
port 8 nsew
<< properties >>
string GDS_END 97990350
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97530348
string path 244.575 122.025 244.575 130.950 
<< end >>
