magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 10 143 2258 2195
<< mvnnmos >>
rect 271 169 1071 2169
rect 1197 169 1997 2169
<< mvndiff >>
rect 176 2119 271 2169
rect 176 2085 191 2119
rect 225 2085 271 2119
rect 176 2051 271 2085
rect 176 2017 191 2051
rect 225 2017 271 2051
rect 176 1983 271 2017
rect 176 1949 191 1983
rect 225 1949 271 1983
rect 176 1915 271 1949
rect 176 1881 191 1915
rect 225 1881 271 1915
rect 176 1847 271 1881
rect 176 1813 191 1847
rect 225 1813 271 1847
rect 176 1779 271 1813
rect 176 1745 191 1779
rect 225 1745 271 1779
rect 176 1711 271 1745
rect 176 1677 191 1711
rect 225 1677 271 1711
rect 176 1643 271 1677
rect 176 1609 191 1643
rect 225 1609 271 1643
rect 176 1575 271 1609
rect 176 1541 191 1575
rect 225 1541 271 1575
rect 176 1507 271 1541
rect 176 1473 191 1507
rect 225 1473 271 1507
rect 176 1439 271 1473
rect 176 1405 191 1439
rect 225 1405 271 1439
rect 176 1371 271 1405
rect 176 1337 191 1371
rect 225 1337 271 1371
rect 176 1303 271 1337
rect 176 1269 191 1303
rect 225 1269 271 1303
rect 176 1235 271 1269
rect 176 1201 191 1235
rect 225 1201 271 1235
rect 176 1167 271 1201
rect 176 1133 191 1167
rect 225 1133 271 1167
rect 176 1099 271 1133
rect 176 1065 191 1099
rect 225 1065 271 1099
rect 176 1031 271 1065
rect 176 997 191 1031
rect 225 997 271 1031
rect 176 963 271 997
rect 176 929 191 963
rect 225 929 271 963
rect 176 895 271 929
rect 176 861 191 895
rect 225 861 271 895
rect 176 827 271 861
rect 176 793 191 827
rect 225 793 271 827
rect 176 759 271 793
rect 176 725 191 759
rect 225 725 271 759
rect 176 691 271 725
rect 176 657 191 691
rect 225 657 271 691
rect 176 623 271 657
rect 176 589 191 623
rect 225 589 271 623
rect 176 555 271 589
rect 176 521 191 555
rect 225 521 271 555
rect 176 487 271 521
rect 176 453 191 487
rect 225 453 271 487
rect 176 419 271 453
rect 176 385 191 419
rect 225 385 271 419
rect 176 351 271 385
rect 176 317 191 351
rect 225 317 271 351
rect 176 283 271 317
rect 176 249 191 283
rect 225 249 271 283
rect 176 215 271 249
rect 176 181 191 215
rect 225 181 271 215
rect 176 169 271 181
rect 1071 2119 1197 2169
rect 1071 2085 1117 2119
rect 1151 2085 1197 2119
rect 1071 2051 1197 2085
rect 1071 2017 1117 2051
rect 1151 2017 1197 2051
rect 1071 1983 1197 2017
rect 1071 1949 1117 1983
rect 1151 1949 1197 1983
rect 1071 1915 1197 1949
rect 1071 1881 1117 1915
rect 1151 1881 1197 1915
rect 1071 1847 1197 1881
rect 1071 1813 1117 1847
rect 1151 1813 1197 1847
rect 1071 1779 1197 1813
rect 1071 1745 1117 1779
rect 1151 1745 1197 1779
rect 1071 1711 1197 1745
rect 1071 1677 1117 1711
rect 1151 1677 1197 1711
rect 1071 1643 1197 1677
rect 1071 1609 1117 1643
rect 1151 1609 1197 1643
rect 1071 1575 1197 1609
rect 1071 1541 1117 1575
rect 1151 1541 1197 1575
rect 1071 1507 1197 1541
rect 1071 1473 1117 1507
rect 1151 1473 1197 1507
rect 1071 1439 1197 1473
rect 1071 1405 1117 1439
rect 1151 1405 1197 1439
rect 1071 1371 1197 1405
rect 1071 1337 1117 1371
rect 1151 1337 1197 1371
rect 1071 1303 1197 1337
rect 1071 1269 1117 1303
rect 1151 1269 1197 1303
rect 1071 1235 1197 1269
rect 1071 1201 1117 1235
rect 1151 1201 1197 1235
rect 1071 1167 1197 1201
rect 1071 1133 1117 1167
rect 1151 1133 1197 1167
rect 1071 1099 1197 1133
rect 1071 1065 1117 1099
rect 1151 1065 1197 1099
rect 1071 1031 1197 1065
rect 1071 997 1117 1031
rect 1151 997 1197 1031
rect 1071 963 1197 997
rect 1071 929 1117 963
rect 1151 929 1197 963
rect 1071 895 1197 929
rect 1071 861 1117 895
rect 1151 861 1197 895
rect 1071 827 1197 861
rect 1071 793 1117 827
rect 1151 793 1197 827
rect 1071 759 1197 793
rect 1071 725 1117 759
rect 1151 725 1197 759
rect 1071 691 1197 725
rect 1071 657 1117 691
rect 1151 657 1197 691
rect 1071 623 1197 657
rect 1071 589 1117 623
rect 1151 589 1197 623
rect 1071 555 1197 589
rect 1071 521 1117 555
rect 1151 521 1197 555
rect 1071 487 1197 521
rect 1071 453 1117 487
rect 1151 453 1197 487
rect 1071 419 1197 453
rect 1071 385 1117 419
rect 1151 385 1197 419
rect 1071 351 1197 385
rect 1071 317 1117 351
rect 1151 317 1197 351
rect 1071 283 1197 317
rect 1071 249 1117 283
rect 1151 249 1197 283
rect 1071 215 1197 249
rect 1071 181 1117 215
rect 1151 181 1197 215
rect 1071 169 1197 181
rect 1997 2119 2092 2169
rect 1997 2085 2043 2119
rect 2077 2085 2092 2119
rect 1997 2051 2092 2085
rect 1997 2017 2043 2051
rect 2077 2017 2092 2051
rect 1997 1983 2092 2017
rect 1997 1949 2043 1983
rect 2077 1949 2092 1983
rect 1997 1915 2092 1949
rect 1997 1881 2043 1915
rect 2077 1881 2092 1915
rect 1997 1847 2092 1881
rect 1997 1813 2043 1847
rect 2077 1813 2092 1847
rect 1997 1779 2092 1813
rect 1997 1745 2043 1779
rect 2077 1745 2092 1779
rect 1997 1711 2092 1745
rect 1997 1677 2043 1711
rect 2077 1677 2092 1711
rect 1997 1643 2092 1677
rect 1997 1609 2043 1643
rect 2077 1609 2092 1643
rect 1997 1575 2092 1609
rect 1997 1541 2043 1575
rect 2077 1541 2092 1575
rect 1997 1507 2092 1541
rect 1997 1473 2043 1507
rect 2077 1473 2092 1507
rect 1997 1439 2092 1473
rect 1997 1405 2043 1439
rect 2077 1405 2092 1439
rect 1997 1371 2092 1405
rect 1997 1337 2043 1371
rect 2077 1337 2092 1371
rect 1997 1303 2092 1337
rect 1997 1269 2043 1303
rect 2077 1269 2092 1303
rect 1997 1235 2092 1269
rect 1997 1201 2043 1235
rect 2077 1201 2092 1235
rect 1997 1167 2092 1201
rect 1997 1133 2043 1167
rect 2077 1133 2092 1167
rect 1997 1099 2092 1133
rect 1997 1065 2043 1099
rect 2077 1065 2092 1099
rect 1997 1031 2092 1065
rect 1997 997 2043 1031
rect 2077 997 2092 1031
rect 1997 963 2092 997
rect 1997 929 2043 963
rect 2077 929 2092 963
rect 1997 895 2092 929
rect 1997 861 2043 895
rect 2077 861 2092 895
rect 1997 827 2092 861
rect 1997 793 2043 827
rect 2077 793 2092 827
rect 1997 759 2092 793
rect 1997 725 2043 759
rect 2077 725 2092 759
rect 1997 691 2092 725
rect 1997 657 2043 691
rect 2077 657 2092 691
rect 1997 623 2092 657
rect 1997 589 2043 623
rect 2077 589 2092 623
rect 1997 555 2092 589
rect 1997 521 2043 555
rect 2077 521 2092 555
rect 1997 487 2092 521
rect 1997 453 2043 487
rect 2077 453 2092 487
rect 1997 419 2092 453
rect 1997 385 2043 419
rect 2077 385 2092 419
rect 1997 351 2092 385
rect 1997 317 2043 351
rect 2077 317 2092 351
rect 1997 283 2092 317
rect 1997 249 2043 283
rect 2077 249 2092 283
rect 1997 215 2092 249
rect 1997 181 2043 215
rect 2077 181 2092 215
rect 1997 169 2092 181
<< mvndiffc >>
rect 191 2085 225 2119
rect 191 2017 225 2051
rect 191 1949 225 1983
rect 191 1881 225 1915
rect 191 1813 225 1847
rect 191 1745 225 1779
rect 191 1677 225 1711
rect 191 1609 225 1643
rect 191 1541 225 1575
rect 191 1473 225 1507
rect 191 1405 225 1439
rect 191 1337 225 1371
rect 191 1269 225 1303
rect 191 1201 225 1235
rect 191 1133 225 1167
rect 191 1065 225 1099
rect 191 997 225 1031
rect 191 929 225 963
rect 191 861 225 895
rect 191 793 225 827
rect 191 725 225 759
rect 191 657 225 691
rect 191 589 225 623
rect 191 521 225 555
rect 191 453 225 487
rect 191 385 225 419
rect 191 317 225 351
rect 191 249 225 283
rect 191 181 225 215
rect 1117 2085 1151 2119
rect 1117 2017 1151 2051
rect 1117 1949 1151 1983
rect 1117 1881 1151 1915
rect 1117 1813 1151 1847
rect 1117 1745 1151 1779
rect 1117 1677 1151 1711
rect 1117 1609 1151 1643
rect 1117 1541 1151 1575
rect 1117 1473 1151 1507
rect 1117 1405 1151 1439
rect 1117 1337 1151 1371
rect 1117 1269 1151 1303
rect 1117 1201 1151 1235
rect 1117 1133 1151 1167
rect 1117 1065 1151 1099
rect 1117 997 1151 1031
rect 1117 929 1151 963
rect 1117 861 1151 895
rect 1117 793 1151 827
rect 1117 725 1151 759
rect 1117 657 1151 691
rect 1117 589 1151 623
rect 1117 521 1151 555
rect 1117 453 1151 487
rect 1117 385 1151 419
rect 1117 317 1151 351
rect 1117 249 1151 283
rect 1117 181 1151 215
rect 2043 2085 2077 2119
rect 2043 2017 2077 2051
rect 2043 1949 2077 1983
rect 2043 1881 2077 1915
rect 2043 1813 2077 1847
rect 2043 1745 2077 1779
rect 2043 1677 2077 1711
rect 2043 1609 2077 1643
rect 2043 1541 2077 1575
rect 2043 1473 2077 1507
rect 2043 1405 2077 1439
rect 2043 1337 2077 1371
rect 2043 1269 2077 1303
rect 2043 1201 2077 1235
rect 2043 1133 2077 1167
rect 2043 1065 2077 1099
rect 2043 997 2077 1031
rect 2043 929 2077 963
rect 2043 861 2077 895
rect 2043 793 2077 827
rect 2043 725 2077 759
rect 2043 657 2077 691
rect 2043 589 2077 623
rect 2043 521 2077 555
rect 2043 453 2077 487
rect 2043 385 2077 419
rect 2043 317 2077 351
rect 2043 249 2077 283
rect 2043 181 2077 215
<< mvpsubdiff >>
rect 36 2131 176 2169
rect 36 2097 123 2131
rect 157 2097 176 2131
rect 36 2063 176 2097
rect 36 2029 123 2063
rect 157 2029 176 2063
rect 36 1995 176 2029
rect 36 1961 123 1995
rect 157 1961 176 1995
rect 36 1927 176 1961
rect 36 1893 123 1927
rect 157 1893 176 1927
rect 36 1859 176 1893
rect 36 1825 123 1859
rect 157 1825 176 1859
rect 36 1791 176 1825
rect 36 1757 123 1791
rect 157 1757 176 1791
rect 36 1723 176 1757
rect 36 1689 123 1723
rect 157 1689 176 1723
rect 36 1655 176 1689
rect 36 1621 123 1655
rect 157 1621 176 1655
rect 36 1587 176 1621
rect 36 1553 123 1587
rect 157 1553 176 1587
rect 36 1519 176 1553
rect 36 1485 123 1519
rect 157 1485 176 1519
rect 36 1451 176 1485
rect 36 1417 123 1451
rect 157 1417 176 1451
rect 36 1383 176 1417
rect 36 1349 123 1383
rect 157 1349 176 1383
rect 36 1315 176 1349
rect 36 1281 123 1315
rect 157 1281 176 1315
rect 36 1247 176 1281
rect 36 1213 123 1247
rect 157 1213 176 1247
rect 36 1179 176 1213
rect 36 1145 123 1179
rect 157 1145 176 1179
rect 36 1111 176 1145
rect 36 1077 123 1111
rect 157 1077 176 1111
rect 36 1043 176 1077
rect 36 1009 123 1043
rect 157 1009 176 1043
rect 36 975 176 1009
rect 36 941 123 975
rect 157 941 176 975
rect 36 907 176 941
rect 36 873 123 907
rect 157 873 176 907
rect 36 839 176 873
rect 36 805 123 839
rect 157 805 176 839
rect 36 771 176 805
rect 36 737 123 771
rect 157 737 176 771
rect 36 703 176 737
rect 36 669 123 703
rect 157 669 176 703
rect 36 635 176 669
rect 36 601 123 635
rect 157 601 176 635
rect 36 567 176 601
rect 36 533 123 567
rect 157 533 176 567
rect 36 499 176 533
rect 36 465 123 499
rect 157 465 176 499
rect 36 431 176 465
rect 36 397 123 431
rect 157 397 176 431
rect 36 363 176 397
rect 36 329 123 363
rect 157 329 176 363
rect 36 295 176 329
rect 36 261 123 295
rect 157 261 176 295
rect 36 227 176 261
rect 36 193 123 227
rect 157 193 176 227
rect 36 169 176 193
rect 2092 2131 2232 2169
rect 2092 2097 2111 2131
rect 2145 2097 2232 2131
rect 2092 2063 2232 2097
rect 2092 2029 2111 2063
rect 2145 2029 2232 2063
rect 2092 1995 2232 2029
rect 2092 1961 2111 1995
rect 2145 1961 2232 1995
rect 2092 1927 2232 1961
rect 2092 1893 2111 1927
rect 2145 1893 2232 1927
rect 2092 1859 2232 1893
rect 2092 1825 2111 1859
rect 2145 1825 2232 1859
rect 2092 1791 2232 1825
rect 2092 1757 2111 1791
rect 2145 1757 2232 1791
rect 2092 1723 2232 1757
rect 2092 1689 2111 1723
rect 2145 1689 2232 1723
rect 2092 1655 2232 1689
rect 2092 1621 2111 1655
rect 2145 1621 2232 1655
rect 2092 1587 2232 1621
rect 2092 1553 2111 1587
rect 2145 1553 2232 1587
rect 2092 1519 2232 1553
rect 2092 1485 2111 1519
rect 2145 1485 2232 1519
rect 2092 1451 2232 1485
rect 2092 1417 2111 1451
rect 2145 1417 2232 1451
rect 2092 1383 2232 1417
rect 2092 1349 2111 1383
rect 2145 1349 2232 1383
rect 2092 1315 2232 1349
rect 2092 1281 2111 1315
rect 2145 1281 2232 1315
rect 2092 1247 2232 1281
rect 2092 1213 2111 1247
rect 2145 1213 2232 1247
rect 2092 1179 2232 1213
rect 2092 1145 2111 1179
rect 2145 1145 2232 1179
rect 2092 1111 2232 1145
rect 2092 1077 2111 1111
rect 2145 1077 2232 1111
rect 2092 1043 2232 1077
rect 2092 1009 2111 1043
rect 2145 1009 2232 1043
rect 2092 975 2232 1009
rect 2092 941 2111 975
rect 2145 941 2232 975
rect 2092 907 2232 941
rect 2092 873 2111 907
rect 2145 873 2232 907
rect 2092 839 2232 873
rect 2092 805 2111 839
rect 2145 805 2232 839
rect 2092 771 2232 805
rect 2092 737 2111 771
rect 2145 737 2232 771
rect 2092 703 2232 737
rect 2092 669 2111 703
rect 2145 669 2232 703
rect 2092 635 2232 669
rect 2092 601 2111 635
rect 2145 601 2232 635
rect 2092 567 2232 601
rect 2092 533 2111 567
rect 2145 533 2232 567
rect 2092 499 2232 533
rect 2092 465 2111 499
rect 2145 465 2232 499
rect 2092 431 2232 465
rect 2092 397 2111 431
rect 2145 397 2232 431
rect 2092 363 2232 397
rect 2092 329 2111 363
rect 2145 329 2232 363
rect 2092 295 2232 329
rect 2092 261 2111 295
rect 2145 261 2232 295
rect 2092 227 2232 261
rect 2092 193 2111 227
rect 2145 193 2232 227
rect 2092 169 2232 193
<< mvpsubdiffcont >>
rect 123 2097 157 2131
rect 123 2029 157 2063
rect 123 1961 157 1995
rect 123 1893 157 1927
rect 123 1825 157 1859
rect 123 1757 157 1791
rect 123 1689 157 1723
rect 123 1621 157 1655
rect 123 1553 157 1587
rect 123 1485 157 1519
rect 123 1417 157 1451
rect 123 1349 157 1383
rect 123 1281 157 1315
rect 123 1213 157 1247
rect 123 1145 157 1179
rect 123 1077 157 1111
rect 123 1009 157 1043
rect 123 941 157 975
rect 123 873 157 907
rect 123 805 157 839
rect 123 737 157 771
rect 123 669 157 703
rect 123 601 157 635
rect 123 533 157 567
rect 123 465 157 499
rect 123 397 157 431
rect 123 329 157 363
rect 123 261 157 295
rect 123 193 157 227
rect 2111 2097 2145 2131
rect 2111 2029 2145 2063
rect 2111 1961 2145 1995
rect 2111 1893 2145 1927
rect 2111 1825 2145 1859
rect 2111 1757 2145 1791
rect 2111 1689 2145 1723
rect 2111 1621 2145 1655
rect 2111 1553 2145 1587
rect 2111 1485 2145 1519
rect 2111 1417 2145 1451
rect 2111 1349 2145 1383
rect 2111 1281 2145 1315
rect 2111 1213 2145 1247
rect 2111 1145 2145 1179
rect 2111 1077 2145 1111
rect 2111 1009 2145 1043
rect 2111 941 2145 975
rect 2111 873 2145 907
rect 2111 805 2145 839
rect 2111 737 2145 771
rect 2111 669 2145 703
rect 2111 601 2145 635
rect 2111 533 2145 567
rect 2111 465 2145 499
rect 2111 397 2145 431
rect 2111 329 2145 363
rect 2111 261 2145 295
rect 2111 193 2145 227
<< poly >>
rect 271 2271 1997 2287
rect 271 2237 291 2271
rect 325 2237 359 2271
rect 393 2237 427 2271
rect 461 2237 495 2271
rect 529 2237 563 2271
rect 597 2237 631 2271
rect 665 2237 699 2271
rect 733 2237 767 2271
rect 801 2237 835 2271
rect 869 2237 903 2271
rect 937 2237 971 2271
rect 1005 2237 1039 2271
rect 1073 2237 1107 2271
rect 1141 2237 1175 2271
rect 1209 2237 1243 2271
rect 1277 2237 1311 2271
rect 1345 2237 1379 2271
rect 1413 2237 1447 2271
rect 1481 2237 1515 2271
rect 1549 2237 1583 2271
rect 1617 2237 1651 2271
rect 1685 2237 1719 2271
rect 1753 2237 1787 2271
rect 1821 2237 1855 2271
rect 1889 2237 1923 2271
rect 1957 2237 1997 2271
rect 271 2221 1997 2237
rect 271 2169 1071 2221
rect 1197 2169 1997 2221
rect 271 117 1071 169
rect 1197 117 1997 169
rect 271 101 1997 117
rect 271 67 291 101
rect 325 67 359 101
rect 393 67 427 101
rect 461 67 495 101
rect 529 67 563 101
rect 597 67 631 101
rect 665 67 699 101
rect 733 67 767 101
rect 801 67 835 101
rect 869 67 903 101
rect 937 67 971 101
rect 1005 67 1039 101
rect 1073 67 1107 101
rect 1141 67 1175 101
rect 1209 67 1243 101
rect 1277 67 1311 101
rect 1345 67 1379 101
rect 1413 67 1447 101
rect 1481 67 1515 101
rect 1549 67 1583 101
rect 1617 67 1651 101
rect 1685 67 1719 101
rect 1753 67 1787 101
rect 1821 67 1855 101
rect 1889 67 1923 101
rect 1957 67 1997 101
rect 271 51 1997 67
<< polycont >>
rect 291 2237 325 2271
rect 359 2237 393 2271
rect 427 2237 461 2271
rect 495 2237 529 2271
rect 563 2237 597 2271
rect 631 2237 665 2271
rect 699 2237 733 2271
rect 767 2237 801 2271
rect 835 2237 869 2271
rect 903 2237 937 2271
rect 971 2237 1005 2271
rect 1039 2237 1073 2271
rect 1107 2237 1141 2271
rect 1175 2237 1209 2271
rect 1243 2237 1277 2271
rect 1311 2237 1345 2271
rect 1379 2237 1413 2271
rect 1447 2237 1481 2271
rect 1515 2237 1549 2271
rect 1583 2237 1617 2271
rect 1651 2237 1685 2271
rect 1719 2237 1753 2271
rect 1787 2237 1821 2271
rect 1855 2237 1889 2271
rect 1923 2237 1957 2271
rect 291 67 325 101
rect 359 67 393 101
rect 427 67 461 101
rect 495 67 529 101
rect 563 67 597 101
rect 631 67 665 101
rect 699 67 733 101
rect 767 67 801 101
rect 835 67 869 101
rect 903 67 937 101
rect 971 67 1005 101
rect 1039 67 1073 101
rect 1107 67 1141 101
rect 1175 67 1209 101
rect 1243 67 1277 101
rect 1311 67 1345 101
rect 1379 67 1413 101
rect 1447 67 1481 101
rect 1515 67 1549 101
rect 1583 67 1617 101
rect 1651 67 1685 101
rect 1719 67 1753 101
rect 1787 67 1821 101
rect 1855 67 1889 101
rect 1923 67 1957 101
<< locali >>
rect 271 2271 1996 2280
rect 271 2237 283 2271
rect 325 2237 355 2271
rect 393 2237 427 2271
rect 461 2237 495 2271
rect 533 2237 563 2271
rect 605 2237 631 2271
rect 677 2237 699 2271
rect 749 2237 767 2271
rect 821 2237 835 2271
rect 893 2237 903 2271
rect 965 2237 971 2271
rect 1037 2237 1039 2271
rect 1073 2237 1075 2271
rect 1141 2237 1147 2271
rect 1209 2237 1219 2271
rect 1277 2237 1291 2271
rect 1345 2237 1363 2271
rect 1413 2237 1435 2271
rect 1481 2237 1507 2271
rect 1549 2237 1579 2271
rect 1617 2237 1651 2271
rect 1685 2237 1719 2271
rect 1757 2237 1787 2271
rect 1829 2237 1855 2271
rect 1901 2237 1923 2271
rect 1973 2237 1997 2271
rect 271 2228 1996 2237
rect 93 2131 2175 2147
rect 93 2097 123 2131
rect 157 2119 2111 2131
rect 157 2109 191 2119
rect 225 2109 1117 2119
rect 93 2063 129 2097
rect 235 2085 1117 2109
rect 1151 2109 2043 2119
rect 2077 2109 2111 2119
rect 1151 2085 2033 2109
rect 2145 2097 2175 2131
rect 93 2029 123 2063
rect 235 2051 2033 2085
rect 2139 2063 2175 2097
rect 93 1995 129 2029
rect 235 2031 1117 2051
rect 235 1997 319 2031
rect 353 1997 391 2031
rect 425 1997 463 2031
rect 497 1997 535 2031
rect 569 1997 607 2031
rect 641 1997 679 2031
rect 713 1997 751 2031
rect 785 1997 823 2031
rect 857 1997 895 2031
rect 929 1997 967 2031
rect 1001 2017 1117 2031
rect 1151 2031 2033 2051
rect 1151 2017 1267 2031
rect 1001 1997 1267 2017
rect 1301 1997 1339 2031
rect 1373 1997 1411 2031
rect 1445 1997 1483 2031
rect 1517 1997 1555 2031
rect 1589 1997 1627 2031
rect 1661 1997 1699 2031
rect 1733 1997 1771 2031
rect 1805 1997 1843 2031
rect 1877 1997 1915 2031
rect 1949 1997 2033 2031
rect 2145 2029 2175 2063
rect 93 1961 123 1995
rect 235 1987 2033 1997
rect 2139 1995 2175 2029
rect 93 1927 129 1961
rect 93 1893 123 1927
rect 93 1859 129 1893
rect 93 1825 123 1859
rect 93 1791 129 1825
rect 93 1757 123 1791
rect 93 1723 129 1757
rect 93 1689 123 1723
rect 93 1655 129 1689
rect 93 1621 123 1655
rect 93 1587 129 1621
rect 93 1553 123 1587
rect 93 1519 129 1553
rect 93 1485 123 1519
rect 93 1451 129 1485
rect 93 1417 123 1451
rect 93 1383 129 1417
rect 93 1349 123 1383
rect 93 1315 129 1349
rect 93 1281 123 1315
rect 93 1247 129 1281
rect 93 1213 123 1247
rect 93 1179 129 1213
rect 93 1145 123 1179
rect 93 1111 129 1145
rect 93 1077 123 1111
rect 93 1043 129 1077
rect 93 1009 123 1043
rect 93 975 129 1009
rect 93 941 123 975
rect 93 907 129 941
rect 93 873 123 907
rect 93 839 129 873
rect 93 805 123 839
rect 93 771 129 805
rect 93 737 123 771
rect 93 703 129 737
rect 93 669 123 703
rect 93 635 129 669
rect 93 601 123 635
rect 93 567 129 601
rect 93 533 123 567
rect 93 499 129 533
rect 93 465 123 499
rect 93 431 129 465
rect 93 397 123 431
rect 93 363 129 397
rect 93 329 123 363
rect 290 1219 324 1953
rect 360 1253 394 1987
rect 430 1219 464 1953
rect 500 1253 534 1987
rect 570 1219 604 1953
rect 640 1253 674 1987
rect 710 1219 744 1953
rect 780 1253 814 1987
rect 850 1219 884 1953
rect 920 1253 954 1987
rect 1060 1983 1208 1987
rect 990 1219 1024 1953
rect 1060 1949 1117 1983
rect 1151 1949 1208 1983
rect 1060 1915 1208 1949
rect 1060 1881 1117 1915
rect 1151 1881 1208 1915
rect 1060 1847 1208 1881
rect 1060 1813 1117 1847
rect 1151 1813 1208 1847
rect 1060 1779 1208 1813
rect 1060 1745 1117 1779
rect 1151 1745 1208 1779
rect 1060 1711 1208 1745
rect 1060 1677 1117 1711
rect 1151 1677 1208 1711
rect 1060 1643 1208 1677
rect 1060 1609 1117 1643
rect 1151 1609 1208 1643
rect 1060 1575 1208 1609
rect 1060 1541 1117 1575
rect 1151 1541 1208 1575
rect 1060 1507 1208 1541
rect 1060 1473 1117 1507
rect 1151 1473 1208 1507
rect 1060 1439 1208 1473
rect 1060 1405 1117 1439
rect 1151 1405 1208 1439
rect 1060 1371 1208 1405
rect 1060 1337 1117 1371
rect 1151 1337 1208 1371
rect 1060 1303 1208 1337
rect 1060 1269 1117 1303
rect 1151 1269 1208 1303
rect 1060 1256 1208 1269
rect 1060 1255 1180 1256
rect 1088 1235 1180 1255
rect 290 1209 1052 1219
rect 290 1103 344 1209
rect 1026 1103 1052 1209
rect 290 1093 1052 1103
rect 1088 1201 1117 1235
rect 1151 1201 1180 1235
rect 1244 1219 1278 1953
rect 1314 1253 1348 1987
rect 1384 1219 1418 1953
rect 1454 1253 1488 1987
rect 1524 1219 1558 1953
rect 1594 1253 1628 1987
rect 1664 1219 1698 1953
rect 1734 1253 1768 1987
rect 1804 1219 1838 1953
rect 1874 1253 1908 1987
rect 1944 1219 1978 1953
rect 1088 1167 1180 1201
rect 1088 1133 1117 1167
rect 1151 1133 1180 1167
rect 1088 1099 1180 1133
rect 290 359 324 1093
rect 93 295 129 329
rect 360 325 394 1059
rect 430 359 464 1093
rect 500 325 534 1059
rect 570 359 604 1093
rect 640 325 674 1059
rect 710 359 744 1093
rect 780 325 814 1059
rect 850 359 884 1093
rect 920 325 954 1059
rect 990 359 1024 1093
rect 1088 1065 1117 1099
rect 1151 1065 1180 1099
rect 1216 1209 1978 1219
rect 1216 1103 1242 1209
rect 1924 1103 1978 1209
rect 1216 1093 1978 1103
rect 1088 1057 1180 1065
rect 1060 1031 1208 1057
rect 1060 997 1117 1031
rect 1151 997 1208 1031
rect 1060 963 1208 997
rect 1060 929 1117 963
rect 1151 929 1208 963
rect 1060 895 1208 929
rect 1060 861 1117 895
rect 1151 861 1208 895
rect 1060 827 1208 861
rect 1060 793 1117 827
rect 1151 793 1208 827
rect 1060 759 1208 793
rect 1060 725 1117 759
rect 1151 725 1208 759
rect 1060 691 1208 725
rect 1060 657 1117 691
rect 1151 657 1208 691
rect 1060 623 1208 657
rect 1060 589 1117 623
rect 1151 589 1208 623
rect 1060 555 1208 589
rect 1060 521 1117 555
rect 1151 521 1208 555
rect 1060 487 1208 521
rect 1060 453 1117 487
rect 1151 453 1208 487
rect 1060 419 1208 453
rect 1060 385 1117 419
rect 1151 385 1208 419
rect 1060 351 1208 385
rect 1244 359 1278 1093
rect 1060 325 1117 351
rect 235 317 1117 325
rect 1151 325 1208 351
rect 1314 325 1348 1059
rect 1384 359 1418 1093
rect 1454 325 1488 1059
rect 1524 359 1558 1093
rect 1594 325 1628 1059
rect 1664 359 1698 1093
rect 1734 325 1768 1059
rect 1804 359 1838 1093
rect 1874 325 1908 1059
rect 1944 359 1978 1093
rect 2145 1961 2175 1995
rect 2139 1927 2175 1961
rect 2145 1893 2175 1927
rect 2139 1859 2175 1893
rect 2145 1825 2175 1859
rect 2139 1791 2175 1825
rect 2145 1757 2175 1791
rect 2139 1723 2175 1757
rect 2145 1689 2175 1723
rect 2139 1655 2175 1689
rect 2145 1621 2175 1655
rect 2139 1587 2175 1621
rect 2145 1553 2175 1587
rect 2139 1519 2175 1553
rect 2145 1485 2175 1519
rect 2139 1451 2175 1485
rect 2145 1417 2175 1451
rect 2139 1383 2175 1417
rect 2145 1349 2175 1383
rect 2139 1315 2175 1349
rect 2145 1281 2175 1315
rect 2139 1247 2175 1281
rect 2145 1213 2175 1247
rect 2139 1179 2175 1213
rect 2145 1145 2175 1179
rect 2139 1111 2175 1145
rect 2145 1077 2175 1111
rect 2139 1043 2175 1077
rect 2145 1009 2175 1043
rect 2139 975 2175 1009
rect 2145 941 2175 975
rect 2139 907 2175 941
rect 2145 873 2175 907
rect 2139 839 2175 873
rect 2145 805 2175 839
rect 2139 771 2175 805
rect 2145 737 2175 771
rect 2139 703 2175 737
rect 2145 669 2175 703
rect 2139 635 2175 669
rect 2145 601 2175 635
rect 2139 567 2175 601
rect 2145 533 2175 567
rect 2139 499 2175 533
rect 2145 465 2175 499
rect 2139 431 2175 465
rect 2145 397 2175 431
rect 2139 363 2175 397
rect 1151 317 2033 325
rect 2145 329 2175 363
rect 235 315 2033 317
rect 93 261 123 295
rect 93 227 129 261
rect 235 281 319 315
rect 353 281 391 315
rect 425 281 463 315
rect 497 281 535 315
rect 569 281 607 315
rect 641 281 679 315
rect 713 281 751 315
rect 785 281 823 315
rect 857 281 895 315
rect 929 281 967 315
rect 1001 283 1267 315
rect 1001 281 1117 283
rect 235 249 1117 281
rect 1151 281 1267 283
rect 1301 281 1339 315
rect 1373 281 1411 315
rect 1445 281 1483 315
rect 1517 281 1555 315
rect 1589 281 1627 315
rect 1661 281 1699 315
rect 1733 281 1771 315
rect 1805 281 1843 315
rect 1877 281 1915 315
rect 1949 281 2033 315
rect 2139 295 2175 329
rect 1151 249 2033 281
rect 2145 261 2175 295
rect 93 193 123 227
rect 235 215 2033 249
rect 2139 227 2175 261
rect 235 203 1117 215
rect 157 193 191 203
rect 93 181 191 193
rect 225 181 1117 203
rect 1151 203 2033 215
rect 1151 181 2043 203
rect 2077 193 2111 203
rect 2145 193 2175 227
rect 2077 181 2175 193
rect 93 165 2175 181
rect 271 101 1996 110
rect 271 67 283 101
rect 325 67 355 101
rect 393 67 427 101
rect 461 67 495 101
rect 533 67 563 101
rect 605 67 631 101
rect 677 67 699 101
rect 749 67 767 101
rect 821 67 835 101
rect 893 67 903 101
rect 965 67 971 101
rect 1037 67 1039 101
rect 1073 67 1075 101
rect 1141 67 1147 101
rect 1209 67 1219 101
rect 1277 67 1291 101
rect 1345 67 1363 101
rect 1413 67 1435 101
rect 1481 67 1507 101
rect 1549 67 1579 101
rect 1617 67 1651 101
rect 1685 67 1719 101
rect 1757 67 1787 101
rect 1829 67 1855 101
rect 1901 67 1923 101
rect 1973 67 1997 101
rect 271 58 1996 67
<< viali >>
rect 283 2237 291 2271
rect 291 2237 317 2271
rect 355 2237 359 2271
rect 359 2237 389 2271
rect 427 2237 461 2271
rect 499 2237 529 2271
rect 529 2237 533 2271
rect 571 2237 597 2271
rect 597 2237 605 2271
rect 643 2237 665 2271
rect 665 2237 677 2271
rect 715 2237 733 2271
rect 733 2237 749 2271
rect 787 2237 801 2271
rect 801 2237 821 2271
rect 859 2237 869 2271
rect 869 2237 893 2271
rect 931 2237 937 2271
rect 937 2237 965 2271
rect 1003 2237 1005 2271
rect 1005 2237 1037 2271
rect 1075 2237 1107 2271
rect 1107 2237 1109 2271
rect 1147 2237 1175 2271
rect 1175 2237 1181 2271
rect 1219 2237 1243 2271
rect 1243 2237 1253 2271
rect 1291 2237 1311 2271
rect 1311 2237 1325 2271
rect 1363 2237 1379 2271
rect 1379 2237 1397 2271
rect 1435 2237 1447 2271
rect 1447 2237 1469 2271
rect 1507 2237 1515 2271
rect 1515 2237 1541 2271
rect 1579 2237 1583 2271
rect 1583 2237 1613 2271
rect 1651 2237 1685 2271
rect 1723 2237 1753 2271
rect 1753 2237 1757 2271
rect 1795 2237 1821 2271
rect 1821 2237 1829 2271
rect 1867 2237 1889 2271
rect 1889 2237 1901 2271
rect 1939 2237 1957 2271
rect 1957 2237 1973 2271
rect 129 2097 157 2109
rect 157 2097 191 2109
rect 129 2085 191 2097
rect 191 2085 225 2109
rect 225 2085 235 2109
rect 2033 2085 2043 2109
rect 2043 2085 2077 2109
rect 2077 2097 2111 2109
rect 2111 2097 2139 2109
rect 2077 2085 2139 2097
rect 129 2063 235 2085
rect 129 2029 157 2063
rect 157 2051 235 2063
rect 2033 2063 2139 2085
rect 2033 2051 2111 2063
rect 157 2029 191 2051
rect 129 2017 191 2029
rect 191 2017 225 2051
rect 225 2017 235 2051
rect 129 1995 235 2017
rect 319 1997 353 2031
rect 391 1997 425 2031
rect 463 1997 497 2031
rect 535 1997 569 2031
rect 607 1997 641 2031
rect 679 1997 713 2031
rect 751 1997 785 2031
rect 823 1997 857 2031
rect 895 1997 929 2031
rect 967 1997 1001 2031
rect 1267 1997 1301 2031
rect 1339 1997 1373 2031
rect 1411 1997 1445 2031
rect 1483 1997 1517 2031
rect 1555 1997 1589 2031
rect 1627 1997 1661 2031
rect 1699 1997 1733 2031
rect 1771 1997 1805 2031
rect 1843 1997 1877 2031
rect 1915 1997 1949 2031
rect 2033 2017 2043 2051
rect 2043 2017 2077 2051
rect 2077 2029 2111 2051
rect 2111 2029 2139 2063
rect 2077 2017 2139 2029
rect 129 1961 157 1995
rect 157 1983 235 1995
rect 2033 1995 2139 2017
rect 157 1961 191 1983
rect 129 1949 191 1961
rect 191 1949 225 1983
rect 225 1949 235 1983
rect 129 1927 235 1949
rect 129 1893 157 1927
rect 157 1915 235 1927
rect 157 1893 191 1915
rect 129 1881 191 1893
rect 191 1881 225 1915
rect 225 1881 235 1915
rect 129 1859 235 1881
rect 129 1825 157 1859
rect 157 1847 235 1859
rect 157 1825 191 1847
rect 129 1813 191 1825
rect 191 1813 225 1847
rect 225 1813 235 1847
rect 129 1791 235 1813
rect 129 1757 157 1791
rect 157 1779 235 1791
rect 157 1757 191 1779
rect 129 1745 191 1757
rect 191 1745 225 1779
rect 225 1745 235 1779
rect 129 1723 235 1745
rect 129 1689 157 1723
rect 157 1711 235 1723
rect 157 1689 191 1711
rect 129 1677 191 1689
rect 191 1677 225 1711
rect 225 1677 235 1711
rect 129 1655 235 1677
rect 129 1621 157 1655
rect 157 1643 235 1655
rect 157 1621 191 1643
rect 129 1609 191 1621
rect 191 1609 225 1643
rect 225 1609 235 1643
rect 129 1587 235 1609
rect 129 1553 157 1587
rect 157 1575 235 1587
rect 157 1553 191 1575
rect 129 1541 191 1553
rect 191 1541 225 1575
rect 225 1541 235 1575
rect 129 1519 235 1541
rect 129 1485 157 1519
rect 157 1507 235 1519
rect 157 1485 191 1507
rect 129 1473 191 1485
rect 191 1473 225 1507
rect 225 1473 235 1507
rect 129 1451 235 1473
rect 129 1417 157 1451
rect 157 1439 235 1451
rect 157 1417 191 1439
rect 129 1405 191 1417
rect 191 1405 225 1439
rect 225 1405 235 1439
rect 129 1383 235 1405
rect 129 1349 157 1383
rect 157 1371 235 1383
rect 157 1349 191 1371
rect 129 1337 191 1349
rect 191 1337 225 1371
rect 225 1337 235 1371
rect 129 1315 235 1337
rect 129 1281 157 1315
rect 157 1303 235 1315
rect 157 1281 191 1303
rect 129 1269 191 1281
rect 191 1269 225 1303
rect 225 1269 235 1303
rect 129 1247 235 1269
rect 129 1213 157 1247
rect 157 1235 235 1247
rect 157 1213 191 1235
rect 129 1201 191 1213
rect 191 1201 225 1235
rect 225 1201 235 1235
rect 129 1179 235 1201
rect 129 1145 157 1179
rect 157 1167 235 1179
rect 157 1145 191 1167
rect 129 1133 191 1145
rect 191 1133 225 1167
rect 225 1133 235 1167
rect 129 1111 235 1133
rect 129 1077 157 1111
rect 157 1099 235 1111
rect 157 1077 191 1099
rect 129 1065 191 1077
rect 191 1065 225 1099
rect 225 1065 235 1099
rect 129 1043 235 1065
rect 129 1009 157 1043
rect 157 1031 235 1043
rect 157 1009 191 1031
rect 129 997 191 1009
rect 191 997 225 1031
rect 225 997 235 1031
rect 129 975 235 997
rect 129 941 157 975
rect 157 963 235 975
rect 157 941 191 963
rect 129 929 191 941
rect 191 929 225 963
rect 225 929 235 963
rect 129 907 235 929
rect 129 873 157 907
rect 157 895 235 907
rect 157 873 191 895
rect 129 861 191 873
rect 191 861 225 895
rect 225 861 235 895
rect 129 839 235 861
rect 129 805 157 839
rect 157 827 235 839
rect 157 805 191 827
rect 129 793 191 805
rect 191 793 225 827
rect 225 793 235 827
rect 129 771 235 793
rect 129 737 157 771
rect 157 759 235 771
rect 157 737 191 759
rect 129 725 191 737
rect 191 725 225 759
rect 225 725 235 759
rect 129 703 235 725
rect 129 669 157 703
rect 157 691 235 703
rect 157 669 191 691
rect 129 657 191 669
rect 191 657 225 691
rect 225 657 235 691
rect 129 635 235 657
rect 129 601 157 635
rect 157 623 235 635
rect 157 601 191 623
rect 129 589 191 601
rect 191 589 225 623
rect 225 589 235 623
rect 129 567 235 589
rect 129 533 157 567
rect 157 555 235 567
rect 157 533 191 555
rect 129 521 191 533
rect 191 521 225 555
rect 225 521 235 555
rect 129 499 235 521
rect 129 465 157 499
rect 157 487 235 499
rect 157 465 191 487
rect 129 453 191 465
rect 191 453 225 487
rect 225 453 235 487
rect 129 431 235 453
rect 129 397 157 431
rect 157 419 235 431
rect 157 397 191 419
rect 129 385 191 397
rect 191 385 225 419
rect 225 385 235 419
rect 129 363 235 385
rect 129 329 157 363
rect 157 351 235 363
rect 344 1103 1026 1209
rect 2033 1983 2111 1995
rect 157 329 191 351
rect 129 317 191 329
rect 191 317 225 351
rect 225 317 235 351
rect 1242 1103 1924 1209
rect 2033 1949 2043 1983
rect 2043 1949 2077 1983
rect 2077 1961 2111 1983
rect 2111 1961 2139 1995
rect 2077 1949 2139 1961
rect 2033 1927 2139 1949
rect 2033 1915 2111 1927
rect 2033 1881 2043 1915
rect 2043 1881 2077 1915
rect 2077 1893 2111 1915
rect 2111 1893 2139 1927
rect 2077 1881 2139 1893
rect 2033 1859 2139 1881
rect 2033 1847 2111 1859
rect 2033 1813 2043 1847
rect 2043 1813 2077 1847
rect 2077 1825 2111 1847
rect 2111 1825 2139 1859
rect 2077 1813 2139 1825
rect 2033 1791 2139 1813
rect 2033 1779 2111 1791
rect 2033 1745 2043 1779
rect 2043 1745 2077 1779
rect 2077 1757 2111 1779
rect 2111 1757 2139 1791
rect 2077 1745 2139 1757
rect 2033 1723 2139 1745
rect 2033 1711 2111 1723
rect 2033 1677 2043 1711
rect 2043 1677 2077 1711
rect 2077 1689 2111 1711
rect 2111 1689 2139 1723
rect 2077 1677 2139 1689
rect 2033 1655 2139 1677
rect 2033 1643 2111 1655
rect 2033 1609 2043 1643
rect 2043 1609 2077 1643
rect 2077 1621 2111 1643
rect 2111 1621 2139 1655
rect 2077 1609 2139 1621
rect 2033 1587 2139 1609
rect 2033 1575 2111 1587
rect 2033 1541 2043 1575
rect 2043 1541 2077 1575
rect 2077 1553 2111 1575
rect 2111 1553 2139 1587
rect 2077 1541 2139 1553
rect 2033 1519 2139 1541
rect 2033 1507 2111 1519
rect 2033 1473 2043 1507
rect 2043 1473 2077 1507
rect 2077 1485 2111 1507
rect 2111 1485 2139 1519
rect 2077 1473 2139 1485
rect 2033 1451 2139 1473
rect 2033 1439 2111 1451
rect 2033 1405 2043 1439
rect 2043 1405 2077 1439
rect 2077 1417 2111 1439
rect 2111 1417 2139 1451
rect 2077 1405 2139 1417
rect 2033 1383 2139 1405
rect 2033 1371 2111 1383
rect 2033 1337 2043 1371
rect 2043 1337 2077 1371
rect 2077 1349 2111 1371
rect 2111 1349 2139 1383
rect 2077 1337 2139 1349
rect 2033 1315 2139 1337
rect 2033 1303 2111 1315
rect 2033 1269 2043 1303
rect 2043 1269 2077 1303
rect 2077 1281 2111 1303
rect 2111 1281 2139 1315
rect 2077 1269 2139 1281
rect 2033 1247 2139 1269
rect 2033 1235 2111 1247
rect 2033 1201 2043 1235
rect 2043 1201 2077 1235
rect 2077 1213 2111 1235
rect 2111 1213 2139 1247
rect 2077 1201 2139 1213
rect 2033 1179 2139 1201
rect 2033 1167 2111 1179
rect 2033 1133 2043 1167
rect 2043 1133 2077 1167
rect 2077 1145 2111 1167
rect 2111 1145 2139 1179
rect 2077 1133 2139 1145
rect 2033 1111 2139 1133
rect 2033 1099 2111 1111
rect 2033 1065 2043 1099
rect 2043 1065 2077 1099
rect 2077 1077 2111 1099
rect 2111 1077 2139 1111
rect 2077 1065 2139 1077
rect 2033 1043 2139 1065
rect 2033 1031 2111 1043
rect 2033 997 2043 1031
rect 2043 997 2077 1031
rect 2077 1009 2111 1031
rect 2111 1009 2139 1043
rect 2077 997 2139 1009
rect 2033 975 2139 997
rect 2033 963 2111 975
rect 2033 929 2043 963
rect 2043 929 2077 963
rect 2077 941 2111 963
rect 2111 941 2139 975
rect 2077 929 2139 941
rect 2033 907 2139 929
rect 2033 895 2111 907
rect 2033 861 2043 895
rect 2043 861 2077 895
rect 2077 873 2111 895
rect 2111 873 2139 907
rect 2077 861 2139 873
rect 2033 839 2139 861
rect 2033 827 2111 839
rect 2033 793 2043 827
rect 2043 793 2077 827
rect 2077 805 2111 827
rect 2111 805 2139 839
rect 2077 793 2139 805
rect 2033 771 2139 793
rect 2033 759 2111 771
rect 2033 725 2043 759
rect 2043 725 2077 759
rect 2077 737 2111 759
rect 2111 737 2139 771
rect 2077 725 2139 737
rect 2033 703 2139 725
rect 2033 691 2111 703
rect 2033 657 2043 691
rect 2043 657 2077 691
rect 2077 669 2111 691
rect 2111 669 2139 703
rect 2077 657 2139 669
rect 2033 635 2139 657
rect 2033 623 2111 635
rect 2033 589 2043 623
rect 2043 589 2077 623
rect 2077 601 2111 623
rect 2111 601 2139 635
rect 2077 589 2139 601
rect 2033 567 2139 589
rect 2033 555 2111 567
rect 2033 521 2043 555
rect 2043 521 2077 555
rect 2077 533 2111 555
rect 2111 533 2139 567
rect 2077 521 2139 533
rect 2033 499 2139 521
rect 2033 487 2111 499
rect 2033 453 2043 487
rect 2043 453 2077 487
rect 2077 465 2111 487
rect 2111 465 2139 499
rect 2077 453 2139 465
rect 2033 431 2139 453
rect 2033 419 2111 431
rect 2033 385 2043 419
rect 2043 385 2077 419
rect 2077 397 2111 419
rect 2111 397 2139 431
rect 2077 385 2139 397
rect 2033 363 2139 385
rect 2033 351 2111 363
rect 2033 317 2043 351
rect 2043 317 2077 351
rect 2077 329 2111 351
rect 2111 329 2139 363
rect 2077 317 2139 329
rect 129 295 235 317
rect 129 261 157 295
rect 157 283 235 295
rect 157 261 191 283
rect 129 249 191 261
rect 191 249 225 283
rect 225 249 235 283
rect 319 281 353 315
rect 391 281 425 315
rect 463 281 497 315
rect 535 281 569 315
rect 607 281 641 315
rect 679 281 713 315
rect 751 281 785 315
rect 823 281 857 315
rect 895 281 929 315
rect 967 281 1001 315
rect 1267 281 1301 315
rect 1339 281 1373 315
rect 1411 281 1445 315
rect 1483 281 1517 315
rect 1555 281 1589 315
rect 1627 281 1661 315
rect 1699 281 1733 315
rect 1771 281 1805 315
rect 1843 281 1877 315
rect 1915 281 1949 315
rect 2033 295 2139 317
rect 2033 283 2111 295
rect 2033 249 2043 283
rect 2043 249 2077 283
rect 2077 261 2111 283
rect 2111 261 2139 295
rect 2077 249 2139 261
rect 129 227 235 249
rect 129 203 157 227
rect 157 215 235 227
rect 2033 227 2139 249
rect 2033 215 2111 227
rect 157 203 191 215
rect 191 203 225 215
rect 225 203 235 215
rect 2033 203 2043 215
rect 2043 203 2077 215
rect 2077 203 2111 215
rect 2111 203 2139 227
rect 283 67 291 101
rect 291 67 317 101
rect 355 67 359 101
rect 359 67 389 101
rect 427 67 461 101
rect 499 67 529 101
rect 529 67 533 101
rect 571 67 597 101
rect 597 67 605 101
rect 643 67 665 101
rect 665 67 677 101
rect 715 67 733 101
rect 733 67 749 101
rect 787 67 801 101
rect 801 67 821 101
rect 859 67 869 101
rect 869 67 893 101
rect 931 67 937 101
rect 937 67 965 101
rect 1003 67 1005 101
rect 1005 67 1037 101
rect 1075 67 1107 101
rect 1107 67 1109 101
rect 1147 67 1175 101
rect 1175 67 1181 101
rect 1219 67 1243 101
rect 1243 67 1253 101
rect 1291 67 1311 101
rect 1311 67 1325 101
rect 1363 67 1379 101
rect 1379 67 1397 101
rect 1435 67 1447 101
rect 1447 67 1469 101
rect 1507 67 1515 101
rect 1515 67 1541 101
rect 1579 67 1583 101
rect 1583 67 1613 101
rect 1651 67 1685 101
rect 1723 67 1753 101
rect 1753 67 1757 101
rect 1795 67 1821 101
rect 1821 67 1829 101
rect 1867 67 1889 101
rect 1889 67 1901 101
rect 1939 67 1957 101
rect 1957 67 1973 101
<< metal1 >>
rect 93 2308 2175 2338
rect 93 2109 243 2308
rect 93 203 129 2109
rect 235 2041 243 2109
rect 271 2228 277 2280
rect 329 2228 341 2280
rect 393 2228 405 2280
rect 457 2271 469 2280
rect 521 2271 533 2280
rect 585 2271 597 2280
rect 649 2271 661 2280
rect 713 2271 725 2280
rect 777 2271 789 2280
rect 461 2237 469 2271
rect 713 2237 715 2271
rect 777 2237 787 2271
rect 457 2228 469 2237
rect 521 2228 533 2237
rect 585 2228 597 2237
rect 649 2228 661 2237
rect 713 2228 725 2237
rect 777 2228 789 2237
rect 841 2228 853 2280
rect 905 2228 917 2280
rect 969 2228 981 2280
rect 1033 2271 1045 2280
rect 1097 2271 1109 2280
rect 1161 2271 1173 2280
rect 1225 2271 1237 2280
rect 1289 2271 1301 2280
rect 1353 2271 1365 2280
rect 1037 2237 1045 2271
rect 1289 2237 1291 2271
rect 1353 2237 1363 2271
rect 1033 2228 1045 2237
rect 1097 2228 1109 2237
rect 1161 2228 1173 2237
rect 1225 2228 1237 2237
rect 1289 2228 1301 2237
rect 1353 2228 1365 2237
rect 1417 2228 1429 2280
rect 1481 2228 1493 2280
rect 1545 2228 1557 2280
rect 1609 2271 1621 2280
rect 1673 2271 1685 2280
rect 1737 2271 1749 2280
rect 1801 2271 1813 2280
rect 1865 2271 1877 2280
rect 1929 2271 1996 2280
rect 1613 2237 1621 2271
rect 1865 2237 1867 2271
rect 1929 2237 1939 2271
rect 1973 2237 1996 2271
rect 1609 2228 1621 2237
rect 1673 2228 1685 2237
rect 1737 2228 1749 2237
rect 1801 2228 1813 2237
rect 1865 2228 1877 2237
rect 1929 2228 1996 2237
rect 271 2071 1996 2228
rect 2024 2109 2175 2308
rect 235 2040 1024 2041
rect 235 2031 326 2040
rect 235 1997 319 2031
rect 235 1988 326 1997
rect 378 1988 390 2040
rect 442 1988 454 2040
rect 506 1988 518 2040
rect 570 1988 582 2040
rect 634 2031 646 2040
rect 698 2031 710 2040
rect 762 2031 774 2040
rect 826 2031 838 2040
rect 890 2031 902 2040
rect 641 1997 646 2031
rect 890 1997 895 2031
rect 634 1988 646 1997
rect 698 1988 710 1997
rect 762 1988 774 1997
rect 826 1988 838 1997
rect 890 1988 902 1997
rect 954 1988 966 2040
rect 1018 1988 1024 2040
rect 235 1987 1024 1988
rect 235 1933 262 1987
rect 1052 1953 1216 2071
rect 2024 2041 2033 2109
rect 1244 2040 2033 2041
rect 1244 1988 1250 2040
rect 1302 1988 1314 2040
rect 1366 2031 1378 2040
rect 1430 2031 1442 2040
rect 1494 2031 1506 2040
rect 1558 2031 1570 2040
rect 1622 2031 1634 2040
rect 1373 1997 1378 2031
rect 1622 1997 1627 2031
rect 1366 1988 1378 1997
rect 1430 1988 1442 1997
rect 1494 1988 1506 1997
rect 1558 1988 1570 1997
rect 1622 1988 1634 1997
rect 1686 1988 1698 2040
rect 1750 1988 1762 2040
rect 1814 1988 1826 2040
rect 1878 1988 1890 2040
rect 1942 2031 2033 2040
rect 1949 1997 2033 2031
rect 1942 1988 2033 1997
rect 1244 1987 2033 1988
rect 256 1897 262 1933
rect 290 1933 1978 1953
rect 290 1925 1058 1933
rect 256 1881 1024 1897
rect 235 1869 1024 1881
rect 1052 1881 1058 1925
rect 1110 1881 1158 1933
rect 1210 1925 1978 1933
rect 2006 1933 2033 1987
rect 1210 1881 1216 1925
rect 2006 1897 2012 1933
rect 1052 1869 1216 1881
rect 1244 1881 2012 1897
rect 1244 1869 2033 1881
rect 256 1817 262 1869
rect 1052 1841 1058 1869
rect 235 1805 262 1817
rect 290 1817 1058 1841
rect 1110 1817 1158 1869
rect 1210 1841 1216 1869
rect 1210 1817 1978 1841
rect 290 1813 1978 1817
rect 2006 1817 2012 1869
rect 256 1785 262 1805
rect 1052 1805 1216 1813
rect 256 1757 1024 1785
rect 256 1753 262 1757
rect 235 1741 262 1753
rect 256 1689 262 1741
rect 1052 1753 1058 1805
rect 1110 1753 1158 1805
rect 1210 1753 1216 1805
rect 2006 1805 2033 1817
rect 2006 1785 2012 1805
rect 1244 1757 2012 1785
rect 1052 1741 1216 1753
rect 1052 1729 1058 1741
rect 290 1701 1058 1729
rect 235 1677 262 1689
rect 256 1673 262 1677
rect 1052 1689 1058 1701
rect 1110 1689 1158 1741
rect 1210 1729 1216 1741
rect 2006 1753 2012 1757
rect 2006 1741 2033 1753
rect 1210 1701 1978 1729
rect 1210 1689 1216 1701
rect 1052 1677 1216 1689
rect 256 1645 1024 1673
rect 256 1625 262 1645
rect 235 1613 262 1625
rect 1052 1625 1058 1677
rect 1110 1625 1158 1677
rect 1210 1625 1216 1677
rect 2006 1689 2012 1741
rect 2006 1677 2033 1689
rect 2006 1673 2012 1677
rect 1244 1645 2012 1673
rect 1052 1617 1216 1625
rect 2006 1625 2012 1645
rect 256 1561 262 1613
rect 290 1613 1978 1617
rect 290 1589 1058 1613
rect 1052 1561 1058 1589
rect 1110 1561 1158 1613
rect 1210 1589 1978 1613
rect 2006 1613 2033 1625
rect 1210 1561 1216 1589
rect 2006 1561 2012 1613
rect 235 1549 1024 1561
rect 256 1533 1024 1549
rect 1052 1549 1216 1561
rect 256 1497 262 1533
rect 1052 1505 1058 1549
rect 235 1485 262 1497
rect 256 1449 262 1485
rect 290 1497 1058 1505
rect 1110 1497 1158 1549
rect 1210 1505 1216 1549
rect 1244 1549 2033 1561
rect 1244 1533 2012 1549
rect 1210 1497 1978 1505
rect 290 1485 1978 1497
rect 290 1477 1058 1485
rect 256 1433 1024 1449
rect 235 1421 1024 1433
rect 1052 1433 1058 1477
rect 1110 1433 1158 1485
rect 1210 1477 1978 1485
rect 2006 1497 2012 1533
rect 2006 1485 2033 1497
rect 1210 1433 1216 1477
rect 2006 1449 2012 1485
rect 1052 1421 1216 1433
rect 1244 1433 2012 1449
rect 1244 1421 2033 1433
rect 256 1369 262 1421
rect 1052 1393 1058 1421
rect 235 1357 262 1369
rect 290 1369 1058 1393
rect 1110 1369 1158 1421
rect 1210 1393 1216 1421
rect 1210 1369 1978 1393
rect 290 1365 1978 1369
rect 2006 1369 2012 1421
rect 256 1337 262 1357
rect 1052 1357 1216 1365
rect 256 1309 1024 1337
rect 256 1305 262 1309
rect 235 1293 262 1305
rect 256 1241 262 1293
rect 1052 1305 1058 1357
rect 1110 1305 1158 1357
rect 1210 1305 1216 1357
rect 2006 1357 2033 1369
rect 2006 1337 2012 1357
rect 1244 1309 2012 1337
rect 1052 1293 1216 1305
rect 1052 1281 1058 1293
rect 290 1253 1058 1281
rect 235 1071 262 1241
rect 1052 1241 1058 1253
rect 1110 1241 1158 1293
rect 1210 1281 1216 1293
rect 2006 1305 2012 1309
rect 2006 1293 2033 1305
rect 1210 1253 1978 1281
rect 1210 1241 1216 1253
rect 1052 1219 1216 1241
rect 2006 1241 2012 1293
rect 290 1218 1978 1219
rect 290 1166 307 1218
rect 359 1209 371 1218
rect 423 1209 435 1218
rect 487 1209 499 1218
rect 551 1209 563 1218
rect 615 1209 627 1218
rect 679 1209 691 1218
rect 743 1209 755 1218
rect 807 1209 819 1218
rect 871 1209 883 1218
rect 935 1209 947 1218
rect 999 1209 1011 1218
rect 1063 1166 1205 1218
rect 1257 1209 1269 1218
rect 1321 1209 1333 1218
rect 1385 1209 1397 1218
rect 1449 1209 1461 1218
rect 1513 1209 1525 1218
rect 1577 1209 1589 1218
rect 1641 1209 1653 1218
rect 1705 1209 1717 1218
rect 1769 1209 1781 1218
rect 1833 1209 1845 1218
rect 1897 1209 1909 1218
rect 1961 1166 1978 1218
rect 290 1146 344 1166
rect 1026 1146 1242 1166
rect 1924 1146 1978 1166
rect 290 1094 307 1146
rect 359 1094 371 1103
rect 423 1094 435 1103
rect 487 1094 499 1103
rect 551 1094 563 1103
rect 615 1094 627 1103
rect 679 1094 691 1103
rect 743 1094 755 1103
rect 807 1094 819 1103
rect 871 1094 883 1103
rect 935 1094 947 1103
rect 999 1094 1011 1103
rect 1063 1094 1205 1146
rect 1257 1094 1269 1103
rect 1321 1094 1333 1103
rect 1385 1094 1397 1103
rect 1449 1094 1461 1103
rect 1513 1094 1525 1103
rect 1577 1094 1589 1103
rect 1641 1094 1653 1103
rect 1705 1094 1717 1103
rect 1769 1094 1781 1103
rect 1833 1094 1845 1103
rect 1897 1094 1909 1103
rect 1961 1094 1978 1146
rect 290 1093 1978 1094
rect 256 1019 262 1071
rect 1052 1071 1216 1093
rect 1052 1059 1058 1071
rect 290 1031 1058 1059
rect 235 1007 262 1019
rect 256 1003 262 1007
rect 1052 1019 1058 1031
rect 1110 1019 1158 1071
rect 1210 1059 1216 1071
rect 2006 1071 2033 1241
rect 1210 1031 1978 1059
rect 1210 1019 1216 1031
rect 1052 1007 1216 1019
rect 256 975 1024 1003
rect 256 955 262 975
rect 235 943 262 955
rect 1052 955 1058 1007
rect 1110 955 1158 1007
rect 1210 955 1216 1007
rect 2006 1019 2012 1071
rect 2006 1007 2033 1019
rect 2006 1003 2012 1007
rect 1244 975 2012 1003
rect 1052 947 1216 955
rect 2006 955 2012 975
rect 256 891 262 943
rect 290 943 1978 947
rect 290 919 1058 943
rect 1052 891 1058 919
rect 1110 891 1158 943
rect 1210 919 1978 943
rect 2006 943 2033 955
rect 1210 891 1216 919
rect 2006 891 2012 943
rect 235 879 1024 891
rect 256 863 1024 879
rect 1052 879 1216 891
rect 256 827 262 863
rect 1052 835 1058 879
rect 235 815 262 827
rect 256 779 262 815
rect 290 827 1058 835
rect 1110 827 1158 879
rect 1210 835 1216 879
rect 1244 879 2033 891
rect 1244 863 2012 879
rect 1210 827 1978 835
rect 290 815 1978 827
rect 290 807 1058 815
rect 256 763 1024 779
rect 235 751 1024 763
rect 1052 763 1058 807
rect 1110 763 1158 815
rect 1210 807 1978 815
rect 2006 827 2012 863
rect 2006 815 2033 827
rect 1210 763 1216 807
rect 2006 779 2012 815
rect 1052 751 1216 763
rect 1244 763 2012 779
rect 1244 751 2033 763
rect 256 699 262 751
rect 1052 723 1058 751
rect 235 687 262 699
rect 290 699 1058 723
rect 1110 699 1158 751
rect 1210 723 1216 751
rect 1210 699 1978 723
rect 290 695 1978 699
rect 2006 699 2012 751
rect 256 667 262 687
rect 1052 687 1216 695
rect 256 639 1024 667
rect 256 635 262 639
rect 235 623 262 635
rect 256 571 262 623
rect 1052 635 1058 687
rect 1110 635 1158 687
rect 1210 635 1216 687
rect 2006 687 2033 699
rect 2006 667 2012 687
rect 1244 639 2012 667
rect 1052 623 1216 635
rect 1052 611 1058 623
rect 290 583 1058 611
rect 235 559 262 571
rect 256 555 262 559
rect 1052 571 1058 583
rect 1110 571 1158 623
rect 1210 611 1216 623
rect 2006 635 2012 639
rect 2006 623 2033 635
rect 1210 583 1978 611
rect 1210 571 1216 583
rect 1052 559 1216 571
rect 256 527 1024 555
rect 256 507 262 527
rect 235 495 262 507
rect 1052 507 1058 559
rect 1110 507 1158 559
rect 1210 507 1216 559
rect 2006 571 2012 623
rect 2006 559 2033 571
rect 2006 555 2012 559
rect 1244 527 2012 555
rect 1052 499 1216 507
rect 2006 507 2012 527
rect 256 443 262 495
rect 290 495 1978 499
rect 290 471 1058 495
rect 1052 443 1058 471
rect 1110 443 1158 495
rect 1210 471 1978 495
rect 2006 495 2033 507
rect 1210 443 1216 471
rect 2006 443 2012 495
rect 235 431 1024 443
rect 256 415 1024 431
rect 1052 431 1216 443
rect 256 379 262 415
rect 1052 387 1058 431
rect 235 325 262 379
rect 290 379 1058 387
rect 1110 379 1158 431
rect 1210 387 1216 431
rect 1244 431 2033 443
rect 1244 415 2012 431
rect 1210 379 1978 387
rect 290 359 1978 379
rect 2006 379 2012 415
rect 235 324 1024 325
rect 235 315 326 324
rect 235 281 319 315
rect 235 272 326 281
rect 378 272 390 324
rect 442 272 454 324
rect 506 272 518 324
rect 570 272 582 324
rect 634 315 646 324
rect 698 315 710 324
rect 762 315 774 324
rect 826 315 838 324
rect 890 315 902 324
rect 641 281 646 315
rect 890 281 895 315
rect 634 272 646 281
rect 698 272 710 281
rect 762 272 774 281
rect 826 272 838 281
rect 890 272 902 281
rect 954 272 966 324
rect 1018 272 1024 324
rect 235 271 1024 272
rect 235 203 243 271
rect 1052 241 1216 359
rect 2006 325 2033 379
rect 1244 324 2033 325
rect 1244 272 1250 324
rect 1302 272 1314 324
rect 1366 315 1378 324
rect 1430 315 1442 324
rect 1494 315 1506 324
rect 1558 315 1570 324
rect 1622 315 1634 324
rect 1373 281 1378 315
rect 1622 281 1627 315
rect 1366 272 1378 281
rect 1430 272 1442 281
rect 1494 272 1506 281
rect 1558 272 1570 281
rect 1622 272 1634 281
rect 1686 272 1698 324
rect 1750 272 1762 324
rect 1814 272 1826 324
rect 1878 272 1890 324
rect 1942 315 2033 324
rect 1949 281 2033 315
rect 1942 272 2033 281
rect 1244 271 2033 272
rect 93 30 243 203
rect 271 110 1996 241
rect 271 58 277 110
rect 329 58 341 110
rect 393 58 405 110
rect 457 101 469 110
rect 521 101 533 110
rect 585 101 597 110
rect 649 101 661 110
rect 713 101 725 110
rect 777 101 789 110
rect 461 67 469 101
rect 713 67 715 101
rect 777 67 787 101
rect 457 58 469 67
rect 521 58 533 67
rect 585 58 597 67
rect 649 58 661 67
rect 713 58 725 67
rect 777 58 789 67
rect 841 58 853 110
rect 905 58 917 110
rect 969 58 981 110
rect 1033 101 1045 110
rect 1097 101 1109 110
rect 1161 101 1173 110
rect 1225 101 1237 110
rect 1289 101 1301 110
rect 1353 101 1365 110
rect 1037 67 1045 101
rect 1289 67 1291 101
rect 1353 67 1363 101
rect 1033 58 1045 67
rect 1097 58 1109 67
rect 1161 58 1173 67
rect 1225 58 1237 67
rect 1289 58 1301 67
rect 1353 58 1365 67
rect 1417 58 1429 110
rect 1481 58 1493 110
rect 1545 58 1557 110
rect 1609 101 1621 110
rect 1673 101 1685 110
rect 1737 101 1749 110
rect 1801 101 1813 110
rect 1865 101 1877 110
rect 1929 101 1996 110
rect 1613 67 1621 101
rect 1865 67 1867 101
rect 1929 67 1939 101
rect 1973 67 1996 101
rect 1609 58 1621 67
rect 1673 58 1685 67
rect 1737 58 1749 67
rect 1801 58 1813 67
rect 1865 58 1877 67
rect 1929 58 1996 67
rect 2024 203 2033 271
rect 2139 203 2175 2109
rect 2024 30 2175 203
rect 93 0 2175 30
<< via1 >>
rect 277 2271 329 2280
rect 277 2237 283 2271
rect 283 2237 317 2271
rect 317 2237 329 2271
rect 277 2228 329 2237
rect 341 2271 393 2280
rect 341 2237 355 2271
rect 355 2237 389 2271
rect 389 2237 393 2271
rect 341 2228 393 2237
rect 405 2271 457 2280
rect 469 2271 521 2280
rect 533 2271 585 2280
rect 597 2271 649 2280
rect 661 2271 713 2280
rect 725 2271 777 2280
rect 789 2271 841 2280
rect 405 2237 427 2271
rect 427 2237 457 2271
rect 469 2237 499 2271
rect 499 2237 521 2271
rect 533 2237 571 2271
rect 571 2237 585 2271
rect 597 2237 605 2271
rect 605 2237 643 2271
rect 643 2237 649 2271
rect 661 2237 677 2271
rect 677 2237 713 2271
rect 725 2237 749 2271
rect 749 2237 777 2271
rect 789 2237 821 2271
rect 821 2237 841 2271
rect 405 2228 457 2237
rect 469 2228 521 2237
rect 533 2228 585 2237
rect 597 2228 649 2237
rect 661 2228 713 2237
rect 725 2228 777 2237
rect 789 2228 841 2237
rect 853 2271 905 2280
rect 853 2237 859 2271
rect 859 2237 893 2271
rect 893 2237 905 2271
rect 853 2228 905 2237
rect 917 2271 969 2280
rect 917 2237 931 2271
rect 931 2237 965 2271
rect 965 2237 969 2271
rect 917 2228 969 2237
rect 981 2271 1033 2280
rect 1045 2271 1097 2280
rect 1109 2271 1161 2280
rect 1173 2271 1225 2280
rect 1237 2271 1289 2280
rect 1301 2271 1353 2280
rect 1365 2271 1417 2280
rect 981 2237 1003 2271
rect 1003 2237 1033 2271
rect 1045 2237 1075 2271
rect 1075 2237 1097 2271
rect 1109 2237 1147 2271
rect 1147 2237 1161 2271
rect 1173 2237 1181 2271
rect 1181 2237 1219 2271
rect 1219 2237 1225 2271
rect 1237 2237 1253 2271
rect 1253 2237 1289 2271
rect 1301 2237 1325 2271
rect 1325 2237 1353 2271
rect 1365 2237 1397 2271
rect 1397 2237 1417 2271
rect 981 2228 1033 2237
rect 1045 2228 1097 2237
rect 1109 2228 1161 2237
rect 1173 2228 1225 2237
rect 1237 2228 1289 2237
rect 1301 2228 1353 2237
rect 1365 2228 1417 2237
rect 1429 2271 1481 2280
rect 1429 2237 1435 2271
rect 1435 2237 1469 2271
rect 1469 2237 1481 2271
rect 1429 2228 1481 2237
rect 1493 2271 1545 2280
rect 1493 2237 1507 2271
rect 1507 2237 1541 2271
rect 1541 2237 1545 2271
rect 1493 2228 1545 2237
rect 1557 2271 1609 2280
rect 1621 2271 1673 2280
rect 1685 2271 1737 2280
rect 1749 2271 1801 2280
rect 1813 2271 1865 2280
rect 1877 2271 1929 2280
rect 1557 2237 1579 2271
rect 1579 2237 1609 2271
rect 1621 2237 1651 2271
rect 1651 2237 1673 2271
rect 1685 2237 1723 2271
rect 1723 2237 1737 2271
rect 1749 2237 1757 2271
rect 1757 2237 1795 2271
rect 1795 2237 1801 2271
rect 1813 2237 1829 2271
rect 1829 2237 1865 2271
rect 1877 2237 1901 2271
rect 1901 2237 1929 2271
rect 1557 2228 1609 2237
rect 1621 2228 1673 2237
rect 1685 2228 1737 2237
rect 1749 2228 1801 2237
rect 1813 2228 1865 2237
rect 1877 2228 1929 2237
rect 326 2031 378 2040
rect 326 1997 353 2031
rect 353 1997 378 2031
rect 326 1988 378 1997
rect 390 2031 442 2040
rect 390 1997 391 2031
rect 391 1997 425 2031
rect 425 1997 442 2031
rect 390 1988 442 1997
rect 454 2031 506 2040
rect 454 1997 463 2031
rect 463 1997 497 2031
rect 497 1997 506 2031
rect 454 1988 506 1997
rect 518 2031 570 2040
rect 518 1997 535 2031
rect 535 1997 569 2031
rect 569 1997 570 2031
rect 518 1988 570 1997
rect 582 2031 634 2040
rect 646 2031 698 2040
rect 710 2031 762 2040
rect 774 2031 826 2040
rect 838 2031 890 2040
rect 902 2031 954 2040
rect 582 1997 607 2031
rect 607 1997 634 2031
rect 646 1997 679 2031
rect 679 1997 698 2031
rect 710 1997 713 2031
rect 713 1997 751 2031
rect 751 1997 762 2031
rect 774 1997 785 2031
rect 785 1997 823 2031
rect 823 1997 826 2031
rect 838 1997 857 2031
rect 857 1997 890 2031
rect 902 1997 929 2031
rect 929 1997 954 2031
rect 582 1988 634 1997
rect 646 1988 698 1997
rect 710 1988 762 1997
rect 774 1988 826 1997
rect 838 1988 890 1997
rect 902 1988 954 1997
rect 966 2031 1018 2040
rect 966 1997 967 2031
rect 967 1997 1001 2031
rect 1001 1997 1018 2031
rect 966 1988 1018 1997
rect 1250 2031 1302 2040
rect 1250 1997 1267 2031
rect 1267 1997 1301 2031
rect 1301 1997 1302 2031
rect 1250 1988 1302 1997
rect 1314 2031 1366 2040
rect 1378 2031 1430 2040
rect 1442 2031 1494 2040
rect 1506 2031 1558 2040
rect 1570 2031 1622 2040
rect 1634 2031 1686 2040
rect 1314 1997 1339 2031
rect 1339 1997 1366 2031
rect 1378 1997 1411 2031
rect 1411 1997 1430 2031
rect 1442 1997 1445 2031
rect 1445 1997 1483 2031
rect 1483 1997 1494 2031
rect 1506 1997 1517 2031
rect 1517 1997 1555 2031
rect 1555 1997 1558 2031
rect 1570 1997 1589 2031
rect 1589 1997 1622 2031
rect 1634 1997 1661 2031
rect 1661 1997 1686 2031
rect 1314 1988 1366 1997
rect 1378 1988 1430 1997
rect 1442 1988 1494 1997
rect 1506 1988 1558 1997
rect 1570 1988 1622 1997
rect 1634 1988 1686 1997
rect 1698 2031 1750 2040
rect 1698 1997 1699 2031
rect 1699 1997 1733 2031
rect 1733 1997 1750 2031
rect 1698 1988 1750 1997
rect 1762 2031 1814 2040
rect 1762 1997 1771 2031
rect 1771 1997 1805 2031
rect 1805 1997 1814 2031
rect 1762 1988 1814 1997
rect 1826 2031 1878 2040
rect 1826 1997 1843 2031
rect 1843 1997 1877 2031
rect 1877 1997 1878 2031
rect 1826 1988 1878 1997
rect 1890 2031 1942 2040
rect 1890 1997 1915 2031
rect 1915 1997 1942 2031
rect 1890 1988 1942 1997
rect 204 1881 235 1933
rect 235 1881 256 1933
rect 1058 1881 1110 1933
rect 1158 1881 1210 1933
rect 2012 1881 2033 1933
rect 2033 1881 2064 1933
rect 204 1817 235 1869
rect 235 1817 256 1869
rect 1058 1817 1110 1869
rect 1158 1817 1210 1869
rect 2012 1817 2033 1869
rect 2033 1817 2064 1869
rect 204 1753 235 1805
rect 235 1753 256 1805
rect 204 1689 235 1741
rect 235 1689 256 1741
rect 1058 1753 1110 1805
rect 1158 1753 1210 1805
rect 204 1625 235 1677
rect 235 1625 256 1677
rect 1058 1689 1110 1741
rect 1158 1689 1210 1741
rect 2012 1753 2033 1805
rect 2033 1753 2064 1805
rect 1058 1625 1110 1677
rect 1158 1625 1210 1677
rect 2012 1689 2033 1741
rect 2033 1689 2064 1741
rect 2012 1625 2033 1677
rect 2033 1625 2064 1677
rect 204 1561 235 1613
rect 235 1561 256 1613
rect 1058 1561 1110 1613
rect 1158 1561 1210 1613
rect 2012 1561 2033 1613
rect 2033 1561 2064 1613
rect 204 1497 235 1549
rect 235 1497 256 1549
rect 204 1433 235 1485
rect 235 1433 256 1485
rect 1058 1497 1110 1549
rect 1158 1497 1210 1549
rect 1058 1433 1110 1485
rect 1158 1433 1210 1485
rect 2012 1497 2033 1549
rect 2033 1497 2064 1549
rect 2012 1433 2033 1485
rect 2033 1433 2064 1485
rect 204 1369 235 1421
rect 235 1369 256 1421
rect 1058 1369 1110 1421
rect 1158 1369 1210 1421
rect 2012 1369 2033 1421
rect 2033 1369 2064 1421
rect 204 1305 235 1357
rect 235 1305 256 1357
rect 204 1241 235 1293
rect 235 1241 256 1293
rect 1058 1305 1110 1357
rect 1158 1305 1210 1357
rect 1058 1241 1110 1293
rect 1158 1241 1210 1293
rect 2012 1305 2033 1357
rect 2033 1305 2064 1357
rect 2012 1241 2033 1293
rect 2033 1241 2064 1293
rect 307 1209 359 1218
rect 371 1209 423 1218
rect 435 1209 487 1218
rect 499 1209 551 1218
rect 563 1209 615 1218
rect 627 1209 679 1218
rect 691 1209 743 1218
rect 755 1209 807 1218
rect 819 1209 871 1218
rect 883 1209 935 1218
rect 947 1209 999 1218
rect 1011 1209 1063 1218
rect 307 1166 344 1209
rect 344 1166 359 1209
rect 371 1166 423 1209
rect 435 1166 487 1209
rect 499 1166 551 1209
rect 563 1166 615 1209
rect 627 1166 679 1209
rect 691 1166 743 1209
rect 755 1166 807 1209
rect 819 1166 871 1209
rect 883 1166 935 1209
rect 947 1166 999 1209
rect 1011 1166 1026 1209
rect 1026 1166 1063 1209
rect 1205 1209 1257 1218
rect 1269 1209 1321 1218
rect 1333 1209 1385 1218
rect 1397 1209 1449 1218
rect 1461 1209 1513 1218
rect 1525 1209 1577 1218
rect 1589 1209 1641 1218
rect 1653 1209 1705 1218
rect 1717 1209 1769 1218
rect 1781 1209 1833 1218
rect 1845 1209 1897 1218
rect 1909 1209 1961 1218
rect 1205 1166 1242 1209
rect 1242 1166 1257 1209
rect 1269 1166 1321 1209
rect 1333 1166 1385 1209
rect 1397 1166 1449 1209
rect 1461 1166 1513 1209
rect 1525 1166 1577 1209
rect 1589 1166 1641 1209
rect 1653 1166 1705 1209
rect 1717 1166 1769 1209
rect 1781 1166 1833 1209
rect 1845 1166 1897 1209
rect 1909 1166 1924 1209
rect 1924 1166 1961 1209
rect 307 1103 344 1146
rect 344 1103 359 1146
rect 371 1103 423 1146
rect 435 1103 487 1146
rect 499 1103 551 1146
rect 563 1103 615 1146
rect 627 1103 679 1146
rect 691 1103 743 1146
rect 755 1103 807 1146
rect 819 1103 871 1146
rect 883 1103 935 1146
rect 947 1103 999 1146
rect 1011 1103 1026 1146
rect 1026 1103 1063 1146
rect 307 1094 359 1103
rect 371 1094 423 1103
rect 435 1094 487 1103
rect 499 1094 551 1103
rect 563 1094 615 1103
rect 627 1094 679 1103
rect 691 1094 743 1103
rect 755 1094 807 1103
rect 819 1094 871 1103
rect 883 1094 935 1103
rect 947 1094 999 1103
rect 1011 1094 1063 1103
rect 1205 1103 1242 1146
rect 1242 1103 1257 1146
rect 1269 1103 1321 1146
rect 1333 1103 1385 1146
rect 1397 1103 1449 1146
rect 1461 1103 1513 1146
rect 1525 1103 1577 1146
rect 1589 1103 1641 1146
rect 1653 1103 1705 1146
rect 1717 1103 1769 1146
rect 1781 1103 1833 1146
rect 1845 1103 1897 1146
rect 1909 1103 1924 1146
rect 1924 1103 1961 1146
rect 1205 1094 1257 1103
rect 1269 1094 1321 1103
rect 1333 1094 1385 1103
rect 1397 1094 1449 1103
rect 1461 1094 1513 1103
rect 1525 1094 1577 1103
rect 1589 1094 1641 1103
rect 1653 1094 1705 1103
rect 1717 1094 1769 1103
rect 1781 1094 1833 1103
rect 1845 1094 1897 1103
rect 1909 1094 1961 1103
rect 204 1019 235 1071
rect 235 1019 256 1071
rect 204 955 235 1007
rect 235 955 256 1007
rect 1058 1019 1110 1071
rect 1158 1019 1210 1071
rect 1058 955 1110 1007
rect 1158 955 1210 1007
rect 2012 1019 2033 1071
rect 2033 1019 2064 1071
rect 2012 955 2033 1007
rect 2033 955 2064 1007
rect 204 891 235 943
rect 235 891 256 943
rect 1058 891 1110 943
rect 1158 891 1210 943
rect 2012 891 2033 943
rect 2033 891 2064 943
rect 204 827 235 879
rect 235 827 256 879
rect 204 763 235 815
rect 235 763 256 815
rect 1058 827 1110 879
rect 1158 827 1210 879
rect 1058 763 1110 815
rect 1158 763 1210 815
rect 2012 827 2033 879
rect 2033 827 2064 879
rect 2012 763 2033 815
rect 2033 763 2064 815
rect 204 699 235 751
rect 235 699 256 751
rect 1058 699 1110 751
rect 1158 699 1210 751
rect 2012 699 2033 751
rect 2033 699 2064 751
rect 204 635 235 687
rect 235 635 256 687
rect 204 571 235 623
rect 235 571 256 623
rect 1058 635 1110 687
rect 1158 635 1210 687
rect 204 507 235 559
rect 235 507 256 559
rect 1058 571 1110 623
rect 1158 571 1210 623
rect 2012 635 2033 687
rect 2033 635 2064 687
rect 1058 507 1110 559
rect 1158 507 1210 559
rect 2012 571 2033 623
rect 2033 571 2064 623
rect 2012 507 2033 559
rect 2033 507 2064 559
rect 204 443 235 495
rect 235 443 256 495
rect 1058 443 1110 495
rect 1158 443 1210 495
rect 2012 443 2033 495
rect 2033 443 2064 495
rect 204 379 235 431
rect 235 379 256 431
rect 1058 379 1110 431
rect 1158 379 1210 431
rect 2012 379 2033 431
rect 2033 379 2064 431
rect 326 315 378 324
rect 326 281 353 315
rect 353 281 378 315
rect 326 272 378 281
rect 390 315 442 324
rect 390 281 391 315
rect 391 281 425 315
rect 425 281 442 315
rect 390 272 442 281
rect 454 315 506 324
rect 454 281 463 315
rect 463 281 497 315
rect 497 281 506 315
rect 454 272 506 281
rect 518 315 570 324
rect 518 281 535 315
rect 535 281 569 315
rect 569 281 570 315
rect 518 272 570 281
rect 582 315 634 324
rect 646 315 698 324
rect 710 315 762 324
rect 774 315 826 324
rect 838 315 890 324
rect 902 315 954 324
rect 582 281 607 315
rect 607 281 634 315
rect 646 281 679 315
rect 679 281 698 315
rect 710 281 713 315
rect 713 281 751 315
rect 751 281 762 315
rect 774 281 785 315
rect 785 281 823 315
rect 823 281 826 315
rect 838 281 857 315
rect 857 281 890 315
rect 902 281 929 315
rect 929 281 954 315
rect 582 272 634 281
rect 646 272 698 281
rect 710 272 762 281
rect 774 272 826 281
rect 838 272 890 281
rect 902 272 954 281
rect 966 315 1018 324
rect 966 281 967 315
rect 967 281 1001 315
rect 1001 281 1018 315
rect 966 272 1018 281
rect 1250 315 1302 324
rect 1250 281 1267 315
rect 1267 281 1301 315
rect 1301 281 1302 315
rect 1250 272 1302 281
rect 1314 315 1366 324
rect 1378 315 1430 324
rect 1442 315 1494 324
rect 1506 315 1558 324
rect 1570 315 1622 324
rect 1634 315 1686 324
rect 1314 281 1339 315
rect 1339 281 1366 315
rect 1378 281 1411 315
rect 1411 281 1430 315
rect 1442 281 1445 315
rect 1445 281 1483 315
rect 1483 281 1494 315
rect 1506 281 1517 315
rect 1517 281 1555 315
rect 1555 281 1558 315
rect 1570 281 1589 315
rect 1589 281 1622 315
rect 1634 281 1661 315
rect 1661 281 1686 315
rect 1314 272 1366 281
rect 1378 272 1430 281
rect 1442 272 1494 281
rect 1506 272 1558 281
rect 1570 272 1622 281
rect 1634 272 1686 281
rect 1698 315 1750 324
rect 1698 281 1699 315
rect 1699 281 1733 315
rect 1733 281 1750 315
rect 1698 272 1750 281
rect 1762 315 1814 324
rect 1762 281 1771 315
rect 1771 281 1805 315
rect 1805 281 1814 315
rect 1762 272 1814 281
rect 1826 315 1878 324
rect 1826 281 1843 315
rect 1843 281 1877 315
rect 1877 281 1878 315
rect 1826 272 1878 281
rect 1890 315 1942 324
rect 1890 281 1915 315
rect 1915 281 1942 315
rect 1890 272 1942 281
rect 277 101 329 110
rect 277 67 283 101
rect 283 67 317 101
rect 317 67 329 101
rect 277 58 329 67
rect 341 101 393 110
rect 341 67 355 101
rect 355 67 389 101
rect 389 67 393 101
rect 341 58 393 67
rect 405 101 457 110
rect 469 101 521 110
rect 533 101 585 110
rect 597 101 649 110
rect 661 101 713 110
rect 725 101 777 110
rect 789 101 841 110
rect 405 67 427 101
rect 427 67 457 101
rect 469 67 499 101
rect 499 67 521 101
rect 533 67 571 101
rect 571 67 585 101
rect 597 67 605 101
rect 605 67 643 101
rect 643 67 649 101
rect 661 67 677 101
rect 677 67 713 101
rect 725 67 749 101
rect 749 67 777 101
rect 789 67 821 101
rect 821 67 841 101
rect 405 58 457 67
rect 469 58 521 67
rect 533 58 585 67
rect 597 58 649 67
rect 661 58 713 67
rect 725 58 777 67
rect 789 58 841 67
rect 853 101 905 110
rect 853 67 859 101
rect 859 67 893 101
rect 893 67 905 101
rect 853 58 905 67
rect 917 101 969 110
rect 917 67 931 101
rect 931 67 965 101
rect 965 67 969 101
rect 917 58 969 67
rect 981 101 1033 110
rect 1045 101 1097 110
rect 1109 101 1161 110
rect 1173 101 1225 110
rect 1237 101 1289 110
rect 1301 101 1353 110
rect 1365 101 1417 110
rect 981 67 1003 101
rect 1003 67 1033 101
rect 1045 67 1075 101
rect 1075 67 1097 101
rect 1109 67 1147 101
rect 1147 67 1161 101
rect 1173 67 1181 101
rect 1181 67 1219 101
rect 1219 67 1225 101
rect 1237 67 1253 101
rect 1253 67 1289 101
rect 1301 67 1325 101
rect 1325 67 1353 101
rect 1365 67 1397 101
rect 1397 67 1417 101
rect 981 58 1033 67
rect 1045 58 1097 67
rect 1109 58 1161 67
rect 1173 58 1225 67
rect 1237 58 1289 67
rect 1301 58 1353 67
rect 1365 58 1417 67
rect 1429 101 1481 110
rect 1429 67 1435 101
rect 1435 67 1469 101
rect 1469 67 1481 101
rect 1429 58 1481 67
rect 1493 101 1545 110
rect 1493 67 1507 101
rect 1507 67 1541 101
rect 1541 67 1545 101
rect 1493 58 1545 67
rect 1557 101 1609 110
rect 1621 101 1673 110
rect 1685 101 1737 110
rect 1749 101 1801 110
rect 1813 101 1865 110
rect 1877 101 1929 110
rect 1557 67 1579 101
rect 1579 67 1609 101
rect 1621 67 1651 101
rect 1651 67 1673 101
rect 1685 67 1723 101
rect 1723 67 1737 101
rect 1749 67 1757 101
rect 1757 67 1795 101
rect 1795 67 1801 101
rect 1813 67 1829 101
rect 1829 67 1865 101
rect 1877 67 1901 101
rect 1901 67 1929 101
rect 1557 58 1609 67
rect 1621 58 1673 67
rect 1685 58 1737 67
rect 1749 58 1801 67
rect 1813 58 1865 67
rect 1877 58 1929 67
<< metal2 >>
rect 65 2300 2203 2323
rect 121 2280 2147 2300
rect 121 2244 277 2280
rect 65 2228 277 2244
rect 329 2228 341 2280
rect 393 2228 405 2280
rect 457 2228 469 2280
rect 521 2228 533 2280
rect 585 2228 597 2280
rect 649 2228 661 2280
rect 713 2228 725 2280
rect 777 2228 789 2280
rect 841 2228 853 2280
rect 905 2228 917 2280
rect 969 2228 981 2280
rect 1033 2228 1045 2280
rect 1097 2228 1109 2280
rect 1161 2228 1173 2280
rect 1225 2228 1237 2280
rect 1289 2228 1301 2280
rect 1353 2228 1365 2280
rect 1417 2228 1429 2280
rect 1481 2228 1493 2280
rect 1545 2228 1557 2280
rect 1609 2228 1621 2280
rect 1673 2228 1685 2280
rect 1737 2228 1749 2280
rect 1801 2228 1813 2280
rect 1865 2228 1877 2280
rect 1929 2244 2147 2280
rect 1929 2228 2203 2244
rect 65 2220 2203 2228
rect 121 2164 2147 2220
rect 65 2141 2203 2164
rect 65 2140 1106 2141
rect 121 2085 1106 2140
rect 1162 2140 2203 2141
rect 1162 2085 2147 2140
rect 121 2084 2147 2085
rect 65 2071 2203 2084
rect 65 2060 169 2071
rect 121 2004 169 2060
rect 1052 2061 1216 2071
rect 65 1980 169 2004
rect 121 1924 169 1980
rect 65 1900 169 1924
rect 121 1844 169 1900
rect 65 1820 169 1844
rect 121 1764 169 1820
rect 65 1740 169 1764
rect 121 1684 169 1740
rect 65 1660 169 1684
rect 121 1604 169 1660
rect 65 1580 169 1604
rect 121 1524 169 1580
rect 65 1500 169 1524
rect 121 1444 169 1500
rect 65 1420 169 1444
rect 121 1364 169 1420
rect 65 1340 169 1364
rect 121 1284 169 1340
rect 65 1260 169 1284
rect 121 1204 169 1260
rect 65 1180 169 1204
rect 121 1124 169 1180
rect 65 1100 169 1124
rect 121 1044 169 1100
rect 65 1020 169 1044
rect 121 964 169 1020
rect 65 940 169 964
rect 121 884 169 940
rect 65 860 169 884
rect 121 804 169 860
rect 65 780 169 804
rect 121 724 169 780
rect 65 700 169 724
rect 121 644 169 700
rect 65 620 169 644
rect 121 564 169 620
rect 65 540 169 564
rect 121 484 169 540
rect 65 460 169 484
rect 121 404 169 460
rect 65 380 169 404
rect 121 324 169 380
rect 65 300 169 324
rect 121 244 169 300
rect 198 2040 1024 2041
rect 198 2021 326 2040
rect 254 1988 326 2021
rect 378 1988 390 2040
rect 442 1988 454 2040
rect 506 1988 518 2040
rect 570 1988 582 2040
rect 634 1988 646 2040
rect 698 1988 710 2040
rect 762 1988 774 2040
rect 826 1988 838 2040
rect 890 1988 902 2040
rect 954 1988 966 2040
rect 1018 1988 1024 2040
rect 254 1987 1024 1988
rect 1052 2005 1106 2061
rect 1162 2005 1216 2061
rect 2098 2060 2203 2071
rect 254 1965 262 1987
rect 198 1953 262 1965
rect 1052 1981 1216 2005
rect 1244 2040 2070 2041
rect 1244 1988 1250 2040
rect 1302 1988 1314 2040
rect 1366 1988 1378 2040
rect 1430 1988 1442 2040
rect 1494 1988 1506 2040
rect 1558 1988 1570 2040
rect 1622 1988 1634 2040
rect 1686 1988 1698 2040
rect 1750 1988 1762 2040
rect 1814 1988 1826 2040
rect 1878 1988 1890 2040
rect 1942 2021 2070 2040
rect 1942 1988 2014 2021
rect 1244 1987 2014 1988
rect 198 1941 1024 1953
rect 254 1933 1024 1941
rect 256 1925 1024 1933
rect 1052 1933 1106 1981
rect 1162 1933 1216 1981
rect 2006 1965 2014 1987
rect 2006 1953 2070 1965
rect 198 1881 204 1885
rect 256 1881 262 1925
rect 1052 1897 1058 1933
rect 1110 1901 1158 1925
rect 198 1869 262 1881
rect 290 1881 1058 1897
rect 1210 1897 1216 1933
rect 1244 1941 2070 1953
rect 1244 1933 2014 1941
rect 1244 1925 2012 1933
rect 1210 1881 1978 1897
rect 290 1869 1106 1881
rect 1162 1869 1978 1881
rect 2006 1881 2012 1925
rect 2064 1881 2070 1885
rect 2006 1869 2070 1881
rect 198 1861 204 1869
rect 256 1841 262 1869
rect 256 1817 1024 1841
rect 254 1813 1024 1817
rect 1052 1817 1058 1869
rect 1110 1821 1158 1845
rect 1210 1817 1216 1869
rect 2006 1841 2012 1869
rect 2064 1861 2070 1869
rect 254 1805 262 1813
rect 198 1781 204 1805
rect 256 1753 262 1805
rect 1052 1805 1106 1817
rect 1162 1805 1216 1817
rect 1244 1817 2012 1841
rect 1244 1813 2014 1817
rect 1052 1785 1058 1805
rect 290 1757 1058 1785
rect 1210 1785 1216 1805
rect 2006 1805 2014 1813
rect 254 1741 262 1753
rect 256 1729 262 1741
rect 1052 1753 1058 1757
rect 1110 1753 1158 1765
rect 1210 1757 1978 1785
rect 1210 1753 1216 1757
rect 1052 1741 1216 1753
rect 198 1701 204 1725
rect 256 1701 1024 1729
rect 256 1689 262 1701
rect 254 1677 262 1689
rect 198 1625 204 1645
rect 256 1625 262 1677
rect 1052 1689 1058 1741
rect 1210 1689 1216 1741
rect 2006 1753 2012 1805
rect 2064 1781 2070 1805
rect 2006 1741 2014 1753
rect 2006 1729 2012 1741
rect 1244 1701 2012 1729
rect 2064 1701 2070 1725
rect 1052 1685 1106 1689
rect 1162 1685 1216 1689
rect 1052 1677 1216 1685
rect 1052 1673 1058 1677
rect 290 1645 1058 1673
rect 1110 1661 1158 1677
rect 1210 1673 1216 1677
rect 2006 1689 2012 1701
rect 2006 1677 2014 1689
rect 198 1621 262 1625
rect 254 1617 262 1621
rect 1052 1625 1058 1645
rect 1210 1645 1978 1673
rect 1210 1625 1216 1645
rect 254 1613 1024 1617
rect 256 1589 1024 1613
rect 1052 1613 1106 1625
rect 1162 1613 1216 1625
rect 2006 1625 2012 1677
rect 2064 1625 2070 1645
rect 2006 1621 2070 1625
rect 2006 1617 2014 1621
rect 198 1561 204 1565
rect 256 1561 262 1589
rect 1052 1561 1058 1613
rect 1110 1581 1158 1605
rect 1210 1561 1216 1613
rect 1244 1613 2014 1617
rect 1244 1589 2012 1613
rect 2006 1561 2012 1589
rect 2064 1561 2070 1565
rect 198 1549 262 1561
rect 198 1541 204 1549
rect 256 1505 262 1549
rect 290 1549 1106 1561
rect 1162 1549 1978 1561
rect 290 1533 1058 1549
rect 256 1497 1024 1505
rect 254 1485 1024 1497
rect 198 1461 204 1485
rect 256 1477 1024 1485
rect 1052 1497 1058 1533
rect 1210 1533 1978 1549
rect 2006 1549 2070 1561
rect 1110 1501 1158 1525
rect 1210 1497 1216 1533
rect 2006 1505 2012 1549
rect 2064 1541 2070 1549
rect 1052 1485 1106 1497
rect 1162 1485 1216 1497
rect 256 1433 262 1477
rect 1052 1449 1058 1485
rect 254 1421 262 1433
rect 290 1433 1058 1449
rect 1210 1449 1216 1485
rect 1244 1497 2012 1505
rect 1244 1485 2014 1497
rect 1244 1477 2012 1485
rect 1110 1433 1158 1445
rect 1210 1433 1978 1449
rect 290 1421 1978 1433
rect 2006 1433 2012 1477
rect 2064 1461 2070 1485
rect 2006 1421 2014 1433
rect 198 1381 204 1405
rect 256 1393 262 1421
rect 256 1369 1024 1393
rect 254 1365 1024 1369
rect 1052 1369 1058 1421
rect 1210 1369 1216 1421
rect 2006 1393 2012 1421
rect 1052 1365 1106 1369
rect 1162 1365 1216 1369
rect 1244 1369 2012 1393
rect 2064 1381 2070 1405
rect 1244 1365 2014 1369
rect 254 1357 262 1365
rect 198 1305 204 1325
rect 256 1305 262 1357
rect 1052 1357 1216 1365
rect 1052 1337 1058 1357
rect 1110 1341 1158 1357
rect 290 1309 1058 1337
rect 198 1301 262 1305
rect 254 1293 262 1301
rect 256 1281 262 1293
rect 1052 1305 1058 1309
rect 1210 1337 1216 1357
rect 2006 1357 2014 1365
rect 1210 1309 1978 1337
rect 1210 1305 1216 1309
rect 1052 1293 1106 1305
rect 1162 1293 1216 1305
rect 256 1253 1024 1281
rect 198 1241 204 1245
rect 256 1241 262 1253
rect 198 1221 262 1241
rect 254 1165 262 1221
rect 1052 1241 1058 1293
rect 1110 1261 1158 1285
rect 1210 1241 1216 1293
rect 2006 1305 2012 1357
rect 2064 1305 2070 1325
rect 2006 1301 2070 1305
rect 2006 1293 2014 1301
rect 2006 1281 2012 1293
rect 1244 1253 2012 1281
rect 1052 1219 1106 1241
rect 198 1141 262 1165
rect 254 1085 262 1141
rect 290 1218 1106 1219
rect 290 1166 307 1218
rect 359 1181 371 1218
rect 423 1181 435 1218
rect 487 1181 499 1218
rect 551 1166 563 1218
rect 615 1181 627 1218
rect 679 1181 691 1218
rect 743 1181 755 1218
rect 807 1181 819 1218
rect 620 1166 627 1181
rect 871 1166 883 1218
rect 935 1181 947 1218
rect 999 1181 1011 1218
rect 1063 1205 1106 1218
rect 1162 1219 1216 1241
rect 2006 1241 2012 1253
rect 2064 1241 2070 1245
rect 2006 1221 2070 1241
rect 1162 1218 1978 1219
rect 1162 1205 1205 1218
rect 1063 1181 1205 1205
rect 1257 1181 1269 1218
rect 1321 1181 1333 1218
rect 940 1166 947 1181
rect 1063 1166 1106 1181
rect 290 1146 324 1166
rect 380 1146 404 1166
rect 460 1146 484 1166
rect 540 1146 564 1166
rect 620 1146 644 1166
rect 700 1146 724 1166
rect 780 1146 804 1166
rect 860 1146 884 1166
rect 940 1146 964 1166
rect 1020 1146 1106 1166
rect 290 1094 307 1146
rect 359 1094 371 1125
rect 423 1094 435 1125
rect 487 1094 499 1125
rect 551 1094 563 1146
rect 620 1125 627 1146
rect 615 1094 627 1125
rect 679 1094 691 1125
rect 743 1094 755 1125
rect 807 1094 819 1125
rect 871 1094 883 1146
rect 940 1125 947 1146
rect 1063 1125 1106 1146
rect 1162 1166 1205 1181
rect 1321 1166 1328 1181
rect 1385 1166 1397 1218
rect 1449 1181 1461 1218
rect 1513 1181 1525 1218
rect 1577 1181 1589 1218
rect 1641 1181 1653 1218
rect 1641 1166 1648 1181
rect 1705 1166 1717 1218
rect 1769 1181 1781 1218
rect 1833 1181 1845 1218
rect 1897 1181 1909 1218
rect 1961 1166 1978 1218
rect 1162 1146 1248 1166
rect 1304 1146 1328 1166
rect 1384 1146 1408 1166
rect 1464 1146 1488 1166
rect 1544 1146 1568 1166
rect 1624 1146 1648 1166
rect 1704 1146 1728 1166
rect 1784 1146 1808 1166
rect 1864 1146 1888 1166
rect 1944 1146 1978 1166
rect 1162 1125 1205 1146
rect 1321 1125 1328 1146
rect 935 1094 947 1125
rect 999 1094 1011 1125
rect 1063 1101 1205 1125
rect 1063 1094 1106 1101
rect 290 1093 1106 1094
rect 198 1071 262 1085
rect 198 1061 204 1071
rect 256 1059 262 1071
rect 1052 1071 1106 1093
rect 1162 1094 1205 1101
rect 1257 1094 1269 1125
rect 1321 1094 1333 1125
rect 1385 1094 1397 1146
rect 1641 1125 1648 1146
rect 1449 1094 1461 1125
rect 1513 1094 1525 1125
rect 1577 1094 1589 1125
rect 1641 1094 1653 1125
rect 1705 1094 1717 1146
rect 1769 1094 1781 1125
rect 1833 1094 1845 1125
rect 1897 1094 1909 1125
rect 1961 1094 1978 1146
rect 1162 1093 1978 1094
rect 2006 1165 2014 1221
rect 2006 1141 2070 1165
rect 1162 1071 1216 1093
rect 256 1031 1024 1059
rect 256 1019 262 1031
rect 254 1007 262 1019
rect 198 981 204 1005
rect 256 955 262 1007
rect 1052 1019 1058 1071
rect 1110 1021 1158 1045
rect 1210 1019 1216 1071
rect 2006 1085 2014 1141
rect 2006 1071 2070 1085
rect 2006 1059 2012 1071
rect 2064 1061 2070 1071
rect 1244 1031 2012 1059
rect 1052 1007 1106 1019
rect 1162 1007 1216 1019
rect 1052 1003 1058 1007
rect 290 975 1058 1003
rect 254 947 262 955
rect 1052 955 1058 975
rect 1210 1003 1216 1007
rect 2006 1019 2012 1031
rect 2006 1007 2014 1019
rect 1210 975 1978 1003
rect 1110 955 1158 965
rect 1210 955 1216 975
rect 254 943 1024 947
rect 198 901 204 925
rect 256 919 1024 943
rect 1052 943 1216 955
rect 2006 955 2012 1007
rect 2064 981 2070 1005
rect 2006 947 2014 955
rect 256 891 262 919
rect 1052 891 1058 943
rect 1110 941 1158 943
rect 1210 891 1216 943
rect 1244 943 2014 947
rect 1244 919 2012 943
rect 2006 891 2012 919
rect 2064 901 2070 925
rect 254 879 262 891
rect 198 827 204 845
rect 256 835 262 879
rect 290 885 1106 891
rect 1162 885 1978 891
rect 290 879 1978 885
rect 290 863 1058 879
rect 256 827 1024 835
rect 198 821 1024 827
rect 254 815 1024 821
rect 256 807 1024 815
rect 1052 827 1058 863
rect 1110 861 1158 879
rect 1210 863 1978 879
rect 2006 879 2014 891
rect 1210 827 1216 863
rect 2006 835 2012 879
rect 1052 815 1106 827
rect 1162 815 1216 827
rect 198 763 204 765
rect 256 763 262 807
rect 1052 779 1058 815
rect 1110 781 1158 805
rect 198 751 262 763
rect 290 763 1058 779
rect 1210 779 1216 815
rect 1244 827 2012 835
rect 2064 827 2070 845
rect 1244 821 2070 827
rect 1244 815 2014 821
rect 1244 807 2012 815
rect 1210 763 1978 779
rect 290 751 1106 763
rect 1162 751 1978 763
rect 2006 763 2012 807
rect 2064 763 2070 765
rect 2006 751 2070 763
rect 198 741 204 751
rect 256 723 262 751
rect 256 699 1024 723
rect 254 695 1024 699
rect 1052 699 1058 751
rect 1110 701 1158 725
rect 1210 699 1216 751
rect 2006 723 2012 751
rect 2064 741 2070 751
rect 254 687 262 695
rect 198 661 204 685
rect 256 635 262 687
rect 1052 687 1106 699
rect 1162 687 1216 699
rect 1244 699 2012 723
rect 1244 695 2014 699
rect 1052 667 1058 687
rect 290 639 1058 667
rect 1210 667 1216 687
rect 2006 687 2014 695
rect 254 623 262 635
rect 256 611 262 623
rect 1052 635 1058 639
rect 1110 635 1158 645
rect 1210 639 1978 667
rect 1210 635 1216 639
rect 1052 623 1216 635
rect 198 581 204 605
rect 256 583 1024 611
rect 256 571 262 583
rect 254 559 262 571
rect 198 507 204 525
rect 256 507 262 559
rect 1052 571 1058 623
rect 1110 621 1158 623
rect 1210 571 1216 623
rect 2006 635 2012 687
rect 2064 661 2070 685
rect 2006 623 2014 635
rect 2006 611 2012 623
rect 1244 583 2012 611
rect 1052 565 1106 571
rect 1162 565 1216 571
rect 1052 559 1216 565
rect 1052 555 1058 559
rect 290 527 1058 555
rect 1110 541 1158 559
rect 1210 555 1216 559
rect 2006 571 2012 583
rect 2064 581 2070 605
rect 2006 559 2014 571
rect 198 501 262 507
rect 254 499 262 501
rect 1052 507 1058 527
rect 1210 527 1978 555
rect 1210 507 1216 527
rect 254 495 1024 499
rect 256 471 1024 495
rect 1052 495 1106 507
rect 1162 495 1216 507
rect 2006 507 2012 559
rect 2064 507 2070 525
rect 2006 501 2070 507
rect 2006 499 2014 501
rect 198 443 204 445
rect 256 443 262 471
rect 1052 443 1058 495
rect 1110 461 1158 485
rect 1210 443 1216 495
rect 1244 495 2014 499
rect 1244 471 2012 495
rect 2006 443 2012 471
rect 2064 443 2070 445
rect 198 431 262 443
rect 198 421 204 431
rect 256 387 262 431
rect 290 431 1106 443
rect 1162 431 1978 443
rect 290 415 1058 431
rect 256 379 1024 387
rect 254 365 1024 379
rect 198 359 1024 365
rect 1052 379 1058 415
rect 1210 415 1978 431
rect 2006 431 2070 443
rect 1110 381 1158 405
rect 1210 379 1216 415
rect 2006 387 2012 431
rect 2064 421 2070 431
rect 198 341 262 359
rect 254 325 262 341
rect 1052 325 1106 379
rect 1162 325 1216 379
rect 1244 379 2012 387
rect 1244 365 2014 379
rect 1244 359 2070 365
rect 2006 341 2070 359
rect 2006 325 2014 341
rect 254 324 1024 325
rect 254 285 326 324
rect 198 272 326 285
rect 378 272 390 324
rect 442 272 454 324
rect 506 272 518 324
rect 570 272 582 324
rect 634 272 646 324
rect 698 272 710 324
rect 762 272 774 324
rect 826 272 838 324
rect 890 272 902 324
rect 954 272 966 324
rect 1018 272 1024 324
rect 198 271 1024 272
rect 1052 301 1216 325
rect 65 241 169 244
rect 1052 245 1106 301
rect 1162 245 1216 301
rect 1244 324 2014 325
rect 1244 272 1250 324
rect 1302 272 1314 324
rect 1366 272 1378 324
rect 1430 272 1442 324
rect 1494 272 1506 324
rect 1558 272 1570 324
rect 1622 272 1634 324
rect 1686 272 1698 324
rect 1750 272 1762 324
rect 1814 272 1826 324
rect 1878 272 1890 324
rect 1942 285 2014 324
rect 1942 272 2070 285
rect 1244 271 2070 272
rect 2098 2004 2147 2060
rect 2098 1980 2203 2004
rect 2098 1924 2147 1980
rect 2098 1900 2203 1924
rect 2098 1844 2147 1900
rect 2098 1820 2203 1844
rect 2098 1764 2147 1820
rect 2098 1740 2203 1764
rect 2098 1684 2147 1740
rect 2098 1660 2203 1684
rect 2098 1604 2147 1660
rect 2098 1580 2203 1604
rect 2098 1524 2147 1580
rect 2098 1500 2203 1524
rect 2098 1444 2147 1500
rect 2098 1420 2203 1444
rect 2098 1364 2147 1420
rect 2098 1340 2203 1364
rect 2098 1284 2147 1340
rect 2098 1260 2203 1284
rect 2098 1204 2147 1260
rect 2098 1180 2203 1204
rect 2098 1124 2147 1180
rect 2098 1100 2203 1124
rect 2098 1044 2147 1100
rect 2098 1020 2203 1044
rect 2098 964 2147 1020
rect 2098 940 2203 964
rect 2098 884 2147 940
rect 2098 860 2203 884
rect 2098 804 2147 860
rect 2098 780 2203 804
rect 2098 724 2147 780
rect 2098 700 2203 724
rect 2098 644 2147 700
rect 2098 620 2203 644
rect 2098 564 2147 620
rect 2098 540 2203 564
rect 2098 484 2147 540
rect 2098 460 2203 484
rect 2098 404 2147 460
rect 2098 380 2203 404
rect 2098 324 2147 380
rect 2098 300 2203 324
rect 1052 241 1216 245
rect 2098 244 2147 300
rect 2098 241 2203 244
rect 65 221 2203 241
rect 65 220 1106 221
rect 121 165 1106 220
rect 1162 220 2203 221
rect 1162 165 2147 220
rect 121 164 2147 165
rect 65 140 2203 164
rect 121 110 2147 140
rect 121 84 277 110
rect 65 58 277 84
rect 329 58 341 110
rect 393 58 405 110
rect 457 58 469 110
rect 521 58 533 110
rect 585 58 597 110
rect 649 58 661 110
rect 713 58 725 110
rect 777 58 789 110
rect 841 58 853 110
rect 905 58 917 110
rect 969 58 981 110
rect 1033 58 1045 110
rect 1097 58 1109 110
rect 1161 58 1173 110
rect 1225 58 1237 110
rect 1289 58 1301 110
rect 1353 58 1365 110
rect 1417 58 1429 110
rect 1481 58 1493 110
rect 1545 58 1557 110
rect 1609 58 1621 110
rect 1673 58 1685 110
rect 1737 58 1749 110
rect 1801 58 1813 110
rect 1865 58 1877 110
rect 1929 84 2147 110
rect 1929 58 2203 84
rect 65 15 2203 58
<< via2 >>
rect 65 2244 121 2300
rect 2147 2244 2203 2300
rect 65 2164 121 2220
rect 2147 2164 2203 2220
rect 65 2084 121 2140
rect 1106 2085 1162 2141
rect 2147 2084 2203 2140
rect 65 2004 121 2060
rect 65 1924 121 1980
rect 65 1844 121 1900
rect 65 1764 121 1820
rect 65 1684 121 1740
rect 65 1604 121 1660
rect 65 1524 121 1580
rect 65 1444 121 1500
rect 65 1364 121 1420
rect 65 1284 121 1340
rect 65 1204 121 1260
rect 65 1124 121 1180
rect 65 1044 121 1100
rect 65 964 121 1020
rect 65 884 121 940
rect 65 804 121 860
rect 65 724 121 780
rect 65 644 121 700
rect 65 564 121 620
rect 65 484 121 540
rect 65 404 121 460
rect 65 324 121 380
rect 65 244 121 300
rect 198 1965 254 2021
rect 1106 2005 1162 2061
rect 198 1933 254 1941
rect 198 1885 204 1933
rect 204 1885 254 1933
rect 1106 1933 1162 1981
rect 2014 1965 2070 2021
rect 1106 1925 1110 1933
rect 1110 1925 1158 1933
rect 1158 1925 1162 1933
rect 1106 1881 1110 1901
rect 1110 1881 1158 1901
rect 1158 1881 1162 1901
rect 2014 1933 2070 1941
rect 1106 1869 1162 1881
rect 2014 1885 2064 1933
rect 2064 1885 2070 1933
rect 198 1817 204 1861
rect 204 1817 254 1861
rect 198 1805 254 1817
rect 1106 1845 1110 1869
rect 1110 1845 1158 1869
rect 1158 1845 1162 1869
rect 1106 1817 1110 1821
rect 1110 1817 1158 1821
rect 1158 1817 1162 1821
rect 198 1753 204 1781
rect 204 1753 254 1781
rect 1106 1805 1162 1817
rect 2014 1817 2064 1861
rect 2064 1817 2070 1861
rect 1106 1765 1110 1805
rect 1110 1765 1158 1805
rect 1158 1765 1162 1805
rect 2014 1805 2070 1817
rect 198 1741 254 1753
rect 198 1725 204 1741
rect 204 1725 254 1741
rect 198 1689 204 1701
rect 204 1689 254 1701
rect 198 1677 254 1689
rect 198 1645 204 1677
rect 204 1645 254 1677
rect 1106 1689 1110 1741
rect 1110 1689 1158 1741
rect 1158 1689 1162 1741
rect 2014 1753 2064 1781
rect 2064 1753 2070 1781
rect 2014 1741 2070 1753
rect 2014 1725 2064 1741
rect 2064 1725 2070 1741
rect 1106 1685 1162 1689
rect 2014 1689 2064 1701
rect 2064 1689 2070 1701
rect 2014 1677 2070 1689
rect 198 1613 254 1621
rect 1106 1625 1110 1661
rect 1110 1625 1158 1661
rect 1158 1625 1162 1661
rect 198 1565 204 1613
rect 204 1565 254 1613
rect 1106 1613 1162 1625
rect 2014 1645 2064 1677
rect 2064 1645 2070 1677
rect 1106 1605 1110 1613
rect 1110 1605 1158 1613
rect 1158 1605 1162 1613
rect 1106 1561 1110 1581
rect 1110 1561 1158 1581
rect 1158 1561 1162 1581
rect 2014 1613 2070 1621
rect 2014 1565 2064 1613
rect 2064 1565 2070 1613
rect 198 1497 204 1541
rect 204 1497 254 1541
rect 1106 1549 1162 1561
rect 198 1485 254 1497
rect 1106 1525 1110 1549
rect 1110 1525 1158 1549
rect 1158 1525 1162 1549
rect 1106 1497 1110 1501
rect 1110 1497 1158 1501
rect 1158 1497 1162 1501
rect 1106 1485 1162 1497
rect 198 1433 204 1461
rect 204 1433 254 1461
rect 198 1421 254 1433
rect 1106 1445 1110 1485
rect 1110 1445 1158 1485
rect 1158 1445 1162 1485
rect 2014 1497 2064 1541
rect 2064 1497 2070 1541
rect 2014 1485 2070 1497
rect 2014 1433 2064 1461
rect 2064 1433 2070 1461
rect 2014 1421 2070 1433
rect 198 1405 204 1421
rect 204 1405 254 1421
rect 198 1369 204 1381
rect 204 1369 254 1381
rect 198 1357 254 1369
rect 1106 1369 1110 1421
rect 1110 1369 1158 1421
rect 1158 1369 1162 1421
rect 2014 1405 2064 1421
rect 2064 1405 2070 1421
rect 1106 1365 1162 1369
rect 2014 1369 2064 1381
rect 2064 1369 2070 1381
rect 198 1325 204 1357
rect 204 1325 254 1357
rect 198 1293 254 1301
rect 198 1245 204 1293
rect 204 1245 254 1293
rect 1106 1305 1110 1341
rect 1110 1305 1158 1341
rect 1158 1305 1162 1341
rect 2014 1357 2070 1369
rect 1106 1293 1162 1305
rect 198 1165 254 1221
rect 1106 1285 1110 1293
rect 1110 1285 1158 1293
rect 1158 1285 1162 1293
rect 1106 1241 1110 1261
rect 1110 1241 1158 1261
rect 1158 1241 1162 1261
rect 2014 1325 2064 1357
rect 2064 1325 2070 1357
rect 2014 1293 2070 1301
rect 198 1085 254 1141
rect 324 1166 359 1181
rect 359 1166 371 1181
rect 371 1166 380 1181
rect 404 1166 423 1181
rect 423 1166 435 1181
rect 435 1166 460 1181
rect 484 1166 487 1181
rect 487 1166 499 1181
rect 499 1166 540 1181
rect 564 1166 615 1181
rect 615 1166 620 1181
rect 644 1166 679 1181
rect 679 1166 691 1181
rect 691 1166 700 1181
rect 724 1166 743 1181
rect 743 1166 755 1181
rect 755 1166 780 1181
rect 804 1166 807 1181
rect 807 1166 819 1181
rect 819 1166 860 1181
rect 1106 1205 1162 1241
rect 2014 1245 2064 1293
rect 2064 1245 2070 1293
rect 884 1166 935 1181
rect 935 1166 940 1181
rect 964 1166 999 1181
rect 999 1166 1011 1181
rect 1011 1166 1020 1181
rect 324 1146 380 1166
rect 404 1146 460 1166
rect 484 1146 540 1166
rect 564 1146 620 1166
rect 644 1146 700 1166
rect 724 1146 780 1166
rect 804 1146 860 1166
rect 884 1146 940 1166
rect 964 1146 1020 1166
rect 324 1125 359 1146
rect 359 1125 371 1146
rect 371 1125 380 1146
rect 404 1125 423 1146
rect 423 1125 435 1146
rect 435 1125 460 1146
rect 484 1125 487 1146
rect 487 1125 499 1146
rect 499 1125 540 1146
rect 564 1125 615 1146
rect 615 1125 620 1146
rect 644 1125 679 1146
rect 679 1125 691 1146
rect 691 1125 700 1146
rect 724 1125 743 1146
rect 743 1125 755 1146
rect 755 1125 780 1146
rect 804 1125 807 1146
rect 807 1125 819 1146
rect 819 1125 860 1146
rect 884 1125 935 1146
rect 935 1125 940 1146
rect 964 1125 999 1146
rect 999 1125 1011 1146
rect 1011 1125 1020 1146
rect 1106 1125 1162 1181
rect 1248 1166 1257 1181
rect 1257 1166 1269 1181
rect 1269 1166 1304 1181
rect 1328 1166 1333 1181
rect 1333 1166 1384 1181
rect 1408 1166 1449 1181
rect 1449 1166 1461 1181
rect 1461 1166 1464 1181
rect 1488 1166 1513 1181
rect 1513 1166 1525 1181
rect 1525 1166 1544 1181
rect 1568 1166 1577 1181
rect 1577 1166 1589 1181
rect 1589 1166 1624 1181
rect 1648 1166 1653 1181
rect 1653 1166 1704 1181
rect 1728 1166 1769 1181
rect 1769 1166 1781 1181
rect 1781 1166 1784 1181
rect 1808 1166 1833 1181
rect 1833 1166 1845 1181
rect 1845 1166 1864 1181
rect 1888 1166 1897 1181
rect 1897 1166 1909 1181
rect 1909 1166 1944 1181
rect 1248 1146 1304 1166
rect 1328 1146 1384 1166
rect 1408 1146 1464 1166
rect 1488 1146 1544 1166
rect 1568 1146 1624 1166
rect 1648 1146 1704 1166
rect 1728 1146 1784 1166
rect 1808 1146 1864 1166
rect 1888 1146 1944 1166
rect 1248 1125 1257 1146
rect 1257 1125 1269 1146
rect 1269 1125 1304 1146
rect 1328 1125 1333 1146
rect 1333 1125 1384 1146
rect 198 1019 204 1061
rect 204 1019 254 1061
rect 1106 1071 1162 1101
rect 1408 1125 1449 1146
rect 1449 1125 1461 1146
rect 1461 1125 1464 1146
rect 1488 1125 1513 1146
rect 1513 1125 1525 1146
rect 1525 1125 1544 1146
rect 1568 1125 1577 1146
rect 1577 1125 1589 1146
rect 1589 1125 1624 1146
rect 1648 1125 1653 1146
rect 1653 1125 1704 1146
rect 1728 1125 1769 1146
rect 1769 1125 1781 1146
rect 1781 1125 1784 1146
rect 1808 1125 1833 1146
rect 1833 1125 1845 1146
rect 1845 1125 1864 1146
rect 1888 1125 1897 1146
rect 1897 1125 1909 1146
rect 1909 1125 1944 1146
rect 2014 1165 2070 1221
rect 198 1007 254 1019
rect 198 1005 204 1007
rect 204 1005 254 1007
rect 198 955 204 981
rect 204 955 254 981
rect 1106 1045 1110 1071
rect 1110 1045 1158 1071
rect 1158 1045 1162 1071
rect 1106 1019 1110 1021
rect 1110 1019 1158 1021
rect 1158 1019 1162 1021
rect 2014 1085 2070 1141
rect 1106 1007 1162 1019
rect 198 943 254 955
rect 1106 965 1110 1007
rect 1110 965 1158 1007
rect 1158 965 1162 1007
rect 2014 1019 2064 1061
rect 2064 1019 2070 1061
rect 2014 1007 2070 1019
rect 198 925 204 943
rect 204 925 254 943
rect 2014 1005 2064 1007
rect 2064 1005 2070 1007
rect 2014 955 2064 981
rect 2064 955 2070 981
rect 198 891 204 901
rect 204 891 254 901
rect 1106 891 1110 941
rect 1110 891 1158 941
rect 1158 891 1162 941
rect 2014 943 2070 955
rect 2014 925 2064 943
rect 2064 925 2070 943
rect 2014 891 2064 901
rect 2064 891 2070 901
rect 198 879 254 891
rect 198 845 204 879
rect 204 845 254 879
rect 1106 885 1162 891
rect 198 815 254 821
rect 198 765 204 815
rect 204 765 254 815
rect 2014 879 2070 891
rect 1106 827 1110 861
rect 1110 827 1158 861
rect 1158 827 1162 861
rect 2014 845 2064 879
rect 2064 845 2070 879
rect 1106 815 1162 827
rect 1106 805 1110 815
rect 1110 805 1158 815
rect 1158 805 1162 815
rect 1106 763 1110 781
rect 1110 763 1158 781
rect 1158 763 1162 781
rect 2014 815 2070 821
rect 1106 751 1162 763
rect 2014 765 2064 815
rect 2064 765 2070 815
rect 198 699 204 741
rect 204 699 254 741
rect 198 687 254 699
rect 1106 725 1110 751
rect 1110 725 1158 751
rect 1158 725 1162 751
rect 1106 699 1110 701
rect 1110 699 1158 701
rect 1158 699 1162 701
rect 198 685 204 687
rect 204 685 254 687
rect 198 635 204 661
rect 204 635 254 661
rect 1106 687 1162 699
rect 2014 699 2064 741
rect 2064 699 2070 741
rect 1106 645 1110 687
rect 1110 645 1158 687
rect 1158 645 1162 687
rect 2014 687 2070 699
rect 198 623 254 635
rect 198 605 204 623
rect 204 605 254 623
rect 198 571 204 581
rect 204 571 254 581
rect 198 559 254 571
rect 198 525 204 559
rect 204 525 254 559
rect 1106 571 1110 621
rect 1110 571 1158 621
rect 1158 571 1162 621
rect 2014 685 2064 687
rect 2064 685 2070 687
rect 2014 635 2064 661
rect 2064 635 2070 661
rect 2014 623 2070 635
rect 2014 605 2064 623
rect 2064 605 2070 623
rect 1106 565 1162 571
rect 2014 571 2064 581
rect 2064 571 2070 581
rect 2014 559 2070 571
rect 198 495 254 501
rect 1106 507 1110 541
rect 1110 507 1158 541
rect 1158 507 1162 541
rect 198 445 204 495
rect 204 445 254 495
rect 1106 495 1162 507
rect 2014 525 2064 559
rect 2064 525 2070 559
rect 1106 485 1110 495
rect 1110 485 1158 495
rect 1158 485 1162 495
rect 1106 443 1110 461
rect 1110 443 1158 461
rect 1158 443 1162 461
rect 2014 495 2070 501
rect 2014 445 2064 495
rect 2064 445 2070 495
rect 198 379 204 421
rect 204 379 254 421
rect 1106 431 1162 443
rect 198 365 254 379
rect 1106 405 1110 431
rect 1110 405 1158 431
rect 1158 405 1162 431
rect 1106 379 1110 381
rect 1110 379 1158 381
rect 1158 379 1162 381
rect 198 285 254 341
rect 1106 325 1162 379
rect 2014 379 2064 421
rect 2064 379 2070 421
rect 2014 365 2070 379
rect 1106 245 1162 301
rect 2014 285 2070 341
rect 2147 2004 2203 2060
rect 2147 1924 2203 1980
rect 2147 1844 2203 1900
rect 2147 1764 2203 1820
rect 2147 1684 2203 1740
rect 2147 1604 2203 1660
rect 2147 1524 2203 1580
rect 2147 1444 2203 1500
rect 2147 1364 2203 1420
rect 2147 1284 2203 1340
rect 2147 1204 2203 1260
rect 2147 1124 2203 1180
rect 2147 1044 2203 1100
rect 2147 964 2203 1020
rect 2147 884 2203 940
rect 2147 804 2203 860
rect 2147 724 2203 780
rect 2147 644 2203 700
rect 2147 564 2203 620
rect 2147 484 2203 540
rect 2147 404 2203 460
rect 2147 324 2203 380
rect 2147 244 2203 300
rect 65 164 121 220
rect 1106 165 1162 221
rect 2147 164 2203 220
rect 65 84 121 140
rect 2147 84 2203 140
<< metal3 >>
rect 60 2304 126 2323
rect 60 2240 61 2304
rect 125 2240 126 2304
rect 2142 2304 2208 2323
rect 60 2224 126 2240
rect 60 2160 61 2224
rect 125 2160 126 2224
rect 60 2144 126 2160
rect 60 2080 61 2144
rect 125 2080 126 2144
rect 60 2064 126 2080
rect 60 2000 61 2064
rect 125 2000 126 2064
rect 60 1984 126 2000
rect 60 1920 61 1984
rect 125 1920 126 1984
rect 60 1904 126 1920
rect 60 1840 61 1904
rect 125 1840 126 1904
rect 60 1824 126 1840
rect 60 1760 61 1824
rect 125 1760 126 1824
rect 60 1744 126 1760
rect 60 1680 61 1744
rect 125 1680 126 1744
rect 60 1664 126 1680
rect 60 1600 61 1664
rect 125 1600 126 1664
rect 60 1584 126 1600
rect 60 1520 61 1584
rect 125 1520 126 1584
rect 60 1504 126 1520
rect 60 1440 61 1504
rect 125 1440 126 1504
rect 60 1424 126 1440
rect 60 1360 61 1424
rect 125 1360 126 1424
rect 60 1344 126 1360
rect 60 1280 61 1344
rect 125 1280 126 1344
rect 60 1264 126 1280
rect 60 1200 61 1264
rect 125 1200 126 1264
rect 60 1184 126 1200
rect 60 1120 61 1184
rect 125 1120 126 1184
rect 60 1104 126 1120
rect 60 1040 61 1104
rect 125 1040 126 1104
rect 60 1024 126 1040
rect 60 960 61 1024
rect 125 960 126 1024
rect 60 944 126 960
rect 60 880 61 944
rect 125 880 126 944
rect 60 864 126 880
rect 60 800 61 864
rect 125 800 126 864
rect 60 784 126 800
rect 60 720 61 784
rect 125 720 126 784
rect 60 704 126 720
rect 60 640 61 704
rect 125 640 126 704
rect 60 624 126 640
rect 60 560 61 624
rect 125 560 126 624
rect 60 544 126 560
rect 60 480 61 544
rect 125 480 126 544
rect 60 464 126 480
rect 60 400 61 464
rect 125 400 126 464
rect 60 384 126 400
rect 60 320 61 384
rect 125 320 126 384
rect 60 304 126 320
rect 60 240 61 304
rect 125 240 126 304
rect 60 224 126 240
rect 60 160 61 224
rect 125 160 126 224
rect 60 144 126 160
rect 60 80 61 144
rect 125 80 126 144
rect 60 15 126 80
rect 193 2271 2075 2272
rect 193 2207 262 2271
rect 326 2207 342 2271
rect 406 2207 422 2271
rect 486 2207 502 2271
rect 566 2207 582 2271
rect 646 2207 662 2271
rect 726 2207 742 2271
rect 806 2207 822 2271
rect 886 2207 902 2271
rect 966 2207 982 2271
rect 1046 2207 1062 2271
rect 1126 2207 1142 2271
rect 1206 2207 1222 2271
rect 1286 2207 1302 2271
rect 1366 2207 1382 2271
rect 1446 2207 1462 2271
rect 1526 2207 1542 2271
rect 1606 2207 1622 2271
rect 1686 2207 1702 2271
rect 1766 2207 1782 2271
rect 1846 2207 1862 2271
rect 1926 2207 1942 2271
rect 2006 2207 2075 2271
rect 193 2206 2075 2207
rect 193 2185 259 2206
rect 193 2121 194 2185
rect 258 2121 259 2185
rect 2009 2185 2075 2206
rect 193 2105 259 2121
rect 193 2041 194 2105
rect 258 2041 259 2105
rect 319 2145 1949 2146
rect 319 2086 1102 2145
rect 193 2026 259 2041
rect 1101 2081 1102 2086
rect 1166 2086 1949 2145
rect 2009 2121 2010 2185
rect 2074 2121 2075 2185
rect 2009 2105 2075 2121
rect 1166 2081 1167 2086
rect 1101 2065 1167 2081
rect 193 2025 1041 2026
rect 193 1961 194 2025
rect 258 1966 1041 2025
rect 1101 2001 1102 2065
rect 1166 2001 1167 2065
rect 2009 2041 2010 2105
rect 2074 2041 2075 2105
rect 2009 2026 2075 2041
rect 1101 1985 1167 2001
rect 258 1961 259 1966
rect 193 1945 259 1961
rect 193 1881 194 1945
rect 258 1881 259 1945
rect 1101 1921 1102 1985
rect 1166 1921 1167 1985
rect 1227 2025 2075 2026
rect 1227 1966 2010 2025
rect 1101 1906 1167 1921
rect 2009 1961 2010 1966
rect 2074 1961 2075 2025
rect 2009 1945 2075 1961
rect 193 1865 259 1881
rect 193 1801 194 1865
rect 258 1801 259 1865
rect 319 1905 1949 1906
rect 319 1846 1102 1905
rect 193 1786 259 1801
rect 1101 1841 1102 1846
rect 1166 1846 1949 1905
rect 2009 1881 2010 1945
rect 2074 1881 2075 1945
rect 2009 1865 2075 1881
rect 1166 1841 1167 1846
rect 1101 1825 1167 1841
rect 193 1785 1041 1786
rect 193 1721 194 1785
rect 258 1726 1041 1785
rect 1101 1761 1102 1825
rect 1166 1761 1167 1825
rect 2009 1801 2010 1865
rect 2074 1801 2075 1865
rect 2009 1786 2075 1801
rect 1101 1745 1167 1761
rect 258 1721 259 1726
rect 193 1705 259 1721
rect 193 1641 194 1705
rect 258 1641 259 1705
rect 1101 1681 1102 1745
rect 1166 1681 1167 1745
rect 1227 1785 2075 1786
rect 1227 1726 2010 1785
rect 1101 1666 1167 1681
rect 2009 1721 2010 1726
rect 2074 1721 2075 1785
rect 2009 1705 2075 1721
rect 193 1625 259 1641
rect 193 1561 194 1625
rect 258 1561 259 1625
rect 319 1665 1949 1666
rect 319 1606 1102 1665
rect 193 1546 259 1561
rect 1101 1601 1102 1606
rect 1166 1606 1949 1665
rect 2009 1641 2010 1705
rect 2074 1641 2075 1705
rect 2009 1625 2075 1641
rect 1166 1601 1167 1606
rect 1101 1585 1167 1601
rect 193 1545 1041 1546
rect 193 1481 194 1545
rect 258 1486 1041 1545
rect 1101 1521 1102 1585
rect 1166 1521 1167 1585
rect 2009 1561 2010 1625
rect 2074 1561 2075 1625
rect 2009 1546 2075 1561
rect 1101 1505 1167 1521
rect 258 1481 259 1486
rect 193 1465 259 1481
rect 193 1401 194 1465
rect 258 1401 259 1465
rect 1101 1441 1102 1505
rect 1166 1441 1167 1505
rect 1227 1545 2075 1546
rect 1227 1486 2010 1545
rect 1101 1426 1167 1441
rect 2009 1481 2010 1486
rect 2074 1481 2075 1545
rect 2009 1465 2075 1481
rect 193 1385 259 1401
rect 193 1321 194 1385
rect 258 1321 259 1385
rect 319 1425 1949 1426
rect 319 1366 1102 1425
rect 193 1306 259 1321
rect 1101 1361 1102 1366
rect 1166 1366 1949 1425
rect 2009 1401 2010 1465
rect 2074 1401 2075 1465
rect 2009 1385 2075 1401
rect 1166 1361 1167 1366
rect 1101 1345 1167 1361
rect 193 1305 1041 1306
rect 193 1241 194 1305
rect 258 1246 1041 1305
rect 1101 1281 1102 1345
rect 1166 1281 1167 1345
rect 2009 1321 2010 1385
rect 2074 1321 2075 1385
rect 2009 1306 2075 1321
rect 1101 1265 1167 1281
rect 258 1241 259 1246
rect 193 1225 259 1241
rect 193 1161 194 1225
rect 258 1161 259 1225
rect 1101 1201 1102 1265
rect 1166 1201 1167 1265
rect 1227 1305 2075 1306
rect 1227 1246 2010 1305
rect 1101 1186 1167 1201
rect 2009 1241 2010 1246
rect 2074 1241 2075 1305
rect 2009 1225 2075 1241
rect 193 1145 259 1161
rect 193 1081 194 1145
rect 258 1081 259 1145
rect 319 1185 1949 1186
rect 319 1181 325 1185
rect 389 1181 405 1185
rect 469 1181 485 1185
rect 549 1181 565 1185
rect 629 1181 645 1185
rect 709 1181 725 1185
rect 789 1181 805 1185
rect 869 1181 885 1185
rect 949 1181 965 1185
rect 319 1125 324 1181
rect 389 1125 404 1181
rect 469 1125 484 1181
rect 549 1125 564 1181
rect 629 1125 644 1181
rect 709 1125 724 1181
rect 789 1125 804 1181
rect 869 1125 884 1181
rect 949 1125 964 1181
rect 319 1121 325 1125
rect 389 1121 405 1125
rect 469 1121 485 1125
rect 549 1121 565 1125
rect 629 1121 645 1125
rect 709 1121 725 1125
rect 789 1121 805 1125
rect 869 1121 885 1125
rect 949 1121 965 1125
rect 1029 1121 1102 1185
rect 1166 1121 1239 1185
rect 1303 1181 1319 1185
rect 1383 1181 1399 1185
rect 1463 1181 1479 1185
rect 1543 1181 1559 1185
rect 1623 1181 1639 1185
rect 1703 1181 1719 1185
rect 1783 1181 1799 1185
rect 1863 1181 1879 1185
rect 1943 1181 1949 1185
rect 1304 1125 1319 1181
rect 1384 1125 1399 1181
rect 1464 1125 1479 1181
rect 1544 1125 1559 1181
rect 1624 1125 1639 1181
rect 1704 1125 1719 1181
rect 1784 1125 1799 1181
rect 1864 1125 1879 1181
rect 1944 1125 1949 1181
rect 1303 1121 1319 1125
rect 1383 1121 1399 1125
rect 1463 1121 1479 1125
rect 1543 1121 1559 1125
rect 1623 1121 1639 1125
rect 1703 1121 1719 1125
rect 1783 1121 1799 1125
rect 1863 1121 1879 1125
rect 1943 1121 1949 1125
rect 319 1120 1949 1121
rect 2009 1161 2010 1225
rect 2074 1161 2075 1225
rect 2009 1145 2075 1161
rect 193 1065 259 1081
rect 193 1001 194 1065
rect 258 1060 259 1065
rect 1101 1105 1167 1120
rect 258 1001 1041 1060
rect 193 1000 1041 1001
rect 1101 1041 1102 1105
rect 1166 1041 1167 1105
rect 2009 1081 2010 1145
rect 2074 1081 2075 1145
rect 2009 1065 2075 1081
rect 2009 1060 2010 1065
rect 1101 1025 1167 1041
rect 193 985 259 1000
rect 193 921 194 985
rect 258 921 259 985
rect 1101 961 1102 1025
rect 1166 961 1167 1025
rect 1227 1001 2010 1060
rect 2074 1001 2075 1065
rect 1227 1000 2075 1001
rect 1101 945 1167 961
rect 1101 940 1102 945
rect 193 905 259 921
rect 193 841 194 905
rect 258 841 259 905
rect 319 881 1102 940
rect 1166 940 1167 945
rect 2009 985 2075 1000
rect 1166 881 1949 940
rect 319 880 1949 881
rect 2009 921 2010 985
rect 2074 921 2075 985
rect 2009 905 2075 921
rect 193 825 259 841
rect 193 761 194 825
rect 258 820 259 825
rect 1101 865 1167 880
rect 258 761 1041 820
rect 193 760 1041 761
rect 1101 801 1102 865
rect 1166 801 1167 865
rect 2009 841 2010 905
rect 2074 841 2075 905
rect 2009 825 2075 841
rect 2009 820 2010 825
rect 1101 785 1167 801
rect 193 745 259 760
rect 193 681 194 745
rect 258 681 259 745
rect 1101 721 1102 785
rect 1166 721 1167 785
rect 1227 761 2010 820
rect 2074 761 2075 825
rect 1227 760 2075 761
rect 1101 705 1167 721
rect 1101 700 1102 705
rect 193 665 259 681
rect 193 601 194 665
rect 258 601 259 665
rect 319 641 1102 700
rect 1166 700 1167 705
rect 2009 745 2075 760
rect 1166 641 1949 700
rect 319 640 1949 641
rect 2009 681 2010 745
rect 2074 681 2075 745
rect 2009 665 2075 681
rect 193 585 259 601
rect 193 521 194 585
rect 258 580 259 585
rect 1101 625 1167 640
rect 258 521 1041 580
rect 193 520 1041 521
rect 1101 561 1102 625
rect 1166 561 1167 625
rect 2009 601 2010 665
rect 2074 601 2075 665
rect 2009 585 2075 601
rect 2009 580 2010 585
rect 1101 545 1167 561
rect 193 505 259 520
rect 193 441 194 505
rect 258 441 259 505
rect 1101 481 1102 545
rect 1166 481 1167 545
rect 1227 521 2010 580
rect 2074 521 2075 585
rect 1227 520 2075 521
rect 1101 465 1167 481
rect 1101 460 1102 465
rect 193 425 259 441
rect 193 361 194 425
rect 258 361 259 425
rect 319 401 1102 460
rect 1166 460 1167 465
rect 2009 505 2075 520
rect 1166 401 1949 460
rect 319 400 1949 401
rect 2009 441 2010 505
rect 2074 441 2075 505
rect 2009 425 2075 441
rect 193 345 259 361
rect 193 281 194 345
rect 258 340 259 345
rect 1101 385 1167 400
rect 258 281 1041 340
rect 193 280 1041 281
rect 1101 321 1102 385
rect 1166 321 1167 385
rect 2009 361 2010 425
rect 2074 361 2075 425
rect 2009 345 2075 361
rect 2009 340 2010 345
rect 1101 305 1167 321
rect 193 265 259 280
rect 193 201 194 265
rect 258 201 259 265
rect 1101 241 1102 305
rect 1166 241 1167 305
rect 1227 281 2010 340
rect 2074 281 2075 345
rect 1227 280 2075 281
rect 1101 225 1167 241
rect 1101 220 1102 225
rect 193 185 259 201
rect 193 121 194 185
rect 258 121 259 185
rect 319 161 1102 220
rect 1166 220 1167 225
rect 2009 265 2075 280
rect 1166 161 1949 220
rect 319 160 1949 161
rect 2009 201 2010 265
rect 2074 201 2075 265
rect 2009 185 2075 201
rect 193 100 259 121
rect 2009 121 2010 185
rect 2074 121 2075 185
rect 2009 100 2075 121
rect 193 99 2075 100
rect 193 35 262 99
rect 326 35 342 99
rect 406 35 422 99
rect 486 35 502 99
rect 566 35 582 99
rect 646 35 662 99
rect 726 35 742 99
rect 806 35 822 99
rect 886 35 902 99
rect 966 35 982 99
rect 1046 35 1062 99
rect 1126 35 1142 99
rect 1206 35 1222 99
rect 1286 35 1302 99
rect 1366 35 1382 99
rect 1446 35 1462 99
rect 1526 35 1542 99
rect 1606 35 1622 99
rect 1686 35 1702 99
rect 1766 35 1782 99
rect 1846 35 1862 99
rect 1926 35 1942 99
rect 2006 35 2075 99
rect 193 34 2075 35
rect 2142 2240 2143 2304
rect 2207 2240 2208 2304
rect 2142 2224 2208 2240
rect 2142 2160 2143 2224
rect 2207 2160 2208 2224
rect 2142 2144 2208 2160
rect 2142 2080 2143 2144
rect 2207 2080 2208 2144
rect 2142 2064 2208 2080
rect 2142 2000 2143 2064
rect 2207 2000 2208 2064
rect 2142 1984 2208 2000
rect 2142 1920 2143 1984
rect 2207 1920 2208 1984
rect 2142 1904 2208 1920
rect 2142 1840 2143 1904
rect 2207 1840 2208 1904
rect 2142 1824 2208 1840
rect 2142 1760 2143 1824
rect 2207 1760 2208 1824
rect 2142 1744 2208 1760
rect 2142 1680 2143 1744
rect 2207 1680 2208 1744
rect 2142 1664 2208 1680
rect 2142 1600 2143 1664
rect 2207 1600 2208 1664
rect 2142 1584 2208 1600
rect 2142 1520 2143 1584
rect 2207 1520 2208 1584
rect 2142 1504 2208 1520
rect 2142 1440 2143 1504
rect 2207 1440 2208 1504
rect 2142 1424 2208 1440
rect 2142 1360 2143 1424
rect 2207 1360 2208 1424
rect 2142 1344 2208 1360
rect 2142 1280 2143 1344
rect 2207 1280 2208 1344
rect 2142 1264 2208 1280
rect 2142 1200 2143 1264
rect 2207 1200 2208 1264
rect 2142 1184 2208 1200
rect 2142 1120 2143 1184
rect 2207 1120 2208 1184
rect 2142 1104 2208 1120
rect 2142 1040 2143 1104
rect 2207 1040 2208 1104
rect 2142 1024 2208 1040
rect 2142 960 2143 1024
rect 2207 960 2208 1024
rect 2142 944 2208 960
rect 2142 880 2143 944
rect 2207 880 2208 944
rect 2142 864 2208 880
rect 2142 800 2143 864
rect 2207 800 2208 864
rect 2142 784 2208 800
rect 2142 720 2143 784
rect 2207 720 2208 784
rect 2142 704 2208 720
rect 2142 640 2143 704
rect 2207 640 2208 704
rect 2142 624 2208 640
rect 2142 560 2143 624
rect 2207 560 2208 624
rect 2142 544 2208 560
rect 2142 480 2143 544
rect 2207 480 2208 544
rect 2142 464 2208 480
rect 2142 400 2143 464
rect 2207 400 2208 464
rect 2142 384 2208 400
rect 2142 320 2143 384
rect 2207 320 2208 384
rect 2142 304 2208 320
rect 2142 240 2143 304
rect 2207 240 2208 304
rect 2142 224 2208 240
rect 2142 160 2143 224
rect 2207 160 2208 224
rect 2142 144 2208 160
rect 2142 80 2143 144
rect 2207 80 2208 144
rect 2142 15 2208 80
<< via3 >>
rect 61 2300 125 2304
rect 61 2244 65 2300
rect 65 2244 121 2300
rect 121 2244 125 2300
rect 61 2240 125 2244
rect 61 2220 125 2224
rect 61 2164 65 2220
rect 65 2164 121 2220
rect 121 2164 125 2220
rect 61 2160 125 2164
rect 61 2140 125 2144
rect 61 2084 65 2140
rect 65 2084 121 2140
rect 121 2084 125 2140
rect 61 2080 125 2084
rect 61 2060 125 2064
rect 61 2004 65 2060
rect 65 2004 121 2060
rect 121 2004 125 2060
rect 61 2000 125 2004
rect 61 1980 125 1984
rect 61 1924 65 1980
rect 65 1924 121 1980
rect 121 1924 125 1980
rect 61 1920 125 1924
rect 61 1900 125 1904
rect 61 1844 65 1900
rect 65 1844 121 1900
rect 121 1844 125 1900
rect 61 1840 125 1844
rect 61 1820 125 1824
rect 61 1764 65 1820
rect 65 1764 121 1820
rect 121 1764 125 1820
rect 61 1760 125 1764
rect 61 1740 125 1744
rect 61 1684 65 1740
rect 65 1684 121 1740
rect 121 1684 125 1740
rect 61 1680 125 1684
rect 61 1660 125 1664
rect 61 1604 65 1660
rect 65 1604 121 1660
rect 121 1604 125 1660
rect 61 1600 125 1604
rect 61 1580 125 1584
rect 61 1524 65 1580
rect 65 1524 121 1580
rect 121 1524 125 1580
rect 61 1520 125 1524
rect 61 1500 125 1504
rect 61 1444 65 1500
rect 65 1444 121 1500
rect 121 1444 125 1500
rect 61 1440 125 1444
rect 61 1420 125 1424
rect 61 1364 65 1420
rect 65 1364 121 1420
rect 121 1364 125 1420
rect 61 1360 125 1364
rect 61 1340 125 1344
rect 61 1284 65 1340
rect 65 1284 121 1340
rect 121 1284 125 1340
rect 61 1280 125 1284
rect 61 1260 125 1264
rect 61 1204 65 1260
rect 65 1204 121 1260
rect 121 1204 125 1260
rect 61 1200 125 1204
rect 61 1180 125 1184
rect 61 1124 65 1180
rect 65 1124 121 1180
rect 121 1124 125 1180
rect 61 1120 125 1124
rect 61 1100 125 1104
rect 61 1044 65 1100
rect 65 1044 121 1100
rect 121 1044 125 1100
rect 61 1040 125 1044
rect 61 1020 125 1024
rect 61 964 65 1020
rect 65 964 121 1020
rect 121 964 125 1020
rect 61 960 125 964
rect 61 940 125 944
rect 61 884 65 940
rect 65 884 121 940
rect 121 884 125 940
rect 61 880 125 884
rect 61 860 125 864
rect 61 804 65 860
rect 65 804 121 860
rect 121 804 125 860
rect 61 800 125 804
rect 61 780 125 784
rect 61 724 65 780
rect 65 724 121 780
rect 121 724 125 780
rect 61 720 125 724
rect 61 700 125 704
rect 61 644 65 700
rect 65 644 121 700
rect 121 644 125 700
rect 61 640 125 644
rect 61 620 125 624
rect 61 564 65 620
rect 65 564 121 620
rect 121 564 125 620
rect 61 560 125 564
rect 61 540 125 544
rect 61 484 65 540
rect 65 484 121 540
rect 121 484 125 540
rect 61 480 125 484
rect 61 460 125 464
rect 61 404 65 460
rect 65 404 121 460
rect 121 404 125 460
rect 61 400 125 404
rect 61 380 125 384
rect 61 324 65 380
rect 65 324 121 380
rect 121 324 125 380
rect 61 320 125 324
rect 61 300 125 304
rect 61 244 65 300
rect 65 244 121 300
rect 121 244 125 300
rect 61 240 125 244
rect 61 220 125 224
rect 61 164 65 220
rect 65 164 121 220
rect 121 164 125 220
rect 61 160 125 164
rect 61 140 125 144
rect 61 84 65 140
rect 65 84 121 140
rect 121 84 125 140
rect 61 80 125 84
rect 262 2207 326 2271
rect 342 2207 406 2271
rect 422 2207 486 2271
rect 502 2207 566 2271
rect 582 2207 646 2271
rect 662 2207 726 2271
rect 742 2207 806 2271
rect 822 2207 886 2271
rect 902 2207 966 2271
rect 982 2207 1046 2271
rect 1062 2207 1126 2271
rect 1142 2207 1206 2271
rect 1222 2207 1286 2271
rect 1302 2207 1366 2271
rect 1382 2207 1446 2271
rect 1462 2207 1526 2271
rect 1542 2207 1606 2271
rect 1622 2207 1686 2271
rect 1702 2207 1766 2271
rect 1782 2207 1846 2271
rect 1862 2207 1926 2271
rect 1942 2207 2006 2271
rect 194 2121 258 2185
rect 194 2041 258 2105
rect 1102 2141 1166 2145
rect 1102 2085 1106 2141
rect 1106 2085 1162 2141
rect 1162 2085 1166 2141
rect 2010 2121 2074 2185
rect 1102 2081 1166 2085
rect 194 2021 258 2025
rect 194 1965 198 2021
rect 198 1965 254 2021
rect 254 1965 258 2021
rect 1102 2061 1166 2065
rect 1102 2005 1106 2061
rect 1106 2005 1162 2061
rect 1162 2005 1166 2061
rect 1102 2001 1166 2005
rect 2010 2041 2074 2105
rect 194 1961 258 1965
rect 194 1941 258 1945
rect 194 1885 198 1941
rect 198 1885 254 1941
rect 254 1885 258 1941
rect 194 1881 258 1885
rect 1102 1981 1166 1985
rect 1102 1925 1106 1981
rect 1106 1925 1162 1981
rect 1162 1925 1166 1981
rect 1102 1921 1166 1925
rect 2010 2021 2074 2025
rect 2010 1965 2014 2021
rect 2014 1965 2070 2021
rect 2070 1965 2074 2021
rect 2010 1961 2074 1965
rect 194 1861 258 1865
rect 194 1805 198 1861
rect 198 1805 254 1861
rect 254 1805 258 1861
rect 194 1801 258 1805
rect 1102 1901 1166 1905
rect 1102 1845 1106 1901
rect 1106 1845 1162 1901
rect 1162 1845 1166 1901
rect 2010 1941 2074 1945
rect 2010 1885 2014 1941
rect 2014 1885 2070 1941
rect 2070 1885 2074 1941
rect 2010 1881 2074 1885
rect 1102 1841 1166 1845
rect 194 1781 258 1785
rect 194 1725 198 1781
rect 198 1725 254 1781
rect 254 1725 258 1781
rect 1102 1821 1166 1825
rect 1102 1765 1106 1821
rect 1106 1765 1162 1821
rect 1162 1765 1166 1821
rect 1102 1761 1166 1765
rect 2010 1861 2074 1865
rect 2010 1805 2014 1861
rect 2014 1805 2070 1861
rect 2070 1805 2074 1861
rect 2010 1801 2074 1805
rect 194 1721 258 1725
rect 194 1701 258 1705
rect 194 1645 198 1701
rect 198 1645 254 1701
rect 254 1645 258 1701
rect 194 1641 258 1645
rect 1102 1741 1166 1745
rect 1102 1685 1106 1741
rect 1106 1685 1162 1741
rect 1162 1685 1166 1741
rect 1102 1681 1166 1685
rect 2010 1781 2074 1785
rect 2010 1725 2014 1781
rect 2014 1725 2070 1781
rect 2070 1725 2074 1781
rect 2010 1721 2074 1725
rect 194 1621 258 1625
rect 194 1565 198 1621
rect 198 1565 254 1621
rect 254 1565 258 1621
rect 194 1561 258 1565
rect 1102 1661 1166 1665
rect 1102 1605 1106 1661
rect 1106 1605 1162 1661
rect 1162 1605 1166 1661
rect 2010 1701 2074 1705
rect 2010 1645 2014 1701
rect 2014 1645 2070 1701
rect 2070 1645 2074 1701
rect 2010 1641 2074 1645
rect 1102 1601 1166 1605
rect 194 1541 258 1545
rect 194 1485 198 1541
rect 198 1485 254 1541
rect 254 1485 258 1541
rect 1102 1581 1166 1585
rect 1102 1525 1106 1581
rect 1106 1525 1162 1581
rect 1162 1525 1166 1581
rect 1102 1521 1166 1525
rect 2010 1621 2074 1625
rect 2010 1565 2014 1621
rect 2014 1565 2070 1621
rect 2070 1565 2074 1621
rect 2010 1561 2074 1565
rect 194 1481 258 1485
rect 194 1461 258 1465
rect 194 1405 198 1461
rect 198 1405 254 1461
rect 254 1405 258 1461
rect 194 1401 258 1405
rect 1102 1501 1166 1505
rect 1102 1445 1106 1501
rect 1106 1445 1162 1501
rect 1162 1445 1166 1501
rect 1102 1441 1166 1445
rect 2010 1541 2074 1545
rect 2010 1485 2014 1541
rect 2014 1485 2070 1541
rect 2070 1485 2074 1541
rect 2010 1481 2074 1485
rect 194 1381 258 1385
rect 194 1325 198 1381
rect 198 1325 254 1381
rect 254 1325 258 1381
rect 194 1321 258 1325
rect 1102 1421 1166 1425
rect 1102 1365 1106 1421
rect 1106 1365 1162 1421
rect 1162 1365 1166 1421
rect 2010 1461 2074 1465
rect 2010 1405 2014 1461
rect 2014 1405 2070 1461
rect 2070 1405 2074 1461
rect 2010 1401 2074 1405
rect 1102 1361 1166 1365
rect 194 1301 258 1305
rect 194 1245 198 1301
rect 198 1245 254 1301
rect 254 1245 258 1301
rect 1102 1341 1166 1345
rect 1102 1285 1106 1341
rect 1106 1285 1162 1341
rect 1162 1285 1166 1341
rect 1102 1281 1166 1285
rect 2010 1381 2074 1385
rect 2010 1325 2014 1381
rect 2014 1325 2070 1381
rect 2070 1325 2074 1381
rect 2010 1321 2074 1325
rect 194 1241 258 1245
rect 194 1221 258 1225
rect 194 1165 198 1221
rect 198 1165 254 1221
rect 254 1165 258 1221
rect 194 1161 258 1165
rect 1102 1261 1166 1265
rect 1102 1205 1106 1261
rect 1106 1205 1162 1261
rect 1162 1205 1166 1261
rect 1102 1201 1166 1205
rect 2010 1301 2074 1305
rect 2010 1245 2014 1301
rect 2014 1245 2070 1301
rect 2070 1245 2074 1301
rect 2010 1241 2074 1245
rect 194 1141 258 1145
rect 194 1085 198 1141
rect 198 1085 254 1141
rect 254 1085 258 1141
rect 194 1081 258 1085
rect 325 1181 389 1185
rect 405 1181 469 1185
rect 485 1181 549 1185
rect 565 1181 629 1185
rect 645 1181 709 1185
rect 725 1181 789 1185
rect 805 1181 869 1185
rect 885 1181 949 1185
rect 965 1181 1029 1185
rect 325 1125 380 1181
rect 380 1125 389 1181
rect 405 1125 460 1181
rect 460 1125 469 1181
rect 485 1125 540 1181
rect 540 1125 549 1181
rect 565 1125 620 1181
rect 620 1125 629 1181
rect 645 1125 700 1181
rect 700 1125 709 1181
rect 725 1125 780 1181
rect 780 1125 789 1181
rect 805 1125 860 1181
rect 860 1125 869 1181
rect 885 1125 940 1181
rect 940 1125 949 1181
rect 965 1125 1020 1181
rect 1020 1125 1029 1181
rect 325 1121 389 1125
rect 405 1121 469 1125
rect 485 1121 549 1125
rect 565 1121 629 1125
rect 645 1121 709 1125
rect 725 1121 789 1125
rect 805 1121 869 1125
rect 885 1121 949 1125
rect 965 1121 1029 1125
rect 1102 1181 1166 1185
rect 1102 1125 1106 1181
rect 1106 1125 1162 1181
rect 1162 1125 1166 1181
rect 1102 1121 1166 1125
rect 1239 1181 1303 1185
rect 1319 1181 1383 1185
rect 1399 1181 1463 1185
rect 1479 1181 1543 1185
rect 1559 1181 1623 1185
rect 1639 1181 1703 1185
rect 1719 1181 1783 1185
rect 1799 1181 1863 1185
rect 1879 1181 1943 1185
rect 1239 1125 1248 1181
rect 1248 1125 1303 1181
rect 1319 1125 1328 1181
rect 1328 1125 1383 1181
rect 1399 1125 1408 1181
rect 1408 1125 1463 1181
rect 1479 1125 1488 1181
rect 1488 1125 1543 1181
rect 1559 1125 1568 1181
rect 1568 1125 1623 1181
rect 1639 1125 1648 1181
rect 1648 1125 1703 1181
rect 1719 1125 1728 1181
rect 1728 1125 1783 1181
rect 1799 1125 1808 1181
rect 1808 1125 1863 1181
rect 1879 1125 1888 1181
rect 1888 1125 1943 1181
rect 1239 1121 1303 1125
rect 1319 1121 1383 1125
rect 1399 1121 1463 1125
rect 1479 1121 1543 1125
rect 1559 1121 1623 1125
rect 1639 1121 1703 1125
rect 1719 1121 1783 1125
rect 1799 1121 1863 1125
rect 1879 1121 1943 1125
rect 2010 1221 2074 1225
rect 2010 1165 2014 1221
rect 2014 1165 2070 1221
rect 2070 1165 2074 1221
rect 2010 1161 2074 1165
rect 194 1061 258 1065
rect 194 1005 198 1061
rect 198 1005 254 1061
rect 254 1005 258 1061
rect 194 1001 258 1005
rect 1102 1101 1166 1105
rect 1102 1045 1106 1101
rect 1106 1045 1162 1101
rect 1162 1045 1166 1101
rect 1102 1041 1166 1045
rect 2010 1141 2074 1145
rect 2010 1085 2014 1141
rect 2014 1085 2070 1141
rect 2070 1085 2074 1141
rect 2010 1081 2074 1085
rect 2010 1061 2074 1065
rect 194 981 258 985
rect 194 925 198 981
rect 198 925 254 981
rect 254 925 258 981
rect 194 921 258 925
rect 1102 1021 1166 1025
rect 1102 965 1106 1021
rect 1106 965 1162 1021
rect 1162 965 1166 1021
rect 1102 961 1166 965
rect 2010 1005 2014 1061
rect 2014 1005 2070 1061
rect 2070 1005 2074 1061
rect 2010 1001 2074 1005
rect 1102 941 1166 945
rect 194 901 258 905
rect 194 845 198 901
rect 198 845 254 901
rect 254 845 258 901
rect 194 841 258 845
rect 1102 885 1106 941
rect 1106 885 1162 941
rect 1162 885 1166 941
rect 1102 881 1166 885
rect 2010 981 2074 985
rect 2010 925 2014 981
rect 2014 925 2070 981
rect 2070 925 2074 981
rect 2010 921 2074 925
rect 194 821 258 825
rect 194 765 198 821
rect 198 765 254 821
rect 254 765 258 821
rect 194 761 258 765
rect 1102 861 1166 865
rect 1102 805 1106 861
rect 1106 805 1162 861
rect 1162 805 1166 861
rect 1102 801 1166 805
rect 2010 901 2074 905
rect 2010 845 2014 901
rect 2014 845 2070 901
rect 2070 845 2074 901
rect 2010 841 2074 845
rect 2010 821 2074 825
rect 194 741 258 745
rect 194 685 198 741
rect 198 685 254 741
rect 254 685 258 741
rect 194 681 258 685
rect 1102 781 1166 785
rect 1102 725 1106 781
rect 1106 725 1162 781
rect 1162 725 1166 781
rect 1102 721 1166 725
rect 2010 765 2014 821
rect 2014 765 2070 821
rect 2070 765 2074 821
rect 2010 761 2074 765
rect 1102 701 1166 705
rect 194 661 258 665
rect 194 605 198 661
rect 198 605 254 661
rect 254 605 258 661
rect 194 601 258 605
rect 1102 645 1106 701
rect 1106 645 1162 701
rect 1162 645 1166 701
rect 1102 641 1166 645
rect 2010 741 2074 745
rect 2010 685 2014 741
rect 2014 685 2070 741
rect 2070 685 2074 741
rect 2010 681 2074 685
rect 194 581 258 585
rect 194 525 198 581
rect 198 525 254 581
rect 254 525 258 581
rect 194 521 258 525
rect 1102 621 1166 625
rect 1102 565 1106 621
rect 1106 565 1162 621
rect 1162 565 1166 621
rect 1102 561 1166 565
rect 2010 661 2074 665
rect 2010 605 2014 661
rect 2014 605 2070 661
rect 2070 605 2074 661
rect 2010 601 2074 605
rect 2010 581 2074 585
rect 194 501 258 505
rect 194 445 198 501
rect 198 445 254 501
rect 254 445 258 501
rect 194 441 258 445
rect 1102 541 1166 545
rect 1102 485 1106 541
rect 1106 485 1162 541
rect 1162 485 1166 541
rect 1102 481 1166 485
rect 2010 525 2014 581
rect 2014 525 2070 581
rect 2070 525 2074 581
rect 2010 521 2074 525
rect 1102 461 1166 465
rect 194 421 258 425
rect 194 365 198 421
rect 198 365 254 421
rect 254 365 258 421
rect 194 361 258 365
rect 1102 405 1106 461
rect 1106 405 1162 461
rect 1162 405 1166 461
rect 1102 401 1166 405
rect 2010 501 2074 505
rect 2010 445 2014 501
rect 2014 445 2070 501
rect 2070 445 2074 501
rect 2010 441 2074 445
rect 194 341 258 345
rect 194 285 198 341
rect 198 285 254 341
rect 254 285 258 341
rect 194 281 258 285
rect 1102 381 1166 385
rect 1102 325 1106 381
rect 1106 325 1162 381
rect 1162 325 1166 381
rect 1102 321 1166 325
rect 2010 421 2074 425
rect 2010 365 2014 421
rect 2014 365 2070 421
rect 2070 365 2074 421
rect 2010 361 2074 365
rect 2010 341 2074 345
rect 194 201 258 265
rect 1102 301 1166 305
rect 1102 245 1106 301
rect 1106 245 1162 301
rect 1162 245 1166 301
rect 1102 241 1166 245
rect 2010 285 2014 341
rect 2014 285 2070 341
rect 2070 285 2074 341
rect 2010 281 2074 285
rect 1102 221 1166 225
rect 194 121 258 185
rect 1102 165 1106 221
rect 1106 165 1162 221
rect 1162 165 1166 221
rect 1102 161 1166 165
rect 2010 201 2074 265
rect 2010 121 2074 185
rect 262 35 326 99
rect 342 35 406 99
rect 422 35 486 99
rect 502 35 566 99
rect 582 35 646 99
rect 662 35 726 99
rect 742 35 806 99
rect 822 35 886 99
rect 902 35 966 99
rect 982 35 1046 99
rect 1062 35 1126 99
rect 1142 35 1206 99
rect 1222 35 1286 99
rect 1302 35 1366 99
rect 1382 35 1446 99
rect 1462 35 1526 99
rect 1542 35 1606 99
rect 1622 35 1686 99
rect 1702 35 1766 99
rect 1782 35 1846 99
rect 1862 35 1926 99
rect 1942 35 2006 99
rect 2143 2300 2207 2304
rect 2143 2244 2147 2300
rect 2147 2244 2203 2300
rect 2203 2244 2207 2300
rect 2143 2240 2207 2244
rect 2143 2220 2207 2224
rect 2143 2164 2147 2220
rect 2147 2164 2203 2220
rect 2203 2164 2207 2220
rect 2143 2160 2207 2164
rect 2143 2140 2207 2144
rect 2143 2084 2147 2140
rect 2147 2084 2203 2140
rect 2203 2084 2207 2140
rect 2143 2080 2207 2084
rect 2143 2060 2207 2064
rect 2143 2004 2147 2060
rect 2147 2004 2203 2060
rect 2203 2004 2207 2060
rect 2143 2000 2207 2004
rect 2143 1980 2207 1984
rect 2143 1924 2147 1980
rect 2147 1924 2203 1980
rect 2203 1924 2207 1980
rect 2143 1920 2207 1924
rect 2143 1900 2207 1904
rect 2143 1844 2147 1900
rect 2147 1844 2203 1900
rect 2203 1844 2207 1900
rect 2143 1840 2207 1844
rect 2143 1820 2207 1824
rect 2143 1764 2147 1820
rect 2147 1764 2203 1820
rect 2203 1764 2207 1820
rect 2143 1760 2207 1764
rect 2143 1740 2207 1744
rect 2143 1684 2147 1740
rect 2147 1684 2203 1740
rect 2203 1684 2207 1740
rect 2143 1680 2207 1684
rect 2143 1660 2207 1664
rect 2143 1604 2147 1660
rect 2147 1604 2203 1660
rect 2203 1604 2207 1660
rect 2143 1600 2207 1604
rect 2143 1580 2207 1584
rect 2143 1524 2147 1580
rect 2147 1524 2203 1580
rect 2203 1524 2207 1580
rect 2143 1520 2207 1524
rect 2143 1500 2207 1504
rect 2143 1444 2147 1500
rect 2147 1444 2203 1500
rect 2203 1444 2207 1500
rect 2143 1440 2207 1444
rect 2143 1420 2207 1424
rect 2143 1364 2147 1420
rect 2147 1364 2203 1420
rect 2203 1364 2207 1420
rect 2143 1360 2207 1364
rect 2143 1340 2207 1344
rect 2143 1284 2147 1340
rect 2147 1284 2203 1340
rect 2203 1284 2207 1340
rect 2143 1280 2207 1284
rect 2143 1260 2207 1264
rect 2143 1204 2147 1260
rect 2147 1204 2203 1260
rect 2203 1204 2207 1260
rect 2143 1200 2207 1204
rect 2143 1180 2207 1184
rect 2143 1124 2147 1180
rect 2147 1124 2203 1180
rect 2203 1124 2207 1180
rect 2143 1120 2207 1124
rect 2143 1100 2207 1104
rect 2143 1044 2147 1100
rect 2147 1044 2203 1100
rect 2203 1044 2207 1100
rect 2143 1040 2207 1044
rect 2143 1020 2207 1024
rect 2143 964 2147 1020
rect 2147 964 2203 1020
rect 2203 964 2207 1020
rect 2143 960 2207 964
rect 2143 940 2207 944
rect 2143 884 2147 940
rect 2147 884 2203 940
rect 2203 884 2207 940
rect 2143 880 2207 884
rect 2143 860 2207 864
rect 2143 804 2147 860
rect 2147 804 2203 860
rect 2203 804 2207 860
rect 2143 800 2207 804
rect 2143 780 2207 784
rect 2143 724 2147 780
rect 2147 724 2203 780
rect 2203 724 2207 780
rect 2143 720 2207 724
rect 2143 700 2207 704
rect 2143 644 2147 700
rect 2147 644 2203 700
rect 2203 644 2207 700
rect 2143 640 2207 644
rect 2143 620 2207 624
rect 2143 564 2147 620
rect 2147 564 2203 620
rect 2203 564 2207 620
rect 2143 560 2207 564
rect 2143 540 2207 544
rect 2143 484 2147 540
rect 2147 484 2203 540
rect 2203 484 2207 540
rect 2143 480 2207 484
rect 2143 460 2207 464
rect 2143 404 2147 460
rect 2147 404 2203 460
rect 2203 404 2207 460
rect 2143 400 2207 404
rect 2143 380 2207 384
rect 2143 324 2147 380
rect 2147 324 2203 380
rect 2203 324 2207 380
rect 2143 320 2207 324
rect 2143 300 2207 304
rect 2143 244 2147 300
rect 2147 244 2203 300
rect 2203 244 2207 300
rect 2143 240 2207 244
rect 2143 220 2207 224
rect 2143 164 2147 220
rect 2147 164 2203 220
rect 2203 164 2207 220
rect 2143 160 2207 164
rect 2143 140 2207 144
rect 2143 84 2147 140
rect 2147 84 2203 140
rect 2203 84 2207 140
rect 2143 80 2207 84
<< metal4 >>
rect 60 2304 126 2323
rect 60 2240 61 2304
rect 125 2240 126 2304
rect 2142 2304 2208 2323
rect 60 2224 126 2240
rect 60 2160 61 2224
rect 125 2160 126 2224
rect 60 2144 126 2160
rect 60 2080 61 2144
rect 125 2080 126 2144
rect 60 2064 126 2080
rect 60 2000 61 2064
rect 125 2000 126 2064
rect 60 1984 126 2000
rect 60 1920 61 1984
rect 125 1920 126 1984
rect 60 1904 126 1920
rect 60 1840 61 1904
rect 125 1840 126 1904
rect 60 1824 126 1840
rect 60 1760 61 1824
rect 125 1760 126 1824
rect 60 1744 126 1760
rect 60 1680 61 1744
rect 125 1680 126 1744
rect 60 1664 126 1680
rect 60 1600 61 1664
rect 125 1600 126 1664
rect 60 1584 126 1600
rect 60 1520 61 1584
rect 125 1520 126 1584
rect 60 1504 126 1520
rect 60 1440 61 1504
rect 125 1440 126 1504
rect 60 1424 126 1440
rect 60 1360 61 1424
rect 125 1360 126 1424
rect 60 1344 126 1360
rect 60 1280 61 1344
rect 125 1280 126 1344
rect 60 1264 126 1280
rect 60 1200 61 1264
rect 125 1200 126 1264
rect 60 1184 126 1200
rect 60 1120 61 1184
rect 125 1120 126 1184
rect 60 1104 126 1120
rect 60 1040 61 1104
rect 125 1040 126 1104
rect 60 1024 126 1040
rect 60 960 61 1024
rect 125 960 126 1024
rect 60 944 126 960
rect 60 880 61 944
rect 125 880 126 944
rect 60 864 126 880
rect 60 800 61 864
rect 125 800 126 864
rect 60 784 126 800
rect 60 720 61 784
rect 125 720 126 784
rect 60 704 126 720
rect 60 640 61 704
rect 125 640 126 704
rect 60 624 126 640
rect 60 560 61 624
rect 125 560 126 624
rect 60 544 126 560
rect 60 480 61 544
rect 125 480 126 544
rect 60 464 126 480
rect 60 400 61 464
rect 125 400 126 464
rect 60 384 126 400
rect 60 320 61 384
rect 125 320 126 384
rect 60 304 126 320
rect 60 240 61 304
rect 125 240 126 304
rect 60 224 126 240
rect 60 160 61 224
rect 125 160 126 224
rect 60 144 126 160
rect 60 80 61 144
rect 125 80 126 144
rect 60 15 126 80
rect 193 2271 2009 2272
rect 193 2207 262 2271
rect 326 2207 342 2271
rect 406 2207 422 2271
rect 486 2207 502 2271
rect 566 2207 582 2271
rect 646 2207 662 2271
rect 726 2207 742 2271
rect 806 2207 822 2271
rect 886 2207 902 2271
rect 966 2207 982 2271
rect 1046 2207 1062 2271
rect 1126 2207 1142 2271
rect 1206 2207 1222 2271
rect 1286 2207 1302 2271
rect 1366 2207 1382 2271
rect 1446 2207 1462 2271
rect 1526 2207 1542 2271
rect 1606 2207 1622 2271
rect 1686 2207 1702 2271
rect 1766 2207 1782 2271
rect 1846 2207 1862 2271
rect 1926 2207 1942 2271
rect 2006 2266 2009 2271
rect 2006 2207 2075 2266
rect 193 2206 2075 2207
rect 193 2185 259 2206
rect 193 2121 194 2185
rect 258 2121 259 2185
rect 193 2105 259 2121
rect 193 2041 194 2105
rect 258 2041 259 2105
rect 193 2025 259 2041
rect 193 1961 194 2025
rect 258 1961 259 2025
rect 193 1945 259 1961
rect 193 1881 194 1945
rect 258 1881 259 1945
rect 193 1865 259 1881
rect 193 1801 194 1865
rect 258 1801 259 1865
rect 193 1785 259 1801
rect 193 1721 194 1785
rect 258 1721 259 1785
rect 193 1705 259 1721
rect 193 1641 194 1705
rect 258 1641 259 1705
rect 193 1625 259 1641
rect 193 1561 194 1625
rect 258 1561 259 1625
rect 193 1545 259 1561
rect 193 1481 194 1545
rect 258 1481 259 1545
rect 193 1465 259 1481
rect 193 1401 194 1465
rect 258 1401 259 1465
rect 193 1385 259 1401
rect 193 1321 194 1385
rect 258 1321 259 1385
rect 193 1305 259 1321
rect 193 1241 194 1305
rect 258 1241 259 1305
rect 193 1225 259 1241
rect 193 1161 194 1225
rect 258 1161 259 1225
rect 193 1145 259 1161
rect 193 1081 194 1145
rect 258 1081 259 1145
rect 193 1065 259 1081
rect 193 1001 194 1065
rect 258 1001 259 1065
rect 193 985 259 1001
rect 193 921 194 985
rect 258 921 259 985
rect 193 905 259 921
rect 193 841 194 905
rect 258 841 259 905
rect 193 825 259 841
rect 193 761 194 825
rect 258 761 259 825
rect 193 745 259 761
rect 193 681 194 745
rect 258 681 259 745
rect 193 665 259 681
rect 193 601 194 665
rect 258 601 259 665
rect 193 585 259 601
rect 193 521 194 585
rect 258 521 259 585
rect 193 505 259 521
rect 193 441 194 505
rect 258 441 259 505
rect 193 425 259 441
rect 193 361 194 425
rect 258 361 259 425
rect 193 345 259 361
rect 193 281 194 345
rect 258 281 259 345
rect 193 265 259 281
rect 193 201 194 265
rect 258 201 259 265
rect 193 185 259 201
rect 193 121 194 185
rect 258 121 259 185
rect 319 1186 379 2146
rect 439 1246 499 2206
rect 559 1186 619 2146
rect 679 1246 739 2206
rect 799 1186 859 2146
rect 919 1246 1002 2206
rect 1062 2145 1167 2146
rect 1062 2081 1102 2145
rect 1166 2081 1167 2145
rect 1062 2065 1167 2081
rect 1062 2001 1102 2065
rect 1166 2001 1167 2065
rect 1062 1985 1167 2001
rect 1062 1921 1102 1985
rect 1166 1921 1167 1985
rect 1062 1905 1167 1921
rect 1062 1841 1102 1905
rect 1166 1841 1167 1905
rect 1062 1825 1167 1841
rect 1062 1761 1102 1825
rect 1166 1761 1167 1825
rect 1062 1745 1167 1761
rect 1062 1681 1102 1745
rect 1166 1681 1167 1745
rect 1062 1665 1167 1681
rect 1062 1601 1102 1665
rect 1166 1601 1167 1665
rect 1062 1585 1167 1601
rect 1062 1521 1102 1585
rect 1166 1521 1167 1585
rect 1062 1505 1167 1521
rect 1062 1441 1102 1505
rect 1166 1441 1167 1505
rect 1062 1425 1167 1441
rect 1062 1361 1102 1425
rect 1166 1361 1167 1425
rect 1062 1345 1167 1361
rect 1062 1281 1102 1345
rect 1166 1281 1167 1345
rect 1062 1265 1167 1281
rect 1062 1201 1102 1265
rect 1166 1201 1167 1265
rect 1227 1246 1349 2206
rect 1062 1186 1167 1201
rect 1409 1186 1469 2146
rect 1529 1246 1589 2206
rect 1649 1186 1709 2146
rect 1769 1246 1829 2206
rect 2009 2185 2075 2206
rect 1889 1186 1949 2146
rect 319 1185 1949 1186
rect 319 1121 325 1185
rect 389 1121 405 1185
rect 469 1121 485 1185
rect 549 1121 565 1185
rect 629 1121 645 1185
rect 709 1121 725 1185
rect 789 1121 805 1185
rect 869 1121 885 1185
rect 949 1121 965 1185
rect 1029 1121 1102 1185
rect 1166 1121 1239 1185
rect 1303 1121 1319 1185
rect 1383 1121 1399 1185
rect 1463 1121 1479 1185
rect 1543 1121 1559 1185
rect 1623 1121 1639 1185
rect 1703 1121 1719 1185
rect 1783 1121 1799 1185
rect 1863 1121 1879 1185
rect 1943 1121 1949 1185
rect 319 1120 1949 1121
rect 319 160 379 1120
rect 193 100 259 121
rect 439 100 499 1060
rect 559 160 619 1120
rect 679 100 739 1060
rect 799 160 859 1120
rect 1062 1105 1167 1120
rect 919 100 1002 1060
rect 1062 1041 1102 1105
rect 1166 1041 1167 1105
rect 1062 1025 1167 1041
rect 1062 961 1102 1025
rect 1166 961 1167 1025
rect 1062 945 1167 961
rect 1062 881 1102 945
rect 1166 881 1167 945
rect 1062 865 1167 881
rect 1062 801 1102 865
rect 1166 801 1167 865
rect 1062 785 1167 801
rect 1062 721 1102 785
rect 1166 721 1167 785
rect 1062 705 1167 721
rect 1062 641 1102 705
rect 1166 641 1167 705
rect 1062 625 1167 641
rect 1062 561 1102 625
rect 1166 561 1167 625
rect 1062 545 1167 561
rect 1062 481 1102 545
rect 1166 481 1167 545
rect 1062 465 1167 481
rect 1062 401 1102 465
rect 1166 401 1167 465
rect 1062 385 1167 401
rect 1062 321 1102 385
rect 1166 321 1167 385
rect 1062 305 1167 321
rect 1062 241 1102 305
rect 1166 241 1167 305
rect 1062 225 1167 241
rect 1062 161 1102 225
rect 1166 161 1167 225
rect 1062 160 1167 161
rect 1227 100 1349 1060
rect 1409 160 1469 1120
rect 1529 100 1589 1060
rect 1649 160 1709 1120
rect 1769 100 1829 1060
rect 1889 160 1949 1120
rect 2009 2121 2010 2185
rect 2074 2121 2075 2185
rect 2009 2105 2075 2121
rect 2009 2041 2010 2105
rect 2074 2041 2075 2105
rect 2009 2025 2075 2041
rect 2009 1961 2010 2025
rect 2074 1961 2075 2025
rect 2009 1945 2075 1961
rect 2009 1881 2010 1945
rect 2074 1881 2075 1945
rect 2009 1865 2075 1881
rect 2009 1801 2010 1865
rect 2074 1801 2075 1865
rect 2009 1785 2075 1801
rect 2009 1721 2010 1785
rect 2074 1721 2075 1785
rect 2009 1705 2075 1721
rect 2009 1641 2010 1705
rect 2074 1641 2075 1705
rect 2009 1625 2075 1641
rect 2009 1561 2010 1625
rect 2074 1561 2075 1625
rect 2009 1545 2075 1561
rect 2009 1481 2010 1545
rect 2074 1481 2075 1545
rect 2009 1465 2075 1481
rect 2009 1401 2010 1465
rect 2074 1401 2075 1465
rect 2009 1385 2075 1401
rect 2009 1321 2010 1385
rect 2074 1321 2075 1385
rect 2009 1305 2075 1321
rect 2009 1241 2010 1305
rect 2074 1241 2075 1305
rect 2009 1225 2075 1241
rect 2009 1161 2010 1225
rect 2074 1161 2075 1225
rect 2009 1145 2075 1161
rect 2009 1081 2010 1145
rect 2074 1081 2075 1145
rect 2009 1065 2075 1081
rect 2009 1001 2010 1065
rect 2074 1001 2075 1065
rect 2009 985 2075 1001
rect 2009 921 2010 985
rect 2074 921 2075 985
rect 2009 905 2075 921
rect 2009 841 2010 905
rect 2074 841 2075 905
rect 2009 825 2075 841
rect 2009 761 2010 825
rect 2074 761 2075 825
rect 2009 745 2075 761
rect 2009 681 2010 745
rect 2074 681 2075 745
rect 2009 665 2075 681
rect 2009 601 2010 665
rect 2074 601 2075 665
rect 2009 585 2075 601
rect 2009 521 2010 585
rect 2074 521 2075 585
rect 2009 505 2075 521
rect 2009 441 2010 505
rect 2074 441 2075 505
rect 2009 425 2075 441
rect 2009 361 2010 425
rect 2074 361 2075 425
rect 2009 345 2075 361
rect 2009 281 2010 345
rect 2074 281 2075 345
rect 2009 265 2075 281
rect 2009 201 2010 265
rect 2074 201 2075 265
rect 2009 185 2075 201
rect 2009 121 2010 185
rect 2074 121 2075 185
rect 2009 100 2075 121
rect 193 99 2075 100
rect 193 35 262 99
rect 326 35 342 99
rect 406 35 422 99
rect 486 35 502 99
rect 566 35 582 99
rect 646 35 662 99
rect 726 35 742 99
rect 806 35 822 99
rect 886 35 902 99
rect 966 35 982 99
rect 1046 35 1062 99
rect 1126 35 1142 99
rect 1206 35 1222 99
rect 1286 35 1302 99
rect 1366 35 1382 99
rect 1446 35 1462 99
rect 1526 35 1542 99
rect 1606 35 1622 99
rect 1686 35 1702 99
rect 1766 35 1782 99
rect 1846 35 1862 99
rect 1926 35 1942 99
rect 2006 35 2075 99
rect 193 34 2075 35
rect 2142 2240 2143 2304
rect 2207 2240 2208 2304
rect 2142 2224 2208 2240
rect 2142 2160 2143 2224
rect 2207 2160 2208 2224
rect 2142 2144 2208 2160
rect 2142 2080 2143 2144
rect 2207 2080 2208 2144
rect 2142 2064 2208 2080
rect 2142 2000 2143 2064
rect 2207 2000 2208 2064
rect 2142 1984 2208 2000
rect 2142 1920 2143 1984
rect 2207 1920 2208 1984
rect 2142 1904 2208 1920
rect 2142 1840 2143 1904
rect 2207 1840 2208 1904
rect 2142 1824 2208 1840
rect 2142 1760 2143 1824
rect 2207 1760 2208 1824
rect 2142 1744 2208 1760
rect 2142 1680 2143 1744
rect 2207 1680 2208 1744
rect 2142 1664 2208 1680
rect 2142 1600 2143 1664
rect 2207 1600 2208 1664
rect 2142 1584 2208 1600
rect 2142 1520 2143 1584
rect 2207 1520 2208 1584
rect 2142 1504 2208 1520
rect 2142 1440 2143 1504
rect 2207 1440 2208 1504
rect 2142 1424 2208 1440
rect 2142 1360 2143 1424
rect 2207 1360 2208 1424
rect 2142 1344 2208 1360
rect 2142 1280 2143 1344
rect 2207 1280 2208 1344
rect 2142 1264 2208 1280
rect 2142 1200 2143 1264
rect 2207 1200 2208 1264
rect 2142 1184 2208 1200
rect 2142 1120 2143 1184
rect 2207 1120 2208 1184
rect 2142 1104 2208 1120
rect 2142 1040 2143 1104
rect 2207 1040 2208 1104
rect 2142 1024 2208 1040
rect 2142 960 2143 1024
rect 2207 960 2208 1024
rect 2142 944 2208 960
rect 2142 880 2143 944
rect 2207 880 2208 944
rect 2142 864 2208 880
rect 2142 800 2143 864
rect 2207 800 2208 864
rect 2142 784 2208 800
rect 2142 720 2143 784
rect 2207 720 2208 784
rect 2142 704 2208 720
rect 2142 640 2143 704
rect 2207 640 2208 704
rect 2142 624 2208 640
rect 2142 560 2143 624
rect 2207 560 2208 624
rect 2142 544 2208 560
rect 2142 480 2143 544
rect 2207 480 2208 544
rect 2142 464 2208 480
rect 2142 400 2143 464
rect 2207 400 2208 464
rect 2142 384 2208 400
rect 2142 320 2143 384
rect 2207 320 2208 384
rect 2142 304 2208 320
rect 2142 240 2143 304
rect 2207 240 2208 304
rect 2142 224 2208 240
rect 2142 160 2143 224
rect 2207 160 2208 224
rect 2142 144 2208 160
rect 2142 80 2143 144
rect 2207 80 2208 144
rect 2142 15 2208 80
<< metal5 >>
rect 0 0 2268 2338
<< labels >>
flabel metal1 s 145 2287 175 2315 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel metal2 s 156 2223 198 2259 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel comment s 1037 1548 1037 1548 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1436 1037 1436 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1324 1037 1324 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1772 1037 1772 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1660 1037 1660 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1940 1037 1940 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1828 1037 1828 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1716 1037 1716 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1604 1037 1604 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1492 1037 1492 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1380 1037 1380 0 FreeSans 200 90 0 0 A
flabel comment s 1037 1268 1037 1268 0 FreeSans 200 90 0 0 A
flabel comment s 277 1881 277 1881 0 FreeSans 200 90 0 0 B
flabel comment s 277 1769 277 1769 0 FreeSans 200 90 0 0 B
flabel comment s 277 1657 277 1657 0 FreeSans 200 90 0 0 B
flabel comment s 277 1545 277 1545 0 FreeSans 200 90 0 0 B
flabel comment s 277 1433 277 1433 0 FreeSans 200 90 0 0 B
flabel comment s 277 1321 277 1321 0 FreeSans 200 90 0 0 B
flabel comment s 1037 1884 1037 1884 0 FreeSans 200 90 0 0 A
flabel comment s 1612 1972 1612 1972 0 FreeSans 200 270 0 0 B
flabel comment s 1332 1972 1332 1972 0 FreeSans 200 270 0 0 B
flabel comment s 1472 1972 1472 1972 0 FreeSans 200 270 0 0 B
flabel comment s 1892 1972 1892 1972 0 FreeSans 200 270 0 0 B
flabel comment s 1752 1972 1752 1972 0 FreeSans 200 270 0 0 B
flabel comment s 1822 1228 1822 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1402 1228 1402 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1962 1228 1962 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1262 1228 1262 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1542 1228 1542 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1682 1228 1682 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1991 1268 1991 1268 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1380 1991 1380 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1492 1991 1492 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1604 1991 1604 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1716 1991 1716 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1828 1991 1828 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1940 1991 1940 0 FreeSans 200 90 0 0 B
flabel comment s 1231 1884 1231 1884 0 FreeSans 200 90 0 0 A
flabel comment s 1991 1321 1991 1321 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1433 1991 1433 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1545 1991 1545 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1657 1991 1657 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1769 1991 1769 0 FreeSans 200 90 0 0 B
flabel comment s 1991 1881 1991 1881 0 FreeSans 200 90 0 0 B
flabel comment s 1231 1268 1231 1268 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1380 1231 1380 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1492 1231 1492 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1604 1231 1604 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1716 1231 1716 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1828 1231 1828 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1940 1231 1940 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1660 1231 1660 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1772 1231 1772 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1324 1231 1324 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1436 1231 1436 0 FreeSans 200 90 0 0 A
flabel comment s 1231 1548 1231 1548 0 FreeSans 200 90 0 0 A
flabel comment s 656 340 656 340 0 FreeSans 200 90 0 0 B
flabel comment s 936 340 936 340 0 FreeSans 200 90 0 0 B
flabel comment s 796 340 796 340 0 FreeSans 200 90 0 0 B
flabel comment s 376 340 376 340 0 FreeSans 200 90 0 0 B
flabel comment s 516 340 516 340 0 FreeSans 200 90 0 0 B
flabel comment s 446 1084 446 1084 0 FreeSans 200 270 0 0 A
flabel comment s 866 1084 866 1084 0 FreeSans 200 270 0 0 A
flabel comment s 306 1084 306 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1006 1084 1006 1084 0 FreeSans 200 270 0 0 A
flabel comment s 726 1084 726 1084 0 FreeSans 200 270 0 0 A
flabel comment s 586 1084 586 1084 0 FreeSans 200 270 0 0 A
flabel comment s 277 1044 277 1044 0 FreeSans 200 270 0 0 B
flabel comment s 277 932 277 932 0 FreeSans 200 270 0 0 B
flabel comment s 277 820 277 820 0 FreeSans 200 270 0 0 B
flabel comment s 277 708 277 708 0 FreeSans 200 270 0 0 B
flabel comment s 277 596 277 596 0 FreeSans 200 270 0 0 B
flabel comment s 277 484 277 484 0 FreeSans 200 270 0 0 B
flabel comment s 277 372 277 372 0 FreeSans 200 270 0 0 B
flabel comment s 1037 428 1037 428 0 FreeSans 200 270 0 0 A
flabel comment s 277 991 277 991 0 FreeSans 200 270 0 0 B
flabel comment s 277 879 277 879 0 FreeSans 200 270 0 0 B
flabel comment s 277 767 277 767 0 FreeSans 200 270 0 0 B
flabel comment s 277 655 277 655 0 FreeSans 200 270 0 0 B
flabel comment s 277 543 277 543 0 FreeSans 200 270 0 0 B
flabel comment s 277 431 277 431 0 FreeSans 200 270 0 0 B
flabel comment s 1037 1044 1037 1044 0 FreeSans 200 270 0 0 A
flabel comment s 1037 932 1037 932 0 FreeSans 200 270 0 0 A
flabel comment s 1037 820 1037 820 0 FreeSans 200 270 0 0 A
flabel comment s 1037 708 1037 708 0 FreeSans 200 270 0 0 A
flabel comment s 1037 596 1037 596 0 FreeSans 200 270 0 0 A
flabel comment s 1037 484 1037 484 0 FreeSans 200 270 0 0 A
flabel comment s 1037 372 1037 372 0 FreeSans 200 270 0 0 A
flabel comment s 1037 652 1037 652 0 FreeSans 200 270 0 0 A
flabel comment s 1037 540 1037 540 0 FreeSans 200 270 0 0 A
flabel comment s 1037 988 1037 988 0 FreeSans 200 270 0 0 A
flabel comment s 1037 876 1037 876 0 FreeSans 200 270 0 0 A
flabel comment s 1037 764 1037 764 0 FreeSans 200 270 0 0 A
flabel comment s 1612 340 1612 340 0 FreeSans 200 90 0 0 B
flabel comment s 1332 340 1332 340 0 FreeSans 200 90 0 0 B
flabel comment s 1472 340 1472 340 0 FreeSans 200 90 0 0 B
flabel comment s 1892 340 1892 340 0 FreeSans 200 90 0 0 B
flabel comment s 1752 340 1752 340 0 FreeSans 200 90 0 0 B
flabel comment s 1822 1084 1822 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1402 1084 1402 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1962 1084 1962 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1262 1084 1262 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1542 1084 1542 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1682 1084 1682 1084 0 FreeSans 200 270 0 0 A
flabel comment s 1991 1044 1991 1044 0 FreeSans 200 270 0 0 B
flabel comment s 1991 932 1991 932 0 FreeSans 200 270 0 0 B
flabel comment s 1991 820 1991 820 0 FreeSans 200 270 0 0 B
flabel comment s 1991 708 1991 708 0 FreeSans 200 270 0 0 B
flabel comment s 1991 596 1991 596 0 FreeSans 200 270 0 0 B
flabel comment s 1991 484 1991 484 0 FreeSans 200 270 0 0 B
flabel comment s 1991 372 1991 372 0 FreeSans 200 270 0 0 B
flabel comment s 1231 428 1231 428 0 FreeSans 200 270 0 0 A
flabel comment s 1991 991 1991 991 0 FreeSans 200 270 0 0 B
flabel comment s 1991 879 1991 879 0 FreeSans 200 270 0 0 B
flabel comment s 1991 767 1991 767 0 FreeSans 200 270 0 0 B
flabel comment s 1991 655 1991 655 0 FreeSans 200 270 0 0 B
flabel comment s 1991 543 1991 543 0 FreeSans 200 270 0 0 B
flabel comment s 1991 431 1991 431 0 FreeSans 200 270 0 0 B
flabel comment s 1231 1044 1231 1044 0 FreeSans 200 270 0 0 A
flabel comment s 1231 932 1231 932 0 FreeSans 200 270 0 0 A
flabel comment s 1231 820 1231 820 0 FreeSans 200 270 0 0 A
flabel comment s 1231 708 1231 708 0 FreeSans 200 270 0 0 A
flabel comment s 1231 596 1231 596 0 FreeSans 200 270 0 0 A
flabel comment s 1231 484 1231 484 0 FreeSans 200 270 0 0 A
flabel comment s 1231 372 1231 372 0 FreeSans 200 270 0 0 A
flabel comment s 1231 652 1231 652 0 FreeSans 200 270 0 0 A
flabel comment s 1231 540 1231 540 0 FreeSans 200 270 0 0 A
flabel comment s 1231 988 1231 988 0 FreeSans 200 270 0 0 A
flabel comment s 1231 876 1231 876 0 FreeSans 200 270 0 0 A
flabel comment s 1231 764 1231 764 0 FreeSans 200 270 0 0 A
flabel comment s 2094 1156 2094 1156 0 FreeSans 300 0 0 0 S
flabel comment s 1134 1150 1134 1150 0 FreeSans 300 0 0 0 D
flabel comment s 174 1156 174 1156 0 FreeSans 300 0 0 0 S
flabel comment s 277 1940 277 1940 0 FreeSans 200 90 0 0 B
flabel comment s 277 1828 277 1828 0 FreeSans 200 90 0 0 B
flabel comment s 277 1716 277 1716 0 FreeSans 200 90 0 0 B
flabel comment s 277 1604 277 1604 0 FreeSans 200 90 0 0 B
flabel comment s 277 1492 277 1492 0 FreeSans 200 90 0 0 B
flabel comment s 277 1380 277 1380 0 FreeSans 200 90 0 0 B
flabel comment s 277 1268 277 1268 0 FreeSans 200 90 0 0 B
flabel comment s 586 1228 586 1228 0 FreeSans 200 90 0 0 A
flabel comment s 726 1228 726 1228 0 FreeSans 200 90 0 0 A
flabel comment s 1006 1228 1006 1228 0 FreeSans 200 90 0 0 A
flabel comment s 306 1228 306 1228 0 FreeSans 200 90 0 0 A
flabel comment s 866 1228 866 1228 0 FreeSans 200 90 0 0 A
flabel comment s 446 1228 446 1228 0 FreeSans 200 90 0 0 A
flabel comment s 516 1972 516 1972 0 FreeSans 200 270 0 0 B
flabel comment s 376 1972 376 1972 0 FreeSans 200 270 0 0 B
flabel comment s 796 1972 796 1972 0 FreeSans 200 270 0 0 B
flabel comment s 936 1972 936 1972 0 FreeSans 200 270 0 0 B
flabel comment s 656 1972 656 1972 0 FreeSans 200 270 0 0 B
flabel comment s 1196 2309 1196 2309 0 FreeSans 280 180 0 0 FOR TILE ALIGMENT USE Y OFFSET OF 11.54
flabel comment s 93 1157 93 1157 0 FreeSans 500 90 0 0 FOR TILE ALIGNMENT USE X OFFSET OF 10.41
flabel comment s 2175 1157 2175 1157 0 FreeSans 500 90 0 0 FOR TILE ALIGNMENT USE X OFFSET OF 10.41
flabel comment s 1196 1 1196 1 0 FreeSans 280 180 0 0 FOR TILE ALIGMENT USE Y OFFSET OF 11.54
flabel metal5 s 1578 590 1665 685 0 FreeSans 200 0 0 0 MET5
port 4 nsew
<< properties >>
string GDS_END 441236
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 337490
string path 6.775 56.350 49.925 56.350 
string device primitive
<< end >>
