magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 157 439 203
rect 1538 157 2006 203
rect 1 21 2006 157
rect 30 -17 64 21
<< locali >>
rect 103 317 169 489
rect 287 390 329 493
rect 280 356 329 390
rect 280 317 314 356
rect 17 283 314 317
rect 650 314 868 348
rect 17 181 87 283
rect 17 147 305 181
rect 103 51 169 147
rect 271 97 305 147
rect 650 255 684 314
rect 610 221 684 255
rect 834 250 868 314
rect 1319 337 1369 391
rect 1044 303 1369 337
rect 1044 287 1116 303
rect 1044 250 1078 287
rect 1319 271 1369 303
rect 1664 393 1698 493
rect 1664 359 1714 393
rect 834 193 1078 250
rect 1680 317 1714 359
rect 1832 317 1898 485
rect 1680 283 2007 317
rect 271 63 337 97
rect 1940 181 2007 283
rect 1680 147 2007 181
rect 1680 97 1730 147
rect 1664 51 1730 97
rect 1832 54 1898 147
<< obsli1 >>
rect 0 527 2024 561
rect 35 359 69 527
rect 203 359 237 527
rect 363 455 429 527
rect 547 416 634 493
rect 428 382 634 416
rect 668 421 702 493
rect 736 455 802 527
rect 836 421 883 493
rect 668 387 883 421
rect 924 383 990 527
rect 1024 421 1058 493
rect 1092 455 1158 527
rect 1192 421 1226 493
rect 1282 425 1522 493
rect 1563 455 1629 527
rect 1024 387 1226 421
rect 1488 421 1522 425
rect 428 333 462 382
rect 355 320 462 333
rect 348 299 462 320
rect 348 286 389 299
rect 496 289 616 338
rect 348 249 382 286
rect 121 215 382 249
rect 35 17 69 113
rect 203 17 237 113
rect 348 165 382 215
rect 416 255 468 265
rect 416 199 536 255
rect 722 206 800 272
rect 916 287 999 349
rect 1488 387 1621 421
rect 1415 289 1552 347
rect 1587 328 1621 387
rect 1748 359 1782 527
rect 1587 294 1645 328
rect 1129 191 1201 255
rect 1235 191 1372 225
rect 1406 199 1577 255
rect 1611 249 1645 294
rect 1932 359 1966 527
rect 1611 215 1889 249
rect 570 165 618 187
rect 348 131 618 165
rect 371 17 437 93
rect 474 51 618 131
rect 668 123 870 157
rect 668 51 702 123
rect 736 17 802 89
rect 836 51 870 123
rect 1024 123 1226 157
rect 1269 153 1372 191
rect 1611 165 1645 215
rect 924 17 990 98
rect 1024 51 1058 123
rect 1092 17 1158 89
rect 1192 51 1226 123
rect 1461 131 1645 165
rect 1293 101 1327 119
rect 1461 101 1495 131
rect 1293 51 1495 101
rect 1541 17 1607 89
rect 1764 17 1798 113
rect 1932 17 1966 113
rect 0 -17 2024 17
<< metal1 >>
rect 0 496 2024 592
rect 570 320 628 329
rect 942 320 1000 329
rect 1494 320 1552 329
rect 570 292 1552 320
rect 570 283 628 292
rect 942 283 1000 292
rect 1494 283 1552 292
rect 478 252 536 261
rect 754 252 812 261
rect 1126 252 1184 261
rect 1402 252 1460 261
rect 478 224 1460 252
rect 478 215 536 224
rect 754 215 812 224
rect 1126 215 1184 224
rect 1402 215 1460 224
rect 0 -48 2024 48
<< obsm1 >>
rect 570 184 628 193
rect 1310 184 1368 193
rect 570 156 1368 184
rect 570 147 628 156
rect 1310 147 1368 156
<< labels >>
rlabel metal1 s 1402 215 1460 224 6 A
port 1 nsew signal input
rlabel metal1 s 1126 215 1184 224 6 A
port 1 nsew signal input
rlabel metal1 s 754 215 812 224 6 A
port 1 nsew signal input
rlabel metal1 s 478 215 536 224 6 A
port 1 nsew signal input
rlabel metal1 s 478 224 1460 252 6 A
port 1 nsew signal input
rlabel metal1 s 1402 252 1460 261 6 A
port 1 nsew signal input
rlabel metal1 s 1126 252 1184 261 6 A
port 1 nsew signal input
rlabel metal1 s 754 252 812 261 6 A
port 1 nsew signal input
rlabel metal1 s 478 252 536 261 6 A
port 1 nsew signal input
rlabel metal1 s 1494 283 1552 292 6 B
port 2 nsew signal input
rlabel metal1 s 942 283 1000 292 6 B
port 2 nsew signal input
rlabel metal1 s 570 283 628 292 6 B
port 2 nsew signal input
rlabel metal1 s 570 292 1552 320 6 B
port 2 nsew signal input
rlabel metal1 s 1494 320 1552 329 6 B
port 2 nsew signal input
rlabel metal1 s 942 320 1000 329 6 B
port 2 nsew signal input
rlabel metal1 s 570 320 628 329 6 B
port 2 nsew signal input
rlabel locali s 834 193 1078 250 6 CIN
port 3 nsew signal input
rlabel locali s 1319 271 1369 303 6 CIN
port 3 nsew signal input
rlabel locali s 1044 250 1078 287 6 CIN
port 3 nsew signal input
rlabel locali s 1044 287 1116 303 6 CIN
port 3 nsew signal input
rlabel locali s 1044 303 1369 337 6 CIN
port 3 nsew signal input
rlabel locali s 834 250 868 314 6 CIN
port 3 nsew signal input
rlabel locali s 610 221 684 255 6 CIN
port 3 nsew signal input
rlabel locali s 650 255 684 314 6 CIN
port 3 nsew signal input
rlabel locali s 1319 337 1369 391 6 CIN
port 3 nsew signal input
rlabel locali s 650 314 868 348 6 CIN
port 3 nsew signal input
rlabel metal1 s 0 -48 2024 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2006 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1538 157 2006 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 157 439 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2062 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2024 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 271 63 337 97 6 COUT
port 8 nsew signal output
rlabel locali s 271 97 305 147 6 COUT
port 8 nsew signal output
rlabel locali s 103 51 169 147 6 COUT
port 8 nsew signal output
rlabel locali s 17 147 305 181 6 COUT
port 8 nsew signal output
rlabel locali s 17 181 87 283 6 COUT
port 8 nsew signal output
rlabel locali s 17 283 314 317 6 COUT
port 8 nsew signal output
rlabel locali s 280 317 314 356 6 COUT
port 8 nsew signal output
rlabel locali s 280 356 329 390 6 COUT
port 8 nsew signal output
rlabel locali s 287 390 329 493 6 COUT
port 8 nsew signal output
rlabel locali s 103 317 169 489 6 COUT
port 8 nsew signal output
rlabel locali s 1832 54 1898 147 6 SUM
port 9 nsew signal output
rlabel locali s 1664 51 1730 97 6 SUM
port 9 nsew signal output
rlabel locali s 1680 97 1730 147 6 SUM
port 9 nsew signal output
rlabel locali s 1680 147 2007 181 6 SUM
port 9 nsew signal output
rlabel locali s 1940 181 2007 283 6 SUM
port 9 nsew signal output
rlabel locali s 1680 283 2007 317 6 SUM
port 9 nsew signal output
rlabel locali s 1832 317 1898 485 6 SUM
port 9 nsew signal output
rlabel locali s 1680 317 1714 359 6 SUM
port 9 nsew signal output
rlabel locali s 1664 359 1714 393 6 SUM
port 9 nsew signal output
rlabel locali s 1664 393 1698 493 6 SUM
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2024 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2093974
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2078288
<< end >>
