magic
tech sky130B
timestamp 1704896540
<< properties >>
string GDS_END 7564366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7563978
<< end >>
