magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -79 -26 199 110
<< mvnmos >>
rect 0 0 120 84
<< mvndiff >>
rect -53 46 0 84
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 120 46 173 84
rect 120 12 131 46
rect 165 12 173 46
rect 120 0 173 12
<< mvndiffc >>
rect -45 12 -11 46
rect 131 12 165 46
<< poly >>
rect 0 84 120 110
rect 0 -26 120 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 131 46 165 62
rect 131 -4 165 12
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_1
timestamp 1704896540
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 148 29 148 29 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87932390
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87931500
<< end >>
