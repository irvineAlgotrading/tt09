magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< locali >>
rect -2738 11533 -2704 11603
rect -2276 11533 -2242 11603
rect -1924 11533 -1890 11603
rect -1572 11533 -1538 11603
rect -648 11533 -614 11603
rect -296 11533 -262 11603
rect 56 11533 90 11603
rect 408 11533 442 11603
rect 760 11533 794 11603
rect 1112 11533 1146 11603
rect 1464 11533 1498 11603
rect 1816 11533 1850 11603
rect 2168 11533 2202 11603
rect 2520 11533 2554 11603
rect 11410 8898 11444 8968
rect 11762 8356 11881 8968
rect 11762 7452 11881 8002
rect 11762 6616 11881 7228
<< metal1 >>
rect 12128 14692 12448 14738
rect -1256 14201 -937 14247
rect -371 12528 -51 12576
rect -459 12110 -139 12158
rect 7753 10254 8073 10300
rect 287 9059 535 9065
rect -4289 8981 -4124 8987
rect 287 8815 289 9059
rect 533 8815 535 9059
tri 11668 8956 11674 8962 ne
rect 11674 8956 11680 9008
rect 11732 8956 11744 9008
rect 11796 8956 11802 9008
tri 11802 8956 11808 8962 nw
rect 287 8802 535 8815
rect 287 8750 289 8802
rect 341 8750 353 8802
rect 405 8750 417 8802
rect 469 8750 481 8802
rect 533 8750 535 8802
rect 287 8737 535 8750
rect -1229 8659 -1223 8711
rect -1171 8659 -1159 8711
rect -1107 8659 -1101 8711
rect 287 8685 289 8737
rect 341 8685 353 8737
rect 405 8685 417 8737
rect 469 8685 481 8737
rect 533 8685 535 8737
rect 287 8672 535 8685
rect 287 8620 289 8672
rect 341 8620 353 8672
rect 405 8620 417 8672
rect 469 8620 481 8672
rect 533 8620 535 8672
rect 287 8607 535 8620
rect 287 8555 289 8607
rect 341 8555 353 8607
rect 405 8555 417 8607
rect 469 8555 481 8607
rect 533 8555 535 8607
rect 287 8549 535 8555
tri -3566 8342 -3549 8359 se
rect -3549 8342 -3314 8359
rect -3890 8307 -3314 8342
rect -1229 8307 -1223 8359
rect -1171 8307 -1159 8359
rect -1107 8307 -1101 8359
rect -3890 8290 -3544 8307
tri -3544 8290 -3527 8307 nw
tri -3464 8290 -3447 8307 ne
rect -3447 8290 -3385 8307
tri -3890 8263 -3863 8290 nw
tri -3447 8282 -3439 8290 ne
tri -3515 8017 -3439 8093 se
rect -3439 8071 -3385 8290
tri -3385 8282 -3360 8307 nw
rect -1647 8217 -1641 8269
rect -1589 8217 -1577 8269
rect -1525 8217 -1513 8269
rect -1461 8217 -1449 8269
rect -1397 8217 -1391 8269
rect -684 8208 -211 8362
tri -3439 8017 -3385 8071 nw
tri 11827 8144 11875 8192 se
tri 11180 8017 11202 8039 sw
tri -3517 8015 -3515 8017 se
rect -3515 8015 -3495 8017
rect -3936 7961 -3495 8015
tri -3495 7961 -3439 8017 nw
rect 11180 8014 11202 8017
tri 11202 8014 11205 8017 sw
rect -3936 7888 -3650 7961
tri -3650 7936 -3625 7961 nw
rect -2668 7919 -1798 7930
rect -2668 7867 -2657 7919
rect -2605 7867 -2585 7919
rect -2533 7867 -2514 7919
rect -2462 7867 -2443 7919
rect -2391 7867 -2372 7919
rect -2320 7867 -2301 7919
rect -2249 7867 -2230 7919
rect -2178 7867 -1798 7919
rect 11143 7884 11315 8014
rect -2668 7859 -1798 7867
tri -1872 7831 -1844 7859 ne
rect -1844 7856 -1798 7859
rect -4099 7713 -4073 7755
rect 11180 7440 11244 7884
tri 11180 7415 11205 7440 nw
rect 11827 7406 11875 8144
tri 11827 7396 11837 7406 ne
rect 11837 7396 11875 7406
tri -1527 7386 -1517 7396 se
tri 11837 7386 11847 7396 ne
rect 11847 7386 11875 7396
rect -1636 7334 -1516 7386
tri 11847 7358 11875 7386 ne
tri -1542 7309 -1517 7334 ne
tri -1542 7034 -1517 7059 se
rect -4700 6992 -4666 7029
rect -1636 6982 -1516 7034
tri -1542 6957 -1517 6982 ne
rect 4837 6874 5157 6922
tri -3310 6805 -3285 6830 se
rect -3893 6804 -3285 6805
rect -3893 6793 -3236 6804
rect -3893 6741 -3495 6793
rect -3443 6741 -3428 6793
rect -3376 6741 -3362 6793
rect -3310 6741 -3236 6793
rect 11802 6765 11875 7200
rect -3893 6729 -3236 6741
tri 11842 6732 11875 6765 ne
rect -3893 6677 -3495 6729
rect -3443 6677 -3428 6729
rect -3376 6677 -3362 6729
rect -3310 6677 -3236 6729
rect -3893 6666 -3236 6677
tri -3310 6641 -3285 6666 ne
tri -1542 6492 -1517 6517 se
rect -1636 6440 -1516 6492
tri -1542 6415 -1517 6440 ne
rect -955 6360 -949 6412
rect -897 6360 -868 6412
rect -816 6360 -788 6412
rect -736 6360 -708 6412
rect -656 6360 -650 6412
rect -607 6360 -601 6412
rect -549 6360 -520 6412
rect -468 6360 -440 6412
rect -388 6360 -360 6412
rect -308 6360 -302 6412
rect 13513 6346 13565 6397
rect -5733 5610 -5605 5611
rect -5733 5558 -5727 5610
rect -5675 5558 -5663 5610
rect -5611 5558 -5605 5610
rect -5733 5536 -5605 5558
rect -5733 5484 -5727 5536
rect -5675 5484 -5663 5536
rect -5611 5484 -5605 5536
rect -5733 5462 -5605 5484
rect -5733 5410 -5727 5462
rect -5675 5410 -5663 5462
rect -5611 5410 -5605 5462
rect -5733 5409 -5605 5410
rect -5733 5170 -5605 5171
rect -5733 5118 -5727 5170
rect -5675 5118 -5663 5170
rect -5611 5118 -5605 5170
rect -5733 5096 -5605 5118
rect -5733 5044 -5727 5096
rect -5675 5044 -5663 5096
rect -5611 5044 -5605 5096
rect -4526 5074 -4324 5093
rect -5733 5022 -5605 5044
rect -5733 4970 -5727 5022
rect -5675 4970 -5663 5022
rect -5611 4970 -5605 5022
rect -5733 4969 -5605 4970
rect -5025 4884 -4971 5070
tri -4971 4884 -4785 5070 sw
rect -4526 5022 -4520 5074
rect -4468 5022 -4451 5074
rect -4399 5022 -4382 5074
rect -4330 5022 -4324 5074
rect -4526 5010 -4324 5022
rect -4526 4958 -4520 5010
rect -4468 4958 -4451 5010
rect -4399 4958 -4382 5010
rect -4330 4958 -4324 5010
rect -4526 4939 -4324 4958
rect -5025 4876 -4703 4884
rect -5025 4870 -4768 4876
tri -4961 4745 -4836 4870 ne
rect -4836 4824 -4768 4870
rect -4716 4824 -4703 4876
rect -4836 4805 -4703 4824
rect -4836 4753 -4768 4805
rect -4716 4753 -4703 4805
rect -4836 4745 -4703 4753
tri -5168 4547 -5107 4608 se
rect -5107 4606 -5074 4608
rect -5064 4606 -5061 4711
tri -5061 4606 -4956 4711 sw
rect -5107 4600 -4705 4606
rect -5107 4548 -4768 4600
rect -4716 4548 -4705 4600
rect -5107 4547 -4705 4548
rect -5212 4531 -4705 4547
rect -5212 4522 -4768 4531
tri -5212 4335 -5025 4522 ne
rect -5025 4479 -4768 4522
rect -4716 4479 -4705 4531
rect -5025 4462 -4705 4479
rect -5025 4410 -4768 4462
rect -4716 4410 -4705 4462
rect -5025 4392 -4705 4410
rect -5025 4340 -4768 4392
rect -4716 4340 -4705 4392
rect -5025 4322 -4705 4340
rect -5025 4270 -4768 4322
rect -4716 4270 -4705 4322
rect -5025 4252 -4705 4270
rect -3433 4578 -3183 4584
rect -3433 4526 -3430 4578
rect -3378 4526 -3366 4578
rect -3314 4526 -3302 4578
rect -3250 4526 -3238 4578
rect -3186 4526 -3183 4578
rect -3433 4513 -3183 4526
rect -3433 4461 -3430 4513
rect -3378 4461 -3366 4513
rect -3314 4461 -3302 4513
rect -3250 4461 -3238 4513
rect -3186 4461 -3183 4513
rect -3433 4448 -3183 4461
rect -3433 4396 -3430 4448
rect -3378 4396 -3366 4448
rect -3314 4396 -3302 4448
rect -3250 4396 -3238 4448
rect -3186 4396 -3183 4448
rect -3433 4382 -3183 4396
rect -3433 4330 -3430 4382
rect -3378 4330 -3366 4382
rect -3314 4330 -3302 4382
rect -3250 4330 -3238 4382
rect -3186 4330 -3183 4382
rect -3433 4316 -3183 4330
rect -3433 4264 -3430 4316
rect -3378 4264 -3366 4316
rect -3314 4264 -3302 4316
rect -3250 4264 -3238 4316
rect -3186 4264 -3183 4316
rect -3433 4258 -3183 4264
rect -2648 4466 -2596 4472
rect -2648 4400 -2596 4414
rect -2648 4334 -2596 4348
rect -2648 4268 -2596 4282
rect -5025 4200 -4768 4252
rect -4716 4200 -4705 4252
rect -5025 4182 -4705 4200
rect -5025 4130 -4768 4182
rect -4716 4130 -4705 4182
rect -5025 4124 -4705 4130
rect -2648 4202 -2596 4216
rect -2648 4136 -2596 4150
rect -2648 4070 -2596 4084
rect -2648 4004 -2596 4018
rect -2648 3938 -2596 3952
rect -5025 3870 -4703 3878
rect -5025 3818 -4768 3870
rect -4716 3818 -4703 3870
rect -5025 3799 -4703 3818
rect -5025 3747 -4768 3799
rect -4716 3747 -4703 3799
rect -5025 3743 -4703 3747
tri -4888 3739 -4884 3743 ne
rect -4884 3739 -4703 3743
rect -2648 3872 -2596 3886
rect -2648 3806 -2596 3820
rect -2648 3740 -2596 3754
rect -410 3772 -276 3778
rect -358 3720 -346 3772
rect -294 3732 -276 3772
rect -410 3714 -294 3720
tri -294 3714 -276 3732 nw
rect 8654 3707 8809 3759
rect -2648 3675 -2596 3688
rect -2648 3617 -2596 3623
rect -4783 3086 -4755 3120
rect -4867 3024 -4813 3058
rect -4779 2816 -4705 2822
rect -4779 2764 -4768 2816
rect -4716 2764 -4705 2816
rect -4779 2745 -4705 2764
rect -4779 2693 -4768 2745
rect -4716 2693 -4705 2745
tri -1978 2784 -1952 2810 sw
tri -1864 2784 -1838 2810 se
rect -1978 2738 -1838 2784
tri -1838 2738 -1812 2764 nw
rect -4779 2687 -4705 2693
rect -4982 2587 -4944 2633
tri -5058 2130 -5025 2163 se
rect -5025 2155 -4709 2163
rect -5025 2130 -4772 2155
rect -5222 2103 -4772 2130
rect -4720 2103 -4709 2155
rect -5222 2084 -4709 2103
rect -5222 2078 -4772 2084
tri -5079 2024 -5025 2078 ne
rect -5025 2032 -4772 2078
rect -4720 2032 -4709 2084
rect -5025 2024 -4709 2032
rect -4704 1956 -4667 1996
rect -2195 1569 -2189 1685
rect -2009 1569 -2003 1685
<< via1 >>
rect 289 8815 533 9059
rect 11680 8956 11732 9008
rect 11744 8956 11796 9008
rect 289 8750 341 8802
rect 353 8750 405 8802
rect 417 8750 469 8802
rect 481 8750 533 8802
rect -1223 8659 -1171 8711
rect -1159 8659 -1107 8711
rect 289 8685 341 8737
rect 353 8685 405 8737
rect 417 8685 469 8737
rect 481 8685 533 8737
rect 289 8620 341 8672
rect 353 8620 405 8672
rect 417 8620 469 8672
rect 481 8620 533 8672
rect 289 8555 341 8607
rect 353 8555 405 8607
rect 417 8555 469 8607
rect 481 8555 533 8607
rect -1223 8307 -1171 8359
rect -1159 8307 -1107 8359
rect -1641 8217 -1589 8269
rect -1577 8217 -1525 8269
rect -1513 8217 -1461 8269
rect -1449 8217 -1397 8269
rect -2657 7867 -2605 7919
rect -2585 7867 -2533 7919
rect -2514 7867 -2462 7919
rect -2443 7867 -2391 7919
rect -2372 7867 -2320 7919
rect -2301 7867 -2249 7919
rect -2230 7867 -2178 7919
rect -3495 6741 -3443 6793
rect -3428 6741 -3376 6793
rect -3362 6741 -3310 6793
rect -3495 6677 -3443 6729
rect -3428 6677 -3376 6729
rect -3362 6677 -3310 6729
rect -949 6360 -897 6412
rect -868 6360 -816 6412
rect -788 6360 -736 6412
rect -708 6360 -656 6412
rect -601 6360 -549 6412
rect -520 6360 -468 6412
rect -440 6360 -388 6412
rect -360 6360 -308 6412
rect -5727 5558 -5675 5610
rect -5663 5558 -5611 5610
rect -5727 5484 -5675 5536
rect -5663 5484 -5611 5536
rect -5727 5410 -5675 5462
rect -5663 5410 -5611 5462
rect -5727 5118 -5675 5170
rect -5663 5118 -5611 5170
rect -5727 5044 -5675 5096
rect -5663 5044 -5611 5096
rect -5727 4970 -5675 5022
rect -5663 4970 -5611 5022
rect -4520 5022 -4468 5074
rect -4451 5022 -4399 5074
rect -4382 5022 -4330 5074
rect -4520 4958 -4468 5010
rect -4451 4958 -4399 5010
rect -4382 4958 -4330 5010
rect -4768 4824 -4716 4876
rect -4768 4753 -4716 4805
rect -4768 4548 -4716 4600
rect -4768 4479 -4716 4531
rect -4768 4410 -4716 4462
rect -4768 4340 -4716 4392
rect -4768 4270 -4716 4322
rect -3430 4526 -3378 4578
rect -3366 4526 -3314 4578
rect -3302 4526 -3250 4578
rect -3238 4526 -3186 4578
rect -3430 4461 -3378 4513
rect -3366 4461 -3314 4513
rect -3302 4461 -3250 4513
rect -3238 4461 -3186 4513
rect -3430 4396 -3378 4448
rect -3366 4396 -3314 4448
rect -3302 4396 -3250 4448
rect -3238 4396 -3186 4448
rect -3430 4330 -3378 4382
rect -3366 4330 -3314 4382
rect -3302 4330 -3250 4382
rect -3238 4330 -3186 4382
rect -3430 4264 -3378 4316
rect -3366 4264 -3314 4316
rect -3302 4264 -3250 4316
rect -3238 4264 -3186 4316
rect -2648 4414 -2596 4466
rect -2648 4348 -2596 4400
rect -2648 4282 -2596 4334
rect -4768 4200 -4716 4252
rect -4768 4130 -4716 4182
rect -2648 4216 -2596 4268
rect -2648 4150 -2596 4202
rect -2648 4084 -2596 4136
rect -2648 4018 -2596 4070
rect -2648 3952 -2596 4004
rect -2648 3886 -2596 3938
rect -4768 3818 -4716 3870
rect -4768 3747 -4716 3799
rect -2648 3820 -2596 3872
rect -2648 3754 -2596 3806
rect -2648 3688 -2596 3740
rect -410 3720 -358 3772
rect -346 3720 -294 3772
rect -2648 3623 -2596 3675
rect -4768 2764 -4716 2816
rect -4768 2693 -4716 2745
rect -4772 2103 -4720 2155
rect -4772 2032 -4720 2084
rect -2189 1569 -2009 1685
<< metal2 >>
rect -2311 10380 -1991 11376
rect -302 10380 546 11752
rect 9068 11640 9542 11734
rect 11057 11640 11377 11734
rect 13155 11691 13506 11734
rect -4041 9915 -3721 9961
rect -3565 9915 -3245 9961
rect 287 9059 535 9065
rect 287 8815 289 9059
rect 533 8815 535 9059
rect 11674 8956 11680 9008
rect 11732 8956 11744 9008
rect 11796 8956 11802 9008
rect 287 8802 535 8815
rect 287 8750 289 8802
rect 341 8750 353 8802
rect 405 8750 417 8802
rect 469 8750 481 8802
rect 533 8750 535 8802
rect 287 8737 535 8750
rect -1229 8659 -1223 8711
rect -1171 8659 -1159 8711
rect -1107 8659 -1101 8711
rect 287 8685 289 8737
rect 341 8685 353 8737
rect 405 8685 417 8737
rect 469 8685 481 8737
rect 533 8685 535 8737
rect 287 8672 535 8685
tri 10356 8819 10381 8844 sw
rect 10356 8714 10578 8819
tri 10578 8714 10683 8819 sw
rect 10356 8677 10683 8714
rect 287 8620 289 8672
rect 341 8620 353 8672
rect 405 8620 417 8672
rect 469 8620 481 8672
rect 533 8620 535 8672
rect 287 8607 535 8620
tri 10491 8613 10555 8677 ne
rect 287 8555 289 8607
rect 341 8555 353 8607
rect 405 8555 417 8607
rect 469 8555 481 8607
rect 533 8555 535 8607
rect 287 8549 535 8555
rect -1229 8307 -1223 8359
rect -1171 8307 -1159 8359
rect -1107 8307 -1101 8359
rect -1647 8217 -1641 8269
rect -1589 8217 -1577 8269
rect -1525 8217 -1513 8269
rect -1461 8217 -1449 8269
rect -1397 8217 -1391 8269
rect -2663 7919 -2172 7926
rect -2663 7867 -2657 7919
rect -2605 7867 -2585 7919
rect -2533 7867 -2514 7919
rect -2462 7867 -2443 7919
rect -2391 7867 -2372 7919
rect -2320 7867 -2301 7919
rect -2249 7867 -2230 7919
rect -2178 7867 -2172 7919
rect -2663 7860 -2172 7867
rect -4526 7812 -4324 7821
rect -4526 7756 -4493 7812
rect -4437 7756 -4413 7812
rect -4357 7756 -4324 7812
rect -4526 7728 -4324 7756
rect -4526 7672 -4493 7728
rect -4437 7672 -4413 7728
rect -4357 7672 -4324 7728
rect -4526 7644 -4324 7672
rect -4526 7588 -4493 7644
rect -4437 7588 -4413 7644
rect -4357 7588 -4324 7644
rect -4526 7559 -4324 7588
rect -4526 7503 -4493 7559
rect -4437 7503 -4413 7559
rect -4357 7503 -4324 7559
rect -2667 7507 -2167 7555
rect -1864 7507 -1545 7555
rect -4526 7474 -4324 7503
rect -4526 7418 -4493 7474
rect -4437 7418 -4413 7474
rect -4357 7418 -4324 7474
rect -4526 7389 -4324 7418
rect 10555 7412 10683 8677
rect 11673 8173 11805 8182
rect 11673 8117 11711 8173
rect 11767 8117 11805 8173
rect 11673 8080 11805 8117
rect 11673 8024 11711 8080
rect 11767 8024 11805 8080
rect 11673 7987 11805 8024
rect 11673 7931 11711 7987
rect 11767 7931 11805 7987
rect 11673 7894 11805 7931
rect 11673 7838 11711 7894
rect 11767 7838 11805 7894
rect 11673 7800 11805 7838
rect 11673 7744 11711 7800
rect 11767 7744 11805 7800
rect 11673 7706 11805 7744
rect 11673 7650 11711 7706
rect 11767 7650 11805 7706
rect 11673 7641 11805 7650
rect 11631 7602 11687 7611
rect 11631 7497 11687 7546
rect -4526 7333 -4493 7389
rect -4437 7333 -4413 7389
rect -4357 7333 -4324 7389
rect -4526 7324 -4324 7333
rect 11631 7392 11687 7441
rect 11631 7327 11687 7336
rect -3501 6793 -3304 6801
rect -3501 6741 -3495 6793
rect -3443 6741 -3428 6793
rect -3376 6741 -3362 6793
rect -3310 6741 -3304 6793
rect -3501 6729 -3304 6741
rect -3501 6677 -3495 6729
rect -3443 6677 -3428 6729
rect -3376 6677 -3362 6729
rect -3310 6677 -3304 6729
rect -962 6697 -642 6745
rect -614 6697 -294 6745
rect 762 6683 1082 6745
rect -3501 6669 -3304 6677
rect 1430 6651 1729 6746
rect 2349 6651 3040 6745
rect 3148 6651 3720 6745
rect 3975 6651 4343 6745
rect 4399 6651 5082 6745
rect 5193 6651 6150 6745
rect 6378 6651 7035 6745
rect 7498 6651 7891 6745
rect 8132 6651 8330 6745
rect 8489 6651 8809 6745
rect -955 6360 -949 6412
rect -897 6360 -868 6412
rect -816 6360 -788 6412
rect -736 6360 -708 6412
rect -656 6360 -650 6412
rect -607 6360 -601 6412
rect -549 6360 -520 6412
rect -468 6360 -440 6412
rect -388 6360 -360 6412
rect -308 6360 -302 6412
rect 78 6399 134 6408
tri 53 6335 78 6360 ne
rect 78 6316 134 6343
rect 78 6233 134 6260
rect 78 6150 134 6177
rect 78 6067 134 6094
rect 78 5984 134 6011
rect 78 5919 134 5928
tri 78 5915 82 5919 ne
rect 82 5915 134 5919
rect 1761 5879 1813 6117
rect -5733 5610 -5605 5611
rect -5733 5558 -5727 5610
rect -5675 5558 -5663 5610
rect -5611 5558 -5605 5610
rect -5733 5536 -5605 5558
rect -5733 5484 -5727 5536
rect -5675 5484 -5663 5536
rect -5611 5484 -5605 5536
rect -5733 5462 -5605 5484
rect -5733 5410 -5727 5462
rect -5675 5410 -5663 5462
rect -5611 5410 -5605 5462
rect -5733 5409 -5605 5410
rect -4526 5370 -4324 5379
rect -4526 5314 -4493 5370
rect -4437 5314 -4413 5370
rect -4357 5314 -4324 5370
rect -4526 5285 -4324 5314
rect -4526 5229 -4493 5285
rect -4437 5229 -4413 5285
rect -4357 5229 -4324 5285
rect -4526 5200 -4324 5229
rect -5733 5170 -5605 5171
rect -5733 5118 -5727 5170
rect -5675 5118 -5663 5170
rect -5611 5118 -5605 5170
rect -5733 5096 -5605 5118
rect -5733 5044 -5727 5096
rect -5675 5044 -5663 5096
rect -5611 5044 -5605 5096
rect -5733 5022 -5605 5044
rect -5733 4970 -5727 5022
rect -5675 4970 -5663 5022
rect -5611 4970 -5605 5022
rect -5733 4969 -5605 4970
rect -4526 5144 -4493 5200
rect -4437 5144 -4413 5200
rect -4357 5144 -4324 5200
rect -4526 5114 -4324 5144
rect -4526 5074 -4493 5114
rect -4437 5074 -4413 5114
rect -4357 5074 -4324 5114
rect -4526 5022 -4520 5074
rect -4468 5028 -4451 5058
rect -4399 5028 -4382 5058
rect -4330 5022 -4324 5074
rect -4526 5010 -4493 5022
rect -4437 5010 -4413 5022
rect -4357 5010 -4324 5022
rect -4526 4958 -4520 5010
rect -4468 4958 -4451 4972
rect -4399 4958 -4382 4972
rect -4330 4958 -4324 5010
rect -4526 4942 -4324 4958
rect -4526 4886 -4493 4942
rect -4437 4886 -4413 4942
rect -4357 4886 -4324 4942
rect -4779 4876 -4705 4882
rect -4779 4824 -4768 4876
rect -4716 4824 -4705 4876
rect -4779 4805 -4705 4824
rect -4779 4753 -4768 4805
rect -4716 4753 -4705 4805
rect -4779 4747 -4705 4753
rect -4526 4856 -4324 4886
rect -4526 4800 -4493 4856
rect -4437 4800 -4413 4856
rect -4357 4800 -4324 4856
rect -4526 4770 -4324 4800
rect -4526 4714 -4493 4770
rect -4437 4714 -4413 4770
rect -4357 4714 -4324 4770
rect -4526 4684 -4324 4714
rect -4526 4628 -4493 4684
rect -4437 4628 -4413 4684
rect -4357 4628 -4324 4684
rect -4779 4600 -4705 4606
rect -4779 4548 -4768 4600
rect -4716 4548 -4705 4600
rect -4779 4531 -4705 4548
rect -4526 4598 -4324 4628
rect -4526 4542 -4493 4598
rect -4437 4542 -4413 4598
rect -4357 4542 -4324 4598
rect 1841 5378 1903 5387
rect 1841 5322 1844 5378
rect 1900 5322 1903 5378
rect 1841 5291 1903 5322
rect 1841 5235 1844 5291
rect 1900 5235 1903 5291
rect 1841 5204 1903 5235
rect 1841 5148 1844 5204
rect 1900 5148 1903 5204
rect 1841 5117 1903 5148
rect 1841 5061 1844 5117
rect 1900 5061 1903 5117
rect 1841 5030 1903 5061
rect 3980 5361 4338 5381
rect 3980 5305 3989 5361
rect 4045 5305 4084 5361
rect 4140 5305 4179 5361
rect 4235 5305 4273 5361
rect 4329 5305 4338 5361
rect 3980 5281 4338 5305
rect 3980 5225 3989 5281
rect 4045 5225 4084 5281
rect 4140 5225 4179 5281
rect 4235 5225 4273 5281
rect 4329 5225 4338 5281
rect 3980 5201 4338 5225
rect 3980 5145 3989 5201
rect 4045 5145 4084 5201
rect 4140 5145 4179 5201
rect 4235 5145 4273 5201
rect 4329 5145 4338 5201
rect 3980 5121 4338 5145
rect 3980 5065 3989 5121
rect 4045 5065 4084 5121
rect 4140 5065 4179 5121
rect 4235 5065 4273 5121
rect 4329 5065 4338 5121
rect 3980 5045 4338 5065
rect 6473 5378 6553 5387
rect 6473 5322 6485 5378
rect 6541 5322 6553 5378
rect 8240 5371 8364 5380
rect 6473 5291 6553 5322
rect 6473 5235 6485 5291
rect 6541 5235 6553 5291
rect 6473 5204 6553 5235
rect 6473 5148 6485 5204
rect 6541 5148 6553 5204
rect 6473 5117 6553 5148
rect 6473 5061 6485 5117
rect 6541 5061 6553 5117
rect 1841 4974 1844 5030
rect 1900 4974 1903 5030
rect 1841 4943 1903 4974
rect 1841 4887 1844 4943
rect 1900 4887 1903 4943
rect 1841 4856 1903 4887
rect 1841 4800 1844 4856
rect 1900 4800 1903 4856
rect 1841 4769 1903 4800
rect 1841 4713 1844 4769
rect 1900 4713 1903 4769
rect 1841 4682 1903 4713
rect 1841 4626 1844 4682
rect 1900 4626 1903 4682
rect 1841 4594 1903 4626
rect -4526 4533 -4324 4542
rect -3433 4578 -3183 4584
rect -4779 4479 -4768 4531
rect -4716 4479 -4705 4531
rect -4779 4462 -4705 4479
rect -4779 4410 -4768 4462
rect -4716 4410 -4705 4462
rect -4779 4392 -4705 4410
rect -4779 4340 -4768 4392
rect -4716 4340 -4705 4392
rect -4779 4322 -4705 4340
rect -4779 4270 -4768 4322
rect -4716 4270 -4705 4322
rect -4779 4252 -4705 4270
rect -3433 4526 -3430 4578
rect -3378 4526 -3366 4578
rect -3314 4526 -3302 4578
rect -3250 4526 -3238 4578
rect -3186 4526 -3183 4578
rect 1841 4538 1844 4594
rect 1900 4538 1903 4594
rect 1841 4529 1903 4538
rect 6473 5030 6553 5061
rect 6473 4974 6485 5030
rect 6541 4974 6553 5030
rect 6473 4943 6553 4974
rect 6473 4887 6485 4943
rect 6541 4887 6553 4943
rect 6473 4856 6553 4887
rect 6473 4800 6485 4856
rect 6541 4800 6553 4856
rect 6473 4769 6553 4800
rect 6473 4713 6485 4769
rect 6541 4713 6553 4769
rect 6473 4682 6553 4713
rect 6473 4626 6485 4682
rect 6541 4626 6553 4682
rect 6473 4594 6553 4626
rect 6473 4538 6485 4594
rect 6541 4538 6553 4594
rect 6473 4529 6553 4538
rect 7594 5338 8075 5346
rect 7594 5282 7603 5338
rect 7659 5282 7685 5338
rect 7741 5282 7767 5338
rect 7823 5282 7848 5338
rect 7904 5282 7929 5338
rect 7985 5282 8010 5338
rect 8066 5282 8075 5338
rect 7594 5256 8075 5282
rect 7594 5200 7603 5256
rect 7659 5200 7685 5256
rect 7741 5200 7767 5256
rect 7823 5200 7848 5256
rect 7904 5200 7929 5256
rect 7985 5200 8010 5256
rect 8066 5200 8075 5256
rect 7594 5174 8075 5200
rect 7594 5118 7603 5174
rect 7659 5118 7685 5174
rect 7741 5118 7767 5174
rect 7823 5118 7848 5174
rect 7904 5118 7929 5174
rect 7985 5118 8010 5174
rect 8066 5118 8075 5174
rect 7594 5092 8075 5118
rect 7594 5036 7603 5092
rect 7659 5036 7685 5092
rect 7741 5036 7767 5092
rect 7823 5036 7848 5092
rect 7904 5036 7929 5092
rect 7985 5036 8010 5092
rect 8066 5036 8075 5092
rect 7594 5010 8075 5036
rect 7594 4954 7603 5010
rect 7659 4954 7685 5010
rect 7741 4954 7767 5010
rect 7823 4954 7848 5010
rect 7904 4954 7929 5010
rect 7985 4954 8010 5010
rect 8066 4954 8075 5010
rect 7594 4928 8075 4954
rect 7594 4872 7603 4928
rect 7659 4872 7685 4928
rect 7741 4872 7767 4928
rect 7823 4872 7848 4928
rect 7904 4872 7929 4928
rect 7985 4872 8010 4928
rect 8066 4872 8075 4928
rect 7594 4846 8075 4872
rect 7594 4790 7603 4846
rect 7659 4790 7685 4846
rect 7741 4790 7767 4846
rect 7823 4790 7848 4846
rect 7904 4790 7929 4846
rect 7985 4790 8010 4846
rect 8066 4790 8075 4846
rect 7594 4764 8075 4790
rect 7594 4708 7603 4764
rect 7659 4708 7685 4764
rect 7741 4708 7767 4764
rect 7823 4708 7848 4764
rect 7904 4708 7929 4764
rect 7985 4708 8010 4764
rect 8066 4708 8075 4764
rect 7594 4682 8075 4708
rect 7594 4626 7603 4682
rect 7659 4626 7685 4682
rect 7741 4626 7767 4682
rect 7823 4626 7848 4682
rect 7904 4626 7929 4682
rect 7985 4626 8010 4682
rect 8066 4626 8075 4682
rect 8240 5315 8274 5371
rect 8330 5315 8364 5371
rect 8240 5291 8364 5315
rect 8240 5235 8274 5291
rect 8330 5235 8364 5291
rect 8240 5211 8364 5235
rect 8240 5155 8274 5211
rect 8330 5155 8364 5211
rect 8240 5131 8364 5155
rect 8240 5075 8274 5131
rect 8330 5075 8364 5131
rect 8240 5051 8364 5075
rect 8240 4995 8274 5051
rect 8330 4995 8364 5051
rect 8240 4971 8364 4995
rect 8240 4915 8274 4971
rect 8330 4915 8364 4971
rect 8240 4891 8364 4915
rect 8240 4835 8274 4891
rect 8330 4835 8364 4891
rect 8240 4810 8364 4835
rect 8240 4754 8274 4810
rect 8330 4754 8364 4810
rect 8240 4729 8364 4754
rect 8240 4673 8274 4729
rect 8330 4673 8364 4729
rect 8240 4664 8364 4673
rect 8652 5371 8776 5380
rect 8652 5315 8686 5371
rect 8742 5315 8776 5371
rect 8652 5291 8776 5315
rect 8652 5235 8686 5291
rect 8742 5235 8776 5291
rect 8652 5211 8776 5235
rect 8652 5155 8686 5211
rect 8742 5155 8776 5211
rect 8652 5131 8776 5155
rect 8652 5075 8686 5131
rect 8742 5075 8776 5131
rect 8652 5051 8776 5075
rect 8652 4995 8686 5051
rect 8742 4995 8776 5051
rect 8652 4971 8776 4995
rect 8652 4915 8686 4971
rect 8742 4915 8776 4971
rect 8652 4891 8776 4915
rect 8652 4835 8686 4891
rect 8742 4835 8776 4891
rect 8652 4810 8776 4835
rect 8652 4754 8686 4810
rect 8742 4754 8776 4810
rect 8652 4729 8776 4754
rect 8652 4673 8686 4729
rect 8742 4673 8776 4729
rect 8652 4664 8776 4673
rect 7594 4600 8075 4626
rect 7594 4544 7603 4600
rect 7659 4544 7685 4600
rect 7741 4544 7767 4600
rect 7823 4544 7848 4600
rect 7904 4544 7929 4600
rect 7985 4544 8010 4600
rect 8066 4544 8075 4600
rect 7594 4536 8075 4544
rect -3433 4513 -3183 4526
rect -3433 4461 -3430 4513
rect -3378 4461 -3366 4513
rect -3314 4461 -3302 4513
rect -3250 4461 -3238 4513
rect -3186 4461 -3183 4513
rect -3433 4448 -3183 4461
rect -3433 4396 -3430 4448
rect -3378 4396 -3366 4448
rect -3314 4396 -3302 4448
rect -3250 4396 -3238 4448
rect -3186 4396 -3183 4448
rect -3433 4382 -3183 4396
rect -3433 4330 -3430 4382
rect -3378 4330 -3366 4382
rect -3314 4330 -3302 4382
rect -3250 4330 -3238 4382
rect -3186 4330 -3183 4382
rect -3433 4316 -3183 4330
rect -3433 4264 -3430 4316
rect -3378 4264 -3366 4316
rect -3314 4264 -3302 4316
rect -3250 4264 -3238 4316
rect -3186 4264 -3183 4316
rect -3433 4258 -3183 4264
rect -2648 4466 -2596 4472
rect -2648 4400 -2596 4414
rect -2648 4334 -2596 4348
rect -2648 4268 -2596 4282
rect -4779 4200 -4768 4252
rect -4716 4200 -4705 4252
rect -4779 4182 -4705 4200
rect -4779 4130 -4768 4182
rect -4716 4130 -4705 4182
rect -4779 4124 -4705 4130
rect -2648 4202 -2596 4216
rect -2648 4136 -2596 4150
rect -2648 4070 -2596 4084
rect -2664 4018 -2648 4025
rect -2596 4018 -2354 4025
rect -2664 4016 -2354 4018
rect -2664 3960 -2657 4016
rect -2601 4004 -2577 4016
rect -2596 3960 -2577 4004
rect -2521 3960 -2497 4016
rect -2441 3960 -2417 4016
rect -2361 3960 -2354 4016
rect -2664 3952 -2648 3960
rect -2596 3952 -2354 3960
rect -2664 3938 -2354 3952
rect -2664 3930 -2648 3938
rect -2596 3930 -2354 3938
rect -4779 3870 -4705 3876
rect -4779 3818 -4768 3870
rect -4716 3818 -4705 3870
rect -4779 3799 -4705 3818
rect -4779 3747 -4768 3799
rect -4716 3747 -4705 3799
rect -4779 3741 -4705 3747
rect -2664 3874 -2657 3930
rect -2596 3886 -2577 3930
rect -2601 3874 -2577 3886
rect -2521 3874 -2497 3930
rect -2441 3874 -2417 3930
rect -2361 3874 -2354 3930
rect -2664 3872 -2354 3874
rect -2664 3844 -2648 3872
rect -2596 3844 -2354 3872
rect -2664 3788 -2657 3844
rect -2596 3820 -2577 3844
rect -2601 3806 -2577 3820
rect -2596 3788 -2577 3806
rect -2521 3788 -2497 3844
rect -2441 3788 -2417 3844
rect -2361 3788 -2354 3844
rect -2664 3758 -2648 3788
rect -2596 3758 -2354 3788
rect -2664 3702 -2657 3758
rect -2596 3754 -2577 3758
rect -2601 3740 -2577 3754
rect -2596 3702 -2577 3740
rect -2521 3702 -2497 3758
rect -2441 3702 -2417 3758
rect -2361 3702 -2354 3758
rect -410 3772 -294 3778
rect -358 3720 -346 3772
rect -410 3714 -294 3720
rect -2664 3688 -2648 3702
rect -2596 3688 -2354 3702
rect -2664 3675 -2354 3688
rect -2664 3672 -2648 3675
rect -2596 3672 -2354 3675
rect -2664 3616 -2657 3672
rect -2596 3623 -2577 3672
rect -2601 3616 -2577 3623
rect -2521 3616 -2497 3672
rect -2441 3616 -2417 3672
rect -2361 3616 -2354 3672
rect -2664 3586 -2354 3616
rect -2664 3530 -2657 3586
rect -2601 3530 -2577 3586
rect -2521 3530 -2497 3586
rect -2441 3530 -2417 3586
rect -2361 3530 -2354 3586
rect -2664 3500 -2354 3530
rect -2664 3444 -2657 3500
rect -2601 3444 -2577 3500
rect -2521 3444 -2497 3500
rect -2441 3444 -2417 3500
rect -2361 3444 -2354 3500
rect -2664 3414 -2354 3444
rect -2664 3358 -2657 3414
rect -2601 3358 -2577 3414
rect -2521 3358 -2497 3414
rect -2441 3358 -2417 3414
rect -2361 3358 -2354 3414
rect -2664 3327 -2354 3358
rect -2664 3271 -2657 3327
rect -2601 3271 -2577 3327
rect -2521 3271 -2497 3327
rect -2441 3271 -2417 3327
rect -2361 3271 -2354 3327
rect -2664 3240 -2354 3271
rect -2664 3184 -2657 3240
rect -2601 3184 -2577 3240
rect -2521 3184 -2497 3240
rect -2441 3184 -2417 3240
rect -2361 3184 -2354 3240
rect -2664 3175 -2354 3184
rect -4779 2816 -4705 2822
rect -4779 2764 -4768 2816
rect -4716 2764 -4705 2816
rect -4779 2745 -4705 2764
rect -4779 2693 -4768 2745
rect -4716 2693 -4705 2745
rect -4779 2687 -4705 2693
rect -3979 2629 -3927 2633
tri -3927 2629 -3923 2633 sw
rect -4783 2155 -4709 2161
rect -4783 2103 -4772 2155
rect -4720 2103 -4709 2155
rect -4783 2084 -4709 2103
rect -4783 2032 -4772 2084
rect -4720 2032 -4709 2084
rect -4783 2026 -4709 2032
rect -3979 1835 -3923 2629
rect -3979 1831 -3927 1835
tri -3927 1831 -3923 1835 nw
rect -3075 942 -3023 2928
rect -2195 1569 -2189 1685
rect -2009 1569 -2003 1685
<< via2 >>
rect -4493 7756 -4437 7812
rect -4413 7756 -4357 7812
rect -4493 7672 -4437 7728
rect -4413 7672 -4357 7728
rect -4493 7588 -4437 7644
rect -4413 7588 -4357 7644
rect -4493 7503 -4437 7559
rect -4413 7503 -4357 7559
rect -4493 7418 -4437 7474
rect -4413 7418 -4357 7474
rect 11711 8117 11767 8173
rect 11711 8024 11767 8080
rect 11711 7931 11767 7987
rect 11711 7838 11767 7894
rect 11711 7744 11767 7800
rect 11711 7650 11767 7706
rect 11631 7546 11687 7602
rect 11631 7441 11687 7497
rect -4493 7333 -4437 7389
rect -4413 7333 -4357 7389
rect 11631 7336 11687 7392
rect 78 6343 134 6399
rect 78 6260 134 6316
rect 78 6177 134 6233
rect 78 6094 134 6150
rect 78 6011 134 6067
rect 78 5928 134 5984
rect -4493 5314 -4437 5370
rect -4413 5314 -4357 5370
rect -4493 5229 -4437 5285
rect -4413 5229 -4357 5285
rect -4493 5144 -4437 5200
rect -4413 5144 -4357 5200
rect -4493 5074 -4437 5114
rect -4413 5074 -4357 5114
rect -4493 5058 -4468 5074
rect -4468 5058 -4451 5074
rect -4451 5058 -4437 5074
rect -4413 5058 -4399 5074
rect -4399 5058 -4382 5074
rect -4382 5058 -4357 5074
rect -4493 5022 -4468 5028
rect -4468 5022 -4451 5028
rect -4451 5022 -4437 5028
rect -4413 5022 -4399 5028
rect -4399 5022 -4382 5028
rect -4382 5022 -4357 5028
rect -4493 5010 -4437 5022
rect -4413 5010 -4357 5022
rect -4493 4972 -4468 5010
rect -4468 4972 -4451 5010
rect -4451 4972 -4437 5010
rect -4413 4972 -4399 5010
rect -4399 4972 -4382 5010
rect -4382 4972 -4357 5010
rect -4493 4886 -4437 4942
rect -4413 4886 -4357 4942
rect -4493 4800 -4437 4856
rect -4413 4800 -4357 4856
rect -4493 4714 -4437 4770
rect -4413 4714 -4357 4770
rect -4493 4628 -4437 4684
rect -4413 4628 -4357 4684
rect -4493 4542 -4437 4598
rect -4413 4542 -4357 4598
rect 1844 5322 1900 5378
rect 1844 5235 1900 5291
rect 1844 5148 1900 5204
rect 1844 5061 1900 5117
rect 3989 5305 4045 5361
rect 4084 5305 4140 5361
rect 4179 5305 4235 5361
rect 4273 5305 4329 5361
rect 3989 5225 4045 5281
rect 4084 5225 4140 5281
rect 4179 5225 4235 5281
rect 4273 5225 4329 5281
rect 3989 5145 4045 5201
rect 4084 5145 4140 5201
rect 4179 5145 4235 5201
rect 4273 5145 4329 5201
rect 3989 5065 4045 5121
rect 4084 5065 4140 5121
rect 4179 5065 4235 5121
rect 4273 5065 4329 5121
rect 6485 5322 6541 5378
rect 6485 5235 6541 5291
rect 6485 5148 6541 5204
rect 6485 5061 6541 5117
rect 1844 4974 1900 5030
rect 1844 4887 1900 4943
rect 1844 4800 1900 4856
rect 1844 4713 1900 4769
rect 1844 4626 1900 4682
rect 1844 4538 1900 4594
rect 6485 4974 6541 5030
rect 6485 4887 6541 4943
rect 6485 4800 6541 4856
rect 6485 4713 6541 4769
rect 6485 4626 6541 4682
rect 6485 4538 6541 4594
rect 7603 5282 7659 5338
rect 7685 5282 7741 5338
rect 7767 5282 7823 5338
rect 7848 5282 7904 5338
rect 7929 5282 7985 5338
rect 8010 5282 8066 5338
rect 7603 5200 7659 5256
rect 7685 5200 7741 5256
rect 7767 5200 7823 5256
rect 7848 5200 7904 5256
rect 7929 5200 7985 5256
rect 8010 5200 8066 5256
rect 7603 5118 7659 5174
rect 7685 5118 7741 5174
rect 7767 5118 7823 5174
rect 7848 5118 7904 5174
rect 7929 5118 7985 5174
rect 8010 5118 8066 5174
rect 7603 5036 7659 5092
rect 7685 5036 7741 5092
rect 7767 5036 7823 5092
rect 7848 5036 7904 5092
rect 7929 5036 7985 5092
rect 8010 5036 8066 5092
rect 7603 4954 7659 5010
rect 7685 4954 7741 5010
rect 7767 4954 7823 5010
rect 7848 4954 7904 5010
rect 7929 4954 7985 5010
rect 8010 4954 8066 5010
rect 7603 4872 7659 4928
rect 7685 4872 7741 4928
rect 7767 4872 7823 4928
rect 7848 4872 7904 4928
rect 7929 4872 7985 4928
rect 8010 4872 8066 4928
rect 7603 4790 7659 4846
rect 7685 4790 7741 4846
rect 7767 4790 7823 4846
rect 7848 4790 7904 4846
rect 7929 4790 7985 4846
rect 8010 4790 8066 4846
rect 7603 4708 7659 4764
rect 7685 4708 7741 4764
rect 7767 4708 7823 4764
rect 7848 4708 7904 4764
rect 7929 4708 7985 4764
rect 8010 4708 8066 4764
rect 7603 4626 7659 4682
rect 7685 4626 7741 4682
rect 7767 4626 7823 4682
rect 7848 4626 7904 4682
rect 7929 4626 7985 4682
rect 8010 4626 8066 4682
rect 8274 5315 8330 5371
rect 8274 5235 8330 5291
rect 8274 5155 8330 5211
rect 8274 5075 8330 5131
rect 8274 4995 8330 5051
rect 8274 4915 8330 4971
rect 8274 4835 8330 4891
rect 8274 4754 8330 4810
rect 8274 4673 8330 4729
rect 8686 5315 8742 5371
rect 8686 5235 8742 5291
rect 8686 5155 8742 5211
rect 8686 5075 8742 5131
rect 8686 4995 8742 5051
rect 8686 4915 8742 4971
rect 8686 4835 8742 4891
rect 8686 4754 8742 4810
rect 8686 4673 8742 4729
rect 7603 4544 7659 4600
rect 7685 4544 7741 4600
rect 7767 4544 7823 4600
rect 7848 4544 7904 4600
rect 7929 4544 7985 4600
rect 8010 4544 8066 4600
rect -2657 4004 -2601 4016
rect -2657 3960 -2648 4004
rect -2648 3960 -2601 4004
rect -2577 3960 -2521 4016
rect -2497 3960 -2441 4016
rect -2417 3960 -2361 4016
rect -2657 3886 -2648 3930
rect -2648 3886 -2601 3930
rect -2657 3874 -2601 3886
rect -2577 3874 -2521 3930
rect -2497 3874 -2441 3930
rect -2417 3874 -2361 3930
rect -2657 3820 -2648 3844
rect -2648 3820 -2601 3844
rect -2657 3806 -2601 3820
rect -2657 3788 -2648 3806
rect -2648 3788 -2601 3806
rect -2577 3788 -2521 3844
rect -2497 3788 -2441 3844
rect -2417 3788 -2361 3844
rect -2657 3754 -2648 3758
rect -2648 3754 -2601 3758
rect -2657 3740 -2601 3754
rect -2657 3702 -2648 3740
rect -2648 3702 -2601 3740
rect -2577 3702 -2521 3758
rect -2497 3702 -2441 3758
rect -2417 3702 -2361 3758
rect -2657 3623 -2648 3672
rect -2648 3623 -2601 3672
rect -2657 3616 -2601 3623
rect -2577 3616 -2521 3672
rect -2497 3616 -2441 3672
rect -2417 3616 -2361 3672
rect -2657 3530 -2601 3586
rect -2577 3530 -2521 3586
rect -2497 3530 -2441 3586
rect -2417 3530 -2361 3586
rect -2657 3444 -2601 3500
rect -2577 3444 -2521 3500
rect -2497 3444 -2441 3500
rect -2417 3444 -2361 3500
rect -2657 3358 -2601 3414
rect -2577 3358 -2521 3414
rect -2497 3358 -2441 3414
rect -2417 3358 -2361 3414
rect -2657 3271 -2601 3327
rect -2577 3271 -2521 3327
rect -2497 3271 -2441 3327
rect -2417 3271 -2361 3327
rect -2657 3184 -2601 3240
rect -2577 3184 -2521 3240
rect -2497 3184 -2441 3240
rect -2417 3184 -2361 3240
<< metal3 >>
rect 11668 8173 11810 8178
rect 11668 8117 11711 8173
rect 11767 8117 11810 8173
rect 11668 8080 11810 8117
rect 11668 8024 11711 8080
rect 11767 8024 11810 8080
rect 11668 7987 11810 8024
rect 11668 7931 11711 7987
rect 11767 7931 11810 7987
rect 11668 7894 11810 7931
rect 11668 7838 11711 7894
rect 11767 7838 11810 7894
rect -4531 7812 -4319 7817
rect -4531 7756 -4493 7812
rect -4437 7756 -4413 7812
rect -4357 7756 -4319 7812
rect -4531 7728 -4319 7756
rect 11668 7800 11810 7838
rect 11668 7744 11711 7800
rect 11767 7744 11810 7800
rect -4531 7672 -4493 7728
rect -4437 7672 -4413 7728
rect -4357 7672 -4319 7728
tri 11634 7706 11668 7740 se
rect 11668 7706 11810 7744
rect -4531 7644 -4319 7672
rect -4531 7588 -4493 7644
rect -4437 7588 -4413 7644
rect -4357 7588 -4319 7644
rect -4531 7559 -4319 7588
rect -4531 7503 -4493 7559
rect -4437 7503 -4413 7559
rect -4357 7503 -4319 7559
rect -4531 7474 -4319 7503
rect -4531 7418 -4493 7474
rect -4437 7418 -4413 7474
rect -4357 7418 -4319 7474
rect -4531 7389 -4319 7418
rect -4531 7333 -4493 7389
rect -4437 7333 -4413 7389
rect -4357 7333 -4319 7389
rect -4531 7328 -4319 7333
tri 11626 7698 11634 7706 se
rect 11634 7698 11711 7706
rect 11626 7650 11711 7698
rect 11767 7650 11810 7706
rect 11626 7645 11810 7650
rect 11626 7602 11692 7645
tri 11692 7607 11730 7645 nw
rect 11626 7546 11631 7602
rect 11687 7546 11692 7602
rect 11626 7497 11692 7546
rect 11626 7441 11631 7497
rect 11687 7441 11692 7497
rect 11626 7392 11692 7441
rect 11626 7336 11631 7392
rect 11687 7336 11692 7392
rect 11626 7331 11692 7336
rect 73 6399 139 6404
rect 73 6343 78 6399
rect 134 6343 139 6399
rect 73 6316 139 6343
rect 73 6260 78 6316
rect 134 6260 139 6316
rect 73 6233 139 6260
rect 73 6177 78 6233
rect 134 6177 139 6233
rect 73 6150 139 6177
rect 73 6094 78 6150
rect 134 6094 139 6150
rect 73 6067 139 6094
rect 73 6011 78 6067
rect 134 6011 139 6067
rect 73 5984 139 6011
rect 73 5928 78 5984
rect 134 5928 139 5984
rect 73 5923 139 5928
rect 1836 5378 1908 5383
rect -4531 5370 -4319 5375
rect -4531 5314 -4493 5370
rect -4437 5314 -4413 5370
rect -4357 5314 -4319 5370
rect -4531 5285 -4319 5314
rect -4531 5229 -4493 5285
rect -4437 5229 -4413 5285
rect -4357 5229 -4319 5285
rect -4531 5200 -4319 5229
rect -4531 5144 -4493 5200
rect -4437 5144 -4413 5200
rect -4357 5144 -4319 5200
rect -4531 5114 -4319 5144
rect -4531 5058 -4493 5114
rect -4437 5058 -4413 5114
rect -4357 5058 -4319 5114
rect -4531 5028 -4319 5058
rect -4531 4972 -4493 5028
rect -4437 4972 -4413 5028
rect -4357 4972 -4319 5028
rect -4531 4942 -4319 4972
rect -4531 4886 -4493 4942
rect -4437 4886 -4413 4942
rect -4357 4886 -4319 4942
rect -4531 4856 -4319 4886
rect -4531 4800 -4493 4856
rect -4437 4800 -4413 4856
rect -4357 4800 -4319 4856
rect -4531 4770 -4319 4800
rect -4531 4714 -4493 4770
rect -4437 4714 -4413 4770
rect -4357 4714 -4319 4770
rect -4531 4684 -4319 4714
rect -4531 4628 -4493 4684
rect -4437 4628 -4413 4684
rect -4357 4628 -4319 4684
rect -4531 4598 -4319 4628
rect -4531 4542 -4493 4598
rect -4437 4542 -4413 4598
rect -4357 4542 -4319 4598
rect -4531 4537 -4319 4542
rect 1836 5322 1844 5378
rect 1900 5322 1908 5378
rect 1836 5291 1908 5322
rect 1836 5235 1844 5291
rect 1900 5235 1908 5291
rect 1836 5204 1908 5235
rect 1836 5148 1844 5204
rect 1900 5148 1908 5204
rect 1836 5117 1908 5148
rect 1836 5061 1844 5117
rect 1900 5061 1908 5117
rect 1836 5030 1908 5061
rect 3984 5361 4334 5386
rect 3984 5305 3989 5361
rect 4045 5305 4084 5361
rect 4140 5305 4179 5361
rect 4235 5305 4273 5361
rect 4329 5305 4334 5361
rect 3984 5281 4334 5305
rect 3984 5225 3989 5281
rect 4045 5225 4084 5281
rect 4140 5225 4179 5281
rect 4235 5225 4273 5281
rect 4329 5225 4334 5281
rect 3984 5201 4334 5225
rect 3984 5145 3989 5201
rect 4045 5145 4084 5201
rect 4140 5145 4179 5201
rect 4235 5145 4273 5201
rect 4329 5145 4334 5201
rect 3984 5121 4334 5145
rect 3984 5065 3989 5121
rect 4045 5065 4084 5121
rect 4140 5065 4179 5121
rect 4235 5065 4273 5121
rect 4329 5065 4334 5121
rect 3984 5040 4334 5065
rect 6468 5378 6558 5383
rect 6468 5322 6485 5378
rect 6541 5322 6558 5378
rect 8235 5371 8369 5376
rect 6468 5291 6558 5322
rect 6468 5235 6485 5291
rect 6541 5235 6558 5291
rect 6468 5204 6558 5235
rect 6468 5148 6485 5204
rect 6541 5148 6558 5204
rect 6468 5117 6558 5148
rect 6468 5061 6485 5117
rect 6541 5061 6558 5117
rect 1836 4974 1844 5030
rect 1900 4974 1908 5030
rect 1836 4943 1908 4974
rect 1836 4887 1844 4943
rect 1900 4887 1908 4943
rect 1836 4856 1908 4887
rect 1836 4800 1844 4856
rect 1900 4800 1908 4856
rect 1836 4769 1908 4800
rect 1836 4713 1844 4769
rect 1900 4713 1908 4769
rect 1836 4682 1908 4713
rect 1836 4626 1844 4682
rect 1900 4626 1908 4682
rect 1836 4594 1908 4626
rect 1836 4538 1844 4594
rect 1900 4538 1908 4594
rect 1836 4533 1908 4538
rect 6468 5030 6558 5061
rect 6468 4974 6485 5030
rect 6541 4974 6558 5030
rect 6468 4943 6558 4974
rect 6468 4887 6485 4943
rect 6541 4887 6558 4943
rect 6468 4856 6558 4887
rect 6468 4800 6485 4856
rect 6541 4800 6558 4856
rect 6468 4769 6558 4800
rect 6468 4713 6485 4769
rect 6541 4713 6558 4769
rect 6468 4682 6558 4713
rect 6468 4626 6485 4682
rect 6541 4626 6558 4682
rect 6468 4594 6558 4626
rect 6468 4538 6485 4594
rect 6541 4538 6558 4594
rect 6468 4533 6558 4538
rect 7598 5338 8071 5351
rect 7598 5282 7603 5338
rect 7659 5282 7685 5338
rect 7741 5282 7767 5338
rect 7823 5282 7848 5338
rect 7904 5282 7929 5338
rect 7985 5282 8010 5338
rect 8066 5282 8071 5338
rect 7598 5256 8071 5282
rect 7598 5200 7603 5256
rect 7659 5200 7685 5256
rect 7741 5200 7767 5256
rect 7823 5200 7848 5256
rect 7904 5200 7929 5256
rect 7985 5200 8010 5256
rect 8066 5200 8071 5256
rect 7598 5174 8071 5200
rect 7598 5118 7603 5174
rect 7659 5118 7685 5174
rect 7741 5118 7767 5174
rect 7823 5118 7848 5174
rect 7904 5118 7929 5174
rect 7985 5118 8010 5174
rect 8066 5118 8071 5174
rect 7598 5092 8071 5118
rect 7598 5036 7603 5092
rect 7659 5036 7685 5092
rect 7741 5036 7767 5092
rect 7823 5036 7848 5092
rect 7904 5036 7929 5092
rect 7985 5036 8010 5092
rect 8066 5036 8071 5092
rect 7598 5010 8071 5036
rect 7598 4954 7603 5010
rect 7659 4954 7685 5010
rect 7741 4954 7767 5010
rect 7823 4954 7848 5010
rect 7904 4954 7929 5010
rect 7985 4954 8010 5010
rect 8066 4954 8071 5010
rect 7598 4928 8071 4954
rect 7598 4872 7603 4928
rect 7659 4872 7685 4928
rect 7741 4872 7767 4928
rect 7823 4872 7848 4928
rect 7904 4872 7929 4928
rect 7985 4872 8010 4928
rect 8066 4872 8071 4928
rect 7598 4846 8071 4872
rect 7598 4790 7603 4846
rect 7659 4790 7685 4846
rect 7741 4790 7767 4846
rect 7823 4790 7848 4846
rect 7904 4790 7929 4846
rect 7985 4790 8010 4846
rect 8066 4790 8071 4846
rect 7598 4764 8071 4790
rect 7598 4708 7603 4764
rect 7659 4708 7685 4764
rect 7741 4708 7767 4764
rect 7823 4708 7848 4764
rect 7904 4708 7929 4764
rect 7985 4708 8010 4764
rect 8066 4708 8071 4764
rect 7598 4682 8071 4708
rect 7598 4626 7603 4682
rect 7659 4626 7685 4682
rect 7741 4626 7767 4682
rect 7823 4626 7848 4682
rect 7904 4626 7929 4682
rect 7985 4626 8010 4682
rect 8066 4626 8071 4682
rect 8235 5315 8274 5371
rect 8330 5315 8369 5371
rect 8235 5291 8369 5315
rect 8235 5235 8274 5291
rect 8330 5235 8369 5291
rect 8235 5211 8369 5235
rect 8235 5155 8274 5211
rect 8330 5155 8369 5211
rect 8235 5131 8369 5155
rect 8235 5075 8274 5131
rect 8330 5075 8369 5131
rect 8235 5051 8369 5075
rect 8235 4995 8274 5051
rect 8330 4995 8369 5051
rect 8235 4971 8369 4995
rect 8235 4915 8274 4971
rect 8330 4915 8369 4971
rect 8235 4891 8369 4915
rect 8235 4835 8274 4891
rect 8330 4835 8369 4891
rect 8235 4810 8369 4835
rect 8235 4754 8274 4810
rect 8330 4754 8369 4810
rect 8235 4729 8369 4754
rect 8235 4673 8274 4729
rect 8330 4673 8369 4729
rect 8235 4668 8369 4673
rect 8647 5371 8781 5376
rect 8647 5315 8686 5371
rect 8742 5315 8781 5371
rect 8647 5291 8781 5315
rect 8647 5235 8686 5291
rect 8742 5235 8781 5291
rect 8647 5211 8781 5235
rect 8647 5155 8686 5211
rect 8742 5155 8781 5211
rect 8647 5131 8781 5155
rect 8647 5075 8686 5131
rect 8742 5075 8781 5131
rect 8647 5051 8781 5075
rect 8647 4995 8686 5051
rect 8742 4995 8781 5051
rect 8647 4971 8781 4995
rect 8647 4915 8686 4971
rect 8742 4915 8781 4971
rect 8647 4891 8781 4915
rect 8647 4835 8686 4891
rect 8742 4835 8781 4891
rect 8647 4810 8781 4835
rect 8647 4754 8686 4810
rect 8742 4754 8781 4810
rect 8647 4729 8781 4754
rect 8647 4673 8686 4729
rect 8742 4673 8781 4729
rect 8647 4668 8781 4673
rect 7598 4600 8071 4626
rect 7598 4544 7603 4600
rect 7659 4544 7685 4600
rect 7741 4544 7767 4600
rect 7823 4544 7848 4600
rect 7904 4544 7929 4600
rect 7985 4544 8010 4600
rect 8066 4544 8071 4600
rect 7598 4531 8071 4544
rect -2669 4016 -2349 4021
rect -2669 3960 -2657 4016
rect -2601 3960 -2577 4016
rect -2521 3960 -2497 4016
rect -2441 3960 -2417 4016
rect -2361 3960 -2349 4016
rect -2669 3930 -2349 3960
rect -2669 3874 -2657 3930
rect -2601 3874 -2577 3930
rect -2521 3874 -2497 3930
rect -2441 3874 -2417 3930
rect -2361 3874 -2349 3930
rect -2669 3844 -2349 3874
rect -2669 3788 -2657 3844
rect -2601 3788 -2577 3844
rect -2521 3788 -2497 3844
rect -2441 3788 -2417 3844
rect -2361 3788 -2349 3844
rect -2669 3758 -2349 3788
rect -2669 3702 -2657 3758
rect -2601 3702 -2577 3758
rect -2521 3702 -2497 3758
rect -2441 3702 -2417 3758
rect -2361 3702 -2349 3758
rect -2669 3672 -2349 3702
rect -2669 3616 -2657 3672
rect -2601 3616 -2577 3672
rect -2521 3616 -2497 3672
rect -2441 3616 -2417 3672
rect -2361 3616 -2349 3672
rect -2669 3586 -2349 3616
rect -2669 3530 -2657 3586
rect -2601 3530 -2577 3586
rect -2521 3530 -2497 3586
rect -2441 3530 -2417 3586
rect -2361 3530 -2349 3586
rect -2669 3500 -2349 3530
rect -2669 3444 -2657 3500
rect -2601 3444 -2577 3500
rect -2521 3444 -2497 3500
rect -2441 3444 -2417 3500
rect -2361 3444 -2349 3500
rect -2669 3414 -2349 3444
rect -2669 3358 -2657 3414
rect -2601 3358 -2577 3414
rect -2521 3358 -2497 3414
rect -2441 3358 -2417 3414
rect -2361 3358 -2349 3414
rect -2669 3327 -2349 3358
rect -2669 3271 -2657 3327
rect -2601 3271 -2577 3327
rect -2521 3271 -2497 3327
rect -2441 3271 -2417 3327
rect -2361 3271 -2349 3327
rect -2669 3240 -2349 3271
rect -2669 3184 -2657 3240
rect -2601 3184 -2577 3240
rect -2521 3184 -2497 3240
rect -2441 3184 -2417 3240
rect -2361 3184 -2349 3240
rect -2669 3179 -2349 3184
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 1 0 -1229 0 1 8659
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 1 0 -1229 0 1 8307
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 1 0 11674 0 1 8956
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1704896540
transform 1 0 -2195 0 1 1569
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1704896540
transform 1 0 -646 0 1 8230
box 0 0 320 116
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1704896540
transform 1 0 -1647 0 1 8217
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform 0 1 -410 1 0 3714
box 0 0 1 1
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_0
timestamp 1704896540
transform 1 0 -3217 0 1 11394
box 0 0 384 180
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_0
timestamp 1704896540
transform 1 0 8983 0 1 4559
box -5 0 301 794
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_1
timestamp 1704896540
transform 1 0 9667 0 1 7358
box -5 0 301 794
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_2
timestamp 1704896540
transform 1 0 220 0 1 7358
box -5 0 301 794
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_3
timestamp 1704896540
transform 1 0 217 0 1 4563
box -5 0 301 794
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_4
timestamp 1704896540
transform 1 0 10338 0 1 4559
box -5 0 301 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_0
timestamp 1704896540
transform 1 0 -3979 0 1 1835
box -5 0 61 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_0
timestamp 1704896540
transform 1 0 11879 0 1 7354
box -5 0 141 794
use M2M3_CDNS_524688791851238  M2M3_CDNS_524688791851238_0
timestamp 1704896540
transform 1 0 -1485 0 1 7674
box -5 0 221 314
use sky130_fd_io__sio_in_diff  sky130_fd_io__sio_in_diff_0
timestamp 1704896540
transform 1 0 -2988 0 1 1240
box -87 -593 16858 13583
use sky130_fd_io__sio_in_diff_ctlblk_tsg4  sky130_fd_io__sio_in_diff_ctlblk_tsg4_0
timestamp 1704896540
transform 1 0 -4671 0 1 1052
box -1642 112 5255 9328
<< labels >>
flabel metal1 s -371 12528 -51 12576 0 FreeSans 400 180 0 0 vcc_io
port 2 nsew
flabel metal1 s -459 12110 -139 12158 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal1 s 4837 6874 5157 6922 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal1 s 7753 10254 8073 10300 0 FreeSans 400 0 0 0 vpwr_ka
port 4 nsew
flabel metal1 s 12128 14692 12448 14738 0 FreeSans 400 0 0 0 vpwr_ka
port 4 nsew
flabel metal1 s -4704 1956 -4667 1996 7 FreeSans 400 0 0 0 out_n
port 6 nsew
flabel metal1 s -4982 2587 -4944 2633 7 FreeSans 400 0 0 0 out_h_n
port 5 nsew
flabel metal1 s -4867 3024 -4813 3058 3 FreeSans 200 0 0 0 ie_diff_sel_h_n
port 7 nsew
flabel metal1 s -4783 3086 -4755 3120 3 FreeSans 200 0 0 0 ie_diff_sel_h
port 8 nsew
flabel metal1 s 13513 6346 13565 6397 0 FreeSans 400 180 0 0 vinref
port 9 nsew
flabel metal1 s -4700 6992 -4666 7029 7 FreeSans 200 180 0 0 sio_diff_hyst_en_h
port 10 nsew
flabel metal1 s -1256 14201 -937 14247 0 FreeSans 400 0 0 0 vpwr_ka
port 4 nsew
flabel metal1 s -4099 7713 -4073 7755 3 FreeSans 200 0 0 0 ie_diff_sel_n
port 11 nsew
flabel metal1 s -283 8208 -211 8362 0 FreeSans 400 180 0 0 pad_esd
port 12 nsew
flabel metal2 s -4041 9915 -3721 9961 0 FreeSans 400 0 0 0 vpwr_ka
port 4 nsew
flabel metal2 s -3565 9915 -3245 9961 0 FreeSans 400 0 0 0 vpb_ka
port 13 nsew
flabel metal2 s 8489 6651 8809 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s -1864 7507 -1545 7555 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 8132 6651 8330 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 7498 6651 7891 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 6378 6651 7035 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 5193 6651 6150 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 4399 6651 5082 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 3975 6651 4343 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 3148 6651 3720 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 2349 6651 3040 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s 762 6683 1082 6745 0 FreeSans 400 180 0 0 vgnd
port 3 nsew
flabel metal2 s -614 6697 -294 6745 0 FreeSans 400 180 0 0 vcc_ioq
port 14 nsew
flabel metal2 s -962 6697 -642 6745 0 FreeSans 400 180 0 0 vcc_ioq
port 14 nsew
flabel metal2 s -2667 7507 -2167 7555 0 FreeSans 400 180 0 0 vcc_ioq
port 14 nsew
flabel metal2 s 11057 11640 11377 11734 0 FreeSans 400 180 0 0 vcc_ioq
port 14 nsew
flabel metal2 s 1430 6651 1729 6746 0 FreeSans 400 180 0 0 vcc_io
port 2 nsew
flabel metal2 s 9068 11640 9542 11734 0 FreeSans 400 180 0 0 vcc_io
port 2 nsew
flabel metal2 s -4526 7795 -4324 7821 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal2 s 13155 11691 13506 11734 0 FreeSans 400 0 0 0 vpwr_ka
port 4 nsew
<< properties >>
string GDS_END 87493054
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87459488
string path 291.475 183.275 291.475 190.175 
<< end >>
