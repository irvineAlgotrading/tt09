magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 10 66 1016 720
<< mvnmos >>
rect 228 92 328 694
rect 384 92 484 694
rect 540 92 640 694
rect 696 92 796 694
<< mvndiff >>
rect 172 682 228 694
rect 172 648 183 682
rect 217 648 228 682
rect 172 614 228 648
rect 172 580 183 614
rect 217 580 228 614
rect 172 546 228 580
rect 172 512 183 546
rect 217 512 228 546
rect 172 478 228 512
rect 172 444 183 478
rect 217 444 228 478
rect 172 410 228 444
rect 172 376 183 410
rect 217 376 228 410
rect 172 342 228 376
rect 172 308 183 342
rect 217 308 228 342
rect 172 274 228 308
rect 172 240 183 274
rect 217 240 228 274
rect 172 206 228 240
rect 172 172 183 206
rect 217 172 228 206
rect 172 138 228 172
rect 172 104 183 138
rect 217 104 228 138
rect 172 92 228 104
rect 328 682 384 694
rect 328 648 339 682
rect 373 648 384 682
rect 328 614 384 648
rect 328 580 339 614
rect 373 580 384 614
rect 328 546 384 580
rect 328 512 339 546
rect 373 512 384 546
rect 328 478 384 512
rect 328 444 339 478
rect 373 444 384 478
rect 328 410 384 444
rect 328 376 339 410
rect 373 376 384 410
rect 328 342 384 376
rect 328 308 339 342
rect 373 308 384 342
rect 328 274 384 308
rect 328 240 339 274
rect 373 240 384 274
rect 328 206 384 240
rect 328 172 339 206
rect 373 172 384 206
rect 328 138 384 172
rect 328 104 339 138
rect 373 104 384 138
rect 328 92 384 104
rect 484 682 540 694
rect 484 648 495 682
rect 529 648 540 682
rect 484 614 540 648
rect 484 580 495 614
rect 529 580 540 614
rect 484 546 540 580
rect 484 512 495 546
rect 529 512 540 546
rect 484 478 540 512
rect 484 444 495 478
rect 529 444 540 478
rect 484 410 540 444
rect 484 376 495 410
rect 529 376 540 410
rect 484 342 540 376
rect 484 308 495 342
rect 529 308 540 342
rect 484 274 540 308
rect 484 240 495 274
rect 529 240 540 274
rect 484 206 540 240
rect 484 172 495 206
rect 529 172 540 206
rect 484 138 540 172
rect 484 104 495 138
rect 529 104 540 138
rect 484 92 540 104
rect 640 682 696 694
rect 640 648 651 682
rect 685 648 696 682
rect 640 614 696 648
rect 640 580 651 614
rect 685 580 696 614
rect 640 546 696 580
rect 640 512 651 546
rect 685 512 696 546
rect 640 478 696 512
rect 640 444 651 478
rect 685 444 696 478
rect 640 410 696 444
rect 640 376 651 410
rect 685 376 696 410
rect 640 342 696 376
rect 640 308 651 342
rect 685 308 696 342
rect 640 274 696 308
rect 640 240 651 274
rect 685 240 696 274
rect 640 206 696 240
rect 640 172 651 206
rect 685 172 696 206
rect 640 138 696 172
rect 640 104 651 138
rect 685 104 696 138
rect 640 92 696 104
rect 796 682 852 694
rect 796 648 807 682
rect 841 648 852 682
rect 796 614 852 648
rect 796 580 807 614
rect 841 580 852 614
rect 796 546 852 580
rect 796 512 807 546
rect 841 512 852 546
rect 796 478 852 512
rect 796 444 807 478
rect 841 444 852 478
rect 796 410 852 444
rect 796 376 807 410
rect 841 376 852 410
rect 796 342 852 376
rect 796 308 807 342
rect 841 308 852 342
rect 796 274 852 308
rect 796 240 807 274
rect 841 240 852 274
rect 796 206 852 240
rect 796 172 807 206
rect 841 172 852 206
rect 796 138 852 172
rect 796 104 807 138
rect 841 104 852 138
rect 796 92 852 104
<< mvndiffc >>
rect 183 648 217 682
rect 183 580 217 614
rect 183 512 217 546
rect 183 444 217 478
rect 183 376 217 410
rect 183 308 217 342
rect 183 240 217 274
rect 183 172 217 206
rect 183 104 217 138
rect 339 648 373 682
rect 339 580 373 614
rect 339 512 373 546
rect 339 444 373 478
rect 339 376 373 410
rect 339 308 373 342
rect 339 240 373 274
rect 339 172 373 206
rect 339 104 373 138
rect 495 648 529 682
rect 495 580 529 614
rect 495 512 529 546
rect 495 444 529 478
rect 495 376 529 410
rect 495 308 529 342
rect 495 240 529 274
rect 495 172 529 206
rect 495 104 529 138
rect 651 648 685 682
rect 651 580 685 614
rect 651 512 685 546
rect 651 444 685 478
rect 651 376 685 410
rect 651 308 685 342
rect 651 240 685 274
rect 651 172 685 206
rect 651 104 685 138
rect 807 648 841 682
rect 807 580 841 614
rect 807 512 841 546
rect 807 444 841 478
rect 807 376 841 410
rect 807 308 841 342
rect 807 240 841 274
rect 807 172 841 206
rect 807 104 841 138
<< mvpsubdiff >>
rect 36 648 94 694
rect 36 614 48 648
rect 82 614 94 648
rect 36 580 94 614
rect 36 546 48 580
rect 82 546 94 580
rect 36 512 94 546
rect 36 478 48 512
rect 82 478 94 512
rect 36 444 94 478
rect 36 410 48 444
rect 82 410 94 444
rect 36 376 94 410
rect 36 342 48 376
rect 82 342 94 376
rect 36 308 94 342
rect 36 274 48 308
rect 82 274 94 308
rect 36 240 94 274
rect 36 206 48 240
rect 82 206 94 240
rect 36 172 94 206
rect 36 138 48 172
rect 82 138 94 172
rect 36 92 94 138
rect 932 648 990 694
rect 932 614 944 648
rect 978 614 990 648
rect 932 580 990 614
rect 932 546 944 580
rect 978 546 990 580
rect 932 512 990 546
rect 932 478 944 512
rect 978 478 990 512
rect 932 444 990 478
rect 932 410 944 444
rect 978 410 990 444
rect 932 376 990 410
rect 932 342 944 376
rect 978 342 990 376
rect 932 308 990 342
rect 932 274 944 308
rect 978 274 990 308
rect 932 240 990 274
rect 932 206 944 240
rect 978 206 990 240
rect 932 172 990 206
rect 932 138 944 172
rect 978 138 990 172
rect 932 92 990 138
<< mvpsubdiffcont >>
rect 48 614 82 648
rect 48 546 82 580
rect 48 478 82 512
rect 48 410 82 444
rect 48 342 82 376
rect 48 274 82 308
rect 48 206 82 240
rect 48 138 82 172
rect 944 614 978 648
rect 944 546 978 580
rect 944 478 978 512
rect 944 410 978 444
rect 944 342 978 376
rect 944 274 978 308
rect 944 206 978 240
rect 944 138 978 172
<< poly >>
rect 207 766 817 786
rect 207 732 223 766
rect 257 732 291 766
rect 325 732 359 766
rect 393 732 427 766
rect 461 732 495 766
rect 529 732 563 766
rect 597 732 631 766
rect 665 732 699 766
rect 733 732 767 766
rect 801 732 817 766
rect 207 716 817 732
rect 228 694 328 716
rect 384 694 484 716
rect 540 694 640 716
rect 696 694 796 716
rect 228 70 328 92
rect 384 70 484 92
rect 540 70 640 92
rect 696 70 796 92
rect 207 54 817 70
rect 207 20 223 54
rect 257 20 291 54
rect 325 20 359 54
rect 393 20 427 54
rect 461 20 495 54
rect 529 20 563 54
rect 597 20 631 54
rect 665 20 699 54
rect 733 20 767 54
rect 801 20 817 54
rect 207 0 817 20
<< polycont >>
rect 223 732 257 766
rect 291 732 325 766
rect 359 732 393 766
rect 427 732 461 766
rect 495 732 529 766
rect 563 732 597 766
rect 631 732 665 766
rect 699 732 733 766
rect 767 732 801 766
rect 223 20 257 54
rect 291 20 325 54
rect 359 20 393 54
rect 427 20 461 54
rect 495 20 529 54
rect 563 20 597 54
rect 631 20 665 54
rect 699 20 733 54
rect 767 20 801 54
<< locali >>
rect 207 732 223 766
rect 277 732 291 766
rect 349 732 359 766
rect 421 732 427 766
rect 493 732 495 766
rect 529 732 531 766
rect 597 732 603 766
rect 665 732 675 766
rect 733 732 747 766
rect 801 732 817 766
rect 183 682 217 698
rect 48 662 82 664
rect 48 590 82 614
rect 48 518 82 546
rect 48 446 82 478
rect 48 376 82 410
rect 48 308 82 340
rect 48 240 82 268
rect 48 172 82 196
rect 48 122 82 124
rect 183 614 217 628
rect 183 546 217 556
rect 183 478 217 484
rect 183 410 217 412
rect 183 374 217 376
rect 183 302 217 308
rect 183 230 217 240
rect 183 158 217 172
rect 183 88 217 104
rect 339 682 373 698
rect 339 614 373 628
rect 339 546 373 556
rect 339 478 373 484
rect 339 410 373 412
rect 339 374 373 376
rect 339 302 373 308
rect 339 230 373 240
rect 339 158 373 172
rect 339 88 373 104
rect 495 682 529 698
rect 495 614 529 628
rect 495 546 529 556
rect 495 478 529 484
rect 495 410 529 412
rect 495 374 529 376
rect 495 302 529 308
rect 495 230 529 240
rect 495 158 529 172
rect 495 88 529 104
rect 651 682 685 698
rect 651 614 685 628
rect 651 546 685 556
rect 651 478 685 484
rect 651 410 685 412
rect 651 374 685 376
rect 651 302 685 308
rect 651 230 685 240
rect 651 158 685 172
rect 651 88 685 104
rect 807 682 841 698
rect 807 614 841 628
rect 807 546 841 556
rect 807 478 841 484
rect 807 410 841 412
rect 807 374 841 376
rect 807 302 841 308
rect 807 230 841 240
rect 807 158 841 172
rect 944 662 978 664
rect 944 590 978 614
rect 944 518 978 546
rect 944 446 978 478
rect 944 376 978 410
rect 944 308 978 340
rect 944 240 978 268
rect 944 172 978 196
rect 944 122 978 124
rect 807 88 841 104
rect 207 20 223 54
rect 277 20 291 54
rect 349 20 359 54
rect 421 20 427 54
rect 493 20 495 54
rect 529 20 531 54
rect 597 20 603 54
rect 665 20 675 54
rect 733 20 747 54
rect 801 20 817 54
<< viali >>
rect 243 732 257 766
rect 257 732 277 766
rect 315 732 325 766
rect 325 732 349 766
rect 387 732 393 766
rect 393 732 421 766
rect 459 732 461 766
rect 461 732 493 766
rect 531 732 563 766
rect 563 732 565 766
rect 603 732 631 766
rect 631 732 637 766
rect 675 732 699 766
rect 699 732 709 766
rect 747 732 767 766
rect 767 732 781 766
rect 48 648 82 662
rect 48 628 82 648
rect 48 580 82 590
rect 48 556 82 580
rect 48 512 82 518
rect 48 484 82 512
rect 48 444 82 446
rect 48 412 82 444
rect 48 342 82 374
rect 48 340 82 342
rect 48 274 82 302
rect 48 268 82 274
rect 48 206 82 230
rect 48 196 82 206
rect 48 138 82 158
rect 48 124 82 138
rect 183 648 217 662
rect 183 628 217 648
rect 183 580 217 590
rect 183 556 217 580
rect 183 512 217 518
rect 183 484 217 512
rect 183 444 217 446
rect 183 412 217 444
rect 183 342 217 374
rect 183 340 217 342
rect 183 274 217 302
rect 183 268 217 274
rect 183 206 217 230
rect 183 196 217 206
rect 183 138 217 158
rect 183 124 217 138
rect 339 648 373 662
rect 339 628 373 648
rect 339 580 373 590
rect 339 556 373 580
rect 339 512 373 518
rect 339 484 373 512
rect 339 444 373 446
rect 339 412 373 444
rect 339 342 373 374
rect 339 340 373 342
rect 339 274 373 302
rect 339 268 373 274
rect 339 206 373 230
rect 339 196 373 206
rect 339 138 373 158
rect 339 124 373 138
rect 495 648 529 662
rect 495 628 529 648
rect 495 580 529 590
rect 495 556 529 580
rect 495 512 529 518
rect 495 484 529 512
rect 495 444 529 446
rect 495 412 529 444
rect 495 342 529 374
rect 495 340 529 342
rect 495 274 529 302
rect 495 268 529 274
rect 495 206 529 230
rect 495 196 529 206
rect 495 138 529 158
rect 495 124 529 138
rect 651 648 685 662
rect 651 628 685 648
rect 651 580 685 590
rect 651 556 685 580
rect 651 512 685 518
rect 651 484 685 512
rect 651 444 685 446
rect 651 412 685 444
rect 651 342 685 374
rect 651 340 685 342
rect 651 274 685 302
rect 651 268 685 274
rect 651 206 685 230
rect 651 196 685 206
rect 651 138 685 158
rect 651 124 685 138
rect 807 648 841 662
rect 807 628 841 648
rect 807 580 841 590
rect 807 556 841 580
rect 807 512 841 518
rect 807 484 841 512
rect 807 444 841 446
rect 807 412 841 444
rect 807 342 841 374
rect 807 340 841 342
rect 807 274 841 302
rect 807 268 841 274
rect 807 206 841 230
rect 807 196 841 206
rect 807 138 841 158
rect 807 124 841 138
rect 944 648 978 662
rect 944 628 978 648
rect 944 580 978 590
rect 944 556 978 580
rect 944 512 978 518
rect 944 484 978 512
rect 944 444 978 446
rect 944 412 978 444
rect 944 342 978 374
rect 944 340 978 342
rect 944 274 978 302
rect 944 268 978 274
rect 944 206 978 230
rect 944 196 978 206
rect 944 138 978 158
rect 944 124 978 138
rect 243 20 257 54
rect 257 20 277 54
rect 315 20 325 54
rect 325 20 349 54
rect 387 20 393 54
rect 393 20 421 54
rect 459 20 461 54
rect 461 20 493 54
rect 531 20 563 54
rect 563 20 565 54
rect 603 20 631 54
rect 631 20 637 54
rect 675 20 699 54
rect 699 20 709 54
rect 747 20 767 54
rect 767 20 781 54
<< metal1 >>
rect 231 766 793 786
rect 231 732 243 766
rect 277 732 315 766
rect 349 732 387 766
rect 421 732 459 766
rect 493 732 531 766
rect 565 732 603 766
rect 637 732 675 766
rect 709 732 747 766
rect 781 732 793 766
rect 231 720 793 732
rect 36 662 94 674
rect 36 628 48 662
rect 82 628 94 662
rect 36 590 94 628
rect 36 556 48 590
rect 82 556 94 590
rect 36 518 94 556
rect 36 484 48 518
rect 82 484 94 518
rect 36 446 94 484
rect 36 412 48 446
rect 82 412 94 446
rect 36 374 94 412
rect 36 340 48 374
rect 82 340 94 374
rect 36 302 94 340
rect 36 268 48 302
rect 82 268 94 302
rect 36 230 94 268
rect 36 196 48 230
rect 82 196 94 230
rect 36 158 94 196
rect 36 124 48 158
rect 82 124 94 158
rect 36 112 94 124
rect 174 662 226 674
rect 174 628 183 662
rect 217 628 226 662
rect 174 590 226 628
rect 174 556 183 590
rect 217 556 226 590
rect 174 518 226 556
rect 174 484 183 518
rect 217 484 226 518
rect 174 446 226 484
rect 174 412 183 446
rect 217 412 226 446
rect 174 374 226 412
rect 174 362 183 374
rect 217 362 226 374
rect 174 302 226 310
rect 174 298 183 302
rect 217 298 226 302
rect 174 234 226 246
rect 174 170 226 182
rect 174 112 226 118
rect 330 668 382 674
rect 330 604 382 616
rect 330 540 382 552
rect 330 484 339 488
rect 373 484 382 488
rect 330 476 382 484
rect 330 412 339 424
rect 373 412 382 424
rect 330 374 382 412
rect 330 340 339 374
rect 373 340 382 374
rect 330 302 382 340
rect 330 268 339 302
rect 373 268 382 302
rect 330 230 382 268
rect 330 196 339 230
rect 373 196 382 230
rect 330 158 382 196
rect 330 124 339 158
rect 373 124 382 158
rect 330 112 382 124
rect 486 662 538 674
rect 486 628 495 662
rect 529 628 538 662
rect 486 590 538 628
rect 486 556 495 590
rect 529 556 538 590
rect 486 518 538 556
rect 486 484 495 518
rect 529 484 538 518
rect 486 446 538 484
rect 486 412 495 446
rect 529 412 538 446
rect 486 374 538 412
rect 486 362 495 374
rect 529 362 538 374
rect 486 302 538 310
rect 486 298 495 302
rect 529 298 538 302
rect 486 234 538 246
rect 486 170 538 182
rect 486 112 538 118
rect 642 668 694 674
rect 642 604 694 616
rect 642 540 694 552
rect 642 484 651 488
rect 685 484 694 488
rect 642 476 694 484
rect 642 412 651 424
rect 685 412 694 424
rect 642 374 694 412
rect 642 340 651 374
rect 685 340 694 374
rect 642 302 694 340
rect 642 268 651 302
rect 685 268 694 302
rect 642 230 694 268
rect 642 196 651 230
rect 685 196 694 230
rect 642 158 694 196
rect 642 124 651 158
rect 685 124 694 158
rect 642 112 694 124
rect 798 662 850 674
rect 798 628 807 662
rect 841 628 850 662
rect 798 590 850 628
rect 798 556 807 590
rect 841 556 850 590
rect 798 518 850 556
rect 798 484 807 518
rect 841 484 850 518
rect 798 446 850 484
rect 798 412 807 446
rect 841 412 850 446
rect 798 374 850 412
rect 798 362 807 374
rect 841 362 850 374
rect 798 302 850 310
rect 798 298 807 302
rect 841 298 850 302
rect 798 234 850 246
rect 798 170 850 182
rect 798 112 850 118
rect 932 662 990 674
rect 932 628 944 662
rect 978 628 990 662
rect 932 590 990 628
rect 932 556 944 590
rect 978 556 990 590
rect 932 518 990 556
rect 932 484 944 518
rect 978 484 990 518
rect 932 446 990 484
rect 932 412 944 446
rect 978 412 990 446
rect 932 374 990 412
rect 932 340 944 374
rect 978 340 990 374
rect 932 302 990 340
rect 932 268 944 302
rect 978 268 990 302
rect 932 230 990 268
rect 932 196 944 230
rect 978 196 990 230
rect 932 158 990 196
rect 932 124 944 158
rect 978 124 990 158
rect 932 112 990 124
rect 231 54 793 66
rect 231 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 793 54
rect 231 0 793 20
<< via1 >>
rect 174 340 183 362
rect 183 340 217 362
rect 217 340 226 362
rect 174 310 226 340
rect 174 268 183 298
rect 183 268 217 298
rect 217 268 226 298
rect 174 246 226 268
rect 174 230 226 234
rect 174 196 183 230
rect 183 196 217 230
rect 217 196 226 230
rect 174 182 226 196
rect 174 158 226 170
rect 174 124 183 158
rect 183 124 217 158
rect 217 124 226 158
rect 174 118 226 124
rect 330 662 382 668
rect 330 628 339 662
rect 339 628 373 662
rect 373 628 382 662
rect 330 616 382 628
rect 330 590 382 604
rect 330 556 339 590
rect 339 556 373 590
rect 373 556 382 590
rect 330 552 382 556
rect 330 518 382 540
rect 330 488 339 518
rect 339 488 373 518
rect 373 488 382 518
rect 330 446 382 476
rect 330 424 339 446
rect 339 424 373 446
rect 373 424 382 446
rect 486 340 495 362
rect 495 340 529 362
rect 529 340 538 362
rect 486 310 538 340
rect 486 268 495 298
rect 495 268 529 298
rect 529 268 538 298
rect 486 246 538 268
rect 486 230 538 234
rect 486 196 495 230
rect 495 196 529 230
rect 529 196 538 230
rect 486 182 538 196
rect 486 158 538 170
rect 486 124 495 158
rect 495 124 529 158
rect 529 124 538 158
rect 486 118 538 124
rect 642 662 694 668
rect 642 628 651 662
rect 651 628 685 662
rect 685 628 694 662
rect 642 616 694 628
rect 642 590 694 604
rect 642 556 651 590
rect 651 556 685 590
rect 685 556 694 590
rect 642 552 694 556
rect 642 518 694 540
rect 642 488 651 518
rect 651 488 685 518
rect 685 488 694 518
rect 642 446 694 476
rect 642 424 651 446
rect 651 424 685 446
rect 685 424 694 446
rect 798 340 807 362
rect 807 340 841 362
rect 841 340 850 362
rect 798 310 850 340
rect 798 268 807 298
rect 807 268 841 298
rect 841 268 850 298
rect 798 246 850 268
rect 798 230 850 234
rect 798 196 807 230
rect 807 196 841 230
rect 841 196 850 230
rect 798 182 850 196
rect 798 158 850 170
rect 798 124 807 158
rect 807 124 841 158
rect 841 124 850 158
rect 798 118 850 124
<< metal2 >>
rect 10 668 1016 674
rect 10 616 330 668
rect 382 616 642 668
rect 694 616 1016 668
rect 10 604 1016 616
rect 10 552 330 604
rect 382 552 642 604
rect 694 552 1016 604
rect 10 540 1016 552
rect 10 488 330 540
rect 382 488 642 540
rect 694 488 1016 540
rect 10 476 1016 488
rect 10 424 330 476
rect 382 424 642 476
rect 694 424 1016 476
rect 10 418 1016 424
rect 10 362 1016 368
rect 10 310 174 362
rect 226 310 486 362
rect 538 310 798 362
rect 850 310 1016 362
rect 10 298 1016 310
rect 10 246 174 298
rect 226 246 486 298
rect 538 246 798 298
rect 850 246 1016 298
rect 10 234 1016 246
rect 10 182 174 234
rect 226 182 486 234
rect 538 182 798 234
rect 850 182 1016 234
rect 10 170 1016 182
rect 10 118 174 170
rect 226 118 486 170
rect 538 118 798 170
rect 850 118 1016 170
rect 10 112 1016 118
<< labels >>
flabel comment s 200 393 200 393 0 FreeSans 300 0 0 0 S
flabel comment s 356 393 356 393 0 FreeSans 300 0 0 0 S
flabel comment s 512 393 512 393 0 FreeSans 300 0 0 0 S
flabel comment s 668 393 668 393 0 FreeSans 300 0 0 0 S
flabel comment s 200 393 200 393 0 FreeSans 300 0 0 0 S
flabel comment s 356 393 356 393 0 FreeSans 300 0 0 0 D
flabel comment s 512 393 512 393 0 FreeSans 300 0 0 0 S
flabel comment s 668 393 668 393 0 FreeSans 300 0 0 0 D
flabel comment s 824 393 824 393 0 FreeSans 300 0 0 0 S
flabel metal2 s 32 217 62 321 0 FreeSans 200 0 0 0 SOURCE
port 2 nsew
flabel metal2 s 31 506 66 603 0 FreeSans 200 0 0 0 DRAIN
port 3 nsew
flabel metal1 s 459 730 560 770 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 461 16 559 50 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 951 327 980 433 0 FreeSans 200 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 53 333 81 430 0 FreeSans 200 90 0 0 SUBSTRATE
port 5 nsew
<< properties >>
string GDS_END 7271672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7254022
<< end >>
