magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect 119 369 219 392
rect 119 335 152 369
rect 186 335 219 369
rect 119 274 219 335
rect 119 240 152 274
rect 186 240 219 274
rect 119 218 219 240
rect 275 369 375 392
rect 275 335 309 369
rect 343 335 375 369
rect 275 274 375 335
rect 275 240 309 274
rect 343 240 375 274
rect 275 218 375 240
rect 431 369 531 392
rect 431 335 466 369
rect 500 335 531 369
rect 431 274 531 335
rect 431 240 466 274
rect 500 240 531 274
rect 431 218 531 240
<< polycont >>
rect 152 335 186 369
rect 152 240 186 274
rect 309 335 343 369
rect 309 240 343 274
rect 466 335 500 369
rect 466 240 500 274
<< locali >>
rect 74 556 108 594
rect 386 556 420 594
rect 230 472 264 510
rect 542 472 576 510
rect 152 369 186 385
rect 152 285 186 323
rect 152 224 186 240
rect 309 369 343 385
rect 309 285 343 323
rect 309 224 343 240
rect 466 369 500 385
rect 466 285 500 323
rect 466 224 500 240
rect 542 138 576 176
rect 72 24 110 58
<< viali >>
rect 74 594 108 628
rect 74 522 108 556
rect 386 594 420 628
rect 230 510 264 544
rect 386 522 420 556
rect 230 438 264 472
rect 542 510 576 544
rect 542 438 576 472
rect 152 335 186 357
rect 152 323 186 335
rect 152 274 186 285
rect 152 251 186 274
rect 309 335 343 357
rect 309 323 343 335
rect 309 274 343 285
rect 309 251 343 274
rect 466 335 500 357
rect 466 323 500 335
rect 466 274 500 285
rect 466 251 500 274
rect 542 176 576 210
rect 542 104 576 138
rect 38 24 72 58
rect 110 24 144 58
<< metal1 >>
rect 69 640 426 690
rect 68 628 426 640
rect 68 594 74 628
rect 108 594 386 628
rect 420 594 426 628
rect 68 590 426 594
rect 68 556 114 590
tri 114 556 148 590 nw
tri 346 556 380 590 ne
rect 380 556 426 590
rect 68 522 74 556
rect 108 522 114 556
rect 68 510 114 522
rect 224 544 270 556
rect 224 510 230 544
rect 264 510 270 544
rect 380 522 386 556
rect 420 522 426 556
tri 270 510 272 512 sw
rect 380 510 426 522
rect 536 544 582 556
tri 534 510 536 512 se
rect 536 510 542 544
rect 576 510 582 544
rect 224 478 272 510
tri 272 478 304 510 sw
tri 502 478 534 510 se
rect 534 478 582 510
rect 224 472 582 478
rect 224 438 230 472
rect 264 438 542 472
rect 576 438 582 472
rect 224 426 582 438
tri 502 392 536 426 ne
rect 146 357 192 369
rect 146 323 152 357
rect 186 323 192 357
rect 146 285 192 323
rect 146 251 152 285
rect 186 251 192 285
rect 146 239 192 251
rect 303 357 349 369
rect 303 323 309 357
rect 343 323 349 357
rect 303 285 349 323
rect 303 251 309 285
rect 343 251 349 285
rect 303 239 349 251
rect 460 357 506 369
rect 460 323 466 357
rect 500 323 506 357
rect 460 285 506 323
rect 460 251 466 285
rect 500 251 506 285
rect 460 239 506 251
rect 536 210 582 426
rect 536 176 542 210
rect 576 176 582 210
rect 536 138 582 176
rect 536 104 542 138
rect 576 104 582 138
rect 536 92 582 104
rect 26 58 578 64
rect 26 24 38 58
rect 72 24 110 58
rect 144 24 578 58
rect 26 0 578 24
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_0
timestamp 1704896540
transform 1 0 119 0 1 36
box -82 -32 182 182
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_1
timestamp 1704896540
transform 1 0 275 0 1 36
box -82 -32 182 182
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_2
timestamp 1704896540
transform 1 0 431 0 1 36
box -82 -32 182 182
use pfet_CDNS_52468879185725  pfet_CDNS_52468879185725_0
timestamp 1704896540
transform 1 0 275 0 -1 624
box -119 -66 219 266
use pfet_CDNS_52468879185725  pfet_CDNS_52468879185725_1
timestamp 1704896540
transform 1 0 119 0 -1 624
box -119 -66 219 266
use pfet_CDNS_52468879185725  pfet_CDNS_52468879185725_2
timestamp 1704896540
transform 1 0 431 0 -1 624
box -119 -66 219 266
<< properties >>
string GDS_END 25729876
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25726092
string path 2.275 12.750 2.275 16.000 
<< end >>
