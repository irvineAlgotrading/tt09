magic
tech sky130A
timestamp 1704896540
<< locali >>
rect 0 233 17 252
rect 0 197 17 216
rect 0 161 17 180
rect 0 125 17 144
rect 0 89 17 108
rect 0 53 17 72
rect 0 17 17 36
<< viali >>
rect 0 252 17 269
rect 0 216 17 233
rect 0 180 17 197
rect 0 144 17 161
rect 0 108 17 125
rect 0 72 17 89
rect 0 36 17 53
rect 0 0 17 17
<< metal1 >>
rect -6 269 23 272
rect -6 252 0 269
rect 17 252 23 269
rect -6 233 23 252
rect -6 216 0 233
rect 17 216 23 233
rect -6 197 23 216
rect -6 180 0 197
rect 17 180 23 197
rect -6 161 23 180
rect -6 144 0 161
rect 17 144 23 161
rect -6 125 23 144
rect -6 108 0 125
rect 17 108 23 125
rect -6 89 23 108
rect -6 72 0 89
rect 17 72 23 89
rect -6 53 23 72
rect -6 36 0 53
rect 17 36 23 53
rect -6 17 23 36
rect -6 0 0 17
rect 17 0 23 17
rect -6 -3 23 0
<< properties >>
string GDS_END 95661996
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95661352
<< end >>
