magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< metal1 >>
rect 78 0 114 395
rect 150 0 186 395
rect 222 79 258 420
rect 294 0 330 395
rect 366 0 402 395
rect 846 0 882 395
rect 918 0 954 395
rect 990 79 1026 420
rect 1062 0 1098 395
rect 1134 0 1170 395
rect 1326 0 1362 395
rect 1398 0 1434 395
rect 1470 79 1506 420
rect 1542 0 1578 395
rect 1614 0 1650 395
rect 2094 0 2130 395
rect 2166 0 2202 395
rect 2238 79 2274 420
rect 2310 0 2346 395
rect 2382 0 2418 395
rect 2574 0 2610 395
rect 2646 0 2682 395
rect 2718 79 2754 420
rect 2790 0 2826 395
rect 2862 0 2898 395
rect 3342 0 3378 395
rect 3414 0 3450 395
rect 3486 79 3522 420
rect 3558 0 3594 395
rect 3630 0 3666 395
rect 3822 0 3858 395
rect 3894 0 3930 395
rect 3966 79 4002 420
rect 4038 0 4074 395
rect 4110 0 4146 395
rect 4590 0 4626 395
rect 4662 0 4698 395
rect 4734 79 4770 420
rect 4806 0 4842 395
rect 4878 0 4914 395
rect 5070 0 5106 395
rect 5142 0 5178 395
rect 5214 79 5250 420
rect 5286 0 5322 395
rect 5358 0 5394 395
rect 5838 0 5874 395
rect 5910 0 5946 395
rect 5982 79 6018 420
rect 6054 0 6090 395
rect 6126 0 6162 395
rect 6318 0 6354 395
rect 6390 0 6426 395
rect 6462 79 6498 420
rect 6534 0 6570 395
rect 6606 0 6642 395
rect 7086 0 7122 395
rect 7158 0 7194 395
rect 7230 79 7266 420
rect 7302 0 7338 395
rect 7374 0 7410 395
rect 7566 0 7602 395
rect 7638 0 7674 395
rect 7710 79 7746 420
rect 7782 0 7818 395
rect 7854 0 7890 395
rect 8334 0 8370 395
rect 8406 0 8442 395
rect 8478 79 8514 420
rect 8550 0 8586 395
rect 8622 0 8658 395
rect 8814 0 8850 395
rect 8886 0 8922 395
rect 8958 79 8994 420
rect 9030 0 9066 395
rect 9102 0 9138 395
rect 9582 0 9618 395
rect 9654 0 9690 395
rect 9726 79 9762 420
rect 9798 0 9834 395
rect 9870 0 9906 395
rect 10062 0 10098 395
rect 10134 0 10170 395
rect 10206 79 10242 420
rect 10278 0 10314 395
rect 10350 0 10386 395
rect 10830 0 10866 395
rect 10902 0 10938 395
rect 10974 79 11010 420
rect 11046 0 11082 395
rect 11118 0 11154 395
rect 11310 0 11346 395
rect 11382 0 11418 395
rect 11454 79 11490 420
rect 11526 0 11562 395
rect 11598 0 11634 395
rect 12078 0 12114 395
rect 12150 0 12186 395
rect 12222 79 12258 420
rect 12294 0 12330 395
rect 12366 0 12402 395
rect 12558 0 12594 395
rect 12630 0 12666 395
rect 12702 79 12738 420
rect 12774 0 12810 395
rect 12846 0 12882 395
rect 13326 0 13362 395
rect 13398 0 13434 395
rect 13470 79 13506 420
rect 13542 0 13578 395
rect 13614 0 13650 395
rect 13806 0 13842 395
rect 13878 0 13914 395
rect 13950 79 13986 420
rect 14022 0 14058 395
rect 14094 0 14130 395
rect 14574 0 14610 395
rect 14646 0 14682 395
rect 14718 79 14754 420
rect 14790 0 14826 395
rect 14862 0 14898 395
rect 15054 0 15090 395
rect 15126 0 15162 395
rect 15198 79 15234 420
rect 15270 0 15306 395
rect 15342 0 15378 395
rect 15822 0 15858 395
rect 15894 0 15930 395
rect 15966 79 16002 420
rect 16038 0 16074 395
rect 16110 0 16146 395
rect 16302 0 16338 395
rect 16374 0 16410 395
rect 16446 79 16482 420
rect 16518 0 16554 395
rect 16590 0 16626 395
rect 17070 0 17106 395
rect 17142 0 17178 395
rect 17214 79 17250 420
rect 17286 0 17322 395
rect 17358 0 17394 395
rect 17550 0 17586 395
rect 17622 0 17658 395
rect 17694 79 17730 420
rect 17766 0 17802 395
rect 17838 0 17874 395
rect 18318 0 18354 395
rect 18390 0 18426 395
rect 18462 79 18498 420
rect 18534 0 18570 395
rect 18606 0 18642 395
rect 18798 0 18834 395
rect 18870 0 18906 395
rect 18942 79 18978 420
rect 19014 0 19050 395
rect 19086 0 19122 395
rect 19566 0 19602 395
rect 19638 0 19674 395
rect 19710 79 19746 420
rect 19782 0 19818 395
rect 19854 0 19890 395
rect 20046 0 20082 395
rect 20118 0 20154 395
rect 20190 79 20226 420
rect 20262 0 20298 395
rect 20334 0 20370 395
rect 20814 0 20850 395
rect 20886 0 20922 395
rect 20958 79 20994 420
rect 21030 0 21066 395
rect 21102 0 21138 395
rect 21294 0 21330 395
rect 21366 0 21402 395
rect 21438 79 21474 420
rect 21510 0 21546 395
rect 21582 0 21618 395
rect 22062 0 22098 395
rect 22134 0 22170 395
rect 22206 79 22242 420
rect 22278 0 22314 395
rect 22350 0 22386 395
rect 22542 0 22578 395
rect 22614 0 22650 395
rect 22686 79 22722 420
rect 22758 0 22794 395
rect 22830 0 22866 395
rect 23310 0 23346 395
rect 23382 0 23418 395
rect 23454 79 23490 420
rect 23526 0 23562 395
rect 23598 0 23634 395
rect 23790 0 23826 395
rect 23862 0 23898 395
rect 23934 79 23970 420
rect 24006 0 24042 395
rect 24078 0 24114 395
rect 24558 0 24594 395
rect 24630 0 24666 395
rect 24702 79 24738 420
rect 24774 0 24810 395
rect 24846 0 24882 395
rect 25038 0 25074 395
rect 25110 0 25146 395
rect 25182 79 25218 420
rect 25254 0 25290 395
rect 25326 0 25362 395
rect 25806 0 25842 395
rect 25878 0 25914 395
rect 25950 79 25986 420
rect 26022 0 26058 395
rect 26094 0 26130 395
rect 26286 0 26322 395
rect 26358 0 26394 395
rect 26430 79 26466 420
rect 26502 0 26538 395
rect 26574 0 26610 395
rect 27054 0 27090 395
rect 27126 0 27162 395
rect 27198 79 27234 420
rect 27270 0 27306 395
rect 27342 0 27378 395
rect 27534 0 27570 395
rect 27606 0 27642 395
rect 27678 79 27714 420
rect 27750 0 27786 395
rect 27822 0 27858 395
rect 28302 0 28338 395
rect 28374 0 28410 395
rect 28446 79 28482 420
rect 28518 0 28554 395
rect 28590 0 28626 395
rect 28782 0 28818 395
rect 28854 0 28890 395
rect 28926 79 28962 420
rect 28998 0 29034 395
rect 29070 0 29106 395
rect 29550 0 29586 395
rect 29622 0 29658 395
rect 29694 79 29730 420
rect 29766 0 29802 395
rect 29838 0 29874 395
rect 30030 0 30066 395
rect 30102 0 30138 395
rect 30174 79 30210 420
rect 30246 0 30282 395
rect 30318 0 30354 395
rect 30798 0 30834 395
rect 30870 0 30906 395
rect 30942 79 30978 420
rect 31014 0 31050 395
rect 31086 0 31122 395
rect 31278 0 31314 395
rect 31350 0 31386 395
rect 31422 79 31458 420
rect 31494 0 31530 395
rect 31566 0 31602 395
rect 32046 0 32082 395
rect 32118 0 32154 395
rect 32190 79 32226 420
rect 32262 0 32298 395
rect 32334 0 32370 395
rect 32526 0 32562 395
rect 32598 0 32634 395
rect 32670 79 32706 420
rect 32742 0 32778 395
rect 32814 0 32850 395
rect 33294 0 33330 395
rect 33366 0 33402 395
rect 33438 79 33474 420
rect 33510 0 33546 395
rect 33582 0 33618 395
rect 33774 0 33810 395
rect 33846 0 33882 395
rect 33918 79 33954 420
rect 33990 0 34026 395
rect 34062 0 34098 395
rect 34542 0 34578 395
rect 34614 0 34650 395
rect 34686 79 34722 420
rect 34758 0 34794 395
rect 34830 0 34866 395
rect 35022 0 35058 395
rect 35094 0 35130 395
rect 35166 79 35202 420
rect 35238 0 35274 395
rect 35310 0 35346 395
rect 35790 0 35826 395
rect 35862 0 35898 395
rect 35934 79 35970 420
rect 36006 0 36042 395
rect 36078 0 36114 395
rect 36270 0 36306 395
rect 36342 0 36378 395
rect 36414 79 36450 420
rect 36486 0 36522 395
rect 36558 0 36594 395
rect 37038 0 37074 395
rect 37110 0 37146 395
rect 37182 79 37218 420
rect 37254 0 37290 395
rect 37326 0 37362 395
rect 37518 0 37554 395
rect 37590 0 37626 395
rect 37662 79 37698 420
rect 37734 0 37770 395
rect 37806 0 37842 395
rect 38286 0 38322 395
rect 38358 0 38394 395
rect 38430 79 38466 420
rect 38502 0 38538 395
rect 38574 0 38610 395
rect 38766 0 38802 395
rect 38838 0 38874 395
rect 38910 79 38946 420
rect 38982 0 39018 395
rect 39054 0 39090 395
rect 39534 0 39570 395
rect 39606 0 39642 395
rect 39678 79 39714 420
rect 39750 0 39786 395
rect 39822 0 39858 395
<< metal2 >>
rect 0 323 39936 371
rect 186 199 294 275
rect 954 199 1062 275
rect 1434 199 1542 275
rect 2202 199 2310 275
rect 2682 199 2790 275
rect 3450 199 3558 275
rect 3930 199 4038 275
rect 4698 199 4806 275
rect 5178 199 5286 275
rect 5946 199 6054 275
rect 6426 199 6534 275
rect 7194 199 7302 275
rect 7674 199 7782 275
rect 8442 199 8550 275
rect 8922 199 9030 275
rect 9690 199 9798 275
rect 10170 199 10278 275
rect 10938 199 11046 275
rect 11418 199 11526 275
rect 12186 199 12294 275
rect 12666 199 12774 275
rect 13434 199 13542 275
rect 13914 199 14022 275
rect 14682 199 14790 275
rect 15162 199 15270 275
rect 15930 199 16038 275
rect 16410 199 16518 275
rect 17178 199 17286 275
rect 17658 199 17766 275
rect 18426 199 18534 275
rect 18906 199 19014 275
rect 19674 199 19782 275
rect 20154 199 20262 275
rect 20922 199 21030 275
rect 21402 199 21510 275
rect 22170 199 22278 275
rect 22650 199 22758 275
rect 23418 199 23526 275
rect 23898 199 24006 275
rect 24666 199 24774 275
rect 25146 199 25254 275
rect 25914 199 26022 275
rect 26394 199 26502 275
rect 27162 199 27270 275
rect 27642 199 27750 275
rect 28410 199 28518 275
rect 28890 199 28998 275
rect 29658 199 29766 275
rect 30138 199 30246 275
rect 30906 199 31014 275
rect 31386 199 31494 275
rect 32154 199 32262 275
rect 32634 199 32742 275
rect 33402 199 33510 275
rect 33882 199 33990 275
rect 34650 199 34758 275
rect 35130 199 35238 275
rect 35898 199 36006 275
rect 36378 199 36486 275
rect 37146 199 37254 275
rect 37626 199 37734 275
rect 38394 199 38502 275
rect 38874 199 38982 275
rect 39642 199 39750 275
rect 0 103 39936 151
rect 186 -55 294 55
rect 954 -55 1062 55
rect 1434 -55 1542 55
rect 2202 -55 2310 55
rect 2682 -55 2790 55
rect 3450 -55 3558 55
rect 3930 -55 4038 55
rect 4698 -55 4806 55
rect 5178 -55 5286 55
rect 5946 -55 6054 55
rect 6426 -55 6534 55
rect 7194 -55 7302 55
rect 7674 -55 7782 55
rect 8442 -55 8550 55
rect 8922 -55 9030 55
rect 9690 -55 9798 55
rect 10170 -55 10278 55
rect 10938 -55 11046 55
rect 11418 -55 11526 55
rect 12186 -55 12294 55
rect 12666 -55 12774 55
rect 13434 -55 13542 55
rect 13914 -55 14022 55
rect 14682 -55 14790 55
rect 15162 -55 15270 55
rect 15930 -55 16038 55
rect 16410 -55 16518 55
rect 17178 -55 17286 55
rect 17658 -55 17766 55
rect 18426 -55 18534 55
rect 18906 -55 19014 55
rect 19674 -55 19782 55
rect 20154 -55 20262 55
rect 20922 -55 21030 55
rect 21402 -55 21510 55
rect 22170 -55 22278 55
rect 22650 -55 22758 55
rect 23418 -55 23526 55
rect 23898 -55 24006 55
rect 24666 -55 24774 55
rect 25146 -55 25254 55
rect 25914 -55 26022 55
rect 26394 -55 26502 55
rect 27162 -55 27270 55
rect 27642 -55 27750 55
rect 28410 -55 28518 55
rect 28890 -55 28998 55
rect 29658 -55 29766 55
rect 30138 -55 30246 55
rect 30906 -55 31014 55
rect 31386 -55 31494 55
rect 32154 -55 32262 55
rect 32634 -55 32742 55
rect 33402 -55 33510 55
rect 33882 -55 33990 55
rect 34650 -55 34758 55
rect 35130 -55 35238 55
rect 35898 -55 36006 55
rect 36378 -55 36486 55
rect 37146 -55 37254 55
rect 37626 -55 37734 55
rect 38394 -55 38502 55
rect 38874 -55 38982 55
rect 39642 -55 39750 55
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_0
timestamp 1704896540
transform -1 0 39936 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_1
timestamp 1704896540
transform 1 0 38688 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_2
timestamp 1704896540
transform -1 0 38688 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_3
timestamp 1704896540
transform 1 0 37440 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_4
timestamp 1704896540
transform -1 0 37440 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_5
timestamp 1704896540
transform 1 0 36192 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_6
timestamp 1704896540
transform -1 0 36192 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_7
timestamp 1704896540
transform 1 0 34944 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_8
timestamp 1704896540
transform -1 0 34944 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_9
timestamp 1704896540
transform 1 0 33696 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_10
timestamp 1704896540
transform -1 0 33696 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_11
timestamp 1704896540
transform 1 0 32448 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_12
timestamp 1704896540
transform -1 0 32448 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_13
timestamp 1704896540
transform 1 0 31200 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_14
timestamp 1704896540
transform -1 0 31200 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_15
timestamp 1704896540
transform 1 0 29952 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_16
timestamp 1704896540
transform -1 0 29952 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_17
timestamp 1704896540
transform 1 0 28704 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_18
timestamp 1704896540
transform -1 0 28704 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_19
timestamp 1704896540
transform 1 0 27456 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_20
timestamp 1704896540
transform -1 0 27456 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_21
timestamp 1704896540
transform 1 0 26208 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_22
timestamp 1704896540
transform -1 0 26208 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_23
timestamp 1704896540
transform 1 0 24960 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_24
timestamp 1704896540
transform -1 0 24960 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_25
timestamp 1704896540
transform 1 0 23712 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_26
timestamp 1704896540
transform -1 0 23712 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_27
timestamp 1704896540
transform 1 0 22464 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_28
timestamp 1704896540
transform -1 0 22464 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_29
timestamp 1704896540
transform 1 0 21216 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_30
timestamp 1704896540
transform -1 0 21216 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_31
timestamp 1704896540
transform 1 0 19968 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_32
timestamp 1704896540
transform -1 0 19968 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_33
timestamp 1704896540
transform 1 0 18720 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_34
timestamp 1704896540
transform -1 0 18720 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_35
timestamp 1704896540
transform 1 0 17472 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_36
timestamp 1704896540
transform -1 0 17472 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_37
timestamp 1704896540
transform 1 0 16224 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_38
timestamp 1704896540
transform -1 0 16224 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_39
timestamp 1704896540
transform 1 0 14976 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_40
timestamp 1704896540
transform -1 0 14976 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_41
timestamp 1704896540
transform 1 0 13728 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_42
timestamp 1704896540
transform -1 0 13728 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_43
timestamp 1704896540
transform 1 0 12480 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_44
timestamp 1704896540
transform -1 0 12480 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_45
timestamp 1704896540
transform 1 0 11232 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_46
timestamp 1704896540
transform -1 0 11232 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_47
timestamp 1704896540
transform 1 0 9984 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_48
timestamp 1704896540
transform -1 0 9984 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_49
timestamp 1704896540
transform 1 0 8736 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_50
timestamp 1704896540
transform -1 0 8736 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_51
timestamp 1704896540
transform 1 0 7488 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_52
timestamp 1704896540
transform -1 0 7488 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_53
timestamp 1704896540
transform 1 0 6240 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_54
timestamp 1704896540
transform -1 0 6240 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_55
timestamp 1704896540
transform 1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_56
timestamp 1704896540
transform -1 0 4992 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_57
timestamp 1704896540
transform 1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_58
timestamp 1704896540
transform -1 0 3744 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_59
timestamp 1704896540
transform 1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_60
timestamp 1704896540
transform -1 0 2496 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_61
timestamp 1704896540
transform 1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_62
timestamp 1704896540
transform -1 0 1248 0 1 0
box -42 -105 650 421
use sky130_fd_bd_sram__openram_dp_cell_dummy_2  sky130_fd_bd_sram__openram_dp_cell_dummy_63
timestamp 1704896540
transform 1 0 0 0 1 0
box -42 -105 650 421
<< labels >>
rlabel metal1 s 34704 249 34704 249 4 vdd
port 1 nsew
rlabel metal1 s 36432 249 36432 249 4 vdd
port 1 nsew
rlabel metal1 s 35952 249 35952 249 4 vdd
port 1 nsew
rlabel metal1 s 30960 249 30960 249 4 vdd
port 1 nsew
rlabel metal1 s 37680 249 37680 249 4 vdd
port 1 nsew
rlabel metal1 s 38928 249 38928 249 4 vdd
port 1 nsew
rlabel metal1 s 22224 249 22224 249 4 vdd
port 1 nsew
rlabel metal1 s 33936 249 33936 249 4 vdd
port 1 nsew
rlabel metal1 s 25200 249 25200 249 4 vdd
port 1 nsew
rlabel metal1 s 28464 249 28464 249 4 vdd
port 1 nsew
rlabel metal1 s 37200 249 37200 249 4 vdd
port 1 nsew
rlabel metal1 s 30192 249 30192 249 4 vdd
port 1 nsew
rlabel metal1 s 31440 249 31440 249 4 vdd
port 1 nsew
rlabel metal1 s 32688 249 32688 249 4 vdd
port 1 nsew
rlabel metal1 s 39696 249 39696 249 4 vdd
port 1 nsew
rlabel metal1 s 22704 249 22704 249 4 vdd
port 1 nsew
rlabel metal1 s 23472 249 23472 249 4 vdd
port 1 nsew
rlabel metal1 s 25968 249 25968 249 4 vdd
port 1 nsew
rlabel metal1 s 27696 249 27696 249 4 vdd
port 1 nsew
rlabel metal1 s 38448 249 38448 249 4 vdd
port 1 nsew
rlabel metal1 s 29712 249 29712 249 4 vdd
port 1 nsew
rlabel metal1 s 27216 249 27216 249 4 vdd
port 1 nsew
rlabel metal1 s 26448 249 26448 249 4 vdd
port 1 nsew
rlabel metal1 s 24720 249 24720 249 4 vdd
port 1 nsew
rlabel metal1 s 35184 249 35184 249 4 vdd
port 1 nsew
rlabel metal1 s 20976 249 20976 249 4 vdd
port 1 nsew
rlabel metal1 s 23952 249 23952 249 4 vdd
port 1 nsew
rlabel metal1 s 21456 249 21456 249 4 vdd
port 1 nsew
rlabel metal1 s 20208 249 20208 249 4 vdd
port 1 nsew
rlabel metal1 s 32208 249 32208 249 4 vdd
port 1 nsew
rlabel metal1 s 28944 249 28944 249 4 vdd
port 1 nsew
rlabel metal1 s 33456 249 33456 249 4 vdd
port 1 nsew
rlabel metal1 s 7728 249 7728 249 4 vdd
port 1 nsew
rlabel metal1 s 18480 249 18480 249 4 vdd
port 1 nsew
rlabel metal1 s 3504 249 3504 249 4 vdd
port 1 nsew
rlabel metal1 s 3984 249 3984 249 4 vdd
port 1 nsew
rlabel metal1 s 13968 249 13968 249 4 vdd
port 1 nsew
rlabel metal1 s 1488 249 1488 249 4 vdd
port 1 nsew
rlabel metal1 s 2256 249 2256 249 4 vdd
port 1 nsew
rlabel metal1 s 15216 249 15216 249 4 vdd
port 1 nsew
rlabel metal1 s 14736 249 14736 249 4 vdd
port 1 nsew
rlabel metal1 s 10992 249 10992 249 4 vdd
port 1 nsew
rlabel metal1 s 2736 249 2736 249 4 vdd
port 1 nsew
rlabel metal1 s 17232 249 17232 249 4 vdd
port 1 nsew
rlabel metal1 s 13488 249 13488 249 4 vdd
port 1 nsew
rlabel metal1 s 11472 249 11472 249 4 vdd
port 1 nsew
rlabel metal1 s 240 249 240 249 4 vdd
port 1 nsew
rlabel metal1 s 8496 249 8496 249 4 vdd
port 1 nsew
rlabel metal1 s 4752 249 4752 249 4 vdd
port 1 nsew
rlabel metal1 s 18960 249 18960 249 4 vdd
port 1 nsew
rlabel metal1 s 16464 249 16464 249 4 vdd
port 1 nsew
rlabel metal1 s 1008 249 1008 249 4 vdd
port 1 nsew
rlabel metal1 s 5232 249 5232 249 4 vdd
port 1 nsew
rlabel metal1 s 12720 249 12720 249 4 vdd
port 1 nsew
rlabel metal1 s 6000 249 6000 249 4 vdd
port 1 nsew
rlabel metal1 s 17712 249 17712 249 4 vdd
port 1 nsew
rlabel metal1 s 6480 249 6480 249 4 vdd
port 1 nsew
rlabel metal1 s 7248 249 7248 249 4 vdd
port 1 nsew
rlabel metal1 s 12240 249 12240 249 4 vdd
port 1 nsew
rlabel metal1 s 9744 249 9744 249 4 vdd
port 1 nsew
rlabel metal1 s 8976 249 8976 249 4 vdd
port 1 nsew
rlabel metal1 s 19728 249 19728 249 4 vdd
port 1 nsew
rlabel metal1 s 10224 249 10224 249 4 vdd
port 1 nsew
rlabel metal1 s 15984 249 15984 249 4 vdd
port 1 nsew
rlabel metal1 s 7104 197 7104 197 4 br1_11
port 308 nsew
rlabel metal1 s 8424 197 8424 197 4 bl1_13
port 315 nsew
rlabel metal1 s 2112 197 2112 197 4 br1_3
port 276 nsew
rlabel metal1 s 5928 197 5928 197 4 bl1_9
port 299 nsew
rlabel metal1 s 168 197 168 197 4 br0_0
port 262 nsew
rlabel metal1 s 4056 197 4056 197 4 bl1_6
port 287 nsew
rlabel metal1 s 2664 197 2664 197 4 br0_4
port 278 nsew
rlabel metal1 s 8568 197 8568 197 4 br0_13
port 314 nsew
rlabel metal1 s 2328 197 2328 197 4 br0_3
port 274 nsew
rlabel metal1 s 3576 197 3576 197 4 br0_5
port 282 nsew
rlabel metal1 s 6072 197 6072 197 4 br0_9
port 298 nsew
rlabel metal1 s 4128 197 4128 197 4 br1_6
port 288 nsew
rlabel metal1 s 1080 197 1080 197 4 br0_1
port 266 nsew
rlabel metal1 s 3360 197 3360 197 4 br1_5
port 284 nsew
rlabel metal1 s 5376 197 5376 197 4 br1_8
port 296 nsew
rlabel metal1 s 2184 197 2184 197 4 bl1_3
port 275 nsew
rlabel metal1 s 9600 197 9600 197 4 br1_15
port 324 nsew
rlabel metal1 s 2808 197 2808 197 4 bl1_4
port 279 nsew
rlabel metal1 s 3912 197 3912 197 4 br0_6
port 286 nsew
rlabel metal1 s 864 197 864 197 4 br1_1
port 268 nsew
rlabel metal1 s 312 197 312 197 4 bl1_0
port 263 nsew
rlabel metal1 s 5304 197 5304 197 4 bl1_8
port 295 nsew
rlabel metal1 s 8352 197 8352 197 4 br1_13
port 316 nsew
rlabel metal1 s 2880 197 2880 197 4 br1_4
port 280 nsew
rlabel metal1 s 1560 197 1560 197 4 bl1_2
port 271 nsew
rlabel metal1 s 9816 197 9816 197 4 br0_15
port 322 nsew
rlabel metal1 s 7584 197 7584 197 4 bl0_12
port 309 nsew
rlabel metal1 s 4680 197 4680 197 4 bl1_7
port 291 nsew
rlabel metal1 s 8640 197 8640 197 4 bl0_13
port 313 nsew
rlabel metal1 s 4824 197 4824 197 4 br0_7
port 290 nsew
rlabel metal1 s 7392 197 7392 197 4 bl0_11
port 305 nsew
rlabel metal1 s 6408 197 6408 197 4 br0_10
port 302 nsew
rlabel metal1 s 7800 197 7800 197 4 bl1_12
port 311 nsew
rlabel metal1 s 5856 197 5856 197 4 br1_9
port 300 nsew
rlabel metal1 s 2592 197 2592 197 4 bl0_4
port 277 nsew
rlabel metal1 s 8904 197 8904 197 4 br0_14
port 318 nsew
rlabel metal1 s 6624 197 6624 197 4 br1_10
port 304 nsew
rlabel metal1 s 384 197 384 197 4 br1_0
port 264 nsew
rlabel metal1 s 3432 197 3432 197 4 bl1_5
port 283 nsew
rlabel metal1 s 7656 197 7656 197 4 br0_12
port 310 nsew
rlabel metal1 s 6552 197 6552 197 4 bl1_10
port 303 nsew
rlabel metal1 s 6336 197 6336 197 4 bl0_10
port 301 nsew
rlabel metal1 s 9672 197 9672 197 4 bl1_15
port 323 nsew
rlabel metal1 s 6144 197 6144 197 4 bl0_9
port 297 nsew
rlabel metal1 s 1632 197 1632 197 4 br1_2
port 272 nsew
rlabel metal1 s 9888 197 9888 197 4 bl0_15
port 321 nsew
rlabel metal1 s 1344 197 1344 197 4 bl0_2
port 269 nsew
rlabel metal1 s 7320 197 7320 197 4 br0_11
port 306 nsew
rlabel metal1 s 5160 197 5160 197 4 br0_8
port 294 nsew
rlabel metal1 s 2400 197 2400 197 4 bl0_3
port 273 nsew
rlabel metal1 s 1416 197 1416 197 4 br0_2
port 270 nsew
rlabel metal1 s 8832 197 8832 197 4 bl0_14
port 317 nsew
rlabel metal1 s 1152 197 1152 197 4 bl0_1
port 265 nsew
rlabel metal1 s 7872 197 7872 197 4 br1_12
port 312 nsew
rlabel metal1 s 5088 197 5088 197 4 bl0_8
port 293 nsew
rlabel metal1 s 7176 197 7176 197 4 bl1_11
port 307 nsew
rlabel metal1 s 96 197 96 197 4 bl0_0
port 261 nsew
rlabel metal1 s 936 197 936 197 4 bl1_1
port 267 nsew
rlabel metal1 s 9048 197 9048 197 4 bl1_14
port 319 nsew
rlabel metal1 s 4608 197 4608 197 4 br1_7
port 292 nsew
rlabel metal1 s 9120 197 9120 197 4 br1_14
port 320 nsew
rlabel metal1 s 4896 197 4896 197 4 bl0_7
port 289 nsew
rlabel metal1 s 3648 197 3648 197 4 bl0_5
port 281 nsew
rlabel metal1 s 3840 197 3840 197 4 bl0_6
port 285 nsew
rlabel metal1 s 17160 197 17160 197 4 bl1_27
port 371 nsew
rlabel metal1 s 18624 197 18624 197 4 bl0_29
port 377 nsew
rlabel metal1 s 14112 197 14112 197 4 br1_22
port 352 nsew
rlabel metal1 s 19872 197 19872 197 4 bl0_31
port 385 nsew
rlabel metal1 s 10920 197 10920 197 4 bl1_17
port 331 nsew
rlabel metal1 s 15288 197 15288 197 4 bl1_24
port 359 nsew
rlabel metal1 s 11544 197 11544 197 4 bl1_18
port 335 nsew
rlabel metal1 s 19104 197 19104 197 4 br1_30
port 384 nsew
rlabel metal1 s 18552 197 18552 197 4 br0_29
port 378 nsew
rlabel metal1 s 19656 197 19656 197 4 bl1_31
port 387 nsew
rlabel metal1 s 16320 197 16320 197 4 bl0_26
port 365 nsew
rlabel metal1 s 16128 197 16128 197 4 bl0_25
port 361 nsew
rlabel metal1 s 14880 197 14880 197 4 bl0_23
port 353 nsew
rlabel metal1 s 13824 197 13824 197 4 bl0_22
port 349 nsew
rlabel metal1 s 12576 197 12576 197 4 bl0_20
port 341 nsew
rlabel metal1 s 14592 197 14592 197 4 br1_23
port 356 nsew
rlabel metal1 s 15840 197 15840 197 4 br1_25
port 364 nsew
rlabel metal1 s 12792 197 12792 197 4 bl1_20
port 343 nsew
rlabel metal1 s 10296 197 10296 197 4 bl1_16
port 327 nsew
rlabel metal1 s 15144 197 15144 197 4 br0_24
port 358 nsew
rlabel metal1 s 12312 197 12312 197 4 br0_19
port 338 nsew
rlabel metal1 s 13632 197 13632 197 4 bl0_21
port 345 nsew
rlabel metal1 s 17376 197 17376 197 4 bl0_27
port 369 nsew
rlabel metal1 s 11616 197 11616 197 4 br1_18
port 336 nsew
rlabel metal1 s 11400 197 11400 197 4 br0_18
port 334 nsew
rlabel metal1 s 11064 197 11064 197 4 br0_17
port 330 nsew
rlabel metal1 s 17304 197 17304 197 4 br0_27
port 370 nsew
rlabel metal1 s 17784 197 17784 197 4 bl1_28
port 375 nsew
rlabel metal1 s 19800 197 19800 197 4 br0_31
port 386 nsew
rlabel metal1 s 18888 197 18888 197 4 br0_30
port 382 nsew
rlabel metal1 s 10080 197 10080 197 4 bl0_16
port 325 nsew
rlabel metal1 s 10152 197 10152 197 4 br0_16
port 326 nsew
rlabel metal1 s 19584 197 19584 197 4 br1_31
port 388 nsew
rlabel metal1 s 13344 197 13344 197 4 br1_21
port 348 nsew
rlabel metal1 s 15072 197 15072 197 4 bl0_24
port 357 nsew
rlabel metal1 s 10848 197 10848 197 4 br1_17
port 332 nsew
rlabel metal1 s 13560 197 13560 197 4 br0_21
port 346 nsew
rlabel metal1 s 16392 197 16392 197 4 br0_26
port 366 nsew
rlabel metal1 s 12384 197 12384 197 4 bl0_19
port 337 nsew
rlabel metal1 s 12168 197 12168 197 4 bl1_19
port 339 nsew
rlabel metal1 s 11136 197 11136 197 4 bl0_17
port 329 nsew
rlabel metal1 s 13896 197 13896 197 4 br0_22
port 350 nsew
rlabel metal1 s 18336 197 18336 197 4 br1_29
port 380 nsew
rlabel metal1 s 18816 197 18816 197 4 bl0_30
port 381 nsew
rlabel metal1 s 19032 197 19032 197 4 bl1_30
port 383 nsew
rlabel metal1 s 15912 197 15912 197 4 bl1_25
port 363 nsew
rlabel metal1 s 12096 197 12096 197 4 br1_19
port 340 nsew
rlabel metal1 s 11328 197 11328 197 4 bl0_18
port 333 nsew
rlabel metal1 s 17088 197 17088 197 4 br1_27
port 372 nsew
rlabel metal1 s 15360 197 15360 197 4 br1_24
port 360 nsew
rlabel metal1 s 16536 197 16536 197 4 bl1_26
port 367 nsew
rlabel metal1 s 14040 197 14040 197 4 bl1_22
port 351 nsew
rlabel metal1 s 17640 197 17640 197 4 br0_28
port 374 nsew
rlabel metal1 s 13416 197 13416 197 4 bl1_21
port 347 nsew
rlabel metal1 s 12648 197 12648 197 4 br0_20
port 342 nsew
rlabel metal1 s 14808 197 14808 197 4 br0_23
port 354 nsew
rlabel metal1 s 17856 197 17856 197 4 br1_28
port 376 nsew
rlabel metal1 s 14664 197 14664 197 4 bl1_23
port 355 nsew
rlabel metal1 s 18408 197 18408 197 4 bl1_29
port 379 nsew
rlabel metal1 s 12864 197 12864 197 4 br1_20
port 344 nsew
rlabel metal1 s 16608 197 16608 197 4 br1_26
port 368 nsew
rlabel metal1 s 10368 197 10368 197 4 br1_16
port 328 nsew
rlabel metal1 s 16056 197 16056 197 4 br0_25
port 362 nsew
rlabel metal1 s 17568 197 17568 197 4 bl0_28
port 373 nsew
rlabel metal1 s 25056 197 25056 197 4 bl0_40
port 421 nsew
rlabel metal1 s 28608 197 28608 197 4 bl0_45
port 441 nsew
rlabel metal1 s 29784 197 29784 197 4 br0_47
port 450 nsew
rlabel metal1 s 27144 197 27144 197 4 bl1_43
port 435 nsew
rlabel metal1 s 22152 197 22152 197 4 bl1_35
port 403 nsew
rlabel metal1 s 20904 197 20904 197 4 bl1_33
port 395 nsew
rlabel metal1 s 25272 197 25272 197 4 bl1_40
port 423 nsew
rlabel metal1 s 20136 197 20136 197 4 br0_32
port 390 nsew
rlabel metal1 s 23616 197 23616 197 4 bl0_37
port 409 nsew
rlabel metal1 s 27840 197 27840 197 4 br1_44
port 440 nsew
rlabel metal1 s 27360 197 27360 197 4 bl0_43
port 433 nsew
rlabel metal1 s 25128 197 25128 197 4 br0_40
port 422 nsew
rlabel metal1 s 22632 197 22632 197 4 br0_36
port 406 nsew
rlabel metal1 s 22080 197 22080 197 4 br1_35
port 404 nsew
rlabel metal1 s 20832 197 20832 197 4 br1_33
port 396 nsew
rlabel metal1 s 25344 197 25344 197 4 br1_40
port 424 nsew
rlabel metal1 s 28536 197 28536 197 4 br0_45
port 442 nsew
rlabel metal1 s 22296 197 22296 197 4 br0_35
port 402 nsew
rlabel metal1 s 21600 197 21600 197 4 br1_34
port 400 nsew
rlabel metal1 s 29856 197 29856 197 4 bl0_47
port 449 nsew
rlabel metal1 s 28320 197 28320 197 4 br1_45
port 444 nsew
rlabel metal1 s 25824 197 25824 197 4 br1_41
port 428 nsew
rlabel metal1 s 26040 197 26040 197 4 br0_41
port 426 nsew
rlabel metal1 s 27288 197 27288 197 4 br0_43
port 434 nsew
rlabel metal1 s 23400 197 23400 197 4 bl1_37
port 411 nsew
rlabel metal1 s 23328 197 23328 197 4 br1_37
port 412 nsew
rlabel metal1 s 28392 197 28392 197 4 bl1_45
port 443 nsew
rlabel metal1 s 24576 197 24576 197 4 br1_39
port 420 nsew
rlabel metal1 s 27768 197 27768 197 4 bl1_44
port 439 nsew
rlabel metal1 s 26520 197 26520 197 4 bl1_42
port 431 nsew
rlabel metal1 s 26592 197 26592 197 4 br1_42
port 432 nsew
rlabel metal1 s 26304 197 26304 197 4 bl0_42
port 429 nsew
rlabel metal1 s 28872 197 28872 197 4 br0_46
port 446 nsew
rlabel metal1 s 23880 197 23880 197 4 br0_38
port 414 nsew
rlabel metal1 s 29640 197 29640 197 4 bl1_47
port 451 nsew
rlabel metal1 s 26376 197 26376 197 4 br0_42
port 430 nsew
rlabel metal1 s 24792 197 24792 197 4 br0_39
port 418 nsew
rlabel metal1 s 24024 197 24024 197 4 bl1_38
port 415 nsew
rlabel metal1 s 22848 197 22848 197 4 br1_36
port 408 nsew
rlabel metal1 s 26112 197 26112 197 4 bl0_41
port 425 nsew
rlabel metal1 s 29568 197 29568 197 4 br1_47
port 452 nsew
rlabel metal1 s 27072 197 27072 197 4 br1_43
port 436 nsew
rlabel metal1 s 29016 197 29016 197 4 bl1_46
port 447 nsew
rlabel metal1 s 27552 197 27552 197 4 bl0_44
port 437 nsew
rlabel metal1 s 21528 197 21528 197 4 bl1_34
port 399 nsew
rlabel metal1 s 24864 197 24864 197 4 bl0_39
port 417 nsew
rlabel metal1 s 23808 197 23808 197 4 bl0_38
port 413 nsew
rlabel metal1 s 24096 197 24096 197 4 br1_38
port 416 nsew
rlabel metal1 s 29088 197 29088 197 4 br1_46
port 448 nsew
rlabel metal1 s 28800 197 28800 197 4 bl0_46
port 445 nsew
rlabel metal1 s 23544 197 23544 197 4 br0_37
port 410 nsew
rlabel metal1 s 27624 197 27624 197 4 br0_44
port 438 nsew
rlabel metal1 s 21312 197 21312 197 4 bl0_34
port 397 nsew
rlabel metal1 s 24648 197 24648 197 4 bl1_39
port 419 nsew
rlabel metal1 s 20064 197 20064 197 4 bl0_32
port 389 nsew
rlabel metal1 s 22368 197 22368 197 4 bl0_35
port 401 nsew
rlabel metal1 s 21048 197 21048 197 4 br0_33
port 394 nsew
rlabel metal1 s 21120 197 21120 197 4 bl0_33
port 393 nsew
rlabel metal1 s 20280 197 20280 197 4 bl1_32
port 391 nsew
rlabel metal1 s 21384 197 21384 197 4 br0_34
port 398 nsew
rlabel metal1 s 22560 197 22560 197 4 bl0_36
port 405 nsew
rlabel metal1 s 20352 197 20352 197 4 br1_32
port 392 nsew
rlabel metal1 s 22776 197 22776 197 4 bl1_36
port 407 nsew
rlabel metal1 s 25896 197 25896 197 4 bl1_41
port 427 nsew
rlabel metal1 s 32544 197 32544 197 4 bl0_52
port 469 nsew
rlabel metal1 s 30048 197 30048 197 4 bl0_48
port 453 nsew
rlabel metal1 s 33600 197 33600 197 4 bl0_53
port 473 nsew
rlabel metal1 s 34080 197 34080 197 4 br1_54
port 480 nsew
rlabel metal1 s 37128 197 37128 197 4 bl1_59
port 499 nsew
rlabel metal1 s 36360 197 36360 197 4 br0_58
port 494 nsew
rlabel metal1 s 31104 197 31104 197 4 bl0_49
port 457 nsew
rlabel metal1 s 38376 197 38376 197 4 bl1_61
port 507 nsew
rlabel metal1 s 30264 197 30264 197 4 bl1_48
port 455 nsew
rlabel metal1 s 32280 197 32280 197 4 br0_51
port 466 nsew
rlabel metal1 s 37824 197 37824 197 4 br1_60
port 504 nsew
rlabel metal1 s 34776 197 34776 197 4 br0_55
port 482 nsew
rlabel metal1 s 39072 197 39072 197 4 br1_62
port 512 nsew
rlabel metal1 s 38520 197 38520 197 4 br0_61
port 506 nsew
rlabel metal1 s 35328 197 35328 197 4 br1_56
port 488 nsew
rlabel metal1 s 38856 197 38856 197 4 br0_62
port 510 nsew
rlabel metal1 s 32760 197 32760 197 4 bl1_52
port 471 nsew
rlabel metal1 s 35040 197 35040 197 4 bl0_56
port 485 nsew
rlabel metal1 s 38592 197 38592 197 4 bl0_61
port 505 nsew
rlabel metal1 s 31368 197 31368 197 4 br0_50
port 462 nsew
rlabel metal1 s 38304 197 38304 197 4 br1_61
port 508 nsew
rlabel metal1 s 35112 197 35112 197 4 br0_56
port 486 nsew
rlabel metal1 s 33384 197 33384 197 4 bl1_53
port 475 nsew
rlabel metal1 s 35808 197 35808 197 4 br1_57
port 492 nsew
rlabel metal1 s 36504 197 36504 197 4 bl1_58
port 495 nsew
rlabel metal1 s 30816 197 30816 197 4 br1_49
port 460 nsew
rlabel metal1 s 32832 197 32832 197 4 br1_52
port 472 nsew
rlabel metal1 s 32352 197 32352 197 4 bl0_51
port 465 nsew
rlabel metal1 s 36576 197 36576 197 4 br1_58
port 496 nsew
rlabel metal1 s 36288 197 36288 197 4 bl0_58
port 493 nsew
rlabel metal1 s 32136 197 32136 197 4 bl1_51
port 467 nsew
rlabel metal1 s 34632 197 34632 197 4 bl1_55
port 483 nsew
rlabel metal1 s 30888 197 30888 197 4 bl1_49
port 459 nsew
rlabel metal1 s 37344 197 37344 197 4 bl0_59
port 497 nsew
rlabel metal1 s 31512 197 31512 197 4 bl1_50
port 463 nsew
rlabel metal1 s 34848 197 34848 197 4 bl0_55
port 481 nsew
rlabel metal1 s 33528 197 33528 197 4 br0_53
port 474 nsew
rlabel metal1 s 36096 197 36096 197 4 bl0_57
port 489 nsew
rlabel metal1 s 33864 197 33864 197 4 br0_54
port 478 nsew
rlabel metal1 s 33792 197 33792 197 4 bl0_54
port 477 nsew
rlabel metal1 s 37536 197 37536 197 4 bl0_60
port 501 nsew
rlabel metal1 s 37752 197 37752 197 4 bl1_60
port 503 nsew
rlabel metal1 s 37056 197 37056 197 4 br1_59
port 500 nsew
rlabel metal1 s 33312 197 33312 197 4 br1_53
port 476 nsew
rlabel metal1 s 32616 197 32616 197 4 br0_52
port 470 nsew
rlabel metal1 s 37608 197 37608 197 4 br0_60
port 502 nsew
rlabel metal1 s 34008 197 34008 197 4 bl1_54
port 479 nsew
rlabel metal1 s 39768 197 39768 197 4 br0_63
port 514 nsew
rlabel metal1 s 39840 197 39840 197 4 bl0_63
port 513 nsew
rlabel metal1 s 38784 197 38784 197 4 bl0_62
port 509 nsew
rlabel metal1 s 39552 197 39552 197 4 br1_63
port 516 nsew
rlabel metal1 s 39000 197 39000 197 4 bl1_62
port 511 nsew
rlabel metal1 s 37272 197 37272 197 4 br0_59
port 498 nsew
rlabel metal1 s 35256 197 35256 197 4 bl1_56
port 487 nsew
rlabel metal1 s 30120 197 30120 197 4 br0_48
port 454 nsew
rlabel metal1 s 39624 197 39624 197 4 bl1_63
port 515 nsew
rlabel metal1 s 31584 197 31584 197 4 br1_50
port 464 nsew
rlabel metal1 s 34560 197 34560 197 4 br1_55
port 484 nsew
rlabel metal1 s 30336 197 30336 197 4 br1_48
port 456 nsew
rlabel metal1 s 36024 197 36024 197 4 br0_57
port 490 nsew
rlabel metal1 s 31296 197 31296 197 4 bl0_50
port 461 nsew
rlabel metal1 s 31032 197 31032 197 4 br0_49
port 458 nsew
rlabel metal1 s 35880 197 35880 197 4 bl1_57
port 491 nsew
rlabel metal1 s 32064 197 32064 197 4 br1_51
port 468 nsew
rlabel metal2 s 27216 237 27216 237 4 gnd
port 2 nsew
rlabel metal2 s 29712 237 29712 237 4 gnd
port 2 nsew
rlabel metal2 s 20976 237 20976 237 4 gnd
port 2 nsew
rlabel metal2 s 25200 237 25200 237 4 gnd
port 2 nsew
rlabel metal2 s 28464 237 28464 237 4 gnd
port 2 nsew
rlabel metal2 s 39696 237 39696 237 4 gnd
port 2 nsew
rlabel metal2 s 27696 237 27696 237 4 gnd
port 2 nsew
rlabel metal2 s 24720 237 24720 237 4 gnd
port 2 nsew
rlabel metal2 s 22224 237 22224 237 4 gnd
port 2 nsew
rlabel metal2 s 30192 237 30192 237 4 gnd
port 2 nsew
rlabel metal2 s 35184 237 35184 237 4 gnd
port 2 nsew
rlabel metal2 s 22704 237 22704 237 4 gnd
port 2 nsew
rlabel metal2 s 32688 237 32688 237 4 gnd
port 2 nsew
rlabel metal2 s 33936 237 33936 237 4 gnd
port 2 nsew
rlabel metal2 s 25968 237 25968 237 4 gnd
port 2 nsew
rlabel metal2 s 36432 237 36432 237 4 gnd
port 2 nsew
rlabel metal2 s 23472 237 23472 237 4 gnd
port 2 nsew
rlabel metal2 s 37680 237 37680 237 4 gnd
port 2 nsew
rlabel metal2 s 38448 237 38448 237 4 gnd
port 2 nsew
rlabel metal2 s 34704 237 34704 237 4 gnd
port 2 nsew
rlabel metal2 s 30960 237 30960 237 4 gnd
port 2 nsew
rlabel metal2 s 20208 237 20208 237 4 gnd
port 2 nsew
rlabel metal2 s 23952 237 23952 237 4 gnd
port 2 nsew
rlabel metal2 s 32208 237 32208 237 4 gnd
port 2 nsew
rlabel metal2 s 33456 237 33456 237 4 gnd
port 2 nsew
rlabel metal2 s 37200 237 37200 237 4 gnd
port 2 nsew
rlabel metal2 s 38928 237 38928 237 4 gnd
port 2 nsew
rlabel metal2 s 28944 237 28944 237 4 gnd
port 2 nsew
rlabel metal2 s 35952 237 35952 237 4 gnd
port 2 nsew
rlabel metal2 s 26448 237 26448 237 4 gnd
port 2 nsew
rlabel metal2 s 31440 237 31440 237 4 gnd
port 2 nsew
rlabel metal2 s 21456 237 21456 237 4 gnd
port 2 nsew
rlabel metal2 s 18480 237 18480 237 4 gnd
port 2 nsew
rlabel metal2 s 9744 237 9744 237 4 gnd
port 2 nsew
rlabel metal2 s 17232 237 17232 237 4 gnd
port 2 nsew
rlabel metal2 s 18960 237 18960 237 4 gnd
port 2 nsew
rlabel metal2 s 12720 237 12720 237 4 gnd
port 2 nsew
rlabel metal2 s 6480 237 6480 237 4 gnd
port 2 nsew
rlabel metal2 s 10224 237 10224 237 4 gnd
port 2 nsew
rlabel metal2 s 15984 237 15984 237 4 gnd
port 2 nsew
rlabel metal2 s 16464 237 16464 237 4 gnd
port 2 nsew
rlabel metal2 s 3504 237 3504 237 4 gnd
port 2 nsew
rlabel metal2 s 13488 237 13488 237 4 gnd
port 2 nsew
rlabel metal2 s 19728 237 19728 237 4 gnd
port 2 nsew
rlabel metal2 s 8976 237 8976 237 4 gnd
port 2 nsew
rlabel metal2 s 14736 237 14736 237 4 gnd
port 2 nsew
rlabel metal2 s 7248 237 7248 237 4 gnd
port 2 nsew
rlabel metal2 s 10992 237 10992 237 4 gnd
port 2 nsew
rlabel metal2 s 5232 237 5232 237 4 gnd
port 2 nsew
rlabel metal2 s 11472 237 11472 237 4 gnd
port 2 nsew
rlabel metal2 s 1008 237 1008 237 4 gnd
port 2 nsew
rlabel metal2 s 17712 237 17712 237 4 gnd
port 2 nsew
rlabel metal2 s 1488 237 1488 237 4 gnd
port 2 nsew
rlabel metal2 s 12240 237 12240 237 4 gnd
port 2 nsew
rlabel metal2 s 3984 237 3984 237 4 gnd
port 2 nsew
rlabel metal2 s 240 237 240 237 4 gnd
port 2 nsew
rlabel metal2 s 8496 237 8496 237 4 gnd
port 2 nsew
rlabel metal2 s 2736 237 2736 237 4 gnd
port 2 nsew
rlabel metal2 s 4752 237 4752 237 4 gnd
port 2 nsew
rlabel metal2 s 2256 237 2256 237 4 gnd
port 2 nsew
rlabel metal2 s 7728 237 7728 237 4 gnd
port 2 nsew
rlabel metal2 s 6000 237 6000 237 4 gnd
port 2 nsew
rlabel metal2 s 13968 237 13968 237 4 gnd
port 2 nsew
rlabel metal2 s 15216 237 15216 237 4 gnd
port 2 nsew
rlabel metal2 s 19968 347 19968 347 4 wl0_0
port 517 nsew
rlabel metal2 s 19968 127 19968 127 4 wl1_0
port 518 nsew
rlabel metal2 s 1008 0 1008 0 4 gnd
port 2 nsew
rlabel metal2 s 1488 0 1488 0 4 gnd
port 2 nsew
rlabel metal2 s 3984 0 3984 0 4 gnd
port 2 nsew
rlabel metal2 s 7728 0 7728 0 4 gnd
port 2 nsew
rlabel metal2 s 17232 0 17232 0 4 gnd
port 2 nsew
rlabel metal2 s 3504 0 3504 0 4 gnd
port 2 nsew
rlabel metal2 s 2256 0 2256 0 4 gnd
port 2 nsew
rlabel metal2 s 13488 0 13488 0 4 gnd
port 2 nsew
rlabel metal2 s 9744 0 9744 0 4 gnd
port 2 nsew
rlabel metal2 s 10224 0 10224 0 4 gnd
port 2 nsew
rlabel metal2 s 4752 0 4752 0 4 gnd
port 2 nsew
rlabel metal2 s 10992 0 10992 0 4 gnd
port 2 nsew
rlabel metal2 s 15984 0 15984 0 4 gnd
port 2 nsew
rlabel metal2 s 8496 0 8496 0 4 gnd
port 2 nsew
rlabel metal2 s 8976 0 8976 0 4 gnd
port 2 nsew
rlabel metal2 s 18960 0 18960 0 4 gnd
port 2 nsew
rlabel metal2 s 18480 0 18480 0 4 gnd
port 2 nsew
rlabel metal2 s 7248 0 7248 0 4 gnd
port 2 nsew
rlabel metal2 s 16464 0 16464 0 4 gnd
port 2 nsew
rlabel metal2 s 6000 0 6000 0 4 gnd
port 2 nsew
rlabel metal2 s 5232 0 5232 0 4 gnd
port 2 nsew
rlabel metal2 s 2736 0 2736 0 4 gnd
port 2 nsew
rlabel metal2 s 13968 0 13968 0 4 gnd
port 2 nsew
rlabel metal2 s 240 0 240 0 4 gnd
port 2 nsew
rlabel metal2 s 19728 0 19728 0 4 gnd
port 2 nsew
rlabel metal2 s 15216 0 15216 0 4 gnd
port 2 nsew
rlabel metal2 s 12720 0 12720 0 4 gnd
port 2 nsew
rlabel metal2 s 6480 0 6480 0 4 gnd
port 2 nsew
rlabel metal2 s 14736 0 14736 0 4 gnd
port 2 nsew
rlabel metal2 s 11472 0 11472 0 4 gnd
port 2 nsew
rlabel metal2 s 12240 0 12240 0 4 gnd
port 2 nsew
rlabel metal2 s 17712 0 17712 0 4 gnd
port 2 nsew
rlabel metal2 s 25968 0 25968 0 4 gnd
port 2 nsew
rlabel metal2 s 28944 0 28944 0 4 gnd
port 2 nsew
rlabel metal2 s 39696 0 39696 0 4 gnd
port 2 nsew
rlabel metal2 s 30192 0 30192 0 4 gnd
port 2 nsew
rlabel metal2 s 20208 0 20208 0 4 gnd
port 2 nsew
rlabel metal2 s 31440 0 31440 0 4 gnd
port 2 nsew
rlabel metal2 s 27216 0 27216 0 4 gnd
port 2 nsew
rlabel metal2 s 21456 0 21456 0 4 gnd
port 2 nsew
rlabel metal2 s 35952 0 35952 0 4 gnd
port 2 nsew
rlabel metal2 s 32208 0 32208 0 4 gnd
port 2 nsew
rlabel metal2 s 33456 0 33456 0 4 gnd
port 2 nsew
rlabel metal2 s 34704 0 34704 0 4 gnd
port 2 nsew
rlabel metal2 s 37200 0 37200 0 4 gnd
port 2 nsew
rlabel metal2 s 38928 0 38928 0 4 gnd
port 2 nsew
rlabel metal2 s 23952 0 23952 0 4 gnd
port 2 nsew
rlabel metal2 s 29712 0 29712 0 4 gnd
port 2 nsew
rlabel metal2 s 25200 0 25200 0 4 gnd
port 2 nsew
rlabel metal2 s 23472 0 23472 0 4 gnd
port 2 nsew
rlabel metal2 s 27696 0 27696 0 4 gnd
port 2 nsew
rlabel metal2 s 20976 0 20976 0 4 gnd
port 2 nsew
rlabel metal2 s 22704 0 22704 0 4 gnd
port 2 nsew
rlabel metal2 s 37680 0 37680 0 4 gnd
port 2 nsew
rlabel metal2 s 35184 0 35184 0 4 gnd
port 2 nsew
rlabel metal2 s 26448 0 26448 0 4 gnd
port 2 nsew
rlabel metal2 s 33936 0 33936 0 4 gnd
port 2 nsew
rlabel metal2 s 24720 0 24720 0 4 gnd
port 2 nsew
rlabel metal2 s 38448 0 38448 0 4 gnd
port 2 nsew
rlabel metal2 s 32688 0 32688 0 4 gnd
port 2 nsew
rlabel metal2 s 36432 0 36432 0 4 gnd
port 2 nsew
rlabel metal2 s 28464 0 28464 0 4 gnd
port 2 nsew
rlabel metal2 s 30960 0 30960 0 4 gnd
port 2 nsew
rlabel metal2 s 22224 0 22224 0 4 gnd
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 39936 395
string GDS_END 4456590
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4396370
<< end >>
