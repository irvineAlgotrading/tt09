magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -122 -66 534 666
<< mvpmos >>
rect 0 0 100 600
rect 156 0 256 600
rect 312 0 412 600
<< mvpdiff >>
rect -50 0 0 600
rect 412 0 462 600
<< poly >>
rect 0 600 100 632
rect 0 -32 100 0
rect 156 600 256 632
rect 156 -32 256 0
rect 312 600 412 632
rect 312 -32 412 0
<< locali >>
rect -45 -4 -11 538
rect 111 -4 145 538
rect 267 -4 301 538
rect 423 -4 457 538
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1704896540
transform 1 0 256 0 1 0
box -36 -36 92 636
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_1
timestamp 1704896540
transform 1 0 100 0 1 0
box -36 -36 92 636
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 92 636
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_1
timestamp 1704896540
transform 1 0 412 0 1 0
box -36 -36 92 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 440 267 440 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85603492
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85601478
<< end >>
