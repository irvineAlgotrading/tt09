magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 6786 897
<< pwell >>
rect 4 43 6706 317
rect -26 -43 6746 43
<< locali >>
rect 44 316 926 363
<< obsli1 >>
rect 0 797 6720 831
rect 22 435 136 751
rect 170 453 232 751
rect 268 489 446 735
rect 480 453 542 751
rect 576 489 754 735
rect 788 453 858 751
rect 892 489 1070 735
rect 1104 453 1166 751
rect 1200 489 1378 735
rect 1412 453 1482 751
rect 170 397 1482 453
rect 1516 447 1696 735
rect 960 282 1482 397
rect 22 85 129 282
rect 163 239 1482 282
rect 163 151 234 239
rect 268 83 446 205
rect 480 146 558 239
rect 592 85 771 205
rect 805 146 854 239
rect 888 85 1066 205
rect 1104 146 1182 239
rect 1216 85 1395 205
rect 1429 146 1478 239
rect 1516 205 1696 279
rect 1512 85 1696 205
rect 1786 158 1852 751
rect 1886 435 2064 751
rect 1904 313 2038 379
rect 1886 85 2064 279
rect 2098 158 2164 751
rect 2198 435 2376 751
rect 2216 313 2350 379
rect 2198 85 2376 279
rect 2410 158 2476 751
rect 2510 435 2688 751
rect 2528 313 2662 379
rect 2510 85 2688 279
rect 2722 158 2788 751
rect 2822 435 3000 751
rect 2840 313 2974 379
rect 2822 85 3000 279
rect 3034 158 3100 751
rect 3134 435 3312 751
rect 3152 313 3286 379
rect 3134 85 3312 279
rect 3346 158 3412 751
rect 3446 435 3624 751
rect 3464 313 3598 379
rect 3446 85 3624 279
rect 3658 158 3724 751
rect 3758 435 3936 751
rect 3776 313 3910 379
rect 3758 85 3936 279
rect 3970 158 4052 751
rect 4086 435 4192 751
rect 4086 313 4220 379
rect 4086 85 4192 279
rect 4282 158 4348 751
rect 4382 435 4560 751
rect 4400 313 4534 379
rect 4382 85 4560 279
rect 4594 158 4660 751
rect 4694 435 4872 751
rect 4712 313 4846 379
rect 4694 85 4872 279
rect 4906 158 4972 751
rect 5006 435 5184 751
rect 5024 313 5158 379
rect 5006 85 5184 279
rect 5218 158 5284 751
rect 5318 435 5496 751
rect 5336 313 5470 379
rect 5318 85 5496 279
rect 5530 158 5596 751
rect 5630 435 5808 751
rect 5648 313 5782 379
rect 5630 85 5808 279
rect 5842 158 5908 751
rect 5942 435 6120 751
rect 5960 313 6094 379
rect 5942 85 6120 279
rect 6154 158 6220 751
rect 6254 435 6432 751
rect 6272 313 6406 379
rect 6254 85 6432 279
rect 6466 158 6548 751
rect 6582 435 6688 751
rect 6582 85 6688 299
rect 0 -17 6720 17
<< metal1 >>
rect 0 791 6720 837
rect 0 689 6720 763
rect 1790 458 6528 504
rect 0 51 6720 125
rect 0 -23 6720 23
<< obsm1 >>
rect 992 310 6418 356
<< labels >>
rlabel locali s 44 316 926 363 6 A
port 1 nsew signal input
rlabel metal1 s 0 51 6720 125 6 VGND
port 2 nsew ground bidirectional
rlabel metal1 s 0 -23 6720 23 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s -26 -43 6746 43 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 4 43 6706 317 6 VNB
port 3 nsew ground bidirectional
rlabel metal1 s 0 791 6720 837 6 VPB
port 4 nsew power bidirectional
rlabel nwell s -66 377 6786 897 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 689 6720 763 6 VPWR
port 5 nsew power bidirectional
rlabel metal1 s 1790 458 6528 504 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 6720 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1091352
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1031596
<< end >>
