magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect -50 -1408 0 -1392
rect -50 -1442 -34 -1408
rect -50 -1458 0 -1442
<< polycont >>
rect -34 16 0 50
rect -34 -1442 0 -1408
<< npolyres >>
rect 0 0 30933 66
rect 30867 -96 30933 0
rect -50 -162 30933 -96
rect -50 -258 16 -162
rect -50 -324 30933 -258
rect 30867 -420 30933 -324
rect -50 -486 30933 -420
rect -50 -582 16 -486
rect -50 -648 30933 -582
rect 30867 -744 30933 -648
rect -50 -810 30933 -744
rect -50 -906 16 -810
rect -50 -972 30933 -906
rect 30867 -1068 30933 -972
rect -50 -1134 30933 -1068
rect -50 -1230 16 -1134
rect -50 -1296 30933 -1230
rect 30867 -1392 30933 -1296
rect 0 -1458 30933 -1392
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect -34 -1408 0 -1392
rect -34 -1458 0 -1442
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform 1 0 -50 0 1 -1458
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform 1 0 -50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 34340492
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34337708
<< end >>
