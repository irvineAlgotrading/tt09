magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 2956 -1894 3007 -1878
rect 2990 -1928 3007 -1894
rect 2956 -1944 3007 -1928
<< polycont >>
rect -34 16 0 50
rect 2956 -1928 2990 -1894
<< npolyres >>
rect 0 0 3007 66
rect 2941 -96 3007 0
rect -50 -162 3007 -96
rect -50 -258 16 -162
rect -50 -324 3007 -258
rect 2941 -420 3007 -324
rect -50 -486 3007 -420
rect -50 -582 16 -486
rect -50 -648 3007 -582
rect 2941 -744 3007 -648
rect -50 -810 3007 -744
rect -50 -906 16 -810
rect -50 -972 3007 -906
rect 2941 -1068 3007 -972
rect -50 -1134 3007 -1068
rect -50 -1230 16 -1134
rect -50 -1296 3007 -1230
rect 2941 -1392 3007 -1296
rect -50 -1458 3007 -1392
rect -50 -1554 16 -1458
rect -50 -1620 3007 -1554
rect 2941 -1716 3007 -1620
rect -50 -1782 3007 -1716
rect -50 -1878 16 -1782
rect -50 -1944 2956 -1878
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 2956 -1894 2991 -1878
rect 2990 -1928 2991 -1894
rect 2956 -1944 2991 -1928
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_0
timestamp 1704896540
transform 1 0 -50 0 1 0
box 0 0 1 1
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_1
timestamp 1704896540
transform 1 0 2940 0 1 -1944
box 0 0 1 1
<< properties >>
string GDS_END 42934138
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42930518
<< end >>
