magic
tech sky130A
timestamp 1704896540
<< pwell >>
rect -13 -13 163 1513
<< nsubdiff >>
rect 0 0 150 1500
use s8_esd_gnd2gnd_strap  s8_esd_gnd2gnd_strap_0
timestamp 1704896540
transform 1 0 0 0 1 0
box 0 0 150 1500
<< properties >>
string GDS_END 42971550
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42971374
<< end >>
