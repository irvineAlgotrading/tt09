magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 0 0 564 534
<< pmos >>
rect 204 102 254 432
rect 310 102 360 432
<< pdiff >>
rect 148 420 204 432
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 254 420 310 432
rect 254 386 265 420
rect 299 386 310 420
rect 254 352 310 386
rect 254 318 265 352
rect 299 318 310 352
rect 254 284 310 318
rect 254 250 265 284
rect 299 250 310 284
rect 254 216 310 250
rect 254 182 265 216
rect 299 182 310 216
rect 254 148 310 182
rect 254 114 265 148
rect 299 114 310 148
rect 254 102 310 114
rect 360 420 416 432
rect 360 386 371 420
rect 405 386 416 420
rect 360 352 416 386
rect 360 318 371 352
rect 405 318 416 352
rect 360 284 416 318
rect 360 250 371 284
rect 405 250 416 284
rect 360 216 416 250
rect 360 182 371 216
rect 405 182 416 216
rect 360 148 416 182
rect 360 114 371 148
rect 405 114 416 148
rect 360 102 416 114
<< pdiffc >>
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 265 386 299 420
rect 265 318 299 352
rect 265 250 299 284
rect 265 182 299 216
rect 265 114 299 148
rect 371 386 405 420
rect 371 318 405 352
rect 371 250 405 284
rect 371 182 405 216
rect 371 114 405 148
<< nsubdiff >>
rect 36 386 94 432
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 470 386 528 432
rect 470 352 482 386
rect 516 352 528 386
rect 470 318 528 352
rect 470 284 482 318
rect 516 284 528 318
rect 470 250 528 284
rect 470 216 482 250
rect 516 216 528 250
rect 470 182 528 216
rect 470 148 482 182
rect 516 148 528 182
rect 470 102 528 148
<< nsubdiffcont >>
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 482 352 516 386
rect 482 284 516 318
rect 482 216 516 250
rect 482 148 516 182
<< poly >>
rect 181 514 383 534
rect 181 480 197 514
rect 231 480 265 514
rect 299 480 333 514
rect 367 480 383 514
rect 181 464 383 480
rect 204 432 254 464
rect 310 432 360 464
rect 204 70 254 102
rect 310 70 360 102
rect 181 54 383 70
rect 181 20 197 54
rect 231 20 265 54
rect 299 20 333 54
rect 367 20 383 54
rect 181 0 383 20
<< polycont >>
rect 197 480 231 514
rect 265 480 299 514
rect 333 480 367 514
rect 197 20 231 54
rect 265 20 299 54
rect 333 20 367 54
<< locali >>
rect 181 480 193 514
rect 231 480 265 514
rect 299 480 333 514
rect 371 480 383 514
rect 159 420 193 436
rect 48 392 82 402
rect 48 320 82 352
rect 48 250 82 284
rect 48 182 82 214
rect 48 132 82 142
rect 159 352 193 358
rect 159 284 193 286
rect 159 248 193 250
rect 159 176 193 182
rect 159 98 193 114
rect 265 420 299 436
rect 265 352 299 358
rect 265 284 299 286
rect 265 248 299 250
rect 265 176 299 182
rect 265 98 299 114
rect 371 420 405 436
rect 371 352 405 358
rect 371 284 405 286
rect 371 248 405 250
rect 371 176 405 182
rect 482 392 516 402
rect 482 320 516 352
rect 482 250 516 284
rect 482 182 516 214
rect 482 132 516 142
rect 371 98 405 114
rect 181 20 193 54
rect 231 20 265 54
rect 299 20 333 54
rect 371 20 383 54
<< viali >>
rect 193 480 197 514
rect 197 480 227 514
rect 265 480 299 514
rect 337 480 367 514
rect 367 480 371 514
rect 48 386 82 392
rect 48 358 82 386
rect 48 318 82 320
rect 48 286 82 318
rect 48 216 82 248
rect 48 214 82 216
rect 48 148 82 176
rect 48 142 82 148
rect 159 386 193 392
rect 159 358 193 386
rect 159 318 193 320
rect 159 286 193 318
rect 159 216 193 248
rect 159 214 193 216
rect 159 148 193 176
rect 159 142 193 148
rect 265 386 299 392
rect 265 358 299 386
rect 265 318 299 320
rect 265 286 299 318
rect 265 216 299 248
rect 265 214 299 216
rect 265 148 299 176
rect 265 142 299 148
rect 371 386 405 392
rect 371 358 405 386
rect 371 318 405 320
rect 371 286 405 318
rect 371 216 405 248
rect 371 214 405 216
rect 371 148 405 176
rect 371 142 405 148
rect 482 386 516 392
rect 482 358 516 386
rect 482 318 516 320
rect 482 286 516 318
rect 482 216 516 248
rect 482 214 516 216
rect 482 148 516 176
rect 482 142 516 148
rect 193 20 197 54
rect 197 20 227 54
rect 265 20 299 54
rect 337 20 367 54
rect 367 20 371 54
<< metal1 >>
rect 181 514 383 534
rect 181 480 193 514
rect 227 480 265 514
rect 299 480 337 514
rect 371 480 383 514
rect 181 468 383 480
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 150 392 202 420
rect 150 358 159 392
rect 193 358 202 392
rect 150 320 202 358
rect 150 286 159 320
rect 193 286 202 320
rect 150 248 202 286
rect 150 236 159 248
rect 193 236 202 248
rect 150 176 202 184
rect 150 172 159 176
rect 193 172 202 176
rect 150 114 202 120
rect 256 414 308 420
rect 256 358 265 362
rect 299 358 308 362
rect 256 350 308 358
rect 256 286 265 298
rect 299 286 308 298
rect 256 248 308 286
rect 256 214 265 248
rect 299 214 308 248
rect 256 176 308 214
rect 256 142 265 176
rect 299 142 308 176
rect 256 114 308 142
rect 362 392 414 420
rect 362 358 371 392
rect 405 358 414 392
rect 362 320 414 358
rect 362 286 371 320
rect 405 286 414 320
rect 362 248 414 286
rect 362 236 371 248
rect 405 236 414 248
rect 362 176 414 184
rect 362 172 371 176
rect 405 172 414 176
rect 362 114 414 120
rect 470 392 528 420
rect 470 358 482 392
rect 516 358 528 392
rect 470 320 528 358
rect 470 286 482 320
rect 516 286 528 320
rect 470 248 528 286
rect 470 214 482 248
rect 516 214 528 248
rect 470 176 528 214
rect 470 142 482 176
rect 516 142 528 176
rect 470 114 528 142
rect 181 54 383 66
rect 181 20 193 54
rect 227 20 265 54
rect 299 20 337 54
rect 371 20 383 54
rect 181 0 383 20
<< via1 >>
rect 150 214 159 236
rect 159 214 193 236
rect 193 214 202 236
rect 150 184 202 214
rect 150 142 159 172
rect 159 142 193 172
rect 193 142 202 172
rect 150 120 202 142
rect 256 392 308 414
rect 256 362 265 392
rect 265 362 299 392
rect 299 362 308 392
rect 256 320 308 350
rect 256 298 265 320
rect 265 298 299 320
rect 299 298 308 320
rect 362 214 371 236
rect 371 214 405 236
rect 405 214 414 236
rect 362 184 414 214
rect 362 142 371 172
rect 371 142 405 172
rect 405 142 414 172
rect 362 120 414 142
<< metal2 >>
rect 10 414 554 420
rect 10 362 256 414
rect 308 362 554 414
rect 10 350 554 362
rect 10 298 256 350
rect 308 298 554 350
rect 10 292 554 298
rect 10 236 554 242
rect 10 184 150 236
rect 202 184 362 236
rect 414 184 554 236
rect 10 172 554 184
rect 10 120 150 172
rect 202 120 362 172
rect 414 120 554 172
rect 10 114 554 120
<< labels >>
flabel metal2 s 10 114 30 242 7 FreeSans 300 180 0 0 SOURCE
port 2 nsew
flabel metal2 s 10 292 30 420 7 FreeSans 300 180 0 0 DRAIN
port 3 nsew
flabel metal1 s 470 114 528 130 3 FreeSans 300 90 0 0 BULK
port 4 nsew
flabel metal1 s 181 0 383 66 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 181 468 383 534 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 36 114 94 130 3 FreeSans 300 90 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9251662
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9244010
<< end >>
