magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -68 -26 948 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 880 50 922 66
rect 914 16 922 50
rect 880 0 922 16
<< ndiffc >>
rect -34 16 0 50
rect 880 16 914 50
<< ndiffres >>
rect 0 0 880 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 880 50 914 66
rect 880 0 914 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 1 0 872 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 97474852
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97474350
<< end >>
