magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -98 -26 282 176
<< mvnmos >>
rect 0 0 200 150
<< mvndiff >>
rect -72 114 0 150
rect -72 80 -61 114
rect -27 80 0 114
rect -72 46 0 80
rect -72 12 -61 46
rect -27 12 0 46
rect -72 0 0 12
rect 200 114 256 150
rect 200 80 211 114
rect 245 80 256 114
rect 200 46 256 80
rect 200 12 211 46
rect 245 12 256 46
rect 200 0 256 12
<< mvndiffc >>
rect -61 80 -27 114
rect -61 12 -27 46
rect 211 80 245 114
rect 211 12 245 46
<< poly >>
rect 0 150 200 182
rect 0 -32 200 0
<< locali >>
rect -61 114 -27 130
rect -61 46 -27 80
rect -61 -4 -27 12
rect 211 114 245 130
rect 211 46 245 80
rect 211 -4 245 12
use hvDFL1sd2_CDNS_52468879185235  hvDFL1sd2_CDNS_52468879185235_0
timestamp 1704896540
transform -1 0 -16 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185235  hvDFL1sd2_CDNS_52468879185235_1
timestamp 1704896540
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -44 63 -44 63 0 FreeSans 300 0 0 0 S
flabel comment s 228 63 228 63 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85638372
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85637414
<< end >>
