magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__dfm1sd2__example_55959141808197  sky130_fd_pr__dfm1sd2__example_55959141808197_0
timestamp 1704896540
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfm1sd2__example_55959141808197  sky130_fd_pr__dfm1sd2__example_55959141808197_1
timestamp 1704896540
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808194  sky130_fd_pr__hvdfl1sd__example_55959141808194_0
timestamp 1704896540
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_0
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_1
timestamp 1704896540
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_2
timestamp 1704896540
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180848  sky130_fd_pr__hvdfm1sd__example_5595914180848_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 68177666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 68174032
<< end >>
