magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 353 0 400
rect -50 319 -34 353
rect -50 285 0 319
rect -50 251 -34 285
rect -50 217 0 251
rect -50 183 -34 217
rect -50 149 0 183
rect -50 115 -34 149
rect -50 81 0 115
rect -50 47 -34 81
rect -50 0 0 47
rect 2000 353 2050 400
rect 2034 319 2050 353
rect 2000 285 2050 319
rect 2034 251 2050 285
rect 2000 217 2050 251
rect 2034 183 2050 217
rect 2000 149 2050 183
rect 2034 115 2050 149
rect 2000 81 2050 115
rect 2034 47 2050 81
rect 2000 0 2050 47
<< polycont >>
rect -34 319 0 353
rect -34 251 0 285
rect -34 183 0 217
rect -34 115 0 149
rect -34 47 0 81
rect 2000 319 2034 353
rect 2000 251 2034 285
rect 2000 183 2034 217
rect 2000 115 2034 149
rect 2000 47 2034 81
<< npolyres >>
rect 0 0 2000 400
<< locali >>
rect -34 353 0 369
rect -34 285 0 319
rect -34 217 0 251
rect -34 149 0 183
rect -34 81 0 115
rect -34 31 0 47
rect 2000 353 2034 369
rect 2000 285 2034 319
rect 2000 217 2034 251
rect 2000 149 2034 183
rect 2000 81 2034 115
rect 2000 31 2034 47
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1704896540
transform -1 0 16 0 1 31
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_1
timestamp 1704896540
transform 1 0 1984 0 1 31
box 0 0 1 1
<< properties >>
string GDS_END 94169472
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94169034
<< end >>
