magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 -36 92 3036
<< pdiff >>
rect 0 2970 56 3000
rect 0 2936 11 2970
rect 45 2936 56 2970
rect 0 2902 56 2936
rect 0 2868 11 2902
rect 45 2868 56 2902
rect 0 2834 56 2868
rect 0 2800 11 2834
rect 45 2800 56 2834
rect 0 2766 56 2800
rect 0 2732 11 2766
rect 45 2732 56 2766
rect 0 2698 56 2732
rect 0 2664 11 2698
rect 45 2664 56 2698
rect 0 2630 56 2664
rect 0 2596 11 2630
rect 45 2596 56 2630
rect 0 2562 56 2596
rect 0 2528 11 2562
rect 45 2528 56 2562
rect 0 2494 56 2528
rect 0 2460 11 2494
rect 45 2460 56 2494
rect 0 2426 56 2460
rect 0 2392 11 2426
rect 45 2392 56 2426
rect 0 2358 56 2392
rect 0 2324 11 2358
rect 45 2324 56 2358
rect 0 2290 56 2324
rect 0 2256 11 2290
rect 45 2256 56 2290
rect 0 2222 56 2256
rect 0 2188 11 2222
rect 45 2188 56 2222
rect 0 2154 56 2188
rect 0 2120 11 2154
rect 45 2120 56 2154
rect 0 2086 56 2120
rect 0 2052 11 2086
rect 45 2052 56 2086
rect 0 2018 56 2052
rect 0 1984 11 2018
rect 45 1984 56 2018
rect 0 1950 56 1984
rect 0 1916 11 1950
rect 45 1916 56 1950
rect 0 1882 56 1916
rect 0 1848 11 1882
rect 45 1848 56 1882
rect 0 1814 56 1848
rect 0 1780 11 1814
rect 45 1780 56 1814
rect 0 1746 56 1780
rect 0 1712 11 1746
rect 45 1712 56 1746
rect 0 1678 56 1712
rect 0 1644 11 1678
rect 45 1644 56 1678
rect 0 1610 56 1644
rect 0 1576 11 1610
rect 45 1576 56 1610
rect 0 1542 56 1576
rect 0 1508 11 1542
rect 45 1508 56 1542
rect 0 1474 56 1508
rect 0 1440 11 1474
rect 45 1440 56 1474
rect 0 1406 56 1440
rect 0 1372 11 1406
rect 45 1372 56 1406
rect 0 1338 56 1372
rect 0 1304 11 1338
rect 45 1304 56 1338
rect 0 1270 56 1304
rect 0 1236 11 1270
rect 45 1236 56 1270
rect 0 1202 56 1236
rect 0 1168 11 1202
rect 45 1168 56 1202
rect 0 1134 56 1168
rect 0 1100 11 1134
rect 45 1100 56 1134
rect 0 1066 56 1100
rect 0 1032 11 1066
rect 45 1032 56 1066
rect 0 998 56 1032
rect 0 964 11 998
rect 45 964 56 998
rect 0 930 56 964
rect 0 896 11 930
rect 45 896 56 930
rect 0 862 56 896
rect 0 828 11 862
rect 45 828 56 862
rect 0 794 56 828
rect 0 760 11 794
rect 45 760 56 794
rect 0 726 56 760
rect 0 692 11 726
rect 45 692 56 726
rect 0 658 56 692
rect 0 624 11 658
rect 45 624 56 658
rect 0 590 56 624
rect 0 556 11 590
rect 45 556 56 590
rect 0 522 56 556
rect 0 488 11 522
rect 45 488 56 522
rect 0 454 56 488
rect 0 420 11 454
rect 45 420 56 454
rect 0 386 56 420
rect 0 352 11 386
rect 45 352 56 386
rect 0 318 56 352
rect 0 284 11 318
rect 45 284 56 318
rect 0 250 56 284
rect 0 216 11 250
rect 45 216 56 250
rect 0 182 56 216
rect 0 148 11 182
rect 45 148 56 182
rect 0 114 56 148
rect 0 80 11 114
rect 45 80 56 114
rect 0 46 56 80
rect 0 12 11 46
rect 45 12 56 46
rect 0 0 56 12
<< pdiffc >>
rect 11 2936 45 2970
rect 11 2868 45 2902
rect 11 2800 45 2834
rect 11 2732 45 2766
rect 11 2664 45 2698
rect 11 2596 45 2630
rect 11 2528 45 2562
rect 11 2460 45 2494
rect 11 2392 45 2426
rect 11 2324 45 2358
rect 11 2256 45 2290
rect 11 2188 45 2222
rect 11 2120 45 2154
rect 11 2052 45 2086
rect 11 1984 45 2018
rect 11 1916 45 1950
rect 11 1848 45 1882
rect 11 1780 45 1814
rect 11 1712 45 1746
rect 11 1644 45 1678
rect 11 1576 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1474
rect 11 1372 45 1406
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 2970 45 2986
rect 11 2902 45 2936
rect 11 2834 45 2868
rect 11 2766 45 2800
rect 11 2698 45 2732
rect 11 2630 45 2664
rect 11 2562 45 2596
rect 11 2494 45 2528
rect 11 2426 45 2460
rect 11 2358 45 2392
rect 11 2290 45 2324
rect 11 2222 45 2256
rect 11 2154 45 2188
rect 11 2086 45 2120
rect 11 2018 45 2052
rect 11 1950 45 1984
rect 11 1882 45 1916
rect 11 1814 45 1848
rect 11 1746 45 1780
rect 11 1678 45 1712
rect 11 1610 45 1644
rect 11 1542 45 1576
rect 11 1474 45 1508
rect 11 1406 45 1440
rect 11 1338 45 1372
rect 11 1270 45 1304
rect 11 1202 45 1236
rect 11 1134 45 1168
rect 11 1066 45 1100
rect 11 998 45 1032
rect 11 930 45 964
rect 11 862 45 896
rect 11 794 45 828
rect 11 726 45 760
rect 11 658 45 692
rect 11 590 45 624
rect 11 522 45 556
rect 11 454 45 488
rect 11 386 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 216
rect 11 114 45 148
rect 11 46 45 80
rect 11 -4 45 12
<< properties >>
string GDS_END 88574060
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88570984
<< end >>
