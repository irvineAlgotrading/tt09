magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 2200 50 2250 66
rect 2234 16 2250 50
rect 2200 0 2250 16
<< polycont >>
rect -34 16 0 50
rect 2200 16 2234 50
<< npolyres >>
rect 0 0 2200 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 2200 50 2234 66
rect 2200 0 2234 16
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform -1 0 16 0 1 0
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform 1 0 2184 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 87731654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87731220
<< end >>
