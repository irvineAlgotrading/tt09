magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect -50 -1732 6 -1716
rect -50 -1766 -28 -1732
rect -50 -1782 6 -1766
<< polycont >>
rect -34 16 0 50
rect -28 -1766 6 -1732
<< npolyres >>
rect 0 0 11598 66
rect 11532 -96 11598 0
rect -50 -162 11598 -96
rect -50 -258 16 -162
rect -50 -324 11598 -258
rect 11532 -420 11598 -324
rect -50 -486 11598 -420
rect -50 -582 16 -486
rect -50 -648 11598 -582
rect 11532 -744 11598 -648
rect -50 -810 11598 -744
rect -50 -906 16 -810
rect -50 -972 11598 -906
rect 11532 -1068 11598 -972
rect -50 -1134 11598 -1068
rect -50 -1230 16 -1134
rect -50 -1296 11598 -1230
rect 11532 -1392 11598 -1296
rect -50 -1458 11598 -1392
rect -50 -1554 16 -1458
rect -50 -1620 11598 -1554
rect 11532 -1716 11598 -1620
rect 6 -1782 11598 -1716
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect -34 -1732 6 -1716
rect -34 -1766 -28 -1732
rect -34 -1782 6 -1766
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform 1 0 -44 0 1 -1782
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform 1 0 -50 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 34413064
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34409768
<< end >>
