* NGSPICE file created from tt_um_audio_player.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

.subckt tt_um_audio_player VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
XTAP_TAPCELL_ROW_17_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1270_ _0953_/X _1342_/B _1154_/X _1269_/X VGND VGND VPWR VPWR _1270_/X sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_14_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1606_ clkload0/A _1606_/D fanout120/X VGND VGND VPWR VPWR _1606_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0985_ _0953_/A _0985_/B VGND VGND VPWR VPWR _1362_/C sky130_fd_sc_hd__nand2b_4
XFILLER_0_14_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1537_ _1229_/A _1357_/A _1562_/B _1542_/B _1236_/B VGND VGND VPWR VPWR _1589_/D
+ sky130_fd_sc_hd__a32o_1
Xfanout116 _0787_/Y VGND VGND VPWR VPWR _1525_/B sky130_fd_sc_hd__buf_2
X_1399_ _1399_/A _1399_/B VGND VGND VPWR VPWR _1399_/Y sky130_fd_sc_hd__nor2_1
Xfanout105 _0851_/D VGND VGND VPWR VPWR _0849_/B sky130_fd_sc_hd__buf_4
XFILLER_0_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1468_ _0996_/A _1467_/Y _1193_/X VGND VGND VPWR VPWR _1468_/Y sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_6_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1322_ _1316_/X _1318_/Y _1321_/X _0843_/Y VGND VGND VPWR VPWR _1322_/X sky130_fd_sc_hd__o31a_1
X_1253_ _0816_/A _0816_/B _1085_/Y _0888_/B _0930_/D VGND VGND VPWR VPWR _1253_/X
+ sky130_fd_sc_hd__a311o_1
X_1184_ _1184_/A _1362_/B _1362_/D VGND VGND VPWR VPWR _1184_/X sky130_fd_sc_hd__or3_1
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0968_ _1035_/A _1036_/A VGND VGND VPWR VPWR _1398_/B sky130_fd_sc_hd__nor2_1
X_0899_ _0900_/A _1539_/A _0900_/C _1236_/B VGND VGND VPWR VPWR _1147_/B sky130_fd_sc_hd__nor4_2
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0822_ _1398_/A _1339_/B VGND VGND VPWR VPWR _1420_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1236_ _1534_/S _1236_/B _1236_/C _1236_/D VGND VGND VPWR VPWR _1237_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1305_ _0854_/X _1339_/D _1043_/B _0953_/A VGND VGND VPWR VPWR _1305_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1098_ _1323_/B _1098_/B VGND VGND VPWR VPWR _1098_/X sky130_fd_sc_hd__or2_1
X_1167_ _1252_/A _1411_/C _1442_/A VGND VGND VPWR VPWR _1167_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1021_ _1190_/B _1021_/B VGND VGND VPWR VPWR _1021_/Y sky130_fd_sc_hd__nor2_1
X_0805_ hold4/A _1605_/Q _1606_/Q VGND VGND VPWR VPWR _0807_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_24_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1219_ _0996_/A _1237_/A _0936_/Y _1218_/Y _0914_/Y VGND VGND VPWR VPWR _1219_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1570_ hold12/A _1570_/B _1570_/C VGND VGND VPWR VPWR _1570_/X sky130_fd_sc_hd__and3_1
XANTENNA_5 _1036_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1004_ _0926_/A _0962_/B _0989_/A VGND VGND VPWR VPWR _1004_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1553_ _0903_/B _1548_/X _1247_/B VGND VGND VPWR VPWR _1554_/B sky130_fd_sc_hd__a21o_1
X_1484_ _1454_/B _1261_/X _1479_/Y _1481_/X _1116_/C VGND VGND VPWR VPWR _1484_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_17_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0984_ _0991_/A _1398_/A VGND VGND VPWR VPWR _1434_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1605_ clkload0/A _1605_/D fanout120/X VGND VGND VPWR VPWR _1605_/Q sky130_fd_sc_hd__dfrtp_1
X_1536_ _1542_/B _1544_/B VGND VGND VPWR VPWR _1562_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_22_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout117 fanout119/X VGND VGND VPWR VPWR fanout117/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout106 _0851_/D VGND VGND VPWR VPWR _1236_/B sky130_fd_sc_hd__buf_4
X_1398_ _1398_/A _1398_/B _1398_/C VGND VGND VPWR VPWR _1398_/X sky130_fd_sc_hd__or3_1
X_1467_ _1146_/B _1343_/C _1028_/X VGND VGND VPWR VPWR _1467_/Y sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_6_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1252_ _1252_/A _1252_/B _1252_/C VGND VGND VPWR VPWR _1252_/X sky130_fd_sc_hd__or3_1
X_1321_ _1135_/B _1299_/Y _1320_/X _1114_/A VGND VGND VPWR VPWR _1321_/X sky130_fd_sc_hd__o211a_1
X_1183_ _1183_/A _1183_/B VGND VGND VPWR VPWR _1183_/Y sky130_fd_sc_hd__nand2_1
X_0967_ _0960_/X _0964_/Y _0966_/X _1560_/A VGND VGND VPWR VPWR _0967_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1519_ _1497_/Y _1517_/Y _1518_/X _1524_/B hold11/X VGND VGND VPWR VPWR _1582_/D
+ sky130_fd_sc_hd__a32o_1
X_0898_ _0844_/X _0887_/X _0897_/X VGND VGND VPWR VPWR _0898_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0821_ _0931_/B _1035_/A _0985_/B VGND VGND VPWR VPWR _1281_/A sky130_fd_sc_hd__nand3_2
XPHY_EDGE_ROW_24_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1166_ _1166_/A _1599_/Q VGND VGND VPWR VPWR _1488_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1235_ _1232_/X _1234_/X _1555_/A VGND VGND VPWR VPWR _1235_/X sky130_fd_sc_hd__o21a_1
X_1304_ _1304_/A1 _1043_/B _1303_/X _1323_/A _1039_/B VGND VGND VPWR VPWR _1304_/X
+ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_22_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1097_ _0953_/X _1029_/Y _1181_/D _1096_/X VGND VGND VPWR VPWR _1098_/B sky130_fd_sc_hd__o22a_1
XFILLER_0_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1020_ _1260_/A _1544_/A VGND VGND VPWR VPWR _1020_/X sky130_fd_sc_hd__or2_1
X_0804_ hold14/X _1605_/Q _0803_/Y VGND VGND VPWR VPWR _1605_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1218_ _1218_/A1 _1037_/A _0869_/A VGND VGND VPWR VPWR _1218_/Y sky130_fd_sc_hd__o21ai_2
X_1149_ _1439_/A _1408_/C _1436_/A _1148_/X _1205_/B VGND VGND VPWR VPWR _1149_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 _1036_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1003_ _0997_/X _1002_/Y _1116_/C VGND VGND VPWR VPWR _1423_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1552_ _1544_/B _1560_/C _1560_/B VGND VGND VPWR VPWR _1555_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1483_ _1483_/A _1483_/B _1483_/C _1483_/D VGND VGND VPWR VPWR _1483_/X sky130_fd_sc_hd__or4_1
XFILLER_0_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0983_ _1339_/B _1212_/B _1339_/C _0978_/X VGND VGND VPWR VPWR _0983_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout118 fanout119/X VGND VGND VPWR VPWR fanout118/X sky130_fd_sc_hd__clkbuf_4
X_1604_ clkload0/A _1604_/D fanout120/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfrtp_2
X_1535_ _1442_/A _0991_/X _1527_/X _1533_/A VGND VGND VPWR VPWR _1544_/B sky130_fd_sc_hd__a31o_2
Xfanout107 _1335_/A VGND VGND VPWR VPWR _0851_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1466_ _1190_/A _1462_/X _1465_/X _1166_/A _1458_/X VGND VGND VPWR VPWR _1466_/X
+ sky130_fd_sc_hd__o311a_1
X_1397_ _0926_/A _0962_/B _1056_/B VGND VGND VPWR VPWR _1398_/C sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ _1323_/A _1320_/B _1320_/C _1320_/D VGND VGND VPWR VPWR _1320_/X sky130_fd_sc_hd__or4_1
X_1251_ _1251_/A _1251_/B _1251_/C VGND VGND VPWR VPWR _1489_/B sky130_fd_sc_hd__or3_1
X_1182_ _1178_/X _1180_/Y _1181_/X _1010_/A VGND VGND VPWR VPWR _1182_/X sky130_fd_sc_hd__a31o_1
X_0966_ _0819_/X _0903_/A _1352_/A _0965_/X VGND VGND VPWR VPWR _0966_/X sky130_fd_sc_hd__a31o_1
X_0897_ _0876_/X _0891_/X _1434_/A _0890_/X VGND VGND VPWR VPWR _0897_/X sky130_fd_sc_hd__o211a_1
X_1518_ hold11/A _1518_/B VGND VGND VPWR VPWR _1518_/X sky130_fd_sc_hd__or2_1
X_1449_ _0926_/A _1420_/C _1420_/D _1082_/Y VGND VGND VPWR VPWR _1449_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap7 _1028_/B VGND VGND VPWR VPWR _1060_/B1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0820_ _1362_/B _0985_/B VGND VGND VPWR VPWR _1114_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1303_ _1319_/B _1029_/B _0888_/B _0928_/B VGND VGND VPWR VPWR _1303_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1234_ _1180_/A _1004_/Y _1233_/Y _0885_/B VGND VGND VPWR VPWR _1234_/X sky130_fd_sc_hd__a22o_1
X_1165_ _1526_/D _1159_/X _1160_/X _1164_/X VGND VGND VPWR VPWR _1165_/X sky130_fd_sc_hd__a31o_1
X_1096_ _1229_/A _1300_/D _1475_/A _0928_/B _0975_/Y VGND VGND VPWR VPWR _1096_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_22_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0949_ _1094_/A _1199_/C VGND VGND VPWR VPWR _1384_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0803_ hold4/A _1605_/Q _1525_/B VGND VGND VPWR VPWR _0803_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1217_ _1180_/A _0947_/Y _1066_/A VGND VGND VPWR VPWR _1217_/Y sky130_fd_sc_hd__a21oi_1
X_1148_ _0816_/B _1304_/A1 _1343_/C wire10/X VGND VGND VPWR VPWR _1148_/X sky130_fd_sc_hd__a31o_1
X_1079_ _0952_/B _0818_/Y _0876_/X _1078_/X _1066_/A VGND VGND VPWR VPWR _1079_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_7 _1183_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1002_ _1218_/A1 _1197_/B _0891_/X _1452_/A VGND VGND VPWR VPWR _1002_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1551_ _1551_/A _1551_/B _1551_/C VGND VGND VPWR VPWR _1560_/C sky130_fd_sc_hd__and3_1
XFILLER_0_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1482_ _0930_/D _1319_/B _0923_/B _1146_/B VGND VGND VPWR VPWR _1483_/D sky130_fd_sc_hd__o22ai_1
XFILLER_0_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0982_ _1339_/B _1339_/C VGND VGND VPWR VPWR _1399_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1603_ clkload1/A _1603_/D fanout117/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfrtp_1
X_1534_ _1533_/Y _1542_/B _1534_/S VGND VGND VPWR VPWR _1588_/D sky130_fd_sc_hd__mux2_1
Xfanout108 _1589_/Q VGND VGND VPWR VPWR _1335_/A sky130_fd_sc_hd__buf_2
Xfanout119 input2/X VGND VGND VPWR VPWR fanout119/X sky130_fd_sc_hd__buf_2
X_1465_ _1258_/A _1464_/X _1217_/Y _1216_/X VGND VGND VPWR VPWR _1465_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1396_ _0960_/X _1393_/X _1395_/X _0964_/Y VGND VGND VPWR VPWR _1396_/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1250_ _1248_/X _1249_/X _1565_/B VGND VGND VPWR VPWR _1251_/C sky130_fd_sc_hd__o21ai_1
X_1181_ _1181_/A _1181_/B _1181_/C _1181_/D VGND VGND VPWR VPWR _1181_/X sky130_fd_sc_hd__or4_1
XFILLER_0_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0896_ _1339_/B _1454_/B VGND VGND VPWR VPWR _1434_/A sky130_fd_sc_hd__nor2_2
X_0965_ _1339_/B _1237_/A _1352_/A VGND VGND VPWR VPWR _0965_/X sky130_fd_sc_hd__and3_1
X_1517_ hold11/A _1518_/B VGND VGND VPWR VPWR _1517_/Y sky130_fd_sc_hd__nand2_1
X_1448_ _1347_/X _1447_/X _1600_/Q VGND VGND VPWR VPWR _1448_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1379_ _1005_/X _1378_/X _0952_/B _0947_/Y VGND VGND VPWR VPWR _1379_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap8 _1039_/B VGND VGND VPWR VPWR _1256_/B sky130_fd_sc_hd__clkbuf_2
Xfanout90 fanout91/X VGND VGND VPWR VPWR _1539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1302_ _0887_/A _0932_/Y _1212_/X _1301_/X _1598_/Q VGND VGND VPWR VPWR _1302_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1233_ _1405_/B _1233_/B VGND VGND VPWR VPWR _1233_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1164_ _1190_/B _1164_/B _1164_/C VGND VGND VPWR VPWR _1164_/X sky130_fd_sc_hd__and3_1
X_1095_ _1100_/A _0849_/B _1362_/B VGND VGND VPWR VPWR _1300_/D sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0948_ _0930_/D _1252_/C _1408_/C _1370_/A _1252_/A _1212_/A VGND VGND VPWR VPWR
+ _0948_/X sky130_fd_sc_hd__mux4_1
X_0879_ _1225_/A _1247_/B VGND VGND VPWR VPWR _0887_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0802_ _1525_/B hold4/X VGND VGND VPWR VPWR _1604_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1216_ _1436_/A _1439_/B _1015_/B _1036_/A VGND VGND VPWR VPWR _1216_/X sky130_fd_sc_hd__a211o_1
X_1147_ _1236_/C _1147_/B VGND VGND VPWR VPWR _1436_/A sky130_fd_sc_hd__nand2_2
X_1078_ _1286_/C _1181_/B VGND VGND VPWR VPWR _1078_/X sky130_fd_sc_hd__or2_1
XFILLER_0_1_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _1398_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1001_ _1405_/A _1001_/B VGND VGND VPWR VPWR _1001_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1550_ _1442_/A _0991_/X _1562_/B _1547_/Y _1181_/A VGND VGND VPWR VPWR _1595_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1481_ _1361_/A _1025_/A _1300_/A _1114_/C _1480_/Y VGND VGND VPWR VPWR _1481_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_27_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ _1199_/C _1094_/A _1335_/A _0991_/A _0932_/A VGND VGND VPWR VPWR _1339_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1602_ clkload1/A _1602_/D fanout117/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1533_ _1533_/A _1542_/B VGND VGND VPWR VPWR _1533_/Y sky130_fd_sc_hd__nor2_1
Xfanout109 _1200_/A1 VGND VGND VPWR VPWR _1072_/B sky130_fd_sc_hd__buf_4
XFILLER_0_22_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1395_ _0966_/X _1394_/X _1225_/A VGND VGND VPWR VPWR _1395_/X sky130_fd_sc_hd__a21o_1
X_1464_ _0869_/A _1237_/A _0936_/Y _1218_/Y _1463_/X VGND VGND VPWR VPWR _1464_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1180_ _1180_/A _1180_/B VGND VGND VPWR VPWR _1180_/Y sky130_fd_sc_hd__nand2_1
X_0964_ _0961_/X _0963_/X _1066_/A VGND VGND VPWR VPWR _0964_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1516_ _1516_/A1 _1514_/Y _1515_/X _1524_/B hold8/X VGND VGND VPWR VPWR _1581_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0895_ _1066_/A _1015_/B VGND VGND VPWR VPWR _1454_/B sky130_fd_sc_hd__or2_4
X_1447_ _1438_/X _1446_/Y _1369_/X VGND VGND VPWR VPWR _1447_/X sky130_fd_sc_hd__a21bo_1
X_1378_ _1378_/A1 _0923_/B _1074_/B _0926_/A VGND VGND VPWR VPWR _1378_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap9 _1259_/B VGND VGND VPWR VPWR _1252_/C sky130_fd_sc_hd__buf_1
Xfanout91 _1591_/Q VGND VGND VPWR VPWR fanout91/X sky130_fd_sc_hd__clkbuf_2
Xfanout80 _1378_/A1 VGND VGND VPWR VPWR _0930_/B sky130_fd_sc_hd__buf_4
XFILLER_0_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1232_ _1323_/A _1228_/X _1230_/X _1231_/Y VGND VGND VPWR VPWR _1232_/X sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_0_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1301_ _1398_/A _1298_/Y _1300_/X _0869_/B VGND VGND VPWR VPWR _1301_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1094_ _1094_/A _1131_/B VGND VGND VPWR VPWR _1181_/D sky130_fd_sc_hd__and2_1
X_1163_ _1029_/B _1110_/Y _1162_/Y _1205_/B _1318_/A VGND VGND VPWR VPWR _1164_/C
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_30_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0947_ _1548_/B _1260_/C VGND VGND VPWR VPWR _0947_/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ _1555_/A _1190_/B VGND VGND VPWR VPWR _0878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clkload0/A VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ _1607_/Q VGND VGND VPWR VPWR _0801_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1146_ _1195_/B _1146_/B VGND VGND VPWR VPWR _1146_/X sky130_fd_sc_hd__or2_1
X_1215_ _1074_/B _1029_/B _1408_/C VGND VGND VPWR VPWR _1439_/B sky130_fd_sc_hd__a21o_1
X_1077_ _0989_/A _0937_/X _1074_/X _1357_/B _0962_/C VGND VGND VPWR VPWR _1077_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 _1593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1000_ _1420_/A _1475_/C VGND VGND VPWR VPWR _1197_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1129_ _1483_/C _1123_/X _1125_/X _1128_/X VGND VGND VPWR VPWR _1129_/X sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _1036_/B _1256_/Y _1135_/X VGND VGND VPWR VPWR _1480_/Y sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _1256_/A _1450_/A VGND VGND VPWR VPWR _0980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1601_ clkload1/A _1601_/D fanout120/X VGND VGND VPWR VPWR _1601_/Q sky130_fd_sc_hd__dfrtp_2
X_1532_ hold10/A input1/X VGND VGND VPWR VPWR _1542_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1394_ _1394_/A _1394_/B _1394_/C VGND VGND VPWR VPWR _1394_/X sky130_fd_sc_hd__or3_1
X_1463_ _1393_/A _1025_/B _1317_/B VGND VGND VPWR VPWR _1463_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_audio_player_140 VGND VGND VPWR VPWR tt_um_audio_player_140/HI uo_out[4] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_11_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0963_ _1074_/A _1074_/C _0963_/C VGND VGND VPWR VPWR _0963_/X sky130_fd_sc_hd__or3_1
X_0894_ _1066_/A _1015_/B VGND VGND VPWR VPWR _1352_/A sky130_fd_sc_hd__nor2_2
X_1515_ _1580_/Q _1513_/C hold8/A VGND VGND VPWR VPWR _1515_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1446_ _1190_/A _1440_/X _1444_/X _1445_/Y _1166_/A VGND VGND VPWR VPWR _1446_/Y
+ sky130_fd_sc_hd__a41oi_2
X_1377_ _1162_/B _1394_/B _1483_/C _1475_/D _0903_/A VGND VGND VPWR VPWR _1377_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout81 _1378_/A1 VGND VGND VPWR VPWR _0814_/B sky130_fd_sc_hd__clkbuf_2
Xfanout70 _0889_/A VGND VGND VPWR VPWR _0930_/D sky130_fd_sc_hd__clkbuf_4
Xfanout92 _1118_/A VGND VGND VPWR VPWR _0873_/A sky130_fd_sc_hd__buf_4
XFILLER_0_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1231_ _1323_/A _0988_/X _0870_/Y VGND VGND VPWR VPWR _1231_/Y sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1162_ _1370_/A _1162_/B VGND VGND VPWR VPWR _1162_/Y sky130_fd_sc_hd__nor2_1
X_1300_ _1300_/A _1300_/B _1362_/C _1300_/D VGND VGND VPWR VPWR _1300_/X sky130_fd_sc_hd__or4_1
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1093_ _1199_/C _1534_/S _1335_/A VGND VGND VPWR VPWR _1131_/B sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_22_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0877_ _1281_/B _0877_/B VGND VGND VPWR VPWR _0877_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0946_ _1408_/C VGND VGND VPWR VPWR _1320_/B sky130_fd_sc_hd__inv_2
X_1429_ _1010_/Y _1426_/X _1428_/Y _1070_/Y VGND VGND VPWR VPWR _1429_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload1 clkload1/A VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0800_ _1010_/B VGND VGND VPWR VPWR _0800_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1214_ _1207_/X _1210_/Y _1213_/X _1560_/A VGND VGND VPWR VPWR _1214_/X sky130_fd_sc_hd__a31o_1
X_1145_ _1015_/B _0921_/Y _0883_/Y VGND VGND VPWR VPWR _1145_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1076_ wire10/X _1233_/B VGND VGND VPWR VPWR _1076_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0929_ _0931_/A _0931_/B _1100_/B VGND VGND VPWR VPWR _1405_/C sky130_fd_sc_hd__or3_4
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1059_ _0926_/A _0962_/B _1036_/A VGND VGND VPWR VPWR _1450_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1128_ _0996_/A _1013_/B _1202_/B _1127_/X _1454_/B VGND VGND VPWR VPWR _1128_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1600_ clkload1/A _1600_/D fanout120/X VGND VGND VPWR VPWR _1600_/Q sky130_fd_sc_hd__dfrtp_4
X_1531_ hold10/A input1/X VGND VGND VPWR VPWR _1560_/B sky130_fd_sc_hd__and2_2
XFILLER_0_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1462_ _1462_/A _1462_/B _1462_/C VGND VGND VPWR VPWR _1462_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1393_ _1393_/A _1393_/B _1411_/C VGND VGND VPWR VPWR _1393_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtt_um_audio_player_130 VGND VGND VPWR VPWR tt_um_audio_player_130/HI uio_out[1] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_141 VGND VGND VPWR VPWR tt_um_audio_player_141/HI uo_out[5] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_36_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0962_ _0989_/A _0962_/B _0962_/C VGND VGND VPWR VPWR _0963_/C sky130_fd_sc_hd__or3_1
X_0893_ _1025_/A _1015_/B VGND VGND VPWR VPWR _1021_/B sky130_fd_sc_hd__or2_1
X_1514_ _1518_/B VGND VGND VPWR VPWR _1514_/Y sky130_fd_sc_hd__inv_2
X_1445_ _0952_/B _1443_/X _1382_/X _1010_/A VGND VGND VPWR VPWR _1445_/Y sky130_fd_sc_hd__o211ai_1
X_1376_ _1010_/A _0962_/C _1411_/C _1057_/B _1597_/Q VGND VGND VPWR VPWR _1376_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout60 _1087_/A2 VGND VGND VPWR VPWR _1443_/S sky130_fd_sc_hd__clkbuf_2
Xfanout93 _0816_/A VGND VGND VPWR VPWR _1118_/A sky130_fd_sc_hd__buf_4
Xfanout82 _0816_/B VGND VGND VPWR VPWR _1378_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout71 _0889_/A VGND VGND VPWR VPWR _1471_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1092_ _0943_/X _0993_/X _1091_/X _0789_/Y VGND VGND VPWR VPWR _1176_/B sky130_fd_sc_hd__o211a_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1161_ _1342_/A _1233_/B _0962_/C VGND VGND VPWR VPWR _1164_/B sky130_fd_sc_hd__a21o_1
X_1230_ _0848_/X _1405_/B _1420_/D _1304_/A1 VGND VGND VPWR VPWR _1230_/X sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0876_ _1281_/B _1205_/A VGND VGND VPWR VPWR _0876_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0945_ _0873_/A _0930_/B _1072_/B _1118_/B _1117_/B VGND VGND VPWR VPWR _1408_/C
+ sky130_fd_sc_hd__a41o_4
X_1428_ _1428_/A _1428_/B VGND VGND VPWR VPWR _1428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1359_ _1015_/B _1483_/A _1442_/A _1357_/Y _1358_/X VGND VGND VPWR VPWR _1359_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload2 clkload2/A VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1213_ _1454_/B _1048_/Y _1212_/X _1211_/X _1111_/B VGND VGND VPWR VPWR _1213_/X
+ sky130_fd_sc_hd__o32a_1
X_1075_ _1075_/A _1260_/C VGND VGND VPWR VPWR _1357_/B sky130_fd_sc_hd__nor2_1
X_1144_ _1166_/A _1137_/X _1139_/X _1140_/X _1143_/X VGND VGND VPWR VPWR _1144_/Y
+ sky130_fd_sc_hd__a32oi_1
XFILLER_0_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0859_ _1236_/C _1548_/B _0858_/B _1394_/A VGND VGND VPWR VPWR _0859_/X sky130_fd_sc_hd__a211o_1
X_0928_ _1199_/D _0928_/B _1252_/A VGND VGND VPWR VPWR _1135_/B sky130_fd_sc_hd__or3_2
Xhold14 hold4/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1058_ _1399_/A _1055_/X _1057_/B _0952_/B fanout6/X VGND VGND VPWR VPWR _1071_/B
+ sky130_fd_sc_hd__o221a_1
X_1127_ _0816_/A _1085_/Y _1362_/C _1300_/B _0816_/B VGND VGND VPWR VPWR _1127_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1392_ _1176_/X _1391_/X _0808_/X VGND VGND VPWR VPWR _1392_/Y sky130_fd_sc_hd__a21oi_1
X_1530_ _1181_/A _1527_/X _1529_/X hold7/A VGND VGND VPWR VPWR _1533_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1461_ _1526_/D _0889_/A _0861_/X _1099_/X VGND VGND VPWR VPWR _1462_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtt_um_audio_player_131 VGND VGND VPWR VPWR tt_um_audio_player_131/HI uio_out[2] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_142 VGND VGND VPWR VPWR tt_um_audio_player_142/HI uo_out[6] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_36_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0961_ _0818_/Y _0827_/X _0883_/Y VGND VGND VPWR VPWR _0961_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0892_ _1057_/A _1181_/A VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__nor2_4
X_1513_ hold8/A _1580_/Q _1513_/C VGND VGND VPWR VPWR _1518_/B sky130_fd_sc_hd__and3_1
X_1444_ _0955_/X _1386_/Y _1442_/Y _1596_/Q VGND VGND VPWR VPWR _1444_/X sky130_fd_sc_hd__a31o_1
X_1375_ _1352_/A _1371_/X _1374_/X _1010_/A VGND VGND VPWR VPWR _1375_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_0_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout61 _1087_/A2 VGND VGND VPWR VPWR _1111_/A sky130_fd_sc_hd__clkbuf_4
Xfanout83 _1591_/Q VGND VGND VPWR VPWR _0816_/B sky130_fd_sc_hd__clkbuf_4
Xfanout94 _1590_/Q VGND VGND VPWR VPWR _0816_/A sky130_fd_sc_hd__clkbuf_4
Xfanout72 _1420_/A VGND VGND VPWR VPWR _0926_/A sky130_fd_sc_hd__clkbuf_4
Xfanout50 _1367_/A1 VGND VGND VPWR VPWR _1317_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1091_ _1424_/A _1023_/X _1052_/X _1090_/X VGND VGND VPWR VPWR _1091_/X sky130_fd_sc_hd__a31o_1
X_1160_ _1111_/A _1319_/B _1073_/Y _1021_/B _1548_/A VGND VGND VPWR VPWR _1160_/X
+ sky130_fd_sc_hd__a311o_1
X_0944_ _1420_/A _0952_/B VGND VGND VPWR VPWR _0944_/Y sky130_fd_sc_hd__nand2_1
X_0875_ _0931_/A _1084_/B _1100_/B VGND VGND VPWR VPWR _1074_/C sky130_fd_sc_hd__nor3_4
XFILLER_0_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1427_ _1548_/B wire10/X _1544_/A _1450_/B VGND VGND VPWR VPWR _1428_/B sky130_fd_sc_hd__or4_1
X_1358_ _1281_/B _1335_/B _1015_/B _1394_/B VGND VGND VPWR VPWR _1358_/X sky130_fd_sc_hd__o211a_1
X_1289_ _0955_/B _1411_/C _1286_/X _1287_/Y _1288_/Y VGND VGND VPWR VPWR _1289_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1212_ _1212_/A _1212_/B VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1143_ _1419_/A _1141_/Y _1142_/Y _1136_/X _1424_/A VGND VGND VPWR VPWR _1143_/X
+ sky130_fd_sc_hd__o221a_1
X_1074_ _1074_/A _1074_/B _1074_/C _1074_/D VGND VGND VPWR VPWR _1074_/X sky130_fd_sc_hd__or4_1
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0927_ _1199_/D _1252_/A VGND VGND VPWR VPWR _0995_/B sky130_fd_sc_hd__nor2_1
X_0789_ _1600_/Q VGND VGND VPWR VPWR _0789_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0858_ _1394_/A _0858_/B VGND VGND VPWR VPWR _0903_/A sky130_fd_sc_hd__or2_2
XFILLER_0_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ _0888_/B _1233_/B _0996_/A VGND VGND VPWR VPWR _1202_/B sky130_fd_sc_hd__a21oi_1
X_1057_ _1057_/A _1057_/B VGND VGND VPWR VPWR _1057_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_17_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1109_ _1111_/A _1025_/Y _0975_/Y VGND VGND VPWR VPWR _1109_/X sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ _1600_/Q _1278_/Y _1347_/X _1390_/Y _1601_/Q VGND VGND VPWR VPWR _1391_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1460_ _1460_/A _1460_/B _0958_/X VGND VGND VPWR VPWR _1462_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1589_ clkload2/A _1589_/D fanout118/X VGND VGND VPWR VPWR _1589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtt_um_audio_player_132 VGND VGND VPWR VPWR tt_um_audio_player_132/HI uio_out[3] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_121 VGND VGND VPWR VPWR tt_um_audio_player_121/HI uio_oe[0] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xtt_um_audio_player_143 VGND VGND VPWR VPWR tt_um_audio_player_143/HI uo_out[7] sky130_fd_sc_hd__conb_1
XFILLER_0_8_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0960_ _1393_/B _0959_/X _1526_/D VGND VGND VPWR VPWR _0960_/X sky130_fd_sc_hd__o21a_1
X_1512_ _1516_/A1 _1510_/X _1511_/Y _1524_/B _1580_/Q VGND VGND VPWR VPWR _1580_/D
+ sky130_fd_sc_hd__a32o_1
X_0891_ _1420_/A _1286_/C _1063_/A VGND VGND VPWR VPWR _0891_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1443_ _0922_/Y _1001_/Y _1443_/S VGND VGND VPWR VPWR _1443_/X sky130_fd_sc_hd__mux2_1
X_1374_ _1180_/A _1054_/Y _1063_/Y _1373_/Y VGND VGND VPWR VPWR _1374_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout40 _1010_/A VGND VGND VPWR VPWR _1066_/A sky130_fd_sc_hd__clkbuf_4
Xfanout73 _0889_/A VGND VGND VPWR VPWR _1420_/A sky130_fd_sc_hd__buf_2
Xfanout51 _1367_/A1 VGND VGND VPWR VPWR _0952_/B sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 _1087_/A2 VGND VGND VPWR VPWR _1218_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout95 _1362_/A VGND VGND VPWR VPWR _0931_/A sky130_fd_sc_hd__buf_4
Xfanout84 fanout91/X VGND VGND VPWR VPWR _1199_/D sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1090_ _1071_/X _1089_/A _1089_/B _1599_/Q VGND VGND VPWR VPWR _1090_/X sky130_fd_sc_hd__a31o_1
X_0943_ _1424_/A _0898_/X _0942_/Y _1563_/S VGND VGND VPWR VPWR _0943_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0874_ _1199_/C _1534_/S VGND VGND VPWR VPWR _1195_/B sky130_fd_sc_hd__or2_2
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1357_ _1357_/A _1357_/B VGND VGND VPWR VPWR _1357_/Y sky130_fd_sc_hd__nand2_1
X_1426_ _0952_/B _1425_/X _1398_/C _0975_/Y VGND VGND VPWR VPWR _1426_/X sky130_fd_sc_hd__o2bb2a_1
X_1288_ _1184_/A _0953_/A _0985_/B _0854_/X VGND VGND VPWR VPWR _1288_/Y sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_21_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1211_ _1211_/A _1475_/D _0827_/X VGND VGND VPWR VPWR _1211_/X sky130_fd_sc_hd__or3b_1
X_1142_ _1010_/Y _1135_/X _1134_/X _1419_/A VGND VGND VPWR VPWR _1142_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1073_ _1074_/B _1074_/D VGND VGND VPWR VPWR _1073_/Y sky130_fd_sc_hd__nor2_1
X_0926_ _0926_/A _1443_/S VGND VGND VPWR VPWR _1260_/C sky130_fd_sc_hd__or2_4
XFILLER_0_15_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0857_ _0931_/A _1100_/A _0849_/B _1035_/A _0931_/B VGND VGND VPWR VPWR _0858_/B
+ sky130_fd_sc_hd__a311oi_4
X_0788_ _1601_/Q VGND VGND VPWR VPWR _1176_/A sky130_fd_sc_hd__inv_2
X_1409_ _1036_/A _0908_/Y _1036_/B _1037_/X _1408_/X VGND VGND VPWR VPWR _1409_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1125_ _0814_/B _0923_/B _0888_/B VGND VGND VPWR VPWR _1125_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ _1063_/A _1056_/B VGND VGND VPWR VPWR _1057_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0909_ _1420_/A _1075_/A VGND VGND VPWR VPWR _1116_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1108_ _0862_/Y _0936_/Y _1063_/Y VGND VGND VPWR VPWR _1108_/X sky130_fd_sc_hd__o21a_1
X_1039_ _1039_/A _1039_/B VGND VGND VPWR VPWR _1039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1390_ _1369_/X _1389_/X _1600_/Q VGND VGND VPWR VPWR _1390_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1588_ clkload2/A _1588_/D fanout118/X VGND VGND VPWR VPWR _1588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_audio_player_133 VGND VGND VPWR VPWR tt_um_audio_player_133/HI uio_out[4] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_122 VGND VGND VPWR VPWR tt_um_audio_player_122/HI uio_oe[1] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload0/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0890_ _1218_/A1 _1260_/A _0861_/X _0877_/Y _0889_/Y VGND VGND VPWR VPWR _0890_/X
+ sky130_fd_sc_hd__a32o_1
X_1511_ _1580_/Q _1513_/C VGND VGND VPWR VPWR _1511_/Y sky130_fd_sc_hd__nand2_1
X_1442_ _1442_/A _1442_/B VGND VGND VPWR VPWR _1442_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1373_ _0877_/Y _1399_/B _1281_/C VGND VGND VPWR VPWR _1373_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout63 _1593_/Q VGND VGND VPWR VPWR _1087_/A2 sky130_fd_sc_hd__buf_2
Xfanout85 fanout91/X VGND VGND VPWR VPWR _1094_/A sky130_fd_sc_hd__buf_1
Xfanout52 _1367_/A1 VGND VGND VPWR VPWR _1452_/A sky130_fd_sc_hd__clkbuf_2
Xfanout41 _1596_/Q VGND VGND VPWR VPWR _1010_/A sky130_fd_sc_hd__clkbuf_4
Xfanout96 _1362_/A VGND VGND VPWR VPWR _0836_/A sky130_fd_sc_hd__buf_1
Xfanout30 _1211_/A VGND VGND VPWR VPWR _1394_/A sky130_fd_sc_hd__clkbuf_4
Xfanout74 _1035_/A VGND VGND VPWR VPWR _0953_/A sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0942_ _0920_/Y _0941_/X _1560_/A VGND VGND VPWR VPWR _0942_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0873_ _0873_/A _0930_/B _1117_/B VGND VGND VPWR VPWR _1205_/A sky130_fd_sc_hd__nor3_2
X_1425_ _1075_/A _0980_/Y _1055_/X VGND VGND VPWR VPWR _1425_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ _0851_/A _1384_/A _1236_/D VGND VGND VPWR VPWR _1287_/Y sky130_fd_sc_hd__a21oi_1
X_1356_ _1419_/A _1356_/B _1356_/C _1356_/D VGND VGND VPWR VPWR _1356_/X sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_21_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1210_ _1210_/A _1210_/B VGND VGND VPWR VPWR _1210_/Y sky130_fd_sc_hd__nand2_1
X_1141_ _1352_/A _1115_/X _1116_/X VGND VGND VPWR VPWR _1141_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1072_ _0930_/B _1072_/B VGND VGND VPWR VPWR _1074_/D sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_23_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0787_ input1/X VGND VGND VPWR VPWR _0787_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0925_ _1117_/B _1256_/A VGND VGND VPWR VPWR _1233_/B sky130_fd_sc_hd__nor2_2
X_0856_ _0873_/A _1072_/B _1118_/B _0930_/B VGND VGND VPWR VPWR _0888_/B sky130_fd_sc_hd__a31oi_4
XFILLER_0_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1408_ _1483_/A wire10/A _1408_/C VGND VGND VPWR VPWR _1408_/X sky130_fd_sc_hd__or3_1
X_1339_ _1361_/A _1339_/B _1339_/C _1339_/D VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__or4_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1055_ _0827_/X _1119_/A _1063_/B _0989_/A VGND VGND VPWR VPWR _1055_/X sky130_fd_sc_hd__o211a_1
X_1124_ _1362_/B _1300_/B VGND VGND VPWR VPWR _1124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0839_ _1118_/A _0913_/A2 _1420_/A _1378_/A1 VGND VGND VPWR VPWR _1037_/A sky130_fd_sc_hd__o211a_2
X_0908_ _1074_/A wire10/X VGND VGND VPWR VPWR _0908_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1107_ _0885_/C _1180_/A _1247_/B VGND VGND VPWR VPWR _1107_/Y sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ _1454_/B _1038_/B _1038_/C _1037_/X VGND VGND VPWR VPWR _1038_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1587_ clkload1/A _1587_/D fanout117/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_audio_player_134 VGND VGND VPWR VPWR tt_um_audio_player_134/HI uio_out[5] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_123 VGND VGND VPWR VPWR tt_um_audio_player_123/HI uio_oe[2] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1441_ _1420_/A _1475_/A _1548_/B _1037_/A _1111_/A VGND VGND VPWR VPWR _1442_/B
+ sky130_fd_sc_hd__a2111o_1
X_1510_ _1580_/Q _1513_/C VGND VGND VPWR VPWR _1510_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1372_ _1548_/A _1286_/C _1434_/C _1420_/C VGND VGND VPWR VPWR _1399_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout42 _1596_/Q VGND VGND VPWR VPWR _1526_/D sky130_fd_sc_hd__clkbuf_4
Xfanout20 _0828_/X VGND VGND VPWR VPWR _1551_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout86 _1106_/A VGND VGND VPWR VPWR _1362_/B sky130_fd_sc_hd__buf_2
Xfanout53 _1135_/A VGND VGND VPWR VPWR _1114_/A sky130_fd_sc_hd__buf_2
Xfanout97 _0900_/A VGND VGND VPWR VPWR _1362_/A sky130_fd_sc_hd__clkbuf_4
Xfanout75 _0928_/B VGND VGND VPWR VPWR _1035_/A sky130_fd_sc_hd__clkbuf_4
Xfanout64 _1398_/A VGND VGND VPWR VPWR _1252_/A sky130_fd_sc_hd__buf_2
XFILLER_0_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout31 _1304_/A1 VGND VGND VPWR VPWR _1074_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ _1112_/A _1452_/C _0939_/Y _0935_/X _1010_/A VGND VGND VPWR VPWR _0941_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0872_ _0900_/C _1236_/B VGND VGND VPWR VPWR _1357_/A sky130_fd_sc_hd__or2_2
XFILLER_0_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1424_ _1424_/A _1424_/B _1424_/C VGND VGND VPWR VPWR _1424_/X sky130_fd_sc_hd__and3_1
X_1355_ _1116_/C _1348_/X _1354_/X _1010_/Y VGND VGND VPWR VPWR _1356_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_2_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1286_ _1405_/A _1420_/C _1286_/C VGND VGND VPWR VPWR _1286_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1071_ _1190_/A _1071_/B _1428_/A _1071_/D VGND VGND VPWR VPWR _1071_/X sky130_fd_sc_hd__or4_1
X_1140_ _1112_/X _1113_/X _0887_/A VGND VGND VPWR VPWR _1140_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0924_ _1361_/A _1074_/A _1037_/A _1195_/B _1218_/A1 VGND VGND VPWR VPWR _0924_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0855_ _0851_/A _0900_/C _1236_/B _1236_/D VGND VGND VPWR VPWR _1286_/C sky130_fd_sc_hd__a31o_2
XFILLER_0_11_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1338_ _1131_/B _1394_/A _1361_/A VGND VGND VPWR VPWR _1338_/X sky130_fd_sc_hd__and3b_1
X_1407_ _1032_/X _1406_/X fanout6/X VGND VGND VPWR VPWR _1415_/A sky130_fd_sc_hd__o21a_1
X_1269_ _1304_/A1 _1323_/A _1420_/C _1212_/A VGND VGND VPWR VPWR _1269_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1123_ _1236_/D _1361_/B _1181_/B _1544_/A _1057_/A VGND VGND VPWR VPWR _1123_/X
+ sky130_fd_sc_hd__o32a_1
X_1054_ _1054_/A VGND VGND VPWR VPWR _1054_/Y sky130_fd_sc_hd__inv_2
X_0907_ _1200_/A1 _0913_/A2 _1118_/A _1378_/A1 VGND VGND VPWR VPWR _1075_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0838_ _0851_/A _1236_/B _1236_/D VGND VGND VPWR VPWR _1420_/C sky130_fd_sc_hd__o21ai_4
XFILLER_0_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1106_ _1106_/A _1323_/B _1300_/B _1181_/B VGND VGND VPWR VPWR _1106_/X sky130_fd_sc_hd__or4_1
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1037_ _1037_/A _1037_/B _1056_/B VGND VGND VPWR VPWR _1037_/X sky130_fd_sc_hd__or3_1
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1586_ _1597_/CLK _1586_/D fanout117/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_audio_player_135 VGND VGND VPWR VPWR tt_um_audio_player_135/HI uio_out[6] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_124 VGND VGND VPWR VPWR tt_um_audio_player_124/HI uio_oe[3] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_36_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1440_ _1379_/X _1439_/Y _1010_/Y VGND VGND VPWR VPWR _1440_/X sky130_fd_sc_hd__a21o_1
X_1371_ _1260_/A _1420_/B _0862_/Y _1318_/B _1370_/Y VGND VGND VPWR VPWR _1371_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1569_ _1176_/A _1562_/B _1565_/X _1568_/X VGND VGND VPWR VPWR _1601_/D sky130_fd_sc_hd__a31o_1
Xfanout21 _1294_/A VGND VGND VPWR VPWR _1036_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout98 _0900_/A VGND VGND VPWR VPWR _0851_/A sky130_fd_sc_hd__buf_4
Xfanout43 _1596_/Q VGND VGND VPWR VPWR _1247_/B sky130_fd_sc_hd__clkbuf_2
Xfanout65 _0932_/A VGND VGND VPWR VPWR _1398_/A sky130_fd_sc_hd__buf_2
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout32 _1304_/A1 VGND VGND VPWR VPWR _1405_/A sky130_fd_sc_hd__clkbuf_4
Xfanout87 _1106_/A VGND VGND VPWR VPWR _0931_/B sky130_fd_sc_hd__buf_4
Xfanout76 _0889_/A VGND VGND VPWR VPWR _0928_/B sky130_fd_sc_hd__buf_2
Xfanout54 _1367_/A1 VGND VGND VPWR VPWR _1135_/A sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0940_ _1548_/A _1420_/D VGND VGND VPWR VPWR _0940_/Y sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_30_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0871_ _1100_/A _1100_/B VGND VGND VPWR VPWR _1281_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1285_ _1282_/X _1284_/Y _1526_/D VGND VGND VPWR VPWR _1285_/Y sky130_fd_sc_hd__a21oi_1
X_1423_ _1423_/A _1423_/B _1423_/C _1423_/D VGND VGND VPWR VPWR _1424_/C sky130_fd_sc_hd__or4_1
X_1354_ _0936_/Y _0975_/Y _1353_/X VGND VGND VPWR VPWR _1354_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1070_ _1190_/A _1071_/D VGND VGND VPWR VPWR _1070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0923_ _1111_/B _0923_/B VGND VGND VPWR VPWR _0923_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0854_ _1362_/B _1084_/B VGND VGND VPWR VPWR _0854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1337_ _1333_/Y _1334_/Y _1336_/X _1210_/A VGND VGND VPWR VPWR _1345_/A sky130_fd_sc_hd__o31a_1
X_1406_ _0922_/Y _1405_/X _1267_/A VGND VGND VPWR VPWR _1406_/X sky130_fd_sc_hd__o21a_1
X_1268_ _1266_/X _1267_/Y _1116_/C VGND VGND VPWR VPWR _1268_/Y sky130_fd_sc_hd__a21oi_1
X_1199_ _1335_/A _0928_/B _1199_/C _1199_/D VGND VGND VPWR VPWR _1283_/C sky130_fd_sc_hd__and4bb_1
XFILLER_0_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ _1236_/D _1361_/B VGND VGND VPWR VPWR _1342_/B sky130_fd_sc_hd__nor2_1
X_1053_ _0827_/X _1119_/A _1398_/A VGND VGND VPWR VPWR _1054_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0837_ _1362_/A _0849_/B _1199_/D VGND VGND VPWR VPWR _1035_/B sky130_fd_sc_hd__o21a_1
X_0906_ _1072_/B _1118_/B _0873_/A _0930_/B VGND VGND VPWR VPWR wire10/A sky130_fd_sc_hd__a211oi_1
XFILLER_0_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1105_ _1114_/A _1237_/A _0940_/Y _1104_/X VGND VGND VPWR VPWR _1105_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1036_ _1036_/A _1036_/B VGND VGND VPWR VPWR _1038_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1585_ _1597_/CLK _1585_/D fanout117/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1019_ _1074_/B _1038_/B _1018_/Y _1210_/A VGND VGND VPWR VPWR _1419_/B sky130_fd_sc_hd__o211a_1
Xtt_um_audio_player_136 VGND VGND VPWR VPWR tt_um_audio_player_136/HI uio_out[7] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_125 VGND VGND VPWR VPWR tt_um_audio_player_125/HI uio_oe[4] sky130_fd_sc_hd__conb_1
XFILLER_0_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1370_ _1370_/A _1450_/A VGND VGND VPWR VPWR _1370_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1499_ _1516_/A1 _1525_/B _1576_/Q VGND VGND VPWR VPWR _1576_/D sky130_fd_sc_hd__mux2_1
X_1568_ _1601_/Q _1568_/B VGND VGND VPWR VPWR _1568_/X sky130_fd_sc_hd__and2_1
Xfanout55 _1367_/A1 VGND VGND VPWR VPWR _1339_/B sky130_fd_sc_hd__clkbuf_4
Xfanout44 _1010_/B VGND VGND VPWR VPWR _1015_/B sky130_fd_sc_hd__clkbuf_4
Xfanout22 _0811_/X VGND VGND VPWR VPWR _1111_/B sky130_fd_sc_hd__buf_4
Xfanout33 _0797_/Y VGND VGND VPWR VPWR _1304_/A1 sky130_fd_sc_hd__buf_2
Xfanout77 _0991_/A VGND VGND VPWR VPWR _1236_/C sky130_fd_sc_hd__clkbuf_4
Xfanout99 _1199_/C VGND VGND VPWR VPWR _0900_/A sky130_fd_sc_hd__buf_2
Xfanout66 _0932_/A VGND VGND VPWR VPWR _0955_/B sky130_fd_sc_hd__buf_2
Xfanout88 fanout91/X VGND VGND VPWR VPWR _1106_/A sky130_fd_sc_hd__buf_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0870_ _1057_/A _1181_/A VGND VGND VPWR VPWR _0870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1422_ _1006_/Y _1421_/X _1352_/A VGND VGND VPWR VPWR _1423_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1353_ _1184_/A _1072_/B _1118_/B _1111_/B _1036_/A VGND VGND VPWR VPWR _1353_/X
+ sky130_fd_sc_hd__a41o_1
X_1284_ _1260_/C _1241_/Y _1283_/Y _0933_/Y _1442_/A VGND VGND VPWR VPWR _1284_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0999_ _1362_/A _1084_/B _0849_/B _1362_/B VGND VGND VPWR VPWR _1001_/B sky130_fd_sc_hd__o31ai_2
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0853_ _1405_/A _1542_/A VGND VGND VPWR VPWR _1551_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0922_ _1370_/A _1300_/B VGND VGND VPWR VPWR _0922_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1405_ _1405_/A _1405_/B _1405_/C VGND VGND VPWR VPWR _1405_/X sky130_fd_sc_hd__and3_1
XFILLER_0_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 ena VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_2
X_1336_ _0928_/B _1335_/Y _1146_/X _1205_/B VGND VGND VPWR VPWR _1336_/X sky130_fd_sc_hd__o211a_1
X_1198_ _1025_/A _0819_/X _1197_/X _1196_/X VGND VGND VPWR VPWR _1198_/X sky130_fd_sc_hd__a31o_1
X_1267_ _1267_/A _1267_/B VGND VGND VPWR VPWR _1267_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ _0962_/C _0915_/Y _1005_/X _1120_/X VGND VGND VPWR VPWR _1121_/X sky130_fd_sc_hd__a31o_1
X_1052_ _1033_/X _1038_/X _1051_/X _1190_/A VGND VGND VPWR VPWR _1052_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0905_ _1084_/B _0849_/B _1362_/A VGND VGND VPWR VPWR _1300_/B sky130_fd_sc_hd__a21oi_4
X_0836_ _0836_/A _1100_/B VGND VGND VPWR VPWR _1319_/B sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_19_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _1361_/A _1319_/B VGND VGND VPWR VPWR _1320_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1104_ _0869_/B _1102_/B _1475_/A _0962_/C VGND VGND VPWR VPWR _1104_/X sky130_fd_sc_hd__o31a_1
X_1035_ _1035_/A _1035_/B VGND VGND VPWR VPWR _1036_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ _1111_/B _1300_/A _1252_/A VGND VGND VPWR VPWR _0819_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1584_ clkload1/A _1584_/D fanout117/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_audio_player_126 VGND VGND VPWR VPWR tt_um_audio_player_126/HI uio_oe[5] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_137 VGND VGND VPWR VPWR tt_um_audio_player_137/HI uo_out[1] sky130_fd_sc_hd__conb_1
X_1018_ _1074_/B _1181_/B VGND VGND VPWR VPWR _1018_/Y sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1567_ _1567_/A _1568_/B VGND VGND VPWR VPWR _1600_/D sky130_fd_sc_hd__and2_1
X_1498_ hold10/X input1/X _1497_/Y VGND VGND VPWR VPWR _1574_/D sky130_fd_sc_hd__o21ba_1
Xfanout34 _1225_/A VGND VGND VPWR VPWR _1190_/A sky130_fd_sc_hd__clkbuf_4
Xfanout89 fanout91/X VGND VGND VPWR VPWR _1236_/D sky130_fd_sc_hd__clkbuf_4
Xfanout56 _1367_/A1 VGND VGND VPWR VPWR _1057_/A sky130_fd_sc_hd__buf_2
Xfanout78 _0889_/A VGND VGND VPWR VPWR _0991_/A sky130_fd_sc_hd__buf_2
Xfanout23 _0800_/Y VGND VGND VPWR VPWR _1258_/A sky130_fd_sc_hd__clkbuf_4
Xfanout67 _0932_/A VGND VGND VPWR VPWR _0985_/B sky130_fd_sc_hd__clkbuf_4
Xfanout12 _1460_/B VGND VGND VPWR VPWR _1281_/C sky130_fd_sc_hd__clkbuf_4
Xfanout45 _1318_/A VGND VGND VPWR VPWR _1323_/B sky130_fd_sc_hd__buf_2
XFILLER_0_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1421_ _1439_/A _0864_/B _1001_/Y _1420_/X VGND VGND VPWR VPWR _1421_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1352_ _1352_/A _1352_/B VGND VGND VPWR VPWR _1356_/C sky130_fd_sc_hd__nand2_1
X_1283_ _1534_/S _1398_/A _1283_/C VGND VGND VPWR VPWR _1283_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0998_ _0816_/A _1200_/A1 _1040_/B _0816_/B VGND VGND VPWR VPWR _1475_/C sky130_fd_sc_hd__o31a_1
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0921_ _1339_/B _1195_/A VGND VGND VPWR VPWR _0921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0852_ _0900_/A _1539_/A _0900_/C _1236_/B VGND VGND VPWR VPWR _1542_/A sky130_fd_sc_hd__nand4_4
XFILLER_0_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1404_ _1560_/A _1401_/X _1403_/X _1166_/A _1396_/X VGND VGND VPWR VPWR _1404_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_1_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1335_ _1335_/A _1335_/B VGND VGND VPWR VPWR _1335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 rst_n VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_1
X_1197_ _1197_/A _1197_/B VGND VGND VPWR VPWR _1197_/X sky130_fd_sc_hd__or2_1
X_1266_ _1111_/A _1001_/Y _1265_/X _1212_/A VGND VGND VPWR VPWR _1266_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1120_ _1066_/A _0914_/Y _1004_/Y _1119_/X VGND VGND VPWR VPWR _1120_/X sky130_fd_sc_hd__o31a_1
X_1051_ _1210_/A _1414_/B _1046_/Y _1050_/X VGND VGND VPWR VPWR _1051_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0904_ _1072_/B _1118_/B _0873_/A VGND VGND VPWR VPWR _0923_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0835_ _0953_/A _0985_/B VGND VGND VPWR VPWR _1102_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1318_ _1318_/A _1318_/B VGND VGND VPWR VPWR _1318_/Y sky130_fd_sc_hd__nor2_1
X_1249_ _1013_/B _0962_/C _1442_/A _1212_/B VGND VGND VPWR VPWR _1249_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_19_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1103_ _0903_/C _1102_/X _1281_/C VGND VGND VPWR VPWR _1103_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1034_ _1405_/A _1420_/C VGND VGND VPWR VPWR _1267_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0818_ _1111_/B _1300_/A _0989_/A VGND VGND VPWR VPWR _0818_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1583_ _1597_/CLK _1583_/D fanout118/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xtt_um_audio_player_127 VGND VGND VPWR VPWR tt_um_audio_player_127/HI uio_oe[6] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_138 VGND VGND VPWR VPWR tt_um_audio_player_138/HI uo_out[2] sky130_fd_sc_hd__conb_1
X_1017_ _1483_/A _1408_/C VGND VGND VPWR VPWR _1038_/B sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1497_ hold6/A hold5/A _1497_/C _1497_/D VGND VGND VPWR VPWR _1497_/Y sky130_fd_sc_hd__nor4_2
X_1566_ _1544_/B _1565_/X _1560_/B VGND VGND VPWR VPWR _1568_/B sky130_fd_sc_hd__o21ai_1
Xfanout35 _0790_/Y VGND VGND VPWR VPWR _1225_/A sky130_fd_sc_hd__buf_2
Xfanout79 _1592_/Q VGND VGND VPWR VPWR _0889_/A sky130_fd_sc_hd__buf_2
Xfanout24 _0800_/Y VGND VGND VPWR VPWR _0869_/B sky130_fd_sc_hd__buf_2
Xfanout57 _1594_/Q VGND VGND VPWR VPWR _1367_/A1 sky130_fd_sc_hd__buf_2
Xfanout68 _1593_/Q VGND VGND VPWR VPWR _0932_/A sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout46 _1010_/B VGND VGND VPWR VPWR _1318_/A sky130_fd_sc_hd__buf_2
XFILLER_0_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1420_ _1420_/A _1420_/B _1420_/C _1420_/D VGND VGND VPWR VPWR _1420_/X sky130_fd_sc_hd__and4_1
X_1351_ _0817_/Y _1037_/B _1350_/Y _1112_/C _0996_/A VGND VGND VPWR VPWR _1352_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1282_ _1282_/A _1282_/B _1282_/C VGND VGND VPWR VPWR _1282_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0997_ _1218_/A1 _0877_/Y _1063_/B _0996_/Y VGND VGND VPWR VPWR _0997_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1549_ _1057_/A _1548_/X _1547_/Y VGND VGND VPWR VPWR _1594_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_17_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0920_ _0920_/A _0920_/B _0920_/C VGND VGND VPWR VPWR _0920_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0851_ _0851_/A _1236_/D _0900_/C _0851_/D VGND VGND VPWR VPWR _1548_/B sky130_fd_sc_hd__and4_4
XFILLER_0_23_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1403_ _0972_/X _1015_/Y _1398_/X _1402_/Y fanout6/X VGND VGND VPWR VPWR _1403_/X
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1334_ _1334_/A _1334_/B VGND VGND VPWR VPWR _1334_/Y sky130_fd_sc_hd__nor2_1
X_1265_ _1370_/A _1265_/B VGND VGND VPWR VPWR _1265_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1196_ _1212_/A _1195_/Y _1454_/B VGND VGND VPWR VPWR _1196_/X sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _1439_/A _1411_/C _1116_/C VGND VGND VPWR VPWR _1050_/X sky130_fd_sc_hd__a21o_1
X_0903_ _0903_/A _0903_/B _0903_/C VGND VGND VPWR VPWR _0920_/A sky130_fd_sc_hd__and3_1
XFILLER_0_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0834_ _1117_/B _1111_/A VGND VGND VPWR VPWR _0933_/B sky130_fd_sc_hd__and2_2
XFILLER_0_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1248_ _0962_/B _1548_/A _1180_/A _0887_/A VGND VGND VPWR VPWR _1248_/X sky130_fd_sc_hd__a31o_1
X_1317_ _1317_/A _1317_/B VGND VGND VPWR VPWR _1318_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1260_/A _1114_/C _1135_/B VGND VGND VPWR VPWR _1180_/B sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_19_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1102_ _1539_/A _1102_/B _1309_/B VGND VGND VPWR VPWR _1102_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1033_ _1039_/A _1267_/A _1010_/Y _1032_/X VGND VGND VPWR VPWR _1033_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0817_ _1074_/A _0817_/B VGND VGND VPWR VPWR _0817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1582_ _1597_/CLK _1582_/D fanout118/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xtt_um_audio_player_128 VGND VGND VPWR VPWR tt_um_audio_player_128/HI uio_oe[7] sky130_fd_sc_hd__conb_1
Xtt_um_audio_player_139 VGND VGND VPWR VPWR tt_um_audio_player_139/HI uo_out[3] sky130_fd_sc_hd__conb_1
X_1016_ _1066_/A _1258_/A VGND VGND VPWR VPWR _1016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1496_ hold2/A hold3/A _1524_/B VGND VGND VPWR VPWR _1497_/D sky130_fd_sc_hd__or3_1
X_1565_ _1600_/Q _1565_/B _1570_/C VGND VGND VPWR VPWR _1565_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_24_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout36 _1598_/Q VGND VGND VPWR VPWR _1424_/A sky130_fd_sc_hd__clkbuf_4
Xfanout47 _1010_/B VGND VGND VPWR VPWR _1181_/A sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout58 _1087_/A2 VGND VGND VPWR VPWR _1256_/A sky130_fd_sc_hd__clkbuf_4
Xfanout14 _0870_/Y VGND VGND VPWR VPWR _0962_/C sky130_fd_sc_hd__clkbuf_4
Xfanout69 _0930_/D VGND VGND VPWR VPWR _1117_/B sky130_fd_sc_hd__buf_4
Xfanout25 _0869_/A VGND VGND VPWR VPWR _0996_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1281_ _1281_/A _1281_/B _1281_/C _1043_/B VGND VGND VPWR VPWR _1282_/C sky130_fd_sc_hd__or4b_1
X_1350_ _1475_/A _1362_/D _0988_/X VGND VGND VPWR VPWR _1350_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0996_ _0996_/A _1135_/B VGND VGND VPWR VPWR _0996_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1548_ _1548_/A _1548_/B _1560_/B VGND VGND VPWR VPWR _1548_/X sky130_fd_sc_hd__and3_1
X_1479_ _0915_/Y _1478_/Y _1317_/A VGND VGND VPWR VPWR _1479_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0850_ _1184_/A _1370_/A VGND VGND VPWR VPWR _1197_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1402_ _1063_/A _1197_/A _1394_/B _0973_/X VGND VGND VPWR VPWR _1402_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1333_ _1450_/A _1332_/X _0975_/Y VGND VGND VPWR VPWR _1333_/Y sky130_fd_sc_hd__a21oi_1
X_1264_ _1010_/A _1258_/X _1263_/X _1255_/Y VGND VGND VPWR VPWR _1277_/B sky130_fd_sc_hd__o211a_1
Xclkbuf_2_1__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload1/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1195_ _1195_/A _1195_/B VGND VGND VPWR VPWR _1195_/Y sky130_fd_sc_hd__nand2_2
X_0979_ _1548_/A _1286_/C VGND VGND VPWR VPWR _1212_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0902_ _1452_/A _0903_/C VGND VGND VPWR VPWR _0902_/Y sky130_fd_sc_hd__nand2_1
X_0833_ _0869_/A _0819_/X _1281_/A _0832_/X VGND VGND VPWR VPWR _0833_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1247_ _1560_/A _1247_/B _1247_/C _1247_/D VGND VGND VPWR VPWR _1251_/B sky130_fd_sc_hd__and4_1
X_1178_ _1304_/A1 _1475_/C _1177_/X _1218_/A1 _0962_/C VGND VGND VPWR VPWR _1178_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1316_ _1394_/A _1313_/Y _1315_/X _0885_/B VGND VGND VPWR VPWR _1316_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap11 _1147_/B VGND VGND VPWR VPWR _1342_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ _1339_/D _1101_/B VGND VGND VPWR VPWR _1309_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1032_ _1036_/A _1025_/Y _0858_/B _0819_/X VGND VGND VPWR VPWR _1032_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_16_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0816_ _0816_/A _0816_/B _1040_/B VGND VGND VPWR VPWR _0817_/B sky130_fd_sc_hd__nand3_1
X_1581_ _1597_/CLK _1581_/D fanout119/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1015_ _1190_/B _1015_/B VGND VGND VPWR VPWR _1015_/Y sky130_fd_sc_hd__nor2_2
Xtt_um_audio_player_129 VGND VGND VPWR VPWR tt_um_audio_player_129/HI uio_out[0] sky130_fd_sc_hd__conb_1
XFILLER_0_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1564_ _1565_/B _1560_/X _1600_/Q VGND VGND VPWR VPWR _1567_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1495_ _1577_/Q _1494_/X hold11/A hold13/A VGND VGND VPWR VPWR _1497_/C sky130_fd_sc_hd__o211a_1
Xfanout37 _1597_/Q VGND VGND VPWR VPWR _1419_/A sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout26 _0869_/A VGND VGND VPWR VPWR _1212_/A sky130_fd_sc_hd__clkbuf_4
Xfanout15 _1102_/B VGND VGND VPWR VPWR _1114_/C sky130_fd_sc_hd__clkbuf_4
Xfanout48 _1595_/Q VGND VGND VPWR VPWR _1010_/B sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout59 _1443_/S VGND VGND VPWR VPWR _0989_/A sky130_fd_sc_hd__buf_2
XFILLER_0_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1280_ _1339_/D _1101_/B _1539_/A _0955_/X VGND VGND VPWR VPWR _1282_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_25_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0995_ _1135_/A _0995_/B VGND VGND VPWR VPWR _0995_/Y sky130_fd_sc_hd__nor2_1
X_1547_ _1560_/B _1547_/B VGND VGND VPWR VPWR _1547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1478_ _1117_/B _1125_/X _1112_/C VGND VGND VPWR VPWR _1478_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1401_ _0990_/X _0991_/X _1400_/X _1190_/B VGND VGND VPWR VPWR _1401_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1194_ _1111_/A _1025_/Y _1193_/X VGND VGND VPWR VPWR _1194_/Y sky130_fd_sc_hd__o21ai_1
X_1332_ _1035_/B _1085_/Y _0888_/B VGND VGND VPWR VPWR _1332_/X sky130_fd_sc_hd__a21o_1
X_1263_ _0914_/Y _1261_/X _1262_/X _1259_/X VGND VGND VPWR VPWR _1263_/X sky130_fd_sc_hd__o31a_1
X_0978_ _0991_/A _1420_/D _1405_/B _1205_/B _1181_/A VGND VGND VPWR VPWR _0978_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0832_ _1420_/B _0827_/X _1551_/A _1131_/A _0869_/B VGND VGND VPWR VPWR _0832_/X
+ sky130_fd_sc_hd__a221o_1
X_0901_ _1236_/C _1420_/D _0955_/B VGND VGND VPWR VPWR _0903_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1315_ _1025_/B _1334_/B _1314_/Y _1252_/B VGND VGND VPWR VPWR _1315_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1246_ _1394_/A _0923_/Y _0962_/C VGND VGND VPWR VPWR _1247_/D sky130_fd_sc_hd__a21o_1
X_1177_ _1361_/A _1300_/A _1281_/B _1335_/B _1420_/A VGND VGND VPWR VPWR _1177_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1031_ _1025_/Y _1028_/X _1029_/Y _1181_/B _1030_/Y VGND VGND VPWR VPWR _1414_/B
+ sky130_fd_sc_hd__o221a_1
X_1100_ _1100_/A _1100_/B _0836_/A VGND VGND VPWR VPWR _1101_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0815_ _1199_/C _1094_/A _1335_/A VGND VGND VPWR VPWR _0933_/A sky130_fd_sc_hd__and3_1
XFILLER_0_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1229_ _1229_/A _1393_/A VGND VGND VPWR VPWR _1334_/B sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1597_/CLK _1580_/D fanout118/X VGND VGND VPWR VPWR _1580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1014_ _1011_/X _1013_/Y fanout6/X VGND VGND VPWR VPWR _1023_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1494_ hold9/A _1578_/Q hold8/A _1580_/Q VGND VGND VPWR VPWR _1494_/X sky130_fd_sc_hd__or4_1
X_1563_ _1559_/Y _1562_/X _1563_/S VGND VGND VPWR VPWR _1599_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout38 _1555_/A VGND VGND VPWR VPWR _1560_/A sky130_fd_sc_hd__buf_2
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout49 _1317_/A VGND VGND VPWR VPWR _1025_/A sky130_fd_sc_hd__clkbuf_4
Xfanout27 _0799_/Y VGND VGND VPWR VPWR _0869_/A sky130_fd_sc_hd__clkbuf_4
Xfanout16 _0933_/B VGND VGND VPWR VPWR _1548_/A sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0994_ _1190_/B _1015_/B VGND VGND VPWR VPWR _1116_/C sky130_fd_sc_hd__nand2_2
X_1477_ _1204_/B _1472_/X _1476_/X _1466_/X _1599_/Q VGND VGND VPWR VPWR _1489_/C
+ sky130_fd_sc_hd__a311o_1
X_1546_ _1551_/A _1551_/B _1533_/A VGND VGND VPWR VPWR _1547_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1400_ _1020_/X _1399_/Y _0978_/X VGND VGND VPWR VPWR _1400_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1331_ _0878_/Y _1327_/X _1330_/X _1598_/Q VGND VGND VPWR VPWR _1331_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1193_ _1025_/A _1452_/C _1192_/Y fanout6/X VGND VGND VPWR VPWR _1193_/X sky130_fd_sc_hd__o31a_1
X_1262_ _0888_/B _1233_/B _1454_/B VGND VGND VPWR VPWR _1262_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0977_ _1318_/A _0972_/X _0976_/Y _0878_/Y VGND VGND VPWR VPWR _0977_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1529_ hold12/A _1570_/B VGND VGND VPWR VPWR _1529_/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0900_/A _1539_/A _0900_/C _1236_/B VGND VGND VPWR VPWR _1420_/D sky130_fd_sc_hd__or4_4
XFILLER_0_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0831_ _1236_/C _1236_/D VGND VGND VPWR VPWR _1131_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ _1339_/D _1101_/B _1114_/B VGND VGND VPWR VPWR _1314_/Y sky130_fd_sc_hd__a21oi_1
X_1176_ _1176_/A _1176_/B _1176_/C VGND VGND VPWR VPWR _1176_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1245_ _1135_/A _1244_/X _1242_/X _1323_/B VGND VGND VPWR VPWR _1247_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_11 _0883_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap13 _1205_/A VGND VGND VPWR VPWR _0877_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1030_ _1087_/A2 _1256_/B _1362_/C _1548_/B _0996_/A VGND VGND VPWR VPWR _1030_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_33_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ _0873_/A _0814_/B VGND VGND VPWR VPWR _1260_/A sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_16_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1228_ _1074_/C _1227_/X _0928_/B _1542_/A VGND VGND VPWR VPWR _1228_/X sky130_fd_sc_hd__o211a_1
X_1159_ _1159_/A _1159_/B _1157_/X VGND VGND VPWR VPWR _1159_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1013_ _1025_/A _1013_/B VGND VGND VPWR VPWR _1013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1493_ _1392_/Y _1490_/Y _1492_/X VGND VGND VPWR VPWR _1608_/D sky130_fd_sc_hd__o21ba_1
X_1562_ _1598_/Q _1562_/B _1570_/C VGND VGND VPWR VPWR _1562_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout39 _1597_/Q VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 _1211_/A VGND VGND VPWR VPWR _1063_/A sky130_fd_sc_hd__clkbuf_4
Xfanout17 _0829_/Y VGND VGND VPWR VPWR _1483_/A sky130_fd_sc_hd__buf_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0993_ _0967_/X _0977_/X _0992_/X _1166_/A VGND VGND VPWR VPWR _0993_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1545_ _0955_/B _1541_/Y _1542_/Y _1544_/Y VGND VGND VPWR VPWR _1593_/D sky130_fd_sc_hd__a22o_1
X_1476_ _1182_/X _1211_/X _1474_/X _1475_/X _1190_/A VGND VGND VPWR VPWR _1476_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1261_ _1114_/C _1286_/C _1074_/C _1260_/X _1025_/A VGND VGND VPWR VPWR _1261_/X
+ sky130_fd_sc_hd__o311a_1
X_1330_ _1324_/Y _1326_/Y _1329_/X _1114_/A VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_36_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1192_ _1357_/A _1260_/C VGND VGND VPWR VPWR _1192_/Y sky130_fd_sc_hd__nor2_1
X_0976_ _1394_/B _0975_/Y _0973_/X _1318_/A VGND VGND VPWR VPWR _0976_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1528_ _1601_/Q _1600_/Q _1565_/B VGND VGND VPWR VPWR _1570_/B sky130_fd_sc_hd__and3_1
X_1459_ _1147_/B _0957_/Y _1039_/B _1323_/A VGND VGND VPWR VPWR _1460_/A sky130_fd_sc_hd__o211a_1
XFILLER_0_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ _1361_/A _0930_/D VGND VGND VPWR VPWR _1483_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1313_ _1025_/B _1334_/B _1252_/B VGND VGND VPWR VPWR _1313_/Y sky130_fd_sc_hd__a21oi_1
X_1244_ _1548_/A _1241_/Y _1243_/Y _1199_/D VGND VGND VPWR VPWR _1244_/X sky130_fd_sc_hd__a22o_1
X_1175_ _1599_/Q _1144_/Y _1153_/Y _1174_/X VGND VGND VPWR VPWR _1176_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_12 _1590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0959_ _0962_/B _1260_/C _0958_/X _0903_/B VGND VGND VPWR VPWR _0959_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0813_ _0873_/A _1118_/B VGND VGND VPWR VPWR _1300_/A sky130_fd_sc_hd__and2_2
XFILLER_0_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1227_ _0836_/A _1106_/A _1100_/A _1100_/B VGND VGND VPWR VPWR _1227_/X sky130_fd_sc_hd__o211a_1
X_1158_ _1037_/B _1146_/X _1318_/A _1162_/B VGND VGND VPWR VPWR _1159_/B sky130_fd_sc_hd__o211ai_1
X_1089_ _1089_/A _1089_/B VGND VGND VPWR VPWR _1089_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1012_ _1471_/A1 _1548_/B _1111_/A VGND VGND VPWR VPWR _1013_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1492_ _1176_/X _1391_/X _1491_/X _1525_/B VGND VGND VPWR VPWR _1492_/X sky130_fd_sc_hd__a31o_1
X_1561_ _1424_/A _1560_/X _1559_/Y VGND VGND VPWR VPWR _1598_/D sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout18 _0829_/Y VGND VGND VPWR VPWR _1162_/B sky130_fd_sc_hd__clkbuf_2
Xfanout29 _1394_/A VGND VGND VPWR VPWR _1323_/A sky130_fd_sc_hd__buf_2
XFILLER_0_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0992_ _0990_/X _0991_/X _0843_/Y _0983_/X VGND VGND VPWR VPWR _0992_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1544_ _1544_/A _1544_/B VGND VGND VPWR VPWR _1544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1475_ _1475_/A _1544_/A _1475_/C _1475_/D VGND VGND VPWR VPWR _1475_/X sky130_fd_sc_hd__or4_1
XFILLER_0_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1191_ _1189_/X _1190_/X _1424_/A VGND VGND VPWR VPWR _1204_/B sky130_fd_sc_hd__o21a_1
X_1260_ _1260_/A _1357_/A _1260_/C VGND VGND VPWR VPWR _1260_/X sky130_fd_sc_hd__or3_1
XFILLER_0_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0975_ _1317_/A _1256_/A VGND VGND VPWR VPWR _0975_/Y sky130_fd_sc_hd__nand2b_4
X_1527_ hold12/A _1488_/A _1527_/C _1601_/Q VGND VGND VPWR VPWR _1527_/X sky130_fd_sc_hd__and4bb_1
X_1389_ _1375_/Y _1376_/X _1377_/X _1388_/X VGND VGND VPWR VPWR _1389_/X sky130_fd_sc_hd__a31o_1
X_1458_ _1451_/X _1454_/X _1457_/X _1419_/A VGND VGND VPWR VPWR _1458_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_9_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1312_ _1312_/A _1312_/B _1302_/X VGND VGND VPWR VPWR _1312_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1174_ _1555_/A _1165_/X _1488_/A _1173_/Y VGND VGND VPWR VPWR _1174_/X sky130_fd_sc_hd__a211o_1
X_1243_ _1362_/C _1339_/D VGND VGND VPWR VPWR _1243_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_13 _1591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0958_ _1405_/A _1405_/B _1323_/A VGND VGND VPWR VPWR _0958_/X sky130_fd_sc_hd__a21o_1
X_0889_ _0889_/A _1286_/C VGND VGND VPWR VPWR _0889_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0812_ _0816_/B _0930_/D VGND VGND VPWR VPWR _1370_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_35_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1226_ _1166_/A _1214_/X _1225_/X _1599_/Q VGND VGND VPWR VPWR _1226_/X sky130_fd_sc_hd__a31o_1
X_1157_ _1199_/D _1300_/B _0953_/X VGND VGND VPWR VPWR _1157_/X sky130_fd_sc_hd__a21o_1
X_1088_ _0843_/Y _1083_/X _1087_/X _1424_/A VGND VGND VPWR VPWR _1089_/B sky130_fd_sc_hd__a31oi_1
XFILLER_0_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1011_ _1111_/A _1394_/C _1252_/C _0940_/Y _1367_/A1 VGND VGND VPWR VPWR _1011_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ _0869_/A _0933_/Y _1076_/Y _1208_/X _1162_/Y VGND VGND VPWR VPWR _1210_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1560_ _1560_/A _1560_/B _1560_/C VGND VGND VPWR VPWR _1560_/X sky130_fd_sc_hd__and3_1
X_1491_ _1605_/Q _1606_/Q _1607_/Q VGND VGND VPWR VPWR _1491_/X sky130_fd_sc_hd__or3_1
Xfanout19 _0828_/X VGND VGND VPWR VPWR _1439_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0991_ _0991_/A _1398_/A _1548_/B VGND VGND VPWR VPWR _0991_/X sky130_fd_sc_hd__and3_1
XFILLER_0_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1543_ _1236_/C _1542_/Y _1541_/Y VGND VGND VPWR VPWR _1592_/D sky130_fd_sc_hd__o21a_1
X_1474_ _1185_/X _1473_/X _1016_/Y VGND VGND VPWR VPWR _1474_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1190_ _1190_/A _1190_/B _1258_/A _0944_/Y VGND VGND VPWR VPWR _1190_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0974_ _1063_/A _1025_/A VGND VGND VPWR VPWR _1267_/A sky130_fd_sc_hd__nor2_2
X_1526_ _1600_/Q hold7/A _1560_/A _1526_/D VGND VGND VPWR VPWR _1527_/C sky130_fd_sc_hd__and4_1
X_1457_ _1210_/A _1456_/X _1211_/X _1111_/B VGND VGND VPWR VPWR _1457_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1388_ _1190_/A _1380_/X _1383_/Y _1387_/X _1166_/A VGND VGND VPWR VPWR _1388_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1311_ _1307_/X _1310_/Y _0843_/Y VGND VGND VPWR VPWR _1312_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_2_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1242_ _1252_/A _1111_/B _0877_/B _1205_/B _1110_/Y VGND VGND VPWR VPWR _1242_/X
+ sky130_fd_sc_hd__o32a_1
X_1173_ _1169_/X _1172_/Y _1555_/A VGND VGND VPWR VPWR _1173_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0957_ _1405_/A _1405_/B VGND VGND VPWR VPWR _0957_/Y sky130_fd_sc_hd__nand2_1
X_0888_ _1074_/A _0888_/B VGND VGND VPWR VPWR _1394_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1509_ _1516_/A1 _1506_/X _1508_/Y _1524_/B hold9/X VGND VGND VPWR VPWR _1579_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0811_ _1362_/B _0953_/A VGND VGND VPWR VPWR _0811_/X sky130_fd_sc_hd__and2_1
XFILLER_0_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1225_ _1225_/A _1225_/B _1225_/C VGND VGND VPWR VPWR _1225_/X sky130_fd_sc_hd__or3_1
X_1156_ _1154_/X _1320_/C _0953_/A _1114_/A _1405_/C VGND VGND VPWR VPWR _1159_/A
+ sky130_fd_sc_hd__o2111a_1
X_1087_ _0814_/B _1087_/A2 _1086_/Y _0883_/Y VGND VGND VPWR VPWR _1087_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ _1010_/A _1010_/B VGND VGND VPWR VPWR _1010_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1208_ _1420_/A _1394_/A _1475_/A _1393_/A VGND VGND VPWR VPWR _1208_/X sky130_fd_sc_hd__or4_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ _1098_/X _1099_/X _1103_/X _1138_/X VGND VGND VPWR VPWR _1139_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_7_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1490_ _1176_/A _1448_/X _1489_/Y hold4/A _1432_/X VGND VGND VPWR VPWR _1490_/Y sky130_fd_sc_hd__a311oi_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0990_ _1281_/C _0986_/Y _0989_/Y _1452_/C _0962_/C VGND VGND VPWR VPWR _0990_/X
+ sky130_fd_sc_hd__o32a_1
X_1542_ _1542_/A _1542_/B VGND VGND VPWR VPWR _1542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_22_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1473_ _1074_/C _0944_/Y _1029_/Y _0876_/X _1483_/A VGND VGND VPWR VPWR _1473_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0973_ _0817_/Y _1483_/A _0936_/Y _0862_/Y _1036_/A VGND VGND VPWR VPWR _0973_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1525_ hold2/X _1525_/B VGND VGND VPWR VPWR _1587_/D sky130_fd_sc_hd__and2_1
X_1387_ _1112_/A _0947_/Y _0955_/X _1386_/Y _0843_/Y VGND VGND VPWR VPWR _1387_/X
+ sky130_fd_sc_hd__o2111a_1
X_1456_ _1212_/A _0933_/Y _1208_/X _1455_/X _1162_/Y VGND VGND VPWR VPWR _1456_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ _1181_/A _1218_/Y _1309_/X _1112_/A VGND VGND VPWR VPWR _1310_/Y sky130_fd_sc_hd__o22ai_1
X_1241_ _0854_/X _1343_/C VGND VGND VPWR VPWR _1241_/Y sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_19_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1172_ fanout6/X _1135_/X _1171_/X VGND VGND VPWR VPWR _1172_/Y sky130_fd_sc_hd__a21oi_1
X_0956_ _1258_/A _0948_/X _1384_/B _0954_/Y VGND VGND VPWR VPWR _1393_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0887_ _0887_/A _0887_/B _0868_/X VGND VGND VPWR VPWR _0887_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_2_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1439_ _1439_/A _1439_/B VGND VGND VPWR VPWR _1439_/Y sky130_fd_sc_hd__nand2_1
X_1508_ _1513_/C VGND VGND VPWR VPWR _1508_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0810_ hold4/X _0808_/X _0809_/X VGND VGND VPWR VPWR _1607_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1224_ _1281_/C _1223_/X _1462_/A _1099_/X VGND VGND VPWR VPWR _1225_/C sky130_fd_sc_hd__o211a_1
X_1086_ _1184_/A _1362_/D VGND VGND VPWR VPWR _1086_/Y sky130_fd_sc_hd__nand2_1
X_1155_ _1362_/B _1362_/D VGND VGND VPWR VPWR _1320_/C sky130_fd_sc_hd__nor2_1
X_0939_ _1114_/C _1342_/A VGND VGND VPWR VPWR _0939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_2__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload2/A sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1207_ _1205_/Y _1206_/X _1010_/Y VGND VGND VPWR VPWR _1207_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1069_ _0940_/Y _1064_/X _1183_/B _1068_/Y _1352_/A VGND VGND VPWR VPWR _1071_/D
+ sky130_fd_sc_hd__a32o_1
X_1138_ _1105_/X _1106_/X _1107_/Y _1555_/A VGND VGND VPWR VPWR _1138_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1541_ _1551_/B _1533_/A _1560_/B VGND VGND VPWR VPWR _1541_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1472_ _1468_/Y _1470_/X _1471_/X _1419_/A VGND VGND VPWR VPWR _1472_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0972_ _1439_/A _0957_/Y _1256_/B _0971_/X _1398_/B VGND VGND VPWR VPWR _0972_/X
+ sky130_fd_sc_hd__a311o_1
X_1524_ hold3/X _1524_/B VGND VGND VPWR VPWR _1586_/D sky130_fd_sc_hd__and2_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1386_ _1384_/X _1385_/X _0903_/B VGND VGND VPWR VPWR _1386_/Y sky130_fd_sc_hd__o21ai_2
X_1455_ _1074_/A _1420_/C _1075_/A _1443_/S _1111_/B VGND VGND VPWR VPWR _1455_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1240_ _1238_/X _1239_/X _1247_/B _1235_/X VGND VGND VPWR VPWR _1251_/A sky130_fd_sc_hd__a211oi_1
X_1171_ _1135_/A _1054_/A _1170_/Y _1334_/A _1210_/A VGND VGND VPWR VPWR _1171_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_19_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0955_ _1236_/C _0955_/B _1057_/A _1181_/A VGND VGND VPWR VPWR _0955_/X sky130_fd_sc_hd__or4b_4
XFILLER_0_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0886_ _1323_/B _1551_/A _0877_/Y _0885_/X VGND VGND VPWR VPWR _0887_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1507_ _1577_/Q _1576_/Q hold9/A _1578_/Q VGND VGND VPWR VPWR _1513_/C sky130_fd_sc_hd__and4_1
XFILLER_0_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1369_ _1356_/X _1360_/X _1368_/X _1599_/Q VGND VGND VPWR VPWR _1369_/X sky130_fd_sc_hd__o31a_1
X_1438_ _1438_/A _1438_/B _1375_/Y _1376_/X VGND VGND VPWR VPWR _1438_/X sky130_fd_sc_hd__or4bb_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1223_ _0985_/B _1039_/B _0957_/Y VGND VGND VPWR VPWR _1223_/X sky130_fd_sc_hd__o21a_1
X_1154_ _0931_/A _0848_/X _1281_/B _0931_/B VGND VGND VPWR VPWR _1154_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1085_ _1335_/A _1534_/S VGND VGND VPWR VPWR _1085_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0869_ _0869_/A _0869_/B VGND VGND VPWR VPWR _0903_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0938_ _0814_/B _0923_/B _1260_/C VGND VGND VPWR VPWR _1452_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1206_ _1420_/C _0939_/Y _1399_/A VGND VGND VPWR VPWR _1206_/X sky130_fd_sc_hd__a21o_1
X_1137_ _1121_/X _1129_/X _1133_/Y _1190_/A VGND VGND VPWR VPWR _1137_/X sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1068_ _1162_/B _0877_/B _0953_/X VGND VGND VPWR VPWR _1068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ _1361_/Y _1542_/B _1544_/B _1539_/Y VGND VGND VPWR VPWR _1591_/D sky130_fd_sc_hd__o31ai_1
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1471_ _1471_/A1 _0817_/B _1200_/X _1202_/X VGND VGND VPWR VPWR _1471_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0971_ _1197_/A _0885_/C _1212_/A VGND VGND VPWR VPWR _0971_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1523_ hold6/X _1524_/B VGND VGND VPWR VPWR _1585_/D sky130_fd_sc_hd__and2_1
X_1454_ _1454_/A _1454_/B _1452_/X VGND VGND VPWR VPWR _1454_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1385_ _0991_/A _1393_/A _0864_/B _1394_/A VGND VGND VPWR VPWR _1385_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_9_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1170_ _1195_/B _1085_/Y _1199_/D VGND VGND VPWR VPWR _1170_/Y sky130_fd_sc_hd__a21oi_1
X_0954_ _1281_/C _1260_/C VGND VGND VPWR VPWR _0954_/Y sky130_fd_sc_hd__nor2_1
X_0885_ _1237_/A _0885_/B _0885_/C VGND VGND VPWR VPWR _0885_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1506_ _1577_/Q _1576_/Q _1578_/Q hold9/A VGND VGND VPWR VPWR _1506_/X sky130_fd_sc_hd__a31o_1
X_1437_ _1551_/A _1210_/A _1436_/Y _1433_/X VGND VGND VPWR VPWR _1438_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1368_ _1281_/C _0932_/Y _1364_/Y _1367_/X _0878_/Y VGND VGND VPWR VPWR _1368_/X
+ sky130_fd_sc_hd__o2111a_1
X_1299_ _1300_/A _1300_/B VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1153_ _1150_/X _1565_/B _1152_/X _0789_/Y VGND VGND VPWR VPWR _1153_/Y sky130_fd_sc_hd__a31oi_1
X_1222_ _1035_/A _1154_/X _1195_/Y _1221_/X _1323_/B VGND VGND VPWR VPWR _1462_/A
+ sky130_fd_sc_hd__o2111ai_2
X_1084_ _0849_/B _1084_/B VGND VGND VPWR VPWR _1362_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0868_ _1339_/B _0859_/X _1183_/A _0867_/Y _1181_/A VGND VGND VPWR VPWR _0868_/X
+ sky130_fd_sc_hd__a311o_1
X_0937_ _1378_/A1 _0923_/B _0926_/A VGND VGND VPWR VPWR _0937_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0799_ _1317_/A VGND VGND VPWR VPWR _0799_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1205_ _1205_/A _1205_/B VGND VGND VPWR VPWR _1205_/Y sky130_fd_sc_hd__nand2_1
X_1136_ _0980_/Y _1021_/Y _1135_/X _1210_/A VGND VGND VPWR VPWR _1136_/X sky130_fd_sc_hd__a22o_1
X_1067_ _1483_/A _1205_/A VGND VGND VPWR VPWR _1067_/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _1119_/A _1475_/D _1146_/B _1343_/C VGND VGND VPWR VPWR _1119_/X sky130_fd_sc_hd__or4_1
XFILLER_0_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ _1439_/A _1197_/X _1469_/Y _1196_/X VGND VGND VPWR VPWR _1470_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1599_ clkload0/A _1599_/D fanout120/X VGND VGND VPWR VPWR _1599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0970_ _0931_/A _1100_/A _1100_/B _0953_/A _0931_/B VGND VGND VPWR VPWR _1039_/B
+ sky130_fd_sc_hd__o311ai_4
X_1522_ hold5/X _1524_/B VGND VGND VPWR VPWR _1584_/D sky130_fd_sc_hd__and2_1
X_1453_ _1074_/A _0952_/B _1125_/X _1452_/C _1548_/A VGND VGND VPWR VPWR _1454_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1384_ _1384_/A _1384_/B _1434_/C VGND VGND VPWR VPWR _1384_/X sky130_fd_sc_hd__and3_1
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0884_ _0836_/A _0931_/B _0928_/B _0985_/B VGND VGND VPWR VPWR _0885_/C sky130_fd_sc_hd__o31ai_2
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0953_ _0953_/A _0985_/B _1114_/A VGND VGND VPWR VPWR _0953_/X sky130_fd_sc_hd__or3_2
XFILLER_0_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1505_ _1516_/A1 _1503_/X _1504_/Y _1524_/B _1578_/Q VGND VGND VPWR VPWR _1578_/D
+ sky130_fd_sc_hd__a32o_1
X_1436_ _1436_/A _1436_/B VGND VGND VPWR VPWR _1436_/Y sky130_fd_sc_hd__nand2_1
X_1367_ _1367_/A1 _1195_/Y _1366_/X VGND VGND VPWR VPWR _1367_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1298_ _0928_/B wire10/X _1283_/C VGND VGND VPWR VPWR _1298_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1221_ _1035_/A _1135_/A _1286_/C _1001_/B _1439_/A VGND VGND VPWR VPWR _1221_/X
+ sky130_fd_sc_hd__a41o_1
X_1083_ _1081_/X _1082_/Y _1010_/B VGND VGND VPWR VPWR _1083_/X sky130_fd_sc_hd__a21o_1
X_1152_ _1405_/C _1048_/Y _1131_/B _1225_/A VGND VGND VPWR VPWR _1152_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0936_ _0930_/B _0923_/B _0930_/D VGND VGND VPWR VPWR _0936_/Y sky130_fd_sc_hd__a21oi_4
X_0867_ _0955_/B _1450_/A _1339_/B VGND VGND VPWR VPWR _0867_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0798_ _0985_/B VGND VGND VPWR VPWR _1211_/A sky130_fd_sc_hd__inv_2
X_1419_ _1419_/A _1419_/B _1419_/C VGND VGND VPWR VPWR _1423_/C sky130_fd_sc_hd__or3_1
XFILLER_0_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1204_ _1204_/A _1204_/B _1204_/C VGND VGND VPWR VPWR _1204_/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1066_ _1066_/A _1452_/A _1015_/B VGND VGND VPWR VPWR _1475_/D sky130_fd_sc_hd__or3b_2
X_1135_ _1135_/A _1135_/B VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__and2_1
X_0919_ _0858_/B _1180_/A _0918_/Y _1526_/D VGND VGND VPWR VPWR _0920_/C sky130_fd_sc_hd__a31o_1
XFILLER_0_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1118_ _1118_/A _1118_/B VGND VGND VPWR VPWR _1343_/C sky130_fd_sc_hd__xnor2_4
X_1049_ _1074_/B _1029_/B _1074_/A VGND VGND VPWR VPWR _1411_/C sky130_fd_sc_hd__a21oi_4
XFILLER_0_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1598_ clkload1/A _1598_/D fanout120/X VGND VGND VPWR VPWR _1598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1521_ hold11/X _1497_/Y _1518_/B _1520_/X VGND VGND VPWR VPWR _1583_/D sky130_fd_sc_hd__a31o_1
X_1383_ _0922_/Y _1037_/B _1382_/X VGND VGND VPWR VPWR _1383_/Y sky130_fd_sc_hd__o21ai_1
X_1452_ _1452_/A _1548_/A _1452_/C VGND VGND VPWR VPWR _1452_/X sky130_fd_sc_hd__or3_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0952_ _0989_/A _0952_/B VGND VGND VPWR VPWR _1037_/B sky130_fd_sc_hd__or2_2
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1504_ _1577_/Q _1576_/Q _1578_/Q VGND VGND VPWR VPWR _1504_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0883_ _1114_/C _0885_/B VGND VGND VPWR VPWR _0883_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1435_ _1405_/A _1548_/B _1450_/A VGND VGND VPWR VPWR _1436_/B sky130_fd_sc_hd__o21ai_1
X_1366_ _1212_/A _0933_/B _1365_/X _1323_/B VGND VGND VPWR VPWR _1366_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1297_ _1285_/Y _1290_/X _1292_/X _1296_/X _1560_/A VGND VGND VPWR VPWR _1312_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1151_ _1166_/A _1563_/S VGND VGND VPWR VPWR _1565_/B sky130_fd_sc_hd__nor2_2
X_1220_ _1258_/A _1219_/X _1217_/Y _1216_/X VGND VGND VPWR VPWR _1225_/B sky130_fd_sc_hd__o211a_1
X_1082_ _0827_/X _1119_/A _1439_/A VGND VGND VPWR VPWR _1082_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0935_ _0921_/Y _0924_/X _0934_/X _1452_/A _1258_/A VGND VGND VPWR VPWR _0935_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0866_ _0873_/A _0930_/B _1118_/B _1117_/B VGND VGND VPWR VPWR _1450_/A sky130_fd_sc_hd__a31o_4
XFILLER_0_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0797_ _0953_/A VGND VGND VPWR VPWR _0797_/Y sky130_fd_sc_hd__inv_2
X_1418_ _1256_/A _1260_/A _1210_/A _0996_/A _0930_/D VGND VGND VPWR VPWR _1419_/C
+ sky130_fd_sc_hd__o2111a_1
X_1349_ _0923_/Y _1205_/B _1483_/C _1067_/Y VGND VGND VPWR VPWR _1356_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1134_ _1442_/A _1063_/Y _0954_/Y _1010_/A VGND VGND VPWR VPWR _1134_/X sky130_fd_sc_hd__a211o_1
X_1203_ _1194_/Y _1198_/X _1202_/X _1419_/A VGND VGND VPWR VPWR _1204_/C sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1065_ _1526_/D _1281_/C VGND VGND VPWR VPWR _1183_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0918_ _0932_/A _1229_/A VGND VGND VPWR VPWR _0918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0849_ _1084_/B _0849_/B VGND VGND VPWR VPWR _1229_/A sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_3_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1117_ _0814_/B _1117_/B VGND VGND VPWR VPWR _1146_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1048_ _1334_/A VGND VGND VPWR VPWR _1048_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1597_ _1597_/CLK _1597_/D fanout119/X VGND VGND VPWR VPWR _1597_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1520_ _1525_/B _1497_/Y hold13/X VGND VGND VPWR VPWR _1520_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1451_ _1205_/Y _1449_/X _1450_/Y _1010_/Y VGND VGND VPWR VPWR _1451_/X sky130_fd_sc_hd__a31o_1
X_1382_ _1063_/A _1258_/A _1381_/X _1180_/A VGND VGND VPWR VPWR _1382_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0951_ _1256_/A _1317_/A VGND VGND VPWR VPWR _1205_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0882_ _1114_/A _1318_/A VGND VGND VPWR VPWR _1460_/B sky130_fd_sc_hd__nand2b_1
X_1503_ _1577_/Q _1576_/Q _1578_/Q VGND VGND VPWR VPWR _1503_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1434_ _1434_/A wire10/X _1434_/C VGND VGND VPWR VPWR _1438_/A sky130_fd_sc_hd__and3_1
X_1296_ _1294_/Y _1295_/X _1015_/Y VGND VGND VPWR VPWR _1296_/X sky130_fd_sc_hd__o21a_1
X_1365_ _1229_/A _0861_/X _1357_/A _1035_/B VGND VGND VPWR VPWR _1365_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1150_ _1010_/Y _1149_/X _1145_/Y _1190_/B VGND VGND VPWR VPWR _1150_/X sky130_fd_sc_hd__a2bb2o_1
X_1081_ _0926_/A _1548_/B _1037_/B VGND VGND VPWR VPWR _1081_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0865_ _0991_/A _0933_/A VGND VGND VPWR VPWR _1394_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0934_ _0817_/B _1114_/C _1420_/D _1260_/C VGND VGND VPWR VPWR _0934_/X sky130_fd_sc_hd__o22a_1
X_0796_ _1335_/A VGND VGND VPWR VPWR _1384_/A sky130_fd_sc_hd__inv_2
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1417_ _1011_/X _1013_/Y _1416_/X _1197_/B fanout6/X VGND VGND VPWR VPWR _1423_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1279_ _1281_/C _1544_/A _1405_/C _0870_/Y _1195_/A VGND VGND VPWR VPWR _1282_/A
+ sky130_fd_sc_hd__o32a_1
X_1348_ _0936_/Y _0975_/Y _1078_/X VGND VGND VPWR VPWR _1348_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1133_ _0996_/A _1130_/Y _1132_/X fanout6/X VGND VGND VPWR VPWR _1133_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1064_ _1405_/A _1420_/C _1252_/B _1398_/A VGND VGND VPWR VPWR _1064_/X sky130_fd_sc_hd__a211o_1
X_1202_ _1483_/C _1202_/B _1202_/C VGND VGND VPWR VPWR _1202_/X sky130_fd_sc_hd__or3_1
XFILLER_0_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0917_ _1252_/A _0908_/Y _0915_/Y _0885_/B VGND VGND VPWR VPWR _0920_/B sky130_fd_sc_hd__o211a_1
X_0848_ _1100_/A _1100_/B VGND VGND VPWR VPWR _0848_/X sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1116_ _1483_/A _1116_/B _1116_/C VGND VGND VPWR VPWR _1116_/X sky130_fd_sc_hd__or3_1
X_1047_ _1135_/A _1548_/A VGND VGND VPWR VPWR _1334_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ _1597_/CLK _1596_/D fanout117/X VGND VGND VPWR VPWR _1596_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1450_ _1450_/A _1450_/B VGND VGND VPWR VPWR _1450_/Y sky130_fd_sc_hd__nand2_1
X_1381_ _0888_/B _1408_/C _1063_/B VGND VGND VPWR VPWR _1381_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1579_ _1597_/CLK _1579_/D fanout118/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0950_ _1199_/D _1199_/C VGND VGND VPWR VPWR _1335_/B sky130_fd_sc_hd__nand2b_1
X_0881_ _1114_/A _1323_/B VGND VGND VPWR VPWR _0885_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1502_ _1516_/A1 _1500_/X _1501_/Y _1524_/B _1577_/Q VGND VGND VPWR VPWR _1577_/D
+ sky130_fd_sc_hd__a32o_1
X_1433_ _0811_/X _1286_/X _1183_/B _0955_/B VGND VGND VPWR VPWR _1433_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1295_ _0957_/Y _1267_/A _1293_/Y _1398_/B _1405_/C VGND VGND VPWR VPWR _1295_/X
+ sky130_fd_sc_hd__a32o_1
X_1364_ _1364_/A _1364_/B VGND VGND VPWR VPWR _1364_/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1080_ fanout6/X _1079_/X _1077_/X _1225_/A VGND VGND VPWR VPWR _1089_/A sky130_fd_sc_hd__o211ai_1
XFILLER_0_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0933_ _0933_/A _0933_/B VGND VGND VPWR VPWR _0933_/Y sky130_fd_sc_hd__nand2_2
X_0864_ _1394_/A _0864_/B VGND VGND VPWR VPWR _1183_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0795_ _0931_/B VGND VGND VPWR VPWR _1361_/A sky130_fd_sc_hd__inv_2
XFILLER_0_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1347_ _1312_/X _1346_/X _1599_/Q VGND VGND VPWR VPWR _1347_/X sky130_fd_sc_hd__a21o_1
X_1416_ _1025_/A _0940_/Y _1394_/C _1063_/A VGND VGND VPWR VPWR _1416_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1278_ _1204_/X _1226_/X _1489_/B _1277_/X VGND VGND VPWR VPWR _1278_/Y sky130_fd_sc_hd__o211ai_1
Xwire10 wire10/A VGND VGND VPWR VPWR wire10/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1201_ _1111_/A _1197_/B _1200_/X VGND VGND VPWR VPWR _1202_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1132_ _0989_/A _1116_/B _1131_/Y _0952_/B _0989_/Y VGND VGND VPWR VPWR _1132_/X
+ sky130_fd_sc_hd__a221o_1
X_1063_ _1063_/A _1063_/B VGND VGND VPWR VPWR _1063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0916_ _0932_/A _0991_/A VGND VGND VPWR VPWR _1544_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0847_ _0851_/A _0900_/C _1236_/B VGND VGND VPWR VPWR _1361_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1046_ _1039_/Y _1044_/X _1045_/X VGND VGND VPWR VPWR _1046_/Y sky130_fd_sc_hd__a21oi_2
X_1115_ _0817_/Y _1267_/A _1114_/X VGND VGND VPWR VPWR _1115_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_28_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1595_ clkload2/A _1595_/D fanout117/X VGND VGND VPWR VPWR _1595_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1029_ _1074_/B _1029_/B VGND VGND VPWR VPWR _1029_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1380_ _1066_/A _1483_/A _1379_/X _1210_/A VGND VGND VPWR VPWR _1380_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1578_ clkload2/A _1578_/D fanout118/X VGND VGND VPWR VPWR _1578_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ _0851_/A _1236_/D _1236_/C _0955_/B VGND VGND VPWR VPWR _1237_/A sky130_fd_sc_hd__a31o_2
XFILLER_0_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1432_ _1176_/C _1431_/X _1601_/Q VGND VGND VPWR VPWR _1432_/X sky130_fd_sc_hd__o21a_1
X_1501_ _1577_/Q _1576_/Q VGND VGND VPWR VPWR _1501_/Y sky130_fd_sc_hd__nand2_1
X_1363_ _0955_/B _0923_/Y _1361_/Y _1102_/B _0903_/B VGND VGND VPWR VPWR _1364_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1294_ _1294_/A _1436_/A VGND VGND VPWR VPWR _1294_/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0932_ _0932_/A _1039_/A VGND VGND VPWR VPWR _0932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0863_ _0851_/A _1236_/D _1236_/C VGND VGND VPWR VPWR _0864_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0794_ _1362_/A VGND VGND VPWR VPWR _1184_/A sky130_fd_sc_hd__inv_2
X_1346_ _1555_/A _1345_/X _1331_/X _1322_/X VGND VGND VPWR VPWR _1346_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1415_ _1415_/A _1415_/B _1415_/C _1415_/D VGND VGND VPWR VPWR _1424_/B sky130_fd_sc_hd__or4_1
XFILLER_0_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1277_ _1488_/A _1277_/B _1276_/X VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__or3b_1
Xfanout120 input2/X VGND VGND VPWR VPWR fanout120/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1200_ _1200_/A1 _0996_/A _1283_/C _1205_/B VGND VGND VPWR VPWR _1200_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1131_ _1131_/A _1131_/B VGND VGND VPWR VPWR _1131_/Y sky130_fd_sc_hd__nor2_1
X_1062_ _1060_/X _1061_/X _1483_/C VGND VGND VPWR VPWR _1428_/A sky130_fd_sc_hd__a21oi_1
X_0915_ _1252_/A _1252_/B VGND VGND VPWR VPWR _0915_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0846_ _1118_/A _1072_/B VGND VGND VPWR VPWR _1029_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1329_ _1114_/C _1320_/D _1328_/X _1323_/B VGND VGND VPWR VPWR _1329_/X sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_34_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1114_ _1114_/A _1114_/B _1114_/C VGND VGND VPWR VPWR _1114_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1045_ _0985_/B _1039_/A _1039_/B _1114_/A VGND VGND VPWR VPWR _1045_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0829_ _1256_/A _1317_/A VGND VGND VPWR VPWR _0829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1594_ clkload2/A _1594_/D fanout117/X VGND VGND VPWR VPWR _1594_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1028_ _1063_/A _1028_/B VGND VGND VPWR VPWR _1028_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1577_ clkload2/A _1577_/D fanout118/X VGND VGND VPWR VPWR _1577_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1500_ _1577_/Q _1576_/Q VGND VGND VPWR VPWR _1500_/X sky130_fd_sc_hd__or2_1
XFILLER_0_2_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1431_ _0943_/X _1404_/X _1424_/X _1430_/Y _0789_/Y VGND VGND VPWR VPWR _1431_/X
+ sky130_fd_sc_hd__o221a_1
X_1293_ _1111_/B _1119_/A _1237_/B VGND VGND VPWR VPWR _1293_/Y sky130_fd_sc_hd__a21oi_1
X_1362_ _1362_/A _1362_/B _1362_/C _1362_/D VGND VGND VPWR VPWR _1364_/A sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _0931_/A _0931_/B _1100_/B _1035_/A VGND VGND VPWR VPWR _1039_/A sky130_fd_sc_hd__or4_4
X_0862_ _1074_/A _1475_/A VGND VGND VPWR VPWR _0862_/Y sky130_fd_sc_hd__nor2_1
X_0793_ _1599_/Q VGND VGND VPWR VPWR _1563_/S sky130_fd_sc_hd__inv_2
XFILLER_0_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1345_ _1345_/A _1345_/B _1345_/C _1345_/D VGND VGND VPWR VPWR _1345_/X sky130_fd_sc_hd__or4_1
XFILLER_0_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1414_ _1483_/C _1414_/B _1414_/C VGND VGND VPWR VPWR _1415_/D sky130_fd_sc_hd__nor3_1
X_1276_ _1471_/A1 _1434_/A _1268_/Y _1275_/Y VGND VGND VPWR VPWR _1276_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout110 _1588_/Q VGND VGND VPWR VPWR _1200_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1130_ _0989_/A _1116_/B _0989_/Y VGND VGND VPWR VPWR _1130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1061_ _1256_/A _1450_/A _1233_/B _0888_/B _1317_/A VGND VGND VPWR VPWR _1061_/X
+ sky130_fd_sc_hd__a221o_1
X_0845_ _1118_/A _1072_/B VGND VGND VPWR VPWR _1119_/A sky130_fd_sc_hd__and2_2
X_0914_ _1063_/A _1063_/B VGND VGND VPWR VPWR _0914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1259_ _1483_/A _1259_/B _1483_/C VGND VGND VPWR VPWR _1259_/X sky130_fd_sc_hd__or3_1
X_1328_ _0931_/A _0848_/X _1281_/B _1361_/A VGND VGND VPWR VPWR _1328_/X sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_34_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1044_ _1339_/D _1043_/B _1323_/A VGND VGND VPWR VPWR _1044_/X sky130_fd_sc_hd__a21o_1
X_1113_ _1258_/A _1109_/X _1110_/Y _1021_/B _1108_/X VGND VGND VPWR VPWR _1113_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0828_ _1398_/A _1339_/B VGND VGND VPWR VPWR _0828_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1593_ clkload2/A _1593_/D fanout119/X VGND VGND VPWR VPWR _1593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ _1063_/A _1028_/B VGND VGND VPWR VPWR _1317_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1576_ _1597_/CLK _1576_/D fanout118/X VGND VGND VPWR VPWR _1576_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1430_ _1089_/Y _1429_/X _1563_/S VGND VGND VPWR VPWR _1430_/Y sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1361_ _1361_/A _1361_/B VGND VGND VPWR VPWR _1361_/Y sky130_fd_sc_hd__xnor2_1
X_1292_ _1551_/C _1292_/B VGND VGND VPWR VPWR _1292_/X sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1559_ _1560_/B _1559_/B VGND VGND VPWR VPWR _1559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0792_ _1424_/A VGND VGND VPWR VPWR _1166_/A sky130_fd_sc_hd__inv_2
XFILLER_0_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0930_ _1118_/A _0930_/B _1118_/B _0930_/D VGND VGND VPWR VPWR _1259_/B sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_15_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0861_ _1362_/A _1106_/A VGND VGND VPWR VPWR _0861_/X sky130_fd_sc_hd__or2_2
XFILLER_0_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1413_ _1025_/Y _1028_/X _1029_/Y _1181_/B _0980_/Y VGND VGND VPWR VPWR _1414_/C
+ sky130_fd_sc_hd__o221a_1
X_1344_ _1434_/A _1308_/X _1343_/X _1342_/X _1183_/B VGND VGND VPWR VPWR _1345_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1275_ _1483_/C _1270_/X _1272_/X _1274_/X VGND VGND VPWR VPWR _1275_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout100 _1590_/Q VGND VGND VPWR VPWR _1199_/C sky130_fd_sc_hd__buf_2
Xfanout111 _0900_/C VGND VGND VPWR VPWR _1084_/B sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _0930_/D _0962_/B _1060_/B1 _1036_/A VGND VGND VPWR VPWR _1060_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0844_ _1195_/A _1442_/A _1560_/A _1526_/D _0833_/Y VGND VGND VPWR VPWR _0844_/X
+ sky130_fd_sc_hd__a2111o_1
X_0913_ _1072_/B _0913_/A2 _1117_/B _1378_/A1 _1118_/A VGND VGND VPWR VPWR _1063_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1189_ _1443_/S _0922_/Y _1188_/X _0933_/Y _1200_/A1 VGND VGND VPWR VPWR _1189_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_26_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1327_ _1405_/A _1195_/B _1074_/C _1037_/B _1029_/Y VGND VGND VPWR VPWR _1327_/X
+ sky130_fd_sc_hd__a2111o_1
X_1258_ _1258_/A _1258_/B VGND VGND VPWR VPWR _1258_/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1043_ _1339_/D _1043_/B VGND VGND VPWR VPWR _1181_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1112_ _1112_/A _1317_/B _1112_/C VGND VGND VPWR VPWR _1112_/X sky130_fd_sc_hd__or3_1
XFILLER_0_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0827_ _1199_/C _1335_/A _0991_/A _1094_/A VGND VGND VPWR VPWR _0827_/X sky130_fd_sc_hd__a211o_2
XFILLER_0_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1592_ clkload2/A _1592_/D fanout119/X VGND VGND VPWR VPWR _1592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1026_ _1072_/B _1118_/B _1117_/B _0930_/B _0873_/A VGND VGND VPWR VPWR _1028_/B
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1575_ clkload1/A hold1/X fanout120/X VGND VGND VPWR VPWR uo_out[0] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1190_/B _1258_/A VGND VGND VPWR VPWR _1551_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1360_ _0843_/Y _1359_/X _1424_/A VGND VGND VPWR VPWR _1360_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1291_ _0908_/Y _0995_/Y _1001_/B _1076_/Y _1135_/A VGND VGND VPWR VPWR _1292_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_18_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1558_ _1424_/A _1570_/C _1544_/B VGND VGND VPWR VPWR _1559_/B sky130_fd_sc_hd__a21o_1
X_1489_ _1600_/Q _1489_/B _1489_/C _1489_/D VGND VGND VPWR VPWR _1489_/Y sky130_fd_sc_hd__nand4_1
XFILLER_0_17_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ _1066_/A VGND VGND VPWR VPWR _1190_/B sky130_fd_sc_hd__inv_2
XFILLER_0_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0860_ _0931_/A _0931_/B VGND VGND VPWR VPWR _1475_/A sky130_fd_sc_hd__nor2_4
X_1343_ _1384_/B _1362_/C _1343_/C VGND VGND VPWR VPWR _1343_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1412_ _1046_/Y _1411_/X _1116_/C VGND VGND VPWR VPWR _1415_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1274_ _1454_/B _1273_/X _1555_/A VGND VGND VPWR VPWR _1274_/X sky130_fd_sc_hd__o21a_1
X_0989_ _0989_/A _1056_/B VGND VGND VPWR VPWR _0989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout101 _0913_/A2 VGND VGND VPWR VPWR _1118_/B sky130_fd_sc_hd__buf_4
Xfanout112 _0900_/C VGND VGND VPWR VPWR _1100_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0912_ _1084_/B _0849_/B _0953_/A _1362_/B _1362_/A VGND VGND VPWR VPWR _1252_/B
+ sky130_fd_sc_hd__o2111a_1
X_0843_ _1597_/Q _1010_/A VGND VGND VPWR VPWR _0843_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1326_ _1398_/B _1325_/Y _0869_/B VGND VGND VPWR VPWR _1326_/Y sky130_fd_sc_hd__a21oi_1
X_1188_ _0827_/X _1119_/A _0864_/B VGND VGND VPWR VPWR _1188_/X sky130_fd_sc_hd__o21a_1
X_1257_ _1439_/A _1256_/B _1267_/B _1281_/A _1212_/A VGND VGND VPWR VPWR _1258_/B
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1111_ _1111_/A _1111_/B VGND VGND VPWR VPWR _1112_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1042_ _1084_/B _0851_/D _0836_/A VGND VGND VPWR VPWR _1043_/B sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_31_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0826_ _1199_/D _0928_/B VGND VGND VPWR VPWR _1110_/B sky130_fd_sc_hd__or2_1
X_1309_ _1308_/X _1309_/B VGND VGND VPWR VPWR _1309_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1591_ clkload2/A _1591_/D fanout119/X VGND VGND VPWR VPWR _1591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1025_ _1025_/A _1025_/B VGND VGND VPWR VPWR _1025_/Y sky130_fd_sc_hd__nand2_2
X_0809_ _0801_/Y _0807_/C _1525_/B VGND VGND VPWR VPWR _0809_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 _1112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1574_ _1597_/CLK _1574_/D fanout117/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1006_/Y _1007_/X _1352_/A VGND VGND VPWR VPWR _1023_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1290_ _1289_/X _1434_/A VGND VGND VPWR VPWR _1290_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1488_ _1488_/A _1488_/B VGND VGND VPWR VPWR _1489_/D sky130_fd_sc_hd__or2_1
X_1557_ _1560_/A _1560_/C VGND VGND VPWR VPWR _1570_/C sky130_fd_sc_hd__and2_1
XFILLER_0_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0790_ _1419_/A VGND VGND VPWR VPWR _0790_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1342_ _1342_/A _1342_/B _1057_/B VGND VGND VPWR VPWR _1342_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1273_ _1135_/A _0995_/B _1405_/C _1181_/B VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__o22a_1
X_1411_ _1439_/A _1542_/A _1411_/C VGND VGND VPWR VPWR _1411_/X sky130_fd_sc_hd__and3_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0988_ _0931_/A _0931_/B _1035_/A VGND VGND VPWR VPWR _0988_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout102 _1040_/B VGND VGND VPWR VPWR _0913_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout113 _1534_/S VGND VGND VPWR VPWR _0900_/C sky130_fd_sc_hd__buf_4
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0842_ _1057_/A _0869_/B VGND VGND VPWR VPWR _1112_/A sky130_fd_sc_hd__nand2_2
X_0911_ _0900_/C _1236_/B _0851_/A _1539_/A VGND VGND VPWR VPWR _1405_/B sky130_fd_sc_hd__o211ai_4
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1256_ _1256_/A _1256_/B VGND VGND VPWR VPWR _1256_/Y sky130_fd_sc_hd__nand2_1
X_1325_ _1084_/B _1420_/C _0861_/X VGND VGND VPWR VPWR _1325_/Y sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _1182_/X _1183_/Y _1186_/X _1190_/A VGND VGND VPWR VPWR _1204_/A sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_4_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1110_ _1135_/A _1110_/B VGND VGND VPWR VPWR _1110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1041_ _0931_/A _1084_/B _1100_/B VGND VGND VPWR VPWR _1339_/D sky130_fd_sc_hd__nand3b_4
XTAP_TAPCELL_ROW_31_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0825_ _1118_/A _0913_/A2 _1378_/A1 VGND VGND VPWR VPWR _0962_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1239_ _1010_/B _1057_/Y _0955_/X _1225_/A VGND VGND VPWR VPWR _1239_/X sky130_fd_sc_hd__o211a_1
X_1308_ _1361_/A _1339_/D _1114_/C VGND VGND VPWR VPWR _1308_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1590_ clkload2/A _1590_/D fanout118/X VGND VGND VPWR VPWR _1590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1024_ _0816_/A _0816_/B _1040_/B _1471_/A1 VGND VGND VPWR VPWR _1025_/B sky130_fd_sc_hd__o31ai_4
X_0808_ _1605_/Q _1606_/Q _1607_/Q VGND VGND VPWR VPWR _0808_/X sky130_fd_sc_hd__and3_1
XFILLER_0_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout4 _1016_/Y VGND VGND VPWR VPWR _1483_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 _1357_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1573_ _1562_/B _1570_/X _1571_/Y hold7/X VGND VGND VPWR VPWR _1603_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1114_/C _1475_/A _0903_/C _1452_/A VGND VGND VPWR VPWR _1007_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1556_ _1225_/A _1562_/B _1560_/C _1555_/X VGND VGND VPWR VPWR _1597_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1487_ _1255_/Y _1483_/X _1484_/X _1486_/X VGND VGND VPWR VPWR _1488_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_17_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1410_ _1454_/B _1409_/X _1419_/A VGND VGND VPWR VPWR _1415_/B sky130_fd_sc_hd__o21ai_1
X_1341_ _0888_/B _1001_/Y _0965_/X VGND VGND VPWR VPWR _1345_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1272_ _1212_/A _1271_/X _1114_/X _1010_/Y VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__a211o_1
X_0987_ _1118_/A _1378_/A1 _0926_/A VGND VGND VPWR VPWR _1056_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1608_ clkload0/A _1608_/D fanout120/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfrtp_1
Xfanout103 _1589_/Q VGND VGND VPWR VPWR _1040_/B sky130_fd_sc_hd__buf_2
Xfanout114 _1588_/Q VGND VGND VPWR VPWR _1534_/S sky130_fd_sc_hd__buf_2
X_1539_ _1539_/A _1542_/B VGND VGND VPWR VPWR _1539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0841_ _0869_/A _1181_/A VGND VGND VPWR VPWR _1442_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ _1534_/S _1335_/A _1199_/C _1199_/D VGND VGND VPWR VPWR _1393_/A sky130_fd_sc_hd__o211a_2
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ _0902_/Y _1185_/X _1483_/C VGND VGND VPWR VPWR _1186_/X sky130_fd_sc_hd__a21o_1
X_1255_ _0903_/A _1021_/Y _1252_/X _1254_/Y _1555_/A VGND VGND VPWR VPWR _1255_/Y
+ sky130_fd_sc_hd__a311oi_2
X_1324_ _1229_/A _1300_/D _1305_/Y _1323_/X VGND VGND VPWR VPWR _1324_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap3 _1497_/Y VGND VGND VPWR VPWR _1516_/A1 sky130_fd_sc_hd__clkbuf_2
X_1040_ _0816_/A _1040_/B VGND VGND VPWR VPWR _1265_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0824_ _0873_/A _0913_/A2 _0930_/B VGND VGND VPWR VPWR _1074_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1238_ _0955_/B _0923_/Y _1039_/A _1237_/Y _0870_/Y VGND VGND VPWR VPWR _1238_/X
+ sky130_fd_sc_hd__a311o_1
X_1169_ _0883_/Y _1167_/Y _1168_/X _1526_/D VGND VGND VPWR VPWR _1169_/X sky130_fd_sc_hd__a31o_1
X_1307_ _1114_/A _1054_/A _1304_/X _1306_/X _1323_/B VGND VGND VPWR VPWR _1307_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1023_ _1423_/A _1023_/B _1023_/C _1023_/D VGND VGND VPWR VPWR _1023_/X sky130_fd_sc_hd__or4_1
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0807_ input1/X _0807_/B _0807_/C VGND VGND VPWR VPWR _1606_/D sky130_fd_sc_hd__and3_1
XFILLER_0_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout5 _1015_/Y VGND VGND VPWR VPWR _1210_/A sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1572_ hold12/X _1560_/X _1571_/Y _1529_/X VGND VGND VPWR VPWR _1602_/D sky130_fd_sc_hd__o211a_1
XANTENNA_3 _1205_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _0989_/A _0827_/X _1004_/Y _0952_/B VGND VGND VPWR VPWR _1006_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1555_ _1555_/A _1555_/B VGND VGND VPWR VPWR _1555_/X sky130_fd_sc_hd__and2_1
XFILLER_0_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1486_ _1116_/C _1485_/X _1275_/Y VGND VGND VPWR VPWR _1486_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1340_ _1399_/A _1338_/X _1339_/X fanout6/X VGND VGND VPWR VPWR _1345_/B sky130_fd_sc_hd__o211a_1
XFILLER_0_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1271_ _0816_/B _1195_/B _1265_/B _1260_/C VGND VGND VPWR VPWR _1271_/X sky130_fd_sc_hd__a31o_1
X_0986_ _1420_/D _1362_/C VGND VGND VPWR VPWR _0986_/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1607_ clkload0/A _1607_/D fanout120/X VGND VGND VPWR VPWR _1607_/Q sky130_fd_sc_hd__dfrtp_1
X_1538_ _0851_/A _1542_/B _1562_/B _1181_/C VGND VGND VPWR VPWR _1590_/D sky130_fd_sc_hd__a22o_1
Xfanout115 _1525_/B VGND VGND VPWR VPWR _1524_/B sky130_fd_sc_hd__buf_2
Xfanout104 _0849_/B VGND VGND VPWR VPWR _1100_/B sky130_fd_sc_hd__buf_4
XFILLER_0_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1469_ _1471_/A1 _0817_/B _1420_/D _0877_/B _1036_/A VGND VGND VPWR VPWR _1469_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_0_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ _0851_/A _0851_/D _1236_/C _0955_/B _1539_/A VGND VGND VPWR VPWR _1195_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1323_ _1323_/A _1323_/B _1101_/B VGND VGND VPWR VPWR _1323_/X sky130_fd_sc_hd__or3b_1
X_1254_ _1025_/A _1253_/X _1063_/Y _1010_/Y VGND VGND VPWR VPWR _1254_/Y sky130_fd_sc_hd__a211oi_1
X_1185_ _1124_/Y _1184_/X _0953_/X VGND VGND VPWR VPWR _1185_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0969_ _1117_/B _1256_/A _1317_/A VGND VGND VPWR VPWR _1181_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0823_ _1256_/A _1317_/A VGND VGND VPWR VPWR _1294_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1306_ _0849_/B _1035_/A _1475_/A _1305_/Y _1162_/B VGND VGND VPWR VPWR _1306_/X
+ sky130_fd_sc_hd__a311o_1
X_1237_ _1237_/A _1237_/B VGND VGND VPWR VPWR _1237_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1099_ _1323_/A _1112_/A _1036_/B _1526_/D VGND VGND VPWR VPWR _1099_/X sky130_fd_sc_hd__o31a_1
X_1168_ _1252_/A _1021_/B _1039_/A _1405_/C _1281_/C VGND VGND VPWR VPWR _1168_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _1362_/C _1020_/X _1021_/Y _1419_/B _1419_/A VGND VGND VPWR VPWR _1023_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0806_ hold4/A _1605_/Q _1606_/Q VGND VGND VPWR VPWR _0807_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout6 _1551_/C VGND VGND VPWR VPWR fanout6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1571_ _1544_/B _1570_/X _1560_/B VGND VGND VPWR VPWR _1571_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 _1004_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ _0926_/A _0962_/B _1443_/S VGND VGND VPWR VPWR _1005_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1554_ _1555_/B _1554_/B VGND VGND VPWR VPWR _1596_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1485_ _1256_/B _0975_/Y _1267_/Y _0862_/Y _1266_/X VGND VGND VPWR VPWR _1485_/X
+ sky130_fd_sc_hd__o221a_1
.ends

