magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 154
rect 189 0 192 154
<< via1 >>
rect 3 0 189 154
<< metal2 >>
rect 3 154 189 157
rect 3 -3 189 0
<< properties >>
string GDS_END 91731964
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91729912
<< end >>
