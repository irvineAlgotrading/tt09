magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< metal2 >>
rect 0 785 56 794
rect 0 705 56 729
rect 0 625 56 649
rect 0 545 56 569
rect 0 465 56 489
rect 0 385 56 409
rect 0 305 56 329
rect 0 225 56 249
rect 0 145 56 169
rect 0 65 56 89
rect 0 0 56 9
<< via2 >>
rect 0 729 56 785
rect 0 649 56 705
rect 0 569 56 625
rect 0 489 56 545
rect 0 409 56 465
rect 0 329 56 385
rect 0 249 56 305
rect 0 169 56 225
rect 0 89 56 145
rect 0 9 56 65
<< metal3 >>
rect -5 785 61 790
rect -5 729 0 785
rect 56 729 61 785
rect -5 705 61 729
rect -5 649 0 705
rect 56 649 61 705
rect -5 625 61 649
rect -5 569 0 625
rect 56 569 61 625
rect -5 545 61 569
rect -5 489 0 545
rect 56 489 61 545
rect -5 465 61 489
rect -5 409 0 465
rect 56 409 61 465
rect -5 385 61 409
rect -5 329 0 385
rect 56 329 61 385
rect -5 305 61 329
rect -5 249 0 305
rect 56 249 61 305
rect -5 225 61 249
rect -5 169 0 225
rect 56 169 61 225
rect -5 145 61 169
rect -5 89 0 145
rect 56 89 61 145
rect -5 65 61 89
rect -5 9 0 65
rect 56 9 61 65
rect -5 4 61 9
<< properties >>
string GDS_END 85412886
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85412114
<< end >>
