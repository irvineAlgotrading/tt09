magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 0 0 466 1072
<< pmos >>
rect 89 36 119 1036
rect 175 36 205 1036
rect 261 36 291 1036
rect 347 36 377 1036
<< pdiff >>
rect 36 983 89 1036
rect 36 949 44 983
rect 78 949 89 983
rect 36 911 89 949
rect 36 877 44 911
rect 78 877 89 911
rect 36 839 89 877
rect 36 805 44 839
rect 78 805 89 839
rect 36 767 89 805
rect 36 733 44 767
rect 78 733 89 767
rect 36 695 89 733
rect 36 661 44 695
rect 78 661 89 695
rect 36 623 89 661
rect 36 589 44 623
rect 78 589 89 623
rect 36 551 89 589
rect 36 517 44 551
rect 78 517 89 551
rect 36 479 89 517
rect 36 445 44 479
rect 78 445 89 479
rect 36 407 89 445
rect 36 373 44 407
rect 78 373 89 407
rect 36 335 89 373
rect 36 301 44 335
rect 78 301 89 335
rect 36 263 89 301
rect 36 229 44 263
rect 78 229 89 263
rect 36 191 89 229
rect 36 157 44 191
rect 78 157 89 191
rect 36 119 89 157
rect 36 85 44 119
rect 78 85 89 119
rect 36 36 89 85
rect 119 983 175 1036
rect 119 949 130 983
rect 164 949 175 983
rect 119 911 175 949
rect 119 877 130 911
rect 164 877 175 911
rect 119 839 175 877
rect 119 805 130 839
rect 164 805 175 839
rect 119 767 175 805
rect 119 733 130 767
rect 164 733 175 767
rect 119 695 175 733
rect 119 661 130 695
rect 164 661 175 695
rect 119 623 175 661
rect 119 589 130 623
rect 164 589 175 623
rect 119 551 175 589
rect 119 517 130 551
rect 164 517 175 551
rect 119 479 175 517
rect 119 445 130 479
rect 164 445 175 479
rect 119 407 175 445
rect 119 373 130 407
rect 164 373 175 407
rect 119 335 175 373
rect 119 301 130 335
rect 164 301 175 335
rect 119 263 175 301
rect 119 229 130 263
rect 164 229 175 263
rect 119 191 175 229
rect 119 157 130 191
rect 164 157 175 191
rect 119 119 175 157
rect 119 85 130 119
rect 164 85 175 119
rect 119 36 175 85
rect 205 983 261 1036
rect 205 949 216 983
rect 250 949 261 983
rect 205 911 261 949
rect 205 877 216 911
rect 250 877 261 911
rect 205 839 261 877
rect 205 805 216 839
rect 250 805 261 839
rect 205 767 261 805
rect 205 733 216 767
rect 250 733 261 767
rect 205 695 261 733
rect 205 661 216 695
rect 250 661 261 695
rect 205 623 261 661
rect 205 589 216 623
rect 250 589 261 623
rect 205 551 261 589
rect 205 517 216 551
rect 250 517 261 551
rect 205 479 261 517
rect 205 445 216 479
rect 250 445 261 479
rect 205 407 261 445
rect 205 373 216 407
rect 250 373 261 407
rect 205 335 261 373
rect 205 301 216 335
rect 250 301 261 335
rect 205 263 261 301
rect 205 229 216 263
rect 250 229 261 263
rect 205 191 261 229
rect 205 157 216 191
rect 250 157 261 191
rect 205 119 261 157
rect 205 85 216 119
rect 250 85 261 119
rect 205 36 261 85
rect 291 983 347 1036
rect 291 949 302 983
rect 336 949 347 983
rect 291 911 347 949
rect 291 877 302 911
rect 336 877 347 911
rect 291 839 347 877
rect 291 805 302 839
rect 336 805 347 839
rect 291 767 347 805
rect 291 733 302 767
rect 336 733 347 767
rect 291 695 347 733
rect 291 661 302 695
rect 336 661 347 695
rect 291 623 347 661
rect 291 589 302 623
rect 336 589 347 623
rect 291 551 347 589
rect 291 517 302 551
rect 336 517 347 551
rect 291 479 347 517
rect 291 445 302 479
rect 336 445 347 479
rect 291 407 347 445
rect 291 373 302 407
rect 336 373 347 407
rect 291 335 347 373
rect 291 301 302 335
rect 336 301 347 335
rect 291 263 347 301
rect 291 229 302 263
rect 336 229 347 263
rect 291 191 347 229
rect 291 157 302 191
rect 336 157 347 191
rect 291 119 347 157
rect 291 85 302 119
rect 336 85 347 119
rect 291 36 347 85
rect 377 983 430 1036
rect 377 949 388 983
rect 422 949 430 983
rect 377 911 430 949
rect 377 877 388 911
rect 422 877 430 911
rect 377 839 430 877
rect 377 805 388 839
rect 422 805 430 839
rect 377 767 430 805
rect 377 733 388 767
rect 422 733 430 767
rect 377 695 430 733
rect 377 661 388 695
rect 422 661 430 695
rect 377 623 430 661
rect 377 589 388 623
rect 422 589 430 623
rect 377 551 430 589
rect 377 517 388 551
rect 422 517 430 551
rect 377 479 430 517
rect 377 445 388 479
rect 422 445 430 479
rect 377 407 430 445
rect 377 373 388 407
rect 422 373 430 407
rect 377 335 430 373
rect 377 301 388 335
rect 422 301 430 335
rect 377 263 430 301
rect 377 229 388 263
rect 422 229 430 263
rect 377 191 430 229
rect 377 157 388 191
rect 422 157 430 191
rect 377 119 430 157
rect 377 85 388 119
rect 422 85 430 119
rect 377 36 430 85
<< pdiffc >>
rect 44 949 78 983
rect 44 877 78 911
rect 44 805 78 839
rect 44 733 78 767
rect 44 661 78 695
rect 44 589 78 623
rect 44 517 78 551
rect 44 445 78 479
rect 44 373 78 407
rect 44 301 78 335
rect 44 229 78 263
rect 44 157 78 191
rect 44 85 78 119
rect 130 949 164 983
rect 130 877 164 911
rect 130 805 164 839
rect 130 733 164 767
rect 130 661 164 695
rect 130 589 164 623
rect 130 517 164 551
rect 130 445 164 479
rect 130 373 164 407
rect 130 301 164 335
rect 130 229 164 263
rect 130 157 164 191
rect 130 85 164 119
rect 216 949 250 983
rect 216 877 250 911
rect 216 805 250 839
rect 216 733 250 767
rect 216 661 250 695
rect 216 589 250 623
rect 216 517 250 551
rect 216 445 250 479
rect 216 373 250 407
rect 216 301 250 335
rect 216 229 250 263
rect 216 157 250 191
rect 216 85 250 119
rect 302 949 336 983
rect 302 877 336 911
rect 302 805 336 839
rect 302 733 336 767
rect 302 661 336 695
rect 302 589 336 623
rect 302 517 336 551
rect 302 445 336 479
rect 302 373 336 407
rect 302 301 336 335
rect 302 229 336 263
rect 302 157 336 191
rect 302 85 336 119
rect 388 949 422 983
rect 388 877 422 911
rect 388 805 422 839
rect 388 733 422 767
rect 388 661 422 695
rect 388 589 422 623
rect 388 517 422 551
rect 388 445 422 479
rect 388 373 422 407
rect 388 301 422 335
rect 388 229 422 263
rect 388 157 422 191
rect 388 85 422 119
<< poly >>
rect 89 1119 377 1135
rect 89 1085 114 1119
rect 148 1085 182 1119
rect 216 1085 250 1119
rect 284 1085 318 1119
rect 352 1085 377 1119
rect 89 1062 377 1085
rect 89 1036 119 1062
rect 175 1036 205 1062
rect 261 1036 291 1062
rect 347 1036 377 1062
rect 89 10 119 36
rect 175 10 205 36
rect 261 10 291 36
rect 347 10 377 36
<< polycont >>
rect 114 1085 148 1119
rect 182 1085 216 1119
rect 250 1085 284 1119
rect 318 1085 352 1119
<< locali >>
rect 98 1119 368 1135
rect 98 1085 108 1119
rect 148 1085 180 1119
rect 216 1085 250 1119
rect 286 1085 318 1119
rect 358 1085 368 1119
rect 98 1067 368 1085
rect 44 983 78 1021
rect 44 911 78 949
rect 44 839 78 877
rect 44 767 78 805
rect 44 695 78 733
rect 44 623 78 661
rect 44 551 78 589
rect 44 479 78 517
rect 44 407 78 445
rect 44 335 78 373
rect 44 263 78 301
rect 44 191 78 229
rect 44 119 78 157
rect 44 51 78 85
rect 130 983 164 1021
rect 130 911 164 949
rect 130 839 164 877
rect 130 767 164 805
rect 130 695 164 733
rect 130 623 164 661
rect 130 551 164 589
rect 130 479 164 517
rect 130 407 164 445
rect 130 335 164 373
rect 130 263 164 301
rect 130 191 164 229
rect 130 119 164 157
rect 130 51 164 85
rect 216 983 250 1021
rect 216 911 250 949
rect 216 839 250 877
rect 216 767 250 805
rect 216 695 250 733
rect 216 623 250 661
rect 216 551 250 589
rect 216 479 250 517
rect 216 407 250 445
rect 216 335 250 373
rect 216 263 250 301
rect 216 191 250 229
rect 216 119 250 157
rect 216 51 250 85
rect 302 983 336 1021
rect 302 911 336 949
rect 302 839 336 877
rect 302 767 336 805
rect 302 695 336 733
rect 302 623 336 661
rect 302 551 336 589
rect 302 479 336 517
rect 302 407 336 445
rect 302 335 336 373
rect 302 263 336 301
rect 302 191 336 229
rect 302 119 336 157
rect 302 51 336 85
rect 388 983 422 1021
rect 388 911 422 949
rect 388 839 422 877
rect 388 767 422 805
rect 388 695 422 733
rect 388 623 422 661
rect 388 551 422 589
rect 388 479 422 517
rect 388 407 422 445
rect 388 335 422 373
rect 388 263 422 301
rect 388 191 422 229
rect 388 119 422 157
rect 388 51 422 85
<< viali >>
rect 108 1085 114 1119
rect 114 1085 142 1119
rect 180 1085 182 1119
rect 182 1085 214 1119
rect 252 1085 284 1119
rect 284 1085 286 1119
rect 324 1085 352 1119
rect 352 1085 358 1119
rect 44 949 78 983
rect 44 877 78 911
rect 44 805 78 839
rect 44 733 78 767
rect 44 661 78 695
rect 44 589 78 623
rect 44 517 78 551
rect 44 445 78 479
rect 44 373 78 407
rect 44 301 78 335
rect 44 229 78 263
rect 44 157 78 191
rect 44 85 78 119
rect 130 949 164 983
rect 130 877 164 911
rect 130 805 164 839
rect 130 733 164 767
rect 130 661 164 695
rect 130 589 164 623
rect 130 517 164 551
rect 130 445 164 479
rect 130 373 164 407
rect 130 301 164 335
rect 130 229 164 263
rect 130 157 164 191
rect 130 85 164 119
rect 216 949 250 983
rect 216 877 250 911
rect 216 805 250 839
rect 216 733 250 767
rect 216 661 250 695
rect 216 589 250 623
rect 216 517 250 551
rect 216 445 250 479
rect 216 373 250 407
rect 216 301 250 335
rect 216 229 250 263
rect 216 157 250 191
rect 216 85 250 119
rect 302 949 336 983
rect 302 877 336 911
rect 302 805 336 839
rect 302 733 336 767
rect 302 661 336 695
rect 302 589 336 623
rect 302 517 336 551
rect 302 445 336 479
rect 302 373 336 407
rect 302 301 336 335
rect 302 229 336 263
rect 302 157 336 191
rect 302 85 336 119
rect 388 949 422 983
rect 388 877 422 911
rect 388 805 422 839
rect 388 733 422 767
rect 388 661 422 695
rect 388 589 422 623
rect 388 517 422 551
rect 388 445 422 479
rect 388 373 422 407
rect 388 301 422 335
rect 388 229 422 263
rect 388 157 422 191
rect 388 85 422 119
<< metal1 >>
rect 96 1119 370 1131
rect 96 1085 108 1119
rect 142 1085 180 1119
rect 214 1085 252 1119
rect 286 1085 324 1119
rect 358 1085 370 1119
rect 96 1073 370 1085
rect 38 983 84 1021
rect 38 949 44 983
rect 78 949 84 983
rect 38 911 84 949
rect 38 877 44 911
rect 78 877 84 911
rect 38 839 84 877
rect 38 805 44 839
rect 78 805 84 839
rect 38 767 84 805
rect 38 733 44 767
rect 78 733 84 767
rect 38 695 84 733
rect 38 661 44 695
rect 78 661 84 695
rect 38 623 84 661
rect 38 589 44 623
rect 78 589 84 623
rect 38 551 84 589
rect 38 517 44 551
rect 78 517 84 551
rect 38 479 84 517
rect 38 445 44 479
rect 78 445 84 479
rect 38 407 84 445
rect 38 373 44 407
rect 78 373 84 407
rect 38 335 84 373
rect 38 301 44 335
rect 78 301 84 335
rect 38 263 84 301
rect 38 229 44 263
rect 78 229 84 263
rect 38 191 84 229
rect 38 157 44 191
rect 78 157 84 191
rect 38 119 84 157
rect 38 85 44 119
rect 78 85 84 119
rect 38 -45 84 85
rect 121 1010 173 1021
rect 121 949 130 958
rect 164 949 173 958
rect 121 946 173 949
rect 121 877 130 894
rect 164 877 173 894
rect 121 839 173 877
rect 121 805 130 839
rect 164 805 173 839
rect 121 767 173 805
rect 121 733 130 767
rect 164 733 173 767
rect 121 695 173 733
rect 121 661 130 695
rect 164 661 173 695
rect 121 623 173 661
rect 121 589 130 623
rect 164 589 173 623
rect 121 551 173 589
rect 121 517 130 551
rect 164 517 173 551
rect 121 479 173 517
rect 121 445 130 479
rect 164 445 173 479
rect 121 407 173 445
rect 121 373 130 407
rect 164 373 173 407
rect 121 335 173 373
rect 121 301 130 335
rect 164 301 173 335
rect 121 263 173 301
rect 121 229 130 263
rect 164 229 173 263
rect 121 191 173 229
rect 121 157 130 191
rect 164 157 173 191
rect 121 119 173 157
rect 121 85 130 119
rect 164 85 173 119
rect 121 51 173 85
rect 210 983 256 1021
rect 210 949 216 983
rect 250 949 256 983
rect 210 911 256 949
rect 210 877 216 911
rect 250 877 256 911
rect 210 839 256 877
rect 210 805 216 839
rect 250 805 256 839
rect 210 767 256 805
rect 210 733 216 767
rect 250 733 256 767
rect 210 695 256 733
rect 210 661 216 695
rect 250 661 256 695
rect 210 623 256 661
rect 210 589 216 623
rect 250 589 256 623
rect 210 551 256 589
rect 210 517 216 551
rect 250 517 256 551
rect 210 479 256 517
rect 210 445 216 479
rect 250 445 256 479
rect 210 407 256 445
rect 210 373 216 407
rect 250 373 256 407
rect 210 335 256 373
rect 210 301 216 335
rect 250 301 256 335
rect 210 263 256 301
rect 210 229 216 263
rect 250 229 256 263
rect 210 191 256 229
rect 210 157 216 191
rect 250 157 256 191
rect 210 119 256 157
rect 210 85 216 119
rect 250 85 256 119
rect 210 -45 256 85
rect 293 1010 345 1021
rect 293 949 302 958
rect 336 949 345 958
rect 293 946 345 949
rect 293 877 302 894
rect 336 877 345 894
rect 293 839 345 877
rect 293 805 302 839
rect 336 805 345 839
rect 293 767 345 805
rect 293 733 302 767
rect 336 733 345 767
rect 293 695 345 733
rect 293 661 302 695
rect 336 661 345 695
rect 293 623 345 661
rect 293 589 302 623
rect 336 589 345 623
rect 293 551 345 589
rect 293 517 302 551
rect 336 517 345 551
rect 293 479 345 517
rect 293 445 302 479
rect 336 445 345 479
rect 293 407 345 445
rect 293 373 302 407
rect 336 373 345 407
rect 293 335 345 373
rect 293 301 302 335
rect 336 301 345 335
rect 293 263 345 301
rect 293 229 302 263
rect 336 229 345 263
rect 293 191 345 229
rect 293 157 302 191
rect 336 157 345 191
rect 293 119 345 157
rect 293 85 302 119
rect 336 85 345 119
rect 293 51 345 85
rect 382 983 428 1021
rect 382 949 388 983
rect 422 949 428 983
rect 382 911 428 949
rect 382 877 388 911
rect 422 877 428 911
rect 382 839 428 877
rect 382 805 388 839
rect 422 805 428 839
rect 382 767 428 805
rect 382 733 388 767
rect 422 733 428 767
rect 382 695 428 733
rect 382 661 388 695
rect 422 661 428 695
rect 382 623 428 661
rect 382 589 388 623
rect 422 589 428 623
rect 382 551 428 589
rect 382 517 388 551
rect 422 517 428 551
rect 382 479 428 517
rect 382 445 388 479
rect 422 445 428 479
rect 382 407 428 445
rect 382 373 388 407
rect 422 373 428 407
rect 382 335 428 373
rect 382 301 388 335
rect 422 301 428 335
rect 382 263 428 301
rect 382 229 388 263
rect 422 229 428 263
rect 382 191 428 229
rect 382 157 388 191
rect 422 157 428 191
rect 382 119 428 157
rect 382 85 388 119
rect 422 85 428 119
rect 382 -45 428 85
rect 38 -97 428 -45
<< via1 >>
rect 121 983 173 1010
rect 121 958 130 983
rect 130 958 164 983
rect 164 958 173 983
rect 121 911 173 946
rect 121 894 130 911
rect 130 894 164 911
rect 164 894 173 911
rect 293 983 345 1010
rect 293 958 302 983
rect 302 958 336 983
rect 336 958 345 983
rect 293 911 345 946
rect 293 894 302 911
rect 302 894 336 911
rect 336 894 345 911
<< metal2 >>
rect 114 1020 180 1029
rect 114 964 119 1020
rect 175 964 180 1020
rect 114 958 121 964
rect 173 958 180 964
rect 114 946 180 958
rect 114 940 121 946
rect 173 940 180 946
rect 114 884 119 940
rect 175 884 180 940
rect 114 875 180 884
rect 286 1020 352 1029
rect 286 964 291 1020
rect 347 964 352 1020
rect 286 958 293 964
rect 345 958 352 964
rect 286 946 352 958
rect 286 940 293 946
rect 345 940 352 946
rect 286 884 291 940
rect 347 884 352 940
rect 286 875 352 884
<< via2 >>
rect 119 1010 175 1020
rect 119 964 121 1010
rect 121 964 173 1010
rect 173 964 175 1010
rect 119 894 121 940
rect 121 894 173 940
rect 173 894 175 940
rect 119 884 175 894
rect 291 1010 347 1020
rect 291 964 293 1010
rect 293 964 345 1010
rect 345 964 347 1010
rect 291 894 293 940
rect 293 894 345 940
rect 345 894 347 940
rect 291 884 347 894
<< metal3 >>
rect 114 1020 352 1029
rect 114 964 119 1020
rect 175 964 291 1020
rect 347 964 352 1020
rect 114 963 352 964
rect 114 940 180 963
rect 114 884 119 940
rect 175 884 180 940
rect 114 875 180 884
rect 286 940 352 963
rect 286 884 291 940
rect 347 884 352 940
rect 286 875 352 884
<< labels >>
flabel metal3 s 114 963 352 1029 0 FreeSans 400 0 0 0 DRAIN
port 2 nsew
flabel metal1 s 96 1073 370 1131 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel metal1 s 38 -97 428 -45 0 FreeSans 400 0 0 0 SOURCE
port 4 nsew
flabel nwell s 84 1063 88 1070 0 FreeSans 400 0 0 0 BULK
port 5 nsew
<< properties >>
string GDS_END 9155000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9141280
string path 0.950 -1.775 10.700 -1.775 
<< end >>
