magic
tech sky130A
timestamp 1704896540
<< viali >>
rect 0 0 53 233
<< metal1 >>
rect -6 233 59 236
rect -6 0 0 233
rect 53 0 59 233
rect -6 -3 59 0
<< properties >>
string GDS_END 87998014
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87996986
<< end >>
