magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 14 0 134 118
rect 4166 0 4367 118
rect 4286 -8 4367 0
rect 2654 -134 2774 -8
rect 1774 -252 1894 -134
rect 2526 -252 2774 -134
rect 2526 -260 2574 -252
rect 2446 -378 2574 -260
rect 3406 -378 3654 -8
rect 4286 -126 4446 -8
rect 4286 -378 4406 -126
<< mvndiff >>
rect 40 76 108 92
rect 40 42 48 76
rect 82 42 108 76
rect 40 26 108 42
rect 4192 76 4341 92
rect 4192 42 4218 76
rect 4252 42 4341 76
rect 4192 26 4341 42
rect 2680 -50 2748 -34
rect 2680 -84 2688 -50
rect 2722 -84 2748 -50
rect 2680 -100 2748 -84
rect 3432 -50 3500 -34
rect 3432 -84 3458 -50
rect 3492 -84 3500 -50
rect 3432 -100 3500 -84
rect 3560 -50 3628 -34
rect 3560 -84 3568 -50
rect 3602 -84 3628 -50
rect 3560 -100 3628 -84
rect 4312 -50 4420 -34
rect 4312 -84 4338 -50
rect 4372 -84 4420 -50
rect 4312 -100 4420 -84
rect 1800 -176 1868 -160
rect 1800 -210 1808 -176
rect 1842 -210 1868 -176
rect 1800 -226 1868 -210
rect 2552 -176 2620 -160
rect 2552 -210 2578 -176
rect 2612 -210 2620 -176
rect 2552 -226 2620 -210
rect 2680 -176 2748 -160
rect 2680 -210 2688 -176
rect 2722 -210 2748 -176
rect 2680 -226 2748 -210
rect 3432 -176 3500 -160
rect 3432 -210 3458 -176
rect 3492 -210 3500 -176
rect 3432 -226 3500 -210
rect 3560 -176 3628 -160
rect 3560 -210 3568 -176
rect 3602 -210 3628 -176
rect 3560 -226 3628 -210
rect 4312 -176 4380 -160
rect 4312 -210 4338 -176
rect 4372 -210 4380 -176
rect 4312 -226 4380 -210
rect 2472 -302 2548 -286
rect 2472 -336 2488 -302
rect 2522 -336 2548 -302
rect 2472 -352 2548 -336
rect 3432 -302 3500 -286
rect 3432 -336 3458 -302
rect 3492 -336 3500 -302
rect 3432 -352 3500 -336
rect 3560 -302 3628 -286
rect 3560 -336 3568 -302
rect 3602 -336 3628 -302
rect 3560 -352 3628 -336
rect 4312 -302 4380 -286
rect 4312 -336 4338 -302
rect 4372 -336 4380 -302
rect 4312 -352 4380 -336
<< mvndiffc >>
rect 48 42 82 76
rect 4218 42 4252 76
rect 2688 -84 2722 -50
rect 3458 -84 3492 -50
rect 3568 -84 3602 -50
rect 4338 -84 4372 -50
rect 1808 -210 1842 -176
rect 2578 -210 2612 -176
rect 2688 -210 2722 -176
rect 3458 -210 3492 -176
rect 3568 -210 3602 -176
rect 4338 -210 4372 -176
rect 2488 -336 2522 -302
rect 3458 -336 3492 -302
rect 3568 -336 3602 -302
rect 4338 -336 4372 -302
<< locali >>
rect 48 76 178 92
rect 94 42 132 76
rect 166 42 178 76
rect 48 26 178 42
rect 4122 76 4252 92
rect 4122 42 4134 76
rect 4168 42 4206 76
rect 4122 26 4252 42
rect 2688 -50 2818 -34
rect 2734 -84 2772 -50
rect 2806 -84 2818 -50
rect 2688 -100 2818 -84
rect 3362 -50 3492 -34
rect 3362 -84 3374 -50
rect 3408 -84 3446 -50
rect 3362 -100 3492 -84
rect 3568 -50 3698 -34
rect 3614 -84 3652 -50
rect 3686 -84 3698 -50
rect 3568 -100 3698 -84
rect 4242 -50 4372 -34
rect 4242 -84 4254 -50
rect 4288 -84 4326 -50
rect 4242 -100 4372 -84
rect 1808 -176 1938 -160
rect 2510 -176 2612 -160
rect 1854 -210 1892 -176
rect 1926 -210 1938 -176
rect 2528 -210 2566 -176
rect 1808 -226 1938 -210
rect 2510 -226 2612 -210
rect 2688 -176 2722 -160
rect 3362 -176 3492 -160
rect 2734 -210 2772 -176
rect 3362 -210 3374 -176
rect 3408 -210 3446 -176
rect 2688 -226 2722 -210
rect 3362 -226 3492 -210
rect 3568 -176 3698 -160
rect 4270 -176 4400 -160
rect 3614 -210 3652 -176
rect 3686 -210 3698 -176
rect 4288 -210 4326 -176
rect 4372 -210 4400 -176
rect 3568 -226 3698 -210
rect 4270 -226 4400 -210
rect 2460 -302 2590 -286
rect 3362 -302 3492 -286
rect 2460 -336 2488 -302
rect 2534 -336 2572 -302
rect 3362 -336 3374 -302
rect 3408 -336 3446 -302
rect 2460 -352 2590 -336
rect 3362 -352 3492 -336
rect 3568 -302 3698 -286
rect 3614 -336 3652 -302
rect 3686 -336 3698 -302
rect 3568 -352 3698 -336
rect 4242 -302 4372 -286
rect 4242 -336 4254 -302
rect 4288 -336 4326 -302
rect 4242 -352 4372 -336
<< viali >>
rect 60 42 82 76
rect 82 42 94 76
rect 132 42 166 76
rect 4134 42 4168 76
rect 4206 42 4218 76
rect 4218 42 4240 76
rect 2700 -84 2722 -50
rect 2722 -84 2734 -50
rect 2772 -84 2806 -50
rect 3374 -84 3408 -50
rect 3446 -84 3458 -50
rect 3458 -84 3480 -50
rect 3580 -84 3602 -50
rect 3602 -84 3614 -50
rect 3652 -84 3686 -50
rect 4254 -84 4288 -50
rect 4326 -84 4338 -50
rect 4338 -84 4360 -50
rect 1820 -210 1842 -176
rect 1842 -210 1854 -176
rect 1892 -210 1926 -176
rect 2494 -210 2528 -176
rect 2566 -210 2578 -176
rect 2578 -210 2600 -176
rect 2700 -210 2722 -176
rect 2722 -210 2734 -176
rect 2772 -210 2806 -176
rect 3374 -210 3408 -176
rect 3446 -210 3458 -176
rect 3458 -210 3480 -176
rect 3580 -210 3602 -176
rect 3602 -210 3614 -176
rect 3652 -210 3686 -176
rect 4254 -210 4288 -176
rect 4326 -210 4338 -176
rect 4338 -210 4360 -176
rect 2500 -336 2522 -302
rect 2522 -336 2534 -302
rect 2572 -336 2606 -302
rect 3374 -336 3408 -302
rect 3446 -336 3458 -302
rect 3458 -336 3480 -302
rect 3580 -336 3602 -302
rect 3602 -336 3614 -302
rect 3652 -336 3686 -302
rect 4254 -336 4288 -302
rect 4326 -336 4338 -302
rect 4338 -336 4360 -302
<< metal1 >>
rect 54 80 172 88
tri 172 80 180 88 sw
tri 4120 80 4128 88 se
rect 4128 80 4246 88
rect 54 76 2130 80
rect 54 42 60 76
rect 94 42 132 76
rect 166 42 2130 76
rect 54 38 2130 42
rect 2131 39 2132 79
rect 2168 39 2169 79
rect 2170 76 4246 80
rect 2170 42 4134 76
rect 4168 42 4206 76
rect 4240 42 4246 76
rect 2170 38 4246 42
rect 54 30 172 38
tri 172 30 180 38 nw
tri 4103 30 4111 38 ne
rect 4111 30 4246 38
tri 4111 13 4128 30 ne
tri 4111 -38 4128 -21 se
rect 4128 -38 4246 30
tri 4246 -38 4271 -13 sw
tri 2687 -45 2694 -38 se
rect 2694 -45 2812 -38
rect 2003 -46 2812 -45
tri 2812 -46 2820 -38 sw
tri 3360 -46 3368 -38 se
rect 3368 -46 3692 -38
tri 3692 -46 3700 -38 sw
tri 4103 -46 4111 -38 se
rect 4111 -46 4366 -38
rect 2003 -50 3070 -46
rect 3072 -47 3108 -46
rect 2003 -84 2700 -50
rect 2734 -84 2772 -50
rect 2806 -84 3070 -50
rect 2003 -87 3070 -84
rect 3071 -87 3109 -47
rect 3110 -50 3950 -46
rect 3952 -47 3988 -46
rect 3110 -84 3374 -50
rect 3408 -84 3446 -50
rect 3480 -84 3580 -50
rect 3614 -84 3652 -50
rect 3686 -84 3950 -50
tri 2003 -113 2029 -87 ne
tri 2012 -164 2029 -147 se
rect 2029 -164 2155 -87
tri 2155 -113 2181 -87 nw
tri 2685 -96 2694 -87 ne
rect 2694 -88 3070 -87
rect 3072 -88 3108 -87
rect 3110 -88 3950 -84
rect 3951 -87 3989 -47
rect 3990 -50 4366 -46
rect 3990 -84 4254 -50
rect 4288 -84 4326 -50
rect 4360 -84 4366 -50
rect 3952 -88 3988 -87
rect 3990 -88 4366 -84
rect 2694 -96 2812 -88
tri 2812 -96 2820 -88 nw
tri 3360 -96 3368 -88 ne
rect 3368 -96 3692 -88
tri 3692 -96 3700 -88 nw
tri 4240 -96 4248 -88 ne
rect 4248 -96 4366 -88
rect 1814 -172 1932 -164
tri 1932 -172 1940 -164 sw
tri 2004 -172 2012 -164 se
rect 2012 -172 2155 -164
tri 2155 -172 2180 -147 sw
tri 2480 -172 2488 -164 se
rect 2488 -172 2812 -164
tri 2812 -172 2820 -164 sw
tri 3360 -172 3368 -164 se
rect 3368 -172 3692 -164
tri 3692 -172 3700 -164 sw
tri 4240 -172 4248 -164 se
rect 4248 -172 4366 -164
rect 1814 -176 2233 -172
rect 2235 -173 2271 -172
rect 1814 -210 1820 -176
rect 1854 -210 1892 -176
rect 1926 -210 2233 -176
rect 1814 -214 2233 -210
rect 2234 -213 2272 -173
rect 2273 -176 3070 -172
rect 3072 -173 3108 -172
rect 2273 -210 2494 -176
rect 2528 -210 2566 -176
rect 2600 -210 2700 -176
rect 2734 -210 2772 -176
rect 2806 -210 3070 -176
rect 2235 -214 2271 -213
rect 2273 -214 3070 -210
rect 3071 -213 3109 -173
rect 3110 -176 3950 -172
rect 3952 -173 3988 -172
rect 3110 -210 3374 -176
rect 3408 -210 3446 -176
rect 3480 -210 3580 -176
rect 3614 -210 3652 -176
rect 3686 -210 3950 -176
rect 3072 -214 3108 -213
rect 3110 -214 3950 -210
rect 3951 -213 3989 -173
rect 3990 -176 4366 -172
rect 3990 -210 4254 -176
rect 4288 -210 4326 -176
rect 4360 -210 4366 -176
rect 3952 -214 3988 -213
rect 3990 -214 4366 -210
rect 1814 -222 1932 -214
tri 1932 -222 1940 -214 nw
tri 2480 -222 2488 -214 ne
rect 2488 -222 2812 -214
tri 2812 -222 2820 -214 nw
tri 3360 -222 3368 -214 ne
rect 3368 -222 3692 -214
tri 3692 -222 3700 -214 nw
tri 4223 -222 4231 -214 ne
rect 4231 -222 4366 -214
tri 4231 -239 4248 -222 ne
tri 4231 -290 4248 -273 se
rect 4248 -290 4366 -222
rect 2494 -298 2612 -290
tri 2612 -298 2620 -290 sw
tri 3360 -298 3368 -290 se
rect 3368 -298 3692 -290
tri 3692 -298 3700 -290 sw
tri 4223 -298 4231 -290 se
rect 4231 -298 4366 -290
rect 2494 -302 2970 -298
rect 2972 -299 3008 -298
rect 2494 -336 2500 -302
rect 2534 -336 2572 -302
rect 2606 -336 2970 -302
rect 2494 -340 2970 -336
rect 2971 -339 3009 -299
rect 3010 -302 3950 -298
rect 3952 -299 3988 -298
rect 3010 -336 3374 -302
rect 3408 -336 3446 -302
rect 3480 -336 3580 -302
rect 3614 -336 3652 -302
rect 3686 -336 3950 -302
rect 2972 -340 3008 -339
rect 3010 -340 3950 -336
rect 3951 -339 3989 -299
rect 3990 -302 4366 -298
rect 3990 -336 4254 -302
rect 4288 -336 4326 -302
rect 4360 -336 4366 -302
rect 3952 -340 3988 -339
rect 3990 -340 4366 -336
rect 2494 -348 2612 -340
tri 2612 -348 2620 -340 nw
tri 3360 -348 3368 -340 ne
rect 3368 -348 3692 -340
tri 3692 -348 3700 -340 nw
tri 4240 -348 4248 -340 ne
rect 4248 -348 4366 -340
<< rmetal1 >>
rect 2130 79 2132 80
rect 2130 39 2131 79
rect 2130 38 2132 39
rect 2168 79 2170 80
rect 2169 39 2170 79
rect 2168 38 2170 39
rect 3070 -47 3072 -46
rect 3108 -47 3110 -46
rect 3070 -87 3071 -47
rect 3109 -87 3110 -47
rect 3950 -47 3952 -46
rect 3988 -47 3990 -46
rect 3070 -88 3072 -87
rect 3108 -88 3110 -87
rect 3950 -87 3951 -47
rect 3989 -87 3990 -47
rect 3950 -88 3952 -87
rect 3988 -88 3990 -87
rect 2233 -173 2235 -172
rect 2271 -173 2273 -172
rect 2233 -213 2234 -173
rect 2272 -213 2273 -173
rect 3070 -173 3072 -172
rect 3108 -173 3110 -172
rect 2233 -214 2235 -213
rect 2271 -214 2273 -213
rect 3070 -213 3071 -173
rect 3109 -213 3110 -173
rect 3950 -173 3952 -172
rect 3988 -173 3990 -172
rect 3070 -214 3072 -213
rect 3108 -214 3110 -213
rect 3950 -213 3951 -173
rect 3989 -213 3990 -173
rect 3950 -214 3952 -213
rect 3988 -214 3990 -213
rect 2970 -299 2972 -298
rect 3008 -299 3010 -298
rect 2970 -339 2971 -299
rect 3009 -339 3010 -299
rect 3950 -299 3952 -298
rect 3988 -299 3990 -298
rect 2970 -340 2972 -339
rect 3008 -340 3010 -339
rect 3950 -339 3951 -299
rect 3989 -339 3990 -299
rect 3950 -340 3952 -339
rect 3988 -340 3990 -339
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 3500 0 1 -348
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform -1 0 4380 0 1 -348
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1704896540
transform -1 0 4380 0 1 -222
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1704896540
transform -1 0 4380 0 1 -96
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1704896540
transform -1 0 3500 0 1 -96
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1704896540
transform -1 0 2620 0 1 -222
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_6
timestamp 1704896540
transform -1 0 3500 0 1 -222
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_7
timestamp 1704896540
transform -1 0 4260 0 1 30
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_8
timestamp 1704896540
transform 1 0 2480 0 1 -348
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_9
timestamp 1704896540
transform 1 0 3560 0 1 -348
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_10
timestamp 1704896540
transform 1 0 3560 0 1 -96
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_11
timestamp 1704896540
transform 1 0 2680 0 1 -96
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_12
timestamp 1704896540
transform 1 0 1800 0 1 -222
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_13
timestamp 1704896540
transform 1 0 2680 0 1 -222
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_14
timestamp 1704896540
transform 1 0 3560 0 1 -222
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_15
timestamp 1704896540
transform 1 0 40 0 1 30
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 1 2500 1 0 -336
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 0 1 3580 1 0 -336
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 0 1 60 1 0 42
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 0 1 3580 1 0 -84
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform 0 1 2700 1 0 -84
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform 0 1 1820 1 0 -210
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1704896540
transform 0 1 2700 1 0 -210
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1704896540
transform 0 1 3580 1 0 -210
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1704896540
transform 0 -1 3480 1 0 -336
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1704896540
transform 0 -1 4360 1 0 -336
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1704896540
transform 0 -1 4360 1 0 -210
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1704896540
transform 0 -1 4240 1 0 42
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1704896540
transform 0 -1 4360 1 0 -84
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1704896540
transform 0 -1 3480 1 0 -84
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1704896540
transform 0 -1 2600 1 0 -210
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1704896540
transform 0 -1 3480 1 0 -210
box 0 0 1 1
use nDFres_CDNS_524688791851259  nDFres_CDNS_524688791851259_0
timestamp 1704896540
transform -1 0 3390 0 -1 -286
box -68 -26 868 92
use nDFres_CDNS_524688791851280  nDFres_CDNS_524688791851280_0
timestamp 1704896540
transform -1 0 4270 0 -1 -286
box -68 -26 668 92
use nDFres_CDNS_524688791851280  nDFres_CDNS_524688791851280_1
timestamp 1704896540
transform -1 0 3390 0 -1 -34
box -68 -26 668 92
use nDFres_CDNS_524688791851280  nDFres_CDNS_524688791851280_2
timestamp 1704896540
transform -1 0 4270 0 -1 -34
box -68 -26 668 92
use nDFres_CDNS_524688791851280  nDFres_CDNS_524688791851280_3
timestamp 1704896540
transform 1 0 3670 0 -1 -160
box -68 -26 668 92
use nDFres_CDNS_524688791851280  nDFres_CDNS_524688791851280_4
timestamp 1704896540
transform 1 0 2790 0 -1 -160
box -68 -26 668 92
use nDFres_CDNS_524688791851280  nDFres_CDNS_524688791851280_5
timestamp 1704896540
transform 1 0 1910 0 -1 -160
box -68 -26 668 92
use nDFres_CDNS_524688791851281  nDFres_CDNS_524688791851281_0
timestamp 1704896540
transform 1 0 150 0 -1 92
box -68 -26 4068 92
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_0
timestamp 1704896540
transform 1 0 2078 0 1 38
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_0
timestamp 1704896540
transform -1 0 3062 0 1 -340
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_1
timestamp 1704896540
transform -1 0 4042 0 1 -340
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_2
timestamp 1704896540
transform -1 0 3162 0 1 -88
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_3
timestamp 1704896540
transform -1 0 4042 0 1 -88
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_4
timestamp 1704896540
transform 1 0 3898 0 1 -214
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_5
timestamp 1704896540
transform 1 0 3018 0 1 -214
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_6
timestamp 1704896540
transform 1 0 2181 0 1 -214
box 0 0 1 1
<< labels >>
flabel metal1 s 2494 -348 2534 -290 0 FreeSans 200 0 0 0 r1
port 1 nsew
flabel metal1 s 54 30 94 88 0 FreeSans 200 0 0 0 r0
port 2 nsew
<< properties >>
string GDS_END 86213420
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86205932
<< end >>
