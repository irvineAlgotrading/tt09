magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 536 3883 4076 4051
rect 1224 3242 4076 3883
rect 536 2810 4076 3242
<< pwell >>
rect 867 2495 1480 2535
rect 1726 2495 2378 2502
rect 867 2449 2378 2495
rect 1616 2251 2378 2449
rect 1149 1993 2378 2251
rect 1616 1795 2378 1993
rect 2722 2495 3774 2502
rect 2722 2082 3890 2495
rect 2722 1932 3774 2082
rect 1726 1776 2378 1795
rect 546 175 3098 1227
rect 568 65 3065 175
<< mvnmos >>
rect 1752 2323 2352 2423
rect 2748 2323 3748 2423
rect 1175 2072 1475 2172
rect 1752 2167 2352 2267
rect 2748 2167 3748 2267
rect 1752 2011 2352 2111
rect 2748 2011 3748 2111
rect 1752 1855 2352 1955
rect 625 201 725 1201
rect 781 201 881 1201
rect 937 201 1037 1201
rect 1093 201 1193 1201
rect 1249 201 1349 1201
rect 1405 201 1505 1201
rect 1561 201 1661 1201
rect 1717 201 1817 1201
rect 1983 201 2083 1201
rect 2139 201 2239 1201
rect 2295 201 2395 1201
rect 2451 201 2551 1201
rect 2607 201 2707 1201
rect 2763 201 2863 1201
rect 2919 201 3019 1201
<< mvpmos >>
rect 655 2876 755 3176
rect 811 2876 911 3176
rect 1077 2876 1177 3176
rect 1343 2876 1443 3876
rect 1499 2876 1599 3876
rect 1655 2876 1755 3876
rect 1811 2876 1911 3876
rect 2077 2876 2177 3876
rect 2233 2876 2333 3876
rect 2389 2876 2489 3876
rect 2545 2876 2645 3876
rect 2811 2876 2911 3876
rect 2967 2876 3067 3876
rect 3233 2876 3333 3876
rect 3389 2876 3489 3876
rect 3545 2876 3645 3876
rect 3701 2876 3801 3876
rect 3857 2876 3957 3876
<< mvndiff >>
rect 1752 2468 2352 2476
rect 1752 2434 1764 2468
rect 1798 2434 1832 2468
rect 1866 2434 1900 2468
rect 1934 2434 1968 2468
rect 2002 2434 2036 2468
rect 2070 2434 2104 2468
rect 2138 2434 2172 2468
rect 2206 2434 2240 2468
rect 2274 2434 2352 2468
rect 1752 2423 2352 2434
rect 2748 2468 3748 2476
rect 2748 2434 2818 2468
rect 2852 2434 2886 2468
rect 2920 2434 2954 2468
rect 2988 2434 3022 2468
rect 3056 2434 3090 2468
rect 3124 2434 3158 2468
rect 3192 2434 3226 2468
rect 3260 2434 3294 2468
rect 3328 2434 3362 2468
rect 3396 2434 3430 2468
rect 3464 2434 3498 2468
rect 3532 2434 3566 2468
rect 3600 2434 3634 2468
rect 3668 2434 3702 2468
rect 3736 2434 3748 2468
rect 2748 2423 3748 2434
rect 1752 2312 2352 2323
rect 1752 2278 1764 2312
rect 1798 2278 1832 2312
rect 1866 2278 1900 2312
rect 1934 2278 1968 2312
rect 2002 2278 2036 2312
rect 2070 2278 2104 2312
rect 2138 2278 2172 2312
rect 2206 2278 2240 2312
rect 2274 2278 2352 2312
rect 1752 2267 2352 2278
rect 1175 2217 1475 2225
rect 1175 2183 1187 2217
rect 1221 2183 1255 2217
rect 1289 2183 1323 2217
rect 1357 2183 1391 2217
rect 1425 2183 1475 2217
rect 1175 2172 1475 2183
rect 2748 2312 3748 2323
rect 2748 2278 2818 2312
rect 2852 2278 2886 2312
rect 2920 2278 2954 2312
rect 2988 2278 3022 2312
rect 3056 2278 3090 2312
rect 3124 2278 3158 2312
rect 3192 2278 3226 2312
rect 3260 2278 3294 2312
rect 3328 2278 3362 2312
rect 3396 2278 3430 2312
rect 3464 2278 3498 2312
rect 3532 2278 3566 2312
rect 3600 2278 3634 2312
rect 3668 2278 3702 2312
rect 3736 2278 3748 2312
rect 2748 2267 3748 2278
rect 1752 2156 2352 2167
rect 1752 2122 1764 2156
rect 1798 2122 1832 2156
rect 1866 2122 1900 2156
rect 1934 2122 1968 2156
rect 2002 2122 2036 2156
rect 2070 2122 2104 2156
rect 2138 2122 2172 2156
rect 2206 2122 2240 2156
rect 2274 2122 2352 2156
rect 1752 2111 2352 2122
rect 1175 2061 1475 2072
rect 1175 2027 1187 2061
rect 1221 2027 1255 2061
rect 1289 2027 1323 2061
rect 1357 2027 1391 2061
rect 1425 2027 1475 2061
rect 1175 2019 1475 2027
rect 2748 2156 3748 2167
rect 2748 2122 2818 2156
rect 2852 2122 2886 2156
rect 2920 2122 2954 2156
rect 2988 2122 3022 2156
rect 3056 2122 3090 2156
rect 3124 2122 3158 2156
rect 3192 2122 3226 2156
rect 3260 2122 3294 2156
rect 3328 2122 3362 2156
rect 3396 2122 3430 2156
rect 3464 2122 3498 2156
rect 3532 2122 3566 2156
rect 3600 2122 3634 2156
rect 3668 2122 3702 2156
rect 3736 2122 3748 2156
rect 2748 2111 3748 2122
rect 1752 2000 2352 2011
rect 1752 1966 1764 2000
rect 1798 1966 1832 2000
rect 1866 1966 1900 2000
rect 1934 1966 1968 2000
rect 2002 1966 2036 2000
rect 2070 1966 2104 2000
rect 2138 1966 2172 2000
rect 2206 1966 2240 2000
rect 2274 1966 2352 2000
rect 1752 1955 2352 1966
rect 2748 2000 3748 2011
rect 2748 1966 2818 2000
rect 2852 1966 2886 2000
rect 2920 1966 2954 2000
rect 2988 1966 3022 2000
rect 3056 1966 3090 2000
rect 3124 1966 3158 2000
rect 3192 1966 3226 2000
rect 3260 1966 3294 2000
rect 3328 1966 3362 2000
rect 3396 1966 3430 2000
rect 3464 1966 3498 2000
rect 3532 1966 3566 2000
rect 3600 1966 3634 2000
rect 3668 1966 3702 2000
rect 3736 1966 3748 2000
rect 2748 1958 3748 1966
rect 1752 1844 2352 1855
rect 1752 1810 1764 1844
rect 1798 1810 1832 1844
rect 1866 1810 1900 1844
rect 1934 1810 1968 1844
rect 2002 1810 2036 1844
rect 2070 1810 2104 1844
rect 2138 1810 2172 1844
rect 2206 1810 2240 1844
rect 2274 1810 2352 1844
rect 1752 1802 2352 1810
rect 572 1131 625 1201
rect 572 1097 580 1131
rect 614 1097 625 1131
rect 572 1063 625 1097
rect 572 1029 580 1063
rect 614 1029 625 1063
rect 572 995 625 1029
rect 572 961 580 995
rect 614 961 625 995
rect 572 927 625 961
rect 572 893 580 927
rect 614 893 625 927
rect 572 859 625 893
rect 572 825 580 859
rect 614 825 625 859
rect 572 791 625 825
rect 572 757 580 791
rect 614 757 625 791
rect 572 723 625 757
rect 572 689 580 723
rect 614 689 625 723
rect 572 655 625 689
rect 572 621 580 655
rect 614 621 625 655
rect 572 587 625 621
rect 572 553 580 587
rect 614 553 625 587
rect 572 519 625 553
rect 572 485 580 519
rect 614 485 625 519
rect 572 451 625 485
rect 572 417 580 451
rect 614 417 625 451
rect 572 383 625 417
rect 572 349 580 383
rect 614 349 625 383
rect 572 315 625 349
rect 572 281 580 315
rect 614 281 625 315
rect 572 247 625 281
rect 572 213 580 247
rect 614 213 625 247
rect 572 201 625 213
rect 725 1131 781 1201
rect 725 1097 736 1131
rect 770 1097 781 1131
rect 725 1063 781 1097
rect 725 1029 736 1063
rect 770 1029 781 1063
rect 725 995 781 1029
rect 725 961 736 995
rect 770 961 781 995
rect 725 927 781 961
rect 725 893 736 927
rect 770 893 781 927
rect 725 859 781 893
rect 725 825 736 859
rect 770 825 781 859
rect 725 791 781 825
rect 725 757 736 791
rect 770 757 781 791
rect 725 723 781 757
rect 725 689 736 723
rect 770 689 781 723
rect 725 655 781 689
rect 725 621 736 655
rect 770 621 781 655
rect 725 587 781 621
rect 725 553 736 587
rect 770 553 781 587
rect 725 519 781 553
rect 725 485 736 519
rect 770 485 781 519
rect 725 451 781 485
rect 725 417 736 451
rect 770 417 781 451
rect 725 383 781 417
rect 725 349 736 383
rect 770 349 781 383
rect 725 315 781 349
rect 725 281 736 315
rect 770 281 781 315
rect 725 247 781 281
rect 725 213 736 247
rect 770 213 781 247
rect 725 201 781 213
rect 881 1131 937 1201
rect 881 1097 892 1131
rect 926 1097 937 1131
rect 881 1063 937 1097
rect 881 1029 892 1063
rect 926 1029 937 1063
rect 881 995 937 1029
rect 881 961 892 995
rect 926 961 937 995
rect 881 927 937 961
rect 881 893 892 927
rect 926 893 937 927
rect 881 859 937 893
rect 881 825 892 859
rect 926 825 937 859
rect 881 791 937 825
rect 881 757 892 791
rect 926 757 937 791
rect 881 723 937 757
rect 881 689 892 723
rect 926 689 937 723
rect 881 655 937 689
rect 881 621 892 655
rect 926 621 937 655
rect 881 587 937 621
rect 881 553 892 587
rect 926 553 937 587
rect 881 519 937 553
rect 881 485 892 519
rect 926 485 937 519
rect 881 451 937 485
rect 881 417 892 451
rect 926 417 937 451
rect 881 383 937 417
rect 881 349 892 383
rect 926 349 937 383
rect 881 315 937 349
rect 881 281 892 315
rect 926 281 937 315
rect 881 247 937 281
rect 881 213 892 247
rect 926 213 937 247
rect 881 201 937 213
rect 1037 1131 1093 1201
rect 1037 1097 1048 1131
rect 1082 1097 1093 1131
rect 1037 1063 1093 1097
rect 1037 1029 1048 1063
rect 1082 1029 1093 1063
rect 1037 995 1093 1029
rect 1037 961 1048 995
rect 1082 961 1093 995
rect 1037 927 1093 961
rect 1037 893 1048 927
rect 1082 893 1093 927
rect 1037 859 1093 893
rect 1037 825 1048 859
rect 1082 825 1093 859
rect 1037 791 1093 825
rect 1037 757 1048 791
rect 1082 757 1093 791
rect 1037 723 1093 757
rect 1037 689 1048 723
rect 1082 689 1093 723
rect 1037 655 1093 689
rect 1037 621 1048 655
rect 1082 621 1093 655
rect 1037 587 1093 621
rect 1037 553 1048 587
rect 1082 553 1093 587
rect 1037 519 1093 553
rect 1037 485 1048 519
rect 1082 485 1093 519
rect 1037 451 1093 485
rect 1037 417 1048 451
rect 1082 417 1093 451
rect 1037 383 1093 417
rect 1037 349 1048 383
rect 1082 349 1093 383
rect 1037 315 1093 349
rect 1037 281 1048 315
rect 1082 281 1093 315
rect 1037 247 1093 281
rect 1037 213 1048 247
rect 1082 213 1093 247
rect 1037 201 1093 213
rect 1193 1131 1249 1201
rect 1193 1097 1204 1131
rect 1238 1097 1249 1131
rect 1193 1063 1249 1097
rect 1193 1029 1204 1063
rect 1238 1029 1249 1063
rect 1193 995 1249 1029
rect 1193 961 1204 995
rect 1238 961 1249 995
rect 1193 927 1249 961
rect 1193 893 1204 927
rect 1238 893 1249 927
rect 1193 859 1249 893
rect 1193 825 1204 859
rect 1238 825 1249 859
rect 1193 791 1249 825
rect 1193 757 1204 791
rect 1238 757 1249 791
rect 1193 723 1249 757
rect 1193 689 1204 723
rect 1238 689 1249 723
rect 1193 655 1249 689
rect 1193 621 1204 655
rect 1238 621 1249 655
rect 1193 587 1249 621
rect 1193 553 1204 587
rect 1238 553 1249 587
rect 1193 519 1249 553
rect 1193 485 1204 519
rect 1238 485 1249 519
rect 1193 451 1249 485
rect 1193 417 1204 451
rect 1238 417 1249 451
rect 1193 383 1249 417
rect 1193 349 1204 383
rect 1238 349 1249 383
rect 1193 315 1249 349
rect 1193 281 1204 315
rect 1238 281 1249 315
rect 1193 247 1249 281
rect 1193 213 1204 247
rect 1238 213 1249 247
rect 1193 201 1249 213
rect 1349 1131 1405 1201
rect 1349 1097 1360 1131
rect 1394 1097 1405 1131
rect 1349 1063 1405 1097
rect 1349 1029 1360 1063
rect 1394 1029 1405 1063
rect 1349 995 1405 1029
rect 1349 961 1360 995
rect 1394 961 1405 995
rect 1349 927 1405 961
rect 1349 893 1360 927
rect 1394 893 1405 927
rect 1349 859 1405 893
rect 1349 825 1360 859
rect 1394 825 1405 859
rect 1349 791 1405 825
rect 1349 757 1360 791
rect 1394 757 1405 791
rect 1349 723 1405 757
rect 1349 689 1360 723
rect 1394 689 1405 723
rect 1349 655 1405 689
rect 1349 621 1360 655
rect 1394 621 1405 655
rect 1349 587 1405 621
rect 1349 553 1360 587
rect 1394 553 1405 587
rect 1349 519 1405 553
rect 1349 485 1360 519
rect 1394 485 1405 519
rect 1349 451 1405 485
rect 1349 417 1360 451
rect 1394 417 1405 451
rect 1349 383 1405 417
rect 1349 349 1360 383
rect 1394 349 1405 383
rect 1349 315 1405 349
rect 1349 281 1360 315
rect 1394 281 1405 315
rect 1349 247 1405 281
rect 1349 213 1360 247
rect 1394 213 1405 247
rect 1349 201 1405 213
rect 1505 1131 1561 1201
rect 1505 1097 1516 1131
rect 1550 1097 1561 1131
rect 1505 1063 1561 1097
rect 1505 1029 1516 1063
rect 1550 1029 1561 1063
rect 1505 995 1561 1029
rect 1505 961 1516 995
rect 1550 961 1561 995
rect 1505 927 1561 961
rect 1505 893 1516 927
rect 1550 893 1561 927
rect 1505 859 1561 893
rect 1505 825 1516 859
rect 1550 825 1561 859
rect 1505 791 1561 825
rect 1505 757 1516 791
rect 1550 757 1561 791
rect 1505 723 1561 757
rect 1505 689 1516 723
rect 1550 689 1561 723
rect 1505 655 1561 689
rect 1505 621 1516 655
rect 1550 621 1561 655
rect 1505 587 1561 621
rect 1505 553 1516 587
rect 1550 553 1561 587
rect 1505 519 1561 553
rect 1505 485 1516 519
rect 1550 485 1561 519
rect 1505 451 1561 485
rect 1505 417 1516 451
rect 1550 417 1561 451
rect 1505 383 1561 417
rect 1505 349 1516 383
rect 1550 349 1561 383
rect 1505 315 1561 349
rect 1505 281 1516 315
rect 1550 281 1561 315
rect 1505 247 1561 281
rect 1505 213 1516 247
rect 1550 213 1561 247
rect 1505 201 1561 213
rect 1661 1131 1717 1201
rect 1661 1097 1672 1131
rect 1706 1097 1717 1131
rect 1661 1063 1717 1097
rect 1661 1029 1672 1063
rect 1706 1029 1717 1063
rect 1661 995 1717 1029
rect 1661 961 1672 995
rect 1706 961 1717 995
rect 1661 927 1717 961
rect 1661 893 1672 927
rect 1706 893 1717 927
rect 1661 859 1717 893
rect 1661 825 1672 859
rect 1706 825 1717 859
rect 1661 791 1717 825
rect 1661 757 1672 791
rect 1706 757 1717 791
rect 1661 723 1717 757
rect 1661 689 1672 723
rect 1706 689 1717 723
rect 1661 655 1717 689
rect 1661 621 1672 655
rect 1706 621 1717 655
rect 1661 587 1717 621
rect 1661 553 1672 587
rect 1706 553 1717 587
rect 1661 519 1717 553
rect 1661 485 1672 519
rect 1706 485 1717 519
rect 1661 451 1717 485
rect 1661 417 1672 451
rect 1706 417 1717 451
rect 1661 383 1717 417
rect 1661 349 1672 383
rect 1706 349 1717 383
rect 1661 315 1717 349
rect 1661 281 1672 315
rect 1706 281 1717 315
rect 1661 247 1717 281
rect 1661 213 1672 247
rect 1706 213 1717 247
rect 1661 201 1717 213
rect 1817 1131 1870 1201
rect 1817 1097 1828 1131
rect 1862 1097 1870 1131
rect 1817 1063 1870 1097
rect 1817 1029 1828 1063
rect 1862 1029 1870 1063
rect 1817 995 1870 1029
rect 1817 961 1828 995
rect 1862 961 1870 995
rect 1817 927 1870 961
rect 1817 893 1828 927
rect 1862 893 1870 927
rect 1817 859 1870 893
rect 1817 825 1828 859
rect 1862 825 1870 859
rect 1817 791 1870 825
rect 1817 757 1828 791
rect 1862 757 1870 791
rect 1817 723 1870 757
rect 1817 689 1828 723
rect 1862 689 1870 723
rect 1817 655 1870 689
rect 1817 621 1828 655
rect 1862 621 1870 655
rect 1817 587 1870 621
rect 1817 553 1828 587
rect 1862 553 1870 587
rect 1817 519 1870 553
rect 1817 485 1828 519
rect 1862 485 1870 519
rect 1817 451 1870 485
rect 1817 417 1828 451
rect 1862 417 1870 451
rect 1817 383 1870 417
rect 1817 349 1828 383
rect 1862 349 1870 383
rect 1817 315 1870 349
rect 1817 281 1828 315
rect 1862 281 1870 315
rect 1817 247 1870 281
rect 1817 213 1828 247
rect 1862 213 1870 247
rect 1817 201 1870 213
rect 1930 1131 1983 1201
rect 1930 1097 1938 1131
rect 1972 1097 1983 1131
rect 1930 1063 1983 1097
rect 1930 1029 1938 1063
rect 1972 1029 1983 1063
rect 1930 995 1983 1029
rect 1930 961 1938 995
rect 1972 961 1983 995
rect 1930 927 1983 961
rect 1930 893 1938 927
rect 1972 893 1983 927
rect 1930 859 1983 893
rect 1930 825 1938 859
rect 1972 825 1983 859
rect 1930 791 1983 825
rect 1930 757 1938 791
rect 1972 757 1983 791
rect 1930 723 1983 757
rect 1930 689 1938 723
rect 1972 689 1983 723
rect 1930 655 1983 689
rect 1930 621 1938 655
rect 1972 621 1983 655
rect 1930 587 1983 621
rect 1930 553 1938 587
rect 1972 553 1983 587
rect 1930 519 1983 553
rect 1930 485 1938 519
rect 1972 485 1983 519
rect 1930 451 1983 485
rect 1930 417 1938 451
rect 1972 417 1983 451
rect 1930 383 1983 417
rect 1930 349 1938 383
rect 1972 349 1983 383
rect 1930 315 1983 349
rect 1930 281 1938 315
rect 1972 281 1983 315
rect 1930 247 1983 281
rect 1930 213 1938 247
rect 1972 213 1983 247
rect 1930 201 1983 213
rect 2083 1131 2139 1201
rect 2083 1097 2094 1131
rect 2128 1097 2139 1131
rect 2083 1063 2139 1097
rect 2083 1029 2094 1063
rect 2128 1029 2139 1063
rect 2083 995 2139 1029
rect 2083 961 2094 995
rect 2128 961 2139 995
rect 2083 927 2139 961
rect 2083 893 2094 927
rect 2128 893 2139 927
rect 2083 859 2139 893
rect 2083 825 2094 859
rect 2128 825 2139 859
rect 2083 791 2139 825
rect 2083 757 2094 791
rect 2128 757 2139 791
rect 2083 723 2139 757
rect 2083 689 2094 723
rect 2128 689 2139 723
rect 2083 655 2139 689
rect 2083 621 2094 655
rect 2128 621 2139 655
rect 2083 587 2139 621
rect 2083 553 2094 587
rect 2128 553 2139 587
rect 2083 519 2139 553
rect 2083 485 2094 519
rect 2128 485 2139 519
rect 2083 451 2139 485
rect 2083 417 2094 451
rect 2128 417 2139 451
rect 2083 383 2139 417
rect 2083 349 2094 383
rect 2128 349 2139 383
rect 2083 315 2139 349
rect 2083 281 2094 315
rect 2128 281 2139 315
rect 2083 247 2139 281
rect 2083 213 2094 247
rect 2128 213 2139 247
rect 2083 201 2139 213
rect 2239 1131 2295 1201
rect 2239 1097 2250 1131
rect 2284 1097 2295 1131
rect 2239 1063 2295 1097
rect 2239 1029 2250 1063
rect 2284 1029 2295 1063
rect 2239 995 2295 1029
rect 2239 961 2250 995
rect 2284 961 2295 995
rect 2239 927 2295 961
rect 2239 893 2250 927
rect 2284 893 2295 927
rect 2239 859 2295 893
rect 2239 825 2250 859
rect 2284 825 2295 859
rect 2239 791 2295 825
rect 2239 757 2250 791
rect 2284 757 2295 791
rect 2239 723 2295 757
rect 2239 689 2250 723
rect 2284 689 2295 723
rect 2239 655 2295 689
rect 2239 621 2250 655
rect 2284 621 2295 655
rect 2239 587 2295 621
rect 2239 553 2250 587
rect 2284 553 2295 587
rect 2239 519 2295 553
rect 2239 485 2250 519
rect 2284 485 2295 519
rect 2239 451 2295 485
rect 2239 417 2250 451
rect 2284 417 2295 451
rect 2239 383 2295 417
rect 2239 349 2250 383
rect 2284 349 2295 383
rect 2239 315 2295 349
rect 2239 281 2250 315
rect 2284 281 2295 315
rect 2239 247 2295 281
rect 2239 213 2250 247
rect 2284 213 2295 247
rect 2239 201 2295 213
rect 2395 1131 2451 1201
rect 2395 1097 2406 1131
rect 2440 1097 2451 1131
rect 2395 1063 2451 1097
rect 2395 1029 2406 1063
rect 2440 1029 2451 1063
rect 2395 995 2451 1029
rect 2395 961 2406 995
rect 2440 961 2451 995
rect 2395 927 2451 961
rect 2395 893 2406 927
rect 2440 893 2451 927
rect 2395 859 2451 893
rect 2395 825 2406 859
rect 2440 825 2451 859
rect 2395 791 2451 825
rect 2395 757 2406 791
rect 2440 757 2451 791
rect 2395 723 2451 757
rect 2395 689 2406 723
rect 2440 689 2451 723
rect 2395 655 2451 689
rect 2395 621 2406 655
rect 2440 621 2451 655
rect 2395 587 2451 621
rect 2395 553 2406 587
rect 2440 553 2451 587
rect 2395 519 2451 553
rect 2395 485 2406 519
rect 2440 485 2451 519
rect 2395 451 2451 485
rect 2395 417 2406 451
rect 2440 417 2451 451
rect 2395 383 2451 417
rect 2395 349 2406 383
rect 2440 349 2451 383
rect 2395 315 2451 349
rect 2395 281 2406 315
rect 2440 281 2451 315
rect 2395 247 2451 281
rect 2395 213 2406 247
rect 2440 213 2451 247
rect 2395 201 2451 213
rect 2551 1131 2607 1201
rect 2551 1097 2562 1131
rect 2596 1097 2607 1131
rect 2551 1063 2607 1097
rect 2551 1029 2562 1063
rect 2596 1029 2607 1063
rect 2551 995 2607 1029
rect 2551 961 2562 995
rect 2596 961 2607 995
rect 2551 927 2607 961
rect 2551 893 2562 927
rect 2596 893 2607 927
rect 2551 859 2607 893
rect 2551 825 2562 859
rect 2596 825 2607 859
rect 2551 791 2607 825
rect 2551 757 2562 791
rect 2596 757 2607 791
rect 2551 723 2607 757
rect 2551 689 2562 723
rect 2596 689 2607 723
rect 2551 655 2607 689
rect 2551 621 2562 655
rect 2596 621 2607 655
rect 2551 587 2607 621
rect 2551 553 2562 587
rect 2596 553 2607 587
rect 2551 519 2607 553
rect 2551 485 2562 519
rect 2596 485 2607 519
rect 2551 451 2607 485
rect 2551 417 2562 451
rect 2596 417 2607 451
rect 2551 383 2607 417
rect 2551 349 2562 383
rect 2596 349 2607 383
rect 2551 315 2607 349
rect 2551 281 2562 315
rect 2596 281 2607 315
rect 2551 247 2607 281
rect 2551 213 2562 247
rect 2596 213 2607 247
rect 2551 201 2607 213
rect 2707 1131 2763 1201
rect 2707 1097 2718 1131
rect 2752 1097 2763 1131
rect 2707 1063 2763 1097
rect 2707 1029 2718 1063
rect 2752 1029 2763 1063
rect 2707 995 2763 1029
rect 2707 961 2718 995
rect 2752 961 2763 995
rect 2707 927 2763 961
rect 2707 893 2718 927
rect 2752 893 2763 927
rect 2707 859 2763 893
rect 2707 825 2718 859
rect 2752 825 2763 859
rect 2707 791 2763 825
rect 2707 757 2718 791
rect 2752 757 2763 791
rect 2707 723 2763 757
rect 2707 689 2718 723
rect 2752 689 2763 723
rect 2707 655 2763 689
rect 2707 621 2718 655
rect 2752 621 2763 655
rect 2707 587 2763 621
rect 2707 553 2718 587
rect 2752 553 2763 587
rect 2707 519 2763 553
rect 2707 485 2718 519
rect 2752 485 2763 519
rect 2707 451 2763 485
rect 2707 417 2718 451
rect 2752 417 2763 451
rect 2707 383 2763 417
rect 2707 349 2718 383
rect 2752 349 2763 383
rect 2707 315 2763 349
rect 2707 281 2718 315
rect 2752 281 2763 315
rect 2707 247 2763 281
rect 2707 213 2718 247
rect 2752 213 2763 247
rect 2707 201 2763 213
rect 2863 1131 2919 1201
rect 2863 1097 2874 1131
rect 2908 1097 2919 1131
rect 2863 1063 2919 1097
rect 2863 1029 2874 1063
rect 2908 1029 2919 1063
rect 2863 995 2919 1029
rect 2863 961 2874 995
rect 2908 961 2919 995
rect 2863 927 2919 961
rect 2863 893 2874 927
rect 2908 893 2919 927
rect 2863 859 2919 893
rect 2863 825 2874 859
rect 2908 825 2919 859
rect 2863 791 2919 825
rect 2863 757 2874 791
rect 2908 757 2919 791
rect 2863 723 2919 757
rect 2863 689 2874 723
rect 2908 689 2919 723
rect 2863 655 2919 689
rect 2863 621 2874 655
rect 2908 621 2919 655
rect 2863 587 2919 621
rect 2863 553 2874 587
rect 2908 553 2919 587
rect 2863 519 2919 553
rect 2863 485 2874 519
rect 2908 485 2919 519
rect 2863 451 2919 485
rect 2863 417 2874 451
rect 2908 417 2919 451
rect 2863 383 2919 417
rect 2863 349 2874 383
rect 2908 349 2919 383
rect 2863 315 2919 349
rect 2863 281 2874 315
rect 2908 281 2919 315
rect 2863 247 2919 281
rect 2863 213 2874 247
rect 2908 213 2919 247
rect 2863 201 2919 213
rect 3019 1131 3072 1201
rect 3019 1097 3030 1131
rect 3064 1097 3072 1131
rect 3019 1063 3072 1097
rect 3019 1029 3030 1063
rect 3064 1029 3072 1063
rect 3019 995 3072 1029
rect 3019 961 3030 995
rect 3064 961 3072 995
rect 3019 927 3072 961
rect 3019 893 3030 927
rect 3064 893 3072 927
rect 3019 859 3072 893
rect 3019 825 3030 859
rect 3064 825 3072 859
rect 3019 791 3072 825
rect 3019 757 3030 791
rect 3064 757 3072 791
rect 3019 723 3072 757
rect 3019 689 3030 723
rect 3064 689 3072 723
rect 3019 655 3072 689
rect 3019 621 3030 655
rect 3064 621 3072 655
rect 3019 587 3072 621
rect 3019 553 3030 587
rect 3064 553 3072 587
rect 3019 519 3072 553
rect 3019 485 3030 519
rect 3064 485 3072 519
rect 3019 451 3072 485
rect 3019 417 3030 451
rect 3064 417 3072 451
rect 3019 383 3072 417
rect 3019 349 3030 383
rect 3064 349 3072 383
rect 3019 315 3072 349
rect 3019 281 3030 315
rect 3064 281 3072 315
rect 3019 247 3072 281
rect 3019 213 3030 247
rect 3064 213 3072 247
rect 3019 201 3072 213
<< mvpdiff >>
rect 1290 3864 1343 3876
rect 1290 3830 1298 3864
rect 1332 3830 1343 3864
rect 1290 3796 1343 3830
rect 1290 3762 1298 3796
rect 1332 3762 1343 3796
rect 1290 3728 1343 3762
rect 1290 3694 1298 3728
rect 1332 3694 1343 3728
rect 1290 3660 1343 3694
rect 1290 3626 1298 3660
rect 1332 3626 1343 3660
rect 1290 3592 1343 3626
rect 1290 3558 1298 3592
rect 1332 3558 1343 3592
rect 1290 3524 1343 3558
rect 1290 3490 1298 3524
rect 1332 3490 1343 3524
rect 1290 3456 1343 3490
rect 1290 3422 1298 3456
rect 1332 3422 1343 3456
rect 1290 3388 1343 3422
rect 1290 3354 1298 3388
rect 1332 3354 1343 3388
rect 1290 3320 1343 3354
rect 1290 3286 1298 3320
rect 1332 3286 1343 3320
rect 1290 3252 1343 3286
rect 1290 3218 1298 3252
rect 1332 3218 1343 3252
rect 1290 3184 1343 3218
rect 602 3164 655 3176
rect 602 3130 610 3164
rect 644 3130 655 3164
rect 602 3096 655 3130
rect 602 3062 610 3096
rect 644 3062 655 3096
rect 602 3028 655 3062
rect 602 2994 610 3028
rect 644 2994 655 3028
rect 602 2960 655 2994
rect 602 2926 610 2960
rect 644 2926 655 2960
rect 602 2876 655 2926
rect 755 3164 811 3176
rect 755 3130 766 3164
rect 800 3130 811 3164
rect 755 3096 811 3130
rect 755 3062 766 3096
rect 800 3062 811 3096
rect 755 3028 811 3062
rect 755 2994 766 3028
rect 800 2994 811 3028
rect 755 2960 811 2994
rect 755 2926 766 2960
rect 800 2926 811 2960
rect 755 2876 811 2926
rect 911 3164 964 3176
rect 911 3130 922 3164
rect 956 3130 964 3164
rect 911 3096 964 3130
rect 911 3062 922 3096
rect 956 3062 964 3096
rect 911 3028 964 3062
rect 911 2994 922 3028
rect 956 2994 964 3028
rect 911 2960 964 2994
rect 911 2926 922 2960
rect 956 2926 964 2960
rect 911 2876 964 2926
rect 1024 3164 1077 3176
rect 1024 3130 1032 3164
rect 1066 3130 1077 3164
rect 1024 3096 1077 3130
rect 1024 3062 1032 3096
rect 1066 3062 1077 3096
rect 1024 3028 1077 3062
rect 1024 2994 1032 3028
rect 1066 2994 1077 3028
rect 1024 2960 1077 2994
rect 1024 2926 1032 2960
rect 1066 2926 1077 2960
rect 1024 2876 1077 2926
rect 1177 3164 1230 3176
rect 1177 3130 1188 3164
rect 1222 3130 1230 3164
rect 1177 3096 1230 3130
rect 1177 3062 1188 3096
rect 1222 3062 1230 3096
rect 1177 3028 1230 3062
rect 1177 2994 1188 3028
rect 1222 2994 1230 3028
rect 1177 2960 1230 2994
rect 1177 2926 1188 2960
rect 1222 2926 1230 2960
rect 1177 2876 1230 2926
rect 1290 3150 1298 3184
rect 1332 3150 1343 3184
rect 1290 3116 1343 3150
rect 1290 3082 1298 3116
rect 1332 3082 1343 3116
rect 1290 3048 1343 3082
rect 1290 3014 1298 3048
rect 1332 3014 1343 3048
rect 1290 2980 1343 3014
rect 1290 2946 1298 2980
rect 1332 2946 1343 2980
rect 1290 2876 1343 2946
rect 1443 3864 1499 3876
rect 1443 3830 1454 3864
rect 1488 3830 1499 3864
rect 1443 3796 1499 3830
rect 1443 3762 1454 3796
rect 1488 3762 1499 3796
rect 1443 3728 1499 3762
rect 1443 3694 1454 3728
rect 1488 3694 1499 3728
rect 1443 3660 1499 3694
rect 1443 3626 1454 3660
rect 1488 3626 1499 3660
rect 1443 3592 1499 3626
rect 1443 3558 1454 3592
rect 1488 3558 1499 3592
rect 1443 3524 1499 3558
rect 1443 3490 1454 3524
rect 1488 3490 1499 3524
rect 1443 3456 1499 3490
rect 1443 3422 1454 3456
rect 1488 3422 1499 3456
rect 1443 3388 1499 3422
rect 1443 3354 1454 3388
rect 1488 3354 1499 3388
rect 1443 3320 1499 3354
rect 1443 3286 1454 3320
rect 1488 3286 1499 3320
rect 1443 3252 1499 3286
rect 1443 3218 1454 3252
rect 1488 3218 1499 3252
rect 1443 3184 1499 3218
rect 1443 3150 1454 3184
rect 1488 3150 1499 3184
rect 1443 3116 1499 3150
rect 1443 3082 1454 3116
rect 1488 3082 1499 3116
rect 1443 3048 1499 3082
rect 1443 3014 1454 3048
rect 1488 3014 1499 3048
rect 1443 2980 1499 3014
rect 1443 2946 1454 2980
rect 1488 2946 1499 2980
rect 1443 2876 1499 2946
rect 1599 3864 1655 3876
rect 1599 3830 1610 3864
rect 1644 3830 1655 3864
rect 1599 3796 1655 3830
rect 1599 3762 1610 3796
rect 1644 3762 1655 3796
rect 1599 3728 1655 3762
rect 1599 3694 1610 3728
rect 1644 3694 1655 3728
rect 1599 3660 1655 3694
rect 1599 3626 1610 3660
rect 1644 3626 1655 3660
rect 1599 3592 1655 3626
rect 1599 3558 1610 3592
rect 1644 3558 1655 3592
rect 1599 3524 1655 3558
rect 1599 3490 1610 3524
rect 1644 3490 1655 3524
rect 1599 3456 1655 3490
rect 1599 3422 1610 3456
rect 1644 3422 1655 3456
rect 1599 3388 1655 3422
rect 1599 3354 1610 3388
rect 1644 3354 1655 3388
rect 1599 3320 1655 3354
rect 1599 3286 1610 3320
rect 1644 3286 1655 3320
rect 1599 3252 1655 3286
rect 1599 3218 1610 3252
rect 1644 3218 1655 3252
rect 1599 3184 1655 3218
rect 1599 3150 1610 3184
rect 1644 3150 1655 3184
rect 1599 3116 1655 3150
rect 1599 3082 1610 3116
rect 1644 3082 1655 3116
rect 1599 3048 1655 3082
rect 1599 3014 1610 3048
rect 1644 3014 1655 3048
rect 1599 2980 1655 3014
rect 1599 2946 1610 2980
rect 1644 2946 1655 2980
rect 1599 2876 1655 2946
rect 1755 3864 1811 3876
rect 1755 3830 1766 3864
rect 1800 3830 1811 3864
rect 1755 3796 1811 3830
rect 1755 3762 1766 3796
rect 1800 3762 1811 3796
rect 1755 3728 1811 3762
rect 1755 3694 1766 3728
rect 1800 3694 1811 3728
rect 1755 3660 1811 3694
rect 1755 3626 1766 3660
rect 1800 3626 1811 3660
rect 1755 3592 1811 3626
rect 1755 3558 1766 3592
rect 1800 3558 1811 3592
rect 1755 3524 1811 3558
rect 1755 3490 1766 3524
rect 1800 3490 1811 3524
rect 1755 3456 1811 3490
rect 1755 3422 1766 3456
rect 1800 3422 1811 3456
rect 1755 3388 1811 3422
rect 1755 3354 1766 3388
rect 1800 3354 1811 3388
rect 1755 3320 1811 3354
rect 1755 3286 1766 3320
rect 1800 3286 1811 3320
rect 1755 3252 1811 3286
rect 1755 3218 1766 3252
rect 1800 3218 1811 3252
rect 1755 3184 1811 3218
rect 1755 3150 1766 3184
rect 1800 3150 1811 3184
rect 1755 3116 1811 3150
rect 1755 3082 1766 3116
rect 1800 3082 1811 3116
rect 1755 3048 1811 3082
rect 1755 3014 1766 3048
rect 1800 3014 1811 3048
rect 1755 2980 1811 3014
rect 1755 2946 1766 2980
rect 1800 2946 1811 2980
rect 1755 2876 1811 2946
rect 1911 3864 1964 3876
rect 1911 3830 1922 3864
rect 1956 3830 1964 3864
rect 1911 3796 1964 3830
rect 1911 3762 1922 3796
rect 1956 3762 1964 3796
rect 1911 3728 1964 3762
rect 1911 3694 1922 3728
rect 1956 3694 1964 3728
rect 1911 3660 1964 3694
rect 1911 3626 1922 3660
rect 1956 3626 1964 3660
rect 1911 3592 1964 3626
rect 1911 3558 1922 3592
rect 1956 3558 1964 3592
rect 1911 3524 1964 3558
rect 1911 3490 1922 3524
rect 1956 3490 1964 3524
rect 1911 3456 1964 3490
rect 1911 3422 1922 3456
rect 1956 3422 1964 3456
rect 1911 3388 1964 3422
rect 1911 3354 1922 3388
rect 1956 3354 1964 3388
rect 1911 3320 1964 3354
rect 1911 3286 1922 3320
rect 1956 3286 1964 3320
rect 1911 3252 1964 3286
rect 1911 3218 1922 3252
rect 1956 3218 1964 3252
rect 1911 3184 1964 3218
rect 1911 3150 1922 3184
rect 1956 3150 1964 3184
rect 1911 3116 1964 3150
rect 1911 3082 1922 3116
rect 1956 3082 1964 3116
rect 1911 3048 1964 3082
rect 1911 3014 1922 3048
rect 1956 3014 1964 3048
rect 1911 2980 1964 3014
rect 1911 2946 1922 2980
rect 1956 2946 1964 2980
rect 1911 2876 1964 2946
rect 2024 3864 2077 3876
rect 2024 3830 2032 3864
rect 2066 3830 2077 3864
rect 2024 3796 2077 3830
rect 2024 3762 2032 3796
rect 2066 3762 2077 3796
rect 2024 3728 2077 3762
rect 2024 3694 2032 3728
rect 2066 3694 2077 3728
rect 2024 3660 2077 3694
rect 2024 3626 2032 3660
rect 2066 3626 2077 3660
rect 2024 3592 2077 3626
rect 2024 3558 2032 3592
rect 2066 3558 2077 3592
rect 2024 3524 2077 3558
rect 2024 3490 2032 3524
rect 2066 3490 2077 3524
rect 2024 3456 2077 3490
rect 2024 3422 2032 3456
rect 2066 3422 2077 3456
rect 2024 3388 2077 3422
rect 2024 3354 2032 3388
rect 2066 3354 2077 3388
rect 2024 3320 2077 3354
rect 2024 3286 2032 3320
rect 2066 3286 2077 3320
rect 2024 3252 2077 3286
rect 2024 3218 2032 3252
rect 2066 3218 2077 3252
rect 2024 3184 2077 3218
rect 2024 3150 2032 3184
rect 2066 3150 2077 3184
rect 2024 3116 2077 3150
rect 2024 3082 2032 3116
rect 2066 3082 2077 3116
rect 2024 3048 2077 3082
rect 2024 3014 2032 3048
rect 2066 3014 2077 3048
rect 2024 2980 2077 3014
rect 2024 2946 2032 2980
rect 2066 2946 2077 2980
rect 2024 2876 2077 2946
rect 2177 3864 2233 3876
rect 2177 3830 2188 3864
rect 2222 3830 2233 3864
rect 2177 3796 2233 3830
rect 2177 3762 2188 3796
rect 2222 3762 2233 3796
rect 2177 3728 2233 3762
rect 2177 3694 2188 3728
rect 2222 3694 2233 3728
rect 2177 3660 2233 3694
rect 2177 3626 2188 3660
rect 2222 3626 2233 3660
rect 2177 3592 2233 3626
rect 2177 3558 2188 3592
rect 2222 3558 2233 3592
rect 2177 3524 2233 3558
rect 2177 3490 2188 3524
rect 2222 3490 2233 3524
rect 2177 3456 2233 3490
rect 2177 3422 2188 3456
rect 2222 3422 2233 3456
rect 2177 3388 2233 3422
rect 2177 3354 2188 3388
rect 2222 3354 2233 3388
rect 2177 3320 2233 3354
rect 2177 3286 2188 3320
rect 2222 3286 2233 3320
rect 2177 3252 2233 3286
rect 2177 3218 2188 3252
rect 2222 3218 2233 3252
rect 2177 3184 2233 3218
rect 2177 3150 2188 3184
rect 2222 3150 2233 3184
rect 2177 3116 2233 3150
rect 2177 3082 2188 3116
rect 2222 3082 2233 3116
rect 2177 3048 2233 3082
rect 2177 3014 2188 3048
rect 2222 3014 2233 3048
rect 2177 2980 2233 3014
rect 2177 2946 2188 2980
rect 2222 2946 2233 2980
rect 2177 2876 2233 2946
rect 2333 3864 2389 3876
rect 2333 3830 2344 3864
rect 2378 3830 2389 3864
rect 2333 3796 2389 3830
rect 2333 3762 2344 3796
rect 2378 3762 2389 3796
rect 2333 3728 2389 3762
rect 2333 3694 2344 3728
rect 2378 3694 2389 3728
rect 2333 3660 2389 3694
rect 2333 3626 2344 3660
rect 2378 3626 2389 3660
rect 2333 3592 2389 3626
rect 2333 3558 2344 3592
rect 2378 3558 2389 3592
rect 2333 3524 2389 3558
rect 2333 3490 2344 3524
rect 2378 3490 2389 3524
rect 2333 3456 2389 3490
rect 2333 3422 2344 3456
rect 2378 3422 2389 3456
rect 2333 3388 2389 3422
rect 2333 3354 2344 3388
rect 2378 3354 2389 3388
rect 2333 3320 2389 3354
rect 2333 3286 2344 3320
rect 2378 3286 2389 3320
rect 2333 3252 2389 3286
rect 2333 3218 2344 3252
rect 2378 3218 2389 3252
rect 2333 3184 2389 3218
rect 2333 3150 2344 3184
rect 2378 3150 2389 3184
rect 2333 3116 2389 3150
rect 2333 3082 2344 3116
rect 2378 3082 2389 3116
rect 2333 3048 2389 3082
rect 2333 3014 2344 3048
rect 2378 3014 2389 3048
rect 2333 2980 2389 3014
rect 2333 2946 2344 2980
rect 2378 2946 2389 2980
rect 2333 2876 2389 2946
rect 2489 3864 2545 3876
rect 2489 3830 2500 3864
rect 2534 3830 2545 3864
rect 2489 3796 2545 3830
rect 2489 3762 2500 3796
rect 2534 3762 2545 3796
rect 2489 3728 2545 3762
rect 2489 3694 2500 3728
rect 2534 3694 2545 3728
rect 2489 3660 2545 3694
rect 2489 3626 2500 3660
rect 2534 3626 2545 3660
rect 2489 3592 2545 3626
rect 2489 3558 2500 3592
rect 2534 3558 2545 3592
rect 2489 3524 2545 3558
rect 2489 3490 2500 3524
rect 2534 3490 2545 3524
rect 2489 3456 2545 3490
rect 2489 3422 2500 3456
rect 2534 3422 2545 3456
rect 2489 3388 2545 3422
rect 2489 3354 2500 3388
rect 2534 3354 2545 3388
rect 2489 3320 2545 3354
rect 2489 3286 2500 3320
rect 2534 3286 2545 3320
rect 2489 3252 2545 3286
rect 2489 3218 2500 3252
rect 2534 3218 2545 3252
rect 2489 3184 2545 3218
rect 2489 3150 2500 3184
rect 2534 3150 2545 3184
rect 2489 3116 2545 3150
rect 2489 3082 2500 3116
rect 2534 3082 2545 3116
rect 2489 3048 2545 3082
rect 2489 3014 2500 3048
rect 2534 3014 2545 3048
rect 2489 2980 2545 3014
rect 2489 2946 2500 2980
rect 2534 2946 2545 2980
rect 2489 2876 2545 2946
rect 2645 3864 2698 3876
rect 2645 3830 2656 3864
rect 2690 3830 2698 3864
rect 2645 3796 2698 3830
rect 2645 3762 2656 3796
rect 2690 3762 2698 3796
rect 2645 3728 2698 3762
rect 2645 3694 2656 3728
rect 2690 3694 2698 3728
rect 2645 3660 2698 3694
rect 2645 3626 2656 3660
rect 2690 3626 2698 3660
rect 2645 3592 2698 3626
rect 2645 3558 2656 3592
rect 2690 3558 2698 3592
rect 2645 3524 2698 3558
rect 2645 3490 2656 3524
rect 2690 3490 2698 3524
rect 2645 3456 2698 3490
rect 2645 3422 2656 3456
rect 2690 3422 2698 3456
rect 2645 3388 2698 3422
rect 2645 3354 2656 3388
rect 2690 3354 2698 3388
rect 2645 3320 2698 3354
rect 2645 3286 2656 3320
rect 2690 3286 2698 3320
rect 2645 3252 2698 3286
rect 2645 3218 2656 3252
rect 2690 3218 2698 3252
rect 2645 3184 2698 3218
rect 2645 3150 2656 3184
rect 2690 3150 2698 3184
rect 2645 3116 2698 3150
rect 2645 3082 2656 3116
rect 2690 3082 2698 3116
rect 2645 3048 2698 3082
rect 2645 3014 2656 3048
rect 2690 3014 2698 3048
rect 2645 2980 2698 3014
rect 2645 2946 2656 2980
rect 2690 2946 2698 2980
rect 2645 2876 2698 2946
rect 2758 3864 2811 3876
rect 2758 3830 2766 3864
rect 2800 3830 2811 3864
rect 2758 3796 2811 3830
rect 2758 3762 2766 3796
rect 2800 3762 2811 3796
rect 2758 3728 2811 3762
rect 2758 3694 2766 3728
rect 2800 3694 2811 3728
rect 2758 3660 2811 3694
rect 2758 3626 2766 3660
rect 2800 3626 2811 3660
rect 2758 3592 2811 3626
rect 2758 3558 2766 3592
rect 2800 3558 2811 3592
rect 2758 3524 2811 3558
rect 2758 3490 2766 3524
rect 2800 3490 2811 3524
rect 2758 3456 2811 3490
rect 2758 3422 2766 3456
rect 2800 3422 2811 3456
rect 2758 3388 2811 3422
rect 2758 3354 2766 3388
rect 2800 3354 2811 3388
rect 2758 3320 2811 3354
rect 2758 3286 2766 3320
rect 2800 3286 2811 3320
rect 2758 3252 2811 3286
rect 2758 3218 2766 3252
rect 2800 3218 2811 3252
rect 2758 3184 2811 3218
rect 2758 3150 2766 3184
rect 2800 3150 2811 3184
rect 2758 3116 2811 3150
rect 2758 3082 2766 3116
rect 2800 3082 2811 3116
rect 2758 3048 2811 3082
rect 2758 3014 2766 3048
rect 2800 3014 2811 3048
rect 2758 2980 2811 3014
rect 2758 2946 2766 2980
rect 2800 2946 2811 2980
rect 2758 2876 2811 2946
rect 2911 3864 2967 3876
rect 2911 3830 2922 3864
rect 2956 3830 2967 3864
rect 2911 3796 2967 3830
rect 2911 3762 2922 3796
rect 2956 3762 2967 3796
rect 2911 3728 2967 3762
rect 2911 3694 2922 3728
rect 2956 3694 2967 3728
rect 2911 3660 2967 3694
rect 2911 3626 2922 3660
rect 2956 3626 2967 3660
rect 2911 3592 2967 3626
rect 2911 3558 2922 3592
rect 2956 3558 2967 3592
rect 2911 3524 2967 3558
rect 2911 3490 2922 3524
rect 2956 3490 2967 3524
rect 2911 3456 2967 3490
rect 2911 3422 2922 3456
rect 2956 3422 2967 3456
rect 2911 3388 2967 3422
rect 2911 3354 2922 3388
rect 2956 3354 2967 3388
rect 2911 3320 2967 3354
rect 2911 3286 2922 3320
rect 2956 3286 2967 3320
rect 2911 3252 2967 3286
rect 2911 3218 2922 3252
rect 2956 3218 2967 3252
rect 2911 3184 2967 3218
rect 2911 3150 2922 3184
rect 2956 3150 2967 3184
rect 2911 3116 2967 3150
rect 2911 3082 2922 3116
rect 2956 3082 2967 3116
rect 2911 3048 2967 3082
rect 2911 3014 2922 3048
rect 2956 3014 2967 3048
rect 2911 2980 2967 3014
rect 2911 2946 2922 2980
rect 2956 2946 2967 2980
rect 2911 2876 2967 2946
rect 3067 3864 3120 3876
rect 3067 3830 3078 3864
rect 3112 3830 3120 3864
rect 3067 3796 3120 3830
rect 3067 3762 3078 3796
rect 3112 3762 3120 3796
rect 3067 3728 3120 3762
rect 3067 3694 3078 3728
rect 3112 3694 3120 3728
rect 3067 3660 3120 3694
rect 3067 3626 3078 3660
rect 3112 3626 3120 3660
rect 3067 3592 3120 3626
rect 3067 3558 3078 3592
rect 3112 3558 3120 3592
rect 3067 3524 3120 3558
rect 3067 3490 3078 3524
rect 3112 3490 3120 3524
rect 3067 3456 3120 3490
rect 3067 3422 3078 3456
rect 3112 3422 3120 3456
rect 3067 3388 3120 3422
rect 3067 3354 3078 3388
rect 3112 3354 3120 3388
rect 3067 3320 3120 3354
rect 3067 3286 3078 3320
rect 3112 3286 3120 3320
rect 3067 3252 3120 3286
rect 3067 3218 3078 3252
rect 3112 3218 3120 3252
rect 3067 3184 3120 3218
rect 3067 3150 3078 3184
rect 3112 3150 3120 3184
rect 3067 3116 3120 3150
rect 3067 3082 3078 3116
rect 3112 3082 3120 3116
rect 3067 3048 3120 3082
rect 3067 3014 3078 3048
rect 3112 3014 3120 3048
rect 3067 2980 3120 3014
rect 3067 2946 3078 2980
rect 3112 2946 3120 2980
rect 3067 2876 3120 2946
rect 3180 3864 3233 3876
rect 3180 3830 3188 3864
rect 3222 3830 3233 3864
rect 3180 3796 3233 3830
rect 3180 3762 3188 3796
rect 3222 3762 3233 3796
rect 3180 3728 3233 3762
rect 3180 3694 3188 3728
rect 3222 3694 3233 3728
rect 3180 3660 3233 3694
rect 3180 3626 3188 3660
rect 3222 3626 3233 3660
rect 3180 3592 3233 3626
rect 3180 3558 3188 3592
rect 3222 3558 3233 3592
rect 3180 3524 3233 3558
rect 3180 3490 3188 3524
rect 3222 3490 3233 3524
rect 3180 3456 3233 3490
rect 3180 3422 3188 3456
rect 3222 3422 3233 3456
rect 3180 3388 3233 3422
rect 3180 3354 3188 3388
rect 3222 3354 3233 3388
rect 3180 3320 3233 3354
rect 3180 3286 3188 3320
rect 3222 3286 3233 3320
rect 3180 3252 3233 3286
rect 3180 3218 3188 3252
rect 3222 3218 3233 3252
rect 3180 3184 3233 3218
rect 3180 3150 3188 3184
rect 3222 3150 3233 3184
rect 3180 3116 3233 3150
rect 3180 3082 3188 3116
rect 3222 3082 3233 3116
rect 3180 3048 3233 3082
rect 3180 3014 3188 3048
rect 3222 3014 3233 3048
rect 3180 2980 3233 3014
rect 3180 2946 3188 2980
rect 3222 2946 3233 2980
rect 3180 2876 3233 2946
rect 3333 3864 3389 3876
rect 3333 3830 3344 3864
rect 3378 3830 3389 3864
rect 3333 3796 3389 3830
rect 3333 3762 3344 3796
rect 3378 3762 3389 3796
rect 3333 3728 3389 3762
rect 3333 3694 3344 3728
rect 3378 3694 3389 3728
rect 3333 3660 3389 3694
rect 3333 3626 3344 3660
rect 3378 3626 3389 3660
rect 3333 3592 3389 3626
rect 3333 3558 3344 3592
rect 3378 3558 3389 3592
rect 3333 3524 3389 3558
rect 3333 3490 3344 3524
rect 3378 3490 3389 3524
rect 3333 3456 3389 3490
rect 3333 3422 3344 3456
rect 3378 3422 3389 3456
rect 3333 3388 3389 3422
rect 3333 3354 3344 3388
rect 3378 3354 3389 3388
rect 3333 3320 3389 3354
rect 3333 3286 3344 3320
rect 3378 3286 3389 3320
rect 3333 3252 3389 3286
rect 3333 3218 3344 3252
rect 3378 3218 3389 3252
rect 3333 3184 3389 3218
rect 3333 3150 3344 3184
rect 3378 3150 3389 3184
rect 3333 3116 3389 3150
rect 3333 3082 3344 3116
rect 3378 3082 3389 3116
rect 3333 3048 3389 3082
rect 3333 3014 3344 3048
rect 3378 3014 3389 3048
rect 3333 2980 3389 3014
rect 3333 2946 3344 2980
rect 3378 2946 3389 2980
rect 3333 2876 3389 2946
rect 3489 3864 3545 3876
rect 3489 3830 3500 3864
rect 3534 3830 3545 3864
rect 3489 3796 3545 3830
rect 3489 3762 3500 3796
rect 3534 3762 3545 3796
rect 3489 3728 3545 3762
rect 3489 3694 3500 3728
rect 3534 3694 3545 3728
rect 3489 3660 3545 3694
rect 3489 3626 3500 3660
rect 3534 3626 3545 3660
rect 3489 3592 3545 3626
rect 3489 3558 3500 3592
rect 3534 3558 3545 3592
rect 3489 3524 3545 3558
rect 3489 3490 3500 3524
rect 3534 3490 3545 3524
rect 3489 3456 3545 3490
rect 3489 3422 3500 3456
rect 3534 3422 3545 3456
rect 3489 3388 3545 3422
rect 3489 3354 3500 3388
rect 3534 3354 3545 3388
rect 3489 3320 3545 3354
rect 3489 3286 3500 3320
rect 3534 3286 3545 3320
rect 3489 3252 3545 3286
rect 3489 3218 3500 3252
rect 3534 3218 3545 3252
rect 3489 3184 3545 3218
rect 3489 3150 3500 3184
rect 3534 3150 3545 3184
rect 3489 3116 3545 3150
rect 3489 3082 3500 3116
rect 3534 3082 3545 3116
rect 3489 3048 3545 3082
rect 3489 3014 3500 3048
rect 3534 3014 3545 3048
rect 3489 2980 3545 3014
rect 3489 2946 3500 2980
rect 3534 2946 3545 2980
rect 3489 2876 3545 2946
rect 3645 3864 3701 3876
rect 3645 3830 3656 3864
rect 3690 3830 3701 3864
rect 3645 3796 3701 3830
rect 3645 3762 3656 3796
rect 3690 3762 3701 3796
rect 3645 3728 3701 3762
rect 3645 3694 3656 3728
rect 3690 3694 3701 3728
rect 3645 3660 3701 3694
rect 3645 3626 3656 3660
rect 3690 3626 3701 3660
rect 3645 3592 3701 3626
rect 3645 3558 3656 3592
rect 3690 3558 3701 3592
rect 3645 3524 3701 3558
rect 3645 3490 3656 3524
rect 3690 3490 3701 3524
rect 3645 3456 3701 3490
rect 3645 3422 3656 3456
rect 3690 3422 3701 3456
rect 3645 3388 3701 3422
rect 3645 3354 3656 3388
rect 3690 3354 3701 3388
rect 3645 3320 3701 3354
rect 3645 3286 3656 3320
rect 3690 3286 3701 3320
rect 3645 3252 3701 3286
rect 3645 3218 3656 3252
rect 3690 3218 3701 3252
rect 3645 3184 3701 3218
rect 3645 3150 3656 3184
rect 3690 3150 3701 3184
rect 3645 3116 3701 3150
rect 3645 3082 3656 3116
rect 3690 3082 3701 3116
rect 3645 3048 3701 3082
rect 3645 3014 3656 3048
rect 3690 3014 3701 3048
rect 3645 2980 3701 3014
rect 3645 2946 3656 2980
rect 3690 2946 3701 2980
rect 3645 2876 3701 2946
rect 3801 3864 3857 3876
rect 3801 3830 3812 3864
rect 3846 3830 3857 3864
rect 3801 3796 3857 3830
rect 3801 3762 3812 3796
rect 3846 3762 3857 3796
rect 3801 3728 3857 3762
rect 3801 3694 3812 3728
rect 3846 3694 3857 3728
rect 3801 3660 3857 3694
rect 3801 3626 3812 3660
rect 3846 3626 3857 3660
rect 3801 3592 3857 3626
rect 3801 3558 3812 3592
rect 3846 3558 3857 3592
rect 3801 3524 3857 3558
rect 3801 3490 3812 3524
rect 3846 3490 3857 3524
rect 3801 3456 3857 3490
rect 3801 3422 3812 3456
rect 3846 3422 3857 3456
rect 3801 3388 3857 3422
rect 3801 3354 3812 3388
rect 3846 3354 3857 3388
rect 3801 3320 3857 3354
rect 3801 3286 3812 3320
rect 3846 3286 3857 3320
rect 3801 3252 3857 3286
rect 3801 3218 3812 3252
rect 3846 3218 3857 3252
rect 3801 3184 3857 3218
rect 3801 3150 3812 3184
rect 3846 3150 3857 3184
rect 3801 3116 3857 3150
rect 3801 3082 3812 3116
rect 3846 3082 3857 3116
rect 3801 3048 3857 3082
rect 3801 3014 3812 3048
rect 3846 3014 3857 3048
rect 3801 2980 3857 3014
rect 3801 2946 3812 2980
rect 3846 2946 3857 2980
rect 3801 2876 3857 2946
rect 3957 3864 4010 3876
rect 3957 3830 3968 3864
rect 4002 3830 4010 3864
rect 3957 3796 4010 3830
rect 3957 3762 3968 3796
rect 4002 3762 4010 3796
rect 3957 3728 4010 3762
rect 3957 3694 3968 3728
rect 4002 3694 4010 3728
rect 3957 3660 4010 3694
rect 3957 3626 3968 3660
rect 4002 3626 4010 3660
rect 3957 3592 4010 3626
rect 3957 3558 3968 3592
rect 4002 3558 4010 3592
rect 3957 3524 4010 3558
rect 3957 3490 3968 3524
rect 4002 3490 4010 3524
rect 3957 3456 4010 3490
rect 3957 3422 3968 3456
rect 4002 3422 4010 3456
rect 3957 3388 4010 3422
rect 3957 3354 3968 3388
rect 4002 3354 4010 3388
rect 3957 3320 4010 3354
rect 3957 3286 3968 3320
rect 4002 3286 4010 3320
rect 3957 3252 4010 3286
rect 3957 3218 3968 3252
rect 4002 3218 4010 3252
rect 3957 3184 4010 3218
rect 3957 3150 3968 3184
rect 4002 3150 4010 3184
rect 3957 3116 4010 3150
rect 3957 3082 3968 3116
rect 4002 3082 4010 3116
rect 3957 3048 4010 3082
rect 3957 3014 3968 3048
rect 4002 3014 4010 3048
rect 3957 2980 4010 3014
rect 3957 2946 3968 2980
rect 4002 2946 4010 2980
rect 3957 2876 4010 2946
<< mvndiffc >>
rect 1764 2434 1798 2468
rect 1832 2434 1866 2468
rect 1900 2434 1934 2468
rect 1968 2434 2002 2468
rect 2036 2434 2070 2468
rect 2104 2434 2138 2468
rect 2172 2434 2206 2468
rect 2240 2434 2274 2468
rect 2818 2434 2852 2468
rect 2886 2434 2920 2468
rect 2954 2434 2988 2468
rect 3022 2434 3056 2468
rect 3090 2434 3124 2468
rect 3158 2434 3192 2468
rect 3226 2434 3260 2468
rect 3294 2434 3328 2468
rect 3362 2434 3396 2468
rect 3430 2434 3464 2468
rect 3498 2434 3532 2468
rect 3566 2434 3600 2468
rect 3634 2434 3668 2468
rect 3702 2434 3736 2468
rect 1764 2278 1798 2312
rect 1832 2278 1866 2312
rect 1900 2278 1934 2312
rect 1968 2278 2002 2312
rect 2036 2278 2070 2312
rect 2104 2278 2138 2312
rect 2172 2278 2206 2312
rect 2240 2278 2274 2312
rect 1187 2183 1221 2217
rect 1255 2183 1289 2217
rect 1323 2183 1357 2217
rect 1391 2183 1425 2217
rect 2818 2278 2852 2312
rect 2886 2278 2920 2312
rect 2954 2278 2988 2312
rect 3022 2278 3056 2312
rect 3090 2278 3124 2312
rect 3158 2278 3192 2312
rect 3226 2278 3260 2312
rect 3294 2278 3328 2312
rect 3362 2278 3396 2312
rect 3430 2278 3464 2312
rect 3498 2278 3532 2312
rect 3566 2278 3600 2312
rect 3634 2278 3668 2312
rect 3702 2278 3736 2312
rect 1764 2122 1798 2156
rect 1832 2122 1866 2156
rect 1900 2122 1934 2156
rect 1968 2122 2002 2156
rect 2036 2122 2070 2156
rect 2104 2122 2138 2156
rect 2172 2122 2206 2156
rect 2240 2122 2274 2156
rect 1187 2027 1221 2061
rect 1255 2027 1289 2061
rect 1323 2027 1357 2061
rect 1391 2027 1425 2061
rect 2818 2122 2852 2156
rect 2886 2122 2920 2156
rect 2954 2122 2988 2156
rect 3022 2122 3056 2156
rect 3090 2122 3124 2156
rect 3158 2122 3192 2156
rect 3226 2122 3260 2156
rect 3294 2122 3328 2156
rect 3362 2122 3396 2156
rect 3430 2122 3464 2156
rect 3498 2122 3532 2156
rect 3566 2122 3600 2156
rect 3634 2122 3668 2156
rect 3702 2122 3736 2156
rect 1764 1966 1798 2000
rect 1832 1966 1866 2000
rect 1900 1966 1934 2000
rect 1968 1966 2002 2000
rect 2036 1966 2070 2000
rect 2104 1966 2138 2000
rect 2172 1966 2206 2000
rect 2240 1966 2274 2000
rect 2818 1966 2852 2000
rect 2886 1966 2920 2000
rect 2954 1966 2988 2000
rect 3022 1966 3056 2000
rect 3090 1966 3124 2000
rect 3158 1966 3192 2000
rect 3226 1966 3260 2000
rect 3294 1966 3328 2000
rect 3362 1966 3396 2000
rect 3430 1966 3464 2000
rect 3498 1966 3532 2000
rect 3566 1966 3600 2000
rect 3634 1966 3668 2000
rect 3702 1966 3736 2000
rect 1764 1810 1798 1844
rect 1832 1810 1866 1844
rect 1900 1810 1934 1844
rect 1968 1810 2002 1844
rect 2036 1810 2070 1844
rect 2104 1810 2138 1844
rect 2172 1810 2206 1844
rect 2240 1810 2274 1844
rect 580 1097 614 1131
rect 580 1029 614 1063
rect 580 961 614 995
rect 580 893 614 927
rect 580 825 614 859
rect 580 757 614 791
rect 580 689 614 723
rect 580 621 614 655
rect 580 553 614 587
rect 580 485 614 519
rect 580 417 614 451
rect 580 349 614 383
rect 580 281 614 315
rect 580 213 614 247
rect 736 1097 770 1131
rect 736 1029 770 1063
rect 736 961 770 995
rect 736 893 770 927
rect 736 825 770 859
rect 736 757 770 791
rect 736 689 770 723
rect 736 621 770 655
rect 736 553 770 587
rect 736 485 770 519
rect 736 417 770 451
rect 736 349 770 383
rect 736 281 770 315
rect 736 213 770 247
rect 892 1097 926 1131
rect 892 1029 926 1063
rect 892 961 926 995
rect 892 893 926 927
rect 892 825 926 859
rect 892 757 926 791
rect 892 689 926 723
rect 892 621 926 655
rect 892 553 926 587
rect 892 485 926 519
rect 892 417 926 451
rect 892 349 926 383
rect 892 281 926 315
rect 892 213 926 247
rect 1048 1097 1082 1131
rect 1048 1029 1082 1063
rect 1048 961 1082 995
rect 1048 893 1082 927
rect 1048 825 1082 859
rect 1048 757 1082 791
rect 1048 689 1082 723
rect 1048 621 1082 655
rect 1048 553 1082 587
rect 1048 485 1082 519
rect 1048 417 1082 451
rect 1048 349 1082 383
rect 1048 281 1082 315
rect 1048 213 1082 247
rect 1204 1097 1238 1131
rect 1204 1029 1238 1063
rect 1204 961 1238 995
rect 1204 893 1238 927
rect 1204 825 1238 859
rect 1204 757 1238 791
rect 1204 689 1238 723
rect 1204 621 1238 655
rect 1204 553 1238 587
rect 1204 485 1238 519
rect 1204 417 1238 451
rect 1204 349 1238 383
rect 1204 281 1238 315
rect 1204 213 1238 247
rect 1360 1097 1394 1131
rect 1360 1029 1394 1063
rect 1360 961 1394 995
rect 1360 893 1394 927
rect 1360 825 1394 859
rect 1360 757 1394 791
rect 1360 689 1394 723
rect 1360 621 1394 655
rect 1360 553 1394 587
rect 1360 485 1394 519
rect 1360 417 1394 451
rect 1360 349 1394 383
rect 1360 281 1394 315
rect 1360 213 1394 247
rect 1516 1097 1550 1131
rect 1516 1029 1550 1063
rect 1516 961 1550 995
rect 1516 893 1550 927
rect 1516 825 1550 859
rect 1516 757 1550 791
rect 1516 689 1550 723
rect 1516 621 1550 655
rect 1516 553 1550 587
rect 1516 485 1550 519
rect 1516 417 1550 451
rect 1516 349 1550 383
rect 1516 281 1550 315
rect 1516 213 1550 247
rect 1672 1097 1706 1131
rect 1672 1029 1706 1063
rect 1672 961 1706 995
rect 1672 893 1706 927
rect 1672 825 1706 859
rect 1672 757 1706 791
rect 1672 689 1706 723
rect 1672 621 1706 655
rect 1672 553 1706 587
rect 1672 485 1706 519
rect 1672 417 1706 451
rect 1672 349 1706 383
rect 1672 281 1706 315
rect 1672 213 1706 247
rect 1828 1097 1862 1131
rect 1828 1029 1862 1063
rect 1828 961 1862 995
rect 1828 893 1862 927
rect 1828 825 1862 859
rect 1828 757 1862 791
rect 1828 689 1862 723
rect 1828 621 1862 655
rect 1828 553 1862 587
rect 1828 485 1862 519
rect 1828 417 1862 451
rect 1828 349 1862 383
rect 1828 281 1862 315
rect 1828 213 1862 247
rect 1938 1097 1972 1131
rect 1938 1029 1972 1063
rect 1938 961 1972 995
rect 1938 893 1972 927
rect 1938 825 1972 859
rect 1938 757 1972 791
rect 1938 689 1972 723
rect 1938 621 1972 655
rect 1938 553 1972 587
rect 1938 485 1972 519
rect 1938 417 1972 451
rect 1938 349 1972 383
rect 1938 281 1972 315
rect 1938 213 1972 247
rect 2094 1097 2128 1131
rect 2094 1029 2128 1063
rect 2094 961 2128 995
rect 2094 893 2128 927
rect 2094 825 2128 859
rect 2094 757 2128 791
rect 2094 689 2128 723
rect 2094 621 2128 655
rect 2094 553 2128 587
rect 2094 485 2128 519
rect 2094 417 2128 451
rect 2094 349 2128 383
rect 2094 281 2128 315
rect 2094 213 2128 247
rect 2250 1097 2284 1131
rect 2250 1029 2284 1063
rect 2250 961 2284 995
rect 2250 893 2284 927
rect 2250 825 2284 859
rect 2250 757 2284 791
rect 2250 689 2284 723
rect 2250 621 2284 655
rect 2250 553 2284 587
rect 2250 485 2284 519
rect 2250 417 2284 451
rect 2250 349 2284 383
rect 2250 281 2284 315
rect 2250 213 2284 247
rect 2406 1097 2440 1131
rect 2406 1029 2440 1063
rect 2406 961 2440 995
rect 2406 893 2440 927
rect 2406 825 2440 859
rect 2406 757 2440 791
rect 2406 689 2440 723
rect 2406 621 2440 655
rect 2406 553 2440 587
rect 2406 485 2440 519
rect 2406 417 2440 451
rect 2406 349 2440 383
rect 2406 281 2440 315
rect 2406 213 2440 247
rect 2562 1097 2596 1131
rect 2562 1029 2596 1063
rect 2562 961 2596 995
rect 2562 893 2596 927
rect 2562 825 2596 859
rect 2562 757 2596 791
rect 2562 689 2596 723
rect 2562 621 2596 655
rect 2562 553 2596 587
rect 2562 485 2596 519
rect 2562 417 2596 451
rect 2562 349 2596 383
rect 2562 281 2596 315
rect 2562 213 2596 247
rect 2718 1097 2752 1131
rect 2718 1029 2752 1063
rect 2718 961 2752 995
rect 2718 893 2752 927
rect 2718 825 2752 859
rect 2718 757 2752 791
rect 2718 689 2752 723
rect 2718 621 2752 655
rect 2718 553 2752 587
rect 2718 485 2752 519
rect 2718 417 2752 451
rect 2718 349 2752 383
rect 2718 281 2752 315
rect 2718 213 2752 247
rect 2874 1097 2908 1131
rect 2874 1029 2908 1063
rect 2874 961 2908 995
rect 2874 893 2908 927
rect 2874 825 2908 859
rect 2874 757 2908 791
rect 2874 689 2908 723
rect 2874 621 2908 655
rect 2874 553 2908 587
rect 2874 485 2908 519
rect 2874 417 2908 451
rect 2874 349 2908 383
rect 2874 281 2908 315
rect 2874 213 2908 247
rect 3030 1097 3064 1131
rect 3030 1029 3064 1063
rect 3030 961 3064 995
rect 3030 893 3064 927
rect 3030 825 3064 859
rect 3030 757 3064 791
rect 3030 689 3064 723
rect 3030 621 3064 655
rect 3030 553 3064 587
rect 3030 485 3064 519
rect 3030 417 3064 451
rect 3030 349 3064 383
rect 3030 281 3064 315
rect 3030 213 3064 247
<< mvpdiffc >>
rect 1298 3830 1332 3864
rect 1298 3762 1332 3796
rect 1298 3694 1332 3728
rect 1298 3626 1332 3660
rect 1298 3558 1332 3592
rect 1298 3490 1332 3524
rect 1298 3422 1332 3456
rect 1298 3354 1332 3388
rect 1298 3286 1332 3320
rect 1298 3218 1332 3252
rect 610 3130 644 3164
rect 610 3062 644 3096
rect 610 2994 644 3028
rect 610 2926 644 2960
rect 766 3130 800 3164
rect 766 3062 800 3096
rect 766 2994 800 3028
rect 766 2926 800 2960
rect 922 3130 956 3164
rect 922 3062 956 3096
rect 922 2994 956 3028
rect 922 2926 956 2960
rect 1032 3130 1066 3164
rect 1032 3062 1066 3096
rect 1032 2994 1066 3028
rect 1032 2926 1066 2960
rect 1188 3130 1222 3164
rect 1188 3062 1222 3096
rect 1188 2994 1222 3028
rect 1188 2926 1222 2960
rect 1298 3150 1332 3184
rect 1298 3082 1332 3116
rect 1298 3014 1332 3048
rect 1298 2946 1332 2980
rect 1454 3830 1488 3864
rect 1454 3762 1488 3796
rect 1454 3694 1488 3728
rect 1454 3626 1488 3660
rect 1454 3558 1488 3592
rect 1454 3490 1488 3524
rect 1454 3422 1488 3456
rect 1454 3354 1488 3388
rect 1454 3286 1488 3320
rect 1454 3218 1488 3252
rect 1454 3150 1488 3184
rect 1454 3082 1488 3116
rect 1454 3014 1488 3048
rect 1454 2946 1488 2980
rect 1610 3830 1644 3864
rect 1610 3762 1644 3796
rect 1610 3694 1644 3728
rect 1610 3626 1644 3660
rect 1610 3558 1644 3592
rect 1610 3490 1644 3524
rect 1610 3422 1644 3456
rect 1610 3354 1644 3388
rect 1610 3286 1644 3320
rect 1610 3218 1644 3252
rect 1610 3150 1644 3184
rect 1610 3082 1644 3116
rect 1610 3014 1644 3048
rect 1610 2946 1644 2980
rect 1766 3830 1800 3864
rect 1766 3762 1800 3796
rect 1766 3694 1800 3728
rect 1766 3626 1800 3660
rect 1766 3558 1800 3592
rect 1766 3490 1800 3524
rect 1766 3422 1800 3456
rect 1766 3354 1800 3388
rect 1766 3286 1800 3320
rect 1766 3218 1800 3252
rect 1766 3150 1800 3184
rect 1766 3082 1800 3116
rect 1766 3014 1800 3048
rect 1766 2946 1800 2980
rect 1922 3830 1956 3864
rect 1922 3762 1956 3796
rect 1922 3694 1956 3728
rect 1922 3626 1956 3660
rect 1922 3558 1956 3592
rect 1922 3490 1956 3524
rect 1922 3422 1956 3456
rect 1922 3354 1956 3388
rect 1922 3286 1956 3320
rect 1922 3218 1956 3252
rect 1922 3150 1956 3184
rect 1922 3082 1956 3116
rect 1922 3014 1956 3048
rect 1922 2946 1956 2980
rect 2032 3830 2066 3864
rect 2032 3762 2066 3796
rect 2032 3694 2066 3728
rect 2032 3626 2066 3660
rect 2032 3558 2066 3592
rect 2032 3490 2066 3524
rect 2032 3422 2066 3456
rect 2032 3354 2066 3388
rect 2032 3286 2066 3320
rect 2032 3218 2066 3252
rect 2032 3150 2066 3184
rect 2032 3082 2066 3116
rect 2032 3014 2066 3048
rect 2032 2946 2066 2980
rect 2188 3830 2222 3864
rect 2188 3762 2222 3796
rect 2188 3694 2222 3728
rect 2188 3626 2222 3660
rect 2188 3558 2222 3592
rect 2188 3490 2222 3524
rect 2188 3422 2222 3456
rect 2188 3354 2222 3388
rect 2188 3286 2222 3320
rect 2188 3218 2222 3252
rect 2188 3150 2222 3184
rect 2188 3082 2222 3116
rect 2188 3014 2222 3048
rect 2188 2946 2222 2980
rect 2344 3830 2378 3864
rect 2344 3762 2378 3796
rect 2344 3694 2378 3728
rect 2344 3626 2378 3660
rect 2344 3558 2378 3592
rect 2344 3490 2378 3524
rect 2344 3422 2378 3456
rect 2344 3354 2378 3388
rect 2344 3286 2378 3320
rect 2344 3218 2378 3252
rect 2344 3150 2378 3184
rect 2344 3082 2378 3116
rect 2344 3014 2378 3048
rect 2344 2946 2378 2980
rect 2500 3830 2534 3864
rect 2500 3762 2534 3796
rect 2500 3694 2534 3728
rect 2500 3626 2534 3660
rect 2500 3558 2534 3592
rect 2500 3490 2534 3524
rect 2500 3422 2534 3456
rect 2500 3354 2534 3388
rect 2500 3286 2534 3320
rect 2500 3218 2534 3252
rect 2500 3150 2534 3184
rect 2500 3082 2534 3116
rect 2500 3014 2534 3048
rect 2500 2946 2534 2980
rect 2656 3830 2690 3864
rect 2656 3762 2690 3796
rect 2656 3694 2690 3728
rect 2656 3626 2690 3660
rect 2656 3558 2690 3592
rect 2656 3490 2690 3524
rect 2656 3422 2690 3456
rect 2656 3354 2690 3388
rect 2656 3286 2690 3320
rect 2656 3218 2690 3252
rect 2656 3150 2690 3184
rect 2656 3082 2690 3116
rect 2656 3014 2690 3048
rect 2656 2946 2690 2980
rect 2766 3830 2800 3864
rect 2766 3762 2800 3796
rect 2766 3694 2800 3728
rect 2766 3626 2800 3660
rect 2766 3558 2800 3592
rect 2766 3490 2800 3524
rect 2766 3422 2800 3456
rect 2766 3354 2800 3388
rect 2766 3286 2800 3320
rect 2766 3218 2800 3252
rect 2766 3150 2800 3184
rect 2766 3082 2800 3116
rect 2766 3014 2800 3048
rect 2766 2946 2800 2980
rect 2922 3830 2956 3864
rect 2922 3762 2956 3796
rect 2922 3694 2956 3728
rect 2922 3626 2956 3660
rect 2922 3558 2956 3592
rect 2922 3490 2956 3524
rect 2922 3422 2956 3456
rect 2922 3354 2956 3388
rect 2922 3286 2956 3320
rect 2922 3218 2956 3252
rect 2922 3150 2956 3184
rect 2922 3082 2956 3116
rect 2922 3014 2956 3048
rect 2922 2946 2956 2980
rect 3078 3830 3112 3864
rect 3078 3762 3112 3796
rect 3078 3694 3112 3728
rect 3078 3626 3112 3660
rect 3078 3558 3112 3592
rect 3078 3490 3112 3524
rect 3078 3422 3112 3456
rect 3078 3354 3112 3388
rect 3078 3286 3112 3320
rect 3078 3218 3112 3252
rect 3078 3150 3112 3184
rect 3078 3082 3112 3116
rect 3078 3014 3112 3048
rect 3078 2946 3112 2980
rect 3188 3830 3222 3864
rect 3188 3762 3222 3796
rect 3188 3694 3222 3728
rect 3188 3626 3222 3660
rect 3188 3558 3222 3592
rect 3188 3490 3222 3524
rect 3188 3422 3222 3456
rect 3188 3354 3222 3388
rect 3188 3286 3222 3320
rect 3188 3218 3222 3252
rect 3188 3150 3222 3184
rect 3188 3082 3222 3116
rect 3188 3014 3222 3048
rect 3188 2946 3222 2980
rect 3344 3830 3378 3864
rect 3344 3762 3378 3796
rect 3344 3694 3378 3728
rect 3344 3626 3378 3660
rect 3344 3558 3378 3592
rect 3344 3490 3378 3524
rect 3344 3422 3378 3456
rect 3344 3354 3378 3388
rect 3344 3286 3378 3320
rect 3344 3218 3378 3252
rect 3344 3150 3378 3184
rect 3344 3082 3378 3116
rect 3344 3014 3378 3048
rect 3344 2946 3378 2980
rect 3500 3830 3534 3864
rect 3500 3762 3534 3796
rect 3500 3694 3534 3728
rect 3500 3626 3534 3660
rect 3500 3558 3534 3592
rect 3500 3490 3534 3524
rect 3500 3422 3534 3456
rect 3500 3354 3534 3388
rect 3500 3286 3534 3320
rect 3500 3218 3534 3252
rect 3500 3150 3534 3184
rect 3500 3082 3534 3116
rect 3500 3014 3534 3048
rect 3500 2946 3534 2980
rect 3656 3830 3690 3864
rect 3656 3762 3690 3796
rect 3656 3694 3690 3728
rect 3656 3626 3690 3660
rect 3656 3558 3690 3592
rect 3656 3490 3690 3524
rect 3656 3422 3690 3456
rect 3656 3354 3690 3388
rect 3656 3286 3690 3320
rect 3656 3218 3690 3252
rect 3656 3150 3690 3184
rect 3656 3082 3690 3116
rect 3656 3014 3690 3048
rect 3656 2946 3690 2980
rect 3812 3830 3846 3864
rect 3812 3762 3846 3796
rect 3812 3694 3846 3728
rect 3812 3626 3846 3660
rect 3812 3558 3846 3592
rect 3812 3490 3846 3524
rect 3812 3422 3846 3456
rect 3812 3354 3846 3388
rect 3812 3286 3846 3320
rect 3812 3218 3846 3252
rect 3812 3150 3846 3184
rect 3812 3082 3846 3116
rect 3812 3014 3846 3048
rect 3812 2946 3846 2980
rect 3968 3830 4002 3864
rect 3968 3762 4002 3796
rect 3968 3694 4002 3728
rect 3968 3626 4002 3660
rect 3968 3558 4002 3592
rect 3968 3490 4002 3524
rect 3968 3422 4002 3456
rect 3968 3354 4002 3388
rect 3968 3286 4002 3320
rect 3968 3218 4002 3252
rect 3968 3150 4002 3184
rect 3968 3082 4002 3116
rect 3968 3014 4002 3048
rect 3968 2946 4002 2980
<< psubdiff >>
rect 893 2475 917 2509
rect 951 2475 986 2509
rect 1020 2475 1055 2509
rect 1089 2475 1124 2509
rect 1158 2475 1192 2509
rect 1226 2475 1260 2509
rect 1294 2475 1328 2509
rect 1362 2475 1396 2509
rect 1430 2475 1454 2509
rect 1642 2445 1676 2469
rect 1642 2375 1676 2411
rect 1642 2305 1676 2341
rect 1642 2234 1676 2271
rect 1642 2163 1676 2200
rect 1642 2092 1676 2129
rect 1642 2021 1676 2058
rect 1642 1950 1676 1987
rect 1642 1879 1676 1916
rect 1642 1821 1676 1845
<< mvpsubdiff >>
rect 3830 2445 3864 2469
rect 3830 2376 3864 2411
rect 3830 2306 3864 2342
rect 3830 2236 3864 2272
rect 3830 2166 3864 2202
rect 3830 2108 3864 2132
rect 594 91 618 125
rect 652 91 687 125
rect 721 91 756 125
rect 790 91 825 125
rect 859 91 894 125
rect 928 91 963 125
rect 997 91 1032 125
rect 1066 91 1101 125
rect 1135 91 1170 125
rect 1204 91 1239 125
rect 1273 91 1308 125
rect 1342 91 1377 125
rect 1411 91 1446 125
rect 1480 91 1515 125
rect 1549 91 1584 125
rect 1618 91 1653 125
rect 1687 91 1722 125
rect 1756 91 1791 125
rect 1825 91 1861 125
rect 1895 91 1931 125
rect 1965 91 2001 125
rect 2035 91 2071 125
rect 2105 91 2141 125
rect 2175 91 2211 125
rect 2245 91 2281 125
rect 2315 91 2351 125
rect 2385 91 2421 125
rect 2455 91 2491 125
rect 2525 91 2561 125
rect 2595 91 2631 125
rect 2665 91 2701 125
rect 2735 91 2771 125
rect 2805 91 2841 125
rect 2875 91 2911 125
rect 2945 91 2981 125
rect 3015 91 3039 125
<< mvnsubdiff >>
rect 603 3950 637 3984
rect 671 3950 705 3984
rect 739 3950 773 3984
rect 807 3950 841 3984
rect 875 3950 909 3984
rect 943 3950 977 3984
rect 1011 3950 1045 3984
rect 1079 3950 1113 3984
rect 1147 3950 1181 3984
rect 1215 3950 1249 3984
rect 1283 3950 1317 3984
rect 1351 3950 1385 3984
rect 1419 3950 1453 3984
rect 1487 3950 1521 3984
rect 1555 3950 1589 3984
rect 1623 3950 1657 3984
rect 1691 3950 1725 3984
rect 1759 3950 1793 3984
rect 1827 3950 1861 3984
rect 1895 3950 1929 3984
rect 1963 3950 1997 3984
rect 2031 3950 2065 3984
rect 2099 3950 2133 3984
rect 2167 3950 2201 3984
rect 2235 3950 2269 3984
rect 2303 3950 2337 3984
rect 2371 3950 2405 3984
rect 2439 3950 2473 3984
rect 2507 3950 2541 3984
rect 2575 3950 2609 3984
rect 2643 3950 2677 3984
rect 2711 3950 2745 3984
rect 2779 3950 2813 3984
rect 2847 3950 2881 3984
rect 2915 3950 2949 3984
rect 2983 3950 3017 3984
rect 3051 3950 3085 3984
rect 3119 3950 3153 3984
rect 3187 3950 3221 3984
rect 3255 3950 3289 3984
rect 3323 3950 3357 3984
rect 3391 3950 3425 3984
rect 3459 3950 3493 3984
rect 3527 3950 3561 3984
rect 3595 3950 3629 3984
rect 3663 3950 3697 3984
rect 3731 3950 3765 3984
rect 3799 3950 3833 3984
rect 3867 3950 3901 3984
rect 3935 3950 4009 3984
<< psubdiffcont >>
rect 917 2475 951 2509
rect 986 2475 1020 2509
rect 1055 2475 1089 2509
rect 1124 2475 1158 2509
rect 1192 2475 1226 2509
rect 1260 2475 1294 2509
rect 1328 2475 1362 2509
rect 1396 2475 1430 2509
rect 1642 2411 1676 2445
rect 1642 2341 1676 2375
rect 1642 2271 1676 2305
rect 1642 2200 1676 2234
rect 1642 2129 1676 2163
rect 1642 2058 1676 2092
rect 1642 1987 1676 2021
rect 1642 1916 1676 1950
rect 1642 1845 1676 1879
<< mvpsubdiffcont >>
rect 3830 2411 3864 2445
rect 3830 2342 3864 2376
rect 3830 2272 3864 2306
rect 3830 2202 3864 2236
rect 3830 2132 3864 2166
rect 618 91 652 125
rect 687 91 721 125
rect 756 91 790 125
rect 825 91 859 125
rect 894 91 928 125
rect 963 91 997 125
rect 1032 91 1066 125
rect 1101 91 1135 125
rect 1170 91 1204 125
rect 1239 91 1273 125
rect 1308 91 1342 125
rect 1377 91 1411 125
rect 1446 91 1480 125
rect 1515 91 1549 125
rect 1584 91 1618 125
rect 1653 91 1687 125
rect 1722 91 1756 125
rect 1791 91 1825 125
rect 1861 91 1895 125
rect 1931 91 1965 125
rect 2001 91 2035 125
rect 2071 91 2105 125
rect 2141 91 2175 125
rect 2211 91 2245 125
rect 2281 91 2315 125
rect 2351 91 2385 125
rect 2421 91 2455 125
rect 2491 91 2525 125
rect 2561 91 2595 125
rect 2631 91 2665 125
rect 2701 91 2735 125
rect 2771 91 2805 125
rect 2841 91 2875 125
rect 2911 91 2945 125
rect 2981 91 3015 125
<< mvnsubdiffcont >>
rect 637 3950 671 3984
rect 705 3950 739 3984
rect 773 3950 807 3984
rect 841 3950 875 3984
rect 909 3950 943 3984
rect 977 3950 1011 3984
rect 1045 3950 1079 3984
rect 1113 3950 1147 3984
rect 1181 3950 1215 3984
rect 1249 3950 1283 3984
rect 1317 3950 1351 3984
rect 1385 3950 1419 3984
rect 1453 3950 1487 3984
rect 1521 3950 1555 3984
rect 1589 3950 1623 3984
rect 1657 3950 1691 3984
rect 1725 3950 1759 3984
rect 1793 3950 1827 3984
rect 1861 3950 1895 3984
rect 1929 3950 1963 3984
rect 1997 3950 2031 3984
rect 2065 3950 2099 3984
rect 2133 3950 2167 3984
rect 2201 3950 2235 3984
rect 2269 3950 2303 3984
rect 2337 3950 2371 3984
rect 2405 3950 2439 3984
rect 2473 3950 2507 3984
rect 2541 3950 2575 3984
rect 2609 3950 2643 3984
rect 2677 3950 2711 3984
rect 2745 3950 2779 3984
rect 2813 3950 2847 3984
rect 2881 3950 2915 3984
rect 2949 3950 2983 3984
rect 3017 3950 3051 3984
rect 3085 3950 3119 3984
rect 3153 3950 3187 3984
rect 3221 3950 3255 3984
rect 3289 3950 3323 3984
rect 3357 3950 3391 3984
rect 3425 3950 3459 3984
rect 3493 3950 3527 3984
rect 3561 3950 3595 3984
rect 3629 3950 3663 3984
rect 3697 3950 3731 3984
rect 3765 3950 3799 3984
rect 3833 3950 3867 3984
rect 3901 3950 3935 3984
<< poly >>
rect 1343 3876 1443 3908
rect 1499 3876 1599 3908
rect 1655 3876 1755 3908
rect 1811 3876 1911 3908
rect 2077 3876 2177 3908
rect 2233 3876 2333 3908
rect 2389 3876 2489 3908
rect 2545 3876 2645 3908
rect 2811 3876 2911 3908
rect 2967 3876 3067 3908
rect 3233 3876 3333 3908
rect 3389 3876 3489 3908
rect 3545 3876 3645 3908
rect 3701 3876 3801 3908
rect 3857 3876 3957 3908
rect 655 3176 755 3208
rect 811 3176 911 3208
rect 1077 3176 1177 3208
rect 655 2844 755 2876
rect 621 2828 755 2844
rect 621 2794 637 2828
rect 671 2794 705 2828
rect 739 2794 755 2828
rect 621 2778 755 2794
rect 811 2844 911 2876
rect 1077 2844 1177 2876
rect 811 2828 1177 2844
rect 811 2794 827 2828
rect 861 2794 902 2828
rect 936 2794 977 2828
rect 1011 2794 1052 2828
rect 1086 2794 1127 2828
rect 1161 2794 1177 2828
rect 811 2778 1177 2794
rect 1343 2844 1443 2876
rect 1499 2844 1599 2876
rect 1343 2828 1599 2844
rect 1343 2794 1359 2828
rect 1393 2794 1454 2828
rect 1488 2794 1549 2828
rect 1583 2794 1599 2828
rect 1343 2778 1599 2794
rect 1655 2844 1755 2876
rect 1811 2844 1911 2876
rect 1655 2828 1911 2844
rect 1655 2794 1671 2828
rect 1705 2794 1766 2828
rect 1800 2794 1861 2828
rect 1895 2794 1911 2828
rect 1655 2778 1911 2794
rect 2077 2844 2177 2876
rect 2233 2844 2333 2876
rect 2077 2828 2333 2844
rect 2077 2794 2093 2828
rect 2127 2794 2188 2828
rect 2222 2794 2283 2828
rect 2317 2794 2333 2828
rect 2077 2778 2333 2794
rect 2389 2844 2489 2876
rect 2545 2844 2645 2876
rect 2811 2844 2911 2876
rect 2389 2828 2645 2844
rect 2389 2794 2405 2828
rect 2439 2794 2500 2828
rect 2534 2794 2595 2828
rect 2629 2794 2645 2828
rect 2389 2778 2645 2794
rect 2777 2828 2911 2844
rect 2777 2794 2793 2828
rect 2827 2794 2861 2828
rect 2895 2794 2911 2828
rect 2777 2778 2911 2794
rect 2967 2844 3067 2876
rect 3233 2844 3333 2876
rect 3389 2844 3489 2876
rect 3545 2844 3645 2876
rect 3701 2844 3801 2876
rect 3857 2844 3957 2876
rect 2967 2828 3101 2844
rect 2967 2794 2983 2828
rect 3017 2794 3051 2828
rect 3085 2794 3101 2828
rect 2967 2778 3101 2794
rect 3233 2828 3958 2844
rect 3233 2794 3249 2828
rect 3283 2794 3323 2828
rect 3357 2794 3397 2828
rect 3431 2794 3470 2828
rect 3504 2794 3543 2828
rect 3577 2794 3616 2828
rect 3650 2794 3689 2828
rect 3723 2794 3762 2828
rect 3796 2794 3835 2828
rect 3869 2794 3908 2828
rect 3942 2794 3958 2828
rect 3233 2778 3958 2794
rect 1720 2323 1752 2423
rect 2352 2388 2518 2423
rect 2352 2354 2400 2388
rect 2434 2354 2468 2388
rect 2502 2354 2518 2388
rect 2352 2323 2518 2354
rect 2650 2407 2748 2423
rect 2650 2373 2666 2407
rect 2700 2373 2748 2407
rect 2650 2338 2748 2373
rect 2650 2304 2666 2338
rect 2700 2323 2748 2338
rect 3748 2323 3780 2423
rect 2700 2304 2716 2323
rect 2650 2269 2716 2304
rect 1507 2202 1573 2218
rect 1507 2172 1523 2202
rect 1143 2072 1175 2172
rect 1475 2168 1523 2172
rect 1557 2168 1573 2202
rect 1475 2122 1573 2168
rect 1475 2088 1523 2122
rect 1557 2088 1573 2122
rect 1475 2072 1573 2088
rect 1720 2167 1752 2267
rect 2352 2232 2518 2267
rect 2352 2198 2400 2232
rect 2434 2198 2468 2232
rect 2502 2198 2518 2232
rect 2352 2167 2518 2198
rect 2650 2235 2666 2269
rect 2700 2267 2716 2269
rect 2700 2235 2748 2267
rect 2650 2200 2748 2235
rect 2650 2166 2666 2200
rect 2700 2167 2748 2200
rect 3748 2167 3780 2267
rect 2700 2166 2716 2167
rect 2650 2131 2716 2166
rect 1720 2011 1752 2111
rect 2352 2076 2518 2111
rect 2352 2042 2400 2076
rect 2434 2042 2468 2076
rect 2502 2042 2518 2076
rect 2352 2011 2518 2042
rect 2650 2097 2666 2131
rect 2700 2111 2716 2131
rect 2700 2097 2748 2111
rect 2650 2061 2748 2097
rect 2650 2027 2666 2061
rect 2700 2027 2748 2061
rect 2650 2011 2748 2027
rect 3748 2011 3780 2111
rect 1720 1855 1752 1955
rect 2352 1925 2518 1955
rect 2352 1891 2400 1925
rect 2434 1891 2468 1925
rect 2502 1891 2518 1925
rect 2352 1855 2518 1891
rect 591 1283 725 1299
rect 591 1249 607 1283
rect 641 1249 675 1283
rect 709 1249 725 1283
rect 591 1233 725 1249
rect 625 1201 725 1233
rect 781 1283 1193 1299
rect 781 1249 797 1283
rect 831 1249 867 1283
rect 901 1249 936 1283
rect 970 1249 1005 1283
rect 1039 1249 1074 1283
rect 1108 1249 1143 1283
rect 1177 1249 1193 1283
rect 781 1233 1193 1249
rect 781 1201 881 1233
rect 937 1201 1037 1233
rect 1093 1201 1193 1233
rect 1249 1283 1817 1299
rect 1249 1249 1265 1283
rect 1299 1249 1337 1283
rect 1371 1249 1409 1283
rect 1443 1249 1481 1283
rect 1515 1249 1553 1283
rect 1587 1249 1625 1283
rect 1659 1249 1696 1283
rect 1730 1249 1767 1283
rect 1801 1249 1817 1283
rect 1249 1233 1817 1249
rect 1249 1201 1349 1233
rect 1405 1201 1505 1233
rect 1561 1201 1661 1233
rect 1717 1201 1817 1233
rect 1983 1283 2551 1299
rect 1983 1249 1999 1283
rect 2033 1249 2071 1283
rect 2105 1249 2143 1283
rect 2177 1249 2215 1283
rect 2249 1249 2287 1283
rect 2321 1249 2359 1283
rect 2393 1249 2430 1283
rect 2464 1249 2501 1283
rect 2535 1249 2551 1283
rect 1983 1233 2551 1249
rect 1983 1201 2083 1233
rect 2139 1201 2239 1233
rect 2295 1201 2395 1233
rect 2451 1201 2551 1233
rect 2607 1283 3019 1299
rect 2607 1249 2623 1283
rect 2657 1249 2693 1283
rect 2727 1249 2762 1283
rect 2796 1249 2831 1283
rect 2865 1249 2900 1283
rect 2934 1249 2969 1283
rect 3003 1249 3019 1283
rect 2607 1233 3019 1249
rect 2607 1201 2707 1233
rect 2763 1201 2863 1233
rect 2919 1201 3019 1233
rect 625 169 725 201
rect 781 169 881 201
rect 937 169 1037 201
rect 1093 169 1193 201
rect 1249 169 1349 201
rect 1405 169 1505 201
rect 1561 169 1661 201
rect 1717 169 1817 201
rect 1983 169 2083 201
rect 2139 169 2239 201
rect 2295 169 2395 201
rect 2451 169 2551 201
rect 2607 169 2707 201
rect 2763 169 2863 201
rect 2919 169 3019 201
<< polycont >>
rect 637 2794 671 2828
rect 705 2794 739 2828
rect 827 2794 861 2828
rect 902 2794 936 2828
rect 977 2794 1011 2828
rect 1052 2794 1086 2828
rect 1127 2794 1161 2828
rect 1359 2794 1393 2828
rect 1454 2794 1488 2828
rect 1549 2794 1583 2828
rect 1671 2794 1705 2828
rect 1766 2794 1800 2828
rect 1861 2794 1895 2828
rect 2093 2794 2127 2828
rect 2188 2794 2222 2828
rect 2283 2794 2317 2828
rect 2405 2794 2439 2828
rect 2500 2794 2534 2828
rect 2595 2794 2629 2828
rect 2793 2794 2827 2828
rect 2861 2794 2895 2828
rect 2983 2794 3017 2828
rect 3051 2794 3085 2828
rect 3249 2794 3283 2828
rect 3323 2794 3357 2828
rect 3397 2794 3431 2828
rect 3470 2794 3504 2828
rect 3543 2794 3577 2828
rect 3616 2794 3650 2828
rect 3689 2794 3723 2828
rect 3762 2794 3796 2828
rect 3835 2794 3869 2828
rect 3908 2794 3942 2828
rect 2400 2354 2434 2388
rect 2468 2354 2502 2388
rect 2666 2373 2700 2407
rect 2666 2304 2700 2338
rect 1523 2168 1557 2202
rect 1523 2088 1557 2122
rect 2400 2198 2434 2232
rect 2468 2198 2502 2232
rect 2666 2235 2700 2269
rect 2666 2166 2700 2200
rect 2400 2042 2434 2076
rect 2468 2042 2502 2076
rect 2666 2097 2700 2131
rect 2666 2027 2700 2061
rect 2400 1891 2434 1925
rect 2468 1891 2502 1925
rect 607 1249 641 1283
rect 675 1249 709 1283
rect 797 1249 831 1283
rect 867 1249 901 1283
rect 936 1249 970 1283
rect 1005 1249 1039 1283
rect 1074 1249 1108 1283
rect 1143 1249 1177 1283
rect 1265 1249 1299 1283
rect 1337 1249 1371 1283
rect 1409 1249 1443 1283
rect 1481 1249 1515 1283
rect 1553 1249 1587 1283
rect 1625 1249 1659 1283
rect 1696 1249 1730 1283
rect 1767 1249 1801 1283
rect 1999 1249 2033 1283
rect 2071 1249 2105 1283
rect 2143 1249 2177 1283
rect 2215 1249 2249 1283
rect 2287 1249 2321 1283
rect 2359 1249 2393 1283
rect 2430 1249 2464 1283
rect 2501 1249 2535 1283
rect 2623 1249 2657 1283
rect 2693 1249 2727 1283
rect 2762 1249 2796 1283
rect 2831 1249 2865 1283
rect 2900 1249 2934 1283
rect 2969 1249 3003 1283
<< locali >>
rect 671 3950 677 3984
rect 739 3950 751 3984
rect 807 3950 825 3984
rect 875 3950 899 3984
rect 943 3950 973 3984
rect 1011 3950 1045 3984
rect 1081 3950 1113 3984
rect 1155 3950 1181 3984
rect 1229 3950 1249 3984
rect 1303 3950 1317 3984
rect 1377 3950 1385 3984
rect 1451 3950 1453 3984
rect 1487 3950 1491 3984
rect 1555 3950 1565 3984
rect 1623 3950 1639 3984
rect 1691 3950 1712 3984
rect 1759 3950 1785 3984
rect 1827 3950 1858 3984
rect 1895 3950 1929 3984
rect 1965 3950 1997 3984
rect 2038 3950 2065 3984
rect 2111 3950 2133 3984
rect 2184 3950 2201 3984
rect 2257 3950 2269 3984
rect 2330 3950 2337 3984
rect 2403 3950 2405 3984
rect 2439 3950 2442 3984
rect 2507 3950 2515 3984
rect 2575 3950 2588 3984
rect 2643 3950 2661 3984
rect 2711 3950 2734 3984
rect 2779 3950 2807 3984
rect 2847 3950 2880 3984
rect 2915 3950 2949 3984
rect 2987 3950 3017 3984
rect 3060 3950 3085 3984
rect 3133 3950 3153 3984
rect 3206 3950 3221 3984
rect 3279 3950 3289 3984
rect 3352 3950 3357 3984
rect 3459 3950 3464 3984
rect 3527 3950 3537 3984
rect 3595 3950 3610 3984
rect 3663 3950 3683 3984
rect 3731 3950 3756 3984
rect 3799 3950 3829 3984
rect 3867 3950 3901 3984
rect 3936 3950 3975 3984
rect 1298 3864 1332 3880
rect 1298 3796 1332 3830
rect 1298 3728 1332 3762
rect 1298 3660 1332 3677
rect 1298 3592 1332 3603
rect 1298 3524 1332 3529
rect 1298 3489 1332 3490
rect 1298 3414 1332 3422
rect 1298 3339 1332 3354
rect 1298 3264 1332 3286
rect 610 3164 644 3166
rect 610 3096 644 3130
rect 610 3028 644 3036
rect 610 2960 644 2994
rect 610 2910 644 2926
rect 766 3164 800 3166
rect 766 3120 800 3130
rect 766 3040 800 3062
rect 766 2960 800 2994
rect 766 2910 800 2926
rect 922 3164 956 3166
rect 922 3123 956 3130
rect 922 3045 956 3062
rect 922 2960 956 2994
rect 922 2910 956 2926
rect 1298 3189 1332 3218
rect 1032 3164 1066 3166
rect 1032 3112 1066 3130
rect 1032 3028 1066 3062
rect 1032 2960 1066 2989
rect 1032 2910 1066 2926
rect 1188 3164 1222 3180
rect 1188 3096 1222 3130
rect 1188 3028 1222 3031
rect 1188 2960 1222 2994
rect 1298 3116 1332 3150
rect 1298 3048 1332 3080
rect 1298 2980 1332 3005
rect 1454 3864 1488 3880
rect 1454 3796 1488 3830
rect 1454 3728 1488 3762
rect 1454 3660 1488 3677
rect 1454 3592 1488 3603
rect 1454 3524 1488 3529
rect 1454 3489 1488 3490
rect 1454 3415 1488 3422
rect 1454 3340 1488 3354
rect 1454 3265 1488 3286
rect 1454 3190 1488 3218
rect 1454 3116 1488 3150
rect 1454 3048 1488 3081
rect 1454 2980 1488 3006
rect 1454 2930 1488 2946
rect 1610 3864 1644 3880
rect 1610 3796 1644 3830
rect 1610 3728 1644 3762
rect 1610 3660 1644 3677
rect 1610 3592 1644 3603
rect 1610 3524 1644 3529
rect 1610 3489 1644 3490
rect 1610 3414 1644 3422
rect 1610 3339 1644 3354
rect 1610 3264 1644 3286
rect 1610 3189 1644 3218
rect 1610 3116 1644 3150
rect 1610 3048 1644 3080
rect 1610 2980 1644 3005
rect 1766 3804 1800 3830
rect 1766 3728 1800 3762
rect 1766 3660 1800 3694
rect 1766 3592 1800 3618
rect 1766 3524 1800 3542
rect 1766 3456 1800 3466
rect 1766 3388 1800 3390
rect 1766 3348 1800 3354
rect 1766 3271 1800 3286
rect 1766 3194 1800 3218
rect 1766 3117 1800 3150
rect 1766 3048 1800 3082
rect 1766 2980 1800 3006
rect 1766 2930 1800 2946
rect 1922 3864 1956 3880
rect 1922 3796 1956 3830
rect 1922 3728 1956 3762
rect 1922 3660 1956 3677
rect 1922 3592 1956 3603
rect 1922 3524 1956 3529
rect 1922 3489 1956 3490
rect 1922 3414 1956 3422
rect 1922 3339 1956 3354
rect 1922 3264 1956 3286
rect 1922 3189 1956 3218
rect 1922 3116 1956 3150
rect 1922 3048 1956 3080
rect 1922 2980 1956 3005
rect 2032 3864 2066 3880
rect 2032 3796 2066 3830
rect 2032 3728 2066 3762
rect 2032 3660 2066 3677
rect 2032 3592 2066 3603
rect 2032 3524 2066 3529
rect 2032 3489 2066 3490
rect 2032 3414 2066 3422
rect 2032 3339 2066 3354
rect 2032 3264 2066 3286
rect 2032 3189 2066 3218
rect 2032 3116 2066 3150
rect 2032 3048 2066 3080
rect 2032 2980 2066 3005
rect 2188 3804 2222 3830
rect 2188 3728 2222 3762
rect 2188 3660 2222 3694
rect 2188 3592 2222 3618
rect 2188 3524 2222 3542
rect 2188 3456 2222 3466
rect 2188 3388 2222 3390
rect 2188 3348 2222 3354
rect 2188 3271 2222 3286
rect 2188 3194 2222 3218
rect 2188 3117 2222 3150
rect 2188 3048 2222 3082
rect 2188 2980 2222 3006
rect 2188 2930 2222 2946
rect 2344 3864 2378 3880
rect 2344 3796 2378 3830
rect 2344 3728 2378 3762
rect 2344 3660 2378 3677
rect 2344 3592 2378 3603
rect 2344 3524 2378 3529
rect 2344 3489 2378 3490
rect 2344 3414 2378 3422
rect 2344 3339 2378 3354
rect 2344 3264 2378 3286
rect 2344 3189 2378 3218
rect 2344 3116 2378 3150
rect 2344 3048 2378 3080
rect 2344 2980 2378 3005
rect 2500 3864 2534 3880
rect 2500 3796 2534 3830
rect 2500 3728 2534 3762
rect 2500 3660 2534 3677
rect 2500 3592 2534 3603
rect 2500 3524 2534 3529
rect 2500 3489 2534 3490
rect 2500 3415 2534 3422
rect 2500 3340 2534 3354
rect 2500 3265 2534 3286
rect 2500 3190 2534 3218
rect 2500 3116 2534 3150
rect 2500 3048 2534 3081
rect 2500 2980 2534 3006
rect 2500 2930 2534 2946
rect 2656 3864 2690 3880
rect 2656 3796 2690 3830
rect 2656 3728 2690 3762
rect 2656 3660 2690 3677
rect 2656 3592 2690 3603
rect 2656 3524 2690 3529
rect 2656 3489 2690 3490
rect 2656 3414 2690 3422
rect 2656 3339 2690 3354
rect 2656 3264 2690 3286
rect 2656 3189 2690 3218
rect 2656 3116 2690 3150
rect 2656 3048 2690 3080
rect 2656 2980 2690 3005
rect 2766 3864 2800 3880
rect 2766 3796 2800 3830
rect 2766 3728 2800 3762
rect 2766 3660 2800 3677
rect 2766 3592 2800 3603
rect 2766 3524 2800 3529
rect 2766 3489 2800 3490
rect 2766 3415 2800 3422
rect 2766 3340 2800 3354
rect 2766 3265 2800 3286
rect 2766 3190 2800 3218
rect 2766 3116 2800 3150
rect 2766 3048 2800 3081
rect 2766 2980 2800 3006
rect 2766 2930 2800 2946
rect 2922 3864 2956 3880
rect 2922 3796 2956 3830
rect 2922 3728 2956 3762
rect 2922 3660 2956 3677
rect 2922 3592 2956 3603
rect 2922 3524 2956 3529
rect 2922 3489 2956 3490
rect 2922 3415 2956 3422
rect 2922 3340 2956 3354
rect 2922 3265 2956 3286
rect 2922 3190 2956 3218
rect 2922 3116 2956 3150
rect 2922 3048 2956 3081
rect 2922 2980 2956 3006
rect 2922 2930 2956 2946
rect 3078 3803 3112 3830
rect 3078 3728 3112 3762
rect 3078 3660 3112 3691
rect 3078 3592 3112 3613
rect 3078 3524 3112 3535
rect 3078 3456 3112 3457
rect 3078 3413 3112 3422
rect 3078 3335 3112 3354
rect 3078 3257 3112 3286
rect 3078 3184 3112 3218
rect 3078 3116 3112 3145
rect 3078 3048 3112 3067
rect 3078 2980 3112 2989
rect 3078 2930 3112 2946
rect 3188 3864 3222 3880
rect 3188 3796 3222 3830
rect 3188 3728 3222 3762
rect 3188 3660 3222 3677
rect 3188 3592 3222 3603
rect 3188 3524 3222 3529
rect 3188 3488 3222 3490
rect 3188 3413 3222 3422
rect 3188 3338 3222 3354
rect 3188 3263 3222 3286
rect 3188 3188 3222 3218
rect 3188 3116 3222 3150
rect 3188 3048 3222 3079
rect 3188 2980 3222 3004
rect 3344 3805 3378 3830
rect 3344 3730 3378 3762
rect 3344 3660 3378 3694
rect 3344 3592 3378 3621
rect 3344 3524 3378 3546
rect 3344 3456 3378 3471
rect 3344 3388 3378 3396
rect 3344 3320 3378 3321
rect 3344 3280 3378 3286
rect 3344 3204 3378 3218
rect 3344 3128 3378 3150
rect 3344 3052 3378 3082
rect 3344 2980 3378 3014
rect 3344 2930 3378 2946
rect 3500 3864 3534 3880
rect 3500 3796 3534 3830
rect 3500 3728 3534 3762
rect 3500 3660 3534 3677
rect 3500 3592 3534 3603
rect 3500 3524 3534 3529
rect 3500 3488 3534 3490
rect 3500 3413 3534 3422
rect 3500 3338 3534 3354
rect 3500 3263 3534 3286
rect 3500 3188 3534 3218
rect 3500 3116 3534 3150
rect 3500 3048 3534 3079
rect 3500 2980 3534 3004
rect 3656 3805 3690 3830
rect 3656 3730 3690 3762
rect 3656 3660 3690 3694
rect 3656 3592 3690 3621
rect 3656 3524 3690 3546
rect 3656 3456 3690 3471
rect 3656 3388 3690 3396
rect 3656 3320 3690 3321
rect 3656 3280 3690 3286
rect 3656 3204 3690 3218
rect 3656 3128 3690 3150
rect 3656 3052 3690 3082
rect 3656 2980 3690 3014
rect 3656 2930 3690 2946
rect 3812 3864 3846 3880
rect 3812 3796 3846 3830
rect 3812 3728 3846 3762
rect 3812 3660 3846 3677
rect 3812 3592 3846 3603
rect 3812 3524 3846 3529
rect 3812 3488 3846 3490
rect 3812 3413 3846 3422
rect 3812 3338 3846 3354
rect 3812 3263 3846 3286
rect 3812 3188 3846 3218
rect 3812 3116 3846 3150
rect 3812 3048 3846 3079
rect 3812 2980 3846 3004
rect 3968 3805 4002 3830
rect 3968 3730 4002 3762
rect 3968 3660 4002 3694
rect 3968 3592 4002 3621
rect 3968 3524 4002 3546
rect 3968 3456 4002 3471
rect 3968 3388 4002 3396
rect 3968 3320 4002 3321
rect 3968 3280 4002 3286
rect 3968 3204 4002 3218
rect 3968 3128 4002 3150
rect 3968 3052 4002 3082
rect 3968 2980 4002 3014
rect 3968 2930 4002 2946
rect 1188 2910 1222 2926
rect 621 2794 637 2828
rect 671 2794 705 2828
rect 743 2794 755 2828
rect 811 2794 827 2828
rect 861 2794 881 2828
rect 936 2794 970 2828
rect 1011 2794 1052 2828
rect 1092 2794 1127 2828
rect 1161 2794 1177 2828
rect 1343 2794 1359 2828
rect 1402 2794 1454 2828
rect 1489 2794 1542 2828
rect 1583 2794 1599 2828
rect 1655 2794 1671 2828
rect 1721 2794 1766 2828
rect 1803 2794 1850 2828
rect 1895 2794 1911 2828
rect 2077 2794 2092 2828
rect 2127 2794 2181 2828
rect 2222 2794 2270 2828
rect 2317 2794 2333 2828
rect 2389 2794 2405 2828
rect 2446 2794 2499 2828
rect 2534 2794 2586 2828
rect 2629 2794 2645 2828
rect 2777 2794 2791 2828
rect 2827 2794 2861 2828
rect 2897 2794 2911 2828
rect 2967 2794 2979 2828
rect 3017 2794 3051 2828
rect 3085 2794 3101 2828
rect 3233 2794 3249 2828
rect 3283 2794 3289 2828
rect 3357 2794 3362 2828
rect 3396 2794 3397 2828
rect 3431 2794 3435 2828
rect 3469 2794 3470 2828
rect 3504 2794 3508 2828
rect 3542 2794 3543 2828
rect 3577 2794 3581 2828
rect 3615 2794 3616 2828
rect 3650 2794 3654 2828
rect 3688 2794 3689 2828
rect 3723 2794 3727 2828
rect 3761 2794 3762 2828
rect 3796 2794 3800 2828
rect 3834 2794 3835 2828
rect 3869 2794 3873 2828
rect 3907 2794 3908 2828
rect 3942 2794 3958 2828
rect 893 2475 905 2509
rect 951 2475 986 2509
rect 1023 2475 1055 2509
rect 1107 2475 1124 2509
rect 1191 2475 1192 2509
rect 1226 2475 1241 2509
rect 1294 2475 1325 2509
rect 1362 2475 1396 2509
rect 1442 2475 1454 2509
rect 1748 2434 1764 2468
rect 1798 2434 1832 2468
rect 1894 2434 1900 2468
rect 1934 2434 1944 2468
rect 2002 2434 2028 2468
rect 2070 2434 2104 2468
rect 2145 2434 2172 2468
rect 2228 2434 2240 2468
rect 2274 2434 2277 2468
rect 2802 2434 2818 2468
rect 2852 2434 2886 2468
rect 2920 2434 2954 2468
rect 2988 2434 3022 2468
rect 3064 2434 3090 2468
rect 3140 2434 3158 2468
rect 3216 2434 3226 2468
rect 3292 2434 3294 2468
rect 3328 2434 3334 2468
rect 3396 2434 3410 2468
rect 3464 2434 3486 2468
rect 3532 2434 3562 2468
rect 3600 2434 3634 2468
rect 3672 2434 3702 2468
rect 3748 2434 3752 2468
rect 3830 2457 3864 2469
rect 1642 2397 1676 2411
rect 2666 2407 2700 2423
rect 2384 2354 2400 2388
rect 2434 2373 2468 2388
rect 2502 2373 2518 2388
rect 2462 2354 2468 2373
rect 1642 2325 1676 2341
rect 2462 2339 2500 2354
rect 2666 2338 2700 2358
rect 1748 2278 1764 2312
rect 1798 2278 1832 2312
rect 1894 2278 1900 2312
rect 1934 2278 1944 2312
rect 2002 2278 2028 2312
rect 2070 2278 2104 2312
rect 2145 2278 2172 2312
rect 2228 2278 2240 2312
rect 2274 2278 2277 2312
rect 3830 2382 3864 2411
rect 1642 2252 1676 2271
rect 2666 2269 2700 2280
rect 2852 2278 2878 2312
rect 2920 2278 2954 2312
rect 2988 2278 3022 2312
rect 3064 2278 3090 2312
rect 3140 2278 3158 2312
rect 3216 2278 3226 2312
rect 3292 2278 3294 2312
rect 3328 2278 3334 2312
rect 3396 2278 3410 2312
rect 3464 2278 3486 2312
rect 3532 2278 3562 2312
rect 3600 2278 3634 2312
rect 3668 2278 3702 2312
rect 3736 2278 3752 2312
rect 3830 2306 3864 2342
rect 1171 2183 1187 2217
rect 1221 2183 1255 2217
rect 1317 2183 1323 2217
rect 1390 2183 1391 2217
rect 1425 2183 1429 2217
rect 1523 2206 1557 2218
rect 1523 2122 1557 2168
rect 1523 2072 1557 2084
rect 1642 2179 1676 2200
rect 2384 2198 2396 2232
rect 2434 2198 2468 2232
rect 2502 2198 2518 2232
rect 2666 2200 2700 2201
rect 2666 2156 2700 2166
rect 3830 2236 3864 2272
rect 3830 2166 3864 2196
rect 1642 2106 1676 2129
rect 1748 2122 1752 2156
rect 1798 2122 1832 2156
rect 1870 2122 1900 2156
rect 1954 2122 1968 2156
rect 2002 2122 2003 2156
rect 2070 2122 2086 2156
rect 2138 2122 2169 2156
rect 2206 2122 2240 2156
rect 2274 2122 2290 2156
rect 2802 2122 2818 2156
rect 2852 2122 2886 2156
rect 2920 2122 2954 2156
rect 2988 2122 3022 2156
rect 3064 2122 3090 2156
rect 3140 2122 3158 2156
rect 3216 2122 3226 2156
rect 3292 2122 3294 2156
rect 3328 2122 3334 2156
rect 3396 2122 3410 2156
rect 3464 2122 3486 2156
rect 3532 2122 3562 2156
rect 3600 2122 3634 2156
rect 3672 2122 3702 2156
rect 3748 2122 3752 2156
rect 3830 2108 3864 2120
rect 2666 2077 2700 2097
rect 1171 2027 1175 2061
rect 1221 2027 1255 2061
rect 1294 2027 1323 2061
rect 1379 2027 1391 2061
rect 1425 2027 1429 2061
rect 1642 2033 1676 2058
rect 2384 2042 2396 2076
rect 2434 2042 2468 2076
rect 2502 2042 2518 2076
rect 2666 2011 2700 2027
rect 1642 1950 1676 1987
rect 1748 1966 1764 2000
rect 1798 1966 1832 2000
rect 1894 1966 1900 2000
rect 1934 1966 1944 2000
rect 2002 1966 2028 2000
rect 2070 1966 2104 2000
rect 2145 1966 2172 2000
rect 2228 1966 2240 2000
rect 2274 1966 2277 2000
rect 2852 1966 2878 2000
rect 2920 1966 2954 2000
rect 2988 1966 3022 2000
rect 3064 1966 3090 2000
rect 3140 1966 3158 2000
rect 3216 1966 3226 2000
rect 3292 1966 3294 2000
rect 3328 1966 3334 2000
rect 3396 1966 3410 2000
rect 3464 1966 3486 2000
rect 3532 1966 3562 2000
rect 3600 1966 3634 2000
rect 3668 1966 3702 2000
rect 3736 1966 3752 2000
rect 1642 1879 1676 1916
rect 2384 1891 2396 1925
rect 2434 1891 2468 1925
rect 2502 1891 2518 1925
rect 1642 1821 1676 1845
rect 1748 1810 1764 1844
rect 1798 1810 1832 1844
rect 1894 1810 1900 1844
rect 1934 1810 1944 1844
rect 2002 1810 2028 1844
rect 2070 1810 2104 1844
rect 2145 1810 2172 1844
rect 2228 1810 2240 1844
rect 2274 1810 2277 1844
rect 591 1249 607 1283
rect 641 1249 675 1283
rect 713 1249 725 1283
rect 781 1249 797 1283
rect 842 1249 867 1283
rect 923 1249 936 1283
rect 970 1249 971 1283
rect 1039 1249 1053 1283
rect 1108 1249 1135 1283
rect 1177 1249 1193 1283
rect 1249 1249 1265 1283
rect 1310 1249 1337 1283
rect 1384 1249 1409 1283
rect 1458 1249 1481 1283
rect 1532 1249 1553 1283
rect 1606 1249 1625 1283
rect 1680 1249 1696 1283
rect 1755 1249 1767 1283
rect 1801 1249 1817 1283
rect 1983 1249 1999 1283
rect 2048 1249 2071 1283
rect 2127 1249 2143 1283
rect 2206 1249 2215 1283
rect 2249 1249 2251 1283
rect 2285 1249 2287 1283
rect 2321 1249 2330 1283
rect 2393 1249 2410 1283
rect 2464 1249 2490 1283
rect 2535 1249 2551 1283
rect 2607 1249 2623 1283
rect 2671 1249 2693 1283
rect 2749 1249 2762 1283
rect 2827 1249 2831 1283
rect 2865 1249 2872 1283
rect 2934 1249 2951 1283
rect 3003 1249 3019 1283
rect 580 1131 614 1147
rect 580 1077 614 1097
rect 580 1001 614 1029
rect 580 927 614 961
rect 580 859 614 890
rect 580 791 614 813
rect 580 723 614 736
rect 580 655 614 659
rect 580 616 614 621
rect 580 539 614 553
rect 580 462 614 485
rect 580 385 614 417
rect 580 315 614 349
rect 580 247 614 274
rect 736 1131 770 1147
rect 736 1077 770 1097
rect 736 1002 770 1029
rect 736 927 770 961
rect 736 859 770 893
rect 736 791 770 818
rect 736 723 770 743
rect 736 655 770 668
rect 736 587 770 592
rect 736 550 770 553
rect 736 474 770 485
rect 736 398 770 417
rect 736 322 770 349
rect 736 247 770 281
rect 736 197 770 213
rect 892 1131 926 1134
rect 892 1095 926 1097
rect 892 1021 926 1029
rect 892 947 926 961
rect 892 873 926 893
rect 892 799 926 825
rect 892 725 926 757
rect 892 655 926 689
rect 892 587 926 617
rect 892 519 926 543
rect 892 451 926 469
rect 892 383 926 395
rect 892 315 926 349
rect 892 247 926 281
rect 892 197 926 213
rect 1048 1131 1082 1147
rect 1048 1077 1082 1097
rect 1048 1002 1082 1029
rect 1048 927 1082 961
rect 1048 859 1082 893
rect 1048 791 1082 818
rect 1048 723 1082 743
rect 1048 655 1082 668
rect 1048 587 1082 592
rect 1048 550 1082 553
rect 1048 474 1082 485
rect 1048 398 1082 417
rect 1048 322 1082 349
rect 1048 247 1082 281
rect 1048 197 1082 213
rect 1204 1131 1238 1134
rect 1204 1092 1238 1097
rect 1204 1016 1238 1029
rect 1204 940 1238 961
rect 1204 864 1238 893
rect 1204 791 1238 825
rect 1204 723 1238 754
rect 1204 655 1238 677
rect 1204 587 1238 600
rect 1204 519 1238 523
rect 1204 480 1238 485
rect 1204 403 1238 417
rect 1204 326 1238 349
rect 1204 247 1238 281
rect 1204 197 1238 213
rect 1360 1131 1394 1147
rect 1360 1077 1394 1097
rect 1360 1001 1394 1029
rect 1360 927 1394 961
rect 1360 859 1394 890
rect 1360 791 1394 813
rect 1360 723 1394 736
rect 1360 655 1394 659
rect 1360 616 1394 621
rect 1360 539 1394 553
rect 1360 462 1394 485
rect 1360 385 1394 417
rect 1360 315 1394 349
rect 1360 247 1394 274
rect 1516 1131 1550 1134
rect 1516 1092 1550 1097
rect 1516 1016 1550 1029
rect 1516 940 1550 961
rect 1516 864 1550 893
rect 1516 791 1550 825
rect 1516 723 1550 754
rect 1516 655 1550 677
rect 1516 587 1550 600
rect 1516 519 1550 523
rect 1516 480 1550 485
rect 1516 403 1550 417
rect 1516 326 1550 349
rect 1516 247 1550 281
rect 1516 197 1550 213
rect 1672 1131 1706 1147
rect 1672 1077 1706 1097
rect 1672 1001 1706 1029
rect 1672 927 1706 961
rect 1672 859 1706 890
rect 1672 791 1706 813
rect 1672 723 1706 736
rect 1672 655 1706 659
rect 1672 616 1706 621
rect 1672 539 1706 553
rect 1672 462 1706 485
rect 1672 385 1706 417
rect 1672 315 1706 349
rect 1672 247 1706 274
rect 1828 1131 1862 1134
rect 1828 1092 1862 1097
rect 1828 1016 1862 1029
rect 1828 940 1862 961
rect 1828 864 1862 893
rect 1828 791 1862 825
rect 1828 723 1862 754
rect 1828 655 1862 677
rect 1828 587 1862 600
rect 1828 519 1862 523
rect 1828 480 1862 485
rect 1828 403 1862 417
rect 1828 326 1862 349
rect 1828 247 1862 281
rect 1828 197 1862 213
rect 1938 1131 1972 1134
rect 1938 1092 1972 1097
rect 1938 1016 1972 1029
rect 1938 940 1972 961
rect 1938 864 1972 893
rect 1938 791 1972 825
rect 1938 723 1972 754
rect 1938 655 1972 677
rect 1938 587 1972 600
rect 1938 519 1972 523
rect 1938 480 1972 485
rect 1938 403 1972 417
rect 1938 326 1972 349
rect 1938 247 1972 281
rect 1938 197 1972 213
rect 2094 1131 2128 1147
rect 2094 1077 2128 1097
rect 2094 1001 2128 1029
rect 2094 927 2128 961
rect 2094 859 2128 890
rect 2094 791 2128 813
rect 2094 723 2128 736
rect 2094 655 2128 659
rect 2094 616 2128 621
rect 2094 539 2128 553
rect 2094 462 2128 485
rect 2094 385 2128 417
rect 2094 315 2128 349
rect 2094 247 2128 274
rect 2250 1131 2284 1134
rect 2250 1092 2284 1097
rect 2250 1016 2284 1029
rect 2250 940 2284 961
rect 2250 864 2284 893
rect 2250 791 2284 825
rect 2250 723 2284 754
rect 2250 655 2284 677
rect 2250 587 2284 600
rect 2250 519 2284 523
rect 2250 480 2284 485
rect 2250 403 2284 417
rect 2250 326 2284 349
rect 2250 247 2284 281
rect 2250 197 2284 213
rect 2406 1131 2440 1147
rect 2406 1077 2440 1097
rect 2406 1001 2440 1029
rect 2406 927 2440 961
rect 2406 859 2440 890
rect 2406 791 2440 813
rect 2406 723 2440 736
rect 2406 655 2440 659
rect 2406 616 2440 621
rect 2406 539 2440 553
rect 2406 462 2440 485
rect 2406 385 2440 417
rect 2406 315 2440 349
rect 2406 247 2440 274
rect 2562 1131 2596 1134
rect 2562 1092 2596 1097
rect 2562 1016 2596 1029
rect 2562 940 2596 961
rect 2562 864 2596 893
rect 2562 791 2596 825
rect 2562 723 2596 754
rect 2562 655 2596 677
rect 2562 587 2596 600
rect 2562 519 2596 523
rect 2562 480 2596 485
rect 2562 403 2596 417
rect 2562 326 2596 349
rect 2562 247 2596 281
rect 2562 197 2596 213
rect 2718 1131 2752 1147
rect 2718 1077 2752 1097
rect 2718 1002 2752 1029
rect 2718 927 2752 961
rect 2718 859 2752 893
rect 2718 791 2752 818
rect 2718 723 2752 743
rect 2718 655 2752 668
rect 2718 587 2752 593
rect 2718 552 2752 553
rect 2718 477 2752 485
rect 2718 402 2752 417
rect 2718 326 2752 349
rect 2718 247 2752 281
rect 2718 197 2752 213
rect 2874 1131 2908 1134
rect 2874 1095 2908 1097
rect 2874 1022 2908 1029
rect 2874 949 2908 961
rect 2874 876 2908 893
rect 2874 803 2908 825
rect 2874 730 2908 757
rect 2874 657 2908 689
rect 2874 587 2908 621
rect 2874 519 2908 549
rect 2874 451 2908 475
rect 2874 383 2908 401
rect 2874 315 2908 349
rect 2874 247 2908 281
rect 2874 197 2908 213
rect 3030 1131 3064 1147
rect 3030 1077 3064 1097
rect 3030 1002 3064 1029
rect 3030 927 3064 961
rect 3030 859 3064 893
rect 3030 791 3064 818
rect 3030 723 3064 743
rect 3030 655 3064 668
rect 3030 587 3064 593
rect 3030 552 3064 553
rect 3030 477 3064 485
rect 3030 402 3064 417
rect 3030 326 3064 349
rect 3030 247 3064 281
rect 3030 197 3064 213
rect 594 91 616 125
rect 652 91 687 125
rect 723 91 756 125
rect 796 91 825 125
rect 869 91 894 125
rect 942 91 963 125
rect 1015 91 1032 125
rect 1088 91 1101 125
rect 1162 91 1170 125
rect 1236 91 1239 125
rect 1273 91 1276 125
rect 1342 91 1350 125
rect 1411 91 1424 125
rect 1480 91 1498 125
rect 1549 91 1572 125
rect 1618 91 1646 125
rect 1687 91 1720 125
rect 1756 91 1791 125
rect 1828 91 1861 125
rect 1902 91 1931 125
rect 1976 91 2001 125
rect 2050 91 2071 125
rect 2124 91 2141 125
rect 2198 91 2211 125
rect 2272 91 2281 125
rect 2346 91 2351 125
rect 2385 91 2386 125
rect 2420 91 2421 125
rect 2455 91 2460 125
rect 2525 91 2534 125
rect 2595 91 2608 125
rect 2665 91 2682 125
rect 2735 91 2756 125
rect 2805 91 2830 125
rect 2875 91 2904 125
rect 2945 91 2978 125
rect 3015 91 3039 125
<< viali >>
rect 603 3950 637 3984
rect 677 3950 705 3984
rect 705 3950 711 3984
rect 751 3950 773 3984
rect 773 3950 785 3984
rect 825 3950 841 3984
rect 841 3950 859 3984
rect 899 3950 909 3984
rect 909 3950 933 3984
rect 973 3950 977 3984
rect 977 3950 1007 3984
rect 1047 3950 1079 3984
rect 1079 3950 1081 3984
rect 1121 3950 1147 3984
rect 1147 3950 1155 3984
rect 1195 3950 1215 3984
rect 1215 3950 1229 3984
rect 1269 3950 1283 3984
rect 1283 3950 1303 3984
rect 1343 3950 1351 3984
rect 1351 3950 1377 3984
rect 1417 3950 1419 3984
rect 1419 3950 1451 3984
rect 1491 3950 1521 3984
rect 1521 3950 1525 3984
rect 1565 3950 1589 3984
rect 1589 3950 1599 3984
rect 1639 3950 1657 3984
rect 1657 3950 1673 3984
rect 1712 3950 1725 3984
rect 1725 3950 1746 3984
rect 1785 3950 1793 3984
rect 1793 3950 1819 3984
rect 1858 3950 1861 3984
rect 1861 3950 1892 3984
rect 1931 3950 1963 3984
rect 1963 3950 1965 3984
rect 2004 3950 2031 3984
rect 2031 3950 2038 3984
rect 2077 3950 2099 3984
rect 2099 3950 2111 3984
rect 2150 3950 2167 3984
rect 2167 3950 2184 3984
rect 2223 3950 2235 3984
rect 2235 3950 2257 3984
rect 2296 3950 2303 3984
rect 2303 3950 2330 3984
rect 2369 3950 2371 3984
rect 2371 3950 2403 3984
rect 2442 3950 2473 3984
rect 2473 3950 2476 3984
rect 2515 3950 2541 3984
rect 2541 3950 2549 3984
rect 2588 3950 2609 3984
rect 2609 3950 2622 3984
rect 2661 3950 2677 3984
rect 2677 3950 2695 3984
rect 2734 3950 2745 3984
rect 2745 3950 2768 3984
rect 2807 3950 2813 3984
rect 2813 3950 2841 3984
rect 2880 3950 2881 3984
rect 2881 3950 2914 3984
rect 2953 3950 2983 3984
rect 2983 3950 2987 3984
rect 3026 3950 3051 3984
rect 3051 3950 3060 3984
rect 3099 3950 3119 3984
rect 3119 3950 3133 3984
rect 3172 3950 3187 3984
rect 3187 3950 3206 3984
rect 3245 3950 3255 3984
rect 3255 3950 3279 3984
rect 3318 3950 3323 3984
rect 3323 3950 3352 3984
rect 3391 3950 3425 3984
rect 3464 3950 3493 3984
rect 3493 3950 3498 3984
rect 3537 3950 3561 3984
rect 3561 3950 3571 3984
rect 3610 3950 3629 3984
rect 3629 3950 3644 3984
rect 3683 3950 3697 3984
rect 3697 3950 3717 3984
rect 3756 3950 3765 3984
rect 3765 3950 3790 3984
rect 3829 3950 3833 3984
rect 3833 3950 3863 3984
rect 3902 3950 3935 3984
rect 3935 3950 3936 3984
rect 3975 3950 4009 3984
rect 1298 3694 1332 3711
rect 1298 3677 1332 3694
rect 1298 3626 1332 3637
rect 1298 3603 1332 3626
rect 1298 3558 1332 3563
rect 1298 3529 1332 3558
rect 1298 3456 1332 3489
rect 1298 3455 1332 3456
rect 1298 3388 1332 3414
rect 1298 3380 1332 3388
rect 1298 3320 1332 3339
rect 1298 3305 1332 3320
rect 1298 3252 1332 3264
rect 1298 3230 1332 3252
rect 610 3166 644 3200
rect 610 3062 644 3070
rect 610 3036 644 3062
rect 766 3166 800 3200
rect 766 3096 800 3120
rect 766 3086 800 3096
rect 766 3028 800 3040
rect 766 3006 800 3028
rect 922 3166 956 3200
rect 922 3096 956 3123
rect 922 3089 956 3096
rect 922 3028 956 3045
rect 922 3011 956 3028
rect 1032 3166 1066 3200
rect 1298 3184 1332 3189
rect 1032 3096 1066 3112
rect 1032 3078 1066 3096
rect 1032 2994 1066 3023
rect 1032 2989 1066 2994
rect 1188 3130 1222 3164
rect 1188 3062 1222 3065
rect 1188 3031 1222 3062
rect 1298 3155 1332 3184
rect 1298 3082 1332 3114
rect 1298 3080 1332 3082
rect 1298 3014 1332 3039
rect 1298 3005 1332 3014
rect 1298 2946 1332 2964
rect 1298 2930 1332 2946
rect 1454 3694 1488 3711
rect 1454 3677 1488 3694
rect 1454 3626 1488 3637
rect 1454 3603 1488 3626
rect 1454 3558 1488 3563
rect 1454 3529 1488 3558
rect 1454 3456 1488 3489
rect 1454 3455 1488 3456
rect 1454 3388 1488 3415
rect 1454 3381 1488 3388
rect 1454 3320 1488 3340
rect 1454 3306 1488 3320
rect 1454 3252 1488 3265
rect 1454 3231 1488 3252
rect 1454 3184 1488 3190
rect 1454 3156 1488 3184
rect 1454 3082 1488 3115
rect 1454 3081 1488 3082
rect 1454 3014 1488 3040
rect 1454 3006 1488 3014
rect 1610 3694 1644 3711
rect 1610 3677 1644 3694
rect 1610 3626 1644 3637
rect 1610 3603 1644 3626
rect 1610 3558 1644 3563
rect 1610 3529 1644 3558
rect 1610 3456 1644 3489
rect 1610 3455 1644 3456
rect 1610 3388 1644 3414
rect 1610 3380 1644 3388
rect 1610 3320 1644 3339
rect 1610 3305 1644 3320
rect 1610 3252 1644 3264
rect 1610 3230 1644 3252
rect 1610 3184 1644 3189
rect 1610 3155 1644 3184
rect 1610 3082 1644 3114
rect 1610 3080 1644 3082
rect 1610 3014 1644 3039
rect 1610 3005 1644 3014
rect 1610 2946 1644 2964
rect 1610 2930 1644 2946
rect 1766 3864 1800 3880
rect 1766 3846 1800 3864
rect 1766 3796 1800 3804
rect 1766 3770 1800 3796
rect 1766 3694 1800 3728
rect 1766 3626 1800 3652
rect 1766 3618 1800 3626
rect 1766 3558 1800 3576
rect 1766 3542 1800 3558
rect 1766 3490 1800 3500
rect 1766 3466 1800 3490
rect 1766 3422 1800 3424
rect 1766 3390 1800 3422
rect 1766 3320 1800 3348
rect 1766 3314 1800 3320
rect 1766 3252 1800 3271
rect 1766 3237 1800 3252
rect 1766 3184 1800 3194
rect 1766 3160 1800 3184
rect 1766 3116 1800 3117
rect 1766 3083 1800 3116
rect 1766 3014 1800 3040
rect 1766 3006 1800 3014
rect 1922 3694 1956 3711
rect 1922 3677 1956 3694
rect 1922 3626 1956 3637
rect 1922 3603 1956 3626
rect 1922 3558 1956 3563
rect 1922 3529 1956 3558
rect 1922 3456 1956 3489
rect 1922 3455 1956 3456
rect 1922 3388 1956 3414
rect 1922 3380 1956 3388
rect 1922 3320 1956 3339
rect 1922 3305 1956 3320
rect 1922 3252 1956 3264
rect 1922 3230 1956 3252
rect 1922 3184 1956 3189
rect 1922 3155 1956 3184
rect 1922 3082 1956 3114
rect 1922 3080 1956 3082
rect 1922 3014 1956 3039
rect 1922 3005 1956 3014
rect 1922 2946 1956 2964
rect 1922 2930 1956 2946
rect 2032 3694 2066 3711
rect 2032 3677 2066 3694
rect 2032 3626 2066 3637
rect 2032 3603 2066 3626
rect 2032 3558 2066 3563
rect 2032 3529 2066 3558
rect 2032 3456 2066 3489
rect 2032 3455 2066 3456
rect 2032 3388 2066 3414
rect 2032 3380 2066 3388
rect 2032 3320 2066 3339
rect 2032 3305 2066 3320
rect 2032 3252 2066 3264
rect 2032 3230 2066 3252
rect 2032 3184 2066 3189
rect 2032 3155 2066 3184
rect 2032 3082 2066 3114
rect 2032 3080 2066 3082
rect 2032 3014 2066 3039
rect 2032 3005 2066 3014
rect 2032 2946 2066 2964
rect 2032 2930 2066 2946
rect 2188 3864 2222 3880
rect 2188 3846 2222 3864
rect 2188 3796 2222 3804
rect 2188 3770 2222 3796
rect 2188 3694 2222 3728
rect 2188 3626 2222 3652
rect 2188 3618 2222 3626
rect 2188 3558 2222 3576
rect 2188 3542 2222 3558
rect 2188 3490 2222 3500
rect 2188 3466 2222 3490
rect 2188 3422 2222 3424
rect 2188 3390 2222 3422
rect 2188 3320 2222 3348
rect 2188 3314 2222 3320
rect 2188 3252 2222 3271
rect 2188 3237 2222 3252
rect 2188 3184 2222 3194
rect 2188 3160 2222 3184
rect 2188 3116 2222 3117
rect 2188 3083 2222 3116
rect 2188 3014 2222 3040
rect 2188 3006 2222 3014
rect 2344 3694 2378 3711
rect 2344 3677 2378 3694
rect 2344 3626 2378 3637
rect 2344 3603 2378 3626
rect 2344 3558 2378 3563
rect 2344 3529 2378 3558
rect 2344 3456 2378 3489
rect 2344 3455 2378 3456
rect 2344 3388 2378 3414
rect 2344 3380 2378 3388
rect 2344 3320 2378 3339
rect 2344 3305 2378 3320
rect 2344 3252 2378 3264
rect 2344 3230 2378 3252
rect 2344 3184 2378 3189
rect 2344 3155 2378 3184
rect 2344 3082 2378 3114
rect 2344 3080 2378 3082
rect 2344 3014 2378 3039
rect 2344 3005 2378 3014
rect 2344 2946 2378 2964
rect 2344 2930 2378 2946
rect 2500 3694 2534 3711
rect 2500 3677 2534 3694
rect 2500 3626 2534 3637
rect 2500 3603 2534 3626
rect 2500 3558 2534 3563
rect 2500 3529 2534 3558
rect 2500 3456 2534 3489
rect 2500 3455 2534 3456
rect 2500 3388 2534 3415
rect 2500 3381 2534 3388
rect 2500 3320 2534 3340
rect 2500 3306 2534 3320
rect 2500 3252 2534 3265
rect 2500 3231 2534 3252
rect 2500 3184 2534 3190
rect 2500 3156 2534 3184
rect 2500 3082 2534 3115
rect 2500 3081 2534 3082
rect 2500 3014 2534 3040
rect 2500 3006 2534 3014
rect 2656 3694 2690 3711
rect 2656 3677 2690 3694
rect 2656 3626 2690 3637
rect 2656 3603 2690 3626
rect 2656 3558 2690 3563
rect 2656 3529 2690 3558
rect 2656 3456 2690 3489
rect 2656 3455 2690 3456
rect 2656 3388 2690 3414
rect 2656 3380 2690 3388
rect 2656 3320 2690 3339
rect 2656 3305 2690 3320
rect 2656 3252 2690 3264
rect 2656 3230 2690 3252
rect 2656 3184 2690 3189
rect 2656 3155 2690 3184
rect 2656 3082 2690 3114
rect 2656 3080 2690 3082
rect 2656 3014 2690 3039
rect 2656 3005 2690 3014
rect 2656 2946 2690 2964
rect 2656 2930 2690 2946
rect 2766 3694 2800 3711
rect 2766 3677 2800 3694
rect 2766 3626 2800 3637
rect 2766 3603 2800 3626
rect 2766 3558 2800 3563
rect 2766 3529 2800 3558
rect 2766 3456 2800 3489
rect 2766 3455 2800 3456
rect 2766 3388 2800 3415
rect 2766 3381 2800 3388
rect 2766 3320 2800 3340
rect 2766 3306 2800 3320
rect 2766 3252 2800 3265
rect 2766 3231 2800 3252
rect 2766 3184 2800 3190
rect 2766 3156 2800 3184
rect 2766 3082 2800 3115
rect 2766 3081 2800 3082
rect 2766 3014 2800 3040
rect 2766 3006 2800 3014
rect 2922 3694 2956 3711
rect 2922 3677 2956 3694
rect 2922 3626 2956 3637
rect 2922 3603 2956 3626
rect 2922 3558 2956 3563
rect 2922 3529 2956 3558
rect 2922 3456 2956 3489
rect 2922 3455 2956 3456
rect 2922 3388 2956 3415
rect 2922 3381 2956 3388
rect 2922 3320 2956 3340
rect 2922 3306 2956 3320
rect 2922 3252 2956 3265
rect 2922 3231 2956 3252
rect 2922 3184 2956 3190
rect 2922 3156 2956 3184
rect 2922 3082 2956 3115
rect 2922 3081 2956 3082
rect 2922 3014 2956 3040
rect 2922 3006 2956 3014
rect 3078 3864 3112 3880
rect 3078 3846 3112 3864
rect 3078 3796 3112 3803
rect 3078 3769 3112 3796
rect 3078 3694 3112 3725
rect 3078 3691 3112 3694
rect 3078 3626 3112 3647
rect 3078 3613 3112 3626
rect 3078 3558 3112 3569
rect 3078 3535 3112 3558
rect 3078 3490 3112 3491
rect 3078 3457 3112 3490
rect 3078 3388 3112 3413
rect 3078 3379 3112 3388
rect 3078 3320 3112 3335
rect 3078 3301 3112 3320
rect 3078 3252 3112 3257
rect 3078 3223 3112 3252
rect 3078 3150 3112 3179
rect 3078 3145 3112 3150
rect 3078 3082 3112 3101
rect 3078 3067 3112 3082
rect 3078 3014 3112 3023
rect 3078 2989 3112 3014
rect 3188 3694 3222 3711
rect 3188 3677 3222 3694
rect 3188 3626 3222 3637
rect 3188 3603 3222 3626
rect 3188 3558 3222 3563
rect 3188 3529 3222 3558
rect 3188 3456 3222 3488
rect 3188 3454 3222 3456
rect 3188 3388 3222 3413
rect 3188 3379 3222 3388
rect 3188 3320 3222 3338
rect 3188 3304 3222 3320
rect 3188 3252 3222 3263
rect 3188 3229 3222 3252
rect 3188 3184 3222 3188
rect 3188 3154 3222 3184
rect 3188 3082 3222 3113
rect 3188 3079 3222 3082
rect 3188 3014 3222 3038
rect 3188 3004 3222 3014
rect 3188 2946 3222 2963
rect 3188 2929 3222 2946
rect 3344 3864 3378 3880
rect 3344 3846 3378 3864
rect 3344 3796 3378 3805
rect 3344 3771 3378 3796
rect 3344 3728 3378 3730
rect 3344 3696 3378 3728
rect 3344 3626 3378 3655
rect 3344 3621 3378 3626
rect 3344 3558 3378 3580
rect 3344 3546 3378 3558
rect 3344 3490 3378 3505
rect 3344 3471 3378 3490
rect 3344 3422 3378 3430
rect 3344 3396 3378 3422
rect 3344 3354 3378 3355
rect 3344 3321 3378 3354
rect 3344 3252 3378 3280
rect 3344 3246 3378 3252
rect 3344 3184 3378 3204
rect 3344 3170 3378 3184
rect 3344 3116 3378 3128
rect 3344 3094 3378 3116
rect 3344 3048 3378 3052
rect 3344 3018 3378 3048
rect 3500 3694 3534 3711
rect 3500 3677 3534 3694
rect 3500 3626 3534 3637
rect 3500 3603 3534 3626
rect 3500 3558 3534 3563
rect 3500 3529 3534 3558
rect 3500 3456 3534 3488
rect 3500 3454 3534 3456
rect 3500 3388 3534 3413
rect 3500 3379 3534 3388
rect 3500 3320 3534 3338
rect 3500 3304 3534 3320
rect 3500 3252 3534 3263
rect 3500 3229 3534 3252
rect 3500 3184 3534 3188
rect 3500 3154 3534 3184
rect 3500 3082 3534 3113
rect 3500 3079 3534 3082
rect 3500 3014 3534 3038
rect 3500 3004 3534 3014
rect 3500 2946 3534 2963
rect 3500 2929 3534 2946
rect 3656 3864 3690 3880
rect 3656 3846 3690 3864
rect 3656 3796 3690 3805
rect 3656 3771 3690 3796
rect 3656 3728 3690 3730
rect 3656 3696 3690 3728
rect 3656 3626 3690 3655
rect 3656 3621 3690 3626
rect 3656 3558 3690 3580
rect 3656 3546 3690 3558
rect 3656 3490 3690 3505
rect 3656 3471 3690 3490
rect 3656 3422 3690 3430
rect 3656 3396 3690 3422
rect 3656 3354 3690 3355
rect 3656 3321 3690 3354
rect 3656 3252 3690 3280
rect 3656 3246 3690 3252
rect 3656 3184 3690 3204
rect 3656 3170 3690 3184
rect 3656 3116 3690 3128
rect 3656 3094 3690 3116
rect 3656 3048 3690 3052
rect 3656 3018 3690 3048
rect 3812 3694 3846 3711
rect 3812 3677 3846 3694
rect 3812 3626 3846 3637
rect 3812 3603 3846 3626
rect 3812 3558 3846 3563
rect 3812 3529 3846 3558
rect 3812 3456 3846 3488
rect 3812 3454 3846 3456
rect 3812 3388 3846 3413
rect 3812 3379 3846 3388
rect 3812 3320 3846 3338
rect 3812 3304 3846 3320
rect 3812 3252 3846 3263
rect 3812 3229 3846 3252
rect 3812 3184 3846 3188
rect 3812 3154 3846 3184
rect 3812 3082 3846 3113
rect 3812 3079 3846 3082
rect 3812 3014 3846 3038
rect 3812 3004 3846 3014
rect 3812 2946 3846 2963
rect 3812 2929 3846 2946
rect 3968 3864 4002 3880
rect 3968 3846 4002 3864
rect 3968 3796 4002 3805
rect 3968 3771 4002 3796
rect 3968 3728 4002 3730
rect 3968 3696 4002 3728
rect 3968 3626 4002 3655
rect 3968 3621 4002 3626
rect 3968 3558 4002 3580
rect 3968 3546 4002 3558
rect 3968 3490 4002 3505
rect 3968 3471 4002 3490
rect 3968 3422 4002 3430
rect 3968 3396 4002 3422
rect 3968 3354 4002 3355
rect 3968 3321 4002 3354
rect 3968 3252 4002 3280
rect 3968 3246 4002 3252
rect 3968 3184 4002 3204
rect 3968 3170 4002 3184
rect 3968 3116 4002 3128
rect 3968 3094 4002 3116
rect 3968 3048 4002 3052
rect 3968 3018 4002 3048
rect 637 2794 671 2828
rect 709 2794 739 2828
rect 739 2794 743 2828
rect 881 2794 902 2828
rect 902 2794 915 2828
rect 970 2794 977 2828
rect 977 2794 1004 2828
rect 1058 2794 1086 2828
rect 1086 2794 1092 2828
rect 1368 2794 1393 2828
rect 1393 2794 1402 2828
rect 1455 2794 1488 2828
rect 1488 2794 1489 2828
rect 1542 2794 1549 2828
rect 1549 2794 1576 2828
rect 1687 2794 1705 2828
rect 1705 2794 1721 2828
rect 1769 2794 1800 2828
rect 1800 2794 1803 2828
rect 1850 2794 1861 2828
rect 1861 2794 1884 2828
rect 2092 2794 2093 2828
rect 2093 2794 2126 2828
rect 2181 2794 2188 2828
rect 2188 2794 2215 2828
rect 2270 2794 2283 2828
rect 2283 2794 2304 2828
rect 2412 2794 2439 2828
rect 2439 2794 2446 2828
rect 2499 2794 2500 2828
rect 2500 2794 2533 2828
rect 2586 2794 2595 2828
rect 2595 2794 2620 2828
rect 2791 2794 2793 2828
rect 2793 2794 2825 2828
rect 2863 2794 2895 2828
rect 2895 2794 2897 2828
rect 2979 2794 2983 2828
rect 2983 2794 3013 2828
rect 3051 2794 3085 2828
rect 3289 2794 3323 2828
rect 3362 2794 3396 2828
rect 3435 2794 3469 2828
rect 3508 2794 3542 2828
rect 3581 2794 3615 2828
rect 3654 2794 3688 2828
rect 3727 2794 3761 2828
rect 3800 2794 3834 2828
rect 3873 2794 3907 2828
rect 905 2475 917 2509
rect 917 2475 939 2509
rect 989 2475 1020 2509
rect 1020 2475 1023 2509
rect 1073 2475 1089 2509
rect 1089 2475 1107 2509
rect 1157 2475 1158 2509
rect 1158 2475 1191 2509
rect 1241 2475 1260 2509
rect 1260 2475 1275 2509
rect 1325 2475 1328 2509
rect 1328 2475 1359 2509
rect 1408 2475 1430 2509
rect 1430 2475 1442 2509
rect 1642 2445 1676 2469
rect 1642 2435 1676 2445
rect 1860 2434 1866 2468
rect 1866 2434 1894 2468
rect 1944 2434 1968 2468
rect 1968 2434 1978 2468
rect 2028 2434 2036 2468
rect 2036 2434 2062 2468
rect 2111 2434 2138 2468
rect 2138 2434 2145 2468
rect 2194 2434 2206 2468
rect 2206 2434 2228 2468
rect 2277 2434 2311 2468
rect 2954 2434 2988 2468
rect 3030 2434 3056 2468
rect 3056 2434 3064 2468
rect 3106 2434 3124 2468
rect 3124 2434 3140 2468
rect 3182 2434 3192 2468
rect 3192 2434 3216 2468
rect 3258 2434 3260 2468
rect 3260 2434 3292 2468
rect 3334 2434 3362 2468
rect 3362 2434 3368 2468
rect 3410 2434 3430 2468
rect 3430 2434 3444 2468
rect 3486 2434 3498 2468
rect 3498 2434 3520 2468
rect 3562 2434 3566 2468
rect 3566 2434 3596 2468
rect 3638 2434 3668 2468
rect 3668 2434 3672 2468
rect 3714 2434 3736 2468
rect 3736 2434 3748 2468
rect 3830 2445 3864 2457
rect 3830 2423 3864 2445
rect 1642 2375 1676 2397
rect 1642 2363 1676 2375
rect 2666 2373 2700 2392
rect 2428 2354 2434 2373
rect 2434 2354 2462 2373
rect 2500 2354 2502 2373
rect 2502 2354 2534 2373
rect 2428 2339 2462 2354
rect 2500 2339 2534 2354
rect 2666 2358 2700 2373
rect 1642 2305 1676 2325
rect 1642 2291 1676 2305
rect 1860 2278 1866 2312
rect 1866 2278 1894 2312
rect 1944 2278 1968 2312
rect 1968 2278 1978 2312
rect 2028 2278 2036 2312
rect 2036 2278 2062 2312
rect 2111 2278 2138 2312
rect 2138 2278 2145 2312
rect 2194 2278 2206 2312
rect 2206 2278 2228 2312
rect 2277 2278 2311 2312
rect 2666 2304 2700 2314
rect 3830 2376 3864 2382
rect 3830 2348 3864 2376
rect 2666 2280 2700 2304
rect 1642 2234 1676 2252
rect 1642 2218 1676 2234
rect 2802 2278 2818 2312
rect 2818 2278 2836 2312
rect 2878 2278 2886 2312
rect 2886 2278 2912 2312
rect 2954 2278 2988 2312
rect 3030 2278 3056 2312
rect 3056 2278 3064 2312
rect 3106 2278 3124 2312
rect 3124 2278 3140 2312
rect 3182 2278 3192 2312
rect 3192 2278 3216 2312
rect 3258 2278 3260 2312
rect 3260 2278 3292 2312
rect 3334 2278 3362 2312
rect 3362 2278 3368 2312
rect 3410 2278 3430 2312
rect 3430 2278 3444 2312
rect 3486 2278 3498 2312
rect 3498 2278 3520 2312
rect 3562 2278 3566 2312
rect 3566 2278 3596 2312
rect 1283 2183 1289 2217
rect 1289 2183 1317 2217
rect 1356 2183 1357 2217
rect 1357 2183 1390 2217
rect 1429 2183 1463 2217
rect 1523 2202 1557 2206
rect 1523 2172 1557 2202
rect 1523 2088 1557 2118
rect 1523 2084 1557 2088
rect 2396 2198 2400 2232
rect 2400 2198 2430 2232
rect 2468 2198 2502 2232
rect 2666 2201 2700 2235
rect 1642 2163 1676 2179
rect 1642 2145 1676 2163
rect 3830 2272 3864 2306
rect 3830 2202 3864 2230
rect 3830 2196 3864 2202
rect 1752 2122 1764 2156
rect 1764 2122 1786 2156
rect 1836 2122 1866 2156
rect 1866 2122 1870 2156
rect 1920 2122 1934 2156
rect 1934 2122 1954 2156
rect 2003 2122 2036 2156
rect 2036 2122 2037 2156
rect 2086 2122 2104 2156
rect 2104 2122 2120 2156
rect 2169 2122 2172 2156
rect 2172 2122 2203 2156
rect 2666 2131 2700 2156
rect 2666 2122 2700 2131
rect 2954 2122 2988 2156
rect 3030 2122 3056 2156
rect 3056 2122 3064 2156
rect 3106 2122 3124 2156
rect 3124 2122 3140 2156
rect 3182 2122 3192 2156
rect 3192 2122 3216 2156
rect 3258 2122 3260 2156
rect 3260 2122 3292 2156
rect 3334 2122 3362 2156
rect 3362 2122 3368 2156
rect 3410 2122 3430 2156
rect 3430 2122 3444 2156
rect 3486 2122 3498 2156
rect 3498 2122 3520 2156
rect 3562 2122 3566 2156
rect 3566 2122 3596 2156
rect 3638 2122 3668 2156
rect 3668 2122 3672 2156
rect 3714 2122 3736 2156
rect 3736 2122 3748 2156
rect 3830 2132 3864 2154
rect 1642 2092 1676 2106
rect 1642 2072 1676 2092
rect 3830 2120 3864 2132
rect 1175 2027 1187 2061
rect 1187 2027 1209 2061
rect 1260 2027 1289 2061
rect 1289 2027 1294 2061
rect 1345 2027 1357 2061
rect 1357 2027 1379 2061
rect 1429 2027 1463 2061
rect 2396 2042 2400 2076
rect 2400 2042 2430 2076
rect 2468 2042 2502 2076
rect 2666 2061 2700 2077
rect 2666 2043 2700 2061
rect 1642 2021 1676 2033
rect 1642 1999 1676 2021
rect 1860 1966 1866 2000
rect 1866 1966 1894 2000
rect 1944 1966 1968 2000
rect 1968 1966 1978 2000
rect 2028 1966 2036 2000
rect 2036 1966 2062 2000
rect 2111 1966 2138 2000
rect 2138 1966 2145 2000
rect 2194 1966 2206 2000
rect 2206 1966 2228 2000
rect 2277 1966 2311 2000
rect 2802 1966 2818 2000
rect 2818 1966 2836 2000
rect 2878 1966 2886 2000
rect 2886 1966 2912 2000
rect 2954 1966 2988 2000
rect 3030 1966 3056 2000
rect 3056 1966 3064 2000
rect 3106 1966 3124 2000
rect 3124 1966 3140 2000
rect 3182 1966 3192 2000
rect 3192 1966 3216 2000
rect 3258 1966 3260 2000
rect 3260 1966 3292 2000
rect 3334 1966 3362 2000
rect 3362 1966 3368 2000
rect 3410 1966 3430 2000
rect 3430 1966 3444 2000
rect 3486 1966 3498 2000
rect 3498 1966 3520 2000
rect 3562 1966 3566 2000
rect 3566 1966 3596 2000
rect 2396 1891 2400 1925
rect 2400 1891 2430 1925
rect 2468 1891 2502 1925
rect 1860 1810 1866 1844
rect 1866 1810 1894 1844
rect 1944 1810 1968 1844
rect 1968 1810 1978 1844
rect 2028 1810 2036 1844
rect 2036 1810 2062 1844
rect 2111 1810 2138 1844
rect 2138 1810 2145 1844
rect 2194 1810 2206 1844
rect 2206 1810 2228 1844
rect 2277 1810 2311 1844
rect 607 1249 641 1283
rect 679 1249 709 1283
rect 709 1249 713 1283
rect 808 1249 831 1283
rect 831 1249 842 1283
rect 889 1249 901 1283
rect 901 1249 923 1283
rect 971 1249 1005 1283
rect 1053 1249 1074 1283
rect 1074 1249 1087 1283
rect 1135 1249 1143 1283
rect 1143 1249 1169 1283
rect 1276 1249 1299 1283
rect 1299 1249 1310 1283
rect 1350 1249 1371 1283
rect 1371 1249 1384 1283
rect 1424 1249 1443 1283
rect 1443 1249 1458 1283
rect 1498 1249 1515 1283
rect 1515 1249 1532 1283
rect 1572 1249 1587 1283
rect 1587 1249 1606 1283
rect 1646 1249 1659 1283
rect 1659 1249 1680 1283
rect 1721 1249 1730 1283
rect 1730 1249 1755 1283
rect 2014 1249 2033 1283
rect 2033 1249 2048 1283
rect 2093 1249 2105 1283
rect 2105 1249 2127 1283
rect 2172 1249 2177 1283
rect 2177 1249 2206 1283
rect 2251 1249 2285 1283
rect 2330 1249 2359 1283
rect 2359 1249 2364 1283
rect 2410 1249 2430 1283
rect 2430 1249 2444 1283
rect 2490 1249 2501 1283
rect 2501 1249 2524 1283
rect 2637 1249 2657 1283
rect 2657 1249 2671 1283
rect 2715 1249 2727 1283
rect 2727 1249 2749 1283
rect 2793 1249 2796 1283
rect 2796 1249 2827 1283
rect 2872 1249 2900 1283
rect 2900 1249 2906 1283
rect 2951 1249 2969 1283
rect 2969 1249 2985 1283
rect 580 1063 614 1077
rect 580 1043 614 1063
rect 580 995 614 1001
rect 580 967 614 995
rect 580 893 614 924
rect 580 890 614 893
rect 580 825 614 847
rect 580 813 614 825
rect 580 757 614 770
rect 580 736 614 757
rect 580 689 614 693
rect 580 659 614 689
rect 580 587 614 616
rect 580 582 614 587
rect 580 519 614 539
rect 580 505 614 519
rect 580 451 614 462
rect 580 428 614 451
rect 580 383 614 385
rect 580 351 614 383
rect 580 281 614 308
rect 580 274 614 281
rect 580 213 614 231
rect 580 197 614 213
rect 736 1063 770 1077
rect 736 1043 770 1063
rect 736 995 770 1002
rect 736 968 770 995
rect 736 893 770 927
rect 736 825 770 852
rect 736 818 770 825
rect 736 757 770 777
rect 736 743 770 757
rect 736 689 770 702
rect 736 668 770 689
rect 736 621 770 626
rect 736 592 770 621
rect 736 519 770 550
rect 736 516 770 519
rect 736 451 770 474
rect 736 440 770 451
rect 736 383 770 398
rect 736 364 770 383
rect 736 315 770 322
rect 736 288 770 315
rect 892 1134 926 1168
rect 892 1063 926 1095
rect 892 1061 926 1063
rect 892 995 926 1021
rect 892 987 926 995
rect 892 927 926 947
rect 892 913 926 927
rect 892 859 926 873
rect 892 839 926 859
rect 892 791 926 799
rect 892 765 926 791
rect 892 723 926 725
rect 892 691 926 723
rect 892 621 926 651
rect 892 617 926 621
rect 892 553 926 577
rect 892 543 926 553
rect 892 485 926 503
rect 892 469 926 485
rect 892 417 926 429
rect 892 395 926 417
rect 1048 1063 1082 1077
rect 1048 1043 1082 1063
rect 1048 995 1082 1002
rect 1048 968 1082 995
rect 1048 893 1082 927
rect 1048 825 1082 852
rect 1048 818 1082 825
rect 1048 757 1082 777
rect 1048 743 1082 757
rect 1048 689 1082 702
rect 1048 668 1082 689
rect 1048 621 1082 626
rect 1048 592 1082 621
rect 1048 519 1082 550
rect 1048 516 1082 519
rect 1048 451 1082 474
rect 1048 440 1082 451
rect 1048 383 1082 398
rect 1048 364 1082 383
rect 1048 315 1082 322
rect 1048 288 1082 315
rect 1204 1134 1238 1168
rect 1204 1063 1238 1092
rect 1204 1058 1238 1063
rect 1204 995 1238 1016
rect 1204 982 1238 995
rect 1204 927 1238 940
rect 1204 906 1238 927
rect 1204 859 1238 864
rect 1204 830 1238 859
rect 1204 757 1238 788
rect 1204 754 1238 757
rect 1204 689 1238 711
rect 1204 677 1238 689
rect 1204 621 1238 634
rect 1204 600 1238 621
rect 1204 553 1238 557
rect 1204 523 1238 553
rect 1204 451 1238 480
rect 1204 446 1238 451
rect 1204 383 1238 403
rect 1204 369 1238 383
rect 1204 315 1238 326
rect 1204 292 1238 315
rect 1360 1063 1394 1077
rect 1360 1043 1394 1063
rect 1360 995 1394 1001
rect 1360 967 1394 995
rect 1360 893 1394 924
rect 1360 890 1394 893
rect 1360 825 1394 847
rect 1360 813 1394 825
rect 1360 757 1394 770
rect 1360 736 1394 757
rect 1360 689 1394 693
rect 1360 659 1394 689
rect 1360 587 1394 616
rect 1360 582 1394 587
rect 1360 519 1394 539
rect 1360 505 1394 519
rect 1360 451 1394 462
rect 1360 428 1394 451
rect 1360 383 1394 385
rect 1360 351 1394 383
rect 1360 281 1394 308
rect 1360 274 1394 281
rect 1360 213 1394 231
rect 1360 197 1394 213
rect 1516 1134 1550 1168
rect 1516 1063 1550 1092
rect 1516 1058 1550 1063
rect 1516 995 1550 1016
rect 1516 982 1550 995
rect 1516 927 1550 940
rect 1516 906 1550 927
rect 1516 859 1550 864
rect 1516 830 1550 859
rect 1516 757 1550 788
rect 1516 754 1550 757
rect 1516 689 1550 711
rect 1516 677 1550 689
rect 1516 621 1550 634
rect 1516 600 1550 621
rect 1516 553 1550 557
rect 1516 523 1550 553
rect 1516 451 1550 480
rect 1516 446 1550 451
rect 1516 383 1550 403
rect 1516 369 1550 383
rect 1516 315 1550 326
rect 1516 292 1550 315
rect 1672 1063 1706 1077
rect 1672 1043 1706 1063
rect 1672 995 1706 1001
rect 1672 967 1706 995
rect 1672 893 1706 924
rect 1672 890 1706 893
rect 1672 825 1706 847
rect 1672 813 1706 825
rect 1672 757 1706 770
rect 1672 736 1706 757
rect 1672 689 1706 693
rect 1672 659 1706 689
rect 1672 587 1706 616
rect 1672 582 1706 587
rect 1672 519 1706 539
rect 1672 505 1706 519
rect 1672 451 1706 462
rect 1672 428 1706 451
rect 1672 383 1706 385
rect 1672 351 1706 383
rect 1672 281 1706 308
rect 1672 274 1706 281
rect 1672 213 1706 231
rect 1672 197 1706 213
rect 1828 1134 1862 1168
rect 1828 1063 1862 1092
rect 1828 1058 1862 1063
rect 1828 995 1862 1016
rect 1828 982 1862 995
rect 1828 927 1862 940
rect 1828 906 1862 927
rect 1828 859 1862 864
rect 1828 830 1862 859
rect 1828 757 1862 788
rect 1828 754 1862 757
rect 1828 689 1862 711
rect 1828 677 1862 689
rect 1828 621 1862 634
rect 1828 600 1862 621
rect 1828 553 1862 557
rect 1828 523 1862 553
rect 1828 451 1862 480
rect 1828 446 1862 451
rect 1828 383 1862 403
rect 1828 369 1862 383
rect 1828 315 1862 326
rect 1828 292 1862 315
rect 1938 1134 1972 1168
rect 1938 1063 1972 1092
rect 1938 1058 1972 1063
rect 1938 995 1972 1016
rect 1938 982 1972 995
rect 1938 927 1972 940
rect 1938 906 1972 927
rect 1938 859 1972 864
rect 1938 830 1972 859
rect 1938 757 1972 788
rect 1938 754 1972 757
rect 1938 689 1972 711
rect 1938 677 1972 689
rect 1938 621 1972 634
rect 1938 600 1972 621
rect 1938 553 1972 557
rect 1938 523 1972 553
rect 1938 451 1972 480
rect 1938 446 1972 451
rect 1938 383 1972 403
rect 1938 369 1972 383
rect 1938 315 1972 326
rect 1938 292 1972 315
rect 2094 1063 2128 1077
rect 2094 1043 2128 1063
rect 2094 995 2128 1001
rect 2094 967 2128 995
rect 2094 893 2128 924
rect 2094 890 2128 893
rect 2094 825 2128 847
rect 2094 813 2128 825
rect 2094 757 2128 770
rect 2094 736 2128 757
rect 2094 689 2128 693
rect 2094 659 2128 689
rect 2094 587 2128 616
rect 2094 582 2128 587
rect 2094 519 2128 539
rect 2094 505 2128 519
rect 2094 451 2128 462
rect 2094 428 2128 451
rect 2094 383 2128 385
rect 2094 351 2128 383
rect 2094 281 2128 308
rect 2094 274 2128 281
rect 2094 213 2128 231
rect 2094 197 2128 213
rect 2250 1134 2284 1168
rect 2250 1063 2284 1092
rect 2250 1058 2284 1063
rect 2250 995 2284 1016
rect 2250 982 2284 995
rect 2250 927 2284 940
rect 2250 906 2284 927
rect 2250 859 2284 864
rect 2250 830 2284 859
rect 2250 757 2284 788
rect 2250 754 2284 757
rect 2250 689 2284 711
rect 2250 677 2284 689
rect 2250 621 2284 634
rect 2250 600 2284 621
rect 2250 553 2284 557
rect 2250 523 2284 553
rect 2250 451 2284 480
rect 2250 446 2284 451
rect 2250 383 2284 403
rect 2250 369 2284 383
rect 2250 315 2284 326
rect 2250 292 2284 315
rect 2406 1063 2440 1077
rect 2406 1043 2440 1063
rect 2406 995 2440 1001
rect 2406 967 2440 995
rect 2406 893 2440 924
rect 2406 890 2440 893
rect 2406 825 2440 847
rect 2406 813 2440 825
rect 2406 757 2440 770
rect 2406 736 2440 757
rect 2406 689 2440 693
rect 2406 659 2440 689
rect 2406 587 2440 616
rect 2406 582 2440 587
rect 2406 519 2440 539
rect 2406 505 2440 519
rect 2406 451 2440 462
rect 2406 428 2440 451
rect 2406 383 2440 385
rect 2406 351 2440 383
rect 2406 281 2440 308
rect 2406 274 2440 281
rect 2406 213 2440 231
rect 2406 197 2440 213
rect 2562 1134 2596 1168
rect 2562 1063 2596 1092
rect 2562 1058 2596 1063
rect 2562 995 2596 1016
rect 2562 982 2596 995
rect 2562 927 2596 940
rect 2562 906 2596 927
rect 2562 859 2596 864
rect 2562 830 2596 859
rect 2562 757 2596 788
rect 2562 754 2596 757
rect 2562 689 2596 711
rect 2562 677 2596 689
rect 2562 621 2596 634
rect 2562 600 2596 621
rect 2562 553 2596 557
rect 2562 523 2596 553
rect 2562 451 2596 480
rect 2562 446 2596 451
rect 2562 383 2596 403
rect 2562 369 2596 383
rect 2562 315 2596 326
rect 2562 292 2596 315
rect 2718 1063 2752 1077
rect 2718 1043 2752 1063
rect 2718 995 2752 1002
rect 2718 968 2752 995
rect 2718 893 2752 927
rect 2718 825 2752 852
rect 2718 818 2752 825
rect 2718 757 2752 777
rect 2718 743 2752 757
rect 2718 689 2752 702
rect 2718 668 2752 689
rect 2718 621 2752 627
rect 2718 593 2752 621
rect 2718 519 2752 552
rect 2718 518 2752 519
rect 2718 451 2752 477
rect 2718 443 2752 451
rect 2718 383 2752 402
rect 2718 368 2752 383
rect 2718 315 2752 326
rect 2718 292 2752 315
rect 2874 1134 2908 1168
rect 2874 1063 2908 1095
rect 2874 1061 2908 1063
rect 2874 995 2908 1022
rect 2874 988 2908 995
rect 2874 927 2908 949
rect 2874 915 2908 927
rect 2874 859 2908 876
rect 2874 842 2908 859
rect 2874 791 2908 803
rect 2874 769 2908 791
rect 2874 723 2908 730
rect 2874 696 2908 723
rect 2874 655 2908 657
rect 2874 623 2908 655
rect 2874 553 2908 583
rect 2874 549 2908 553
rect 2874 485 2908 509
rect 2874 475 2908 485
rect 2874 417 2908 435
rect 2874 401 2908 417
rect 3030 1063 3064 1077
rect 3030 1043 3064 1063
rect 3030 995 3064 1002
rect 3030 968 3064 995
rect 3030 893 3064 927
rect 3030 825 3064 852
rect 3030 818 3064 825
rect 3030 757 3064 777
rect 3030 743 3064 757
rect 3030 689 3064 702
rect 3030 668 3064 689
rect 3030 621 3064 627
rect 3030 593 3064 621
rect 3030 519 3064 552
rect 3030 518 3064 519
rect 3030 451 3064 477
rect 3030 443 3064 451
rect 3030 383 3064 402
rect 3030 368 3064 383
rect 3030 315 3064 326
rect 3030 292 3064 315
rect 616 91 618 125
rect 618 91 650 125
rect 689 91 721 125
rect 721 91 723 125
rect 762 91 790 125
rect 790 91 796 125
rect 835 91 859 125
rect 859 91 869 125
rect 908 91 928 125
rect 928 91 942 125
rect 981 91 997 125
rect 997 91 1015 125
rect 1054 91 1066 125
rect 1066 91 1088 125
rect 1128 91 1135 125
rect 1135 91 1162 125
rect 1202 91 1204 125
rect 1204 91 1236 125
rect 1276 91 1308 125
rect 1308 91 1310 125
rect 1350 91 1377 125
rect 1377 91 1384 125
rect 1424 91 1446 125
rect 1446 91 1458 125
rect 1498 91 1515 125
rect 1515 91 1532 125
rect 1572 91 1584 125
rect 1584 91 1606 125
rect 1646 91 1653 125
rect 1653 91 1680 125
rect 1720 91 1722 125
rect 1722 91 1754 125
rect 1794 91 1825 125
rect 1825 91 1828 125
rect 1868 91 1895 125
rect 1895 91 1902 125
rect 1942 91 1965 125
rect 1965 91 1976 125
rect 2016 91 2035 125
rect 2035 91 2050 125
rect 2090 91 2105 125
rect 2105 91 2124 125
rect 2164 91 2175 125
rect 2175 91 2198 125
rect 2238 91 2245 125
rect 2245 91 2272 125
rect 2312 91 2315 125
rect 2315 91 2346 125
rect 2386 91 2420 125
rect 2460 91 2491 125
rect 2491 91 2494 125
rect 2534 91 2561 125
rect 2561 91 2568 125
rect 2608 91 2631 125
rect 2631 91 2642 125
rect 2682 91 2701 125
rect 2701 91 2716 125
rect 2756 91 2771 125
rect 2771 91 2790 125
rect 2830 91 2841 125
rect 2841 91 2864 125
rect 2904 91 2911 125
rect 2911 91 2938 125
rect 2978 91 2981 125
rect 2981 91 3012 125
<< metal1 >>
rect 591 3984 4076 4051
rect 591 3950 603 3984
rect 637 3950 677 3984
rect 711 3950 751 3984
rect 785 3950 825 3984
rect 859 3950 899 3984
rect 933 3950 973 3984
rect 1007 3950 1047 3984
rect 1081 3950 1121 3984
rect 1155 3950 1195 3984
rect 1229 3950 1269 3984
rect 1303 3950 1343 3984
rect 1377 3950 1417 3984
rect 1451 3950 1491 3984
rect 1525 3950 1565 3984
rect 1599 3950 1639 3984
rect 1673 3950 1712 3984
rect 1746 3950 1785 3984
rect 1819 3950 1858 3984
rect 1892 3950 1931 3984
rect 1965 3950 2004 3984
rect 2038 3950 2077 3984
rect 2111 3950 2150 3984
rect 2184 3950 2223 3984
rect 2257 3950 2296 3984
rect 2330 3950 2369 3984
rect 2403 3950 2442 3984
rect 2476 3950 2515 3984
rect 2549 3950 2588 3984
rect 2622 3950 2661 3984
rect 2695 3950 2734 3984
rect 2768 3950 2807 3984
rect 2841 3950 2880 3984
rect 2914 3950 2953 3984
rect 2987 3950 3026 3984
rect 3060 3950 3099 3984
rect 3133 3950 3172 3984
rect 3206 3950 3245 3984
rect 3279 3950 3318 3984
rect 3352 3950 3391 3984
rect 3425 3950 3464 3984
rect 3498 3950 3537 3984
rect 3571 3950 3610 3984
rect 3644 3950 3683 3984
rect 3717 3950 3756 3984
rect 3790 3950 3829 3984
rect 3863 3950 3902 3984
rect 3936 3950 3975 3984
rect 4009 3950 4076 3984
rect 591 3880 4076 3950
rect 591 3846 1766 3880
rect 1800 3846 2188 3880
rect 2222 3846 3078 3880
rect 3112 3846 3344 3880
rect 3378 3846 3656 3880
rect 3690 3846 3968 3880
rect 4002 3846 4076 3880
rect 591 3805 4076 3846
rect 591 3804 3344 3805
rect 591 3783 1766 3804
tri 726 3770 739 3783 ne
rect 739 3770 827 3783
tri 827 3770 840 3783 nw
tri 992 3770 1005 3783 ne
rect 1005 3770 1093 3783
tri 1093 3770 1106 3783 nw
tri 1726 3770 1739 3783 ne
rect 1739 3770 1766 3783
rect 1800 3783 2188 3804
rect 1800 3770 1827 3783
tri 1827 3770 1840 3783 nw
tri 2148 3770 2161 3783 ne
rect 2161 3770 2188 3783
rect 2222 3803 3344 3804
rect 2222 3783 3078 3803
rect 2222 3770 2248 3783
tri 739 3769 740 3770 ne
rect 740 3769 826 3770
tri 826 3769 827 3770 nw
tri 1005 3769 1006 3770 ne
rect 1006 3769 1092 3770
tri 1092 3769 1093 3770 nw
tri 1739 3769 1740 3770 ne
rect 1740 3769 1826 3770
tri 1826 3769 1827 3770 nw
tri 2161 3769 2162 3770 ne
rect 2162 3769 2248 3770
tri 2248 3769 2262 3783 nw
tri 3038 3769 3052 3783 ne
rect 3052 3769 3078 3783
rect 3112 3783 3344 3803
rect 3112 3771 3140 3783
tri 3140 3771 3152 3783 nw
tri 3304 3771 3316 3783 ne
rect 3316 3771 3344 3783
rect 3378 3783 3656 3805
rect 3378 3771 3406 3783
tri 3406 3771 3418 3783 nw
tri 3616 3771 3628 3783 ne
rect 3628 3771 3656 3783
rect 3690 3783 3968 3805
rect 3690 3771 3718 3783
tri 3718 3771 3730 3783 nw
tri 3928 3771 3940 3783 ne
rect 3940 3771 3968 3783
rect 4002 3783 4076 3805
rect 4002 3771 4008 3783
rect 3112 3769 3118 3771
tri 740 3749 760 3769 ne
rect 604 3200 650 3212
rect 604 3166 610 3200
rect 644 3166 650 3200
rect 604 3070 650 3166
rect 604 3036 610 3070
rect 644 3036 650 3070
rect 604 2948 650 3036
rect 760 3200 806 3769
tri 806 3749 826 3769 nw
tri 1006 3749 1026 3769 ne
rect 760 3166 766 3200
rect 800 3166 806 3200
rect 760 3120 806 3166
rect 760 3086 766 3120
rect 800 3086 806 3120
rect 760 3040 806 3086
rect 760 3006 766 3040
rect 800 3006 806 3040
rect 760 2994 806 3006
rect 913 3200 965 3212
rect 913 3166 922 3200
rect 956 3166 965 3200
rect 913 3123 965 3166
rect 913 3121 922 3123
rect 956 3121 965 3123
rect 913 3057 965 3069
rect 913 2999 965 3005
rect 1026 3200 1072 3769
tri 1072 3749 1092 3769 nw
tri 1740 3749 1760 3769 ne
rect 1760 3728 1806 3769
tri 1806 3749 1826 3769 nw
tri 2162 3749 2182 3769 ne
rect 1026 3166 1032 3200
rect 1066 3166 1072 3200
rect 1292 3711 1338 3723
rect 1292 3677 1298 3711
rect 1332 3677 1338 3711
rect 1292 3637 1338 3677
rect 1292 3603 1298 3637
rect 1332 3603 1338 3637
rect 1292 3563 1338 3603
rect 1292 3529 1298 3563
rect 1332 3529 1338 3563
rect 1292 3489 1338 3529
rect 1292 3455 1298 3489
rect 1332 3455 1338 3489
rect 1292 3414 1338 3455
rect 1292 3380 1298 3414
rect 1332 3380 1338 3414
rect 1292 3339 1338 3380
rect 1292 3305 1298 3339
rect 1332 3305 1338 3339
rect 1292 3264 1338 3305
rect 1292 3230 1298 3264
rect 1332 3230 1338 3264
rect 1292 3189 1338 3230
rect 1026 3112 1072 3166
rect 1026 3078 1032 3112
rect 1066 3078 1072 3112
rect 1026 3023 1072 3078
rect 1026 2989 1032 3023
rect 1066 2989 1072 3023
rect 1026 2977 1072 2989
rect 1182 3164 1228 3176
rect 1182 3130 1188 3164
rect 1222 3130 1228 3164
rect 1182 3065 1228 3130
rect 1182 3031 1188 3065
rect 1222 3031 1228 3065
tri 650 2948 664 2962 sw
rect 604 2942 664 2948
tri 604 2930 616 2942 ne
rect 616 2930 664 2942
tri 664 2930 682 2948 sw
tri 616 2929 617 2930 ne
rect 617 2929 682 2930
tri 682 2929 683 2930 sw
tri 617 2882 664 2929 ne
rect 664 2928 683 2929
tri 683 2928 684 2929 sw
rect 664 2912 842 2928
tri 842 2912 858 2928 sw
rect 664 2882 858 2912
tri 822 2846 858 2882 ne
tri 858 2846 924 2912 sw
rect 858 2834 924 2846
tri 924 2834 936 2846 sw
rect 1182 2837 1228 3031
rect 1292 3155 1298 3189
rect 1332 3155 1338 3189
rect 1292 3114 1338 3155
rect 1292 3080 1298 3114
rect 1332 3080 1338 3114
rect 1292 3039 1338 3080
rect 1292 3005 1298 3039
rect 1332 3005 1338 3039
rect 1292 2989 1338 3005
rect 1445 3711 1497 3723
rect 1445 3677 1454 3711
rect 1488 3677 1497 3711
rect 1445 3637 1497 3677
rect 1445 3603 1454 3637
rect 1488 3603 1497 3637
rect 1445 3563 1497 3603
rect 1445 3529 1454 3563
rect 1488 3529 1497 3563
rect 1445 3489 1497 3529
rect 1445 3455 1454 3489
rect 1488 3455 1497 3489
rect 1445 3415 1497 3455
rect 1445 3381 1454 3415
rect 1488 3381 1497 3415
rect 1445 3340 1497 3381
rect 1445 3306 1454 3340
rect 1488 3306 1497 3340
rect 1445 3265 1497 3306
rect 1445 3231 1454 3265
rect 1488 3231 1497 3265
rect 1445 3190 1497 3231
rect 1445 3156 1454 3190
rect 1488 3156 1497 3190
rect 1445 3148 1497 3156
rect 1445 3084 1454 3096
rect 1488 3084 1497 3096
rect 1445 3006 1454 3032
rect 1488 3006 1497 3032
tri 1338 2989 1349 3000 sw
rect 1445 2994 1497 3006
rect 1604 3711 1650 3723
rect 1604 3677 1610 3711
rect 1644 3677 1650 3711
rect 1604 3637 1650 3677
rect 1604 3603 1610 3637
rect 1644 3603 1650 3637
rect 1604 3563 1650 3603
rect 1604 3529 1610 3563
rect 1644 3529 1650 3563
rect 1604 3489 1650 3529
rect 1604 3455 1610 3489
rect 1644 3455 1650 3489
rect 1604 3414 1650 3455
rect 1604 3380 1610 3414
rect 1644 3380 1650 3414
rect 1604 3339 1650 3380
rect 1604 3305 1610 3339
rect 1644 3305 1650 3339
rect 1604 3264 1650 3305
rect 1604 3230 1610 3264
rect 1644 3230 1650 3264
rect 1604 3189 1650 3230
rect 1604 3155 1610 3189
rect 1644 3155 1650 3189
rect 1604 3114 1650 3155
rect 1604 3080 1610 3114
rect 1644 3080 1650 3114
rect 1604 3039 1650 3080
rect 1604 3005 1610 3039
rect 1644 3005 1650 3039
tri 1598 2994 1604 3000 se
rect 1604 2994 1650 3005
rect 1760 3694 1766 3728
rect 1800 3694 1806 3728
rect 2182 3728 2228 3769
tri 2228 3749 2248 3769 nw
tri 3052 3749 3072 3769 ne
rect 1760 3652 1806 3694
rect 1760 3618 1766 3652
rect 1800 3618 1806 3652
rect 1760 3576 1806 3618
rect 1760 3542 1766 3576
rect 1800 3542 1806 3576
rect 1760 3500 1806 3542
rect 1760 3466 1766 3500
rect 1800 3466 1806 3500
rect 1760 3424 1806 3466
rect 1760 3390 1766 3424
rect 1800 3390 1806 3424
rect 1760 3348 1806 3390
rect 1760 3314 1766 3348
rect 1800 3314 1806 3348
rect 1760 3271 1806 3314
rect 1760 3237 1766 3271
rect 1800 3237 1806 3271
rect 1760 3194 1806 3237
rect 1760 3160 1766 3194
rect 1800 3160 1806 3194
rect 1760 3117 1806 3160
rect 1760 3083 1766 3117
rect 1800 3083 1806 3117
rect 1760 3040 1806 3083
rect 1760 3006 1766 3040
rect 1800 3006 1806 3040
tri 1593 2989 1598 2994 se
rect 1598 2989 1650 2994
tri 1650 2989 1661 3000 sw
rect 1760 2994 1806 3006
rect 1916 3711 1962 3723
rect 1916 3677 1922 3711
rect 1956 3677 1962 3711
rect 1916 3637 1962 3677
rect 1916 3603 1922 3637
rect 1956 3603 1962 3637
rect 1916 3563 1962 3603
rect 1916 3529 1922 3563
rect 1956 3529 1962 3563
rect 1916 3489 1962 3529
rect 1916 3455 1922 3489
rect 1956 3455 1962 3489
rect 1916 3414 1962 3455
rect 1916 3380 1922 3414
rect 1956 3380 1962 3414
rect 1916 3339 1962 3380
rect 1916 3305 1922 3339
rect 1956 3305 1962 3339
rect 1916 3264 1962 3305
rect 1916 3230 1922 3264
rect 1956 3230 1962 3264
rect 1916 3189 1962 3230
rect 1916 3155 1922 3189
rect 1956 3155 1962 3189
rect 1916 3114 1962 3155
rect 1916 3080 1922 3114
rect 1956 3080 1962 3114
rect 1916 3039 1962 3080
rect 1916 3005 1922 3039
rect 1956 3005 1962 3039
tri 1910 2994 1916 3000 se
rect 1916 2994 1962 3005
tri 1905 2989 1910 2994 se
rect 1910 2989 1962 2994
rect 1292 2966 1349 2989
tri 1349 2966 1372 2989 sw
tri 1570 2966 1593 2989 se
rect 1593 2966 1661 2989
tri 1661 2966 1684 2989 sw
tri 1882 2966 1905 2989 se
rect 1905 2966 1962 2989
rect 1292 2964 1962 2966
rect 1292 2930 1298 2964
rect 1332 2930 1610 2964
rect 1644 2930 1922 2964
rect 1956 2930 1962 2964
tri 1228 2837 1262 2871 sw
rect 1292 2866 1962 2930
rect 2026 3711 2072 3723
rect 2026 3677 2032 3711
rect 2066 3677 2072 3711
rect 2026 3637 2072 3677
rect 2026 3603 2032 3637
rect 2066 3603 2072 3637
rect 2026 3563 2072 3603
rect 2026 3529 2032 3563
rect 2066 3529 2072 3563
rect 2026 3489 2072 3529
rect 2026 3455 2032 3489
rect 2066 3455 2072 3489
rect 2026 3414 2072 3455
rect 2026 3380 2032 3414
rect 2066 3380 2072 3414
rect 2026 3339 2072 3380
rect 2026 3305 2032 3339
rect 2066 3305 2072 3339
rect 2026 3264 2072 3305
rect 2026 3230 2032 3264
rect 2066 3230 2072 3264
rect 2026 3189 2072 3230
rect 2026 3155 2032 3189
rect 2066 3155 2072 3189
rect 2026 3114 2072 3155
rect 2026 3080 2032 3114
rect 2066 3080 2072 3114
rect 2026 3039 2072 3080
rect 2026 3005 2032 3039
rect 2066 3005 2072 3039
rect 2026 2989 2072 3005
rect 2182 3694 2188 3728
rect 2222 3694 2228 3728
rect 3072 3725 3118 3769
tri 3118 3749 3140 3771 nw
tri 3316 3749 3338 3771 ne
rect 2182 3652 2228 3694
rect 2182 3618 2188 3652
rect 2222 3618 2228 3652
rect 2182 3576 2228 3618
rect 2182 3542 2188 3576
rect 2222 3542 2228 3576
rect 2182 3500 2228 3542
rect 2182 3466 2188 3500
rect 2222 3466 2228 3500
rect 2182 3424 2228 3466
rect 2182 3390 2188 3424
rect 2222 3390 2228 3424
rect 2182 3348 2228 3390
rect 2182 3314 2188 3348
rect 2222 3314 2228 3348
rect 2182 3271 2228 3314
rect 2182 3237 2188 3271
rect 2222 3237 2228 3271
rect 2182 3194 2228 3237
rect 2182 3160 2188 3194
rect 2222 3160 2228 3194
rect 2182 3117 2228 3160
rect 2182 3083 2188 3117
rect 2222 3083 2228 3117
rect 2182 3040 2228 3083
rect 2182 3006 2188 3040
rect 2222 3006 2228 3040
tri 2072 2989 2083 3000 sw
rect 2182 2994 2228 3006
rect 2338 3711 2384 3723
rect 2338 3677 2344 3711
rect 2378 3677 2384 3711
rect 2338 3637 2384 3677
rect 2338 3603 2344 3637
rect 2378 3603 2384 3637
rect 2338 3563 2384 3603
rect 2338 3529 2344 3563
rect 2378 3529 2384 3563
rect 2338 3489 2384 3529
rect 2338 3455 2344 3489
rect 2378 3455 2384 3489
rect 2338 3414 2384 3455
rect 2338 3380 2344 3414
rect 2378 3380 2384 3414
rect 2338 3339 2384 3380
rect 2338 3305 2344 3339
rect 2378 3305 2384 3339
rect 2338 3264 2384 3305
rect 2338 3230 2344 3264
rect 2378 3230 2384 3264
rect 2338 3189 2384 3230
rect 2338 3155 2344 3189
rect 2378 3155 2384 3189
rect 2338 3114 2384 3155
rect 2338 3080 2344 3114
rect 2378 3080 2384 3114
rect 2338 3039 2384 3080
rect 2338 3005 2344 3039
rect 2378 3005 2384 3039
tri 2332 2994 2338 3000 se
rect 2338 2994 2384 3005
rect 2492 3711 2544 3723
rect 2492 3677 2500 3711
rect 2534 3677 2544 3711
rect 2492 3637 2544 3677
rect 2492 3603 2500 3637
rect 2534 3603 2544 3637
rect 2492 3563 2544 3603
rect 2492 3529 2500 3563
rect 2534 3529 2544 3563
rect 2492 3489 2544 3529
rect 2492 3455 2500 3489
rect 2534 3455 2544 3489
rect 2492 3415 2544 3455
rect 2492 3381 2500 3415
rect 2534 3381 2544 3415
rect 2492 3340 2544 3381
rect 2492 3306 2500 3340
rect 2534 3306 2544 3340
rect 2492 3265 2544 3306
rect 2492 3231 2500 3265
rect 2534 3231 2544 3265
rect 2492 3190 2544 3231
rect 2492 3156 2500 3190
rect 2534 3156 2544 3190
rect 2492 3148 2544 3156
rect 2492 3084 2500 3096
rect 2534 3084 2544 3096
rect 2492 3006 2500 3032
rect 2534 3006 2544 3032
tri 2327 2989 2332 2994 se
rect 2332 2989 2384 2994
tri 2384 2989 2395 3000 sw
rect 2492 2994 2544 3006
rect 2650 3711 2696 3723
rect 2650 3677 2656 3711
rect 2690 3677 2696 3711
rect 2650 3637 2696 3677
rect 2650 3603 2656 3637
rect 2690 3603 2696 3637
rect 2650 3563 2696 3603
rect 2650 3529 2656 3563
rect 2690 3529 2696 3563
rect 2650 3489 2696 3529
rect 2650 3455 2656 3489
rect 2690 3455 2696 3489
rect 2650 3414 2696 3455
rect 2650 3380 2656 3414
rect 2690 3380 2696 3414
rect 2650 3339 2696 3380
rect 2650 3305 2656 3339
rect 2690 3305 2696 3339
rect 2650 3264 2696 3305
rect 2650 3230 2656 3264
rect 2690 3230 2696 3264
rect 2650 3189 2696 3230
rect 2650 3155 2656 3189
rect 2690 3155 2696 3189
rect 2650 3114 2696 3155
rect 2650 3080 2656 3114
rect 2690 3080 2696 3114
rect 2650 3039 2696 3080
rect 2650 3005 2656 3039
rect 2690 3005 2696 3039
tri 2644 2994 2650 3000 se
rect 2650 2994 2696 3005
rect 2757 3711 2809 3723
rect 2757 3677 2766 3711
rect 2800 3677 2809 3711
rect 2757 3637 2809 3677
rect 2757 3603 2766 3637
rect 2800 3603 2809 3637
rect 2757 3563 2809 3603
rect 2757 3529 2766 3563
rect 2800 3529 2809 3563
rect 2757 3489 2809 3529
rect 2757 3455 2766 3489
rect 2800 3455 2809 3489
rect 2757 3415 2809 3455
rect 2757 3381 2766 3415
rect 2800 3381 2809 3415
rect 2757 3340 2809 3381
rect 2757 3306 2766 3340
rect 2800 3306 2809 3340
rect 2757 3265 2809 3306
rect 2757 3231 2766 3265
rect 2800 3231 2809 3265
rect 2757 3190 2809 3231
rect 2757 3156 2766 3190
rect 2800 3156 2809 3190
rect 2757 3148 2809 3156
rect 2757 3084 2766 3096
rect 2800 3084 2809 3096
rect 2757 3006 2766 3032
rect 2800 3006 2809 3032
rect 2757 2994 2809 3006
rect 2916 3711 2962 3723
rect 2916 3677 2922 3711
rect 2956 3677 2962 3711
rect 2916 3637 2962 3677
rect 2916 3603 2922 3637
rect 2956 3603 2962 3637
rect 2916 3563 2962 3603
rect 2916 3529 2922 3563
rect 2956 3529 2962 3563
rect 2916 3489 2962 3529
rect 2916 3455 2922 3489
rect 2956 3455 2962 3489
rect 2916 3415 2962 3455
rect 2916 3381 2922 3415
rect 2956 3381 2962 3415
rect 2916 3340 2962 3381
rect 2916 3306 2922 3340
rect 2956 3306 2962 3340
rect 2916 3265 2962 3306
rect 2916 3231 2922 3265
rect 2956 3231 2962 3265
rect 2916 3190 2962 3231
rect 2916 3156 2922 3190
rect 2956 3156 2962 3190
rect 2916 3115 2962 3156
rect 2916 3081 2922 3115
rect 2956 3081 2962 3115
rect 2916 3040 2962 3081
rect 2916 3006 2922 3040
rect 2956 3006 2962 3040
rect 2916 2994 2962 3006
rect 3072 3691 3078 3725
rect 3112 3691 3118 3725
rect 3338 3730 3384 3771
tri 3384 3749 3406 3771 nw
tri 3628 3749 3650 3771 ne
rect 3072 3647 3118 3691
rect 3072 3613 3078 3647
rect 3112 3613 3118 3647
rect 3072 3569 3118 3613
rect 3072 3535 3078 3569
rect 3112 3535 3118 3569
rect 3072 3491 3118 3535
rect 3072 3457 3078 3491
rect 3112 3457 3118 3491
rect 3072 3413 3118 3457
rect 3072 3379 3078 3413
rect 3112 3379 3118 3413
rect 3072 3335 3118 3379
rect 3072 3301 3078 3335
rect 3112 3301 3118 3335
rect 3072 3257 3118 3301
rect 3072 3223 3078 3257
rect 3112 3223 3118 3257
rect 3072 3179 3118 3223
rect 3072 3145 3078 3179
rect 3112 3145 3118 3179
rect 3072 3101 3118 3145
rect 3072 3067 3078 3101
rect 3112 3067 3118 3101
rect 3072 3023 3118 3067
tri 2639 2989 2644 2994 se
rect 2644 2989 2696 2994
rect 2026 2966 2083 2989
tri 2083 2966 2106 2989 sw
tri 2304 2966 2327 2989 se
rect 2327 2966 2395 2989
tri 2395 2966 2418 2989 sw
tri 2616 2966 2639 2989 se
rect 2639 2966 2696 2989
rect 3072 2989 3078 3023
rect 3112 2989 3118 3023
rect 3072 2977 3118 2989
rect 3182 3711 3228 3723
rect 3182 3677 3188 3711
rect 3222 3677 3228 3711
rect 3182 3637 3228 3677
rect 3182 3603 3188 3637
rect 3222 3603 3228 3637
rect 3182 3563 3228 3603
rect 3182 3529 3188 3563
rect 3222 3529 3228 3563
rect 3182 3488 3228 3529
rect 3182 3454 3188 3488
rect 3222 3454 3228 3488
rect 3182 3413 3228 3454
rect 3182 3379 3188 3413
rect 3222 3379 3228 3413
rect 3182 3338 3228 3379
rect 3182 3304 3188 3338
rect 3222 3304 3228 3338
rect 3182 3263 3228 3304
rect 3182 3229 3188 3263
rect 3222 3229 3228 3263
rect 3182 3188 3228 3229
rect 3182 3154 3188 3188
rect 3222 3154 3228 3188
rect 3182 3113 3228 3154
rect 3182 3079 3188 3113
rect 3222 3079 3228 3113
rect 3182 3038 3228 3079
rect 3182 3004 3188 3038
rect 3222 3004 3228 3038
rect 3338 3696 3344 3730
rect 3378 3696 3384 3730
rect 3650 3730 3696 3771
tri 3696 3749 3718 3771 nw
tri 3940 3749 3962 3771 ne
rect 3338 3655 3384 3696
rect 3338 3621 3344 3655
rect 3378 3621 3384 3655
rect 3338 3580 3384 3621
rect 3338 3546 3344 3580
rect 3378 3546 3384 3580
rect 3338 3505 3384 3546
rect 3338 3471 3344 3505
rect 3378 3471 3384 3505
rect 3338 3430 3384 3471
rect 3338 3396 3344 3430
rect 3378 3396 3384 3430
rect 3338 3355 3384 3396
rect 3338 3321 3344 3355
rect 3378 3321 3384 3355
rect 3338 3280 3384 3321
rect 3338 3246 3344 3280
rect 3378 3246 3384 3280
rect 3338 3204 3384 3246
rect 3338 3170 3344 3204
rect 3378 3170 3384 3204
rect 3338 3128 3384 3170
rect 3338 3094 3344 3128
rect 3378 3094 3384 3128
rect 3338 3052 3384 3094
rect 3338 3018 3344 3052
rect 3378 3018 3384 3052
tri 3228 3004 3232 3008 sw
rect 3338 3006 3384 3018
rect 3494 3711 3540 3723
rect 3494 3677 3500 3711
rect 3534 3677 3540 3711
rect 3494 3637 3540 3677
rect 3494 3603 3500 3637
rect 3534 3603 3540 3637
rect 3494 3563 3540 3603
rect 3494 3529 3500 3563
rect 3534 3529 3540 3563
rect 3494 3488 3540 3529
rect 3494 3454 3500 3488
rect 3534 3454 3540 3488
rect 3494 3413 3540 3454
rect 3494 3379 3500 3413
rect 3534 3379 3540 3413
rect 3494 3338 3540 3379
rect 3494 3304 3500 3338
rect 3534 3304 3540 3338
rect 3494 3263 3540 3304
rect 3494 3229 3500 3263
rect 3534 3229 3540 3263
rect 3494 3188 3540 3229
rect 3494 3154 3500 3188
rect 3534 3154 3540 3188
rect 3494 3113 3540 3154
rect 3494 3079 3500 3113
rect 3534 3079 3540 3113
rect 3494 3038 3540 3079
tri 3492 3006 3494 3008 se
rect 3494 3006 3500 3038
tri 3490 3004 3492 3006 se
rect 3492 3004 3500 3006
rect 3534 3004 3540 3038
rect 3650 3696 3656 3730
rect 3690 3696 3696 3730
rect 3962 3730 4008 3771
tri 4008 3749 4042 3783 nw
rect 3650 3655 3696 3696
rect 3650 3621 3656 3655
rect 3690 3621 3696 3655
rect 3650 3580 3696 3621
rect 3650 3546 3656 3580
rect 3690 3546 3696 3580
rect 3650 3505 3696 3546
rect 3650 3471 3656 3505
rect 3690 3471 3696 3505
rect 3650 3430 3696 3471
rect 3650 3396 3656 3430
rect 3690 3396 3696 3430
rect 3650 3355 3696 3396
rect 3650 3321 3656 3355
rect 3690 3321 3696 3355
rect 3650 3280 3696 3321
rect 3650 3246 3656 3280
rect 3690 3246 3696 3280
rect 3650 3204 3696 3246
rect 3650 3170 3656 3204
rect 3690 3170 3696 3204
rect 3650 3128 3696 3170
rect 3650 3094 3656 3128
rect 3690 3094 3696 3128
rect 3650 3052 3696 3094
rect 3650 3018 3656 3052
rect 3690 3018 3696 3052
tri 3540 3004 3544 3008 sw
rect 3650 3006 3696 3018
rect 3806 3711 3852 3723
rect 3806 3677 3812 3711
rect 3846 3677 3852 3711
rect 3806 3637 3852 3677
rect 3806 3603 3812 3637
rect 3846 3603 3852 3637
rect 3806 3563 3852 3603
rect 3806 3529 3812 3563
rect 3846 3529 3852 3563
rect 3806 3488 3852 3529
rect 3806 3454 3812 3488
rect 3846 3454 3852 3488
rect 3806 3413 3852 3454
rect 3806 3379 3812 3413
rect 3846 3379 3852 3413
rect 3806 3338 3852 3379
rect 3806 3304 3812 3338
rect 3846 3304 3852 3338
rect 3806 3263 3852 3304
rect 3806 3229 3812 3263
rect 3846 3229 3852 3263
rect 3806 3188 3852 3229
rect 3806 3154 3812 3188
rect 3846 3154 3852 3188
rect 3806 3113 3852 3154
rect 3806 3079 3812 3113
rect 3846 3079 3852 3113
rect 3806 3038 3852 3079
tri 3804 3006 3806 3008 se
rect 3806 3006 3812 3038
tri 3802 3004 3804 3006 se
rect 3804 3004 3812 3006
rect 3846 3004 3852 3038
rect 3962 3696 3968 3730
rect 4002 3696 4008 3730
rect 3962 3655 4008 3696
rect 3962 3621 3968 3655
rect 4002 3621 4008 3655
rect 3962 3580 4008 3621
rect 3962 3546 3968 3580
rect 4002 3546 4008 3580
rect 3962 3505 4008 3546
rect 3962 3471 3968 3505
rect 4002 3471 4008 3505
rect 3962 3430 4008 3471
rect 3962 3396 3968 3430
rect 4002 3396 4008 3430
rect 3962 3355 4008 3396
rect 3962 3321 3968 3355
rect 4002 3321 4008 3355
rect 3962 3280 4008 3321
rect 3962 3246 3968 3280
rect 4002 3246 4008 3280
rect 3962 3204 4008 3246
rect 3962 3170 3968 3204
rect 4002 3170 4008 3204
rect 3962 3128 4008 3170
rect 3962 3094 3968 3128
rect 4002 3094 4008 3128
rect 3962 3052 4008 3094
rect 3962 3018 3968 3052
rect 4002 3018 4008 3052
rect 3962 3006 4008 3018
rect 2026 2964 2696 2966
rect 2026 2930 2032 2964
rect 2066 2930 2344 2964
rect 2378 2930 2656 2964
rect 2690 2930 2696 2964
rect 2026 2866 2696 2930
rect 3182 2974 3232 3004
tri 3232 2974 3262 3004 sw
tri 3460 2974 3490 3004 se
rect 3490 2974 3544 3004
tri 3544 2974 3574 3004 sw
tri 3772 2974 3802 3004 se
rect 3802 2974 3852 3004
rect 3182 2963 3852 2974
rect 3182 2929 3188 2963
rect 3222 2950 3500 2963
rect 3534 2950 3812 2963
rect 3222 2929 3482 2950
rect 3182 2898 3482 2929
rect 3534 2898 3546 2950
rect 3598 2929 3812 2950
rect 3846 2929 3852 2963
rect 3598 2898 3852 2929
rect 3182 2874 3852 2898
rect 625 2832 755 2834
rect 625 2780 633 2832
rect 685 2780 697 2832
rect 749 2780 755 2832
rect 858 2828 1104 2834
rect 858 2794 881 2828
rect 915 2794 970 2828
rect 1004 2794 1058 2828
rect 1092 2794 1104 2828
rect 858 2788 1104 2794
tri 951 2780 959 2788 ne
rect 959 2780 1104 2788
rect 1182 2785 1328 2837
rect 1380 2828 1392 2837
rect 1444 2828 1588 2837
rect 1444 2794 1455 2828
rect 1489 2794 1542 2828
rect 1576 2794 1588 2828
rect 1380 2785 1392 2794
rect 1444 2785 1588 2794
rect 1675 2828 1774 2837
rect 1675 2794 1687 2828
rect 1721 2794 1769 2828
rect 1675 2785 1774 2794
rect 1826 2785 1838 2837
rect 1890 2785 1896 2837
rect 2080 2828 2120 2837
rect 2172 2828 2184 2837
rect 2236 2828 2316 2837
rect 2080 2794 2092 2828
rect 2172 2794 2181 2828
rect 2236 2794 2270 2828
rect 2304 2794 2316 2828
rect 2080 2785 2120 2794
rect 2172 2785 2184 2794
rect 2236 2785 2316 2794
rect 2400 2828 2510 2837
rect 2400 2794 2412 2828
rect 2446 2794 2499 2828
rect 2400 2785 2510 2794
rect 2562 2785 2574 2837
rect 2626 2785 2632 2837
rect 2779 2785 2785 2837
rect 2837 2785 2849 2837
rect 2901 2785 2909 2837
rect 2967 2828 3007 2837
rect 3059 2828 3071 2837
rect 2967 2794 2979 2828
rect 2967 2785 3007 2794
rect 3059 2785 3071 2794
rect 3123 2785 3129 2837
rect 3277 2828 3324 2837
rect 3376 2828 3388 2837
rect 3440 2828 3919 2837
rect 3277 2794 3289 2828
rect 3323 2794 3324 2828
rect 3469 2794 3508 2828
rect 3542 2794 3581 2828
rect 3615 2794 3654 2828
rect 3688 2794 3727 2828
rect 3761 2794 3800 2828
rect 3834 2794 3873 2828
rect 3907 2794 3919 2828
rect 3277 2785 3324 2794
rect 3376 2785 3388 2794
rect 3440 2785 3919 2794
tri 959 2754 985 2780 ne
rect 985 2728 1104 2780
tri 1104 2728 1138 2762 sw
rect 985 2676 1444 2728
rect 1496 2676 1508 2728
rect 1560 2676 1566 2728
rect 2114 2676 2120 2728
rect 2172 2676 2184 2728
rect 2236 2676 4076 2728
rect 595 2642 1774 2648
rect 647 2596 1774 2642
rect 1826 2596 1838 2648
rect 1890 2596 4076 2648
rect 595 2578 647 2590
tri 647 2562 681 2596 nw
rect 595 2520 647 2526
rect 2386 2516 2392 2568
rect 2444 2516 2456 2568
rect 2508 2516 3083 2568
rect 3135 2516 3147 2568
rect 3199 2516 4076 2568
rect 839 2509 1808 2515
rect 839 2475 905 2509
rect 939 2475 989 2509
rect 1023 2475 1073 2509
rect 1107 2475 1157 2509
rect 1191 2475 1241 2509
rect 1275 2475 1325 2509
rect 1359 2475 1408 2509
rect 1442 2475 1808 2509
rect 839 2469 1808 2475
rect 839 2460 1642 2469
rect 839 2344 1047 2460
rect 1163 2435 1642 2460
rect 1676 2435 1808 2469
rect 1163 2397 1808 2435
rect 1848 2468 1930 2477
rect 1848 2434 1860 2468
rect 1894 2434 1930 2468
rect 1848 2425 1930 2434
rect 1982 2425 1994 2477
rect 2046 2468 2706 2477
rect 2062 2434 2111 2468
rect 2145 2434 2194 2468
rect 2228 2434 2277 2468
rect 2311 2434 2706 2468
rect 2046 2425 2706 2434
rect 2942 2468 3890 2474
rect 2942 2434 2954 2468
rect 2988 2434 3030 2468
rect 3064 2434 3106 2468
rect 3140 2434 3182 2468
rect 3216 2434 3258 2468
rect 3292 2434 3334 2468
rect 3368 2434 3410 2468
rect 3444 2434 3486 2468
rect 3520 2434 3562 2468
rect 3596 2434 3638 2468
rect 3672 2434 3704 2468
rect 2942 2428 3704 2434
tri 2626 2423 2628 2425 ne
rect 2628 2423 2706 2425
tri 3652 2423 3657 2428 ne
rect 3657 2423 3704 2428
rect 1163 2363 1642 2397
rect 1676 2363 1808 2397
tri 2628 2392 2659 2423 ne
rect 2659 2392 2706 2423
tri 3657 2394 3686 2423 ne
rect 3686 2416 3704 2423
rect 3756 2416 3768 2468
rect 3820 2457 3832 2468
rect 3820 2423 3830 2457
rect 3820 2416 3832 2423
rect 3884 2416 3890 2468
tri 2659 2391 2660 2392 ne
rect 1163 2344 1808 2363
rect 839 2333 1808 2344
rect 2416 2373 2632 2379
rect 2416 2339 2428 2373
rect 2462 2339 2500 2373
rect 2534 2339 2580 2373
rect 2416 2333 2580 2339
rect 839 2325 965 2333
tri 965 2325 973 2333 nw
tri 1602 2325 1610 2333 ne
rect 1610 2325 1808 2333
rect 839 2084 939 2325
tri 939 2299 965 2325 nw
tri 1610 2299 1636 2325 ne
rect 1636 2291 1642 2325
rect 1676 2291 1808 2325
tri 2546 2318 2561 2333 ne
rect 2561 2321 2580 2333
rect 2561 2318 2632 2321
rect 1636 2252 1808 2291
rect 1848 2312 2323 2318
tri 2561 2314 2565 2318 ne
rect 2565 2314 2632 2318
rect 1848 2278 1860 2312
rect 1894 2278 1944 2312
rect 1978 2278 2028 2312
rect 2062 2278 2111 2312
rect 2145 2278 2194 2312
rect 2228 2278 2277 2312
rect 2311 2278 2323 2312
tri 2565 2299 2580 2314 ne
rect 2580 2309 2632 2314
rect 1848 2272 2323 2278
rect 1246 2174 1252 2226
rect 1304 2217 1316 2226
rect 1368 2217 1475 2226
rect 1390 2183 1429 2217
rect 1463 2183 1475 2217
rect 1304 2174 1316 2183
rect 1368 2174 1475 2183
rect 1514 2206 1566 2222
rect 1514 2204 1523 2206
rect 1557 2204 1566 2206
rect 1514 2140 1566 2152
tri 939 2084 956 2101 sw
rect 1514 2084 1523 2088
rect 1557 2084 1566 2088
rect 839 2072 956 2084
tri 956 2072 968 2084 sw
rect 1514 2072 1566 2084
rect 1636 2218 1642 2252
rect 1676 2218 1808 2252
rect 2580 2251 2632 2257
rect 2660 2358 2666 2392
rect 2700 2358 2706 2392
rect 2660 2314 2706 2358
rect 3686 2386 3890 2416
rect 3686 2334 3704 2386
rect 3756 2334 3768 2386
rect 3820 2382 3832 2386
rect 3820 2348 3830 2382
rect 3820 2334 3832 2348
rect 3884 2334 3890 2386
rect 2660 2280 2666 2314
rect 2700 2280 2706 2314
rect 1636 2179 1808 2218
rect 1636 2145 1642 2179
rect 1676 2162 1808 2179
tri 1808 2162 1842 2196 sw
rect 2384 2187 2392 2239
rect 2444 2187 2456 2239
rect 2508 2187 2514 2239
rect 2660 2235 2706 2280
rect 2660 2201 2666 2235
rect 2700 2201 2706 2235
rect 1676 2156 2215 2162
rect 1676 2145 1752 2156
rect 1636 2122 1752 2145
rect 1786 2122 1836 2156
rect 1870 2122 1920 2156
rect 1954 2122 2003 2156
rect 2037 2122 2086 2156
rect 2120 2122 2169 2156
rect 2203 2122 2215 2156
rect 1636 2116 2215 2122
rect 2660 2156 2706 2201
rect 2660 2122 2666 2156
rect 2700 2122 2706 2156
rect 1636 2106 1808 2116
rect 1636 2072 1642 2106
rect 1676 2072 1808 2106
tri 1808 2082 1842 2116 nw
rect 839 2067 968 2072
tri 968 2067 973 2072 sw
rect 839 2061 1475 2067
rect 839 2027 1175 2061
rect 1209 2027 1260 2061
rect 1294 2027 1345 2061
rect 1379 2027 1429 2061
rect 1463 2027 1475 2061
rect 839 2021 1475 2027
rect 1636 2033 1808 2072
rect 2384 2033 2392 2085
rect 2444 2033 2456 2085
rect 2508 2033 2514 2085
rect 2660 2077 2706 2122
rect 2660 2043 2666 2077
rect 2700 2043 2706 2077
rect 1636 1999 1642 2033
rect 1676 1999 1808 2033
rect 2660 2031 2706 2043
rect 2790 2312 3482 2321
rect 2790 2278 2802 2312
rect 2836 2278 2878 2312
rect 2912 2278 2954 2312
rect 2988 2278 3030 2312
rect 3064 2278 3106 2312
rect 3140 2278 3182 2312
rect 3216 2278 3258 2312
rect 3292 2278 3334 2312
rect 3368 2278 3410 2312
rect 3444 2278 3482 2312
rect 2790 2269 3482 2278
rect 3534 2269 3546 2321
rect 3598 2269 3608 2321
rect 3686 2306 3890 2334
rect 3686 2304 3830 2306
rect 3864 2304 3890 2306
rect 2790 2009 2902 2269
tri 2902 2235 2936 2269 nw
rect 3686 2252 3704 2304
rect 3756 2252 3768 2304
rect 3820 2272 3830 2304
rect 3820 2252 3832 2272
rect 3884 2252 3890 2304
rect 3686 2230 3890 2252
rect 3686 2222 3830 2230
rect 3864 2222 3890 2230
tri 3652 2162 3686 2196 se
rect 3686 2170 3704 2222
rect 3756 2170 3768 2222
rect 3820 2196 3830 2222
rect 3820 2170 3832 2196
rect 3884 2170 3890 2222
rect 3686 2162 3890 2170
rect 2942 2156 3890 2162
rect 2942 2122 2954 2156
rect 2988 2122 3030 2156
rect 3064 2122 3106 2156
rect 3140 2122 3182 2156
rect 3216 2122 3258 2156
rect 3292 2122 3334 2156
rect 3368 2122 3410 2156
rect 3444 2122 3486 2156
rect 3520 2122 3562 2156
rect 3596 2122 3638 2156
rect 3672 2140 3714 2156
rect 3748 2154 3890 2156
rect 3748 2140 3830 2154
rect 3864 2140 3890 2154
rect 3672 2122 3704 2140
rect 2942 2116 3704 2122
tri 3652 2082 3686 2116 ne
rect 3686 2088 3704 2116
rect 3756 2088 3768 2140
rect 3820 2120 3830 2140
rect 3820 2088 3832 2120
rect 3884 2088 3890 2140
rect 3686 2082 3890 2088
tri 2902 2009 2936 2043 sw
rect 1636 1987 1808 1999
rect 1848 2000 2323 2006
rect 1848 1966 1860 2000
rect 1894 1966 1944 2000
rect 1978 1966 2028 2000
rect 2062 1966 2111 2000
rect 2145 1966 2194 2000
rect 2228 1966 2277 2000
rect 2311 1966 2323 2000
rect 1848 1960 2323 1966
rect 2790 2000 3482 2009
rect 2790 1966 2802 2000
rect 2836 1966 2878 2000
rect 2912 1966 2954 2000
rect 2988 1966 3030 2000
rect 3064 1966 3106 2000
rect 3140 1966 3182 2000
rect 3216 1966 3258 2000
rect 3292 1966 3334 2000
rect 3368 1966 3410 2000
rect 3444 1966 3482 2000
rect 2790 1957 3482 1966
rect 3534 1957 3546 2009
rect 3598 1957 3608 2009
rect 1246 1880 1252 1932
rect 1304 1880 1316 1932
rect 1368 1925 2514 1932
rect 1368 1891 2396 1925
rect 2430 1891 2468 1925
rect 2502 1891 2514 1925
rect 1368 1884 2514 1891
rect 1368 1880 1374 1884
tri 1374 1880 1378 1884 nw
rect 1848 1844 1930 1856
rect 1848 1810 1860 1844
rect 1894 1810 1930 1844
rect 1848 1804 1930 1810
rect 1982 1804 1994 1856
rect 2046 1844 2323 1856
rect 2062 1810 2111 1844
rect 2145 1810 2194 1844
rect 2228 1810 2277 1844
rect 2311 1810 2323 1844
rect 2046 1804 2323 1810
rect 621 1724 879 1776
rect 931 1724 943 1776
rect 995 1724 1001 1776
rect 621 1644 2666 1696
rect 2718 1644 2730 1696
rect 2782 1644 2788 1696
rect 1340 1496 1346 1548
rect 1398 1496 1410 1548
rect 1462 1496 2392 1548
rect 2444 1496 2456 1548
rect 2508 1496 2847 1548
rect 2899 1496 2911 1548
rect 2963 1496 3153 1548
rect 565 1416 2586 1468
rect 2638 1416 2650 1468
rect 2702 1416 3153 1468
rect 552 1240 558 1292
rect 610 1283 622 1292
rect 674 1283 725 1292
rect 674 1249 679 1283
rect 713 1249 725 1283
rect 610 1240 622 1249
rect 674 1240 725 1249
rect 796 1283 840 1292
rect 892 1283 904 1292
rect 956 1283 1181 1292
rect 796 1249 808 1283
rect 956 1249 971 1283
rect 1005 1249 1053 1283
rect 1087 1249 1135 1283
rect 1169 1249 1181 1283
rect 796 1240 840 1249
rect 892 1240 904 1249
rect 956 1240 1181 1249
rect 1264 1240 1270 1292
rect 1322 1240 1334 1292
rect 1386 1283 2414 1292
rect 1386 1249 1424 1283
rect 1458 1249 1498 1283
rect 1532 1249 1572 1283
rect 1606 1249 1646 1283
rect 1680 1249 1721 1283
rect 1755 1249 2014 1283
rect 2048 1249 2093 1283
rect 2127 1249 2172 1283
rect 2206 1249 2251 1283
rect 2285 1249 2330 1283
rect 2364 1249 2410 1283
rect 1386 1240 2414 1249
rect 2466 1240 2478 1292
rect 2530 1240 2536 1292
rect 2625 1283 2666 1292
rect 2718 1283 2730 1292
rect 2782 1283 2997 1292
rect 2625 1249 2637 1283
rect 2782 1249 2793 1283
rect 2827 1249 2872 1283
rect 2906 1249 2951 1283
rect 2985 1249 2997 1283
rect 2625 1240 2666 1249
rect 2718 1240 2730 1249
rect 2782 1240 2997 1249
rect 886 1168 1868 1203
rect 886 1134 892 1168
rect 926 1134 1204 1168
rect 1238 1134 1516 1168
rect 1550 1134 1828 1168
rect 1862 1134 1868 1168
rect 886 1123 1868 1134
rect 886 1095 938 1123
tri 938 1095 966 1123 nw
tri 1164 1095 1192 1123 ne
rect 1192 1095 1250 1123
tri 1250 1095 1278 1123 nw
tri 1476 1095 1504 1123 ne
rect 1504 1095 1562 1123
tri 1562 1095 1590 1123 nw
tri 1788 1095 1816 1123 ne
rect 1816 1095 1868 1123
rect 574 1077 620 1089
rect 574 1043 580 1077
rect 614 1043 620 1077
rect 574 1001 620 1043
rect 574 967 580 1001
rect 614 967 620 1001
rect 574 924 620 967
rect 574 890 580 924
rect 614 890 620 924
rect 574 847 620 890
rect 574 813 580 847
rect 614 813 620 847
rect 574 770 620 813
rect 574 736 580 770
rect 614 736 620 770
rect 574 693 620 736
rect 574 659 580 693
rect 614 659 620 693
rect 574 616 620 659
rect 574 582 580 616
rect 614 582 620 616
rect 574 539 620 582
rect 574 505 580 539
rect 614 505 620 539
rect 574 462 620 505
rect 574 428 580 462
rect 614 428 620 462
rect 574 385 620 428
rect 574 351 580 385
rect 614 351 620 385
rect 574 308 620 351
tri 568 274 574 280 se
rect 574 274 580 308
rect 614 274 620 308
rect 730 1077 776 1089
rect 730 1043 736 1077
rect 770 1043 776 1077
rect 730 1002 776 1043
rect 730 968 736 1002
rect 770 968 776 1002
rect 730 927 776 968
rect 730 893 736 927
rect 770 893 776 927
rect 730 852 776 893
rect 730 818 736 852
rect 770 818 776 852
rect 730 777 776 818
rect 730 743 736 777
rect 770 743 776 777
rect 730 702 776 743
rect 730 668 736 702
rect 770 668 776 702
rect 730 626 776 668
rect 730 592 736 626
rect 770 592 776 626
rect 730 550 776 592
rect 730 516 736 550
rect 770 516 776 550
rect 730 474 776 516
rect 730 440 736 474
rect 770 440 776 474
rect 730 398 776 440
rect 730 364 736 398
rect 770 364 776 398
rect 886 1061 892 1095
rect 926 1092 935 1095
tri 935 1092 938 1095 nw
tri 1192 1092 1195 1095 ne
rect 1195 1092 1247 1095
tri 1247 1092 1250 1095 nw
tri 1504 1092 1507 1095 ne
rect 1507 1092 1559 1095
tri 1559 1092 1562 1095 nw
tri 1816 1092 1819 1095 ne
rect 1819 1092 1868 1095
rect 926 1061 932 1092
tri 932 1089 935 1092 nw
tri 1195 1089 1198 1092 ne
rect 886 1021 932 1061
rect 886 987 892 1021
rect 926 987 932 1021
rect 886 947 932 987
rect 886 913 892 947
rect 926 913 932 947
rect 886 873 932 913
rect 886 839 892 873
rect 926 839 932 873
rect 886 799 932 839
rect 886 765 892 799
rect 926 765 932 799
rect 886 725 932 765
rect 886 691 892 725
rect 926 691 932 725
rect 886 651 932 691
rect 886 617 892 651
rect 926 617 932 651
rect 886 577 932 617
rect 886 543 892 577
rect 926 543 932 577
rect 886 503 932 543
rect 886 469 892 503
rect 926 469 932 503
rect 886 429 932 469
rect 886 395 892 429
rect 926 395 932 429
tri 776 364 801 389 sw
rect 886 383 932 395
rect 1042 1077 1088 1089
rect 1042 1043 1048 1077
rect 1082 1043 1088 1077
rect 1042 1002 1088 1043
rect 1042 968 1048 1002
rect 1082 968 1088 1002
rect 1042 927 1088 968
rect 1042 893 1048 927
rect 1082 893 1088 927
rect 1042 852 1088 893
rect 1042 818 1048 852
rect 1082 818 1088 852
rect 1042 777 1088 818
rect 1042 743 1048 777
rect 1082 743 1088 777
rect 1042 702 1088 743
rect 1042 668 1048 702
rect 1082 668 1088 702
rect 1042 626 1088 668
rect 1042 592 1048 626
rect 1082 592 1088 626
rect 1042 550 1088 592
rect 1042 516 1048 550
rect 1082 516 1088 550
rect 1042 474 1088 516
rect 1042 440 1048 474
rect 1082 440 1088 474
rect 1042 398 1088 440
tri 1036 383 1042 389 se
rect 1042 383 1048 398
tri 1017 364 1036 383 se
rect 1036 364 1048 383
rect 1082 364 1088 398
rect 730 355 801 364
tri 801 355 810 364 sw
tri 1008 355 1017 364 se
rect 1017 355 1088 364
rect 730 328 1088 355
tri 620 274 626 280 sw
rect 730 276 736 328
rect 788 276 800 328
rect 852 322 1088 328
rect 852 288 1048 322
rect 1082 288 1088 322
rect 852 276 1088 288
rect 1198 1058 1204 1092
rect 1238 1058 1244 1092
tri 1244 1089 1247 1092 nw
tri 1507 1089 1510 1092 ne
rect 1198 1016 1244 1058
rect 1198 982 1204 1016
rect 1238 982 1244 1016
rect 1198 940 1244 982
rect 1198 906 1204 940
rect 1238 906 1244 940
rect 1198 864 1244 906
rect 1198 830 1204 864
rect 1238 830 1244 864
rect 1198 788 1244 830
rect 1198 754 1204 788
rect 1238 754 1244 788
rect 1198 711 1244 754
rect 1198 677 1204 711
rect 1238 677 1244 711
rect 1198 634 1244 677
rect 1198 600 1204 634
rect 1238 600 1244 634
rect 1198 557 1244 600
rect 1198 523 1204 557
rect 1238 523 1244 557
rect 1198 480 1244 523
rect 1198 446 1204 480
rect 1238 446 1244 480
rect 1198 403 1244 446
rect 1198 369 1204 403
rect 1238 369 1244 403
rect 1198 326 1244 369
rect 1198 292 1204 326
rect 1238 292 1244 326
rect 1198 280 1244 292
rect 1354 1077 1400 1089
rect 1354 1043 1360 1077
rect 1394 1043 1400 1077
rect 1354 1001 1400 1043
rect 1354 967 1360 1001
rect 1394 967 1400 1001
rect 1354 924 1400 967
rect 1354 890 1360 924
rect 1394 890 1400 924
rect 1354 847 1400 890
rect 1354 813 1360 847
rect 1394 813 1400 847
rect 1354 770 1400 813
rect 1354 736 1360 770
rect 1394 736 1400 770
rect 1354 693 1400 736
rect 1354 659 1360 693
rect 1394 659 1400 693
rect 1354 616 1400 659
rect 1354 582 1360 616
rect 1394 582 1400 616
rect 1354 539 1400 582
rect 1354 505 1360 539
rect 1394 505 1400 539
rect 1354 462 1400 505
rect 1354 428 1360 462
rect 1394 428 1400 462
rect 1354 385 1400 428
rect 1354 351 1360 385
rect 1394 351 1400 385
rect 1354 308 1400 351
tri 1350 276 1354 280 se
rect 1354 276 1360 308
tri 1348 274 1350 276 se
rect 1350 274 1360 276
rect 1394 274 1400 308
rect 1510 1058 1516 1092
rect 1550 1058 1556 1092
tri 1556 1089 1559 1092 nw
tri 1819 1089 1822 1092 ne
rect 1510 1016 1556 1058
rect 1510 982 1516 1016
rect 1550 982 1556 1016
rect 1510 940 1556 982
rect 1510 906 1516 940
rect 1550 906 1556 940
rect 1510 864 1556 906
rect 1510 830 1516 864
rect 1550 830 1556 864
rect 1510 788 1556 830
rect 1510 754 1516 788
rect 1550 754 1556 788
rect 1510 711 1556 754
rect 1510 677 1516 711
rect 1550 677 1556 711
rect 1510 634 1556 677
rect 1510 600 1516 634
rect 1550 600 1556 634
rect 1510 557 1556 600
rect 1510 523 1516 557
rect 1550 523 1556 557
rect 1510 480 1556 523
rect 1510 446 1516 480
rect 1550 446 1556 480
rect 1510 403 1556 446
rect 1510 369 1516 403
rect 1550 369 1556 403
rect 1510 326 1556 369
rect 1510 292 1516 326
rect 1550 292 1556 326
rect 1510 280 1556 292
rect 1666 1077 1712 1089
rect 1666 1043 1672 1077
rect 1706 1043 1712 1077
rect 1666 1001 1712 1043
rect 1666 967 1672 1001
rect 1706 967 1712 1001
rect 1666 924 1712 967
rect 1666 890 1672 924
rect 1706 890 1712 924
rect 1666 847 1712 890
rect 1666 813 1672 847
rect 1706 813 1712 847
rect 1666 770 1712 813
rect 1666 736 1672 770
rect 1706 736 1712 770
rect 1666 693 1712 736
rect 1666 659 1672 693
rect 1706 659 1712 693
rect 1666 616 1712 659
rect 1666 582 1672 616
rect 1706 582 1712 616
rect 1666 539 1712 582
rect 1666 505 1672 539
rect 1706 505 1712 539
rect 1666 462 1712 505
rect 1666 428 1672 462
rect 1706 428 1712 462
rect 1666 385 1712 428
rect 1666 351 1672 385
rect 1706 351 1712 385
rect 1666 308 1712 351
tri 1400 274 1406 280 sw
tri 1660 274 1666 280 se
rect 1666 274 1672 308
rect 1706 274 1712 308
rect 1822 1058 1828 1092
rect 1862 1058 1868 1092
rect 1822 1016 1868 1058
rect 1822 982 1828 1016
rect 1862 982 1868 1016
rect 1822 940 1868 982
rect 1822 906 1828 940
rect 1862 906 1868 940
rect 1822 864 1868 906
rect 1822 830 1828 864
rect 1862 830 1868 864
rect 1822 788 1868 830
rect 1822 754 1828 788
rect 1862 754 1868 788
rect 1822 711 1868 754
rect 1822 677 1828 711
rect 1862 677 1868 711
rect 1822 634 1868 677
rect 1822 600 1828 634
rect 1862 600 1868 634
rect 1822 557 1868 600
rect 1822 523 1828 557
rect 1862 523 1868 557
rect 1822 480 1868 523
rect 1822 446 1828 480
rect 1862 446 1868 480
rect 1822 403 1868 446
rect 1822 369 1828 403
rect 1862 369 1868 403
rect 1822 326 1868 369
rect 1822 292 1828 326
rect 1862 292 1868 326
rect 1822 280 1868 292
rect 1932 1168 2914 1203
rect 1932 1134 1938 1168
rect 1972 1134 2250 1168
rect 2284 1134 2562 1168
rect 2596 1134 2874 1168
rect 2908 1134 2914 1168
rect 1932 1123 2914 1134
rect 1932 1095 1984 1123
tri 1984 1095 2012 1123 nw
tri 2210 1095 2238 1123 ne
rect 2238 1095 2296 1123
tri 2296 1095 2324 1123 nw
tri 2522 1095 2550 1123 ne
rect 2550 1095 2608 1123
tri 2608 1095 2636 1123 nw
tri 2834 1095 2862 1123 ne
rect 2862 1095 2914 1123
rect 1932 1092 1981 1095
tri 1981 1092 1984 1095 nw
tri 2238 1092 2241 1095 ne
rect 2241 1092 2293 1095
tri 2293 1092 2296 1095 nw
tri 2550 1092 2553 1095 ne
rect 2553 1092 2602 1095
rect 1932 1058 1938 1092
rect 1972 1058 1978 1092
tri 1978 1089 1981 1092 nw
tri 2241 1089 2244 1092 ne
rect 1932 1016 1978 1058
rect 1932 982 1938 1016
rect 1972 982 1978 1016
rect 1932 940 1978 982
rect 1932 906 1938 940
rect 1972 906 1978 940
rect 1932 864 1978 906
rect 1932 830 1938 864
rect 1972 830 1978 864
rect 1932 788 1978 830
rect 1932 754 1938 788
rect 1972 754 1978 788
rect 1932 711 1978 754
rect 1932 677 1938 711
rect 1972 677 1978 711
rect 1932 634 1978 677
rect 1932 600 1938 634
rect 1972 600 1978 634
rect 1932 557 1978 600
rect 1932 523 1938 557
rect 1972 523 1978 557
rect 1932 480 1978 523
rect 1932 446 1938 480
rect 1972 446 1978 480
rect 1932 403 1978 446
rect 1932 369 1938 403
rect 1972 369 1978 403
rect 1932 326 1978 369
rect 1932 292 1938 326
rect 1972 292 1978 326
rect 1932 280 1978 292
rect 2088 1077 2134 1089
rect 2088 1043 2094 1077
rect 2128 1043 2134 1077
rect 2088 1001 2134 1043
rect 2088 967 2094 1001
rect 2128 967 2134 1001
rect 2088 924 2134 967
rect 2088 890 2094 924
rect 2128 890 2134 924
rect 2088 847 2134 890
rect 2088 813 2094 847
rect 2128 813 2134 847
rect 2088 770 2134 813
rect 2088 736 2094 770
rect 2128 736 2134 770
rect 2088 693 2134 736
rect 2088 659 2094 693
rect 2128 659 2134 693
rect 2088 616 2134 659
rect 2088 582 2094 616
rect 2128 582 2134 616
rect 2088 539 2134 582
rect 2088 505 2094 539
rect 2128 505 2134 539
rect 2088 462 2134 505
rect 2088 428 2094 462
rect 2128 428 2134 462
rect 2088 385 2134 428
rect 2088 351 2094 385
rect 2128 351 2134 385
rect 2088 308 2134 351
tri 1712 274 1718 280 sw
tri 2082 274 2088 280 se
rect 2088 274 2094 308
rect 2128 274 2134 308
rect 2244 1058 2250 1092
rect 2284 1058 2290 1092
tri 2290 1089 2293 1092 nw
tri 2553 1089 2556 1092 ne
rect 2244 1016 2290 1058
rect 2244 982 2250 1016
rect 2284 982 2290 1016
rect 2244 940 2290 982
rect 2244 906 2250 940
rect 2284 906 2290 940
rect 2244 864 2290 906
rect 2244 830 2250 864
rect 2284 830 2290 864
rect 2244 788 2290 830
rect 2244 754 2250 788
rect 2284 754 2290 788
rect 2244 711 2290 754
rect 2244 677 2250 711
rect 2284 677 2290 711
rect 2244 634 2290 677
rect 2244 600 2250 634
rect 2284 600 2290 634
rect 2244 557 2290 600
rect 2244 523 2250 557
rect 2284 523 2290 557
rect 2244 480 2290 523
rect 2244 446 2250 480
rect 2284 446 2290 480
rect 2244 403 2290 446
rect 2244 369 2250 403
rect 2284 369 2290 403
rect 2244 326 2290 369
rect 2244 292 2250 326
rect 2284 292 2290 326
rect 2244 280 2290 292
rect 2400 1077 2446 1089
rect 2400 1043 2406 1077
rect 2440 1043 2446 1077
rect 2400 1001 2446 1043
rect 2400 967 2406 1001
rect 2440 967 2446 1001
rect 2400 924 2446 967
rect 2400 890 2406 924
rect 2440 890 2446 924
rect 2400 847 2446 890
rect 2400 813 2406 847
rect 2440 813 2446 847
rect 2400 770 2446 813
rect 2400 736 2406 770
rect 2440 736 2446 770
rect 2400 693 2446 736
rect 2400 659 2406 693
rect 2440 659 2446 693
rect 2400 616 2446 659
rect 2400 582 2406 616
rect 2440 582 2446 616
rect 2400 539 2446 582
rect 2400 505 2406 539
rect 2440 505 2446 539
rect 2400 462 2446 505
rect 2400 428 2406 462
rect 2440 428 2446 462
rect 2400 385 2446 428
rect 2400 351 2406 385
rect 2440 351 2446 385
rect 2400 308 2446 351
tri 2134 274 2140 280 sw
tri 2394 274 2400 280 se
rect 2400 274 2406 308
rect 2440 274 2446 308
rect 2556 1058 2562 1092
rect 2596 1058 2602 1092
tri 2602 1089 2608 1095 nw
tri 2862 1089 2868 1095 ne
rect 2556 1016 2602 1058
rect 2556 982 2562 1016
rect 2596 982 2602 1016
rect 2556 940 2602 982
rect 2556 906 2562 940
rect 2596 906 2602 940
rect 2556 864 2602 906
rect 2556 830 2562 864
rect 2596 830 2602 864
rect 2556 788 2602 830
rect 2556 754 2562 788
rect 2596 754 2602 788
rect 2556 711 2602 754
rect 2556 677 2562 711
rect 2596 677 2602 711
rect 2556 634 2602 677
rect 2556 600 2562 634
rect 2596 600 2602 634
rect 2556 557 2602 600
rect 2556 523 2562 557
rect 2596 523 2602 557
rect 2556 480 2602 523
rect 2556 446 2562 480
rect 2596 446 2602 480
rect 2556 403 2602 446
rect 2556 369 2562 403
rect 2596 369 2602 403
rect 2556 326 2602 369
rect 2556 292 2562 326
rect 2596 292 2602 326
rect 2556 280 2602 292
rect 2709 1077 2761 1089
rect 2709 1043 2718 1077
rect 2752 1043 2761 1077
rect 2709 1002 2761 1043
rect 2709 982 2718 1002
rect 2752 982 2761 1002
rect 2709 927 2761 930
rect 2709 918 2718 927
rect 2752 918 2761 927
rect 2709 852 2761 866
rect 2709 818 2718 852
rect 2752 818 2761 852
rect 2709 777 2761 818
rect 2709 743 2718 777
rect 2752 743 2761 777
rect 2709 702 2761 743
rect 2709 668 2718 702
rect 2752 668 2761 702
rect 2709 627 2761 668
rect 2709 593 2718 627
rect 2752 593 2761 627
rect 2709 552 2761 593
rect 2709 518 2718 552
rect 2752 518 2761 552
rect 2709 477 2761 518
rect 2709 443 2718 477
rect 2752 443 2761 477
rect 2709 402 2761 443
rect 2709 368 2718 402
rect 2752 368 2761 402
rect 2868 1061 2874 1095
rect 2908 1061 2914 1095
rect 2868 1022 2914 1061
rect 2868 988 2874 1022
rect 2908 988 2914 1022
rect 2868 949 2914 988
rect 2868 915 2874 949
rect 2908 915 2914 949
rect 2868 876 2914 915
rect 2868 842 2874 876
rect 2908 842 2914 876
rect 2868 803 2914 842
rect 2868 769 2874 803
rect 2908 769 2914 803
rect 2868 730 2914 769
rect 2868 696 2874 730
rect 2908 696 2914 730
rect 2868 657 2914 696
rect 2868 623 2874 657
rect 2908 623 2914 657
rect 2868 583 2914 623
rect 2868 549 2874 583
rect 2908 549 2914 583
rect 2868 509 2914 549
rect 2868 475 2874 509
rect 2908 475 2914 509
rect 2868 435 2914 475
rect 2868 401 2874 435
rect 2908 401 2914 435
tri 2761 368 2786 393 sw
rect 2868 389 2914 401
rect 3021 1077 3073 1089
rect 3021 1043 3030 1077
rect 3064 1043 3073 1077
rect 3021 1002 3073 1043
rect 3021 982 3030 1002
rect 3064 982 3073 1002
rect 3021 927 3073 930
rect 3021 918 3030 927
rect 3064 918 3073 927
rect 3021 852 3073 866
rect 3021 818 3030 852
rect 3064 818 3073 852
rect 3021 777 3073 818
rect 3021 743 3030 777
rect 3064 743 3073 777
rect 3021 702 3073 743
rect 3021 668 3030 702
rect 3064 668 3073 702
rect 3021 627 3073 668
rect 3021 593 3030 627
rect 3064 593 3073 627
rect 3021 552 3073 593
rect 3021 518 3030 552
rect 3064 518 3073 552
rect 3021 477 3073 518
rect 3021 443 3030 477
rect 3064 443 3073 477
rect 3021 402 3073 443
tri 3017 389 3021 393 se
rect 3021 389 3030 402
tri 2996 368 3017 389 se
rect 3017 368 3030 389
rect 3064 368 3073 402
rect 2709 359 2786 368
tri 2786 359 2795 368 sw
tri 2987 359 2996 368 se
rect 2996 359 3073 368
rect 2709 326 3073 359
rect 2709 292 2718 326
rect 2752 292 3030 326
rect 3064 292 3073 326
rect 2709 280 3073 292
tri 540 246 568 274 se
rect 568 246 626 274
tri 626 246 654 274 sw
tri 1320 246 1348 274 se
rect 1348 246 1406 274
tri 1406 246 1434 274 sw
tri 1632 246 1660 274 se
rect 1660 246 1718 274
tri 1718 246 1746 274 sw
tri 2054 246 2082 274 se
rect 2082 246 2140 274
tri 2140 246 2168 274 sw
tri 2366 246 2394 274 se
rect 2394 246 2446 274
tri 2446 246 2480 280 sw
rect 536 243 3891 246
rect 536 238 3705 243
rect 536 231 1047 238
rect 536 197 580 231
rect 614 197 1047 231
rect 536 186 1047 197
rect 1099 186 1111 238
rect 1163 231 3705 238
rect 1163 197 1360 231
rect 1394 197 1672 231
rect 1706 197 2094 231
rect 2128 197 2406 231
rect 2440 197 3705 231
rect 1163 191 3705 197
rect 3757 191 3769 243
rect 3821 191 3833 243
rect 3885 191 3891 243
rect 1163 186 3891 191
rect 536 125 3891 186
rect 536 91 616 125
rect 650 91 689 125
rect 723 91 762 125
rect 796 91 835 125
rect 869 91 908 125
rect 942 91 981 125
rect 1015 123 1054 125
rect 1088 123 1128 125
rect 1162 123 1202 125
rect 1015 91 1047 123
rect 536 71 1047 91
rect 1099 71 1111 123
rect 1163 91 1202 123
rect 1236 91 1276 125
rect 1310 91 1350 125
rect 1384 91 1424 125
rect 1458 91 1498 125
rect 1532 91 1572 125
rect 1606 91 1646 125
rect 1680 91 1720 125
rect 1754 91 1794 125
rect 1828 91 1868 125
rect 1902 91 1942 125
rect 1976 91 2016 125
rect 2050 91 2090 125
rect 2124 91 2164 125
rect 2198 91 2238 125
rect 2272 91 2312 125
rect 2346 91 2386 125
rect 2420 91 2460 125
rect 2494 91 2534 125
rect 2568 91 2608 125
rect 2642 91 2682 125
rect 2716 91 2756 125
rect 2790 91 2830 125
rect 2864 91 2904 125
rect 2938 91 2978 125
rect 3012 117 3891 125
rect 3012 91 3705 117
rect 1163 71 3705 91
rect 536 65 3705 71
rect 3757 65 3769 117
rect 3821 65 3833 117
rect 3885 65 3891 117
rect 536 -169 3891 65
<< via1 >>
rect 913 3089 922 3121
rect 922 3089 956 3121
rect 956 3089 965 3121
rect 913 3069 965 3089
rect 913 3045 965 3057
rect 913 3011 922 3045
rect 922 3011 956 3045
rect 956 3011 965 3045
rect 913 3005 965 3011
rect 1445 3115 1497 3148
rect 1445 3096 1454 3115
rect 1454 3096 1488 3115
rect 1488 3096 1497 3115
rect 1445 3081 1454 3084
rect 1454 3081 1488 3084
rect 1488 3081 1497 3084
rect 1445 3040 1497 3081
rect 1445 3032 1454 3040
rect 1454 3032 1488 3040
rect 1488 3032 1497 3040
rect 2492 3115 2544 3148
rect 2492 3096 2500 3115
rect 2500 3096 2534 3115
rect 2534 3096 2544 3115
rect 2492 3081 2500 3084
rect 2500 3081 2534 3084
rect 2534 3081 2544 3084
rect 2492 3040 2544 3081
rect 2492 3032 2500 3040
rect 2500 3032 2534 3040
rect 2534 3032 2544 3040
rect 2757 3115 2809 3148
rect 2757 3096 2766 3115
rect 2766 3096 2800 3115
rect 2800 3096 2809 3115
rect 2757 3081 2766 3084
rect 2766 3081 2800 3084
rect 2800 3081 2809 3084
rect 2757 3040 2809 3081
rect 2757 3032 2766 3040
rect 2766 3032 2800 3040
rect 2800 3032 2809 3040
rect 3482 2929 3500 2950
rect 3500 2929 3534 2950
rect 3482 2898 3534 2929
rect 3546 2898 3598 2950
rect 633 2828 685 2832
rect 633 2794 637 2828
rect 637 2794 671 2828
rect 671 2794 685 2828
rect 633 2780 685 2794
rect 697 2828 749 2832
rect 697 2794 709 2828
rect 709 2794 743 2828
rect 743 2794 749 2828
rect 697 2780 749 2794
rect 1328 2828 1380 2837
rect 1392 2828 1444 2837
rect 1328 2794 1368 2828
rect 1368 2794 1380 2828
rect 1392 2794 1402 2828
rect 1402 2794 1444 2828
rect 1328 2785 1380 2794
rect 1392 2785 1444 2794
rect 1774 2828 1826 2837
rect 1774 2794 1803 2828
rect 1803 2794 1826 2828
rect 1774 2785 1826 2794
rect 1838 2828 1890 2837
rect 1838 2794 1850 2828
rect 1850 2794 1884 2828
rect 1884 2794 1890 2828
rect 1838 2785 1890 2794
rect 2120 2828 2172 2837
rect 2184 2828 2236 2837
rect 2120 2794 2126 2828
rect 2126 2794 2172 2828
rect 2184 2794 2215 2828
rect 2215 2794 2236 2828
rect 2120 2785 2172 2794
rect 2184 2785 2236 2794
rect 2510 2828 2562 2837
rect 2510 2794 2533 2828
rect 2533 2794 2562 2828
rect 2510 2785 2562 2794
rect 2574 2828 2626 2837
rect 2574 2794 2586 2828
rect 2586 2794 2620 2828
rect 2620 2794 2626 2828
rect 2574 2785 2626 2794
rect 2785 2828 2837 2837
rect 2785 2794 2791 2828
rect 2791 2794 2825 2828
rect 2825 2794 2837 2828
rect 2785 2785 2837 2794
rect 2849 2828 2901 2837
rect 2849 2794 2863 2828
rect 2863 2794 2897 2828
rect 2897 2794 2901 2828
rect 2849 2785 2901 2794
rect 3007 2828 3059 2837
rect 3071 2828 3123 2837
rect 3007 2794 3013 2828
rect 3013 2794 3051 2828
rect 3051 2794 3059 2828
rect 3071 2794 3085 2828
rect 3085 2794 3123 2828
rect 3007 2785 3059 2794
rect 3071 2785 3123 2794
rect 3324 2828 3376 2837
rect 3388 2828 3440 2837
rect 3324 2794 3362 2828
rect 3362 2794 3376 2828
rect 3388 2794 3396 2828
rect 3396 2794 3435 2828
rect 3435 2794 3440 2828
rect 3324 2785 3376 2794
rect 3388 2785 3440 2794
rect 1444 2676 1496 2728
rect 1508 2676 1560 2728
rect 2120 2676 2172 2728
rect 2184 2676 2236 2728
rect 595 2590 647 2642
rect 1774 2596 1826 2648
rect 1838 2596 1890 2648
rect 595 2526 647 2578
rect 2392 2516 2444 2568
rect 2456 2516 2508 2568
rect 3083 2516 3135 2568
rect 3147 2516 3199 2568
rect 1047 2344 1163 2460
rect 1930 2468 1982 2477
rect 1930 2434 1944 2468
rect 1944 2434 1978 2468
rect 1978 2434 1982 2468
rect 1930 2425 1982 2434
rect 1994 2468 2046 2477
rect 1994 2434 2028 2468
rect 2028 2434 2046 2468
rect 1994 2425 2046 2434
rect 3704 2434 3714 2468
rect 3714 2434 3748 2468
rect 3748 2434 3756 2468
rect 3704 2416 3756 2434
rect 3768 2416 3820 2468
rect 3832 2457 3884 2468
rect 3832 2423 3864 2457
rect 3864 2423 3884 2457
rect 3832 2416 3884 2423
rect 2580 2321 2632 2373
rect 1252 2217 1304 2226
rect 1316 2217 1368 2226
rect 1252 2183 1283 2217
rect 1283 2183 1304 2217
rect 1316 2183 1317 2217
rect 1317 2183 1356 2217
rect 1356 2183 1368 2217
rect 1252 2174 1304 2183
rect 1316 2174 1368 2183
rect 1514 2172 1523 2204
rect 1523 2172 1557 2204
rect 1557 2172 1566 2204
rect 1514 2152 1566 2172
rect 1514 2118 1566 2140
rect 1514 2088 1523 2118
rect 1523 2088 1557 2118
rect 1557 2088 1566 2118
rect 2580 2257 2632 2309
rect 3704 2334 3756 2386
rect 3768 2334 3820 2386
rect 3832 2382 3884 2386
rect 3832 2348 3864 2382
rect 3864 2348 3884 2382
rect 3832 2334 3884 2348
rect 2392 2232 2444 2239
rect 2392 2198 2396 2232
rect 2396 2198 2430 2232
rect 2430 2198 2444 2232
rect 2392 2187 2444 2198
rect 2456 2232 2508 2239
rect 2456 2198 2468 2232
rect 2468 2198 2502 2232
rect 2502 2198 2508 2232
rect 2456 2187 2508 2198
rect 2392 2076 2444 2085
rect 2392 2042 2396 2076
rect 2396 2042 2430 2076
rect 2430 2042 2444 2076
rect 2392 2033 2444 2042
rect 2456 2076 2508 2085
rect 2456 2042 2468 2076
rect 2468 2042 2502 2076
rect 2502 2042 2508 2076
rect 2456 2033 2508 2042
rect 3482 2312 3534 2321
rect 3482 2278 3486 2312
rect 3486 2278 3520 2312
rect 3520 2278 3534 2312
rect 3482 2269 3534 2278
rect 3546 2312 3598 2321
rect 3546 2278 3562 2312
rect 3562 2278 3596 2312
rect 3596 2278 3598 2312
rect 3546 2269 3598 2278
rect 3704 2252 3756 2304
rect 3768 2252 3820 2304
rect 3832 2272 3864 2304
rect 3864 2272 3884 2304
rect 3832 2252 3884 2272
rect 3704 2170 3756 2222
rect 3768 2170 3820 2222
rect 3832 2196 3864 2222
rect 3864 2196 3884 2222
rect 3832 2170 3884 2196
rect 3704 2122 3714 2140
rect 3714 2122 3748 2140
rect 3748 2122 3756 2140
rect 3704 2088 3756 2122
rect 3768 2088 3820 2140
rect 3832 2120 3864 2140
rect 3864 2120 3884 2140
rect 3832 2088 3884 2120
rect 3482 2000 3534 2009
rect 3482 1966 3486 2000
rect 3486 1966 3520 2000
rect 3520 1966 3534 2000
rect 3482 1957 3534 1966
rect 3546 2000 3598 2009
rect 3546 1966 3562 2000
rect 3562 1966 3596 2000
rect 3596 1966 3598 2000
rect 3546 1957 3598 1966
rect 1252 1880 1304 1932
rect 1316 1880 1368 1932
rect 1930 1844 1982 1856
rect 1930 1810 1944 1844
rect 1944 1810 1978 1844
rect 1978 1810 1982 1844
rect 1930 1804 1982 1810
rect 1994 1844 2046 1856
rect 1994 1810 2028 1844
rect 2028 1810 2046 1844
rect 1994 1804 2046 1810
rect 879 1724 931 1776
rect 943 1724 995 1776
rect 2666 1644 2718 1696
rect 2730 1644 2782 1696
rect 1346 1496 1398 1548
rect 1410 1496 1462 1548
rect 2392 1496 2444 1548
rect 2456 1496 2508 1548
rect 2847 1496 2899 1548
rect 2911 1496 2963 1548
rect 2586 1416 2638 1468
rect 2650 1416 2702 1468
rect 558 1283 610 1292
rect 622 1283 674 1292
rect 558 1249 607 1283
rect 607 1249 610 1283
rect 622 1249 641 1283
rect 641 1249 674 1283
rect 558 1240 610 1249
rect 622 1240 674 1249
rect 840 1283 892 1292
rect 904 1283 956 1292
rect 840 1249 842 1283
rect 842 1249 889 1283
rect 889 1249 892 1283
rect 904 1249 923 1283
rect 923 1249 956 1283
rect 840 1240 892 1249
rect 904 1240 956 1249
rect 1270 1283 1322 1292
rect 1270 1249 1276 1283
rect 1276 1249 1310 1283
rect 1310 1249 1322 1283
rect 1270 1240 1322 1249
rect 1334 1283 1386 1292
rect 2414 1283 2466 1292
rect 1334 1249 1350 1283
rect 1350 1249 1384 1283
rect 1384 1249 1386 1283
rect 2414 1249 2444 1283
rect 2444 1249 2466 1283
rect 1334 1240 1386 1249
rect 2414 1240 2466 1249
rect 2478 1283 2530 1292
rect 2478 1249 2490 1283
rect 2490 1249 2524 1283
rect 2524 1249 2530 1283
rect 2478 1240 2530 1249
rect 2666 1283 2718 1292
rect 2730 1283 2782 1292
rect 2666 1249 2671 1283
rect 2671 1249 2715 1283
rect 2715 1249 2718 1283
rect 2730 1249 2749 1283
rect 2749 1249 2782 1283
rect 2666 1240 2718 1249
rect 2730 1240 2782 1249
rect 736 322 788 328
rect 736 288 770 322
rect 770 288 788 322
rect 736 276 788 288
rect 800 276 852 328
rect 2709 968 2718 982
rect 2718 968 2752 982
rect 2752 968 2761 982
rect 2709 930 2761 968
rect 2709 893 2718 918
rect 2718 893 2752 918
rect 2752 893 2761 918
rect 2709 866 2761 893
rect 3021 968 3030 982
rect 3030 968 3064 982
rect 3064 968 3073 982
rect 3021 930 3073 968
rect 3021 893 3030 918
rect 3030 893 3064 918
rect 3064 893 3073 918
rect 3021 866 3073 893
rect 1047 186 1099 238
rect 1111 186 1163 238
rect 3705 191 3757 243
rect 3769 191 3821 243
rect 3833 191 3885 243
rect 1047 91 1054 123
rect 1054 91 1088 123
rect 1088 91 1099 123
rect 1047 71 1099 91
rect 1111 91 1128 123
rect 1128 91 1162 123
rect 1162 91 1163 123
rect 1111 71 1163 91
rect 3705 65 3757 117
rect 3769 65 3821 117
rect 3833 65 3885 117
<< metal2 >>
rect 1445 3148 3340 3154
rect 913 3121 965 3127
rect 913 3057 965 3069
rect 1497 3096 2492 3148
rect 2544 3096 2757 3148
rect 2809 3096 3340 3148
rect 1445 3084 3340 3096
rect 1497 3032 2492 3084
rect 2544 3032 2757 3084
rect 2809 3048 3340 3084
tri 3340 3048 3446 3154 sw
rect 2809 3032 3446 3048
rect 1445 3026 3446 3032
tri 882 2898 913 2929 se
rect 913 2907 965 3005
tri 1890 2992 1924 3026 ne
rect 913 2898 956 2907
tri 956 2898 965 2907 nw
tri 839 2855 882 2898 se
rect 882 2855 913 2898
tri 913 2855 956 2898 nw
tri 821 2837 839 2855 se
rect 839 2837 895 2855
tri 895 2837 913 2855 nw
tri 816 2832 821 2837 se
rect 821 2832 890 2837
tri 890 2832 895 2837 nw
rect 625 2780 633 2832
rect 685 2780 697 2832
rect 749 2785 843 2832
tri 843 2785 890 2832 nw
rect 1322 2785 1328 2837
rect 1380 2785 1392 2837
rect 1444 2785 1450 2837
rect 1768 2785 1774 2837
rect 1826 2785 1838 2837
rect 1890 2785 1896 2837
rect 749 2780 838 2785
tri 838 2780 843 2785 nw
tri 696 2746 730 2780 ne
rect 595 2642 647 2648
rect 595 2578 647 2590
tri 561 1292 595 1326 se
rect 595 1292 647 2526
tri 647 1292 680 1325 sw
rect 552 1240 558 1292
rect 610 1240 622 1292
rect 674 1240 680 1292
rect 730 328 782 2780
tri 782 2746 816 2780 nw
rect 1047 2460 1163 2466
rect 872 1724 879 1776
rect 931 1724 943 1776
rect 995 1724 1001 1776
rect 872 1696 930 1724
tri 930 1696 958 1724 nw
tri 838 1292 872 1326 se
rect 872 1292 924 1696
tri 924 1690 930 1696 nw
tri 924 1292 958 1326 sw
rect 834 1240 840 1292
rect 892 1240 904 1292
rect 956 1240 962 1292
tri 782 328 816 362 sw
rect 730 276 736 328
rect 788 276 800 328
rect 852 276 858 328
rect 1047 238 1163 2344
tri 1319 2257 1322 2260 se
rect 1322 2257 1374 2785
tri 1374 2751 1408 2785 nw
rect 1438 2676 1444 2728
rect 1496 2676 1508 2728
rect 1560 2676 1566 2728
tri 1480 2648 1508 2676 ne
rect 1508 2648 1566 2676
tri 1508 2642 1514 2648 ne
tri 1314 2252 1319 2257 se
rect 1319 2252 1374 2257
tri 1301 2239 1314 2252 se
rect 1314 2239 1374 2252
tri 1288 2226 1301 2239 se
rect 1301 2226 1374 2239
rect 1246 2174 1252 2226
rect 1304 2174 1316 2226
rect 1368 2174 1374 2226
tri 1288 2152 1310 2174 ne
rect 1310 2152 1374 2174
tri 1310 2140 1322 2152 ne
tri 1313 1957 1322 1966 se
rect 1322 1957 1374 2152
tri 1288 1932 1313 1957 se
rect 1313 1932 1374 1957
rect 1246 1880 1252 1932
rect 1304 1880 1316 1932
rect 1368 1880 1374 1932
rect 1514 2204 1566 2648
rect 1768 2648 1896 2785
rect 1768 2596 1774 2648
rect 1826 2596 1838 2648
rect 1890 2596 1896 2648
rect 1514 2140 1566 2152
rect 1340 1496 1346 1548
rect 1398 1496 1410 1548
rect 1462 1496 1468 1548
rect 1340 1468 1398 1496
tri 1398 1468 1426 1496 nw
tri 1306 1292 1340 1326 se
rect 1340 1292 1392 1468
tri 1392 1462 1398 1468 nw
rect 1264 1240 1270 1292
rect 1322 1240 1334 1292
rect 1386 1240 1392 1292
rect 1514 1071 1566 2088
rect 1924 2477 2052 3026
tri 2052 2992 2086 3026 nw
tri 3286 2994 3318 3026 ne
rect 3318 2837 3446 3026
rect 2114 2785 2120 2837
rect 2172 2785 2184 2837
rect 2236 2785 2242 2837
rect 2504 2785 2510 2837
rect 2562 2785 2574 2837
rect 2626 2785 2632 2837
rect 2779 2785 2785 2837
rect 2837 2785 2849 2837
rect 2901 2785 2907 2837
rect 3001 2785 3007 2837
rect 3059 2785 3071 2837
rect 3123 2785 3129 2837
rect 3318 2785 3324 2837
rect 3376 2785 3388 2837
rect 3440 2785 3446 2837
rect 3476 2950 3604 2974
rect 3476 2898 3482 2950
rect 3534 2898 3546 2950
rect 3598 2898 3604 2950
rect 2114 2728 2242 2785
tri 2546 2751 2580 2785 ne
rect 2114 2676 2120 2728
rect 2172 2676 2184 2728
rect 2236 2676 2242 2728
rect 2386 2516 2392 2568
rect 2444 2516 2456 2568
rect 2508 2516 2514 2568
tri 2428 2482 2462 2516 ne
rect 1924 2425 1930 2477
rect 1982 2425 1994 2477
rect 2046 2425 2052 2477
rect 1924 1856 2052 2425
tri 2446 2257 2462 2273 se
rect 2462 2257 2514 2516
tri 2441 2252 2446 2257 se
rect 2446 2252 2514 2257
tri 2428 2239 2441 2252 se
rect 2441 2239 2514 2252
rect 2386 2187 2392 2239
rect 2444 2187 2456 2239
rect 2508 2187 2514 2239
rect 2580 2373 2632 2785
tri 2807 2751 2841 2785 ne
rect 2580 2309 2632 2321
rect 2386 2033 2392 2085
rect 2444 2033 2456 2085
rect 2508 2033 2514 2085
tri 2428 2009 2452 2033 ne
rect 2452 2009 2514 2033
tri 2452 1999 2462 2009 ne
rect 1924 1804 1930 1856
rect 1982 1804 1994 1856
rect 2046 1804 2052 1856
tri 2428 1548 2462 1582 se
rect 2462 1548 2514 2009
rect 2386 1496 2392 1548
rect 2444 1496 2456 1548
rect 2508 1496 2514 1548
tri 2428 1468 2456 1496 ne
rect 2456 1468 2514 1496
tri 2456 1462 2462 1468 ne
tri 2428 1292 2462 1326 se
rect 2462 1292 2514 1468
rect 2580 1496 2632 2257
rect 2660 1644 2666 1696
rect 2718 1644 2730 1696
rect 2782 1644 2788 1696
tri 2702 1610 2736 1644 ne
tri 2632 1496 2638 1502 sw
rect 2580 1468 2638 1496
tri 2638 1468 2666 1496 sw
rect 2580 1416 2586 1468
rect 2638 1416 2650 1468
rect 2702 1416 2708 1468
tri 2724 1314 2736 1326 se
rect 2736 1314 2788 1644
rect 2841 1548 2893 2785
tri 2893 2771 2907 2785 nw
tri 3043 2771 3057 2785 ne
rect 3057 2771 3129 2785
tri 3057 2751 3077 2771 ne
rect 3077 2568 3129 2771
tri 3129 2568 3163 2602 sw
rect 3077 2516 3083 2568
rect 3135 2516 3147 2568
rect 3199 2516 3205 2568
rect 3476 2321 3604 2898
rect 3476 2269 3482 2321
rect 3534 2269 3546 2321
rect 3598 2269 3604 2321
rect 3476 2009 3604 2269
rect 3476 1957 3482 2009
rect 3534 1957 3546 2009
rect 3598 1957 3604 2009
rect 3699 2468 3891 2474
rect 3699 2416 3704 2468
rect 3756 2416 3768 2468
rect 3820 2416 3832 2468
rect 3884 2416 3891 2468
rect 3699 2386 3891 2416
rect 3699 2334 3704 2386
rect 3756 2334 3768 2386
rect 3820 2334 3832 2386
rect 3884 2334 3891 2386
rect 3699 2304 3891 2334
rect 3699 2252 3704 2304
rect 3756 2252 3768 2304
rect 3820 2252 3832 2304
rect 3884 2252 3891 2304
rect 3699 2222 3891 2252
rect 3699 2170 3704 2222
rect 3756 2170 3768 2222
rect 3820 2170 3832 2222
rect 3884 2170 3891 2222
rect 3699 2140 3891 2170
rect 3699 2088 3704 2140
rect 3756 2088 3768 2140
rect 3820 2088 3832 2140
rect 3884 2088 3891 2140
tri 2893 1548 2927 1582 sw
rect 2841 1496 2847 1548
rect 2899 1496 2911 1548
rect 2963 1496 2969 1548
tri 2514 1292 2536 1314 sw
tri 2702 1292 2724 1314 se
rect 2724 1292 2788 1314
rect 2408 1240 2414 1292
rect 2466 1240 2478 1292
rect 2530 1240 2536 1292
rect 2660 1240 2666 1292
rect 2718 1240 2730 1292
rect 2782 1240 2788 1292
tri 1566 1071 1588 1093 sw
tri 1514 997 1588 1071 ne
tri 1588 1010 1649 1071 sw
rect 1588 997 1649 1010
tri 1588 982 1603 997 ne
rect 1603 988 1649 997
tri 1649 988 1671 1010 sw
rect 1603 982 3073 988
tri 1603 936 1649 982 ne
rect 1649 936 2709 982
tri 2675 930 2681 936 ne
rect 2681 930 2709 936
rect 2761 936 3021 982
rect 2761 930 2789 936
tri 2789 930 2795 936 nw
tri 2987 930 2993 936 ne
rect 2993 930 3021 936
tri 2681 918 2693 930 ne
rect 2693 918 2777 930
tri 2777 918 2789 930 nw
tri 2993 918 3005 930 ne
rect 3005 918 3073 930
tri 2693 902 2709 918 ne
tri 2761 902 2777 918 nw
tri 3005 902 3021 918 ne
rect 2709 860 2761 866
rect 3021 860 3073 866
rect 1099 186 1111 238
rect 1047 123 1163 186
rect 1099 71 1111 123
rect 1047 65 1163 71
rect 3699 243 3891 2088
rect 3699 191 3705 243
rect 3757 191 3769 243
rect 3821 191 3833 243
rect 3885 191 3891 243
rect 3699 117 3891 191
rect 3699 65 3705 117
rect 3757 65 3769 117
rect 3821 65 3833 117
rect 3885 65 3891 117
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_0
timestamp 1704896540
transform 0 1 1752 1 0 1855
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_1
timestamp 1704896540
transform 0 1 1752 1 0 2011
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_2
timestamp 1704896540
transform 0 1 1752 -1 0 2267
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808528  sky130_fd_pr__nfet_01v8__example_55959141808528_3
timestamp 1704896540
transform 0 1 1752 -1 0 2423
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808533  sky130_fd_pr__nfet_01v8__example_55959141808533_0
timestamp 1704896540
transform -1 0 725 0 1 201
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808550  sky130_fd_pr__nfet_01v8__example_55959141808550_0
timestamp 1704896540
transform 1 0 2607 0 1 201
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808550  sky130_fd_pr__nfet_01v8__example_55959141808550_1
timestamp 1704896540
transform 0 -1 3748 1 0 2011
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808550  sky130_fd_pr__nfet_01v8__example_55959141808550_2
timestamp 1704896540
transform -1 0 1193 0 1 201
box -1 0 413 1
use sky130_fd_pr__nfet_01v8__example_55959141808600  sky130_fd_pr__nfet_01v8__example_55959141808600_0
timestamp 1704896540
transform 0 1 1175 1 0 2072
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808607  sky130_fd_pr__nfet_01v8__example_55959141808607_0
timestamp 1704896540
transform 1 0 1983 0 1 201
box -1 0 569 1
use sky130_fd_pr__nfet_01v8__example_55959141808607  sky130_fd_pr__nfet_01v8__example_55959141808607_1
timestamp 1704896540
transform -1 0 1817 0 1 201
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_0
timestamp 1704896540
transform -1 0 1911 0 -1 3876
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_1
timestamp 1704896540
transform -1 0 1599 0 -1 3876
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_2
timestamp 1704896540
transform 1 0 2077 0 -1 3876
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808189  sky130_fd_pr__pfet_01v8__example_55959141808189_3
timestamp 1704896540
transform 1 0 2389 0 -1 3876
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_0
timestamp 1704896540
transform 1 0 1077 0 -1 3176
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_1
timestamp 1704896540
transform -1 0 755 0 -1 3176
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_2
timestamp 1704896540
transform -1 0 911 0 -1 3176
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808537  sky130_fd_pr__pfet_01v8__example_55959141808537_0
timestamp 1704896540
transform 1 0 3233 0 -1 3876
box -1 0 725 1
use sky130_fd_pr__pfet_01v8__example_55959141808548  sky130_fd_pr__pfet_01v8__example_55959141808548_0
timestamp 1704896540
transform -1 0 2911 0 -1 3876
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808548  sky130_fd_pr__pfet_01v8__example_55959141808548_1
timestamp 1704896540
transform -1 0 3067 0 -1 3876
box -1 0 101 1
<< labels >>
flabel metal2 s 3497 2028 3567 2095 3 FreeSans 200 0 0 0 OUT
port 1 nsew
flabel metal2 s 1940 2676 2035 2758 3 FreeSans 200 0 0 0 OUT_B
port 2 nsew
flabel metal1 s 3675 2686 3805 2723 3 FreeSans 200 0 0 0 MODE_NORMAL_N
port 3 nsew
flabel metal1 s 710 1653 851 1689 3 FreeSans 200 0 0 0 IN_VCCHIB
port 4 nsew
flabel metal1 s 696 1738 851 1771 3 FreeSans 200 0 0 0 INB_VCCHIB
port 5 nsew
flabel metal1 s 695 1431 865 1462 3 FreeSans 200 0 0 0 IN_VDDIO
port 6 nsew
flabel metal1 s 3678 2605 3804 2639 3 FreeSans 200 0 0 0 MODE_VCCHIB_N
port 7 nsew
flabel metal1 s 3689 2525 3799 2561 3 FreeSans 200 0 0 0 MODE_NORMAL
port 8 nsew
flabel metal1 s 1621 1510 1785 1539 3 FreeSans 200 0 0 0 MODE_VCCHIB
port 9 nsew
flabel metal1 s 682 3811 1004 4027 3 FreeSans 200 0 0 0 VDDIO_Q
port 10 nsew
flabel metal1 s 599 86 824 210 3 FreeSans 200 0 0 0 VSSD
port 11 nsew
<< properties >>
string GDS_END 17088434
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 16989590
<< end >>
