magic
tech sky130A
timestamp 1704896540
<< properties >>
string GDS_END 58008230
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 58007842
<< end >>
