magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 -36 236 3036
<< pdiff >>
rect 0 2970 60 3000
rect 0 2936 11 2970
rect 45 2936 60 2970
rect 0 2902 60 2936
rect 0 2868 11 2902
rect 45 2868 60 2902
rect 0 2834 60 2868
rect 0 2800 11 2834
rect 45 2800 60 2834
rect 0 2766 60 2800
rect 0 2732 11 2766
rect 45 2732 60 2766
rect 0 2698 60 2732
rect 0 2664 11 2698
rect 45 2664 60 2698
rect 0 2630 60 2664
rect 0 2596 11 2630
rect 45 2596 60 2630
rect 0 2562 60 2596
rect 0 2528 11 2562
rect 45 2528 60 2562
rect 0 2494 60 2528
rect 0 2460 11 2494
rect 45 2460 60 2494
rect 0 2426 60 2460
rect 0 2392 11 2426
rect 45 2392 60 2426
rect 0 2358 60 2392
rect 0 2324 11 2358
rect 45 2324 60 2358
rect 0 2290 60 2324
rect 0 2256 11 2290
rect 45 2256 60 2290
rect 0 2222 60 2256
rect 0 2188 11 2222
rect 45 2188 60 2222
rect 0 2154 60 2188
rect 0 2120 11 2154
rect 45 2120 60 2154
rect 0 2086 60 2120
rect 0 2052 11 2086
rect 45 2052 60 2086
rect 0 2018 60 2052
rect 0 1984 11 2018
rect 45 1984 60 2018
rect 0 1950 60 1984
rect 0 1916 11 1950
rect 45 1916 60 1950
rect 0 1882 60 1916
rect 0 1848 11 1882
rect 45 1848 60 1882
rect 0 1814 60 1848
rect 0 1780 11 1814
rect 45 1780 60 1814
rect 0 1746 60 1780
rect 0 1712 11 1746
rect 45 1712 60 1746
rect 0 1678 60 1712
rect 0 1644 11 1678
rect 45 1644 60 1678
rect 0 1610 60 1644
rect 0 1576 11 1610
rect 45 1576 60 1610
rect 0 1542 60 1576
rect 0 1508 11 1542
rect 45 1508 60 1542
rect 0 1474 60 1508
rect 0 1440 11 1474
rect 45 1440 60 1474
rect 0 1406 60 1440
rect 0 1372 11 1406
rect 45 1372 60 1406
rect 0 1338 60 1372
rect 0 1304 11 1338
rect 45 1304 60 1338
rect 0 1270 60 1304
rect 0 1236 11 1270
rect 45 1236 60 1270
rect 0 1202 60 1236
rect 0 1168 11 1202
rect 45 1168 60 1202
rect 0 1134 60 1168
rect 0 1100 11 1134
rect 45 1100 60 1134
rect 0 1066 60 1100
rect 0 1032 11 1066
rect 45 1032 60 1066
rect 0 998 60 1032
rect 0 964 11 998
rect 45 964 60 998
rect 0 930 60 964
rect 0 896 11 930
rect 45 896 60 930
rect 0 862 60 896
rect 0 828 11 862
rect 45 828 60 862
rect 0 794 60 828
rect 0 760 11 794
rect 45 760 60 794
rect 0 726 60 760
rect 0 692 11 726
rect 45 692 60 726
rect 0 658 60 692
rect 0 624 11 658
rect 45 624 60 658
rect 0 590 60 624
rect 0 556 11 590
rect 45 556 60 590
rect 0 522 60 556
rect 0 488 11 522
rect 45 488 60 522
rect 0 454 60 488
rect 0 420 11 454
rect 45 420 60 454
rect 0 386 60 420
rect 0 352 11 386
rect 45 352 60 386
rect 0 318 60 352
rect 0 284 11 318
rect 45 284 60 318
rect 0 250 60 284
rect 0 216 11 250
rect 45 216 60 250
rect 0 182 60 216
rect 0 148 11 182
rect 45 148 60 182
rect 0 114 60 148
rect 0 80 11 114
rect 45 80 60 114
rect 0 46 60 80
rect 0 12 11 46
rect 45 12 60 46
rect 0 0 60 12
<< pdiffc >>
rect 11 2936 45 2970
rect 11 2868 45 2902
rect 11 2800 45 2834
rect 11 2732 45 2766
rect 11 2664 45 2698
rect 11 2596 45 2630
rect 11 2528 45 2562
rect 11 2460 45 2494
rect 11 2392 45 2426
rect 11 2324 45 2358
rect 11 2256 45 2290
rect 11 2188 45 2222
rect 11 2120 45 2154
rect 11 2052 45 2086
rect 11 1984 45 2018
rect 11 1916 45 1950
rect 11 1848 45 1882
rect 11 1780 45 1814
rect 11 1712 45 1746
rect 11 1644 45 1678
rect 11 1576 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1474
rect 11 1372 45 1406
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< nsubdiff >>
rect 60 2914 200 3000
rect 60 2880 79 2914
rect 113 2880 200 2914
rect 60 2846 200 2880
rect 60 2812 79 2846
rect 113 2812 200 2846
rect 60 2778 200 2812
rect 60 2744 79 2778
rect 113 2744 200 2778
rect 60 2710 200 2744
rect 60 2676 79 2710
rect 113 2676 200 2710
rect 60 2642 200 2676
rect 60 2608 79 2642
rect 113 2608 200 2642
rect 60 2574 200 2608
rect 60 2540 79 2574
rect 113 2540 200 2574
rect 60 2506 200 2540
rect 60 2472 79 2506
rect 113 2472 200 2506
rect 60 2438 200 2472
rect 60 2404 79 2438
rect 113 2404 200 2438
rect 60 2370 200 2404
rect 60 2336 79 2370
rect 113 2336 200 2370
rect 60 2302 200 2336
rect 60 2268 79 2302
rect 113 2268 200 2302
rect 60 2234 200 2268
rect 60 2200 79 2234
rect 113 2200 200 2234
rect 60 2166 200 2200
rect 60 2132 79 2166
rect 113 2132 200 2166
rect 60 2098 200 2132
rect 60 2064 79 2098
rect 113 2064 200 2098
rect 60 2030 200 2064
rect 60 1996 79 2030
rect 113 1996 200 2030
rect 60 1962 200 1996
rect 60 1928 79 1962
rect 113 1928 200 1962
rect 60 1894 200 1928
rect 60 1860 79 1894
rect 113 1860 200 1894
rect 60 1826 200 1860
rect 60 1792 79 1826
rect 113 1792 200 1826
rect 60 1758 200 1792
rect 60 1724 79 1758
rect 113 1724 200 1758
rect 60 1690 200 1724
rect 60 1656 79 1690
rect 113 1656 200 1690
rect 60 1622 200 1656
rect 60 1588 79 1622
rect 113 1588 200 1622
rect 60 1554 200 1588
rect 60 1520 79 1554
rect 113 1520 200 1554
rect 60 1486 200 1520
rect 60 1452 79 1486
rect 113 1452 200 1486
rect 60 1418 200 1452
rect 60 1384 79 1418
rect 113 1384 200 1418
rect 60 1350 200 1384
rect 60 1316 79 1350
rect 113 1316 200 1350
rect 60 1282 200 1316
rect 60 1248 79 1282
rect 113 1248 200 1282
rect 60 1214 200 1248
rect 60 1180 79 1214
rect 113 1180 200 1214
rect 60 1146 200 1180
rect 60 1112 79 1146
rect 113 1112 200 1146
rect 60 1078 200 1112
rect 60 1044 79 1078
rect 113 1044 200 1078
rect 60 1010 200 1044
rect 60 976 79 1010
rect 113 976 200 1010
rect 60 942 200 976
rect 60 908 79 942
rect 113 908 200 942
rect 60 874 200 908
rect 60 840 79 874
rect 113 840 200 874
rect 60 806 200 840
rect 60 772 79 806
rect 113 772 200 806
rect 60 738 200 772
rect 60 704 79 738
rect 113 704 200 738
rect 60 670 200 704
rect 60 636 79 670
rect 113 636 200 670
rect 60 602 200 636
rect 60 568 79 602
rect 113 568 200 602
rect 60 534 200 568
rect 60 500 79 534
rect 113 500 200 534
rect 60 466 200 500
rect 60 432 79 466
rect 113 432 200 466
rect 60 398 200 432
rect 60 364 79 398
rect 113 364 200 398
rect 60 330 200 364
rect 60 296 79 330
rect 113 296 200 330
rect 60 262 200 296
rect 60 228 79 262
rect 113 228 200 262
rect 60 194 200 228
rect 60 160 79 194
rect 113 160 200 194
rect 60 126 200 160
rect 60 92 79 126
rect 113 92 200 126
rect 60 58 200 92
rect 60 24 79 58
rect 113 24 200 58
rect 60 0 200 24
<< nsubdiffcont >>
rect 79 2880 113 2914
rect 79 2812 113 2846
rect 79 2744 113 2778
rect 79 2676 113 2710
rect 79 2608 113 2642
rect 79 2540 113 2574
rect 79 2472 113 2506
rect 79 2404 113 2438
rect 79 2336 113 2370
rect 79 2268 113 2302
rect 79 2200 113 2234
rect 79 2132 113 2166
rect 79 2064 113 2098
rect 79 1996 113 2030
rect 79 1928 113 1962
rect 79 1860 113 1894
rect 79 1792 113 1826
rect 79 1724 113 1758
rect 79 1656 113 1690
rect 79 1588 113 1622
rect 79 1520 113 1554
rect 79 1452 113 1486
rect 79 1384 113 1418
rect 79 1316 113 1350
rect 79 1248 113 1282
rect 79 1180 113 1214
rect 79 1112 113 1146
rect 79 1044 113 1078
rect 79 976 113 1010
rect 79 908 113 942
rect 79 840 113 874
rect 79 772 113 806
rect 79 704 113 738
rect 79 636 113 670
rect 79 568 113 602
rect 79 500 113 534
rect 79 432 113 466
rect 79 364 113 398
rect 79 296 113 330
rect 79 228 113 262
rect 79 160 113 194
rect 79 92 113 126
rect 79 24 113 58
<< locali >>
rect 11 2970 113 2986
rect 45 2936 113 2970
rect 11 2914 113 2936
rect 11 2902 79 2914
rect 45 2880 79 2902
rect 45 2868 113 2880
rect 11 2846 113 2868
rect 11 2834 79 2846
rect 45 2812 79 2834
rect 45 2800 113 2812
rect 11 2778 113 2800
rect 11 2766 79 2778
rect 45 2744 79 2766
rect 45 2732 113 2744
rect 11 2710 113 2732
rect 11 2698 79 2710
rect 45 2676 79 2698
rect 45 2664 113 2676
rect 11 2642 113 2664
rect 11 2630 79 2642
rect 45 2608 79 2630
rect 45 2596 113 2608
rect 11 2574 113 2596
rect 11 2562 79 2574
rect 45 2540 79 2562
rect 45 2528 113 2540
rect 11 2506 113 2528
rect 11 2494 79 2506
rect 45 2472 79 2494
rect 45 2460 113 2472
rect 11 2438 113 2460
rect 11 2426 79 2438
rect 45 2404 79 2426
rect 45 2392 113 2404
rect 11 2370 113 2392
rect 11 2358 79 2370
rect 45 2336 79 2358
rect 45 2324 113 2336
rect 11 2302 113 2324
rect 11 2290 79 2302
rect 45 2268 79 2290
rect 45 2256 113 2268
rect 11 2234 113 2256
rect 11 2222 79 2234
rect 45 2200 79 2222
rect 45 2188 113 2200
rect 11 2166 113 2188
rect 11 2154 79 2166
rect 45 2132 79 2154
rect 45 2120 113 2132
rect 11 2098 113 2120
rect 11 2086 79 2098
rect 45 2064 79 2086
rect 45 2052 113 2064
rect 11 2030 113 2052
rect 11 2018 79 2030
rect 45 1996 79 2018
rect 45 1984 113 1996
rect 11 1962 113 1984
rect 11 1950 79 1962
rect 45 1928 79 1950
rect 45 1916 113 1928
rect 11 1894 113 1916
rect 11 1882 79 1894
rect 45 1860 79 1882
rect 45 1848 113 1860
rect 11 1826 113 1848
rect 11 1814 79 1826
rect 45 1792 79 1814
rect 45 1780 113 1792
rect 11 1758 113 1780
rect 11 1746 79 1758
rect 45 1724 79 1746
rect 45 1712 113 1724
rect 11 1690 113 1712
rect 11 1678 79 1690
rect 45 1656 79 1678
rect 45 1644 113 1656
rect 11 1622 113 1644
rect 11 1610 79 1622
rect 45 1588 79 1610
rect 45 1576 113 1588
rect 11 1554 113 1576
rect 11 1542 79 1554
rect 45 1520 79 1542
rect 45 1508 113 1520
rect 11 1486 113 1508
rect 11 1474 79 1486
rect 45 1452 79 1474
rect 45 1440 113 1452
rect 11 1418 113 1440
rect 11 1406 79 1418
rect 45 1384 79 1406
rect 45 1372 113 1384
rect 11 1350 113 1372
rect 11 1338 79 1350
rect 45 1316 79 1338
rect 45 1304 113 1316
rect 11 1282 113 1304
rect 11 1270 79 1282
rect 45 1248 79 1270
rect 45 1236 113 1248
rect 11 1214 113 1236
rect 11 1202 79 1214
rect 45 1180 79 1202
rect 45 1168 113 1180
rect 11 1146 113 1168
rect 11 1134 79 1146
rect 45 1112 79 1134
rect 45 1100 113 1112
rect 11 1078 113 1100
rect 11 1066 79 1078
rect 45 1044 79 1066
rect 45 1032 113 1044
rect 11 1010 113 1032
rect 11 998 79 1010
rect 45 976 79 998
rect 45 964 113 976
rect 11 942 113 964
rect 11 930 79 942
rect 45 908 79 930
rect 45 896 113 908
rect 11 874 113 896
rect 11 862 79 874
rect 45 840 79 862
rect 45 828 113 840
rect 11 806 113 828
rect 11 794 79 806
rect 45 772 79 794
rect 45 760 113 772
rect 11 738 113 760
rect 11 726 79 738
rect 45 704 79 726
rect 45 692 113 704
rect 11 670 113 692
rect 11 658 79 670
rect 45 636 79 658
rect 45 624 113 636
rect 11 602 113 624
rect 11 590 79 602
rect 45 568 79 590
rect 45 556 113 568
rect 11 534 113 556
rect 11 522 79 534
rect 45 500 79 522
rect 45 488 113 500
rect 11 466 113 488
rect 11 454 79 466
rect 45 432 79 454
rect 45 420 113 432
rect 11 398 113 420
rect 11 386 79 398
rect 45 364 79 386
rect 45 352 113 364
rect 11 330 113 352
rect 11 318 79 330
rect 45 296 79 318
rect 45 284 113 296
rect 11 262 113 284
rect 11 250 79 262
rect 45 228 79 250
rect 45 216 113 228
rect 11 194 113 216
rect 11 182 79 194
rect 45 160 79 182
rect 45 148 113 160
rect 11 126 113 148
rect 11 114 79 126
rect 45 92 79 114
rect 45 80 113 92
rect 11 58 113 80
rect 11 46 79 58
rect 45 24 79 46
rect 45 12 113 24
rect 11 -4 113 12
<< properties >>
string GDS_END 89376642
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89370622
<< end >>
