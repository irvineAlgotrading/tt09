magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 319 266
<< mvpmos >>
rect 0 0 200 200
<< mvpdiff >>
rect -50 0 0 200
rect 200 0 250 200
<< poly >>
rect 0 200 200 226
rect 0 -26 200 0
<< metal1 >>
rect -51 -16 -5 186
rect 205 -16 251 186
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 236
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_1
timestamp 1704896540
transform 1 0 200 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 228 85 228 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85974866
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85973848
<< end >>
