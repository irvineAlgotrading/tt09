magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 721 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 493
rect 271 333 337 493
rect 543 333 609 493
rect 103 289 609 333
rect 18 199 66 265
rect 103 127 169 289
rect 214 215 432 255
rect 494 215 719 255
<< obsli1 >>
rect 0 527 736 561
rect 18 299 69 527
rect 203 367 237 527
rect 371 367 509 527
rect 643 289 719 527
rect 18 93 69 157
rect 271 127 609 181
rect 18 59 421 93
rect 459 17 525 93
rect 643 17 719 177
rect 0 -17 736 17
<< metal1 >>
rect 0 496 736 592
rect 0 -48 736 48
<< labels >>
rlabel locali s 18 199 66 265 6 A
port 1 nsew signal input
rlabel locali s 214 215 432 255 6 B
port 2 nsew signal input
rlabel locali s 494 215 719 255 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 721 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 103 127 169 289 6 Y
port 8 nsew signal output
rlabel locali s 103 289 609 333 6 Y
port 8 nsew signal output
rlabel locali s 543 333 609 493 6 Y
port 8 nsew signal output
rlabel locali s 271 333 337 493 6 Y
port 8 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1827162
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1819936
<< end >>
