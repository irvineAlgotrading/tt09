magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 2511 4522 9109 4552
rect 419 4416 9109 4522
rect 2511 3852 9109 4416
rect 2511 3851 3603 3852
rect 7107 3851 7552 3852
rect 8152 3851 9109 3852
<< pwell >>
rect 2592 3554 9001 3746
rect 2592 3532 8713 3554
rect 417 3446 8713 3532
<< mvnmos >>
rect 2671 3580 2791 3720
rect 2847 3580 2967 3720
rect 3023 3580 3143 3720
rect 3323 3580 3443 3720
rect 3623 3580 3743 3720
rect 3799 3580 3919 3720
rect 3975 3580 4095 3720
rect 4151 3580 4271 3720
rect 4327 3580 4447 3720
rect 4503 3580 4623 3720
rect 4679 3580 4799 3720
rect 4855 3580 4975 3720
rect 5031 3580 5151 3720
rect 5207 3580 5327 3720
rect 5383 3580 5503 3720
rect 5559 3580 5679 3720
rect 5735 3580 5855 3720
rect 5911 3580 6031 3720
rect 6087 3580 6207 3720
rect 6263 3580 6383 3720
rect 6439 3580 6559 3720
rect 6615 3580 6735 3720
rect 6791 3580 6911 3720
rect 6967 3580 7087 3720
rect 7267 3580 7387 3720
rect 7443 3580 7563 3720
rect 7619 3580 7739 3720
rect 7795 3580 7915 3720
rect 7971 3580 8091 3720
rect 8271 3580 8391 3720
rect 8447 3580 8567 3720
rect 8623 3580 8743 3720
rect 8799 3580 8919 3720
<< mvpmos >>
rect 2671 4186 2791 4386
rect 2847 4186 2967 4386
rect 3023 4186 3143 4386
rect 3323 4186 3443 4386
rect 3623 4186 3743 4386
rect 3799 4186 3919 4386
rect 3975 4186 4095 4386
rect 4151 4186 4271 4386
rect 4327 4186 4447 4386
rect 4503 4186 4623 4386
rect 4679 4186 4799 4386
rect 4855 4186 4975 4386
rect 5031 4186 5151 4386
rect 5207 4186 5327 4386
rect 5383 4186 5503 4386
rect 5559 4186 5679 4386
rect 5735 4186 5855 4386
rect 5911 4186 6031 4386
rect 6087 4186 6207 4386
rect 6263 4186 6383 4386
rect 6439 4186 6559 4386
rect 6615 4186 6735 4386
rect 6791 4186 6911 4386
rect 6967 4186 7087 4386
rect 7267 4186 7387 4386
rect 7443 4186 7563 4386
rect 7619 4186 7739 4386
rect 7795 4186 7915 4386
rect 7971 4186 8091 4386
rect 8271 4186 8391 4386
rect 8447 4186 8567 4386
rect 8623 4186 8743 4386
rect 8799 4186 8919 4386
rect 2671 3918 2791 4118
rect 2847 3918 2967 4118
rect 3023 3918 3143 4118
rect 3323 3918 3443 4118
rect 3623 3918 3743 4118
rect 3799 3918 3919 4118
rect 3975 3918 4095 4118
rect 4151 3918 4271 4118
rect 4327 3918 4447 4118
rect 4503 3918 4623 4118
rect 4679 3918 4799 4118
rect 4855 3918 4975 4118
rect 5031 3918 5151 4118
rect 5207 3918 5327 4118
rect 5383 3918 5503 4118
rect 5559 3918 5679 4118
rect 5735 3918 5855 4118
rect 5911 3918 6031 4118
rect 6087 3918 6207 4118
rect 6263 3918 6383 4118
rect 6439 3918 6559 4118
rect 6615 3918 6735 4118
rect 6791 3918 6911 4118
rect 6967 3918 7087 4118
rect 7267 3918 7387 4118
rect 7443 3918 7563 4118
rect 7619 3918 7739 4118
rect 7795 3918 7915 4118
rect 7971 3918 8091 4118
rect 8271 3918 8391 4118
rect 8447 3918 8567 4118
rect 8623 3918 8743 4118
rect 8799 3918 8919 4118
<< mvndiff >>
rect 2618 3708 2671 3720
rect 2618 3674 2626 3708
rect 2660 3674 2671 3708
rect 2618 3640 2671 3674
rect 2618 3606 2626 3640
rect 2660 3606 2671 3640
rect 2618 3580 2671 3606
rect 2791 3708 2847 3720
rect 2791 3674 2802 3708
rect 2836 3674 2847 3708
rect 2791 3640 2847 3674
rect 2791 3606 2802 3640
rect 2836 3606 2847 3640
rect 2791 3580 2847 3606
rect 2967 3580 3023 3720
rect 3143 3708 3196 3720
rect 3143 3674 3154 3708
rect 3188 3674 3196 3708
rect 3143 3640 3196 3674
rect 3143 3606 3154 3640
rect 3188 3606 3196 3640
rect 3143 3580 3196 3606
rect 3270 3708 3323 3720
rect 3270 3674 3278 3708
rect 3312 3674 3323 3708
rect 3270 3640 3323 3674
rect 3270 3606 3278 3640
rect 3312 3606 3323 3640
rect 3270 3580 3323 3606
rect 3443 3708 3496 3720
rect 3443 3674 3454 3708
rect 3488 3674 3496 3708
rect 3443 3640 3496 3674
rect 3443 3606 3454 3640
rect 3488 3606 3496 3640
rect 3443 3580 3496 3606
rect 3570 3708 3623 3720
rect 3570 3674 3578 3708
rect 3612 3674 3623 3708
rect 3570 3640 3623 3674
rect 3570 3606 3578 3640
rect 3612 3606 3623 3640
rect 3570 3580 3623 3606
rect 3743 3708 3799 3720
rect 3743 3674 3754 3708
rect 3788 3674 3799 3708
rect 3743 3640 3799 3674
rect 3743 3606 3754 3640
rect 3788 3606 3799 3640
rect 3743 3580 3799 3606
rect 3919 3708 3975 3720
rect 3919 3674 3930 3708
rect 3964 3674 3975 3708
rect 3919 3640 3975 3674
rect 3919 3606 3930 3640
rect 3964 3606 3975 3640
rect 3919 3580 3975 3606
rect 4095 3708 4151 3720
rect 4095 3674 4106 3708
rect 4140 3674 4151 3708
rect 4095 3640 4151 3674
rect 4095 3606 4106 3640
rect 4140 3606 4151 3640
rect 4095 3580 4151 3606
rect 4271 3708 4327 3720
rect 4271 3674 4282 3708
rect 4316 3674 4327 3708
rect 4271 3640 4327 3674
rect 4271 3606 4282 3640
rect 4316 3606 4327 3640
rect 4271 3580 4327 3606
rect 4447 3708 4503 3720
rect 4447 3674 4458 3708
rect 4492 3674 4503 3708
rect 4447 3640 4503 3674
rect 4447 3606 4458 3640
rect 4492 3606 4503 3640
rect 4447 3580 4503 3606
rect 4623 3708 4679 3720
rect 4623 3674 4634 3708
rect 4668 3674 4679 3708
rect 4623 3640 4679 3674
rect 4623 3606 4634 3640
rect 4668 3606 4679 3640
rect 4623 3580 4679 3606
rect 4799 3708 4855 3720
rect 4799 3674 4810 3708
rect 4844 3674 4855 3708
rect 4799 3640 4855 3674
rect 4799 3606 4810 3640
rect 4844 3606 4855 3640
rect 4799 3580 4855 3606
rect 4975 3708 5031 3720
rect 4975 3674 4986 3708
rect 5020 3674 5031 3708
rect 4975 3640 5031 3674
rect 4975 3606 4986 3640
rect 5020 3606 5031 3640
rect 4975 3580 5031 3606
rect 5151 3708 5207 3720
rect 5151 3674 5162 3708
rect 5196 3674 5207 3708
rect 5151 3640 5207 3674
rect 5151 3606 5162 3640
rect 5196 3606 5207 3640
rect 5151 3580 5207 3606
rect 5327 3708 5383 3720
rect 5327 3674 5338 3708
rect 5372 3674 5383 3708
rect 5327 3640 5383 3674
rect 5327 3606 5338 3640
rect 5372 3606 5383 3640
rect 5327 3580 5383 3606
rect 5503 3708 5559 3720
rect 5503 3674 5514 3708
rect 5548 3674 5559 3708
rect 5503 3640 5559 3674
rect 5503 3606 5514 3640
rect 5548 3606 5559 3640
rect 5503 3580 5559 3606
rect 5679 3708 5735 3720
rect 5679 3674 5690 3708
rect 5724 3674 5735 3708
rect 5679 3640 5735 3674
rect 5679 3606 5690 3640
rect 5724 3606 5735 3640
rect 5679 3580 5735 3606
rect 5855 3708 5911 3720
rect 5855 3674 5866 3708
rect 5900 3674 5911 3708
rect 5855 3640 5911 3674
rect 5855 3606 5866 3640
rect 5900 3606 5911 3640
rect 5855 3580 5911 3606
rect 6031 3708 6087 3720
rect 6031 3674 6042 3708
rect 6076 3674 6087 3708
rect 6031 3640 6087 3674
rect 6031 3606 6042 3640
rect 6076 3606 6087 3640
rect 6031 3580 6087 3606
rect 6207 3708 6263 3720
rect 6207 3674 6218 3708
rect 6252 3674 6263 3708
rect 6207 3640 6263 3674
rect 6207 3606 6218 3640
rect 6252 3606 6263 3640
rect 6207 3580 6263 3606
rect 6383 3708 6439 3720
rect 6383 3674 6394 3708
rect 6428 3674 6439 3708
rect 6383 3640 6439 3674
rect 6383 3606 6394 3640
rect 6428 3606 6439 3640
rect 6383 3580 6439 3606
rect 6559 3708 6615 3720
rect 6559 3674 6570 3708
rect 6604 3674 6615 3708
rect 6559 3640 6615 3674
rect 6559 3606 6570 3640
rect 6604 3606 6615 3640
rect 6559 3580 6615 3606
rect 6735 3708 6791 3720
rect 6735 3674 6746 3708
rect 6780 3674 6791 3708
rect 6735 3640 6791 3674
rect 6735 3606 6746 3640
rect 6780 3606 6791 3640
rect 6735 3580 6791 3606
rect 6911 3708 6967 3720
rect 6911 3674 6922 3708
rect 6956 3674 6967 3708
rect 6911 3640 6967 3674
rect 6911 3606 6922 3640
rect 6956 3606 6967 3640
rect 6911 3580 6967 3606
rect 7087 3708 7140 3720
rect 7087 3674 7098 3708
rect 7132 3674 7140 3708
rect 7087 3640 7140 3674
rect 7087 3606 7098 3640
rect 7132 3606 7140 3640
rect 7087 3580 7140 3606
rect 7214 3708 7267 3720
rect 7214 3674 7222 3708
rect 7256 3674 7267 3708
rect 7214 3640 7267 3674
rect 7214 3606 7222 3640
rect 7256 3606 7267 3640
rect 7214 3580 7267 3606
rect 7387 3708 7443 3720
rect 7387 3674 7398 3708
rect 7432 3674 7443 3708
rect 7387 3640 7443 3674
rect 7387 3606 7398 3640
rect 7432 3606 7443 3640
rect 7387 3580 7443 3606
rect 7563 3708 7619 3720
rect 7563 3674 7574 3708
rect 7608 3674 7619 3708
rect 7563 3640 7619 3674
rect 7563 3606 7574 3640
rect 7608 3606 7619 3640
rect 7563 3580 7619 3606
rect 7739 3708 7795 3720
rect 7739 3674 7750 3708
rect 7784 3674 7795 3708
rect 7739 3640 7795 3674
rect 7739 3606 7750 3640
rect 7784 3606 7795 3640
rect 7739 3580 7795 3606
rect 7915 3708 7971 3720
rect 7915 3674 7926 3708
rect 7960 3674 7971 3708
rect 7915 3640 7971 3674
rect 7915 3606 7926 3640
rect 7960 3606 7971 3640
rect 7915 3580 7971 3606
rect 8091 3708 8144 3720
rect 8091 3674 8102 3708
rect 8136 3674 8144 3708
rect 8091 3640 8144 3674
rect 8091 3606 8102 3640
rect 8136 3606 8144 3640
rect 8091 3580 8144 3606
rect 8215 3708 8271 3720
rect 8215 3674 8226 3708
rect 8260 3674 8271 3708
rect 8215 3640 8271 3674
rect 8215 3606 8226 3640
rect 8260 3606 8271 3640
rect 8215 3580 8271 3606
rect 8391 3708 8447 3720
rect 8391 3674 8402 3708
rect 8436 3674 8447 3708
rect 8391 3640 8447 3674
rect 8391 3606 8402 3640
rect 8436 3606 8447 3640
rect 8391 3580 8447 3606
rect 8567 3708 8623 3720
rect 8567 3674 8578 3708
rect 8612 3674 8623 3708
rect 8567 3640 8623 3674
rect 8567 3606 8578 3640
rect 8612 3606 8623 3640
rect 8567 3580 8623 3606
rect 8743 3708 8799 3720
rect 8743 3674 8754 3708
rect 8788 3674 8799 3708
rect 8743 3640 8799 3674
rect 8743 3606 8754 3640
rect 8788 3606 8799 3640
rect 8743 3580 8799 3606
rect 8919 3708 8975 3720
rect 8919 3674 8930 3708
rect 8964 3674 8975 3708
rect 8919 3640 8975 3674
rect 8919 3606 8930 3640
rect 8964 3606 8975 3640
rect 8919 3580 8975 3606
<< mvpdiff >>
rect 2618 4368 2671 4386
rect 2618 4334 2626 4368
rect 2660 4334 2671 4368
rect 2618 4300 2671 4334
rect 2618 4266 2626 4300
rect 2660 4266 2671 4300
rect 2618 4232 2671 4266
rect 2618 4198 2626 4232
rect 2660 4198 2671 4232
rect 2618 4186 2671 4198
rect 2791 4368 2847 4386
rect 2791 4334 2802 4368
rect 2836 4334 2847 4368
rect 2791 4300 2847 4334
rect 2791 4266 2802 4300
rect 2836 4266 2847 4300
rect 2791 4232 2847 4266
rect 2791 4198 2802 4232
rect 2836 4198 2847 4232
rect 2791 4186 2847 4198
rect 2967 4368 3023 4386
rect 2967 4334 2978 4368
rect 3012 4334 3023 4368
rect 2967 4300 3023 4334
rect 2967 4266 2978 4300
rect 3012 4266 3023 4300
rect 2967 4232 3023 4266
rect 2967 4198 2978 4232
rect 3012 4198 3023 4232
rect 2967 4186 3023 4198
rect 3143 4368 3196 4386
rect 3143 4334 3154 4368
rect 3188 4334 3196 4368
rect 3143 4300 3196 4334
rect 3143 4266 3154 4300
rect 3188 4266 3196 4300
rect 3143 4232 3196 4266
rect 3143 4198 3154 4232
rect 3188 4198 3196 4232
rect 3143 4186 3196 4198
rect 3270 4368 3323 4386
rect 3270 4334 3278 4368
rect 3312 4334 3323 4368
rect 3270 4300 3323 4334
rect 3270 4266 3278 4300
rect 3312 4266 3323 4300
rect 3270 4232 3323 4266
rect 3270 4198 3278 4232
rect 3312 4198 3323 4232
rect 3270 4186 3323 4198
rect 3443 4368 3496 4386
rect 3443 4334 3454 4368
rect 3488 4334 3496 4368
rect 3443 4300 3496 4334
rect 3443 4266 3454 4300
rect 3488 4266 3496 4300
rect 3443 4232 3496 4266
rect 3443 4198 3454 4232
rect 3488 4198 3496 4232
rect 3443 4186 3496 4198
rect 3570 4368 3623 4386
rect 3570 4334 3578 4368
rect 3612 4334 3623 4368
rect 3570 4300 3623 4334
rect 3570 4266 3578 4300
rect 3612 4266 3623 4300
rect 3570 4232 3623 4266
rect 3570 4198 3578 4232
rect 3612 4198 3623 4232
rect 3570 4186 3623 4198
rect 3743 4368 3799 4386
rect 3743 4334 3754 4368
rect 3788 4334 3799 4368
rect 3743 4300 3799 4334
rect 3743 4266 3754 4300
rect 3788 4266 3799 4300
rect 3743 4232 3799 4266
rect 3743 4198 3754 4232
rect 3788 4198 3799 4232
rect 3743 4186 3799 4198
rect 3919 4368 3975 4386
rect 3919 4334 3930 4368
rect 3964 4334 3975 4368
rect 3919 4300 3975 4334
rect 3919 4266 3930 4300
rect 3964 4266 3975 4300
rect 3919 4232 3975 4266
rect 3919 4198 3930 4232
rect 3964 4198 3975 4232
rect 3919 4186 3975 4198
rect 4095 4368 4151 4386
rect 4095 4334 4106 4368
rect 4140 4334 4151 4368
rect 4095 4300 4151 4334
rect 4095 4266 4106 4300
rect 4140 4266 4151 4300
rect 4095 4232 4151 4266
rect 4095 4198 4106 4232
rect 4140 4198 4151 4232
rect 4095 4186 4151 4198
rect 4271 4368 4327 4386
rect 4271 4334 4282 4368
rect 4316 4334 4327 4368
rect 4271 4300 4327 4334
rect 4271 4266 4282 4300
rect 4316 4266 4327 4300
rect 4271 4232 4327 4266
rect 4271 4198 4282 4232
rect 4316 4198 4327 4232
rect 4271 4186 4327 4198
rect 4447 4368 4503 4386
rect 4447 4334 4458 4368
rect 4492 4334 4503 4368
rect 4447 4300 4503 4334
rect 4447 4266 4458 4300
rect 4492 4266 4503 4300
rect 4447 4232 4503 4266
rect 4447 4198 4458 4232
rect 4492 4198 4503 4232
rect 4447 4186 4503 4198
rect 4623 4368 4679 4386
rect 4623 4334 4634 4368
rect 4668 4334 4679 4368
rect 4623 4300 4679 4334
rect 4623 4266 4634 4300
rect 4668 4266 4679 4300
rect 4623 4232 4679 4266
rect 4623 4198 4634 4232
rect 4668 4198 4679 4232
rect 4623 4186 4679 4198
rect 4799 4368 4855 4386
rect 4799 4334 4810 4368
rect 4844 4334 4855 4368
rect 4799 4300 4855 4334
rect 4799 4266 4810 4300
rect 4844 4266 4855 4300
rect 4799 4232 4855 4266
rect 4799 4198 4810 4232
rect 4844 4198 4855 4232
rect 4799 4186 4855 4198
rect 4975 4368 5031 4386
rect 4975 4334 4986 4368
rect 5020 4334 5031 4368
rect 4975 4300 5031 4334
rect 4975 4266 4986 4300
rect 5020 4266 5031 4300
rect 4975 4232 5031 4266
rect 4975 4198 4986 4232
rect 5020 4198 5031 4232
rect 4975 4186 5031 4198
rect 5151 4368 5207 4386
rect 5151 4334 5162 4368
rect 5196 4334 5207 4368
rect 5151 4300 5207 4334
rect 5151 4266 5162 4300
rect 5196 4266 5207 4300
rect 5151 4232 5207 4266
rect 5151 4198 5162 4232
rect 5196 4198 5207 4232
rect 5151 4186 5207 4198
rect 5327 4368 5383 4386
rect 5327 4334 5338 4368
rect 5372 4334 5383 4368
rect 5327 4300 5383 4334
rect 5327 4266 5338 4300
rect 5372 4266 5383 4300
rect 5327 4232 5383 4266
rect 5327 4198 5338 4232
rect 5372 4198 5383 4232
rect 5327 4186 5383 4198
rect 5503 4368 5559 4386
rect 5503 4334 5514 4368
rect 5548 4334 5559 4368
rect 5503 4300 5559 4334
rect 5503 4266 5514 4300
rect 5548 4266 5559 4300
rect 5503 4232 5559 4266
rect 5503 4198 5514 4232
rect 5548 4198 5559 4232
rect 5503 4186 5559 4198
rect 5679 4368 5735 4386
rect 5679 4334 5690 4368
rect 5724 4334 5735 4368
rect 5679 4300 5735 4334
rect 5679 4266 5690 4300
rect 5724 4266 5735 4300
rect 5679 4232 5735 4266
rect 5679 4198 5690 4232
rect 5724 4198 5735 4232
rect 5679 4186 5735 4198
rect 5855 4368 5911 4386
rect 5855 4334 5866 4368
rect 5900 4334 5911 4368
rect 5855 4300 5911 4334
rect 5855 4266 5866 4300
rect 5900 4266 5911 4300
rect 5855 4232 5911 4266
rect 5855 4198 5866 4232
rect 5900 4198 5911 4232
rect 5855 4186 5911 4198
rect 6031 4368 6087 4386
rect 6031 4334 6042 4368
rect 6076 4334 6087 4368
rect 6031 4300 6087 4334
rect 6031 4266 6042 4300
rect 6076 4266 6087 4300
rect 6031 4232 6087 4266
rect 6031 4198 6042 4232
rect 6076 4198 6087 4232
rect 6031 4186 6087 4198
rect 6207 4368 6263 4386
rect 6207 4334 6218 4368
rect 6252 4334 6263 4368
rect 6207 4300 6263 4334
rect 6207 4266 6218 4300
rect 6252 4266 6263 4300
rect 6207 4232 6263 4266
rect 6207 4198 6218 4232
rect 6252 4198 6263 4232
rect 6207 4186 6263 4198
rect 6383 4368 6439 4386
rect 6383 4334 6394 4368
rect 6428 4334 6439 4368
rect 6383 4300 6439 4334
rect 6383 4266 6394 4300
rect 6428 4266 6439 4300
rect 6383 4232 6439 4266
rect 6383 4198 6394 4232
rect 6428 4198 6439 4232
rect 6383 4186 6439 4198
rect 6559 4368 6615 4386
rect 6559 4334 6570 4368
rect 6604 4334 6615 4368
rect 6559 4300 6615 4334
rect 6559 4266 6570 4300
rect 6604 4266 6615 4300
rect 6559 4232 6615 4266
rect 6559 4198 6570 4232
rect 6604 4198 6615 4232
rect 6559 4186 6615 4198
rect 6735 4368 6791 4386
rect 6735 4334 6746 4368
rect 6780 4334 6791 4368
rect 6735 4300 6791 4334
rect 6735 4266 6746 4300
rect 6780 4266 6791 4300
rect 6735 4232 6791 4266
rect 6735 4198 6746 4232
rect 6780 4198 6791 4232
rect 6735 4186 6791 4198
rect 6911 4368 6967 4386
rect 6911 4334 6922 4368
rect 6956 4334 6967 4368
rect 6911 4300 6967 4334
rect 6911 4266 6922 4300
rect 6956 4266 6967 4300
rect 6911 4232 6967 4266
rect 6911 4198 6922 4232
rect 6956 4198 6967 4232
rect 6911 4186 6967 4198
rect 7087 4368 7140 4386
rect 7087 4334 7098 4368
rect 7132 4334 7140 4368
rect 7087 4300 7140 4334
rect 7087 4266 7098 4300
rect 7132 4266 7140 4300
rect 7087 4232 7140 4266
rect 7087 4198 7098 4232
rect 7132 4198 7140 4232
rect 7087 4186 7140 4198
rect 7214 4368 7267 4386
rect 7214 4334 7222 4368
rect 7256 4334 7267 4368
rect 7214 4300 7267 4334
rect 7214 4266 7222 4300
rect 7256 4266 7267 4300
rect 7214 4232 7267 4266
rect 7214 4198 7222 4232
rect 7256 4198 7267 4232
rect 7214 4186 7267 4198
rect 7387 4368 7443 4386
rect 7387 4334 7398 4368
rect 7432 4334 7443 4368
rect 7387 4300 7443 4334
rect 7387 4266 7398 4300
rect 7432 4266 7443 4300
rect 7387 4232 7443 4266
rect 7387 4198 7398 4232
rect 7432 4198 7443 4232
rect 7387 4186 7443 4198
rect 7563 4368 7619 4386
rect 7563 4334 7574 4368
rect 7608 4334 7619 4368
rect 7563 4300 7619 4334
rect 7563 4266 7574 4300
rect 7608 4266 7619 4300
rect 7563 4232 7619 4266
rect 7563 4198 7574 4232
rect 7608 4198 7619 4232
rect 7563 4186 7619 4198
rect 7739 4368 7795 4386
rect 7739 4334 7750 4368
rect 7784 4334 7795 4368
rect 7739 4300 7795 4334
rect 7739 4266 7750 4300
rect 7784 4266 7795 4300
rect 7739 4232 7795 4266
rect 7739 4198 7750 4232
rect 7784 4198 7795 4232
rect 7739 4186 7795 4198
rect 7915 4368 7971 4386
rect 7915 4334 7926 4368
rect 7960 4334 7971 4368
rect 7915 4300 7971 4334
rect 7915 4266 7926 4300
rect 7960 4266 7971 4300
rect 7915 4232 7971 4266
rect 7915 4198 7926 4232
rect 7960 4198 7971 4232
rect 7915 4186 7971 4198
rect 8091 4368 8144 4386
rect 8091 4334 8102 4368
rect 8136 4334 8144 4368
rect 8091 4300 8144 4334
rect 8091 4266 8102 4300
rect 8136 4266 8144 4300
rect 8091 4232 8144 4266
rect 8091 4198 8102 4232
rect 8136 4198 8144 4232
rect 8091 4186 8144 4198
rect 8218 4368 8271 4386
rect 8218 4334 8226 4368
rect 8260 4334 8271 4368
rect 8218 4300 8271 4334
rect 8218 4266 8226 4300
rect 8260 4266 8271 4300
rect 8218 4232 8271 4266
rect 8218 4198 8226 4232
rect 8260 4198 8271 4232
rect 8218 4186 8271 4198
rect 8391 4368 8447 4386
rect 8391 4334 8402 4368
rect 8436 4334 8447 4368
rect 8391 4300 8447 4334
rect 8391 4266 8402 4300
rect 8436 4266 8447 4300
rect 8391 4232 8447 4266
rect 8391 4198 8402 4232
rect 8436 4198 8447 4232
rect 8391 4186 8447 4198
rect 8567 4368 8623 4386
rect 8567 4334 8578 4368
rect 8612 4334 8623 4368
rect 8567 4300 8623 4334
rect 8567 4266 8578 4300
rect 8612 4266 8623 4300
rect 8567 4232 8623 4266
rect 8567 4198 8578 4232
rect 8612 4198 8623 4232
rect 8567 4186 8623 4198
rect 8743 4368 8799 4386
rect 8743 4334 8754 4368
rect 8788 4334 8799 4368
rect 8743 4300 8799 4334
rect 8743 4266 8754 4300
rect 8788 4266 8799 4300
rect 8743 4232 8799 4266
rect 8743 4198 8754 4232
rect 8788 4198 8799 4232
rect 8743 4186 8799 4198
rect 8919 4368 8972 4386
rect 8919 4334 8930 4368
rect 8964 4334 8972 4368
rect 8919 4300 8972 4334
rect 8919 4266 8930 4300
rect 8964 4266 8972 4300
rect 8919 4232 8972 4266
rect 8919 4198 8930 4232
rect 8964 4198 8972 4232
rect 8919 4186 8972 4198
rect 2618 4106 2671 4118
rect 2618 4072 2626 4106
rect 2660 4072 2671 4106
rect 2618 4038 2671 4072
rect 2618 4004 2626 4038
rect 2660 4004 2671 4038
rect 2618 3970 2671 4004
rect 2618 3936 2626 3970
rect 2660 3936 2671 3970
rect 2618 3918 2671 3936
rect 2791 4106 2847 4118
rect 2791 4072 2802 4106
rect 2836 4072 2847 4106
rect 2791 4038 2847 4072
rect 2791 4004 2802 4038
rect 2836 4004 2847 4038
rect 2791 3970 2847 4004
rect 2791 3936 2802 3970
rect 2836 3936 2847 3970
rect 2791 3918 2847 3936
rect 2967 4106 3023 4118
rect 2967 4072 2978 4106
rect 3012 4072 3023 4106
rect 2967 4038 3023 4072
rect 2967 4004 2978 4038
rect 3012 4004 3023 4038
rect 2967 3970 3023 4004
rect 2967 3936 2978 3970
rect 3012 3936 3023 3970
rect 2967 3918 3023 3936
rect 3143 4106 3196 4118
rect 3143 4072 3154 4106
rect 3188 4072 3196 4106
rect 3143 4038 3196 4072
rect 3143 4004 3154 4038
rect 3188 4004 3196 4038
rect 3143 3970 3196 4004
rect 3143 3936 3154 3970
rect 3188 3936 3196 3970
rect 3143 3918 3196 3936
rect 3270 4106 3323 4118
rect 3270 4072 3278 4106
rect 3312 4072 3323 4106
rect 3270 4038 3323 4072
rect 3270 4004 3278 4038
rect 3312 4004 3323 4038
rect 3270 3970 3323 4004
rect 3270 3936 3278 3970
rect 3312 3936 3323 3970
rect 3270 3918 3323 3936
rect 3443 4106 3496 4118
rect 3443 4072 3454 4106
rect 3488 4072 3496 4106
rect 3443 4038 3496 4072
rect 3443 4004 3454 4038
rect 3488 4004 3496 4038
rect 3443 3970 3496 4004
rect 3443 3936 3454 3970
rect 3488 3936 3496 3970
rect 3443 3918 3496 3936
rect 3570 4106 3623 4118
rect 3570 4072 3578 4106
rect 3612 4072 3623 4106
rect 3570 4038 3623 4072
rect 3570 4004 3578 4038
rect 3612 4004 3623 4038
rect 3570 3970 3623 4004
rect 3570 3936 3578 3970
rect 3612 3936 3623 3970
rect 3570 3918 3623 3936
rect 3743 4106 3799 4118
rect 3743 4072 3754 4106
rect 3788 4072 3799 4106
rect 3743 4038 3799 4072
rect 3743 4004 3754 4038
rect 3788 4004 3799 4038
rect 3743 3970 3799 4004
rect 3743 3936 3754 3970
rect 3788 3936 3799 3970
rect 3743 3918 3799 3936
rect 3919 4106 3975 4118
rect 3919 4072 3930 4106
rect 3964 4072 3975 4106
rect 3919 4038 3975 4072
rect 3919 4004 3930 4038
rect 3964 4004 3975 4038
rect 3919 3970 3975 4004
rect 3919 3936 3930 3970
rect 3964 3936 3975 3970
rect 3919 3918 3975 3936
rect 4095 4106 4151 4118
rect 4095 4072 4106 4106
rect 4140 4072 4151 4106
rect 4095 4038 4151 4072
rect 4095 4004 4106 4038
rect 4140 4004 4151 4038
rect 4095 3970 4151 4004
rect 4095 3936 4106 3970
rect 4140 3936 4151 3970
rect 4095 3918 4151 3936
rect 4271 4106 4327 4118
rect 4271 4072 4282 4106
rect 4316 4072 4327 4106
rect 4271 4038 4327 4072
rect 4271 4004 4282 4038
rect 4316 4004 4327 4038
rect 4271 3970 4327 4004
rect 4271 3936 4282 3970
rect 4316 3936 4327 3970
rect 4271 3918 4327 3936
rect 4447 4106 4503 4118
rect 4447 4072 4458 4106
rect 4492 4072 4503 4106
rect 4447 4038 4503 4072
rect 4447 4004 4458 4038
rect 4492 4004 4503 4038
rect 4447 3970 4503 4004
rect 4447 3936 4458 3970
rect 4492 3936 4503 3970
rect 4447 3918 4503 3936
rect 4623 4106 4679 4118
rect 4623 4072 4634 4106
rect 4668 4072 4679 4106
rect 4623 4038 4679 4072
rect 4623 4004 4634 4038
rect 4668 4004 4679 4038
rect 4623 3970 4679 4004
rect 4623 3936 4634 3970
rect 4668 3936 4679 3970
rect 4623 3918 4679 3936
rect 4799 4106 4855 4118
rect 4799 4072 4810 4106
rect 4844 4072 4855 4106
rect 4799 4038 4855 4072
rect 4799 4004 4810 4038
rect 4844 4004 4855 4038
rect 4799 3970 4855 4004
rect 4799 3936 4810 3970
rect 4844 3936 4855 3970
rect 4799 3918 4855 3936
rect 4975 4106 5031 4118
rect 4975 4072 4986 4106
rect 5020 4072 5031 4106
rect 4975 4038 5031 4072
rect 4975 4004 4986 4038
rect 5020 4004 5031 4038
rect 4975 3970 5031 4004
rect 4975 3936 4986 3970
rect 5020 3936 5031 3970
rect 4975 3918 5031 3936
rect 5151 4106 5207 4118
rect 5151 4072 5162 4106
rect 5196 4072 5207 4106
rect 5151 4038 5207 4072
rect 5151 4004 5162 4038
rect 5196 4004 5207 4038
rect 5151 3970 5207 4004
rect 5151 3936 5162 3970
rect 5196 3936 5207 3970
rect 5151 3918 5207 3936
rect 5327 4106 5383 4118
rect 5327 4072 5338 4106
rect 5372 4072 5383 4106
rect 5327 4038 5383 4072
rect 5327 4004 5338 4038
rect 5372 4004 5383 4038
rect 5327 3970 5383 4004
rect 5327 3936 5338 3970
rect 5372 3936 5383 3970
rect 5327 3918 5383 3936
rect 5503 4106 5559 4118
rect 5503 4072 5514 4106
rect 5548 4072 5559 4106
rect 5503 4038 5559 4072
rect 5503 4004 5514 4038
rect 5548 4004 5559 4038
rect 5503 3970 5559 4004
rect 5503 3936 5514 3970
rect 5548 3936 5559 3970
rect 5503 3918 5559 3936
rect 5679 4106 5735 4118
rect 5679 4072 5690 4106
rect 5724 4072 5735 4106
rect 5679 4038 5735 4072
rect 5679 4004 5690 4038
rect 5724 4004 5735 4038
rect 5679 3970 5735 4004
rect 5679 3936 5690 3970
rect 5724 3936 5735 3970
rect 5679 3918 5735 3936
rect 5855 4106 5911 4118
rect 5855 4072 5866 4106
rect 5900 4072 5911 4106
rect 5855 4038 5911 4072
rect 5855 4004 5866 4038
rect 5900 4004 5911 4038
rect 5855 3970 5911 4004
rect 5855 3936 5866 3970
rect 5900 3936 5911 3970
rect 5855 3918 5911 3936
rect 6031 4106 6087 4118
rect 6031 4072 6042 4106
rect 6076 4072 6087 4106
rect 6031 4038 6087 4072
rect 6031 4004 6042 4038
rect 6076 4004 6087 4038
rect 6031 3970 6087 4004
rect 6031 3936 6042 3970
rect 6076 3936 6087 3970
rect 6031 3918 6087 3936
rect 6207 4106 6263 4118
rect 6207 4072 6218 4106
rect 6252 4072 6263 4106
rect 6207 4038 6263 4072
rect 6207 4004 6218 4038
rect 6252 4004 6263 4038
rect 6207 3970 6263 4004
rect 6207 3936 6218 3970
rect 6252 3936 6263 3970
rect 6207 3918 6263 3936
rect 6383 4106 6439 4118
rect 6383 4072 6394 4106
rect 6428 4072 6439 4106
rect 6383 4038 6439 4072
rect 6383 4004 6394 4038
rect 6428 4004 6439 4038
rect 6383 3970 6439 4004
rect 6383 3936 6394 3970
rect 6428 3936 6439 3970
rect 6383 3918 6439 3936
rect 6559 4106 6615 4118
rect 6559 4072 6570 4106
rect 6604 4072 6615 4106
rect 6559 4038 6615 4072
rect 6559 4004 6570 4038
rect 6604 4004 6615 4038
rect 6559 3970 6615 4004
rect 6559 3936 6570 3970
rect 6604 3936 6615 3970
rect 6559 3918 6615 3936
rect 6735 4106 6791 4118
rect 6735 4072 6746 4106
rect 6780 4072 6791 4106
rect 6735 4038 6791 4072
rect 6735 4004 6746 4038
rect 6780 4004 6791 4038
rect 6735 3970 6791 4004
rect 6735 3936 6746 3970
rect 6780 3936 6791 3970
rect 6735 3918 6791 3936
rect 6911 4106 6967 4118
rect 6911 4072 6922 4106
rect 6956 4072 6967 4106
rect 6911 4038 6967 4072
rect 6911 4004 6922 4038
rect 6956 4004 6967 4038
rect 6911 3970 6967 4004
rect 6911 3936 6922 3970
rect 6956 3936 6967 3970
rect 6911 3918 6967 3936
rect 7087 4106 7140 4118
rect 7087 4072 7098 4106
rect 7132 4072 7140 4106
rect 7087 4038 7140 4072
rect 7087 4004 7098 4038
rect 7132 4004 7140 4038
rect 7087 3970 7140 4004
rect 7087 3936 7098 3970
rect 7132 3936 7140 3970
rect 7087 3918 7140 3936
rect 7214 4106 7267 4118
rect 7214 4072 7222 4106
rect 7256 4072 7267 4106
rect 7214 4038 7267 4072
rect 7214 4004 7222 4038
rect 7256 4004 7267 4038
rect 7214 3970 7267 4004
rect 7214 3936 7222 3970
rect 7256 3936 7267 3970
rect 7214 3918 7267 3936
rect 7387 4106 7443 4118
rect 7387 4072 7398 4106
rect 7432 4072 7443 4106
rect 7387 4038 7443 4072
rect 7387 4004 7398 4038
rect 7432 4004 7443 4038
rect 7387 3970 7443 4004
rect 7387 3936 7398 3970
rect 7432 3936 7443 3970
rect 7387 3918 7443 3936
rect 7563 4106 7619 4118
rect 7563 4072 7574 4106
rect 7608 4072 7619 4106
rect 7563 4038 7619 4072
rect 7563 4004 7574 4038
rect 7608 4004 7619 4038
rect 7563 3970 7619 4004
rect 7563 3936 7574 3970
rect 7608 3936 7619 3970
rect 7563 3918 7619 3936
rect 7739 4106 7795 4118
rect 7739 4072 7750 4106
rect 7784 4072 7795 4106
rect 7739 4038 7795 4072
rect 7739 4004 7750 4038
rect 7784 4004 7795 4038
rect 7739 3970 7795 4004
rect 7739 3936 7750 3970
rect 7784 3936 7795 3970
rect 7739 3918 7795 3936
rect 7915 4106 7971 4118
rect 7915 4072 7926 4106
rect 7960 4072 7971 4106
rect 7915 4038 7971 4072
rect 7915 4004 7926 4038
rect 7960 4004 7971 4038
rect 7915 3970 7971 4004
rect 7915 3936 7926 3970
rect 7960 3936 7971 3970
rect 7915 3918 7971 3936
rect 8091 4106 8144 4118
rect 8091 4072 8102 4106
rect 8136 4072 8144 4106
rect 8091 4038 8144 4072
rect 8091 4004 8102 4038
rect 8136 4004 8144 4038
rect 8091 3970 8144 4004
rect 8091 3936 8102 3970
rect 8136 3936 8144 3970
rect 8091 3918 8144 3936
rect 8218 4106 8271 4118
rect 8218 4072 8226 4106
rect 8260 4072 8271 4106
rect 8218 4038 8271 4072
rect 8218 4004 8226 4038
rect 8260 4004 8271 4038
rect 8218 3970 8271 4004
rect 8218 3936 8226 3970
rect 8260 3936 8271 3970
rect 8218 3918 8271 3936
rect 8391 4106 8447 4118
rect 8391 4072 8402 4106
rect 8436 4072 8447 4106
rect 8391 4038 8447 4072
rect 8391 4004 8402 4038
rect 8436 4004 8447 4038
rect 8391 3918 8447 4004
rect 8567 4106 8623 4118
rect 8567 4072 8578 4106
rect 8612 4072 8623 4106
rect 8567 4038 8623 4072
rect 8567 4004 8578 4038
rect 8612 4004 8623 4038
rect 8567 3970 8623 4004
rect 8567 3936 8578 3970
rect 8612 3936 8623 3970
rect 8567 3918 8623 3936
rect 8743 4106 8799 4118
rect 8743 4072 8754 4106
rect 8788 4072 8799 4106
rect 8743 4038 8799 4072
rect 8743 4004 8754 4038
rect 8788 4004 8799 4038
rect 8743 3918 8799 4004
rect 8919 4106 8972 4118
rect 8919 4072 8930 4106
rect 8964 4072 8972 4106
rect 8919 4038 8972 4072
rect 8919 4004 8930 4038
rect 8964 4004 8972 4038
rect 8919 3970 8972 4004
rect 8919 3936 8930 3970
rect 8964 3936 8972 3970
rect 8919 3918 8972 3936
<< mvndiffc >>
rect 2626 3674 2660 3708
rect 2626 3606 2660 3640
rect 2802 3674 2836 3708
rect 2802 3606 2836 3640
rect 3154 3674 3188 3708
rect 3154 3606 3188 3640
rect 3278 3674 3312 3708
rect 3278 3606 3312 3640
rect 3454 3674 3488 3708
rect 3454 3606 3488 3640
rect 3578 3674 3612 3708
rect 3578 3606 3612 3640
rect 3754 3674 3788 3708
rect 3754 3606 3788 3640
rect 3930 3674 3964 3708
rect 3930 3606 3964 3640
rect 4106 3674 4140 3708
rect 4106 3606 4140 3640
rect 4282 3674 4316 3708
rect 4282 3606 4316 3640
rect 4458 3674 4492 3708
rect 4458 3606 4492 3640
rect 4634 3674 4668 3708
rect 4634 3606 4668 3640
rect 4810 3674 4844 3708
rect 4810 3606 4844 3640
rect 4986 3674 5020 3708
rect 4986 3606 5020 3640
rect 5162 3674 5196 3708
rect 5162 3606 5196 3640
rect 5338 3674 5372 3708
rect 5338 3606 5372 3640
rect 5514 3674 5548 3708
rect 5514 3606 5548 3640
rect 5690 3674 5724 3708
rect 5690 3606 5724 3640
rect 5866 3674 5900 3708
rect 5866 3606 5900 3640
rect 6042 3674 6076 3708
rect 6042 3606 6076 3640
rect 6218 3674 6252 3708
rect 6218 3606 6252 3640
rect 6394 3674 6428 3708
rect 6394 3606 6428 3640
rect 6570 3674 6604 3708
rect 6570 3606 6604 3640
rect 6746 3674 6780 3708
rect 6746 3606 6780 3640
rect 6922 3674 6956 3708
rect 6922 3606 6956 3640
rect 7098 3674 7132 3708
rect 7098 3606 7132 3640
rect 7222 3674 7256 3708
rect 7222 3606 7256 3640
rect 7398 3674 7432 3708
rect 7398 3606 7432 3640
rect 7574 3674 7608 3708
rect 7574 3606 7608 3640
rect 7750 3674 7784 3708
rect 7750 3606 7784 3640
rect 7926 3674 7960 3708
rect 7926 3606 7960 3640
rect 8102 3674 8136 3708
rect 8102 3606 8136 3640
rect 8226 3674 8260 3708
rect 8226 3606 8260 3640
rect 8402 3674 8436 3708
rect 8402 3606 8436 3640
rect 8578 3674 8612 3708
rect 8578 3606 8612 3640
rect 8754 3674 8788 3708
rect 8754 3606 8788 3640
rect 8930 3674 8964 3708
rect 8930 3606 8964 3640
<< mvpdiffc >>
rect 2626 4334 2660 4368
rect 2626 4266 2660 4300
rect 2626 4198 2660 4232
rect 2802 4334 2836 4368
rect 2802 4266 2836 4300
rect 2802 4198 2836 4232
rect 2978 4334 3012 4368
rect 2978 4266 3012 4300
rect 2978 4198 3012 4232
rect 3154 4334 3188 4368
rect 3154 4266 3188 4300
rect 3154 4198 3188 4232
rect 3278 4334 3312 4368
rect 3278 4266 3312 4300
rect 3278 4198 3312 4232
rect 3454 4334 3488 4368
rect 3454 4266 3488 4300
rect 3454 4198 3488 4232
rect 3578 4334 3612 4368
rect 3578 4266 3612 4300
rect 3578 4198 3612 4232
rect 3754 4334 3788 4368
rect 3754 4266 3788 4300
rect 3754 4198 3788 4232
rect 3930 4334 3964 4368
rect 3930 4266 3964 4300
rect 3930 4198 3964 4232
rect 4106 4334 4140 4368
rect 4106 4266 4140 4300
rect 4106 4198 4140 4232
rect 4282 4334 4316 4368
rect 4282 4266 4316 4300
rect 4282 4198 4316 4232
rect 4458 4334 4492 4368
rect 4458 4266 4492 4300
rect 4458 4198 4492 4232
rect 4634 4334 4668 4368
rect 4634 4266 4668 4300
rect 4634 4198 4668 4232
rect 4810 4334 4844 4368
rect 4810 4266 4844 4300
rect 4810 4198 4844 4232
rect 4986 4334 5020 4368
rect 4986 4266 5020 4300
rect 4986 4198 5020 4232
rect 5162 4334 5196 4368
rect 5162 4266 5196 4300
rect 5162 4198 5196 4232
rect 5338 4334 5372 4368
rect 5338 4266 5372 4300
rect 5338 4198 5372 4232
rect 5514 4334 5548 4368
rect 5514 4266 5548 4300
rect 5514 4198 5548 4232
rect 5690 4334 5724 4368
rect 5690 4266 5724 4300
rect 5690 4198 5724 4232
rect 5866 4334 5900 4368
rect 5866 4266 5900 4300
rect 5866 4198 5900 4232
rect 6042 4334 6076 4368
rect 6042 4266 6076 4300
rect 6042 4198 6076 4232
rect 6218 4334 6252 4368
rect 6218 4266 6252 4300
rect 6218 4198 6252 4232
rect 6394 4334 6428 4368
rect 6394 4266 6428 4300
rect 6394 4198 6428 4232
rect 6570 4334 6604 4368
rect 6570 4266 6604 4300
rect 6570 4198 6604 4232
rect 6746 4334 6780 4368
rect 6746 4266 6780 4300
rect 6746 4198 6780 4232
rect 6922 4334 6956 4368
rect 6922 4266 6956 4300
rect 6922 4198 6956 4232
rect 7098 4334 7132 4368
rect 7098 4266 7132 4300
rect 7098 4198 7132 4232
rect 7222 4334 7256 4368
rect 7222 4266 7256 4300
rect 7222 4198 7256 4232
rect 7398 4334 7432 4368
rect 7398 4266 7432 4300
rect 7398 4198 7432 4232
rect 7574 4334 7608 4368
rect 7574 4266 7608 4300
rect 7574 4198 7608 4232
rect 7750 4334 7784 4368
rect 7750 4266 7784 4300
rect 7750 4198 7784 4232
rect 7926 4334 7960 4368
rect 7926 4266 7960 4300
rect 7926 4198 7960 4232
rect 8102 4334 8136 4368
rect 8102 4266 8136 4300
rect 8102 4198 8136 4232
rect 8226 4334 8260 4368
rect 8226 4266 8260 4300
rect 8226 4198 8260 4232
rect 8402 4334 8436 4368
rect 8402 4266 8436 4300
rect 8402 4198 8436 4232
rect 8578 4334 8612 4368
rect 8578 4266 8612 4300
rect 8578 4198 8612 4232
rect 8754 4334 8788 4368
rect 8754 4266 8788 4300
rect 8754 4198 8788 4232
rect 8930 4334 8964 4368
rect 8930 4266 8964 4300
rect 8930 4198 8964 4232
rect 2626 4072 2660 4106
rect 2626 4004 2660 4038
rect 2626 3936 2660 3970
rect 2802 4072 2836 4106
rect 2802 4004 2836 4038
rect 2802 3936 2836 3970
rect 2978 4072 3012 4106
rect 2978 4004 3012 4038
rect 2978 3936 3012 3970
rect 3154 4072 3188 4106
rect 3154 4004 3188 4038
rect 3154 3936 3188 3970
rect 3278 4072 3312 4106
rect 3278 4004 3312 4038
rect 3278 3936 3312 3970
rect 3454 4072 3488 4106
rect 3454 4004 3488 4038
rect 3454 3936 3488 3970
rect 3578 4072 3612 4106
rect 3578 4004 3612 4038
rect 3578 3936 3612 3970
rect 3754 4072 3788 4106
rect 3754 4004 3788 4038
rect 3754 3936 3788 3970
rect 3930 4072 3964 4106
rect 3930 4004 3964 4038
rect 3930 3936 3964 3970
rect 4106 4072 4140 4106
rect 4106 4004 4140 4038
rect 4106 3936 4140 3970
rect 4282 4072 4316 4106
rect 4282 4004 4316 4038
rect 4282 3936 4316 3970
rect 4458 4072 4492 4106
rect 4458 4004 4492 4038
rect 4458 3936 4492 3970
rect 4634 4072 4668 4106
rect 4634 4004 4668 4038
rect 4634 3936 4668 3970
rect 4810 4072 4844 4106
rect 4810 4004 4844 4038
rect 4810 3936 4844 3970
rect 4986 4072 5020 4106
rect 4986 4004 5020 4038
rect 4986 3936 5020 3970
rect 5162 4072 5196 4106
rect 5162 4004 5196 4038
rect 5162 3936 5196 3970
rect 5338 4072 5372 4106
rect 5338 4004 5372 4038
rect 5338 3936 5372 3970
rect 5514 4072 5548 4106
rect 5514 4004 5548 4038
rect 5514 3936 5548 3970
rect 5690 4072 5724 4106
rect 5690 4004 5724 4038
rect 5690 3936 5724 3970
rect 5866 4072 5900 4106
rect 5866 4004 5900 4038
rect 5866 3936 5900 3970
rect 6042 4072 6076 4106
rect 6042 4004 6076 4038
rect 6042 3936 6076 3970
rect 6218 4072 6252 4106
rect 6218 4004 6252 4038
rect 6218 3936 6252 3970
rect 6394 4072 6428 4106
rect 6394 4004 6428 4038
rect 6394 3936 6428 3970
rect 6570 4072 6604 4106
rect 6570 4004 6604 4038
rect 6570 3936 6604 3970
rect 6746 4072 6780 4106
rect 6746 4004 6780 4038
rect 6746 3936 6780 3970
rect 6922 4072 6956 4106
rect 6922 4004 6956 4038
rect 6922 3936 6956 3970
rect 7098 4072 7132 4106
rect 7098 4004 7132 4038
rect 7098 3936 7132 3970
rect 7222 4072 7256 4106
rect 7222 4004 7256 4038
rect 7222 3936 7256 3970
rect 7398 4072 7432 4106
rect 7398 4004 7432 4038
rect 7398 3936 7432 3970
rect 7574 4072 7608 4106
rect 7574 4004 7608 4038
rect 7574 3936 7608 3970
rect 7750 4072 7784 4106
rect 7750 4004 7784 4038
rect 7750 3936 7784 3970
rect 7926 4072 7960 4106
rect 7926 4004 7960 4038
rect 7926 3936 7960 3970
rect 8102 4072 8136 4106
rect 8102 4004 8136 4038
rect 8102 3936 8136 3970
rect 8226 4072 8260 4106
rect 8226 4004 8260 4038
rect 8226 3936 8260 3970
rect 8402 4072 8436 4106
rect 8402 4004 8436 4038
rect 8578 4072 8612 4106
rect 8578 4004 8612 4038
rect 8578 3936 8612 3970
rect 8754 4072 8788 4106
rect 8754 4004 8788 4038
rect 8930 4072 8964 4106
rect 8930 4004 8964 4038
rect 8930 3936 8964 3970
<< psubdiff >>
rect 443 3472 519 3506
rect 553 3472 587 3506
rect 621 3472 655 3506
rect 689 3472 723 3506
rect 757 3472 791 3506
rect 825 3472 859 3506
rect 893 3472 927 3506
rect 961 3472 995 3506
rect 1029 3472 1063 3506
rect 1097 3472 1131 3506
rect 1165 3472 1199 3506
rect 1233 3472 1267 3506
rect 1301 3472 1335 3506
rect 1369 3472 1403 3506
rect 1437 3472 1471 3506
rect 1505 3472 1539 3506
rect 1573 3472 1607 3506
rect 1641 3472 1675 3506
rect 1709 3472 1743 3506
rect 1777 3472 1811 3506
rect 1845 3472 1879 3506
rect 1913 3472 1947 3506
rect 1981 3472 2015 3506
rect 2049 3472 2083 3506
rect 2117 3472 2151 3506
rect 2185 3472 2219 3506
rect 2253 3472 2287 3506
rect 2321 3472 2355 3506
rect 2389 3472 2423 3506
rect 2457 3472 2491 3506
<< nsubdiff >>
rect 429 4452 479 4486
rect 513 4452 547 4486
rect 581 4452 615 4486
rect 649 4452 683 4486
rect 717 4452 751 4486
rect 785 4452 819 4486
rect 853 4452 887 4486
rect 921 4452 955 4486
rect 989 4452 1023 4486
rect 1057 4452 1091 4486
rect 1125 4452 1159 4486
rect 1193 4452 1227 4486
rect 1261 4452 1295 4486
rect 1329 4452 1363 4486
rect 1397 4452 1431 4486
rect 1465 4452 1499 4486
rect 1533 4452 1567 4486
rect 1601 4452 1635 4486
rect 1669 4452 1703 4486
rect 1737 4452 1771 4486
rect 1805 4452 1839 4486
rect 1873 4452 1907 4486
rect 1941 4452 1975 4486
rect 2009 4452 2043 4486
rect 2077 4452 2111 4486
rect 2145 4452 2179 4486
rect 2213 4452 2247 4486
rect 2281 4452 2315 4486
rect 2349 4452 2383 4486
rect 2417 4452 2451 4486
rect 2485 4452 2505 4486
<< mvpsubdiff >>
rect 2525 3472 2559 3506
rect 2593 3472 2627 3506
rect 2661 3472 2695 3506
rect 2729 3472 2763 3506
rect 2797 3472 2831 3506
rect 2865 3472 2899 3506
rect 2933 3472 2967 3506
rect 3001 3472 3035 3506
rect 3069 3472 3103 3506
rect 3137 3472 3171 3506
rect 3205 3472 3239 3506
rect 3273 3472 3307 3506
rect 3341 3472 3375 3506
rect 3409 3472 3443 3506
rect 3477 3472 3511 3506
rect 3545 3472 3579 3506
rect 3613 3472 3647 3506
rect 3681 3472 3715 3506
rect 3749 3472 3783 3506
rect 3817 3472 3851 3506
rect 3885 3472 3919 3506
rect 3953 3472 3987 3506
rect 4021 3472 4055 3506
rect 4089 3472 4123 3506
rect 4157 3472 4191 3506
rect 4225 3472 4259 3506
rect 4293 3472 4327 3506
rect 4361 3472 4395 3506
rect 4429 3472 4463 3506
rect 4497 3472 4531 3506
rect 4565 3472 4599 3506
rect 4633 3472 4667 3506
rect 4701 3472 4735 3506
rect 4769 3472 4803 3506
rect 4837 3472 4871 3506
rect 4905 3472 4939 3506
rect 4973 3472 5007 3506
rect 5041 3472 5075 3506
rect 5109 3472 5143 3506
rect 5177 3472 5211 3506
rect 5245 3472 5279 3506
rect 5313 3472 5347 3506
rect 5381 3472 5415 3506
rect 5449 3472 5483 3506
rect 5517 3472 5551 3506
rect 5585 3472 5619 3506
rect 5653 3472 5687 3506
rect 5721 3472 5755 3506
rect 5789 3472 5823 3506
rect 5857 3472 5891 3506
rect 5925 3472 5959 3506
rect 5993 3472 6027 3506
rect 6061 3472 6095 3506
rect 6129 3472 6163 3506
rect 6197 3472 6231 3506
rect 6265 3472 6299 3506
rect 6333 3472 6367 3506
rect 6401 3472 6435 3506
rect 6469 3472 6503 3506
rect 6537 3472 6571 3506
rect 6605 3472 6639 3506
rect 6673 3472 6707 3506
rect 6741 3472 6775 3506
rect 6809 3472 6843 3506
rect 6877 3472 6911 3506
rect 6945 3472 6979 3506
rect 7013 3472 7047 3506
rect 7081 3472 7115 3506
rect 7149 3472 7183 3506
rect 7217 3472 7251 3506
rect 7285 3472 7319 3506
rect 7353 3472 7387 3506
rect 7421 3472 7455 3506
rect 7489 3472 7523 3506
rect 7557 3472 7591 3506
rect 7625 3472 7659 3506
rect 7693 3472 7727 3506
rect 7761 3472 7795 3506
rect 7829 3472 7863 3506
rect 7897 3472 7931 3506
rect 7965 3472 7999 3506
rect 8033 3472 8067 3506
rect 8101 3472 8135 3506
rect 8169 3472 8203 3506
rect 8237 3472 8271 3506
rect 8305 3472 8339 3506
rect 8373 3472 8407 3506
rect 8441 3472 8475 3506
rect 8509 3472 8543 3506
rect 8577 3472 8611 3506
rect 8645 3472 8687 3506
<< mvnsubdiff >>
rect 2505 4452 2519 4486
rect 2553 4452 2587 4486
rect 2621 4452 2655 4486
rect 2689 4452 2723 4486
rect 2757 4452 2791 4486
rect 2825 4452 2859 4486
rect 2893 4452 2927 4486
rect 2961 4452 2995 4486
rect 3029 4452 3063 4486
rect 3097 4452 3131 4486
rect 3165 4452 3199 4486
rect 3233 4452 3267 4486
rect 3301 4452 3335 4486
rect 3369 4452 3403 4486
rect 3437 4452 3471 4486
rect 3505 4452 3539 4486
rect 3573 4452 3607 4486
rect 3641 4452 3675 4486
rect 3709 4452 3743 4486
rect 3777 4452 3811 4486
rect 3845 4452 3879 4486
rect 3913 4452 3947 4486
rect 3981 4452 4015 4486
rect 4049 4452 4083 4486
rect 4117 4452 4151 4486
rect 4185 4452 4219 4486
rect 4253 4452 4287 4486
rect 4321 4452 4355 4486
rect 4389 4452 4423 4486
rect 4457 4452 4491 4486
rect 4525 4452 4559 4486
rect 4593 4452 4627 4486
rect 4661 4452 4695 4486
rect 4729 4452 4763 4486
rect 4797 4452 4831 4486
rect 4865 4452 4899 4486
rect 4933 4452 4967 4486
rect 5001 4452 5035 4486
rect 5069 4452 5103 4486
rect 5137 4452 5171 4486
rect 5205 4452 5239 4486
rect 5273 4452 5307 4486
rect 5341 4452 5375 4486
rect 5409 4452 5443 4486
rect 5477 4452 5511 4486
rect 5545 4452 5579 4486
rect 5613 4452 5647 4486
rect 5681 4452 5715 4486
rect 5749 4452 5783 4486
rect 5817 4452 5851 4486
rect 5885 4452 5919 4486
rect 5953 4452 5987 4486
rect 6021 4452 6055 4486
rect 6089 4452 6123 4486
rect 6157 4452 6191 4486
rect 6225 4452 6259 4486
rect 6293 4452 6327 4486
rect 6361 4452 6395 4486
rect 6429 4452 6463 4486
rect 6497 4452 6531 4486
rect 6565 4452 6599 4486
rect 6633 4452 6667 4486
rect 6701 4452 6735 4486
rect 6769 4452 6803 4486
rect 6837 4452 6871 4486
rect 6905 4452 6939 4486
rect 6973 4452 7007 4486
rect 7041 4452 7075 4486
rect 7109 4452 7143 4486
rect 7177 4452 7211 4486
rect 7245 4452 7279 4486
rect 7313 4452 7347 4486
rect 7381 4452 7415 4486
rect 7449 4452 7483 4486
rect 7517 4452 7551 4486
rect 7585 4452 7619 4486
rect 7653 4452 7687 4486
rect 7721 4452 7755 4486
rect 7789 4452 7823 4486
rect 7857 4452 7891 4486
rect 7925 4452 7959 4486
rect 7993 4452 8027 4486
rect 8061 4452 8095 4486
rect 8129 4452 8163 4486
rect 8197 4452 8231 4486
rect 8265 4452 8299 4486
rect 8333 4452 8367 4486
rect 8401 4452 8435 4486
rect 8469 4452 8503 4486
rect 8537 4452 8571 4486
rect 8605 4452 8639 4486
rect 8673 4452 8707 4486
rect 8741 4452 8775 4486
rect 8809 4452 8843 4486
rect 8877 4452 8911 4486
rect 8945 4452 8972 4486
<< psubdiffcont >>
rect 519 3472 553 3506
rect 587 3472 621 3506
rect 655 3472 689 3506
rect 723 3472 757 3506
rect 791 3472 825 3506
rect 859 3472 893 3506
rect 927 3472 961 3506
rect 995 3472 1029 3506
rect 1063 3472 1097 3506
rect 1131 3472 1165 3506
rect 1199 3472 1233 3506
rect 1267 3472 1301 3506
rect 1335 3472 1369 3506
rect 1403 3472 1437 3506
rect 1471 3472 1505 3506
rect 1539 3472 1573 3506
rect 1607 3472 1641 3506
rect 1675 3472 1709 3506
rect 1743 3472 1777 3506
rect 1811 3472 1845 3506
rect 1879 3472 1913 3506
rect 1947 3472 1981 3506
rect 2015 3472 2049 3506
rect 2083 3472 2117 3506
rect 2151 3472 2185 3506
rect 2219 3472 2253 3506
rect 2287 3472 2321 3506
rect 2355 3472 2389 3506
rect 2423 3472 2457 3506
rect 2491 3472 2505 3506
<< nsubdiffcont >>
rect 479 4452 513 4486
rect 547 4452 581 4486
rect 615 4452 649 4486
rect 683 4452 717 4486
rect 751 4452 785 4486
rect 819 4452 853 4486
rect 887 4452 921 4486
rect 955 4452 989 4486
rect 1023 4452 1057 4486
rect 1091 4452 1125 4486
rect 1159 4452 1193 4486
rect 1227 4452 1261 4486
rect 1295 4452 1329 4486
rect 1363 4452 1397 4486
rect 1431 4452 1465 4486
rect 1499 4452 1533 4486
rect 1567 4452 1601 4486
rect 1635 4452 1669 4486
rect 1703 4452 1737 4486
rect 1771 4452 1805 4486
rect 1839 4452 1873 4486
rect 1907 4452 1941 4486
rect 1975 4452 2009 4486
rect 2043 4452 2077 4486
rect 2111 4452 2145 4486
rect 2179 4452 2213 4486
rect 2247 4452 2281 4486
rect 2315 4452 2349 4486
rect 2383 4452 2417 4486
rect 2451 4452 2485 4486
<< mvpsubdiffcont >>
rect 2505 3472 2525 3506
rect 2559 3472 2593 3506
rect 2627 3472 2661 3506
rect 2695 3472 2729 3506
rect 2763 3472 2797 3506
rect 2831 3472 2865 3506
rect 2899 3472 2933 3506
rect 2967 3472 3001 3506
rect 3035 3472 3069 3506
rect 3103 3472 3137 3506
rect 3171 3472 3205 3506
rect 3239 3472 3273 3506
rect 3307 3472 3341 3506
rect 3375 3472 3409 3506
rect 3443 3472 3477 3506
rect 3511 3472 3545 3506
rect 3579 3472 3613 3506
rect 3647 3472 3681 3506
rect 3715 3472 3749 3506
rect 3783 3472 3817 3506
rect 3851 3472 3885 3506
rect 3919 3472 3953 3506
rect 3987 3472 4021 3506
rect 4055 3472 4089 3506
rect 4123 3472 4157 3506
rect 4191 3472 4225 3506
rect 4259 3472 4293 3506
rect 4327 3472 4361 3506
rect 4395 3472 4429 3506
rect 4463 3472 4497 3506
rect 4531 3472 4565 3506
rect 4599 3472 4633 3506
rect 4667 3472 4701 3506
rect 4735 3472 4769 3506
rect 4803 3472 4837 3506
rect 4871 3472 4905 3506
rect 4939 3472 4973 3506
rect 5007 3472 5041 3506
rect 5075 3472 5109 3506
rect 5143 3472 5177 3506
rect 5211 3472 5245 3506
rect 5279 3472 5313 3506
rect 5347 3472 5381 3506
rect 5415 3472 5449 3506
rect 5483 3472 5517 3506
rect 5551 3472 5585 3506
rect 5619 3472 5653 3506
rect 5687 3472 5721 3506
rect 5755 3472 5789 3506
rect 5823 3472 5857 3506
rect 5891 3472 5925 3506
rect 5959 3472 5993 3506
rect 6027 3472 6061 3506
rect 6095 3472 6129 3506
rect 6163 3472 6197 3506
rect 6231 3472 6265 3506
rect 6299 3472 6333 3506
rect 6367 3472 6401 3506
rect 6435 3472 6469 3506
rect 6503 3472 6537 3506
rect 6571 3472 6605 3506
rect 6639 3472 6673 3506
rect 6707 3472 6741 3506
rect 6775 3472 6809 3506
rect 6843 3472 6877 3506
rect 6911 3472 6945 3506
rect 6979 3472 7013 3506
rect 7047 3472 7081 3506
rect 7115 3472 7149 3506
rect 7183 3472 7217 3506
rect 7251 3472 7285 3506
rect 7319 3472 7353 3506
rect 7387 3472 7421 3506
rect 7455 3472 7489 3506
rect 7523 3472 7557 3506
rect 7591 3472 7625 3506
rect 7659 3472 7693 3506
rect 7727 3472 7761 3506
rect 7795 3472 7829 3506
rect 7863 3472 7897 3506
rect 7931 3472 7965 3506
rect 7999 3472 8033 3506
rect 8067 3472 8101 3506
rect 8135 3472 8169 3506
rect 8203 3472 8237 3506
rect 8271 3472 8305 3506
rect 8339 3472 8373 3506
rect 8407 3472 8441 3506
rect 8475 3472 8509 3506
rect 8543 3472 8577 3506
rect 8611 3472 8645 3506
<< mvnsubdiffcont >>
rect 2519 4452 2553 4486
rect 2587 4452 2621 4486
rect 2655 4452 2689 4486
rect 2723 4452 2757 4486
rect 2791 4452 2825 4486
rect 2859 4452 2893 4486
rect 2927 4452 2961 4486
rect 2995 4452 3029 4486
rect 3063 4452 3097 4486
rect 3131 4452 3165 4486
rect 3199 4452 3233 4486
rect 3267 4452 3301 4486
rect 3335 4452 3369 4486
rect 3403 4452 3437 4486
rect 3471 4452 3505 4486
rect 3539 4452 3573 4486
rect 3607 4452 3641 4486
rect 3675 4452 3709 4486
rect 3743 4452 3777 4486
rect 3811 4452 3845 4486
rect 3879 4452 3913 4486
rect 3947 4452 3981 4486
rect 4015 4452 4049 4486
rect 4083 4452 4117 4486
rect 4151 4452 4185 4486
rect 4219 4452 4253 4486
rect 4287 4452 4321 4486
rect 4355 4452 4389 4486
rect 4423 4452 4457 4486
rect 4491 4452 4525 4486
rect 4559 4452 4593 4486
rect 4627 4452 4661 4486
rect 4695 4452 4729 4486
rect 4763 4452 4797 4486
rect 4831 4452 4865 4486
rect 4899 4452 4933 4486
rect 4967 4452 5001 4486
rect 5035 4452 5069 4486
rect 5103 4452 5137 4486
rect 5171 4452 5205 4486
rect 5239 4452 5273 4486
rect 5307 4452 5341 4486
rect 5375 4452 5409 4486
rect 5443 4452 5477 4486
rect 5511 4452 5545 4486
rect 5579 4452 5613 4486
rect 5647 4452 5681 4486
rect 5715 4452 5749 4486
rect 5783 4452 5817 4486
rect 5851 4452 5885 4486
rect 5919 4452 5953 4486
rect 5987 4452 6021 4486
rect 6055 4452 6089 4486
rect 6123 4452 6157 4486
rect 6191 4452 6225 4486
rect 6259 4452 6293 4486
rect 6327 4452 6361 4486
rect 6395 4452 6429 4486
rect 6463 4452 6497 4486
rect 6531 4452 6565 4486
rect 6599 4452 6633 4486
rect 6667 4452 6701 4486
rect 6735 4452 6769 4486
rect 6803 4452 6837 4486
rect 6871 4452 6905 4486
rect 6939 4452 6973 4486
rect 7007 4452 7041 4486
rect 7075 4452 7109 4486
rect 7143 4452 7177 4486
rect 7211 4452 7245 4486
rect 7279 4452 7313 4486
rect 7347 4452 7381 4486
rect 7415 4452 7449 4486
rect 7483 4452 7517 4486
rect 7551 4452 7585 4486
rect 7619 4452 7653 4486
rect 7687 4452 7721 4486
rect 7755 4452 7789 4486
rect 7823 4452 7857 4486
rect 7891 4452 7925 4486
rect 7959 4452 7993 4486
rect 8027 4452 8061 4486
rect 8095 4452 8129 4486
rect 8163 4452 8197 4486
rect 8231 4452 8265 4486
rect 8299 4452 8333 4486
rect 8367 4452 8401 4486
rect 8435 4452 8469 4486
rect 8503 4452 8537 4486
rect 8571 4452 8605 4486
rect 8639 4452 8673 4486
rect 8707 4452 8741 4486
rect 8775 4452 8809 4486
rect 8843 4452 8877 4486
rect 8911 4452 8945 4486
<< poly >>
rect 2671 4386 2791 4412
rect 2847 4386 2967 4412
rect 3023 4386 3143 4412
rect 3323 4386 3443 4412
rect 3623 4386 3743 4412
rect 3799 4386 3919 4412
rect 3975 4386 4095 4412
rect 4151 4386 4271 4412
rect 4327 4386 4447 4412
rect 4503 4386 4623 4412
rect 4679 4386 4799 4412
rect 4855 4386 4975 4412
rect 5031 4386 5151 4412
rect 5207 4386 5327 4412
rect 5383 4386 5503 4412
rect 5559 4386 5679 4412
rect 5735 4386 5855 4412
rect 5911 4386 6031 4412
rect 6087 4386 6207 4412
rect 6263 4386 6383 4412
rect 6439 4386 6559 4412
rect 6615 4386 6735 4412
rect 6791 4386 6911 4412
rect 6967 4386 7087 4412
rect 7267 4386 7387 4412
rect 7443 4386 7563 4412
rect 7619 4386 7739 4412
rect 7795 4386 7915 4412
rect 7971 4386 8091 4412
rect 8271 4386 8391 4412
rect 8447 4386 8567 4412
rect 8623 4386 8743 4412
rect 8799 4386 8919 4412
rect 2671 4118 2791 4186
rect 2847 4118 2967 4186
rect 3023 4118 3143 4186
rect 3323 4118 3443 4186
rect 3623 4118 3743 4186
rect 3799 4118 3919 4186
rect 3975 4118 4095 4186
rect 4151 4118 4271 4186
rect 4327 4118 4447 4186
rect 4503 4118 4623 4186
rect 4679 4118 4799 4186
rect 4855 4118 4975 4186
rect 5031 4118 5151 4186
rect 5207 4118 5327 4186
rect 5383 4118 5503 4186
rect 5559 4118 5679 4186
rect 5735 4118 5855 4186
rect 5911 4118 6031 4186
rect 6087 4118 6207 4186
rect 6263 4118 6383 4186
rect 6439 4118 6559 4186
rect 6615 4118 6735 4186
rect 6791 4118 6911 4186
rect 6967 4118 7087 4186
rect 7267 4118 7387 4186
rect 7443 4118 7563 4186
rect 7619 4118 7739 4186
rect 7795 4118 7915 4186
rect 7971 4118 8091 4186
rect 8271 4118 8391 4186
rect 8447 4118 8567 4186
rect 8623 4118 8743 4186
rect 8799 4118 8919 4186
rect 2671 3870 2791 3918
rect 2671 3836 2713 3870
rect 2747 3836 2791 3870
rect 2671 3802 2791 3836
rect 2671 3768 2713 3802
rect 2747 3768 2791 3802
rect 2671 3720 2791 3768
rect 2847 3870 2967 3918
rect 2847 3836 2893 3870
rect 2927 3836 2967 3870
rect 2847 3802 2967 3836
rect 2847 3768 2893 3802
rect 2927 3768 2967 3802
rect 2847 3720 2967 3768
rect 3023 3870 3143 3918
rect 3023 3836 3064 3870
rect 3098 3836 3143 3870
rect 3023 3802 3143 3836
rect 3023 3768 3064 3802
rect 3098 3768 3143 3802
rect 3023 3720 3143 3768
rect 3323 3870 3443 3918
rect 3323 3836 3367 3870
rect 3401 3836 3443 3870
rect 3323 3802 3443 3836
rect 3323 3768 3367 3802
rect 3401 3768 3443 3802
rect 3323 3720 3443 3768
rect 3623 3870 3743 3918
rect 3623 3836 3669 3870
rect 3703 3836 3743 3870
rect 3623 3802 3743 3836
rect 3623 3768 3669 3802
rect 3703 3768 3743 3802
rect 3623 3720 3743 3768
rect 3799 3843 3919 3918
rect 3975 3843 4095 3918
rect 3799 3827 4095 3843
rect 3799 3793 3822 3827
rect 3856 3793 3890 3827
rect 3924 3793 3958 3827
rect 3992 3793 4026 3827
rect 4060 3793 4095 3827
rect 3799 3777 4095 3793
rect 3799 3720 3919 3777
rect 3975 3720 4095 3777
rect 4151 3870 4271 3918
rect 4151 3836 4191 3870
rect 4225 3836 4271 3870
rect 4151 3802 4271 3836
rect 4151 3768 4191 3802
rect 4225 3768 4271 3802
rect 4151 3720 4271 3768
rect 4327 3870 4447 3918
rect 4327 3836 4374 3870
rect 4408 3836 4447 3870
rect 4327 3802 4447 3836
rect 4327 3768 4374 3802
rect 4408 3768 4447 3802
rect 4327 3720 4447 3768
rect 4503 3886 4623 3918
rect 4679 3886 4799 3918
rect 4503 3870 4799 3886
rect 4503 3836 4526 3870
rect 4560 3836 4594 3870
rect 4628 3836 4662 3870
rect 4696 3836 4730 3870
rect 4764 3836 4799 3870
rect 4503 3820 4799 3836
rect 4503 3720 4623 3820
rect 4679 3720 4799 3820
rect 4855 3886 4975 3918
rect 5031 3886 5151 3918
rect 4855 3870 5151 3886
rect 4855 3836 4881 3870
rect 4915 3836 4949 3870
rect 4983 3836 5017 3870
rect 5051 3836 5085 3870
rect 5119 3836 5151 3870
rect 4855 3820 5151 3836
rect 4855 3720 4975 3820
rect 5031 3720 5151 3820
rect 5207 3886 5327 3918
rect 5383 3886 5503 3918
rect 5207 3870 5503 3886
rect 5207 3836 5230 3870
rect 5264 3836 5298 3870
rect 5332 3836 5366 3870
rect 5400 3836 5434 3870
rect 5468 3836 5503 3870
rect 5207 3820 5503 3836
rect 5207 3720 5327 3820
rect 5383 3720 5503 3820
rect 5559 3870 5679 3918
rect 5559 3836 5605 3870
rect 5639 3836 5679 3870
rect 5559 3802 5679 3836
rect 5559 3768 5605 3802
rect 5639 3768 5679 3802
rect 5559 3720 5679 3768
rect 5735 3870 5855 3918
rect 5735 3836 5782 3870
rect 5816 3836 5855 3870
rect 5735 3802 5855 3836
rect 5735 3768 5782 3802
rect 5816 3768 5855 3802
rect 5735 3720 5855 3768
rect 5911 3886 6031 3918
rect 6087 3886 6207 3918
rect 5911 3870 6207 3886
rect 5911 3836 5934 3870
rect 5968 3836 6002 3870
rect 6036 3836 6070 3870
rect 6104 3836 6138 3870
rect 6172 3836 6207 3870
rect 5911 3820 6207 3836
rect 5911 3720 6031 3820
rect 6087 3720 6207 3820
rect 6263 3886 6383 3918
rect 6439 3886 6559 3918
rect 6263 3870 6559 3886
rect 6263 3836 6289 3870
rect 6323 3836 6357 3870
rect 6391 3836 6425 3870
rect 6459 3836 6493 3870
rect 6527 3836 6559 3870
rect 6263 3820 6559 3836
rect 6263 3720 6383 3820
rect 6439 3720 6559 3820
rect 6615 3886 6735 3918
rect 6791 3886 6911 3918
rect 6615 3870 6911 3886
rect 6615 3836 6638 3870
rect 6672 3836 6706 3870
rect 6740 3836 6774 3870
rect 6808 3836 6842 3870
rect 6876 3836 6911 3870
rect 6615 3820 6911 3836
rect 6615 3720 6735 3820
rect 6791 3720 6911 3820
rect 6967 3870 7087 3918
rect 6967 3836 7013 3870
rect 7047 3836 7087 3870
rect 6967 3802 7087 3836
rect 6967 3768 7013 3802
rect 7047 3768 7087 3802
rect 6967 3720 7087 3768
rect 7267 3870 7387 3918
rect 7267 3836 7309 3870
rect 7343 3836 7387 3870
rect 7267 3802 7387 3836
rect 7267 3768 7309 3802
rect 7343 3768 7387 3802
rect 7267 3720 7387 3768
rect 7443 3870 7563 3918
rect 7443 3836 7489 3870
rect 7523 3836 7563 3870
rect 7443 3802 7563 3836
rect 7443 3768 7489 3802
rect 7523 3768 7563 3802
rect 7443 3720 7563 3768
rect 7619 3843 7739 3918
rect 7795 3843 7915 3918
rect 7619 3827 7915 3843
rect 7619 3793 7642 3827
rect 7676 3793 7710 3827
rect 7744 3793 7778 3827
rect 7812 3793 7846 3827
rect 7880 3793 7915 3827
rect 7619 3777 7915 3793
rect 7619 3720 7739 3777
rect 7795 3720 7915 3777
rect 7971 3870 8091 3918
rect 7971 3836 8011 3870
rect 8045 3836 8091 3870
rect 7971 3802 8091 3836
rect 7971 3768 8011 3802
rect 8045 3768 8091 3802
rect 7971 3720 8091 3768
rect 8271 3870 8391 3918
rect 8271 3836 8312 3870
rect 8346 3836 8391 3870
rect 8271 3802 8391 3836
rect 8271 3768 8312 3802
rect 8346 3768 8391 3802
rect 8271 3720 8391 3768
rect 8447 3870 8567 3918
rect 8447 3836 8490 3870
rect 8524 3836 8567 3870
rect 8447 3802 8567 3836
rect 8447 3768 8490 3802
rect 8524 3768 8567 3802
rect 8447 3720 8567 3768
rect 8623 3870 8743 3918
rect 8623 3836 8666 3870
rect 8700 3836 8743 3870
rect 8623 3802 8743 3836
rect 8623 3768 8666 3802
rect 8700 3768 8743 3802
rect 8623 3720 8743 3768
rect 8799 3870 8919 3918
rect 8799 3836 8844 3870
rect 8878 3836 8919 3870
rect 8799 3802 8919 3836
rect 8799 3768 8844 3802
rect 8878 3768 8919 3802
rect 8799 3720 8919 3768
rect 2671 3554 2791 3580
rect 2847 3554 2967 3580
rect 3023 3554 3143 3580
rect 3323 3554 3443 3580
rect 3623 3554 3743 3580
rect 3799 3554 3919 3580
rect 3975 3554 4095 3580
rect 4151 3554 4271 3580
rect 4327 3554 4447 3580
rect 4503 3554 4623 3580
rect 4679 3554 4799 3580
rect 4855 3554 4975 3580
rect 5031 3554 5151 3580
rect 5207 3554 5327 3580
rect 5383 3554 5503 3580
rect 5559 3554 5679 3580
rect 5735 3554 5855 3580
rect 5911 3554 6031 3580
rect 6087 3554 6207 3580
rect 6263 3554 6383 3580
rect 6439 3554 6559 3580
rect 6615 3554 6735 3580
rect 6791 3554 6911 3580
rect 6967 3554 7087 3580
rect 7267 3554 7387 3580
rect 7443 3554 7563 3580
rect 7619 3554 7739 3580
rect 7795 3554 7915 3580
rect 7971 3554 8091 3580
rect 8271 3554 8391 3580
rect 8447 3554 8567 3580
rect 8623 3554 8743 3580
rect 8799 3554 8919 3580
<< polycont >>
rect 2713 3836 2747 3870
rect 2713 3768 2747 3802
rect 2893 3836 2927 3870
rect 2893 3768 2927 3802
rect 3064 3836 3098 3870
rect 3064 3768 3098 3802
rect 3367 3836 3401 3870
rect 3367 3768 3401 3802
rect 3669 3836 3703 3870
rect 3669 3768 3703 3802
rect 3822 3793 3856 3827
rect 3890 3793 3924 3827
rect 3958 3793 3992 3827
rect 4026 3793 4060 3827
rect 4191 3836 4225 3870
rect 4191 3768 4225 3802
rect 4374 3836 4408 3870
rect 4374 3768 4408 3802
rect 4526 3836 4560 3870
rect 4594 3836 4628 3870
rect 4662 3836 4696 3870
rect 4730 3836 4764 3870
rect 4881 3836 4915 3870
rect 4949 3836 4983 3870
rect 5017 3836 5051 3870
rect 5085 3836 5119 3870
rect 5230 3836 5264 3870
rect 5298 3836 5332 3870
rect 5366 3836 5400 3870
rect 5434 3836 5468 3870
rect 5605 3836 5639 3870
rect 5605 3768 5639 3802
rect 5782 3836 5816 3870
rect 5782 3768 5816 3802
rect 5934 3836 5968 3870
rect 6002 3836 6036 3870
rect 6070 3836 6104 3870
rect 6138 3836 6172 3870
rect 6289 3836 6323 3870
rect 6357 3836 6391 3870
rect 6425 3836 6459 3870
rect 6493 3836 6527 3870
rect 6638 3836 6672 3870
rect 6706 3836 6740 3870
rect 6774 3836 6808 3870
rect 6842 3836 6876 3870
rect 7013 3836 7047 3870
rect 7013 3768 7047 3802
rect 7309 3836 7343 3870
rect 7309 3768 7343 3802
rect 7489 3836 7523 3870
rect 7489 3768 7523 3802
rect 7642 3793 7676 3827
rect 7710 3793 7744 3827
rect 7778 3793 7812 3827
rect 7846 3793 7880 3827
rect 8011 3836 8045 3870
rect 8011 3768 8045 3802
rect 8312 3836 8346 3870
rect 8312 3768 8346 3802
rect 8490 3836 8524 3870
rect 8490 3768 8524 3802
rect 8666 3836 8700 3870
rect 8666 3768 8700 3802
rect 8844 3836 8878 3870
rect 8844 3768 8878 3802
<< locali >>
rect 429 4452 467 4486
rect 513 4452 539 4486
rect 581 4452 611 4486
rect 649 4452 683 4486
rect 717 4452 751 4486
rect 789 4452 819 4486
rect 861 4452 887 4486
rect 933 4452 955 4486
rect 1005 4452 1023 4486
rect 1077 4452 1091 4486
rect 1149 4452 1159 4486
rect 1221 4452 1227 4486
rect 1293 4452 1295 4486
rect 1329 4452 1331 4486
rect 1397 4452 1403 4486
rect 1465 4452 1475 4486
rect 1533 4452 1547 4486
rect 1601 4452 1619 4486
rect 1669 4452 1691 4486
rect 1737 4452 1763 4486
rect 1805 4452 1835 4486
rect 1873 4452 1907 4486
rect 1941 4452 1975 4486
rect 2013 4452 2043 4486
rect 2085 4452 2111 4486
rect 2157 4452 2179 4486
rect 2229 4452 2247 4486
rect 2301 4452 2315 4486
rect 2373 4452 2383 4486
rect 2445 4452 2451 4486
rect 2517 4452 2519 4486
rect 2553 4452 2555 4486
rect 2621 4452 2627 4486
rect 2689 4452 2699 4486
rect 2757 4452 2771 4486
rect 2825 4452 2843 4486
rect 2893 4452 2915 4486
rect 2961 4452 2987 4486
rect 3029 4452 3059 4486
rect 3097 4452 3131 4486
rect 3165 4452 3199 4486
rect 3237 4452 3267 4486
rect 3309 4452 3335 4486
rect 3381 4452 3403 4486
rect 3453 4452 3471 4486
rect 3525 4452 3539 4486
rect 3597 4452 3607 4486
rect 3669 4452 3675 4486
rect 3741 4452 3743 4486
rect 3777 4452 3779 4486
rect 3845 4452 3851 4486
rect 3913 4452 3923 4486
rect 3981 4452 3995 4486
rect 4049 4452 4067 4486
rect 4117 4452 4139 4486
rect 4185 4452 4211 4486
rect 4253 4452 4283 4486
rect 4321 4452 4355 4486
rect 4389 4452 4423 4486
rect 4461 4452 4491 4486
rect 4533 4452 4559 4486
rect 4605 4452 4627 4486
rect 4677 4452 4695 4486
rect 4749 4452 4763 4486
rect 4821 4452 4831 4486
rect 4893 4452 4899 4486
rect 4965 4452 4967 4486
rect 5001 4452 5003 4486
rect 5069 4452 5075 4486
rect 5137 4452 5147 4486
rect 5205 4452 5219 4486
rect 5273 4452 5291 4486
rect 5341 4452 5363 4486
rect 5409 4452 5435 4486
rect 5477 4452 5507 4486
rect 5545 4452 5579 4486
rect 5613 4452 5647 4486
rect 5685 4452 5715 4486
rect 5757 4452 5783 4486
rect 5829 4452 5851 4486
rect 5901 4452 5919 4486
rect 5973 4452 5987 4486
rect 6045 4452 6055 4486
rect 6117 4452 6123 4486
rect 6189 4452 6191 4486
rect 6225 4452 6227 4486
rect 6293 4452 6299 4486
rect 6361 4452 6371 4486
rect 6429 4452 6443 4486
rect 6497 4452 6515 4486
rect 6565 4452 6587 4486
rect 6633 4452 6659 4486
rect 6701 4452 6731 4486
rect 6769 4452 6803 4486
rect 6837 4452 6871 4486
rect 6909 4452 6939 4486
rect 6981 4452 7007 4486
rect 7053 4452 7075 4486
rect 7125 4452 7143 4486
rect 7197 4452 7211 4486
rect 7269 4452 7279 4486
rect 7341 4452 7347 4486
rect 7413 4452 7415 4486
rect 7449 4452 7451 4486
rect 7517 4452 7523 4486
rect 7585 4452 7595 4486
rect 7653 4452 7667 4486
rect 7721 4452 7739 4486
rect 7789 4452 7811 4486
rect 7857 4452 7883 4486
rect 7925 4452 7955 4486
rect 7993 4452 8027 4486
rect 8061 4452 8095 4486
rect 8133 4452 8163 4486
rect 8205 4452 8231 4486
rect 8277 4452 8299 4486
rect 8349 4452 8367 4486
rect 8421 4452 8435 4486
rect 8493 4452 8503 4486
rect 8565 4452 8571 4486
rect 8637 4452 8639 4486
rect 8673 4452 8675 4486
rect 8741 4452 8747 4486
rect 8809 4452 8819 4486
rect 8877 4452 8891 4486
rect 8945 4452 8972 4486
rect 2626 4368 2660 4386
rect 2626 4300 2660 4334
rect 2626 4232 2660 4266
rect 2659 4164 2660 4198
rect 2625 4126 2660 4164
rect 2659 4106 2660 4126
rect 2626 4038 2660 4072
rect 2626 3970 2660 4004
rect 2626 3743 2660 3936
rect 2802 4368 2836 4380
rect 2802 4300 2836 4308
rect 2802 4232 2836 4266
rect 2802 4106 2836 4198
rect 2802 4038 2836 4072
rect 2802 3970 2836 4004
rect 2802 3920 2836 3936
rect 2978 4368 3012 4386
rect 2978 4300 3012 4334
rect 2978 4232 3012 4266
rect 2978 4106 3012 4198
rect 2978 4038 3012 4072
rect 2978 3970 3012 4004
rect 2696 3870 2889 3885
rect 2923 3870 2943 3885
rect 2696 3836 2713 3870
rect 2747 3862 2889 3870
rect 2747 3836 2893 3862
rect 2927 3836 2943 3870
rect 2696 3824 2943 3836
rect 2696 3802 2889 3824
rect 2923 3802 2943 3824
rect 2696 3768 2713 3802
rect 2747 3790 2889 3802
rect 2747 3768 2893 3790
rect 2927 3768 2943 3802
rect 2588 3709 2626 3743
rect 2978 3726 3012 3936
rect 3154 4368 3188 4380
rect 3154 4300 3188 4308
rect 3154 4232 3188 4266
rect 3154 4106 3188 4198
rect 3154 4038 3188 4072
rect 3154 3970 3188 4004
rect 3154 3920 3188 3936
rect 3278 4368 3312 4380
rect 3278 4300 3312 4308
rect 3278 4232 3312 4266
rect 3278 4106 3312 4198
rect 3454 4368 3488 4386
rect 3454 4300 3488 4334
rect 3454 4232 3488 4266
rect 3454 4155 3488 4198
rect 3578 4368 3612 4380
rect 3578 4300 3612 4308
rect 3578 4232 3612 4266
rect 3417 4121 3455 4155
rect 3278 4038 3312 4072
rect 3278 3970 3312 4004
rect 3278 3920 3312 3936
rect 3454 4106 3488 4121
rect 3454 4038 3488 4072
rect 3454 3970 3488 4004
rect 3454 3870 3488 3936
rect 3578 4106 3612 4198
rect 3578 4038 3612 4072
rect 3578 3970 3612 4004
rect 3754 4368 3788 4386
rect 3754 4300 3788 4334
rect 3754 4232 3788 4266
rect 3754 4106 3788 4198
rect 3754 4038 3788 4072
rect 3754 3970 3788 4004
rect 3578 3920 3612 3936
rect 3753 3936 3754 3955
rect 3930 4368 3964 4380
rect 3930 4300 3964 4308
rect 3930 4232 3964 4266
rect 3930 4106 3964 4198
rect 3930 4038 3964 4072
rect 3930 3970 3964 4004
rect 3788 3936 3791 3955
rect 3753 3921 3791 3936
rect 4106 4368 4140 4386
rect 4106 4300 4140 4334
rect 4106 4232 4140 4266
rect 4106 4106 4140 4198
rect 4106 4038 4140 4072
rect 4106 3970 4140 4004
rect 3048 3843 3061 3870
rect 3048 3836 3064 3843
rect 3098 3836 3114 3870
rect 3048 3805 3114 3836
rect 3048 3771 3061 3805
rect 3095 3802 3114 3805
rect 3048 3768 3064 3771
rect 3098 3768 3114 3802
rect 3154 3836 3367 3870
rect 3401 3836 3417 3870
rect 3154 3802 3417 3836
rect 3154 3768 3367 3802
rect 3401 3768 3417 3802
rect 3454 3869 3669 3870
rect 3703 3869 3719 3870
rect 3454 3835 3466 3869
rect 3500 3835 3538 3869
rect 3572 3835 3614 3869
rect 3648 3836 3669 3869
rect 3648 3835 3686 3836
rect 3454 3802 3719 3835
rect 3454 3768 3669 3802
rect 3703 3768 3719 3802
rect 3154 3726 3232 3768
rect 2626 3708 2660 3709
rect 2626 3640 2660 3674
rect 2626 3590 2660 3606
rect 2802 3708 2836 3724
rect 2802 3663 2836 3674
rect 2802 3591 2836 3606
rect 2978 3708 3232 3726
rect 2978 3674 3154 3708
rect 3188 3674 3232 3708
rect 2978 3640 3232 3674
rect 2978 3606 3154 3640
rect 3188 3606 3232 3640
rect 2978 3589 3232 3606
rect 3278 3708 3312 3724
rect 3278 3663 3312 3674
rect 3278 3591 3312 3606
rect 3454 3708 3488 3768
rect 3454 3640 3488 3674
rect 3454 3590 3488 3606
rect 3578 3708 3612 3724
rect 3578 3663 3612 3674
rect 3578 3591 3612 3606
rect 3754 3708 3788 3921
rect 3930 3920 3964 3936
rect 4104 3936 4106 3955
rect 4282 4368 4316 4380
rect 4282 4300 4316 4308
rect 4282 4232 4316 4266
rect 4282 4106 4316 4198
rect 4282 4038 4316 4072
rect 4282 3970 4316 4004
rect 4140 3936 4142 3955
rect 4104 3921 4142 3936
rect 3822 3835 3823 3843
rect 3857 3835 3925 3869
rect 3959 3835 4026 3869
rect 3822 3827 4060 3835
rect 3856 3793 3890 3827
rect 3924 3793 3958 3827
rect 3992 3793 4026 3827
rect 3822 3777 4060 3793
rect 3754 3640 3788 3674
rect 3754 3590 3788 3606
rect 3930 3708 3964 3724
rect 3930 3663 3964 3674
rect 3930 3591 3964 3606
rect 4106 3708 4140 3921
rect 4282 3920 4316 3936
rect 4458 4368 4492 4386
rect 4458 4300 4492 4334
rect 4458 4232 4492 4266
rect 4458 4106 4492 4198
rect 4458 4038 4492 4072
rect 4458 3970 4492 4004
rect 4634 4368 4668 4380
rect 4634 4300 4668 4308
rect 4634 4232 4668 4266
rect 4634 4106 4668 4198
rect 4634 4038 4668 4072
rect 4634 3970 4668 4004
rect 4492 3921 4530 3955
rect 4810 4368 4844 4386
rect 4810 4300 4844 4334
rect 4810 4232 4844 4266
rect 4810 4106 4844 4198
rect 4810 4038 4844 4072
rect 4810 3970 4844 4004
rect 4175 3836 4191 3870
rect 4227 3836 4241 3870
rect 4358 3869 4374 3870
rect 4408 3869 4424 3870
rect 4175 3802 4241 3836
rect 4352 3836 4374 3869
rect 4352 3835 4390 3836
rect 4175 3768 4191 3802
rect 4225 3798 4241 3802
rect 4227 3768 4241 3798
rect 4358 3802 4424 3835
rect 4358 3768 4374 3802
rect 4408 3768 4424 3802
rect 4106 3640 4140 3674
rect 4106 3590 4140 3606
rect 4282 3708 4316 3724
rect 4282 3663 4316 3674
rect 4282 3591 4316 3606
rect 4458 3708 4492 3921
rect 4634 3920 4668 3936
rect 4808 3936 4810 3955
rect 4986 4368 5020 4380
rect 4986 4300 5020 4308
rect 4986 4232 5020 4266
rect 4986 4106 5020 4198
rect 4986 4038 5020 4072
rect 4986 3970 5020 4004
rect 4844 3936 4846 3955
rect 4808 3921 4846 3936
rect 5162 4368 5196 4386
rect 5162 4300 5196 4334
rect 5162 4232 5196 4266
rect 5162 4106 5196 4198
rect 5162 4038 5196 4072
rect 5162 3970 5196 4004
rect 4526 3870 4764 3886
rect 4560 3869 4594 3870
rect 4561 3836 4594 3869
rect 4628 3869 4662 3870
rect 4628 3836 4629 3869
rect 4696 3836 4730 3870
rect 4526 3835 4527 3836
rect 4561 3835 4629 3836
rect 4663 3835 4730 3836
rect 4526 3820 4764 3835
rect 4458 3640 4492 3674
rect 4458 3590 4492 3606
rect 4634 3708 4668 3724
rect 4634 3663 4668 3674
rect 4634 3591 4668 3606
rect 4810 3708 4844 3921
rect 4986 3920 5020 3936
rect 5160 3936 5162 3955
rect 5338 4368 5372 4380
rect 5338 4300 5372 4308
rect 5338 4232 5372 4266
rect 5338 4106 5372 4198
rect 5338 4038 5372 4072
rect 5338 3970 5372 4004
rect 5196 3936 5198 3955
rect 5160 3921 5198 3936
rect 5514 4368 5548 4386
rect 5514 4300 5548 4334
rect 5514 4232 5548 4266
rect 5514 4106 5548 4198
rect 5514 4038 5548 4072
rect 5514 3970 5548 4004
rect 4881 3870 5119 3886
rect 4915 3869 4949 3870
rect 4920 3836 4949 3869
rect 4983 3869 5017 3870
rect 4881 3835 4886 3836
rect 4920 3835 4983 3836
rect 5051 3869 5085 3870
rect 5051 3836 5080 3869
rect 5017 3835 5080 3836
rect 5114 3835 5119 3836
rect 4881 3820 5119 3835
rect 4810 3640 4844 3674
rect 4810 3590 4844 3606
rect 4986 3708 5020 3724
rect 4986 3663 5020 3674
rect 4986 3591 5020 3606
rect 5162 3708 5196 3921
rect 5338 3920 5372 3936
rect 5513 3936 5514 3955
rect 5690 4368 5724 4380
rect 5690 4300 5724 4308
rect 5690 4232 5724 4266
rect 5690 4106 5724 4198
rect 5690 4038 5724 4072
rect 5690 3970 5724 4004
rect 5548 3936 5551 3955
rect 5513 3921 5551 3936
rect 5866 4368 5900 4386
rect 5866 4300 5900 4334
rect 5866 4232 5900 4266
rect 5866 4106 5900 4198
rect 5866 4038 5900 4072
rect 5866 3970 5900 4004
rect 5230 3870 5468 3886
rect 5264 3869 5298 3870
rect 5265 3836 5298 3869
rect 5332 3869 5366 3870
rect 5332 3836 5333 3869
rect 5400 3836 5434 3870
rect 5230 3835 5231 3836
rect 5265 3835 5333 3836
rect 5367 3835 5434 3836
rect 5230 3820 5468 3835
rect 5162 3640 5196 3674
rect 5162 3590 5196 3606
rect 5338 3708 5372 3724
rect 5338 3663 5372 3674
rect 5338 3591 5372 3606
rect 5514 3708 5548 3921
rect 5690 3920 5724 3936
rect 5865 3936 5866 3955
rect 6042 4368 6076 4380
rect 6042 4300 6076 4308
rect 6042 4232 6076 4266
rect 6042 4106 6076 4198
rect 6042 4038 6076 4072
rect 6042 3970 6076 4004
rect 5900 3936 5903 3955
rect 5865 3921 5903 3936
rect 6218 4368 6252 4386
rect 6218 4300 6252 4334
rect 6218 4232 6252 4266
rect 6218 4106 6252 4198
rect 6218 4038 6252 4072
rect 6218 3970 6252 4004
rect 5589 3869 5605 3870
rect 5639 3869 5655 3870
rect 5766 3869 5782 3870
rect 5816 3869 5832 3870
rect 5639 3836 5654 3869
rect 5616 3835 5654 3836
rect 5760 3836 5782 3869
rect 5760 3835 5798 3836
rect 5589 3802 5655 3835
rect 5589 3768 5605 3802
rect 5639 3768 5655 3802
rect 5766 3802 5832 3835
rect 5766 3768 5782 3802
rect 5816 3768 5832 3802
rect 5514 3640 5548 3674
rect 5514 3590 5548 3606
rect 5690 3708 5724 3724
rect 5690 3663 5724 3674
rect 5690 3591 5724 3606
rect 5866 3708 5900 3921
rect 6042 3920 6076 3936
rect 6216 3936 6218 3955
rect 6394 4368 6428 4380
rect 6394 4300 6428 4308
rect 6394 4232 6428 4266
rect 6394 4106 6428 4198
rect 6394 4038 6428 4072
rect 6394 3970 6428 4004
rect 6252 3936 6254 3955
rect 6216 3921 6254 3936
rect 6570 4368 6604 4386
rect 6570 4300 6604 4334
rect 6570 4232 6604 4266
rect 6570 4106 6604 4198
rect 6570 4038 6604 4072
rect 6570 3970 6604 4004
rect 5934 3870 6172 3886
rect 5968 3869 6002 3870
rect 5969 3836 6002 3869
rect 6036 3869 6070 3870
rect 6036 3836 6037 3869
rect 6104 3836 6138 3870
rect 5934 3835 5935 3836
rect 5969 3835 6037 3836
rect 6071 3835 6138 3836
rect 5934 3820 6172 3835
rect 5866 3640 5900 3674
rect 5866 3590 5900 3606
rect 6042 3708 6076 3724
rect 6042 3663 6076 3674
rect 6042 3591 6076 3606
rect 6218 3708 6252 3921
rect 6394 3920 6428 3936
rect 6568 3936 6570 3955
rect 6746 4368 6780 4380
rect 6746 4300 6780 4308
rect 6746 4232 6780 4266
rect 6746 4106 6780 4198
rect 6746 4038 6780 4072
rect 6746 3970 6780 4004
rect 6604 3936 6606 3955
rect 6568 3921 6606 3936
rect 6922 4368 6956 4386
rect 6922 4300 6956 4334
rect 6922 4232 6956 4266
rect 6922 4106 6956 4198
rect 6922 4038 6956 4072
rect 6922 3970 6956 4004
rect 6289 3870 6527 3886
rect 6323 3869 6357 3870
rect 6328 3836 6357 3869
rect 6391 3869 6425 3870
rect 6289 3835 6294 3836
rect 6328 3835 6391 3836
rect 6459 3869 6493 3870
rect 6459 3836 6488 3869
rect 6425 3835 6488 3836
rect 6522 3835 6527 3836
rect 6289 3820 6527 3835
rect 6218 3640 6252 3674
rect 6218 3590 6252 3606
rect 6394 3708 6428 3724
rect 6394 3663 6428 3674
rect 6394 3591 6428 3606
rect 6570 3708 6604 3921
rect 6746 3920 6780 3936
rect 6921 3936 6922 3955
rect 7098 4368 7132 4380
rect 7098 4300 7132 4308
rect 7098 4232 7132 4266
rect 7098 4106 7132 4198
rect 7098 4038 7132 4072
rect 7098 3970 7132 4004
rect 6956 3936 6959 3955
rect 6921 3921 6959 3936
rect 6638 3870 6876 3886
rect 6672 3869 6706 3870
rect 6673 3836 6706 3869
rect 6740 3869 6774 3870
rect 6740 3836 6741 3869
rect 6808 3836 6842 3870
rect 6638 3835 6639 3836
rect 6673 3835 6741 3836
rect 6775 3835 6842 3836
rect 6638 3820 6876 3835
rect 6570 3640 6604 3674
rect 6570 3590 6604 3606
rect 6746 3708 6780 3724
rect 6746 3663 6780 3674
rect 6746 3591 6780 3606
rect 6922 3708 6956 3921
rect 7098 3920 7132 3936
rect 7222 4368 7256 4386
rect 7222 4300 7256 4334
rect 7222 4232 7256 4266
rect 7222 4106 7256 4198
rect 7398 4368 7432 4380
rect 7398 4300 7432 4308
rect 7398 4232 7432 4266
rect 7222 4038 7256 4072
rect 7222 3970 7256 4004
rect 7222 3931 7256 3936
rect 6997 3869 7013 3870
rect 7047 3869 7063 3870
rect 7047 3836 7062 3869
rect 7024 3835 7062 3836
rect 7222 3859 7256 3897
rect 6997 3802 7063 3835
rect 6997 3768 7013 3802
rect 7047 3768 7063 3802
rect 6922 3640 6956 3674
rect 6922 3590 6956 3606
rect 7098 3708 7132 3724
rect 7098 3663 7132 3674
rect 7098 3591 7132 3606
rect 7222 3708 7256 3825
rect 7293 4074 7359 4156
rect 7293 4040 7308 4074
rect 7342 4040 7359 4074
rect 7293 4002 7359 4040
rect 7293 3968 7308 4002
rect 7342 3968 7359 4002
rect 7293 3870 7359 3968
rect 7398 4106 7432 4198
rect 7398 4038 7432 4072
rect 7398 3970 7432 4004
rect 7574 4368 7608 4386
rect 7574 4300 7608 4334
rect 7574 4232 7608 4266
rect 7574 4106 7608 4198
rect 7574 4038 7608 4072
rect 7574 3970 7608 4004
rect 7398 3920 7432 3936
rect 7573 3936 7574 3955
rect 7750 4368 7784 4380
rect 7750 4300 7784 4308
rect 7750 4232 7784 4266
rect 7750 4106 7784 4198
rect 7750 4038 7784 4072
rect 7750 3970 7784 4004
rect 7608 3936 7611 3955
rect 7573 3921 7611 3936
rect 7926 4368 7960 4386
rect 7926 4300 7960 4334
rect 7926 4232 7960 4266
rect 7926 4106 7960 4198
rect 7926 4038 7960 4072
rect 7926 3970 7960 4004
rect 7293 3836 7309 3870
rect 7343 3836 7359 3870
rect 7473 3869 7489 3870
rect 7523 3869 7539 3870
rect 7293 3802 7359 3836
rect 7468 3836 7489 3869
rect 7468 3835 7506 3836
rect 7293 3768 7309 3802
rect 7343 3768 7359 3802
rect 7473 3802 7539 3835
rect 7473 3768 7489 3802
rect 7523 3768 7539 3802
rect 7222 3640 7256 3674
rect 7222 3590 7256 3606
rect 7398 3708 7432 3724
rect 7398 3663 7432 3674
rect 7398 3591 7432 3606
rect 7574 3708 7608 3921
rect 7750 3920 7784 3936
rect 7924 3936 7926 3955
rect 8102 4368 8136 4380
rect 8102 4300 8136 4308
rect 8102 4232 8136 4266
rect 8102 4106 8136 4198
rect 8102 4038 8136 4072
rect 8102 3970 8136 4004
rect 7960 3936 7962 3955
rect 7924 3921 7962 3936
rect 7642 3835 7643 3843
rect 7677 3835 7745 3869
rect 7779 3835 7846 3869
rect 7642 3827 7880 3835
rect 7676 3793 7710 3827
rect 7744 3793 7778 3827
rect 7812 3793 7846 3827
rect 7642 3777 7880 3793
rect 7574 3640 7608 3674
rect 7574 3590 7608 3606
rect 7750 3708 7784 3724
rect 7750 3663 7784 3674
rect 7750 3591 7784 3606
rect 7926 3708 7960 3921
rect 8102 3920 8136 3936
rect 8226 4368 8260 4414
rect 8226 4300 8260 4334
rect 8226 4232 8260 4266
rect 8226 4106 8260 4198
rect 8226 4038 8260 4072
rect 8226 3970 8260 4004
rect 8402 4368 8436 4384
rect 8402 4300 8436 4334
rect 8402 4232 8436 4266
rect 8402 4106 8436 4198
rect 8402 4038 8436 4072
rect 8578 4368 8612 4380
rect 8578 4300 8612 4308
rect 8578 4232 8612 4266
rect 8578 4106 8612 4198
rect 8754 4368 8788 4384
rect 8754 4300 8788 4334
rect 8754 4232 8788 4266
rect 8578 4038 8612 4072
rect 8402 3988 8436 4004
rect 8474 3992 8540 4019
rect 8474 3958 8486 3992
rect 8520 3958 8540 3992
rect 8260 3936 8436 3954
rect 8226 3920 8436 3936
rect 7995 3836 8011 3870
rect 8047 3836 8061 3870
rect 7995 3802 8061 3836
rect 7995 3768 8011 3802
rect 8045 3798 8061 3802
rect 8047 3768 8061 3798
rect 8226 3864 8260 3920
rect 8226 3792 8260 3830
rect 8296 3836 8312 3870
rect 8346 3836 8362 3870
rect 8296 3802 8362 3836
rect 8296 3768 8312 3802
rect 8346 3768 8362 3802
rect 7926 3640 7960 3674
rect 7926 3590 7960 3606
rect 8102 3708 8136 3724
rect 8102 3663 8136 3674
rect 8102 3591 8136 3606
rect 8226 3708 8260 3724
rect 8226 3663 8260 3674
rect 8226 3591 8260 3606
rect 8402 3708 8436 3920
rect 8474 3920 8540 3958
rect 8578 3970 8612 4004
rect 8578 3920 8612 3936
rect 8650 4149 8716 4161
rect 8650 4115 8666 4149
rect 8700 4115 8716 4149
rect 8650 4077 8716 4115
rect 8650 4043 8666 4077
rect 8700 4043 8716 4077
rect 8474 3886 8486 3920
rect 8520 3886 8540 3920
rect 8474 3870 8540 3886
rect 8474 3836 8490 3870
rect 8524 3836 8540 3870
rect 8474 3802 8540 3836
rect 8474 3768 8490 3802
rect 8524 3768 8540 3802
rect 8650 3870 8716 4043
rect 8754 4106 8788 4198
rect 8754 4038 8788 4072
rect 8754 3988 8788 4004
rect 8930 4368 8964 4414
rect 8930 4300 8964 4334
rect 8930 4232 8964 4266
rect 8930 4106 8964 4198
rect 8930 4038 8964 4072
rect 8930 3970 8964 4004
rect 8650 3836 8666 3870
rect 8700 3836 8716 3870
rect 8650 3802 8716 3836
rect 8650 3768 8666 3802
rect 8700 3768 8716 3802
rect 8754 3936 8930 3954
rect 8754 3920 8964 3936
rect 8998 4230 9064 4242
rect 8998 4196 9014 4230
rect 9048 4196 9064 4230
rect 8998 4158 9064 4196
rect 8998 4124 9014 4158
rect 9048 4124 9064 4158
rect 8754 3872 8788 3920
rect 8998 3870 9064 4124
rect 8754 3800 8788 3838
rect 8828 3836 8844 3870
rect 8878 3836 9064 3870
rect 8828 3802 9064 3836
rect 8828 3768 8844 3802
rect 8878 3768 9064 3802
rect 8402 3640 8436 3674
rect 8402 3590 8436 3606
rect 8578 3708 8612 3724
rect 8578 3663 8612 3674
rect 8578 3591 8612 3606
rect 8754 3708 8788 3766
rect 8754 3640 8788 3674
rect 8754 3590 8788 3606
rect 8930 3708 8964 3724
rect 8930 3663 8964 3674
rect 8930 3591 8964 3606
rect 443 3472 507 3506
rect 553 3472 579 3506
rect 621 3472 651 3506
rect 689 3472 723 3506
rect 757 3472 791 3506
rect 829 3472 859 3506
rect 901 3472 927 3506
rect 973 3472 995 3506
rect 1045 3472 1063 3506
rect 1117 3472 1131 3506
rect 1189 3472 1199 3506
rect 1261 3472 1267 3506
rect 1333 3472 1335 3506
rect 1369 3472 1371 3506
rect 1437 3472 1443 3506
rect 1505 3472 1515 3506
rect 1573 3472 1587 3506
rect 1641 3472 1659 3506
rect 1709 3472 1731 3506
rect 1777 3472 1803 3506
rect 1845 3472 1875 3506
rect 1913 3472 1947 3506
rect 1981 3472 2015 3506
rect 2053 3472 2083 3506
rect 2125 3472 2151 3506
rect 2197 3472 2219 3506
rect 2269 3472 2287 3506
rect 2341 3472 2355 3506
rect 2413 3472 2423 3506
rect 2485 3472 2491 3506
rect 2557 3472 2559 3506
rect 2593 3472 2595 3506
rect 2661 3472 2667 3506
rect 2729 3472 2739 3506
rect 2797 3472 2811 3506
rect 2865 3472 2883 3506
rect 2933 3472 2955 3506
rect 3001 3472 3027 3506
rect 3069 3472 3099 3506
rect 3137 3472 3171 3506
rect 3205 3472 3239 3506
rect 3277 3472 3307 3506
rect 3349 3472 3375 3506
rect 3421 3472 3443 3506
rect 3493 3472 3511 3506
rect 3565 3472 3579 3506
rect 3637 3472 3647 3506
rect 3709 3472 3715 3506
rect 3781 3472 3783 3506
rect 3817 3472 3819 3506
rect 3885 3472 3891 3506
rect 3953 3472 3963 3506
rect 4021 3472 4035 3506
rect 4089 3472 4107 3506
rect 4157 3472 4179 3506
rect 4225 3472 4251 3506
rect 4293 3472 4323 3506
rect 4361 3472 4395 3506
rect 4429 3472 4463 3506
rect 4501 3472 4531 3506
rect 4573 3472 4599 3506
rect 4645 3472 4667 3506
rect 4717 3472 4735 3506
rect 4789 3472 4803 3506
rect 4861 3472 4871 3506
rect 4933 3472 4939 3506
rect 5005 3472 5007 3506
rect 5041 3472 5043 3506
rect 5109 3472 5115 3506
rect 5177 3472 5187 3506
rect 5245 3472 5259 3506
rect 5313 3472 5331 3506
rect 5381 3472 5403 3506
rect 5449 3472 5475 3506
rect 5517 3472 5547 3506
rect 5585 3472 5619 3506
rect 5653 3472 5687 3506
rect 5725 3472 5755 3506
rect 5797 3472 5823 3506
rect 5869 3472 5891 3506
rect 5941 3472 5959 3506
rect 6013 3472 6027 3506
rect 6085 3472 6095 3506
rect 6157 3472 6163 3506
rect 6229 3472 6231 3506
rect 6265 3472 6267 3506
rect 6333 3472 6339 3506
rect 6401 3472 6411 3506
rect 6469 3472 6483 3506
rect 6537 3472 6555 3506
rect 6605 3472 6627 3506
rect 6673 3472 6699 3506
rect 6741 3472 6771 3506
rect 6809 3472 6843 3506
rect 6877 3472 6911 3506
rect 6949 3472 6979 3506
rect 7021 3472 7047 3506
rect 7093 3472 7115 3506
rect 7165 3472 7183 3506
rect 7237 3472 7251 3506
rect 7309 3472 7319 3506
rect 7381 3472 7387 3506
rect 7453 3472 7455 3506
rect 7489 3472 7491 3506
rect 7557 3472 7563 3506
rect 7625 3472 7635 3506
rect 7693 3472 7707 3506
rect 7761 3472 7779 3506
rect 7829 3472 7851 3506
rect 7897 3472 7923 3506
rect 7965 3472 7995 3506
rect 8033 3472 8067 3506
rect 8101 3472 8135 3506
rect 8173 3472 8203 3506
rect 8245 3472 8271 3506
rect 8317 3472 8339 3506
rect 8389 3472 8407 3506
rect 8461 3472 8475 3506
rect 8533 3472 8543 3506
rect 8605 3472 8611 3506
rect 8645 3472 8687 3506
<< viali >>
rect 467 4452 479 4486
rect 479 4452 501 4486
rect 539 4452 547 4486
rect 547 4452 573 4486
rect 611 4452 615 4486
rect 615 4452 645 4486
rect 683 4452 717 4486
rect 755 4452 785 4486
rect 785 4452 789 4486
rect 827 4452 853 4486
rect 853 4452 861 4486
rect 899 4452 921 4486
rect 921 4452 933 4486
rect 971 4452 989 4486
rect 989 4452 1005 4486
rect 1043 4452 1057 4486
rect 1057 4452 1077 4486
rect 1115 4452 1125 4486
rect 1125 4452 1149 4486
rect 1187 4452 1193 4486
rect 1193 4452 1221 4486
rect 1259 4452 1261 4486
rect 1261 4452 1293 4486
rect 1331 4452 1363 4486
rect 1363 4452 1365 4486
rect 1403 4452 1431 4486
rect 1431 4452 1437 4486
rect 1475 4452 1499 4486
rect 1499 4452 1509 4486
rect 1547 4452 1567 4486
rect 1567 4452 1581 4486
rect 1619 4452 1635 4486
rect 1635 4452 1653 4486
rect 1691 4452 1703 4486
rect 1703 4452 1725 4486
rect 1763 4452 1771 4486
rect 1771 4452 1797 4486
rect 1835 4452 1839 4486
rect 1839 4452 1869 4486
rect 1907 4452 1941 4486
rect 1979 4452 2009 4486
rect 2009 4452 2013 4486
rect 2051 4452 2077 4486
rect 2077 4452 2085 4486
rect 2123 4452 2145 4486
rect 2145 4452 2157 4486
rect 2195 4452 2213 4486
rect 2213 4452 2229 4486
rect 2267 4452 2281 4486
rect 2281 4452 2301 4486
rect 2339 4452 2349 4486
rect 2349 4452 2373 4486
rect 2411 4452 2417 4486
rect 2417 4452 2445 4486
rect 2483 4452 2485 4486
rect 2485 4452 2517 4486
rect 2555 4452 2587 4486
rect 2587 4452 2589 4486
rect 2627 4452 2655 4486
rect 2655 4452 2661 4486
rect 2699 4452 2723 4486
rect 2723 4452 2733 4486
rect 2771 4452 2791 4486
rect 2791 4452 2805 4486
rect 2843 4452 2859 4486
rect 2859 4452 2877 4486
rect 2915 4452 2927 4486
rect 2927 4452 2949 4486
rect 2987 4452 2995 4486
rect 2995 4452 3021 4486
rect 3059 4452 3063 4486
rect 3063 4452 3093 4486
rect 3131 4452 3165 4486
rect 3203 4452 3233 4486
rect 3233 4452 3237 4486
rect 3275 4452 3301 4486
rect 3301 4452 3309 4486
rect 3347 4452 3369 4486
rect 3369 4452 3381 4486
rect 3419 4452 3437 4486
rect 3437 4452 3453 4486
rect 3491 4452 3505 4486
rect 3505 4452 3525 4486
rect 3563 4452 3573 4486
rect 3573 4452 3597 4486
rect 3635 4452 3641 4486
rect 3641 4452 3669 4486
rect 3707 4452 3709 4486
rect 3709 4452 3741 4486
rect 3779 4452 3811 4486
rect 3811 4452 3813 4486
rect 3851 4452 3879 4486
rect 3879 4452 3885 4486
rect 3923 4452 3947 4486
rect 3947 4452 3957 4486
rect 3995 4452 4015 4486
rect 4015 4452 4029 4486
rect 4067 4452 4083 4486
rect 4083 4452 4101 4486
rect 4139 4452 4151 4486
rect 4151 4452 4173 4486
rect 4211 4452 4219 4486
rect 4219 4452 4245 4486
rect 4283 4452 4287 4486
rect 4287 4452 4317 4486
rect 4355 4452 4389 4486
rect 4427 4452 4457 4486
rect 4457 4452 4461 4486
rect 4499 4452 4525 4486
rect 4525 4452 4533 4486
rect 4571 4452 4593 4486
rect 4593 4452 4605 4486
rect 4643 4452 4661 4486
rect 4661 4452 4677 4486
rect 4715 4452 4729 4486
rect 4729 4452 4749 4486
rect 4787 4452 4797 4486
rect 4797 4452 4821 4486
rect 4859 4452 4865 4486
rect 4865 4452 4893 4486
rect 4931 4452 4933 4486
rect 4933 4452 4965 4486
rect 5003 4452 5035 4486
rect 5035 4452 5037 4486
rect 5075 4452 5103 4486
rect 5103 4452 5109 4486
rect 5147 4452 5171 4486
rect 5171 4452 5181 4486
rect 5219 4452 5239 4486
rect 5239 4452 5253 4486
rect 5291 4452 5307 4486
rect 5307 4452 5325 4486
rect 5363 4452 5375 4486
rect 5375 4452 5397 4486
rect 5435 4452 5443 4486
rect 5443 4452 5469 4486
rect 5507 4452 5511 4486
rect 5511 4452 5541 4486
rect 5579 4452 5613 4486
rect 5651 4452 5681 4486
rect 5681 4452 5685 4486
rect 5723 4452 5749 4486
rect 5749 4452 5757 4486
rect 5795 4452 5817 4486
rect 5817 4452 5829 4486
rect 5867 4452 5885 4486
rect 5885 4452 5901 4486
rect 5939 4452 5953 4486
rect 5953 4452 5973 4486
rect 6011 4452 6021 4486
rect 6021 4452 6045 4486
rect 6083 4452 6089 4486
rect 6089 4452 6117 4486
rect 6155 4452 6157 4486
rect 6157 4452 6189 4486
rect 6227 4452 6259 4486
rect 6259 4452 6261 4486
rect 6299 4452 6327 4486
rect 6327 4452 6333 4486
rect 6371 4452 6395 4486
rect 6395 4452 6405 4486
rect 6443 4452 6463 4486
rect 6463 4452 6477 4486
rect 6515 4452 6531 4486
rect 6531 4452 6549 4486
rect 6587 4452 6599 4486
rect 6599 4452 6621 4486
rect 6659 4452 6667 4486
rect 6667 4452 6693 4486
rect 6731 4452 6735 4486
rect 6735 4452 6765 4486
rect 6803 4452 6837 4486
rect 6875 4452 6905 4486
rect 6905 4452 6909 4486
rect 6947 4452 6973 4486
rect 6973 4452 6981 4486
rect 7019 4452 7041 4486
rect 7041 4452 7053 4486
rect 7091 4452 7109 4486
rect 7109 4452 7125 4486
rect 7163 4452 7177 4486
rect 7177 4452 7197 4486
rect 7235 4452 7245 4486
rect 7245 4452 7269 4486
rect 7307 4452 7313 4486
rect 7313 4452 7341 4486
rect 7379 4452 7381 4486
rect 7381 4452 7413 4486
rect 7451 4452 7483 4486
rect 7483 4452 7485 4486
rect 7523 4452 7551 4486
rect 7551 4452 7557 4486
rect 7595 4452 7619 4486
rect 7619 4452 7629 4486
rect 7667 4452 7687 4486
rect 7687 4452 7701 4486
rect 7739 4452 7755 4486
rect 7755 4452 7773 4486
rect 7811 4452 7823 4486
rect 7823 4452 7845 4486
rect 7883 4452 7891 4486
rect 7891 4452 7917 4486
rect 7955 4452 7959 4486
rect 7959 4452 7989 4486
rect 8027 4452 8061 4486
rect 8099 4452 8129 4486
rect 8129 4452 8133 4486
rect 8171 4452 8197 4486
rect 8197 4452 8205 4486
rect 8243 4452 8265 4486
rect 8265 4452 8277 4486
rect 8315 4452 8333 4486
rect 8333 4452 8349 4486
rect 8387 4452 8401 4486
rect 8401 4452 8421 4486
rect 8459 4452 8469 4486
rect 8469 4452 8493 4486
rect 8531 4452 8537 4486
rect 8537 4452 8565 4486
rect 8603 4452 8605 4486
rect 8605 4452 8637 4486
rect 8675 4452 8707 4486
rect 8707 4452 8709 4486
rect 8747 4452 8775 4486
rect 8775 4452 8781 4486
rect 8819 4452 8843 4486
rect 8843 4452 8853 4486
rect 8891 4452 8911 4486
rect 8911 4452 8925 4486
rect 2625 4164 2659 4198
rect 2625 4106 2659 4126
rect 2625 4092 2626 4106
rect 2626 4092 2659 4106
rect 2802 4380 2836 4414
rect 2802 4334 2836 4342
rect 2802 4308 2836 4334
rect 2889 3870 2923 3896
rect 2889 3862 2893 3870
rect 2893 3862 2923 3870
rect 2889 3802 2923 3824
rect 2889 3790 2893 3802
rect 2893 3790 2923 3802
rect 2554 3709 2588 3743
rect 2626 3709 2660 3743
rect 3154 4380 3188 4414
rect 3154 4334 3188 4342
rect 3154 4308 3188 4334
rect 3278 4380 3312 4414
rect 3278 4334 3312 4342
rect 3278 4308 3312 4334
rect 3578 4380 3612 4414
rect 3578 4334 3612 4342
rect 3578 4308 3612 4334
rect 3383 4121 3417 4155
rect 3455 4121 3489 4155
rect 3061 3870 3095 3877
rect 3719 3921 3753 3955
rect 3930 4380 3964 4414
rect 3930 4334 3964 4342
rect 3930 4308 3964 4334
rect 3791 3921 3825 3955
rect 3061 3843 3064 3870
rect 3064 3843 3095 3870
rect 3061 3802 3095 3805
rect 3061 3771 3064 3802
rect 3064 3771 3095 3802
rect 3466 3835 3500 3869
rect 3538 3835 3572 3869
rect 3614 3835 3648 3869
rect 3686 3836 3703 3869
rect 3703 3836 3720 3869
rect 3686 3835 3720 3836
rect 2802 3640 2836 3663
rect 2802 3629 2836 3640
rect 2802 3557 2836 3591
rect 3278 3640 3312 3663
rect 3278 3629 3312 3640
rect 3278 3557 3312 3591
rect 3578 3640 3612 3663
rect 3578 3629 3612 3640
rect 3578 3557 3612 3591
rect 4070 3921 4104 3955
rect 4282 4380 4316 4414
rect 4282 4334 4316 4342
rect 4282 4308 4316 4334
rect 4142 3921 4176 3955
rect 3823 3835 3857 3869
rect 3925 3835 3959 3869
rect 4026 3835 4060 3869
rect 3930 3640 3964 3663
rect 3930 3629 3964 3640
rect 3930 3557 3964 3591
rect 4634 4380 4668 4414
rect 4634 4334 4668 4342
rect 4634 4308 4668 4334
rect 4458 3936 4492 3955
rect 4458 3921 4492 3936
rect 4530 3921 4564 3955
rect 4193 3836 4225 3870
rect 4225 3836 4227 3870
rect 4318 3835 4352 3869
rect 4390 3836 4408 3869
rect 4408 3836 4424 3869
rect 4390 3835 4424 3836
rect 4193 3768 4225 3798
rect 4225 3768 4227 3798
rect 4193 3764 4227 3768
rect 4282 3640 4316 3663
rect 4282 3629 4316 3640
rect 4282 3557 4316 3591
rect 4774 3921 4808 3955
rect 4986 4380 5020 4414
rect 4986 4334 5020 4342
rect 4986 4308 5020 4334
rect 4846 3921 4880 3955
rect 4527 3836 4560 3869
rect 4560 3836 4561 3869
rect 4629 3836 4662 3869
rect 4662 3836 4663 3869
rect 4730 3836 4764 3869
rect 4527 3835 4561 3836
rect 4629 3835 4663 3836
rect 4730 3835 4764 3836
rect 4634 3640 4668 3663
rect 4634 3629 4668 3640
rect 4634 3557 4668 3591
rect 5126 3921 5160 3955
rect 5338 4380 5372 4414
rect 5338 4334 5372 4342
rect 5338 4308 5372 4334
rect 5198 3921 5232 3955
rect 4886 3836 4915 3869
rect 4915 3836 4920 3869
rect 4886 3835 4920 3836
rect 4983 3835 5017 3869
rect 5080 3836 5085 3869
rect 5085 3836 5114 3869
rect 5080 3835 5114 3836
rect 4986 3640 5020 3663
rect 4986 3629 5020 3640
rect 4986 3557 5020 3591
rect 5479 3921 5513 3955
rect 5690 4380 5724 4414
rect 5690 4334 5724 4342
rect 5690 4308 5724 4334
rect 5551 3921 5585 3955
rect 5231 3836 5264 3869
rect 5264 3836 5265 3869
rect 5333 3836 5366 3869
rect 5366 3836 5367 3869
rect 5434 3836 5468 3869
rect 5231 3835 5265 3836
rect 5333 3835 5367 3836
rect 5434 3835 5468 3836
rect 5338 3640 5372 3663
rect 5338 3629 5372 3640
rect 5338 3557 5372 3591
rect 5831 3921 5865 3955
rect 6042 4380 6076 4414
rect 6042 4334 6076 4342
rect 6042 4308 6076 4334
rect 5903 3921 5937 3955
rect 5582 3836 5605 3869
rect 5605 3836 5616 3869
rect 5582 3835 5616 3836
rect 5654 3835 5688 3869
rect 5726 3835 5760 3869
rect 5798 3836 5816 3869
rect 5816 3836 5832 3869
rect 5798 3835 5832 3836
rect 5690 3640 5724 3663
rect 5690 3629 5724 3640
rect 5690 3557 5724 3591
rect 6182 3921 6216 3955
rect 6394 4380 6428 4414
rect 6394 4334 6428 4342
rect 6394 4308 6428 4334
rect 6254 3921 6288 3955
rect 5935 3836 5968 3869
rect 5968 3836 5969 3869
rect 6037 3836 6070 3869
rect 6070 3836 6071 3869
rect 6138 3836 6172 3869
rect 5935 3835 5969 3836
rect 6037 3835 6071 3836
rect 6138 3835 6172 3836
rect 6042 3640 6076 3663
rect 6042 3629 6076 3640
rect 6042 3557 6076 3591
rect 6534 3921 6568 3955
rect 6746 4380 6780 4414
rect 6746 4334 6780 4342
rect 6746 4308 6780 4334
rect 6606 3921 6640 3955
rect 6294 3836 6323 3869
rect 6323 3836 6328 3869
rect 6294 3835 6328 3836
rect 6391 3835 6425 3869
rect 6488 3836 6493 3869
rect 6493 3836 6522 3869
rect 6488 3835 6522 3836
rect 6394 3640 6428 3663
rect 6394 3629 6428 3640
rect 6394 3557 6428 3591
rect 6887 3921 6921 3955
rect 7098 4380 7132 4414
rect 7098 4334 7132 4342
rect 7098 4308 7132 4334
rect 6959 3921 6993 3955
rect 6639 3836 6672 3869
rect 6672 3836 6673 3869
rect 6741 3836 6774 3869
rect 6774 3836 6775 3869
rect 6842 3836 6876 3869
rect 6639 3835 6673 3836
rect 6741 3835 6775 3836
rect 6842 3835 6876 3836
rect 6746 3640 6780 3663
rect 6746 3629 6780 3640
rect 6746 3557 6780 3591
rect 7398 4380 7432 4414
rect 7398 4334 7432 4342
rect 7398 4308 7432 4334
rect 7222 3897 7256 3931
rect 6990 3836 7013 3869
rect 7013 3836 7024 3869
rect 6990 3835 7024 3836
rect 7062 3835 7096 3869
rect 7222 3825 7256 3859
rect 7098 3640 7132 3663
rect 7098 3629 7132 3640
rect 7098 3557 7132 3591
rect 7308 4040 7342 4074
rect 7308 3968 7342 4002
rect 7539 3921 7573 3955
rect 7750 4380 7784 4414
rect 7750 4334 7784 4342
rect 7750 4308 7784 4334
rect 7611 3921 7645 3955
rect 7434 3835 7468 3869
rect 7506 3836 7523 3869
rect 7523 3836 7540 3869
rect 7506 3835 7540 3836
rect 7398 3640 7432 3663
rect 7398 3629 7432 3640
rect 7398 3557 7432 3591
rect 7890 3921 7924 3955
rect 8102 4380 8136 4414
rect 8102 4334 8136 4342
rect 8102 4308 8136 4334
rect 7962 3921 7996 3955
rect 7643 3835 7677 3869
rect 7745 3835 7779 3869
rect 7846 3835 7880 3869
rect 7750 3640 7784 3663
rect 7750 3629 7784 3640
rect 7750 3557 7784 3591
rect 8578 4380 8612 4414
rect 8578 4334 8612 4342
rect 8578 4308 8612 4334
rect 8486 3958 8520 3992
rect 8013 3836 8045 3870
rect 8045 3836 8047 3870
rect 8013 3768 8045 3798
rect 8045 3768 8047 3798
rect 8312 3870 8346 3872
rect 8226 3830 8260 3864
rect 8013 3764 8047 3768
rect 8226 3758 8260 3792
rect 8312 3838 8346 3870
rect 8312 3768 8346 3800
rect 8312 3766 8346 3768
rect 8102 3640 8136 3663
rect 8102 3629 8136 3640
rect 8102 3557 8136 3591
rect 8226 3640 8260 3663
rect 8226 3629 8260 3640
rect 8226 3557 8260 3591
rect 8666 4115 8700 4149
rect 8666 4043 8700 4077
rect 8486 3886 8520 3920
rect 9014 4196 9048 4230
rect 9014 4124 9048 4158
rect 8754 3838 8788 3872
rect 8754 3766 8788 3800
rect 8578 3640 8612 3663
rect 8578 3629 8612 3640
rect 8578 3557 8612 3591
rect 8930 3640 8964 3663
rect 8930 3629 8964 3640
rect 8930 3557 8964 3591
rect 507 3472 519 3506
rect 519 3472 541 3506
rect 579 3472 587 3506
rect 587 3472 613 3506
rect 651 3472 655 3506
rect 655 3472 685 3506
rect 723 3472 757 3506
rect 795 3472 825 3506
rect 825 3472 829 3506
rect 867 3472 893 3506
rect 893 3472 901 3506
rect 939 3472 961 3506
rect 961 3472 973 3506
rect 1011 3472 1029 3506
rect 1029 3472 1045 3506
rect 1083 3472 1097 3506
rect 1097 3472 1117 3506
rect 1155 3472 1165 3506
rect 1165 3472 1189 3506
rect 1227 3472 1233 3506
rect 1233 3472 1261 3506
rect 1299 3472 1301 3506
rect 1301 3472 1333 3506
rect 1371 3472 1403 3506
rect 1403 3472 1405 3506
rect 1443 3472 1471 3506
rect 1471 3472 1477 3506
rect 1515 3472 1539 3506
rect 1539 3472 1549 3506
rect 1587 3472 1607 3506
rect 1607 3472 1621 3506
rect 1659 3472 1675 3506
rect 1675 3472 1693 3506
rect 1731 3472 1743 3506
rect 1743 3472 1765 3506
rect 1803 3472 1811 3506
rect 1811 3472 1837 3506
rect 1875 3472 1879 3506
rect 1879 3472 1909 3506
rect 1947 3472 1981 3506
rect 2019 3472 2049 3506
rect 2049 3472 2053 3506
rect 2091 3472 2117 3506
rect 2117 3472 2125 3506
rect 2163 3472 2185 3506
rect 2185 3472 2197 3506
rect 2235 3472 2253 3506
rect 2253 3472 2269 3506
rect 2307 3472 2321 3506
rect 2321 3472 2341 3506
rect 2379 3472 2389 3506
rect 2389 3472 2413 3506
rect 2451 3472 2457 3506
rect 2457 3472 2485 3506
rect 2523 3472 2525 3506
rect 2525 3472 2557 3506
rect 2595 3472 2627 3506
rect 2627 3472 2629 3506
rect 2667 3472 2695 3506
rect 2695 3472 2701 3506
rect 2739 3472 2763 3506
rect 2763 3472 2773 3506
rect 2811 3472 2831 3506
rect 2831 3472 2845 3506
rect 2883 3472 2899 3506
rect 2899 3472 2917 3506
rect 2955 3472 2967 3506
rect 2967 3472 2989 3506
rect 3027 3472 3035 3506
rect 3035 3472 3061 3506
rect 3099 3472 3103 3506
rect 3103 3472 3133 3506
rect 3171 3472 3205 3506
rect 3243 3472 3273 3506
rect 3273 3472 3277 3506
rect 3315 3472 3341 3506
rect 3341 3472 3349 3506
rect 3387 3472 3409 3506
rect 3409 3472 3421 3506
rect 3459 3472 3477 3506
rect 3477 3472 3493 3506
rect 3531 3472 3545 3506
rect 3545 3472 3565 3506
rect 3603 3472 3613 3506
rect 3613 3472 3637 3506
rect 3675 3472 3681 3506
rect 3681 3472 3709 3506
rect 3747 3472 3749 3506
rect 3749 3472 3781 3506
rect 3819 3472 3851 3506
rect 3851 3472 3853 3506
rect 3891 3472 3919 3506
rect 3919 3472 3925 3506
rect 3963 3472 3987 3506
rect 3987 3472 3997 3506
rect 4035 3472 4055 3506
rect 4055 3472 4069 3506
rect 4107 3472 4123 3506
rect 4123 3472 4141 3506
rect 4179 3472 4191 3506
rect 4191 3472 4213 3506
rect 4251 3472 4259 3506
rect 4259 3472 4285 3506
rect 4323 3472 4327 3506
rect 4327 3472 4357 3506
rect 4395 3472 4429 3506
rect 4467 3472 4497 3506
rect 4497 3472 4501 3506
rect 4539 3472 4565 3506
rect 4565 3472 4573 3506
rect 4611 3472 4633 3506
rect 4633 3472 4645 3506
rect 4683 3472 4701 3506
rect 4701 3472 4717 3506
rect 4755 3472 4769 3506
rect 4769 3472 4789 3506
rect 4827 3472 4837 3506
rect 4837 3472 4861 3506
rect 4899 3472 4905 3506
rect 4905 3472 4933 3506
rect 4971 3472 4973 3506
rect 4973 3472 5005 3506
rect 5043 3472 5075 3506
rect 5075 3472 5077 3506
rect 5115 3472 5143 3506
rect 5143 3472 5149 3506
rect 5187 3472 5211 3506
rect 5211 3472 5221 3506
rect 5259 3472 5279 3506
rect 5279 3472 5293 3506
rect 5331 3472 5347 3506
rect 5347 3472 5365 3506
rect 5403 3472 5415 3506
rect 5415 3472 5437 3506
rect 5475 3472 5483 3506
rect 5483 3472 5509 3506
rect 5547 3472 5551 3506
rect 5551 3472 5581 3506
rect 5619 3472 5653 3506
rect 5691 3472 5721 3506
rect 5721 3472 5725 3506
rect 5763 3472 5789 3506
rect 5789 3472 5797 3506
rect 5835 3472 5857 3506
rect 5857 3472 5869 3506
rect 5907 3472 5925 3506
rect 5925 3472 5941 3506
rect 5979 3472 5993 3506
rect 5993 3472 6013 3506
rect 6051 3472 6061 3506
rect 6061 3472 6085 3506
rect 6123 3472 6129 3506
rect 6129 3472 6157 3506
rect 6195 3472 6197 3506
rect 6197 3472 6229 3506
rect 6267 3472 6299 3506
rect 6299 3472 6301 3506
rect 6339 3472 6367 3506
rect 6367 3472 6373 3506
rect 6411 3472 6435 3506
rect 6435 3472 6445 3506
rect 6483 3472 6503 3506
rect 6503 3472 6517 3506
rect 6555 3472 6571 3506
rect 6571 3472 6589 3506
rect 6627 3472 6639 3506
rect 6639 3472 6661 3506
rect 6699 3472 6707 3506
rect 6707 3472 6733 3506
rect 6771 3472 6775 3506
rect 6775 3472 6805 3506
rect 6843 3472 6877 3506
rect 6915 3472 6945 3506
rect 6945 3472 6949 3506
rect 6987 3472 7013 3506
rect 7013 3472 7021 3506
rect 7059 3472 7081 3506
rect 7081 3472 7093 3506
rect 7131 3472 7149 3506
rect 7149 3472 7165 3506
rect 7203 3472 7217 3506
rect 7217 3472 7237 3506
rect 7275 3472 7285 3506
rect 7285 3472 7309 3506
rect 7347 3472 7353 3506
rect 7353 3472 7381 3506
rect 7419 3472 7421 3506
rect 7421 3472 7453 3506
rect 7491 3472 7523 3506
rect 7523 3472 7525 3506
rect 7563 3472 7591 3506
rect 7591 3472 7597 3506
rect 7635 3472 7659 3506
rect 7659 3472 7669 3506
rect 7707 3472 7727 3506
rect 7727 3472 7741 3506
rect 7779 3472 7795 3506
rect 7795 3472 7813 3506
rect 7851 3472 7863 3506
rect 7863 3472 7885 3506
rect 7923 3472 7931 3506
rect 7931 3472 7957 3506
rect 7995 3472 7999 3506
rect 7999 3472 8029 3506
rect 8067 3472 8101 3506
rect 8139 3472 8169 3506
rect 8169 3472 8173 3506
rect 8211 3472 8237 3506
rect 8237 3472 8245 3506
rect 8283 3472 8305 3506
rect 8305 3472 8317 3506
rect 8355 3472 8373 3506
rect 8373 3472 8389 3506
rect 8427 3472 8441 3506
rect 8441 3472 8461 3506
rect 8499 3472 8509 3506
rect 8509 3472 8533 3506
rect 8571 3472 8577 3506
rect 8577 3472 8605 3506
<< metal1 >>
rect 455 4486 9041 4498
rect 455 4452 467 4486
rect 501 4452 539 4486
rect 573 4452 611 4486
rect 645 4452 683 4486
rect 717 4452 755 4486
rect 789 4452 827 4486
rect 861 4452 899 4486
rect 933 4452 971 4486
rect 1005 4452 1043 4486
rect 1077 4452 1115 4486
rect 1149 4452 1187 4486
rect 1221 4452 1259 4486
rect 1293 4452 1331 4486
rect 1365 4452 1403 4486
rect 1437 4452 1475 4486
rect 1509 4452 1547 4486
rect 1581 4452 1619 4486
rect 1653 4452 1691 4486
rect 1725 4452 1763 4486
rect 1797 4452 1835 4486
rect 1869 4452 1907 4486
rect 1941 4452 1979 4486
rect 2013 4452 2051 4486
rect 2085 4452 2123 4486
rect 2157 4452 2195 4486
rect 2229 4452 2267 4486
rect 2301 4452 2339 4486
rect 2373 4452 2411 4486
rect 2445 4452 2483 4486
rect 2517 4452 2555 4486
rect 2589 4452 2627 4486
rect 2661 4452 2699 4486
rect 2733 4452 2771 4486
rect 2805 4452 2843 4486
rect 2877 4452 2915 4486
rect 2949 4452 2987 4486
rect 3021 4452 3059 4486
rect 3093 4452 3131 4486
rect 3165 4452 3203 4486
rect 3237 4452 3275 4486
rect 3309 4452 3347 4486
rect 3381 4452 3419 4486
rect 3453 4452 3491 4486
rect 3525 4452 3563 4486
rect 3597 4452 3635 4486
rect 3669 4452 3707 4486
rect 3741 4452 3779 4486
rect 3813 4452 3851 4486
rect 3885 4452 3923 4486
rect 3957 4452 3995 4486
rect 4029 4452 4067 4486
rect 4101 4452 4139 4486
rect 4173 4452 4211 4486
rect 4245 4452 4283 4486
rect 4317 4452 4355 4486
rect 4389 4452 4427 4486
rect 4461 4452 4499 4486
rect 4533 4452 4571 4486
rect 4605 4452 4643 4486
rect 4677 4452 4715 4486
rect 4749 4452 4787 4486
rect 4821 4452 4859 4486
rect 4893 4452 4931 4486
rect 4965 4452 5003 4486
rect 5037 4452 5075 4486
rect 5109 4452 5147 4486
rect 5181 4452 5219 4486
rect 5253 4452 5291 4486
rect 5325 4452 5363 4486
rect 5397 4452 5435 4486
rect 5469 4452 5507 4486
rect 5541 4452 5579 4486
rect 5613 4452 5651 4486
rect 5685 4452 5723 4486
rect 5757 4452 5795 4486
rect 5829 4452 5867 4486
rect 5901 4452 5939 4486
rect 5973 4452 6011 4486
rect 6045 4452 6083 4486
rect 6117 4452 6155 4486
rect 6189 4452 6227 4486
rect 6261 4452 6299 4486
rect 6333 4452 6371 4486
rect 6405 4452 6443 4486
rect 6477 4452 6515 4486
rect 6549 4452 6587 4486
rect 6621 4452 6659 4486
rect 6693 4452 6731 4486
rect 6765 4452 6803 4486
rect 6837 4452 6875 4486
rect 6909 4452 6947 4486
rect 6981 4452 7019 4486
rect 7053 4452 7091 4486
rect 7125 4452 7163 4486
rect 7197 4452 7235 4486
rect 7269 4452 7307 4486
rect 7341 4452 7379 4486
rect 7413 4452 7451 4486
rect 7485 4452 7523 4486
rect 7557 4452 7595 4486
rect 7629 4452 7667 4486
rect 7701 4452 7739 4486
rect 7773 4452 7811 4486
rect 7845 4452 7883 4486
rect 7917 4452 7955 4486
rect 7989 4452 8027 4486
rect 8061 4452 8099 4486
rect 8133 4452 8171 4486
rect 8205 4452 8243 4486
rect 8277 4452 8315 4486
rect 8349 4452 8387 4486
rect 8421 4452 8459 4486
rect 8493 4452 8531 4486
rect 8565 4452 8603 4486
rect 8637 4452 8675 4486
rect 8709 4452 8747 4486
rect 8781 4452 8819 4486
rect 8853 4452 8891 4486
rect 8925 4452 9041 4486
rect 455 4440 9041 4452
rect 2571 4414 9041 4440
rect 2571 4380 2802 4414
rect 2836 4380 3154 4414
rect 3188 4380 3278 4414
rect 3312 4380 3578 4414
rect 3612 4380 3930 4414
rect 3964 4380 4282 4414
rect 4316 4380 4634 4414
rect 4668 4380 4986 4414
rect 5020 4380 5338 4414
rect 5372 4380 5690 4414
rect 5724 4380 6042 4414
rect 6076 4380 6394 4414
rect 6428 4380 6746 4414
rect 6780 4380 7098 4414
rect 7132 4380 7398 4414
rect 7432 4380 7750 4414
rect 7784 4380 8102 4414
rect 8136 4380 8578 4414
rect 8612 4380 9041 4414
rect 2571 4342 9041 4380
rect 2571 4308 2802 4342
rect 2836 4308 3154 4342
rect 3188 4308 3278 4342
rect 3312 4308 3578 4342
rect 3612 4308 3930 4342
rect 3964 4308 4282 4342
rect 4316 4308 4634 4342
rect 4668 4308 4986 4342
rect 5020 4308 5338 4342
rect 5372 4308 5690 4342
rect 5724 4308 6042 4342
rect 6076 4308 6394 4342
rect 6428 4308 6746 4342
rect 6780 4308 7098 4342
rect 7132 4308 7398 4342
rect 7432 4308 7750 4342
rect 7784 4308 8102 4342
rect 8136 4308 8578 4342
rect 8612 4308 9041 4342
rect 2571 4295 9041 4308
rect 2619 4198 2665 4210
rect 3684 4201 5050 4253
rect 5102 4201 5114 4253
rect 5166 4201 5172 4253
rect 2619 4164 2625 4198
rect 2659 4164 2665 4198
rect 5874 4196 5880 4248
rect 5932 4196 5944 4248
rect 5996 4242 6002 4248
tri 6002 4242 6008 4248 sw
rect 5996 4230 9054 4242
rect 5996 4196 9014 4230
rect 9048 4196 9054 4230
rect 2619 4158 2665 4164
tri 2665 4158 2703 4196 sw
tri 8974 4167 9003 4196 ne
rect 9003 4167 9054 4196
tri 4791 4161 4797 4167 se
rect 4797 4161 4803 4167
rect 2619 4155 2703 4158
tri 2703 4155 2706 4158 sw
rect 3371 4155 4803 4161
rect 2619 4126 2706 4155
rect 2619 4092 2625 4126
rect 2659 4121 2706 4126
tri 2706 4121 2740 4155 sw
rect 3371 4121 3383 4155
rect 3417 4121 3455 4155
rect 3489 4121 4803 4155
rect 2659 4115 2740 4121
tri 2740 4115 2746 4121 sw
rect 3371 4115 4803 4121
rect 4855 4115 4867 4167
rect 4919 4161 4925 4167
tri 4925 4161 4931 4167 sw
tri 9003 4162 9008 4167 ne
rect 4919 4149 8706 4161
rect 4919 4115 8666 4149
rect 8700 4115 8706 4149
rect 2659 4092 2746 4115
rect 2619 4086 2746 4092
tri 2746 4086 2775 4115 sw
tri 8626 4086 8655 4115 ne
rect 8655 4086 8706 4115
rect 9008 4158 9054 4167
rect 9008 4124 9014 4158
rect 9048 4124 9054 4158
rect 9008 4112 9054 4124
rect 2619 4080 7348 4086
tri 8655 4081 8660 4086 ne
tri 2684 4077 2687 4080 ne
rect 2687 4077 7348 4080
tri 2687 4074 2690 4077 ne
rect 2690 4074 7348 4077
tri 2690 4058 2706 4074 ne
rect 2706 4058 7308 4074
tri 7268 4040 7286 4058 ne
rect 7286 4040 7308 4058
rect 7342 4040 7348 4074
tri 7286 4024 7302 4040 ne
rect 7302 4002 7348 4040
rect 8660 4077 8706 4086
rect 8660 4043 8666 4077
rect 8700 4043 8706 4077
rect 8660 4031 8706 4043
rect 7302 3968 7308 4002
rect 7342 3968 7348 4002
tri 8475 3992 8480 3997 se
rect 8480 3992 8526 4004
tri 3553 3961 3559 3967 sw
tri 5658 3961 5664 3967 se
tri 5792 3961 5798 3967 sw
rect 3552 3915 3701 3961
rect 3703 3955 4352 3961
rect 3703 3921 3719 3955
rect 3753 3921 3791 3955
rect 3825 3921 4070 3955
rect 4104 3921 4142 3955
rect 4176 3921 4352 3955
rect 3703 3915 4352 3921
rect 4446 3955 5608 3961
rect 4446 3921 4458 3955
rect 4492 3921 4530 3955
rect 4564 3921 4774 3955
rect 4808 3921 4846 3955
rect 4880 3921 5126 3955
rect 5160 3921 5198 3955
rect 5232 3921 5479 3955
rect 5513 3921 5551 3955
rect 5585 3921 5608 3955
rect 4446 3915 5608 3921
rect 5613 3915 5806 3961
rect 5811 3955 7005 3961
rect 7302 3956 7348 3968
tri 8444 3961 8475 3992 se
rect 8475 3961 8486 3992
rect 7527 3958 8486 3961
rect 8520 3958 8526 3992
rect 5811 3921 5831 3955
rect 5865 3921 5903 3955
rect 5937 3921 6182 3955
rect 6216 3921 6254 3955
rect 6288 3921 6534 3955
rect 6568 3921 6606 3955
rect 6640 3921 6887 3955
rect 6921 3921 6959 3955
rect 6993 3921 7005 3955
rect 7527 3955 8526 3958
rect 5811 3915 7005 3921
rect 7216 3931 7262 3943
tri 4272 3908 4279 3915 ne
rect 4279 3908 4352 3915
rect 2883 3896 2929 3908
tri 4279 3897 4290 3908 ne
rect 4290 3897 4352 3908
tri 4352 3897 4364 3909 sw
rect 7216 3897 7222 3931
rect 7256 3897 7262 3931
rect 7527 3921 7539 3955
rect 7573 3921 7611 3955
rect 7645 3921 7890 3955
rect 7924 3921 7962 3955
rect 7996 3921 8526 3955
rect 7527 3920 8526 3921
rect 2883 3862 2889 3896
rect 2923 3862 2929 3896
tri 4290 3889 4298 3897 ne
rect 4298 3889 4364 3897
rect 2883 3842 2929 3862
rect 2456 3824 2929 3842
rect 2456 3790 2889 3824
rect 2923 3790 2929 3824
rect 2456 3778 2929 3790
rect 3055 3877 3101 3889
tri 4298 3886 4301 3889 ne
rect 4301 3886 4364 3889
tri 4364 3886 4375 3897 sw
rect 7216 3886 7262 3897
tri 7262 3886 7295 3919 sw
rect 7527 3915 8486 3920
tri 8444 3886 8473 3915 ne
rect 8473 3886 8486 3915
rect 8520 3886 8526 3920
tri 4301 3882 4305 3886 ne
rect 4305 3882 4375 3886
rect 3055 3843 3061 3877
rect 3095 3843 3101 3877
tri 4180 3875 4187 3882 se
rect 4187 3875 4233 3882
tri 4305 3881 4306 3882 ne
rect 3055 3805 3101 3843
rect 3454 3870 4233 3875
rect 3454 3869 4193 3870
rect 3454 3835 3466 3869
rect 3500 3835 3538 3869
rect 3572 3835 3614 3869
rect 3648 3835 3686 3869
rect 3720 3835 3823 3869
rect 3857 3835 3925 3869
rect 3959 3835 4026 3869
rect 4060 3836 4193 3869
rect 4227 3836 4233 3870
rect 4060 3835 4233 3836
rect 3454 3829 4233 3835
rect 4306 3875 4375 3882
tri 4375 3875 4386 3886 sw
rect 7216 3875 7295 3886
tri 7295 3875 7306 3886 sw
tri 8473 3884 8475 3886 ne
rect 8475 3884 8526 3886
tri 8001 3876 8007 3882 se
rect 8007 3876 8053 3882
tri 8000 3875 8001 3876 se
rect 8001 3875 8053 3876
rect 4306 3869 7108 3875
rect 4306 3835 4318 3869
rect 4352 3835 4390 3869
rect 4424 3835 4527 3869
rect 4561 3835 4629 3869
rect 4663 3835 4730 3869
rect 4764 3835 4886 3869
rect 4920 3835 4983 3869
rect 5017 3835 5080 3869
rect 5114 3835 5231 3869
rect 5265 3835 5333 3869
rect 5367 3835 5434 3869
rect 5468 3835 5582 3869
rect 5616 3835 5654 3869
rect 5688 3835 5726 3869
rect 5760 3835 5798 3869
rect 5832 3835 5935 3869
rect 5969 3835 6037 3869
rect 6071 3835 6138 3869
rect 6172 3835 6294 3869
rect 6328 3835 6391 3869
rect 6425 3835 6488 3869
rect 6522 3835 6639 3869
rect 6673 3835 6741 3869
rect 6775 3835 6842 3869
rect 6876 3835 6990 3869
rect 7024 3835 7062 3869
rect 7096 3835 7108 3869
rect 4306 3829 7108 3835
rect 7216 3870 8053 3875
rect 7216 3869 8013 3870
rect 7216 3859 7434 3869
tri 4153 3825 4157 3829 ne
rect 4157 3825 4233 3829
tri 4157 3813 4169 3825 ne
rect 4169 3813 4233 3825
rect 7216 3825 7222 3859
rect 7256 3835 7434 3859
rect 7468 3835 7506 3869
rect 7540 3835 7643 3869
rect 7677 3835 7745 3869
rect 7779 3835 7846 3869
rect 7880 3836 8013 3869
rect 8047 3836 8053 3870
rect 7880 3835 8053 3836
rect 7256 3829 8053 3835
rect 7256 3825 7262 3829
rect 7216 3813 7262 3825
tri 7262 3813 7278 3829 nw
tri 7973 3813 7989 3829 ne
rect 7989 3813 8053 3829
rect 2446 3771 2453 3778
tri 2453 3771 2460 3778 nw
rect 3055 3771 3061 3805
rect 3095 3771 3101 3805
tri 4169 3800 4182 3813 ne
rect 4182 3800 4233 3813
tri 7989 3800 8002 3813 ne
rect 8002 3800 8053 3813
tri 4182 3798 4184 3800 ne
rect 4184 3798 4233 3800
tri 8002 3798 8004 3800 ne
rect 8004 3798 8053 3800
tri 4184 3795 4187 3798 ne
rect 2446 3770 2452 3771
tri 2452 3770 2453 3771 nw
rect 3055 3759 3101 3771
rect 4187 3764 4193 3798
rect 4227 3764 4233 3798
tri 8004 3795 8007 3798 ne
tri 3355 3749 3361 3755 se
rect 3361 3749 3968 3755
rect 2542 3743 2672 3749
rect 2542 3709 2554 3743
rect 2588 3709 2626 3743
rect 2660 3731 2672 3743
tri 2672 3731 2690 3749 sw
tri 3337 3731 3355 3749 se
rect 3355 3731 3968 3749
rect 2660 3709 3968 3731
rect 2542 3703 3968 3709
rect 4020 3703 4032 3755
rect 4084 3703 4090 3755
rect 4187 3752 4233 3764
rect 8007 3764 8013 3798
rect 8047 3764 8053 3798
rect 8007 3752 8053 3764
rect 8217 3870 8269 3876
rect 8217 3804 8269 3818
rect 8306 3872 8352 3884
tri 8475 3879 8480 3884 ne
tri 8352 3872 8356 3876 sw
rect 8480 3874 8526 3884
tri 8746 3874 8748 3876 se
rect 8748 3874 8794 3884
tri 8744 3872 8746 3874 se
rect 8746 3872 8794 3874
rect 8306 3838 8312 3872
rect 8346 3842 8356 3872
tri 8356 3842 8386 3872 sw
tri 8714 3842 8744 3872 se
rect 8744 3842 8754 3872
rect 8346 3838 8754 3842
rect 8788 3838 8794 3872
rect 8306 3800 8794 3838
rect 8306 3766 8312 3800
rect 8346 3796 8754 3800
rect 8346 3766 8356 3796
tri 8356 3766 8386 3796 nw
tri 8714 3766 8744 3796 ne
rect 8744 3766 8754 3796
rect 8788 3766 8794 3800
rect 8306 3754 8352 3766
tri 8352 3762 8356 3766 nw
tri 8744 3762 8748 3766 ne
rect 8748 3754 8794 3766
rect 8217 3746 8269 3752
rect 2571 3663 9000 3675
rect 2571 3629 2802 3663
rect 2836 3629 3278 3663
rect 3312 3629 3578 3663
rect 3612 3629 3930 3663
rect 3964 3629 4282 3663
rect 4316 3629 4634 3663
rect 4668 3629 4986 3663
rect 5020 3629 5338 3663
rect 5372 3629 5690 3663
rect 5724 3629 6042 3663
rect 6076 3629 6394 3663
rect 6428 3629 6746 3663
rect 6780 3629 7098 3663
rect 7132 3629 7398 3663
rect 7432 3629 7750 3663
rect 7784 3629 8102 3663
rect 8136 3629 8226 3663
rect 8260 3629 8578 3663
rect 8612 3629 8930 3663
rect 8964 3629 9000 3663
rect 2571 3591 9000 3629
rect 2571 3557 2802 3591
rect 2836 3557 3278 3591
rect 3312 3557 3578 3591
rect 3612 3557 3930 3591
rect 3964 3557 4282 3591
rect 4316 3557 4634 3591
rect 4668 3557 4986 3591
rect 5020 3557 5338 3591
rect 5372 3557 5690 3591
rect 5724 3557 6042 3591
rect 6076 3557 6394 3591
rect 6428 3557 6746 3591
rect 6780 3557 7098 3591
rect 7132 3557 7398 3591
rect 7432 3557 7750 3591
rect 7784 3557 8102 3591
rect 8136 3557 8226 3591
rect 8260 3557 8578 3591
rect 8612 3557 8930 3591
rect 8964 3557 9000 3591
rect 2571 3518 9000 3557
rect 495 3506 9000 3518
rect 495 3472 507 3506
rect 541 3472 579 3506
rect 613 3472 651 3506
rect 685 3472 723 3506
rect 757 3472 795 3506
rect 829 3472 867 3506
rect 901 3472 939 3506
rect 973 3472 1011 3506
rect 1045 3472 1083 3506
rect 1117 3472 1155 3506
rect 1189 3472 1227 3506
rect 1261 3472 1299 3506
rect 1333 3472 1371 3506
rect 1405 3472 1443 3506
rect 1477 3472 1515 3506
rect 1549 3472 1587 3506
rect 1621 3472 1659 3506
rect 1693 3472 1731 3506
rect 1765 3472 1803 3506
rect 1837 3472 1875 3506
rect 1909 3472 1947 3506
rect 1981 3472 2019 3506
rect 2053 3472 2091 3506
rect 2125 3472 2163 3506
rect 2197 3472 2235 3506
rect 2269 3472 2307 3506
rect 2341 3472 2379 3506
rect 2413 3472 2451 3506
rect 2485 3472 2523 3506
rect 2557 3472 2595 3506
rect 2629 3472 2667 3506
rect 2701 3472 2739 3506
rect 2773 3472 2811 3506
rect 2845 3472 2883 3506
rect 2917 3472 2955 3506
rect 2989 3472 3027 3506
rect 3061 3472 3099 3506
rect 3133 3472 3171 3506
rect 3205 3472 3243 3506
rect 3277 3472 3315 3506
rect 3349 3472 3387 3506
rect 3421 3472 3459 3506
rect 3493 3472 3531 3506
rect 3565 3472 3603 3506
rect 3637 3472 3675 3506
rect 3709 3472 3747 3506
rect 3781 3472 3819 3506
rect 3853 3472 3891 3506
rect 3925 3472 3963 3506
rect 3997 3472 4035 3506
rect 4069 3472 4107 3506
rect 4141 3472 4179 3506
rect 4213 3472 4251 3506
rect 4285 3472 4323 3506
rect 4357 3472 4395 3506
rect 4429 3472 4467 3506
rect 4501 3472 4539 3506
rect 4573 3472 4611 3506
rect 4645 3472 4683 3506
rect 4717 3472 4755 3506
rect 4789 3472 4827 3506
rect 4861 3472 4899 3506
rect 4933 3472 4971 3506
rect 5005 3472 5043 3506
rect 5077 3472 5115 3506
rect 5149 3472 5187 3506
rect 5221 3472 5259 3506
rect 5293 3472 5331 3506
rect 5365 3472 5403 3506
rect 5437 3472 5475 3506
rect 5509 3472 5547 3506
rect 5581 3472 5619 3506
rect 5653 3472 5691 3506
rect 5725 3472 5763 3506
rect 5797 3472 5835 3506
rect 5869 3472 5907 3506
rect 5941 3472 5979 3506
rect 6013 3472 6051 3506
rect 6085 3472 6123 3506
rect 6157 3472 6195 3506
rect 6229 3472 6267 3506
rect 6301 3472 6339 3506
rect 6373 3472 6411 3506
rect 6445 3472 6483 3506
rect 6517 3472 6555 3506
rect 6589 3472 6627 3506
rect 6661 3472 6699 3506
rect 6733 3472 6771 3506
rect 6805 3472 6843 3506
rect 6877 3472 6915 3506
rect 6949 3472 6987 3506
rect 7021 3472 7059 3506
rect 7093 3472 7131 3506
rect 7165 3472 7203 3506
rect 7237 3472 7275 3506
rect 7309 3472 7347 3506
rect 7381 3472 7419 3506
rect 7453 3472 7491 3506
rect 7525 3472 7563 3506
rect 7597 3472 7635 3506
rect 7669 3472 7707 3506
rect 7741 3472 7779 3506
rect 7813 3472 7851 3506
rect 7885 3472 7923 3506
rect 7957 3472 7995 3506
rect 8029 3472 8067 3506
rect 8101 3472 8139 3506
rect 8173 3472 8211 3506
rect 8245 3472 8283 3506
rect 8317 3472 8355 3506
rect 8389 3472 8427 3506
rect 8461 3472 8499 3506
rect 8533 3472 8571 3506
rect 8605 3472 9000 3506
rect 495 3460 9000 3472
rect 5044 3215 5050 3267
rect 5102 3215 5114 3267
rect 5166 3215 5172 3267
rect 4118 2623 4170 2629
tri 4082 2553 4118 2589 se
rect 4671 2610 4723 2616
rect 4118 2559 4170 2571
tri 4170 2553 4200 2583 sw
tri 5797 2586 5803 2592 se
rect 4118 2501 4170 2507
rect 4671 2540 4723 2558
rect 5803 2540 5809 2592
rect 5861 2540 5873 2592
rect 5925 2540 5931 2592
tri 5931 2586 5937 2592 sw
rect 4671 2482 4723 2488
tri 4097 1871 4131 1905 ne
rect 4131 1810 4183 1905
tri 4183 1871 4217 1905 nw
tri 4322 1607 4331 1616 se
rect 4331 1607 4377 1648
rect 4088 1601 4140 1607
tri 4300 1585 4322 1607 se
rect 4322 1596 4377 1607
rect 4322 1585 4336 1596
tri 4140 1555 4170 1585 sw
tri 4270 1555 4300 1585 se
rect 4300 1555 4336 1585
tri 4336 1555 4377 1596 nw
rect 4140 1549 4290 1555
rect 4088 1537 4290 1549
rect 4140 1509 4290 1537
tri 4290 1509 4336 1555 nw
rect 4088 1479 4140 1485
tri 4140 1479 4170 1509 nw
rect 4824 1247 5182 1360
<< rmetal1 >>
rect 3701 3915 3703 3961
rect 5608 3915 5613 3961
rect 5806 3915 5811 3961
<< via1 >>
rect 5050 4201 5102 4253
rect 5114 4201 5166 4253
rect 5880 4196 5932 4248
rect 5944 4196 5996 4248
rect 4803 4115 4855 4167
rect 4867 4115 4919 4167
rect 3968 3703 4020 3755
rect 4032 3703 4084 3755
rect 8217 3864 8269 3870
rect 8217 3830 8226 3864
rect 8226 3830 8260 3864
rect 8260 3830 8269 3864
rect 8217 3818 8269 3830
rect 8217 3792 8269 3804
rect 8217 3758 8226 3792
rect 8226 3758 8260 3792
rect 8260 3758 8269 3792
rect 8217 3752 8269 3758
rect 5050 3215 5102 3267
rect 5114 3215 5166 3267
rect 4118 2571 4170 2623
rect 4118 2507 4170 2559
rect 4671 2558 4723 2610
rect 5809 2540 5861 2592
rect 5873 2540 5925 2592
rect 4671 2488 4723 2540
rect 4088 1549 4140 1601
rect 4088 1485 4140 1537
<< metal2 >>
tri 3556 4196 3561 4201 ne
rect 3561 4196 3614 4201
tri 3561 4167 3590 4196 ne
rect 3590 4167 3614 4196
rect 3665 4196 3679 4201
tri 3679 4196 3684 4201 nw
tri 3665 4182 3679 4196 nw
tri 3590 4143 3614 4167 ne
rect 4110 4025 4162 4213
rect 5044 4201 5050 4253
rect 5102 4201 5114 4253
rect 5166 4201 5172 4253
tri 5044 4196 5049 4201 ne
rect 5049 4196 5156 4201
tri 5156 4196 5161 4201 nw
rect 5874 4196 5880 4248
rect 5932 4196 5944 4248
rect 5996 4196 6002 4248
tri 5049 4170 5075 4196 ne
rect 4797 4115 4803 4167
rect 4855 4115 4867 4167
rect 4919 4115 4925 4167
tri 4162 4025 4170 4033 sw
rect 4110 4011 4170 4025
tri 4110 4003 4118 4011 ne
rect 3962 3703 3968 3755
rect 4020 3703 4032 3755
rect 4084 3703 4090 3755
tri 3983 3648 4038 3703 ne
rect 4038 2399 4090 3703
rect 4118 2623 4170 4011
tri 4787 3818 4797 3828 se
rect 4797 3818 4851 4115
tri 4851 4081 4885 4115 nw
tri 4773 3804 4787 3818 se
rect 4787 3804 4851 3818
tri 4744 3775 4773 3804 se
rect 4773 3775 4851 3804
rect 4744 3723 4851 3775
rect 4118 2559 4170 2571
rect 4118 2501 4170 2507
tri 4671 2773 4744 2846 se
rect 4744 2824 4796 3723
tri 4796 3668 4851 3723 nw
tri 5044 3267 5075 3298 se
rect 5075 3267 5127 4196
tri 5127 4167 5156 4196 nw
tri 5875 4167 5904 4196 ne
rect 5904 4167 5962 4196
tri 5904 4161 5910 4167 ne
tri 5127 3267 5161 3301 sw
rect 5044 3215 5050 3267
rect 5102 3215 5114 3267
rect 5166 3215 5172 3267
rect 4744 2773 4745 2824
tri 4745 2773 4796 2824 nw
tri 5844 2857 5910 2923 se
rect 5910 2901 5962 4167
tri 5962 4161 5997 4196 nw
rect 8217 3870 8269 3876
rect 8217 3804 8269 3818
rect 8217 3746 8269 3752
rect 5910 2857 5918 2901
tri 5918 2857 5962 2901 nw
rect 4671 2610 4723 2773
tri 4723 2751 4745 2773 nw
tri 5809 2592 5844 2627 se
rect 5844 2592 5896 2857
tri 5896 2835 5918 2857 nw
tri 5896 2592 5931 2627 sw
rect 4671 2540 4723 2558
rect 5803 2540 5809 2592
rect 5861 2540 5873 2592
rect 5925 2540 5931 2592
rect 4671 2482 4723 2488
tri 4038 2349 4088 2399 ne
rect 4088 2371 4090 2399
tri 4090 2371 4140 2421 sw
rect 4088 1601 4140 2371
rect 4088 1537 4140 1549
rect 4088 1479 4140 1485
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_0
timestamp 1704896540
transform -1 0 6098 0 -1 3226
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1704896540
transform -1 0 2910 0 1 3436
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1704896540
transform -1 0 7506 0 1 3436
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1704896540
transform 1 0 3204 0 1 3436
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x4  sky130_fd_io__hvsbt_inv_x4_0
timestamp 1704896540
transform 1 0 7324 0 1 3436
box 107 226 812 873
use sky130_fd_io__hvsbt_inv_x4  sky130_fd_io__hvsbt_inv_x4_1
timestamp 1704896540
transform 1 0 3504 0 1 3436
box 107 226 812 873
use sky130_fd_io__hvsbt_inv_x8  sky130_fd_io__hvsbt_inv_x8_0
timestamp 1704896540
transform 1 0 5616 0 1 3436
box 107 226 1516 873
use sky130_fd_io__hvsbt_inv_x8v2  sky130_fd_io__hvsbt_inv_x8v2_0
timestamp 1704896540
transform 1 0 4208 0 1 3436
box 107 226 1516 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1704896540
transform 1 0 2728 0 1 3436
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1704896540
transform 1 0 8504 0 1 3436
box 107 226 460 873
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1704896540
transform -1 0 8686 0 1 3436
box 107 226 460 873
<< labels >>
flabel metal2 s 4128 4183 4156 4207 3 FreeSans 520 0 0 0 HLD_OVR
port 1 nsew
flabel metal1 s 5581 2998 5581 2998 0 FreeSans 440 0 0 0 VCC_IO
flabel metal1 s 2709 4335 2832 4438 3 FreeSans 520 0 0 0 VCC_IO
port 3 nsew
flabel metal1 s 2754 3479 2929 3557 3 FreeSans 520 0 0 0 VGND
port 4 nsew
flabel metal1 s 5639 3921 5793 3954 3 FreeSans 520 0 0 0 HLD_I_H_N
port 5 nsew
flabel metal1 s 8026 3927 8091 3951 3 FreeSans 520 0 0 0 OD_I_H
port 6 nsew
flabel metal1 s 5725 1995 5725 1995 0 FreeSans 440 0 0 0 VGND
flabel metal1 s 5699 2830 5699 2830 0 FreeSans 440 0 0 0 VPWR
flabel metal1 s 4824 1247 5182 1360 3 FreeSans 520 0 0 0 VPWR
port 7 nsew
flabel metal1 s 3552 3915 3606 3961 3 FreeSans 520 0 0 0 HLD_I_H
port 8 nsew
<< properties >>
string GDS_END 21655858
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21611784
<< end >>
