magic
tech sky130A
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_0
timestamp 1704896540
transform 1 0 800 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_1
timestamp 1704896540
transform 1 0 2512 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_2
timestamp 1704896540
transform 1 0 4224 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_3
timestamp 1704896540
transform 1 0 5936 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_4
timestamp 1704896540
transform 1 0 7648 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_55959141808666  sky130_fd_pr__dfl1sd2__example_55959141808666_5
timestamp 1704896540
transform 1 0 9360 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_0
timestamp 1704896540
transform 1 0 1656 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_1
timestamp 1704896540
transform 1 0 3368 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_2
timestamp 1704896540
transform 1 0 5080 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_3
timestamp 1704896540
transform 1 0 6792 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808337  sky130_fd_pr__hvdfl1sd2__example_55959141808337_4
timestamp 1704896540
transform 1 0 8504 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808338  sky130_fd_pr__hvdfl1sd__example_55959141808338_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808338  sky130_fd_pr__hvdfl1sd__example_55959141808338_1
timestamp 1704896540
transform 1 0 10216 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 58043050
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 58036310
<< end >>
