magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< comment >>
rect 0 23025 60 23759
rect 14940 23025 15000 23759
rect 0 19801 60 22865
rect 14940 19801 15000 22865
rect 0 18832 60 19641
rect 14940 18832 15000 19641
rect 0 17441 60 18672
rect 14940 17441 15000 18672
rect 0 13739 60 17281
rect 14940 13739 15000 17281
rect 0 12381 60 13579
rect 14940 12381 15000 13579
rect 0 11023 60 12221
rect 14940 11023 15000 12221
rect 0 9665 60 10863
rect 14940 9665 15000 10863
rect 0 8307 60 9505
rect 14940 8307 15000 9505
rect 0 6949 60 8147
rect 14940 6949 15000 8147
rect 0 5512 60 6789
rect 14940 5512 15000 6789
rect 0 4154 60 5352
rect 14940 4154 15000 5352
rect 0 2796 60 3994
rect 14940 2796 15000 3994
rect 0 1438 60 2636
rect 14940 1438 15000 2636
rect 0 80 60 1278
rect 14940 80 15000 1278
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_0
timestamp 1704896540
transform 1 0 14000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_1
timestamp 1704896540
transform 1 0 13000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_2
timestamp 1704896540
transform 1 0 12000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_3
timestamp 1704896540
transform 1 0 11000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_4
timestamp 1704896540
transform 1 0 10000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_5
timestamp 1704896540
transform 1 0 9000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_6
timestamp 1704896540
transform 1 0 8000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_7
timestamp 1704896540
transform 1 0 7000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_8
timestamp 1704896540
transform 1 0 6000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_9
timestamp 1704896540
transform 1 0 15000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_10
timestamp 1704896540
transform 1 0 0 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_11
timestamp 1704896540
transform 1 0 5000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_12
timestamp 1704896540
transform 1 0 4000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_13
timestamp 1704896540
transform 1 0 3000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_14
timestamp 1704896540
transform 1 0 16000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_15
timestamp 1704896540
transform 1 0 2000 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_16
timestamp 1704896540
transform 1 0 1000 0 1 0
box 0 250 1000 13599
<< labels >>
flabel comment s 14940 80 15000 1278 7 FreeSans 4000 0 0 0 vpb_ka
port 1 nsew
flabel comment s 14940 4154 15000 5352 7 FreeSans 4000 0 0 0 vcc_ioq
port 2 nsew
flabel comment s 14940 2796 15000 3994 7 FreeSans 4000 0 0 0 vgnd
port 3 nsew
flabel comment s 14940 1438 15000 2636 7 FreeSans 4000 0 0 0 vpwr_ka
port 4 nsew
flabel comment s 14940 13739 15000 17281 7 FreeSans 4000 0 0 0 vgnd_io
port 5 nsew
flabel comment s 14940 17441 15000 18672 7 FreeSans 4000 0 0 0 vcc_io
port 6 nsew
flabel comment s 14940 12381 15000 13579 7 FreeSans 4000 0 0 0 vcc_io
port 6 nsew
flabel comment s 14940 5512 15000 6789 7 FreeSans 4000 0 0 0 vgnd
port 3 nsew
flabel comment s 0 8307 60 9505 7 FreeSans 4000 180 0 0 vpb
port 7 nsew
flabel comment s 14940 19801 15000 22865 7 FreeSans 4000 0 0 0 vgnd_io
port 5 nsew
flabel comment s 0 6949 60 8147 7 FreeSans 4000 180 0 0 vcc_ioq
port 2 nsew
flabel comment s 0 9665 60 10863 7 FreeSans 4000 180 0 0 vpwr
port 8 nsew
flabel comment s 0 11023 60 12221 7 FreeSans 4000 180 0 0 vgnd
port 3 nsew
flabel comment s 0 19801 60 22865 7 FreeSans 4000 180 0 0 vgnd_io
port 5 nsew
flabel comment s 0 5512 60 6789 7 FreeSans 4000 180 0 0 vgnd
port 3 nsew
flabel comment s 0 13739 60 17281 7 FreeSans 4000 180 0 0 vgnd_io
port 5 nsew
flabel comment s 0 12381 60 13579 7 FreeSans 4000 180 0 0 vcc_io
port 6 nsew
flabel comment s 14940 11023 15000 12221 7 FreeSans 4000 0 0 0 vgnd
port 3 nsew
flabel comment s 0 2796 60 3994 7 FreeSans 4000 180 0 0 vgnd
port 3 nsew
flabel comment s 0 1438 60 2636 7 FreeSans 4000 180 0 0 vpwr_ka
port 4 nsew
flabel comment s 0 4154 60 5352 7 FreeSans 4000 180 0 0 vcc_ioq
port 2 nsew
flabel comment s 0 80 60 1278 7 FreeSans 4000 180 0 0 vpb_ka
port 1 nsew
flabel comment s 0 23025 60 23759 3 FreeSans 4000 0 0 0 vssio_amx
port 9 nsew
flabel comment s 14940 8307 15000 9505 7 FreeSans 4000 0 0 0 vpb
port 7 nsew
flabel comment s 14940 9665 15000 10863 7 FreeSans 4000 0 0 0 vpwr
port 8 nsew
flabel comment s 14940 6949 15000 8147 7 FreeSans 4000 0 0 0 vcc_ioq
port 2 nsew
flabel comment s 14940 23025 15000 23759 7 FreeSans 4000 0 0 0 vssio_amx
port 9 nsew
flabel comment s 14940 18832 15000 19641 7 FreeSans 4000 0 0 0 vio_amx
port 10 nsew
flabel comment s 0 18832 60 19641 3 FreeSans 4000 0 0 0 vio_amx
port 10 nsew
flabel comment s 0 17441 60 18672 7 FreeSans 4000 180 0 0 vcc_io
port 6 nsew
<< properties >>
string GDS_END 85514706
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85509750
<< end >>
