magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -105 -26 607 2026
rect 815 -26 1527 2026
rect 1735 -26 2447 2026
rect 2655 -26 3367 2026
rect 3575 -26 4287 2026
rect 4495 -26 5207 2026
rect 5415 -26 6127 2026
rect 6335 -26 7047 2026
rect 7255 -26 7967 2026
rect 8175 -26 8887 2026
rect 9095 -26 9807 2026
<< mvnmos >>
rect 0 0 100 2000
rect 402 0 502 2000
rect 920 0 1020 2000
rect 1322 0 1422 2000
rect 1840 0 1940 2000
rect 2242 0 2342 2000
rect 2760 0 2860 2000
rect 3162 0 3262 2000
rect 3680 0 3780 2000
rect 4082 0 4182 2000
rect 4600 0 4700 2000
rect 5002 0 5102 2000
rect 5520 0 5620 2000
rect 5922 0 6022 2000
rect 6440 0 6540 2000
rect 6842 0 6942 2000
rect 7360 0 7460 2000
rect 7762 0 7862 2000
rect 8280 0 8380 2000
rect 8682 0 8782 2000
rect 9200 0 9300 2000
rect 9602 0 9702 2000
<< mvndiff >>
rect -79 0 0 2000
rect 100 0 402 2000
rect 502 0 581 2000
rect 841 0 920 2000
rect 1020 0 1322 2000
rect 1422 0 1501 2000
rect 1761 0 1840 2000
rect 1940 0 2242 2000
rect 2342 0 2421 2000
rect 2681 0 2760 2000
rect 2860 0 3162 2000
rect 3262 0 3341 2000
rect 3601 0 3680 2000
rect 3780 0 4082 2000
rect 4182 0 4261 2000
rect 4521 0 4600 2000
rect 4700 0 5002 2000
rect 5102 0 5181 2000
rect 5441 0 5520 2000
rect 5620 0 5922 2000
rect 6022 0 6101 2000
rect 6361 0 6440 2000
rect 6540 0 6842 2000
rect 6942 0 7021 2000
rect 7281 0 7360 2000
rect 7460 0 7762 2000
rect 7862 0 7941 2000
rect 8201 0 8280 2000
rect 8380 0 8682 2000
rect 8782 0 8861 2000
rect 9121 0 9200 2000
rect 9300 0 9602 2000
rect 9702 0 9781 2000
<< poly >>
rect 0 2000 100 2032
rect 402 2000 502 2032
rect 920 2000 1020 2032
rect 1322 2000 1422 2032
rect 1840 2000 1940 2032
rect 2242 2000 2342 2032
rect 2760 2000 2860 2032
rect 3162 2000 3262 2032
rect 3680 2000 3780 2032
rect 4082 2000 4182 2032
rect 4600 2000 4700 2032
rect 5002 2000 5102 2032
rect 5520 2000 5620 2032
rect 5922 2000 6022 2032
rect 6440 2000 6540 2032
rect 6842 2000 6942 2032
rect 7360 2000 7460 2032
rect 7762 2000 7862 2032
rect 8280 2000 8380 2032
rect 8682 2000 8782 2032
rect 9200 2000 9300 2032
rect 9602 2000 9702 2032
rect 0 -32 100 0
rect 402 -32 502 0
rect 920 -32 1020 0
rect 1322 -32 1422 0
rect 1840 -32 1940 0
rect 2242 -32 2342 0
rect 2760 -32 2860 0
rect 3162 -32 3262 0
rect 3680 -32 3780 0
rect 4082 -32 4182 0
rect 4600 -32 4700 0
rect 5002 -32 5102 0
rect 5520 -32 5620 0
rect 5922 -32 6022 0
rect 6440 -32 6540 0
rect 6842 -32 6942 0
rect 7360 -32 7460 0
rect 7762 -32 7862 0
rect 8280 -32 8380 0
rect 8682 -32 8782 0
rect 9200 -32 9300 0
rect 9602 -32 9702 0
<< locali >>
rect -192 -4 -90 1978
rect 592 -4 830 1966
rect 1512 -4 1750 1966
rect 2432 -4 2670 1966
rect 3352 -4 3590 1966
rect 4272 -4 4510 1966
rect 5192 -4 5430 1966
rect 6112 -4 6350 1966
rect 7032 -4 7270 1966
rect 7952 -4 8190 1966
rect 8872 -4 9110 1966
rect 9792 -4 9894 1978
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_0
timestamp 1704896540
transform 1 0 8861 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_1
timestamp 1704896540
transform 1 0 7941 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_2
timestamp 1704896540
transform 1 0 7021 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_3
timestamp 1704896540
transform 1 0 6101 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_4
timestamp 1704896540
transform 1 0 5181 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_5
timestamp 1704896540
transform 1 0 4261 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_6
timestamp 1704896540
transform 1 0 3341 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_7
timestamp 1704896540
transform 1 0 2421 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_8
timestamp 1704896540
transform 1 0 1501 0 1 0
box -26 -26 286 2026
use hvDFTPL1s2_CDNS_52468879185836  hvDFTPL1s2_CDNS_52468879185836_9
timestamp 1704896540
transform 1 0 581 0 1 0
box -26 -26 286 2026
use hvDFTPL1s_CDNS_52468879185835  hvDFTPL1s_CDNS_52468879185835_0
timestamp 1704896540
transform -1 0 -79 0 1 0
box -26 -26 226 2026
use hvDFTPL1s_CDNS_52468879185835  hvDFTPL1s_CDNS_52468879185835_1
timestamp 1704896540
transform 1 0 9781 0 1 0
box -26 -26 226 2026
<< labels >>
flabel comment s -141 987 -141 987 0 FreeSans 300 0 0 0 S
flabel comment s 251 1000 251 1000 0 FreeSans 300 0 0 0 D
flabel comment s 711 981 711 981 0 FreeSans 300 0 0 0 S
flabel comment s 1171 1000 1171 1000 0 FreeSans 300 0 0 0 D
flabel comment s 1631 981 1631 981 0 FreeSans 300 0 0 0 S
flabel comment s 2091 1000 2091 1000 0 FreeSans 300 0 0 0 D
flabel comment s 2551 981 2551 981 0 FreeSans 300 0 0 0 S
flabel comment s 3011 1000 3011 1000 0 FreeSans 300 0 0 0 D
flabel comment s 3471 981 3471 981 0 FreeSans 300 0 0 0 S
flabel comment s 3931 1000 3931 1000 0 FreeSans 300 0 0 0 D
flabel comment s 4391 981 4391 981 0 FreeSans 300 0 0 0 S
flabel comment s 4851 1000 4851 1000 0 FreeSans 300 0 0 0 D
flabel comment s 5311 981 5311 981 0 FreeSans 300 0 0 0 S
flabel comment s 5771 1000 5771 1000 0 FreeSans 300 0 0 0 D
flabel comment s 6231 981 6231 981 0 FreeSans 300 0 0 0 S
flabel comment s 6691 1000 6691 1000 0 FreeSans 300 0 0 0 D
flabel comment s 7151 981 7151 981 0 FreeSans 300 0 0 0 S
flabel comment s 7611 1000 7611 1000 0 FreeSans 300 0 0 0 D
flabel comment s 8071 981 8071 981 0 FreeSans 300 0 0 0 S
flabel comment s 8531 1000 8531 1000 0 FreeSans 300 0 0 0 D
flabel comment s 8991 981 8991 981 0 FreeSans 300 0 0 0 S
flabel comment s 9451 1000 9451 1000 0 FreeSans 300 0 0 0 D
flabel comment s 9843 987 9843 987 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 34362424
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34350920
<< end >>
