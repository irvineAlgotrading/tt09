magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 975 1466
<< mvpmos >>
rect 0 0 400 1400
rect 456 0 856 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 856 0 906 1400
<< poly >>
rect 0 1400 400 1426
rect 0 -26 400 0
rect 456 1400 856 1426
rect 456 -26 856 0
<< locali >>
rect 411 -4 445 1354
<< metal1 >>
rect -51 -16 -5 1410
rect 861 -16 907 1410
use DFM1sd_CDNS_524688791851132  DFM1sd_CDNS_524688791851132_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 1436
use DFM1sd_CDNS_524688791851132  DFM1sd_CDNS_524688791851132_1
timestamp 1704896540
transform 1 0 856 0 1 0
box -36 -36 89 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_0
timestamp 1704896540
transform 1 0 400 0 1 0
box -36 -36 92 1436
<< labels >>
flabel comment s -28 697 -28 697 0 FreeSans 300 0 0 0 S
flabel comment s 428 675 428 675 0 FreeSans 300 0 0 0 D
flabel comment s 884 697 884 697 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 78928318
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78926802
<< end >>
