magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -1422 129 -54 3010
rect 3508 129 3678 681
rect -1422 -41 3678 129
<< pwell >>
rect 3172 2319 4089 2405
rect 3172 1076 3258 2319
rect 4003 1076 4089 2319
rect 3172 990 4089 1076
<< mvpsubdiff >>
rect 3198 2345 3281 2379
rect 3315 2345 3349 2379
rect 3383 2345 3417 2379
rect 3451 2345 3485 2379
rect 3519 2345 3553 2379
rect 3587 2345 3621 2379
rect 3655 2345 3689 2379
rect 3723 2345 3757 2379
rect 3791 2345 3825 2379
rect 3859 2345 3893 2379
rect 3927 2345 3961 2379
rect 3995 2345 4063 2379
rect 3198 2311 3232 2345
rect 3198 2243 3232 2277
rect 4029 2274 4063 2345
rect 3198 2175 3232 2209
rect 3198 2107 3232 2141
rect 3198 2039 3232 2073
rect 3198 1971 3232 2005
rect 3198 1903 3232 1937
rect 3198 1835 3232 1869
rect 3198 1767 3232 1801
rect 3198 1699 3232 1733
rect 3198 1631 3232 1665
rect 3198 1563 3232 1597
rect 3198 1495 3232 1529
rect 3198 1427 3232 1461
rect 3198 1359 3232 1393
rect 3198 1291 3232 1325
rect 3198 1223 3232 1257
rect 3198 1155 3232 1189
rect 4029 2206 4063 2240
rect 4029 2138 4063 2172
rect 4029 2070 4063 2104
rect 4029 2002 4063 2036
rect 4029 1934 4063 1968
rect 4029 1866 4063 1900
rect 4029 1798 4063 1832
rect 4029 1730 4063 1764
rect 4029 1662 4063 1696
rect 4029 1594 4063 1628
rect 4029 1526 4063 1560
rect 4029 1458 4063 1492
rect 4029 1390 4063 1424
rect 4029 1322 4063 1356
rect 4029 1254 4063 1288
rect 4029 1186 4063 1220
rect 3198 1050 3232 1121
rect 4029 1118 4063 1152
rect 4029 1050 4063 1084
rect 3198 1016 3266 1050
rect 3300 1016 3334 1050
rect 3368 1016 3402 1050
rect 3436 1016 3470 1050
rect 3504 1016 3538 1050
rect 3572 1016 3606 1050
rect 3640 1016 3674 1050
rect 3708 1016 3742 1050
rect 3776 1016 3810 1050
rect 3844 1016 3878 1050
rect 3912 1016 4063 1050
<< mvnsubdiff >>
rect -347 2882 -311 2943
rect -347 2848 -346 2882
rect -312 2848 -311 2882
rect -347 2814 -311 2848
rect -347 2780 -346 2814
rect -312 2780 -311 2814
rect -347 2746 -311 2780
rect -347 2712 -346 2746
rect -312 2712 -311 2746
rect -347 2678 -311 2712
rect -347 2644 -346 2678
rect -312 2644 -311 2678
rect -347 2610 -311 2644
rect -347 2576 -346 2610
rect -312 2576 -311 2610
rect -347 2542 -311 2576
rect -347 2508 -346 2542
rect -312 2508 -311 2542
rect -347 2474 -311 2508
rect -347 2440 -346 2474
rect -312 2440 -311 2474
rect -347 2406 -311 2440
rect -347 2372 -346 2406
rect -312 2372 -311 2406
rect -347 2338 -311 2372
rect -347 2304 -346 2338
rect -312 2304 -311 2338
rect -347 2270 -311 2304
rect -347 2236 -346 2270
rect -312 2236 -311 2270
rect -347 2202 -311 2236
rect -347 2168 -346 2202
rect -312 2168 -311 2202
rect -347 2134 -311 2168
rect -347 2100 -346 2134
rect -312 2100 -311 2134
rect -347 2066 -311 2100
rect -347 2032 -346 2066
rect -312 2032 -311 2066
rect -347 1998 -311 2032
rect -347 1964 -346 1998
rect -312 1964 -311 1998
rect -347 1930 -311 1964
rect -347 1896 -346 1930
rect -312 1896 -311 1930
rect -347 1862 -311 1896
rect -347 1828 -346 1862
rect -312 1828 -311 1862
rect -347 1794 -311 1828
rect -347 1760 -346 1794
rect -312 1760 -311 1794
rect -347 1726 -311 1760
rect -347 1692 -346 1726
rect -312 1692 -311 1726
rect -347 1658 -311 1692
rect -347 1624 -346 1658
rect -312 1624 -311 1658
rect -347 1590 -311 1624
rect -347 1556 -346 1590
rect -312 1556 -311 1590
rect -347 1522 -311 1556
rect -347 1488 -346 1522
rect -312 1488 -311 1522
rect -347 1454 -311 1488
rect -347 1420 -346 1454
rect -312 1420 -311 1454
rect -347 1386 -311 1420
rect -347 1352 -346 1386
rect -312 1352 -311 1386
rect -347 1318 -311 1352
rect -347 1284 -346 1318
rect -312 1284 -311 1318
rect -347 1250 -311 1284
rect -347 1216 -346 1250
rect -312 1216 -311 1250
rect -347 1182 -311 1216
rect -347 1148 -346 1182
rect -312 1148 -311 1182
rect -347 1114 -311 1148
rect -347 1080 -346 1114
rect -312 1080 -311 1114
rect -347 1046 -311 1080
rect -347 1012 -346 1046
rect -312 1012 -311 1046
rect -347 978 -311 1012
rect -347 944 -346 978
rect -312 944 -311 978
rect -347 910 -311 944
rect -347 876 -346 910
rect -312 876 -311 910
rect -347 842 -311 876
rect -347 808 -346 842
rect -312 808 -311 842
rect -347 774 -311 808
rect -347 740 -346 774
rect -312 740 -311 774
rect -347 706 -311 740
rect -347 672 -346 706
rect -312 672 -311 706
rect -347 638 -311 672
rect -347 604 -346 638
rect -312 604 -311 638
rect -347 570 -311 604
rect -347 536 -346 570
rect -312 536 -311 570
rect -347 502 -311 536
rect -347 468 -346 502
rect -312 468 -311 502
rect -347 434 -311 468
rect -347 400 -346 434
rect -312 400 -311 434
rect -347 366 -311 400
rect -347 332 -346 366
rect -312 332 -311 366
rect -347 298 -311 332
rect -347 264 -346 298
rect -312 264 -311 298
rect -347 230 -311 264
rect -347 196 -346 230
rect -312 196 -311 230
rect -347 162 -311 196
rect -347 128 -346 162
rect -312 128 -311 162
rect -347 94 -311 128
rect -347 60 -346 94
rect -312 62 -311 94
rect 3575 565 3611 599
rect 3575 531 3576 565
rect 3610 531 3611 565
rect 3575 497 3611 531
rect 3575 463 3576 497
rect 3610 463 3611 497
rect 3575 429 3611 463
rect 3575 395 3576 429
rect 3610 395 3611 429
rect 3575 361 3611 395
rect 3575 327 3576 361
rect 3610 327 3611 361
rect 3575 293 3611 327
rect 3575 259 3576 293
rect 3610 259 3611 293
rect 3575 225 3611 259
rect 3575 191 3576 225
rect 3610 191 3611 225
rect 3575 157 3611 191
rect 3575 123 3576 157
rect 3610 123 3611 157
rect 3575 62 3611 123
rect -312 61 3611 62
rect -312 60 -265 61
rect -347 27 -265 60
rect -231 27 -197 61
rect -163 27 -129 61
rect -95 27 -61 61
rect -27 27 7 61
rect 41 27 75 61
rect 109 27 143 61
rect 177 27 211 61
rect 245 27 279 61
rect 313 27 347 61
rect 381 27 415 61
rect 449 27 483 61
rect 517 27 551 61
rect 585 27 619 61
rect 653 27 687 61
rect 721 27 755 61
rect 789 27 823 61
rect 857 27 891 61
rect 925 27 959 61
rect 993 27 1027 61
rect 1061 27 1095 61
rect 1129 27 1163 61
rect 1197 27 1231 61
rect 1265 27 1299 61
rect 1333 27 1367 61
rect 1401 27 1435 61
rect 1469 27 1503 61
rect 1537 27 1571 61
rect 1605 27 1639 61
rect 1673 27 1707 61
rect 1741 27 1775 61
rect 1809 27 1843 61
rect 1877 27 1911 61
rect 1945 27 1979 61
rect 2013 27 2047 61
rect 2081 27 2115 61
rect 2149 27 2183 61
rect 2217 27 2251 61
rect 2285 27 2319 61
rect 2353 27 2387 61
rect 2421 27 2455 61
rect 2489 27 2523 61
rect 2557 27 2591 61
rect 2625 27 2659 61
rect 2693 27 2727 61
rect 2761 27 2795 61
rect 2829 27 2863 61
rect 2897 27 2931 61
rect 2965 27 2999 61
rect 3033 27 3067 61
rect 3101 27 3135 61
rect 3169 27 3203 61
rect 3237 27 3271 61
rect 3305 27 3339 61
rect 3373 27 3407 61
rect 3441 27 3475 61
rect 3509 27 3543 61
rect 3577 27 3611 61
rect -347 26 3611 27
<< mvpsubdiffcont >>
rect 3281 2345 3315 2379
rect 3349 2345 3383 2379
rect 3417 2345 3451 2379
rect 3485 2345 3519 2379
rect 3553 2345 3587 2379
rect 3621 2345 3655 2379
rect 3689 2345 3723 2379
rect 3757 2345 3791 2379
rect 3825 2345 3859 2379
rect 3893 2345 3927 2379
rect 3961 2345 3995 2379
rect 3198 2277 3232 2311
rect 3198 2209 3232 2243
rect 4029 2240 4063 2274
rect 3198 2141 3232 2175
rect 3198 2073 3232 2107
rect 3198 2005 3232 2039
rect 3198 1937 3232 1971
rect 3198 1869 3232 1903
rect 3198 1801 3232 1835
rect 3198 1733 3232 1767
rect 3198 1665 3232 1699
rect 3198 1597 3232 1631
rect 3198 1529 3232 1563
rect 3198 1461 3232 1495
rect 3198 1393 3232 1427
rect 3198 1325 3232 1359
rect 3198 1257 3232 1291
rect 3198 1189 3232 1223
rect 4029 2172 4063 2206
rect 4029 2104 4063 2138
rect 4029 2036 4063 2070
rect 4029 1968 4063 2002
rect 4029 1900 4063 1934
rect 4029 1832 4063 1866
rect 4029 1764 4063 1798
rect 4029 1696 4063 1730
rect 4029 1628 4063 1662
rect 4029 1560 4063 1594
rect 4029 1492 4063 1526
rect 4029 1424 4063 1458
rect 4029 1356 4063 1390
rect 4029 1288 4063 1322
rect 4029 1220 4063 1254
rect 3198 1121 3232 1155
rect 4029 1152 4063 1186
rect 4029 1084 4063 1118
rect 3266 1016 3300 1050
rect 3334 1016 3368 1050
rect 3402 1016 3436 1050
rect 3470 1016 3504 1050
rect 3538 1016 3572 1050
rect 3606 1016 3640 1050
rect 3674 1016 3708 1050
rect 3742 1016 3776 1050
rect 3810 1016 3844 1050
rect 3878 1016 3912 1050
<< mvnsubdiffcont >>
rect -346 2848 -312 2882
rect -346 2780 -312 2814
rect -346 2712 -312 2746
rect -346 2644 -312 2678
rect -346 2576 -312 2610
rect -346 2508 -312 2542
rect -346 2440 -312 2474
rect -346 2372 -312 2406
rect -346 2304 -312 2338
rect -346 2236 -312 2270
rect -346 2168 -312 2202
rect -346 2100 -312 2134
rect -346 2032 -312 2066
rect -346 1964 -312 1998
rect -346 1896 -312 1930
rect -346 1828 -312 1862
rect -346 1760 -312 1794
rect -346 1692 -312 1726
rect -346 1624 -312 1658
rect -346 1556 -312 1590
rect -346 1488 -312 1522
rect -346 1420 -312 1454
rect -346 1352 -312 1386
rect -346 1284 -312 1318
rect -346 1216 -312 1250
rect -346 1148 -312 1182
rect -346 1080 -312 1114
rect -346 1012 -312 1046
rect -346 944 -312 978
rect -346 876 -312 910
rect -346 808 -312 842
rect -346 740 -312 774
rect -346 672 -312 706
rect -346 604 -312 638
rect -346 536 -312 570
rect -346 468 -312 502
rect -346 400 -312 434
rect -346 332 -312 366
rect -346 264 -312 298
rect -346 196 -312 230
rect -346 128 -312 162
rect -346 60 -312 94
rect 3576 531 3610 565
rect 3576 463 3610 497
rect 3576 395 3610 429
rect 3576 327 3610 361
rect 3576 259 3610 293
rect 3576 191 3610 225
rect 3576 123 3610 157
rect -265 27 -231 61
rect -197 27 -163 61
rect -129 27 -95 61
rect -61 27 -27 61
rect 7 27 41 61
rect 75 27 109 61
rect 143 27 177 61
rect 211 27 245 61
rect 279 27 313 61
rect 347 27 381 61
rect 415 27 449 61
rect 483 27 517 61
rect 551 27 585 61
rect 619 27 653 61
rect 687 27 721 61
rect 755 27 789 61
rect 823 27 857 61
rect 891 27 925 61
rect 959 27 993 61
rect 1027 27 1061 61
rect 1095 27 1129 61
rect 1163 27 1197 61
rect 1231 27 1265 61
rect 1299 27 1333 61
rect 1367 27 1401 61
rect 1435 27 1469 61
rect 1503 27 1537 61
rect 1571 27 1605 61
rect 1639 27 1673 61
rect 1707 27 1741 61
rect 1775 27 1809 61
rect 1843 27 1877 61
rect 1911 27 1945 61
rect 1979 27 2013 61
rect 2047 27 2081 61
rect 2115 27 2149 61
rect 2183 27 2217 61
rect 2251 27 2285 61
rect 2319 27 2353 61
rect 2387 27 2421 61
rect 2455 27 2489 61
rect 2523 27 2557 61
rect 2591 27 2625 61
rect 2659 27 2693 61
rect 2727 27 2761 61
rect 2795 27 2829 61
rect 2863 27 2897 61
rect 2931 27 2965 61
rect 2999 27 3033 61
rect 3067 27 3101 61
rect 3135 27 3169 61
rect 3203 27 3237 61
rect 3271 27 3305 61
rect 3339 27 3373 61
rect 3407 27 3441 61
rect 3475 27 3509 61
rect 3543 27 3577 61
<< poly >>
rect 3930 2199 3996 2215
rect 3930 2165 3946 2199
rect 3980 2165 3996 2199
rect 3930 2130 3996 2165
rect 3930 2096 3946 2130
rect 3980 2096 3996 2130
rect 3930 2061 3996 2096
rect 3930 2027 3946 2061
rect 3980 2027 3996 2061
rect 3930 1992 3996 2027
rect 3930 1958 3946 1992
rect 3980 1958 3996 1992
rect 3930 1923 3996 1958
rect 3930 1889 3946 1923
rect 3980 1889 3996 1923
rect 3930 1854 3996 1889
rect 3930 1820 3946 1854
rect 3980 1820 3996 1854
rect 3930 1785 3996 1820
rect 3930 1751 3946 1785
rect 3980 1751 3996 1785
rect 3930 1716 3996 1751
rect 3930 1682 3946 1716
rect 3980 1682 3996 1716
rect 3930 1647 3996 1682
rect 3930 1613 3946 1647
rect 3980 1613 3996 1647
rect 3930 1578 3996 1613
rect 3930 1544 3946 1578
rect 3980 1544 3996 1578
rect 3930 1509 3996 1544
rect 3930 1475 3946 1509
rect 3980 1475 3996 1509
rect 3930 1439 3996 1475
rect 3930 1405 3946 1439
rect 3980 1405 3996 1439
rect 3930 1369 3996 1405
rect 3930 1335 3946 1369
rect 3980 1335 3996 1369
rect 3930 1299 3996 1335
rect 3930 1265 3946 1299
rect 3980 1265 3996 1299
rect 3930 1229 3996 1265
rect 3930 1195 3946 1229
rect 3980 1195 3996 1229
rect 3930 1179 3996 1195
<< polycont >>
rect 3946 2165 3980 2199
rect 3946 2096 3980 2130
rect 3946 2027 3980 2061
rect 3946 1958 3980 1992
rect 3946 1889 3980 1923
rect 3946 1820 3980 1854
rect 3946 1751 3980 1785
rect 3946 1682 3980 1716
rect 3946 1613 3980 1647
rect 3946 1544 3980 1578
rect 3946 1475 3980 1509
rect 3946 1405 3980 1439
rect 3946 1335 3980 1369
rect 3946 1265 3980 1299
rect 3946 1195 3980 1229
<< locali >>
rect 375 17510 2047 17516
rect 375 17476 407 17510
rect 441 17476 482 17510
rect 516 17476 557 17510
rect 591 17476 632 17510
rect 666 17476 707 17510
rect 741 17476 782 17510
rect 816 17476 857 17510
rect 891 17476 932 17510
rect 966 17476 1007 17510
rect 1041 17476 1082 17510
rect 1116 17476 1157 17510
rect 1191 17476 1232 17510
rect 1266 17476 1307 17510
rect 1341 17476 1382 17510
rect 1416 17476 1457 17510
rect 1491 17476 1532 17510
rect 1566 17476 1607 17510
rect 1641 17476 1682 17510
rect 1716 17476 1757 17510
rect 1791 17476 1832 17510
rect 1866 17476 1907 17510
rect 1941 17476 1981 17510
rect 2015 17476 2047 17510
rect 375 17470 2047 17476
rect 2268 17510 3061 17516
rect 2268 17476 2300 17510
rect 2334 17476 2378 17510
rect 2412 17476 2456 17510
rect 2490 17476 2533 17510
rect 2567 17476 2610 17510
rect 2644 17476 2687 17510
rect 2721 17476 2764 17510
rect 2798 17476 2841 17510
rect 2875 17476 2918 17510
rect 2952 17476 2995 17510
rect 3029 17476 3061 17510
rect 2268 17470 3061 17476
rect 381 17331 415 17369
rect 381 17259 415 17297
rect 381 17187 415 17225
rect 381 17115 415 17153
rect 381 17043 415 17081
rect 381 16971 415 17009
rect 381 16899 415 16937
rect 381 16827 415 16865
rect 381 16755 415 16793
rect 381 16682 415 16721
rect 381 16609 415 16648
rect 381 16536 415 16575
rect 381 16463 415 16502
rect 381 16390 415 16429
rect 381 16317 415 16356
rect 381 16244 415 16283
rect 381 16171 415 16210
rect 381 16098 415 16137
rect 381 16025 415 16064
rect 381 15952 415 15991
rect 381 15879 415 15918
rect 381 15806 415 15845
rect 381 15733 415 15772
rect 381 15660 415 15699
rect 381 15587 415 15626
rect 381 15514 415 15553
rect 381 15441 415 15480
rect 381 15368 415 15407
rect 381 15295 415 15334
rect 381 15222 415 15261
rect 381 15149 415 15188
rect 381 15076 415 15115
rect 381 15003 415 15042
rect 381 14930 415 14969
rect 381 14857 415 14896
rect 381 14784 415 14823
rect 381 14711 415 14750
rect 381 14638 415 14677
rect 381 14565 415 14604
rect 381 14492 415 14531
rect 381 14419 415 14458
rect 381 14346 415 14385
rect 381 14273 415 14312
rect 381 14200 415 14239
rect 381 14127 415 14166
rect 381 14054 415 14093
rect 381 13981 415 14020
rect 381 13908 415 13947
rect 381 13835 415 13874
rect 381 13762 415 13801
rect 381 13689 415 13728
rect 381 13616 415 13655
rect 381 13543 415 13582
rect 381 13470 415 13509
rect 381 13397 415 13436
rect 381 13324 415 13363
rect 381 13251 415 13290
rect 381 13178 415 13217
rect 1701 17321 1735 17360
rect 1701 17248 1735 17287
rect 1701 17175 1735 17214
rect 1701 17102 1735 17141
rect 1701 17029 1735 17068
rect 1701 16956 1735 16995
rect 1701 16883 1735 16922
rect 1701 16810 1735 16849
rect 1701 16737 1735 16776
rect 1701 16664 1735 16703
rect 1701 16591 1735 16630
rect 1701 16518 1735 16557
rect 1701 16445 1735 16484
rect 1701 16372 1735 16411
rect 1701 16299 1735 16338
rect 1701 16226 1735 16265
rect 1701 16153 1735 16192
rect 1701 16080 1735 16119
rect 1701 16007 1735 16046
rect 1701 15934 1735 15973
rect 1701 15861 1735 15900
rect 1701 15788 1735 15827
rect 1701 15715 1735 15754
rect 1701 15642 1735 15681
rect 1701 15569 1735 15608
rect 1701 15496 1735 15535
rect 1701 15423 1735 15462
rect 1701 15350 1735 15389
rect 1701 15277 1735 15316
rect 1701 15204 1735 15243
rect 1701 15131 1735 15170
rect 1701 15058 1735 15097
rect 1701 14985 1735 15024
rect 1701 14912 1735 14951
rect 1701 14839 1735 14878
rect 1701 14766 1735 14805
rect 1701 14693 1735 14732
rect 1701 14620 1735 14659
rect 1701 14547 1735 14586
rect 1701 14474 1735 14513
rect 1701 14401 1735 14440
rect 1701 14328 1735 14367
rect 1701 14255 1735 14294
rect 1701 14182 1735 14221
rect 1701 14109 1735 14148
rect 1701 14036 1735 14075
rect 1701 13963 1735 14002
rect 1701 13890 1735 13929
rect 1701 13817 1735 13856
rect 1701 13744 1735 13783
rect 1701 13671 1735 13710
rect 1701 13598 1735 13637
rect 1701 13524 1735 13564
rect 1701 13450 1735 13490
rect 1701 13376 1735 13416
rect 1701 13302 1735 13342
rect 1701 13228 1735 13268
rect 3021 17356 3055 17395
rect 3021 17283 3055 17322
rect 3021 17210 3055 17249
rect 3021 17137 3055 17176
rect 3021 17064 3055 17103
rect 3021 16991 3055 17030
rect 3021 16918 3055 16957
rect 3021 16845 3055 16884
rect 3021 16772 3055 16811
rect 3021 16699 3055 16738
rect 3021 16626 3055 16665
rect 3021 16553 3055 16592
rect 3021 16480 3055 16519
rect 3021 16407 3055 16446
rect 3021 16334 3055 16373
rect 3021 16261 3055 16300
rect 3021 16188 3055 16227
rect 3021 16115 3055 16154
rect 3021 16042 3055 16081
rect 3021 15969 3055 16008
rect 3021 15896 3055 15935
rect 3021 15823 3055 15862
rect 3021 15750 3055 15789
rect 3021 15677 3055 15716
rect 3021 15604 3055 15643
rect 3021 15531 3055 15570
rect 3021 15458 3055 15497
rect 3021 15385 3055 15424
rect 3021 15312 3055 15351
rect 3021 15239 3055 15278
rect 3021 15166 3055 15205
rect 3021 15093 3055 15132
rect 3021 15020 3055 15059
rect 3021 14947 3055 14986
rect 3021 14874 3055 14913
rect 3021 14801 3055 14840
rect 3021 14728 3055 14767
rect 3021 14655 3055 14694
rect 3021 14582 3055 14621
rect 3021 14509 3055 14548
rect 3021 14436 3055 14475
rect 3021 14363 3055 14402
rect 3021 14290 3055 14329
rect 3021 14217 3055 14256
rect 3021 14144 3055 14183
rect 3021 14071 3055 14110
rect 3021 13998 3055 14037
rect 3021 13925 3055 13964
rect 3021 13852 3055 13891
rect 3021 13779 3055 13818
rect 3021 13706 3055 13745
rect 3021 13633 3055 13672
rect 3021 13560 3055 13599
rect 3021 13487 3055 13526
rect 3021 13414 3055 13453
rect 3021 13341 3055 13380
rect 3021 13268 3055 13307
rect 3021 13195 3055 13234
rect 381 13105 415 13144
rect 381 13032 415 13071
rect 3021 13122 3055 13161
rect 3021 13048 3055 13088
rect 381 12959 415 12998
rect 381 12886 415 12925
rect 381 12813 415 12852
rect 381 12740 415 12779
rect 381 12667 415 12706
rect 381 12594 415 12633
rect 381 12521 415 12560
rect 381 12448 415 12487
rect 381 11512 415 11550
rect 381 11440 415 11478
rect 381 11368 415 11406
rect 381 11296 415 11334
rect 381 11224 415 11262
rect 381 11152 415 11190
rect 381 11080 415 11118
rect 381 11008 415 11046
rect 381 10936 415 10974
rect 381 10864 415 10902
rect 381 10792 415 10830
rect 381 10720 415 10758
rect 381 10648 415 10686
rect 381 10576 415 10614
rect 381 10504 415 10542
rect 381 10432 415 10470
rect 381 10360 415 10398
rect 381 10288 415 10326
rect 381 10216 415 10254
rect 381 10144 415 10182
rect 381 10072 415 10110
rect 381 10000 415 10038
rect 381 9928 415 9966
rect 381 9856 415 9894
rect 381 9784 415 9822
rect 381 9712 415 9750
rect 381 9640 415 9678
rect 381 9568 415 9606
rect 381 9496 415 9534
rect 381 9424 415 9462
rect 381 9352 415 9390
rect 381 9280 415 9318
rect 381 9208 415 9246
rect 381 9136 415 9174
rect 381 9064 415 9102
rect 381 8992 415 9030
rect 381 8920 415 8958
rect 381 8848 415 8886
rect 381 8776 415 8814
rect 381 8704 415 8742
rect 381 8632 415 8670
rect 381 8560 415 8598
rect 381 8488 415 8526
rect 381 8416 415 8454
rect 381 8344 415 8382
rect 381 8272 415 8310
rect 381 8200 415 8238
rect 381 8128 415 8166
rect 381 8056 415 8094
rect 381 7984 415 8022
rect 381 7912 415 7950
rect 381 7840 415 7878
rect 381 7768 415 7806
rect 381 7696 415 7734
rect 381 7624 415 7662
rect 381 7552 415 7590
rect 381 7480 415 7518
rect 381 7408 415 7446
rect 381 7336 415 7374
rect 381 7264 415 7302
rect 381 7192 415 7230
rect 381 7120 415 7158
rect 381 7048 415 7086
rect 381 6976 415 7014
rect 381 6904 415 6942
rect 381 6832 415 6870
rect 381 6760 415 6798
rect 381 6688 415 6726
rect 381 6616 415 6654
rect 381 6544 415 6582
rect 381 6472 415 6510
rect 381 6400 415 6438
rect 381 6328 415 6366
rect 381 6256 415 6294
rect 381 6184 415 6222
rect 381 6112 415 6150
rect 381 6040 415 6078
rect 381 5968 415 6006
rect 381 5896 415 5934
rect 381 5824 415 5862
rect 381 5752 415 5790
rect 381 5680 415 5718
rect 381 5608 415 5646
rect 381 5536 415 5574
rect 381 5464 415 5502
rect 381 5392 415 5430
rect 381 5320 415 5358
rect 381 5248 415 5286
rect 381 5176 415 5214
rect 381 5104 415 5142
rect 381 5032 415 5070
rect 381 4960 415 4998
rect 381 4888 415 4926
rect 381 4816 415 4854
rect 381 4744 415 4782
rect 381 4672 415 4710
rect 381 4600 415 4638
rect 381 4528 415 4566
rect 381 4456 415 4494
rect 381 4384 415 4422
rect 381 4312 415 4350
rect 381 4240 415 4278
rect 381 4168 415 4206
rect 3021 10278 3055 10316
rect 3021 10206 3055 10244
rect 3021 10134 3055 10172
rect 3021 10062 3055 10100
rect 3021 9990 3055 10028
rect 3021 9918 3055 9956
rect 3021 9846 3055 9884
rect 3021 9774 3055 9812
rect 3021 9702 3055 9740
rect 3021 9630 3055 9668
rect 3021 9558 3055 9596
rect 3021 9486 3055 9524
rect 3021 9414 3055 9452
rect 3021 9342 3055 9380
rect 3021 9270 3055 9308
rect 3021 9198 3055 9236
rect 3021 9126 3055 9164
rect 3021 9054 3055 9092
rect 3021 8982 3055 9020
rect 3021 8910 3055 8948
rect 3021 8838 3055 8876
rect 3021 8766 3055 8804
rect 3021 8694 3055 8732
rect 3021 8622 3055 8660
rect 3021 8550 3055 8588
rect 3021 8478 3055 8516
rect 3021 8406 3055 8444
rect 3021 8334 3055 8372
rect 3021 8262 3055 8300
rect 3021 8190 3055 8228
rect 3021 8118 3055 8156
rect 3021 8046 3055 8084
rect 3021 7974 3055 8012
rect 3021 7902 3055 7940
rect 3021 7830 3055 7868
rect 3021 7758 3055 7796
rect 3021 7686 3055 7724
rect 3021 7614 3055 7652
rect 3021 7542 3055 7580
rect 3021 7470 3055 7508
rect 3021 7398 3055 7436
rect 3021 7326 3055 7364
rect 3021 7254 3055 7292
rect 3021 7182 3055 7220
rect 3021 7110 3055 7148
rect 3021 7038 3055 7076
rect 3021 6966 3055 7004
rect 3021 6894 3055 6932
rect 3021 6822 3055 6860
rect 3021 6750 3055 6788
rect 3021 6678 3055 6716
rect 3021 6606 3055 6644
rect 3021 6534 3055 6572
rect 3021 6462 3055 6500
rect 3021 6390 3055 6428
rect 3021 6318 3055 6356
rect 3021 6246 3055 6284
rect 3021 6174 3055 6212
rect 3021 6102 3055 6140
rect 3021 6030 3055 6068
rect 3021 5958 3055 5996
rect 3021 5886 3055 5924
rect 3021 5814 3055 5852
rect 3021 5742 3055 5780
rect 3021 5670 3055 5708
rect 3021 5598 3055 5636
rect 3021 5526 3055 5564
rect 3021 5454 3055 5492
rect 3021 5382 3055 5420
rect 3021 5309 3055 5348
rect 3021 5236 3055 5275
rect 3021 5163 3055 5202
rect 3021 5090 3055 5129
rect 3021 5017 3055 5056
rect 3021 4944 3055 4983
rect 3021 4871 3055 4910
rect 3021 4798 3055 4837
rect 3021 4725 3055 4764
rect 3021 4652 3055 4691
rect 3021 4579 3055 4618
rect 3021 4506 3055 4545
rect 3021 4433 3055 4472
rect 3021 4360 3055 4399
rect 3021 4287 3055 4326
rect 3021 4214 3055 4253
rect 381 4095 415 4134
rect 381 4022 415 4061
rect 381 3949 415 3988
rect 381 3876 415 3915
rect 381 3803 415 3842
rect 381 3730 415 3769
rect 381 3657 415 3696
rect 381 3584 415 3623
rect 381 3511 415 3550
rect 381 3438 415 3477
rect 381 3365 415 3404
rect 381 3292 415 3331
rect 381 3219 415 3258
rect 381 3146 415 3185
rect 381 3073 415 3112
rect 381 3000 415 3039
rect -347 2882 -311 2943
rect -347 2848 -346 2882
rect -312 2848 -311 2882
rect -347 2814 -311 2848
rect -347 2780 -346 2814
rect -312 2780 -311 2814
rect -347 2746 -311 2780
rect -347 2712 -346 2746
rect -312 2712 -311 2746
rect -347 2678 -311 2712
rect -347 2644 -346 2678
rect -312 2644 -311 2678
rect -347 2610 -311 2644
rect -347 2576 -346 2610
rect -312 2576 -311 2610
rect -347 2542 -311 2576
rect -347 2508 -346 2542
rect -312 2508 -311 2542
rect -347 2474 -311 2508
rect -347 2440 -346 2474
rect -312 2440 -311 2474
rect -347 2406 -311 2440
rect -347 2372 -346 2406
rect -312 2372 -311 2406
rect -347 2338 -311 2372
rect -347 2304 -346 2338
rect -312 2304 -311 2338
rect -347 2270 -311 2304
rect -347 2236 -346 2270
rect -312 2236 -311 2270
rect -347 2202 -311 2236
rect -347 2168 -346 2202
rect -312 2168 -311 2202
rect -347 2134 -311 2168
rect -347 2100 -346 2134
rect -312 2100 -311 2134
rect -347 2066 -311 2100
rect -347 2032 -346 2066
rect -312 2032 -311 2066
rect -347 1998 -311 2032
rect -347 1964 -346 1998
rect -312 1964 -311 1998
rect -347 1930 -311 1964
rect -347 1896 -346 1930
rect -312 1896 -311 1930
rect -347 1862 -311 1896
rect -347 1828 -346 1862
rect -312 1828 -311 1862
rect -347 1794 -311 1828
rect -347 1760 -346 1794
rect -312 1760 -311 1794
rect -347 1726 -311 1760
rect -347 1692 -346 1726
rect -312 1692 -311 1726
rect -347 1658 -311 1692
rect -347 1624 -346 1658
rect -312 1624 -311 1658
rect -347 1590 -311 1624
rect -347 1556 -346 1590
rect -312 1556 -311 1590
rect -347 1522 -311 1556
rect -347 1488 -346 1522
rect -312 1488 -311 1522
rect -347 1454 -311 1488
rect -347 1420 -346 1454
rect -312 1420 -311 1454
rect -347 1386 -311 1420
rect -347 1352 -346 1386
rect -312 1352 -311 1386
rect -347 1318 -311 1352
rect -347 1284 -346 1318
rect -312 1284 -311 1318
rect -347 1250 -311 1284
rect -347 1216 -346 1250
rect -312 1216 -311 1250
rect -347 1182 -311 1216
rect -347 1148 -346 1182
rect -312 1148 -311 1182
rect -347 1114 -311 1148
rect -347 1080 -346 1114
rect -312 1080 -311 1114
rect -347 1046 -311 1080
rect -347 1012 -346 1046
rect -312 1012 -311 1046
rect -347 978 -311 1012
rect -347 944 -346 978
rect -312 944 -311 978
rect -347 910 -311 944
rect 381 2927 415 2966
rect 381 2854 415 2893
rect 381 2781 415 2820
rect 381 2708 415 2747
rect 381 2635 415 2674
rect 381 2562 415 2601
rect 381 2489 415 2528
rect 381 2416 415 2455
rect 381 2343 415 2382
rect 381 2270 415 2309
rect 381 2197 415 2236
rect 381 2124 415 2163
rect 381 2051 415 2090
rect 381 1978 415 2017
rect 381 1905 415 1944
rect 381 1832 415 1871
rect 381 1759 415 1798
rect 381 1686 415 1725
rect 381 1613 415 1652
rect 381 1540 415 1579
rect 381 1467 415 1506
rect 381 1394 415 1433
rect 381 1321 415 1360
rect 381 1248 415 1287
rect 381 1175 415 1214
rect 381 1102 415 1141
rect 381 1029 415 1068
rect 381 956 415 995
rect 1695 3642 1741 3674
rect 1695 3608 1701 3642
rect 1735 3608 1741 3642
rect 1695 3570 1741 3608
rect 1695 3536 1701 3570
rect 1735 3536 1741 3570
rect 1695 3498 1741 3536
rect 1695 3464 1701 3498
rect 1735 3464 1741 3498
rect 1695 3426 1741 3464
rect 1695 3392 1701 3426
rect 1735 3392 1741 3426
rect 1695 3354 1741 3392
rect 1695 3320 1701 3354
rect 1735 3320 1741 3354
rect 1695 3282 1741 3320
rect 1695 3248 1701 3282
rect 1735 3248 1741 3282
rect 1695 3210 1741 3248
rect 1695 3176 1701 3210
rect 1735 3176 1741 3210
rect 1695 3138 1741 3176
rect 1695 3104 1701 3138
rect 1735 3104 1741 3138
rect 1695 3066 1741 3104
rect 1695 3032 1701 3066
rect 1735 3032 1741 3066
rect 1695 2994 1741 3032
rect 1695 2960 1701 2994
rect 1735 2960 1741 2994
rect 1695 2922 1741 2960
rect 1695 2888 1701 2922
rect 1735 2888 1741 2922
rect 1695 2850 1741 2888
rect 1695 2816 1701 2850
rect 1735 2816 1741 2850
rect 1695 2778 1741 2816
rect 1695 2744 1701 2778
rect 1735 2744 1741 2778
rect 1695 2706 1741 2744
rect 1695 2672 1701 2706
rect 1735 2672 1741 2706
rect 1695 2634 1741 2672
rect 1695 2600 1701 2634
rect 1735 2600 1741 2634
rect 1695 2562 1741 2600
rect 1695 2528 1701 2562
rect 1735 2528 1741 2562
rect 1695 2490 1741 2528
rect 1695 2456 1701 2490
rect 1735 2456 1741 2490
rect 1695 2418 1741 2456
rect 1695 2384 1701 2418
rect 1735 2384 1741 2418
rect 1695 2346 1741 2384
rect 1695 2312 1701 2346
rect 1735 2312 1741 2346
rect 1695 2274 1741 2312
rect 1695 2240 1701 2274
rect 1735 2240 1741 2274
rect 1695 2202 1741 2240
rect 1695 2168 1701 2202
rect 1735 2168 1741 2202
rect 1695 2130 1741 2168
rect 1695 2096 1701 2130
rect 1735 2096 1741 2130
rect 1695 2058 1741 2096
rect 1695 2024 1701 2058
rect 1735 2024 1741 2058
rect 3189 2379 3414 2388
rect 3189 2345 3201 2379
rect 3235 2345 3273 2379
rect 3315 2345 3345 2379
rect 3383 2345 3417 2379
rect 3451 2345 3485 2379
rect 3519 2345 3553 2379
rect 3587 2345 3621 2379
rect 3655 2345 3689 2379
rect 3723 2345 3757 2379
rect 3791 2345 3825 2379
rect 3859 2345 3893 2379
rect 3927 2345 3961 2379
rect 3995 2345 4063 2379
rect 3189 2336 3414 2345
rect 3189 2311 3241 2336
rect 3189 2271 3198 2311
rect 3232 2271 3241 2311
rect 3189 2243 3241 2271
rect 4029 2274 4063 2345
rect 3189 2199 3198 2243
rect 3232 2199 3241 2243
rect 3384 2226 3422 2260
rect 3456 2226 3494 2260
rect 3528 2226 3566 2260
rect 3600 2226 3638 2260
rect 3189 2175 3241 2199
rect 3189 2127 3198 2175
rect 3232 2127 3241 2175
rect 3189 2107 3241 2127
rect 3189 2055 3198 2107
rect 3232 2055 3241 2107
rect 3946 2159 3980 2165
rect 3661 2070 3699 2104
rect 3733 2070 3771 2104
rect 3805 2070 3843 2104
rect 3189 2043 3241 2055
rect 3946 2061 3980 2096
rect 1695 1986 1741 2024
rect 1695 1952 1701 1986
rect 1735 1952 1741 1986
rect 1695 1914 1741 1952
rect 1695 1880 1701 1914
rect 1735 1880 1741 1914
rect 1695 1842 1741 1880
rect 1695 1808 1701 1842
rect 1735 1808 1741 1842
rect 1695 1770 1741 1808
rect 1695 1736 1701 1770
rect 1735 1736 1741 1770
rect 1695 1698 1741 1736
rect 3198 2039 3232 2043
rect 3198 1971 3232 2005
rect 3946 1992 3980 2027
rect 3198 1903 3232 1937
rect 3384 1914 3422 1948
rect 3456 1914 3494 1948
rect 3528 1914 3566 1948
rect 3600 1914 3638 1948
rect 3946 1923 3980 1958
rect 3198 1835 3232 1869
rect 3198 1767 3232 1801
rect 3946 1854 3980 1889
rect 3618 1758 3656 1792
rect 3690 1758 3728 1792
rect 3762 1758 3800 1792
rect 3834 1758 3872 1792
rect 3946 1785 3980 1820
rect 3198 1730 3232 1733
rect 1695 1664 1701 1698
rect 1735 1664 1741 1698
rect 1695 1626 1741 1664
rect 1695 1592 1701 1626
rect 1735 1592 1741 1626
rect 1695 1554 1741 1592
rect 1695 1520 1701 1554
rect 1735 1520 1741 1554
rect 1695 1482 1741 1520
rect 1695 1448 1701 1482
rect 1735 1448 1741 1482
rect 1695 1410 1741 1448
rect 1695 1376 1701 1410
rect 1735 1376 1741 1410
rect 1695 1338 1741 1376
rect 1695 1304 1701 1338
rect 1735 1304 1741 1338
rect 1695 1266 1741 1304
rect 1695 1232 1701 1266
rect 1735 1232 1741 1266
rect 1695 1194 1741 1232
rect 1695 1160 1701 1194
rect 1735 1160 1741 1194
rect 1695 1122 1741 1160
rect 1695 1088 1701 1122
rect 1735 1088 1741 1122
rect 1695 1050 1741 1088
rect 1695 1016 1701 1050
rect 1735 1016 1741 1050
rect 1695 978 1741 1016
rect 3189 1718 3241 1730
rect 3189 1665 3198 1718
rect 3232 1665 3241 1718
rect 3189 1646 3241 1665
rect 3189 1597 3198 1646
rect 3232 1597 3241 1646
rect 3946 1716 3980 1751
rect 3946 1647 3980 1682
rect 3384 1602 3422 1636
rect 3456 1602 3494 1636
rect 3528 1602 3566 1636
rect 3600 1602 3638 1636
rect 3189 1574 3241 1597
rect 3189 1529 3198 1574
rect 3232 1529 3241 1574
rect 3189 1502 3241 1529
rect 3189 1461 3198 1502
rect 3232 1461 3241 1502
rect 3946 1578 3980 1613
rect 3946 1509 3980 1544
rect 3189 1430 3241 1461
rect 3618 1446 3656 1480
rect 3690 1446 3728 1480
rect 3762 1446 3800 1480
rect 3834 1446 3872 1480
rect 3189 1393 3198 1430
rect 3232 1393 3241 1430
rect 3189 1359 3241 1393
rect 3189 1324 3198 1359
rect 3232 1324 3241 1359
rect 3946 1439 3980 1475
rect 3946 1369 3980 1405
rect 3189 1291 3241 1324
rect 3189 1252 3198 1291
rect 3232 1252 3241 1291
rect 3384 1290 3422 1324
rect 3456 1290 3494 1324
rect 3528 1290 3566 1324
rect 3600 1290 3638 1324
rect 3946 1299 3980 1335
rect 3189 1223 3241 1252
rect 3189 1180 3198 1223
rect 3232 1180 3241 1223
rect 3946 1229 3980 1265
rect 3189 1155 3241 1180
rect 3189 1108 3198 1155
rect 3232 1108 3241 1155
rect 3618 1154 3656 1188
rect 3690 1154 3728 1188
rect 3762 1154 3800 1188
rect 3834 1154 3872 1188
rect 3946 1179 3980 1195
rect 4029 2206 4063 2240
rect 4029 2138 4063 2172
rect 4029 2070 4063 2104
rect 4029 2002 4063 2036
rect 4029 1934 4063 1968
rect 4029 1866 4063 1900
rect 4029 1798 4063 1832
rect 4029 1730 4063 1764
rect 4029 1662 4063 1696
rect 4029 1594 4063 1628
rect 4029 1526 4063 1560
rect 4029 1458 4063 1492
rect 4029 1390 4063 1424
rect 4029 1322 4063 1356
rect 4029 1254 4063 1288
rect 4029 1186 4063 1220
rect 3189 1059 3241 1108
rect 4029 1118 4063 1152
rect 3189 1050 3414 1059
rect 4029 1050 4063 1084
rect 3189 1016 3201 1050
rect 3235 1016 3266 1050
rect 3307 1016 3334 1050
rect 3379 1016 3402 1050
rect 3436 1016 3470 1050
rect 3504 1016 3538 1050
rect 3572 1016 3606 1050
rect 3640 1016 3674 1050
rect 3708 1016 3742 1050
rect 3776 1016 3810 1050
rect 3844 1016 3878 1050
rect 3912 1016 4063 1050
rect 3189 1007 3414 1016
rect 1695 944 1701 978
rect 1735 944 1741 978
rect -347 876 -346 910
rect -312 876 -311 910
rect -347 842 -311 876
rect -347 808 -346 842
rect -312 808 -311 842
rect -347 774 -311 808
rect -347 740 -346 774
rect -312 740 -311 774
rect -347 706 -311 740
rect -347 672 -346 706
rect -312 672 -311 706
rect -347 638 -311 672
rect -347 604 -346 638
rect -312 604 -311 638
rect 1695 906 1741 944
rect 1695 872 1701 906
rect 1735 872 1741 906
rect 1695 834 1741 872
rect 1695 800 1701 834
rect 1735 800 1741 834
rect 1695 762 1741 800
rect 1695 728 1701 762
rect 1735 728 1741 762
rect 1695 690 1741 728
rect 1695 656 1701 690
rect 1735 656 1741 690
rect -347 570 -311 604
rect -347 536 -346 570
rect -312 536 -311 570
rect -347 502 -311 536
rect -347 468 -346 502
rect -312 468 -311 502
rect -347 434 -311 468
rect -347 400 -346 434
rect -312 400 -311 434
rect -347 366 -311 400
rect -347 332 -346 366
rect -312 332 -311 366
rect -347 298 -311 332
rect 381 530 415 584
rect 381 442 415 496
rect 381 353 415 408
rect 1695 617 1741 656
rect 1695 583 1701 617
rect 1735 583 1741 617
rect 1695 544 1741 583
rect 1695 510 1701 544
rect 1735 510 1741 544
rect 1695 471 1741 510
rect 1695 437 1701 471
rect 1735 437 1741 471
rect 1695 398 1741 437
rect 1695 364 1701 398
rect 1735 364 1741 398
rect 1695 332 1741 364
rect 3575 587 3611 599
rect 3575 531 3576 587
rect 3610 531 3611 587
rect 3575 511 3611 531
rect 3575 463 3576 511
rect 3610 463 3611 511
rect 3575 436 3611 463
rect 3575 395 3576 436
rect 3610 395 3611 436
rect 3575 361 3611 395
rect 3575 327 3576 361
rect 3610 327 3611 361
rect -347 264 -346 298
rect -312 264 -311 298
rect -347 230 -311 264
rect 3575 293 3611 327
rect 3575 252 3576 293
rect 3610 252 3611 293
rect -347 196 -346 230
rect -312 196 -311 230
rect 427 216 466 250
rect 500 216 539 250
rect 573 216 612 250
rect 646 216 685 250
rect 719 216 758 250
rect 792 216 831 250
rect 865 216 904 250
rect 938 216 977 250
rect 1011 216 1050 250
rect 1084 216 1123 250
rect 1157 216 1196 250
rect 1230 216 1269 250
rect 1303 216 1342 250
rect 1376 216 1415 250
rect 1449 216 1488 250
rect 1522 216 1561 250
rect 1595 216 1634 250
rect 1668 216 1707 250
rect 1741 216 1780 250
rect 1814 216 1853 250
rect 1887 216 1926 250
rect 1960 216 1999 250
rect 2033 216 2072 250
rect 2106 216 2145 250
rect 2179 216 2217 250
rect 2251 216 2289 250
rect 2323 216 2361 250
rect 2395 216 2433 250
rect 2467 216 2505 250
rect 2539 216 2577 250
rect 2611 216 2649 250
rect 2683 216 2721 250
rect 2755 216 2793 250
rect 2827 216 2865 250
rect 2899 216 2937 250
rect 2971 216 3009 250
rect 3575 225 3611 252
rect -347 162 -311 196
rect -347 128 -346 162
rect -312 128 -311 162
rect -347 94 -311 128
rect -347 60 -346 94
rect -312 62 -311 94
rect 3575 177 3576 225
rect 3610 177 3611 225
rect 3575 157 3611 177
rect 3575 102 3576 157
rect 3610 102 3611 157
rect 3575 62 3611 102
rect -312 61 3611 62
rect -312 60 -265 61
rect -347 27 -265 60
rect -231 27 -197 61
rect -163 27 -129 61
rect -95 27 -61 61
rect -27 27 7 61
rect 41 27 75 61
rect 109 27 143 61
rect 177 27 211 61
rect 245 27 279 61
rect 313 27 347 61
rect 381 27 415 61
rect 449 27 483 61
rect 517 27 551 61
rect 585 27 619 61
rect 653 27 687 61
rect 721 27 755 61
rect 789 27 823 61
rect 857 27 891 61
rect 925 27 959 61
rect 993 27 1027 61
rect 1061 27 1095 61
rect 1129 27 1163 61
rect 1197 27 1231 61
rect 1265 27 1299 61
rect 1333 27 1367 61
rect 1401 27 1435 61
rect 1469 27 1503 61
rect 1537 27 1571 61
rect 1605 27 1639 61
rect 1673 27 1707 61
rect 1741 27 1775 61
rect 1809 27 1843 61
rect 1877 27 1911 61
rect 1945 27 1979 61
rect 2013 27 2047 61
rect 2081 27 2115 61
rect 2149 27 2183 61
rect 2217 27 2251 61
rect 2285 27 2319 61
rect 2353 27 2387 61
rect 2421 27 2455 61
rect 2489 27 2523 61
rect 2557 27 2591 61
rect 2625 27 2659 61
rect 2693 27 2727 61
rect 2761 27 2795 61
rect 2829 27 2863 61
rect 2897 27 2931 61
rect 2965 27 2999 61
rect 3033 27 3067 61
rect 3101 27 3135 61
rect 3169 27 3203 61
rect 3237 27 3271 61
rect 3305 27 3339 61
rect 3373 27 3407 61
rect 3441 27 3475 61
rect 3509 27 3543 61
rect 3610 27 3611 61
rect -347 26 3611 27
<< viali >>
rect 407 17476 441 17510
rect 482 17476 516 17510
rect 557 17476 591 17510
rect 632 17476 666 17510
rect 707 17476 741 17510
rect 782 17476 816 17510
rect 857 17476 891 17510
rect 932 17476 966 17510
rect 1007 17476 1041 17510
rect 1082 17476 1116 17510
rect 1157 17476 1191 17510
rect 1232 17476 1266 17510
rect 1307 17476 1341 17510
rect 1382 17476 1416 17510
rect 1457 17476 1491 17510
rect 1532 17476 1566 17510
rect 1607 17476 1641 17510
rect 1682 17476 1716 17510
rect 1757 17476 1791 17510
rect 1832 17476 1866 17510
rect 1907 17476 1941 17510
rect 1981 17476 2015 17510
rect 2300 17476 2334 17510
rect 2378 17476 2412 17510
rect 2456 17476 2490 17510
rect 2533 17476 2567 17510
rect 2610 17476 2644 17510
rect 2687 17476 2721 17510
rect 2764 17476 2798 17510
rect 2841 17476 2875 17510
rect 2918 17476 2952 17510
rect 2995 17476 3029 17510
rect 381 17369 415 17403
rect 3021 17395 3055 17429
rect 381 17297 415 17331
rect 381 17225 415 17259
rect 381 17153 415 17187
rect 381 17081 415 17115
rect 381 17009 415 17043
rect 381 16937 415 16971
rect 381 16865 415 16899
rect 381 16793 415 16827
rect 381 16721 415 16755
rect 381 16648 415 16682
rect 381 16575 415 16609
rect 381 16502 415 16536
rect 381 16429 415 16463
rect 381 16356 415 16390
rect 381 16283 415 16317
rect 381 16210 415 16244
rect 381 16137 415 16171
rect 381 16064 415 16098
rect 381 15991 415 16025
rect 381 15918 415 15952
rect 381 15845 415 15879
rect 381 15772 415 15806
rect 381 15699 415 15733
rect 381 15626 415 15660
rect 381 15553 415 15587
rect 381 15480 415 15514
rect 381 15407 415 15441
rect 381 15334 415 15368
rect 381 15261 415 15295
rect 381 15188 415 15222
rect 381 15115 415 15149
rect 381 15042 415 15076
rect 381 14969 415 15003
rect 381 14896 415 14930
rect 381 14823 415 14857
rect 381 14750 415 14784
rect 381 14677 415 14711
rect 381 14604 415 14638
rect 381 14531 415 14565
rect 381 14458 415 14492
rect 381 14385 415 14419
rect 381 14312 415 14346
rect 381 14239 415 14273
rect 381 14166 415 14200
rect 381 14093 415 14127
rect 381 14020 415 14054
rect 381 13947 415 13981
rect 381 13874 415 13908
rect 381 13801 415 13835
rect 381 13728 415 13762
rect 381 13655 415 13689
rect 381 13582 415 13616
rect 381 13509 415 13543
rect 381 13436 415 13470
rect 381 13363 415 13397
rect 381 13290 415 13324
rect 381 13217 415 13251
rect 1701 17360 1735 17394
rect 1701 17287 1735 17321
rect 1701 17214 1735 17248
rect 1701 17141 1735 17175
rect 1701 17068 1735 17102
rect 1701 16995 1735 17029
rect 1701 16922 1735 16956
rect 1701 16849 1735 16883
rect 1701 16776 1735 16810
rect 1701 16703 1735 16737
rect 1701 16630 1735 16664
rect 1701 16557 1735 16591
rect 1701 16484 1735 16518
rect 1701 16411 1735 16445
rect 1701 16338 1735 16372
rect 1701 16265 1735 16299
rect 1701 16192 1735 16226
rect 1701 16119 1735 16153
rect 1701 16046 1735 16080
rect 1701 15973 1735 16007
rect 1701 15900 1735 15934
rect 1701 15827 1735 15861
rect 1701 15754 1735 15788
rect 1701 15681 1735 15715
rect 1701 15608 1735 15642
rect 1701 15535 1735 15569
rect 1701 15462 1735 15496
rect 1701 15389 1735 15423
rect 1701 15316 1735 15350
rect 1701 15243 1735 15277
rect 1701 15170 1735 15204
rect 1701 15097 1735 15131
rect 1701 15024 1735 15058
rect 1701 14951 1735 14985
rect 1701 14878 1735 14912
rect 1701 14805 1735 14839
rect 1701 14732 1735 14766
rect 1701 14659 1735 14693
rect 1701 14586 1735 14620
rect 1701 14513 1735 14547
rect 1701 14440 1735 14474
rect 1701 14367 1735 14401
rect 1701 14294 1735 14328
rect 1701 14221 1735 14255
rect 1701 14148 1735 14182
rect 1701 14075 1735 14109
rect 1701 14002 1735 14036
rect 1701 13929 1735 13963
rect 1701 13856 1735 13890
rect 1701 13783 1735 13817
rect 1701 13710 1735 13744
rect 1701 13637 1735 13671
rect 1701 13564 1735 13598
rect 1701 13490 1735 13524
rect 1701 13416 1735 13450
rect 1701 13342 1735 13376
rect 1701 13268 1735 13302
rect 1701 13194 1735 13228
rect 3021 17322 3055 17356
rect 3021 17249 3055 17283
rect 3021 17176 3055 17210
rect 3021 17103 3055 17137
rect 3021 17030 3055 17064
rect 3021 16957 3055 16991
rect 3021 16884 3055 16918
rect 3021 16811 3055 16845
rect 3021 16738 3055 16772
rect 3021 16665 3055 16699
rect 3021 16592 3055 16626
rect 3021 16519 3055 16553
rect 3021 16446 3055 16480
rect 3021 16373 3055 16407
rect 3021 16300 3055 16334
rect 3021 16227 3055 16261
rect 3021 16154 3055 16188
rect 3021 16081 3055 16115
rect 3021 16008 3055 16042
rect 3021 15935 3055 15969
rect 3021 15862 3055 15896
rect 3021 15789 3055 15823
rect 3021 15716 3055 15750
rect 3021 15643 3055 15677
rect 3021 15570 3055 15604
rect 3021 15497 3055 15531
rect 3021 15424 3055 15458
rect 3021 15351 3055 15385
rect 3021 15278 3055 15312
rect 3021 15205 3055 15239
rect 3021 15132 3055 15166
rect 3021 15059 3055 15093
rect 3021 14986 3055 15020
rect 3021 14913 3055 14947
rect 3021 14840 3055 14874
rect 3021 14767 3055 14801
rect 3021 14694 3055 14728
rect 3021 14621 3055 14655
rect 3021 14548 3055 14582
rect 3021 14475 3055 14509
rect 3021 14402 3055 14436
rect 3021 14329 3055 14363
rect 3021 14256 3055 14290
rect 3021 14183 3055 14217
rect 3021 14110 3055 14144
rect 3021 14037 3055 14071
rect 3021 13964 3055 13998
rect 3021 13891 3055 13925
rect 3021 13818 3055 13852
rect 3021 13745 3055 13779
rect 3021 13672 3055 13706
rect 3021 13599 3055 13633
rect 3021 13526 3055 13560
rect 3021 13453 3055 13487
rect 3021 13380 3055 13414
rect 3021 13307 3055 13341
rect 3021 13234 3055 13268
rect 381 13144 415 13178
rect 381 13071 415 13105
rect 381 12998 415 13032
rect 3021 13161 3055 13195
rect 3021 13088 3055 13122
rect 3021 13014 3055 13048
rect 381 12925 415 12959
rect 381 12852 415 12886
rect 381 12779 415 12813
rect 381 12706 415 12740
rect 381 12633 415 12667
rect 381 12560 415 12594
rect 381 12487 415 12521
rect 381 12414 415 12448
rect 381 11550 415 11584
rect 381 11478 415 11512
rect 381 11406 415 11440
rect 381 11334 415 11368
rect 381 11262 415 11296
rect 381 11190 415 11224
rect 381 11118 415 11152
rect 381 11046 415 11080
rect 381 10974 415 11008
rect 381 10902 415 10936
rect 381 10830 415 10864
rect 381 10758 415 10792
rect 381 10686 415 10720
rect 381 10614 415 10648
rect 381 10542 415 10576
rect 381 10470 415 10504
rect 381 10398 415 10432
rect 381 10326 415 10360
rect 381 10254 415 10288
rect 381 10182 415 10216
rect 381 10110 415 10144
rect 381 10038 415 10072
rect 381 9966 415 10000
rect 381 9894 415 9928
rect 381 9822 415 9856
rect 381 9750 415 9784
rect 381 9678 415 9712
rect 381 9606 415 9640
rect 381 9534 415 9568
rect 381 9462 415 9496
rect 381 9390 415 9424
rect 381 9318 415 9352
rect 381 9246 415 9280
rect 381 9174 415 9208
rect 381 9102 415 9136
rect 381 9030 415 9064
rect 381 8958 415 8992
rect 381 8886 415 8920
rect 381 8814 415 8848
rect 381 8742 415 8776
rect 381 8670 415 8704
rect 381 8598 415 8632
rect 381 8526 415 8560
rect 381 8454 415 8488
rect 381 8382 415 8416
rect 381 8310 415 8344
rect 381 8238 415 8272
rect 381 8166 415 8200
rect 381 8094 415 8128
rect 381 8022 415 8056
rect 381 7950 415 7984
rect 381 7878 415 7912
rect 381 7806 415 7840
rect 381 7734 415 7768
rect 381 7662 415 7696
rect 381 7590 415 7624
rect 381 7518 415 7552
rect 381 7446 415 7480
rect 381 7374 415 7408
rect 381 7302 415 7336
rect 381 7230 415 7264
rect 381 7158 415 7192
rect 381 7086 415 7120
rect 381 7014 415 7048
rect 381 6942 415 6976
rect 381 6870 415 6904
rect 381 6798 415 6832
rect 381 6726 415 6760
rect 381 6654 415 6688
rect 381 6582 415 6616
rect 381 6510 415 6544
rect 381 6438 415 6472
rect 381 6366 415 6400
rect 381 6294 415 6328
rect 381 6222 415 6256
rect 381 6150 415 6184
rect 381 6078 415 6112
rect 381 6006 415 6040
rect 381 5934 415 5968
rect 381 5862 415 5896
rect 381 5790 415 5824
rect 381 5718 415 5752
rect 381 5646 415 5680
rect 381 5574 415 5608
rect 381 5502 415 5536
rect 381 5430 415 5464
rect 381 5358 415 5392
rect 381 5286 415 5320
rect 381 5214 415 5248
rect 381 5142 415 5176
rect 381 5070 415 5104
rect 381 4998 415 5032
rect 381 4926 415 4960
rect 381 4854 415 4888
rect 381 4782 415 4816
rect 381 4710 415 4744
rect 381 4638 415 4672
rect 381 4566 415 4600
rect 381 4494 415 4528
rect 381 4422 415 4456
rect 381 4350 415 4384
rect 381 4278 415 4312
rect 381 4206 415 4240
rect 3021 10316 3055 10350
rect 3021 10244 3055 10278
rect 3021 10172 3055 10206
rect 3021 10100 3055 10134
rect 3021 10028 3055 10062
rect 3021 9956 3055 9990
rect 3021 9884 3055 9918
rect 3021 9812 3055 9846
rect 3021 9740 3055 9774
rect 3021 9668 3055 9702
rect 3021 9596 3055 9630
rect 3021 9524 3055 9558
rect 3021 9452 3055 9486
rect 3021 9380 3055 9414
rect 3021 9308 3055 9342
rect 3021 9236 3055 9270
rect 3021 9164 3055 9198
rect 3021 9092 3055 9126
rect 3021 9020 3055 9054
rect 3021 8948 3055 8982
rect 3021 8876 3055 8910
rect 3021 8804 3055 8838
rect 3021 8732 3055 8766
rect 3021 8660 3055 8694
rect 3021 8588 3055 8622
rect 3021 8516 3055 8550
rect 3021 8444 3055 8478
rect 3021 8372 3055 8406
rect 3021 8300 3055 8334
rect 3021 8228 3055 8262
rect 3021 8156 3055 8190
rect 3021 8084 3055 8118
rect 3021 8012 3055 8046
rect 3021 7940 3055 7974
rect 3021 7868 3055 7902
rect 3021 7796 3055 7830
rect 3021 7724 3055 7758
rect 3021 7652 3055 7686
rect 3021 7580 3055 7614
rect 3021 7508 3055 7542
rect 3021 7436 3055 7470
rect 3021 7364 3055 7398
rect 3021 7292 3055 7326
rect 3021 7220 3055 7254
rect 3021 7148 3055 7182
rect 3021 7076 3055 7110
rect 3021 7004 3055 7038
rect 3021 6932 3055 6966
rect 3021 6860 3055 6894
rect 3021 6788 3055 6822
rect 3021 6716 3055 6750
rect 3021 6644 3055 6678
rect 3021 6572 3055 6606
rect 3021 6500 3055 6534
rect 3021 6428 3055 6462
rect 3021 6356 3055 6390
rect 3021 6284 3055 6318
rect 3021 6212 3055 6246
rect 3021 6140 3055 6174
rect 3021 6068 3055 6102
rect 3021 5996 3055 6030
rect 3021 5924 3055 5958
rect 3021 5852 3055 5886
rect 3021 5780 3055 5814
rect 3021 5708 3055 5742
rect 3021 5636 3055 5670
rect 3021 5564 3055 5598
rect 3021 5492 3055 5526
rect 3021 5420 3055 5454
rect 3021 5348 3055 5382
rect 3021 5275 3055 5309
rect 3021 5202 3055 5236
rect 3021 5129 3055 5163
rect 3021 5056 3055 5090
rect 3021 4983 3055 5017
rect 3021 4910 3055 4944
rect 3021 4837 3055 4871
rect 3021 4764 3055 4798
rect 3021 4691 3055 4725
rect 3021 4618 3055 4652
rect 3021 4545 3055 4579
rect 3021 4472 3055 4506
rect 3021 4399 3055 4433
rect 3021 4326 3055 4360
rect 3021 4253 3055 4287
rect 3021 4180 3055 4214
rect 381 4134 415 4168
rect 381 4061 415 4095
rect 381 3988 415 4022
rect 381 3915 415 3949
rect 381 3842 415 3876
rect 381 3769 415 3803
rect 381 3696 415 3730
rect 381 3623 415 3657
rect 381 3550 415 3584
rect 381 3477 415 3511
rect 381 3404 415 3438
rect 381 3331 415 3365
rect 381 3258 415 3292
rect 381 3185 415 3219
rect 381 3112 415 3146
rect 381 3039 415 3073
rect 381 2966 415 3000
rect 381 2893 415 2927
rect 381 2820 415 2854
rect 381 2747 415 2781
rect 381 2674 415 2708
rect 381 2601 415 2635
rect 381 2528 415 2562
rect 381 2455 415 2489
rect 381 2382 415 2416
rect 381 2309 415 2343
rect 381 2236 415 2270
rect 381 2163 415 2197
rect 381 2090 415 2124
rect 381 2017 415 2051
rect 381 1944 415 1978
rect 381 1871 415 1905
rect 381 1798 415 1832
rect 381 1725 415 1759
rect 381 1652 415 1686
rect 381 1579 415 1613
rect 381 1506 415 1540
rect 381 1433 415 1467
rect 381 1360 415 1394
rect 381 1287 415 1321
rect 381 1214 415 1248
rect 381 1141 415 1175
rect 381 1068 415 1102
rect 381 995 415 1029
rect 381 922 415 956
rect 1701 3608 1735 3642
rect 1701 3536 1735 3570
rect 1701 3464 1735 3498
rect 1701 3392 1735 3426
rect 1701 3320 1735 3354
rect 1701 3248 1735 3282
rect 1701 3176 1735 3210
rect 1701 3104 1735 3138
rect 1701 3032 1735 3066
rect 1701 2960 1735 2994
rect 1701 2888 1735 2922
rect 1701 2816 1735 2850
rect 1701 2744 1735 2778
rect 1701 2672 1735 2706
rect 1701 2600 1735 2634
rect 1701 2528 1735 2562
rect 1701 2456 1735 2490
rect 1701 2384 1735 2418
rect 1701 2312 1735 2346
rect 1701 2240 1735 2274
rect 1701 2168 1735 2202
rect 1701 2096 1735 2130
rect 1701 2024 1735 2058
rect 3201 2345 3235 2379
rect 3273 2345 3281 2379
rect 3281 2345 3307 2379
rect 3345 2345 3349 2379
rect 3349 2345 3379 2379
rect 3198 2277 3232 2305
rect 3198 2271 3232 2277
rect 3198 2209 3232 2233
rect 3198 2199 3232 2209
rect 3350 2226 3384 2260
rect 3422 2226 3456 2260
rect 3494 2226 3528 2260
rect 3566 2226 3600 2260
rect 3638 2226 3672 2260
rect 3198 2141 3232 2161
rect 3198 2127 3232 2141
rect 3198 2073 3232 2089
rect 3198 2055 3232 2073
rect 3946 2199 3980 2231
rect 3946 2197 3980 2199
rect 3946 2130 3980 2159
rect 3946 2125 3980 2130
rect 3627 2070 3661 2104
rect 3699 2070 3733 2104
rect 3771 2070 3805 2104
rect 3843 2070 3877 2104
rect 1701 1952 1735 1986
rect 1701 1880 1735 1914
rect 1701 1808 1735 1842
rect 1701 1736 1735 1770
rect 3350 1914 3384 1948
rect 3422 1914 3456 1948
rect 3494 1914 3528 1948
rect 3566 1914 3600 1948
rect 3638 1914 3672 1948
rect 3584 1758 3618 1792
rect 3656 1758 3690 1792
rect 3728 1758 3762 1792
rect 3800 1758 3834 1792
rect 3872 1758 3906 1792
rect 1701 1664 1735 1698
rect 1701 1592 1735 1626
rect 1701 1520 1735 1554
rect 1701 1448 1735 1482
rect 1701 1376 1735 1410
rect 1701 1304 1735 1338
rect 1701 1232 1735 1266
rect 1701 1160 1735 1194
rect 1701 1088 1735 1122
rect 1701 1016 1735 1050
rect 3198 1699 3232 1718
rect 3198 1684 3232 1699
rect 3198 1631 3232 1646
rect 3198 1612 3232 1631
rect 3350 1602 3384 1636
rect 3422 1602 3456 1636
rect 3494 1602 3528 1636
rect 3566 1602 3600 1636
rect 3638 1602 3672 1636
rect 3198 1563 3232 1574
rect 3198 1540 3232 1563
rect 3198 1495 3232 1502
rect 3198 1468 3232 1495
rect 3584 1446 3618 1480
rect 3656 1446 3690 1480
rect 3728 1446 3762 1480
rect 3800 1446 3834 1480
rect 3872 1446 3906 1480
rect 3198 1427 3232 1430
rect 3198 1396 3232 1427
rect 3198 1325 3232 1358
rect 3198 1324 3232 1325
rect 3198 1257 3232 1286
rect 3198 1252 3232 1257
rect 3350 1290 3384 1324
rect 3422 1290 3456 1324
rect 3494 1290 3528 1324
rect 3566 1290 3600 1324
rect 3638 1290 3672 1324
rect 3198 1189 3232 1214
rect 3198 1180 3232 1189
rect 3198 1121 3232 1142
rect 3198 1108 3232 1121
rect 3584 1154 3618 1188
rect 3656 1154 3690 1188
rect 3728 1154 3762 1188
rect 3800 1154 3834 1188
rect 3872 1154 3906 1188
rect 3201 1016 3235 1050
rect 3273 1016 3300 1050
rect 3300 1016 3307 1050
rect 3345 1016 3368 1050
rect 3368 1016 3379 1050
rect 1701 944 1735 978
rect 1701 872 1735 906
rect 1701 800 1735 834
rect 1701 728 1735 762
rect 1701 656 1735 690
rect 381 584 415 618
rect 381 496 415 530
rect 381 408 415 442
rect 381 319 415 353
rect 1701 583 1735 617
rect 1701 510 1735 544
rect 1701 437 1735 471
rect 1701 364 1735 398
rect 3576 565 3610 587
rect 3576 553 3610 565
rect 3576 497 3610 511
rect 3576 477 3610 497
rect 3576 429 3610 436
rect 3576 402 3610 429
rect 3576 327 3610 361
rect 3576 259 3610 286
rect 3576 252 3610 259
rect 393 216 427 250
rect 466 216 500 250
rect 539 216 573 250
rect 612 216 646 250
rect 685 216 719 250
rect 758 216 792 250
rect 831 216 865 250
rect 904 216 938 250
rect 977 216 1011 250
rect 1050 216 1084 250
rect 1123 216 1157 250
rect 1196 216 1230 250
rect 1269 216 1303 250
rect 1342 216 1376 250
rect 1415 216 1449 250
rect 1488 216 1522 250
rect 1561 216 1595 250
rect 1634 216 1668 250
rect 1707 216 1741 250
rect 1780 216 1814 250
rect 1853 216 1887 250
rect 1926 216 1960 250
rect 1999 216 2033 250
rect 2072 216 2106 250
rect 2145 216 2179 250
rect 2217 216 2251 250
rect 2289 216 2323 250
rect 2361 216 2395 250
rect 2433 216 2467 250
rect 2505 216 2539 250
rect 2577 216 2611 250
rect 2649 216 2683 250
rect 2721 216 2755 250
rect 2793 216 2827 250
rect 2865 216 2899 250
rect 2937 216 2971 250
rect 3009 216 3043 250
rect 3576 191 3610 211
rect 3576 177 3610 191
rect 3576 123 3610 136
rect 3576 102 3610 123
rect 3576 27 3577 61
rect 3577 27 3610 61
<< metal1 >>
rect 49 17656 2744 17862
rect 49 17596 2176 17602
rect 49 17550 2124 17596
tri 2096 17522 2124 17550 ne
rect 2124 17532 2176 17544
rect 375 17510 2047 17516
rect 375 17476 407 17510
rect 441 17476 482 17510
rect 516 17476 557 17510
rect 591 17476 632 17510
rect 666 17476 707 17510
rect 741 17476 782 17510
rect 816 17476 857 17510
rect 891 17476 932 17510
rect 966 17476 1007 17510
rect 1041 17476 1082 17510
rect 1116 17476 1157 17510
rect 1191 17476 1232 17510
rect 1266 17476 1307 17510
rect 1341 17476 1382 17510
rect 1416 17476 1457 17510
rect 1491 17476 1532 17510
rect 1566 17476 1607 17510
rect 1641 17476 1682 17510
rect 1716 17476 1757 17510
rect 1791 17476 1832 17510
rect 1866 17476 1907 17510
rect 1941 17476 1981 17510
rect 2015 17476 2047 17510
rect 375 17470 2047 17476
rect 2124 17474 2176 17480
rect 2268 17510 3061 17516
rect 2268 17476 2300 17510
rect 2334 17476 2378 17510
rect 2412 17476 2456 17510
rect 2490 17476 2533 17510
rect 2567 17476 2610 17510
rect 2644 17476 2687 17510
rect 2721 17476 2764 17510
rect 2798 17476 2841 17510
rect 2875 17476 2918 17510
rect 2952 17476 2995 17510
rect 3029 17476 3061 17510
rect 2268 17470 3061 17476
rect 375 17403 421 17470
rect 375 17369 381 17403
rect 415 17369 421 17403
rect 375 17331 421 17369
rect 375 17297 381 17331
rect 415 17297 421 17331
rect 375 17259 421 17297
rect 375 17225 381 17259
rect 415 17225 421 17259
rect 375 17187 421 17225
rect 375 17153 381 17187
rect 415 17153 421 17187
rect 375 17115 421 17153
rect 375 17081 381 17115
rect 415 17081 421 17115
rect 375 17043 421 17081
rect 375 17009 381 17043
rect 415 17009 421 17043
rect 375 16971 421 17009
rect 375 16937 381 16971
rect 415 16937 421 16971
rect 375 16899 421 16937
rect 375 16865 381 16899
rect 415 16865 421 16899
rect 375 16827 421 16865
rect 375 16793 381 16827
rect 415 16793 421 16827
rect 375 16755 421 16793
rect 375 16721 381 16755
rect 415 16721 421 16755
rect 375 16682 421 16721
rect 375 16648 381 16682
rect 415 16648 421 16682
rect 375 16609 421 16648
rect 375 16575 381 16609
rect 415 16575 421 16609
rect 375 16536 421 16575
rect 375 16502 381 16536
rect 415 16502 421 16536
rect 375 16463 421 16502
rect 375 16429 381 16463
rect 415 16429 421 16463
rect 375 16390 421 16429
rect 375 16356 381 16390
rect 415 16356 421 16390
rect 375 16317 421 16356
rect 375 16283 381 16317
rect 415 16283 421 16317
rect 375 16244 421 16283
rect 375 16210 381 16244
rect 415 16210 421 16244
rect 375 16171 421 16210
rect 375 16137 381 16171
rect 415 16137 421 16171
rect 375 16098 421 16137
rect 375 16064 381 16098
rect 415 16064 421 16098
rect 375 16025 421 16064
rect 375 15991 381 16025
rect 415 15991 421 16025
rect 375 15952 421 15991
rect 375 15918 381 15952
rect 415 15918 421 15952
rect 375 15879 421 15918
rect 375 15845 381 15879
rect 415 15845 421 15879
rect 375 15806 421 15845
rect 375 15772 381 15806
rect 415 15772 421 15806
rect 375 15733 421 15772
rect 375 15699 381 15733
rect 415 15699 421 15733
rect 375 15660 421 15699
rect 375 15626 381 15660
rect 415 15626 421 15660
rect 375 15587 421 15626
rect 375 15553 381 15587
rect 415 15553 421 15587
rect 375 15514 421 15553
rect 375 15480 381 15514
rect 415 15480 421 15514
rect 375 15441 421 15480
rect 375 15407 381 15441
rect 415 15407 421 15441
rect 375 15368 421 15407
rect 375 15334 381 15368
rect 415 15334 421 15368
rect 375 15295 421 15334
rect 375 15261 381 15295
rect 415 15261 421 15295
rect 375 15222 421 15261
rect 375 15188 381 15222
rect 415 15188 421 15222
rect 375 15149 421 15188
rect 375 15115 381 15149
rect 415 15115 421 15149
rect 375 15076 421 15115
rect 375 15042 381 15076
rect 415 15042 421 15076
rect 375 15003 421 15042
rect 375 14969 381 15003
rect 415 14969 421 15003
rect 375 14930 421 14969
rect 375 14896 381 14930
rect 415 14896 421 14930
rect 375 14857 421 14896
rect 375 14823 381 14857
rect 415 14823 421 14857
rect 375 14784 421 14823
rect 375 14750 381 14784
rect 415 14750 421 14784
rect 375 14711 421 14750
rect 375 14677 381 14711
rect 415 14677 421 14711
rect 375 14638 421 14677
rect 375 14604 381 14638
rect 415 14604 421 14638
rect 375 14565 421 14604
rect 375 14531 381 14565
rect 415 14531 421 14565
rect 375 14492 421 14531
rect 375 14458 381 14492
rect 415 14458 421 14492
rect 375 14419 421 14458
rect 375 14385 381 14419
rect 415 14385 421 14419
rect 375 14346 421 14385
rect 375 14312 381 14346
rect 415 14312 421 14346
rect 375 14273 421 14312
rect 375 14239 381 14273
rect 415 14239 421 14273
rect 375 14200 421 14239
rect 375 14166 381 14200
rect 415 14166 421 14200
rect 375 14127 421 14166
rect 375 14093 381 14127
rect 415 14093 421 14127
rect 375 14054 421 14093
rect 375 14020 381 14054
rect 415 14020 421 14054
rect 375 13981 421 14020
rect 375 13947 381 13981
rect 415 13947 421 13981
rect 375 13908 421 13947
rect 375 13874 381 13908
rect 415 13874 421 13908
rect 375 13835 421 13874
rect 375 13801 381 13835
rect 415 13801 421 13835
rect 375 13762 421 13801
rect 375 13728 381 13762
rect 415 13728 421 13762
rect 375 13689 421 13728
rect 375 13655 381 13689
rect 415 13655 421 13689
rect 375 13616 421 13655
rect 375 13582 381 13616
rect 415 13582 421 13616
rect 375 13543 421 13582
rect 375 13509 381 13543
rect 415 13509 421 13543
rect 375 13470 421 13509
rect 375 13436 381 13470
rect 415 13436 421 13470
rect 375 13397 421 13436
rect 375 13363 381 13397
rect 415 13363 421 13397
rect 375 13324 421 13363
rect 375 13290 381 13324
rect 415 13290 421 13324
rect 375 13251 421 13290
rect 375 13217 381 13251
rect 415 13217 421 13251
rect 375 13178 421 13217
rect 1695 17394 1741 17470
rect 1695 17360 1701 17394
rect 1735 17360 1741 17394
rect 1695 17321 1741 17360
rect 1695 17287 1701 17321
rect 1735 17287 1741 17321
rect 1695 17248 1741 17287
rect 1695 17214 1701 17248
rect 1735 17214 1741 17248
rect 1695 17175 1741 17214
rect 1695 17141 1701 17175
rect 1735 17141 1741 17175
rect 1695 17102 1741 17141
rect 1695 17068 1701 17102
rect 1735 17068 1741 17102
rect 1695 17029 1741 17068
rect 1695 16995 1701 17029
rect 1735 16995 1741 17029
rect 1695 16956 1741 16995
rect 1695 16922 1701 16956
rect 1735 16922 1741 16956
rect 1695 16883 1741 16922
rect 1695 16849 1701 16883
rect 1735 16849 1741 16883
rect 1695 16810 1741 16849
rect 1695 16776 1701 16810
rect 1735 16776 1741 16810
rect 1695 16737 1741 16776
rect 1695 16703 1701 16737
rect 1735 16703 1741 16737
rect 1695 16664 1741 16703
rect 1695 16630 1701 16664
rect 1735 16630 1741 16664
rect 1695 16591 1741 16630
rect 1695 16557 1701 16591
rect 1735 16557 1741 16591
rect 1695 16518 1741 16557
rect 1695 16484 1701 16518
rect 1735 16484 1741 16518
rect 1695 16445 1741 16484
rect 1695 16411 1701 16445
rect 1735 16411 1741 16445
rect 1695 16372 1741 16411
rect 1695 16338 1701 16372
rect 1735 16338 1741 16372
rect 1695 16299 1741 16338
rect 1695 16265 1701 16299
rect 1735 16265 1741 16299
rect 1695 16226 1741 16265
rect 1695 16192 1701 16226
rect 1735 16192 1741 16226
rect 1695 16153 1741 16192
rect 1695 16119 1701 16153
rect 1735 16119 1741 16153
rect 1695 16080 1741 16119
rect 1695 16046 1701 16080
rect 1735 16046 1741 16080
rect 1695 16007 1741 16046
rect 1695 15973 1701 16007
rect 1735 15973 1741 16007
rect 1695 15934 1741 15973
rect 1695 15900 1701 15934
rect 1735 15900 1741 15934
rect 1695 15861 1741 15900
rect 1695 15827 1701 15861
rect 1735 15827 1741 15861
rect 1695 15788 1741 15827
rect 1695 15754 1701 15788
rect 1735 15754 1741 15788
rect 1695 15715 1741 15754
rect 1695 15681 1701 15715
rect 1735 15681 1741 15715
rect 1695 15642 1741 15681
rect 1695 15608 1701 15642
rect 1735 15608 1741 15642
rect 1695 15569 1741 15608
rect 1695 15535 1701 15569
rect 1735 15535 1741 15569
rect 1695 15496 1741 15535
rect 1695 15462 1701 15496
rect 1735 15462 1741 15496
rect 1695 15423 1741 15462
rect 1695 15389 1701 15423
rect 1735 15389 1741 15423
rect 1695 15350 1741 15389
rect 1695 15316 1701 15350
rect 1735 15316 1741 15350
rect 1695 15277 1741 15316
rect 1695 15243 1701 15277
rect 1735 15243 1741 15277
rect 1695 15204 1741 15243
rect 1695 15170 1701 15204
rect 1735 15170 1741 15204
rect 1695 15131 1741 15170
rect 1695 15097 1701 15131
rect 1735 15097 1741 15131
rect 1695 15058 1741 15097
rect 1695 15024 1701 15058
rect 1735 15024 1741 15058
rect 1695 14985 1741 15024
rect 1695 14951 1701 14985
rect 1735 14951 1741 14985
rect 1695 14912 1741 14951
rect 1695 14878 1701 14912
rect 1735 14878 1741 14912
rect 1695 14839 1741 14878
rect 1695 14805 1701 14839
rect 1735 14805 1741 14839
rect 1695 14766 1741 14805
rect 1695 14732 1701 14766
rect 1735 14732 1741 14766
rect 1695 14693 1741 14732
rect 1695 14659 1701 14693
rect 1735 14659 1741 14693
rect 1695 14620 1741 14659
rect 1695 14586 1701 14620
rect 1735 14586 1741 14620
rect 1695 14547 1741 14586
rect 1695 14513 1701 14547
rect 1735 14513 1741 14547
rect 1695 14474 1741 14513
rect 1695 14440 1701 14474
rect 1735 14440 1741 14474
rect 1695 14401 1741 14440
rect 1695 14367 1701 14401
rect 1735 14367 1741 14401
rect 1695 14328 1741 14367
rect 1695 14294 1701 14328
rect 1735 14294 1741 14328
rect 1695 14255 1741 14294
rect 1695 14221 1701 14255
rect 1735 14221 1741 14255
rect 1695 14182 1741 14221
rect 1695 14148 1701 14182
rect 1735 14148 1741 14182
rect 1695 14109 1741 14148
rect 1695 14075 1701 14109
rect 1735 14075 1741 14109
rect 1695 14036 1741 14075
rect 1695 14002 1701 14036
rect 1735 14002 1741 14036
rect 1695 13963 1741 14002
rect 1695 13929 1701 13963
rect 1735 13929 1741 13963
rect 1695 13890 1741 13929
rect 1695 13856 1701 13890
rect 1735 13856 1741 13890
rect 1695 13817 1741 13856
rect 1695 13783 1701 13817
rect 1735 13783 1741 13817
rect 1695 13744 1741 13783
rect 1695 13710 1701 13744
rect 1735 13710 1741 13744
rect 1695 13671 1741 13710
rect 1695 13637 1701 13671
rect 1735 13637 1741 13671
rect 1695 13598 1741 13637
rect 1695 13564 1701 13598
rect 1735 13564 1741 13598
rect 1695 13524 1741 13564
rect 1695 13490 1701 13524
rect 1735 13490 1741 13524
rect 1695 13450 1741 13490
rect 1695 13416 1701 13450
rect 1735 13416 1741 13450
rect 1695 13376 1741 13416
rect 1695 13342 1701 13376
rect 1735 13342 1741 13376
rect 1695 13302 1741 13342
rect 1695 13268 1701 13302
rect 1735 13268 1741 13302
rect 1695 13228 1741 13268
rect 1695 13194 1701 13228
rect 1735 13194 1741 13228
rect 1695 13182 1741 13194
rect 3015 17429 3061 17470
rect 3015 17395 3021 17429
rect 3055 17395 3061 17429
rect 3015 17356 3061 17395
rect 3015 17322 3021 17356
rect 3055 17322 3061 17356
rect 3015 17283 3061 17322
rect 3015 17249 3021 17283
rect 3055 17249 3061 17283
rect 3015 17210 3061 17249
rect 3015 17176 3021 17210
rect 3055 17176 3061 17210
rect 3015 17137 3061 17176
rect 3015 17103 3021 17137
rect 3055 17103 3061 17137
rect 3015 17064 3061 17103
rect 3015 17030 3021 17064
rect 3055 17030 3061 17064
rect 3015 16991 3061 17030
rect 3015 16957 3021 16991
rect 3055 16957 3061 16991
rect 3015 16918 3061 16957
rect 3015 16884 3021 16918
rect 3055 16884 3061 16918
rect 3015 16845 3061 16884
rect 3015 16811 3021 16845
rect 3055 16811 3061 16845
rect 3015 16772 3061 16811
rect 3015 16738 3021 16772
rect 3055 16738 3061 16772
rect 3015 16699 3061 16738
rect 3015 16665 3021 16699
rect 3055 16665 3061 16699
rect 3015 16626 3061 16665
rect 3015 16592 3021 16626
rect 3055 16592 3061 16626
rect 3015 16553 3061 16592
rect 3015 16519 3021 16553
rect 3055 16519 3061 16553
rect 3015 16480 3061 16519
rect 3015 16446 3021 16480
rect 3055 16446 3061 16480
rect 3015 16407 3061 16446
rect 3015 16373 3021 16407
rect 3055 16373 3061 16407
rect 3015 16334 3061 16373
rect 3015 16300 3021 16334
rect 3055 16300 3061 16334
rect 3015 16261 3061 16300
rect 3015 16227 3021 16261
rect 3055 16227 3061 16261
rect 3015 16188 3061 16227
rect 3015 16154 3021 16188
rect 3055 16154 3061 16188
rect 3015 16115 3061 16154
rect 3015 16081 3021 16115
rect 3055 16081 3061 16115
rect 3015 16042 3061 16081
rect 3015 16008 3021 16042
rect 3055 16008 3061 16042
rect 3015 15969 3061 16008
rect 3015 15935 3021 15969
rect 3055 15935 3061 15969
rect 3015 15896 3061 15935
rect 3015 15862 3021 15896
rect 3055 15862 3061 15896
rect 3015 15823 3061 15862
rect 3015 15789 3021 15823
rect 3055 15789 3061 15823
rect 3015 15750 3061 15789
rect 3015 15716 3021 15750
rect 3055 15716 3061 15750
rect 3015 15677 3061 15716
rect 3015 15643 3021 15677
rect 3055 15643 3061 15677
rect 3015 15604 3061 15643
rect 3015 15570 3021 15604
rect 3055 15570 3061 15604
rect 3015 15531 3061 15570
rect 3015 15497 3021 15531
rect 3055 15497 3061 15531
rect 3015 15458 3061 15497
rect 3015 15424 3021 15458
rect 3055 15424 3061 15458
rect 3015 15385 3061 15424
rect 3015 15351 3021 15385
rect 3055 15351 3061 15385
rect 3015 15312 3061 15351
rect 3015 15278 3021 15312
rect 3055 15278 3061 15312
rect 3015 15239 3061 15278
rect 3015 15205 3021 15239
rect 3055 15205 3061 15239
rect 3015 15166 3061 15205
rect 3015 15132 3021 15166
rect 3055 15132 3061 15166
rect 3015 15093 3061 15132
rect 3015 15059 3021 15093
rect 3055 15059 3061 15093
rect 3015 15020 3061 15059
rect 3015 14986 3021 15020
rect 3055 14986 3061 15020
rect 3015 14947 3061 14986
rect 3015 14913 3021 14947
rect 3055 14913 3061 14947
rect 3015 14874 3061 14913
rect 3015 14840 3021 14874
rect 3055 14840 3061 14874
rect 3015 14801 3061 14840
rect 3015 14767 3021 14801
rect 3055 14767 3061 14801
rect 3015 14728 3061 14767
rect 3015 14694 3021 14728
rect 3055 14694 3061 14728
rect 3015 14655 3061 14694
rect 3015 14621 3021 14655
rect 3055 14621 3061 14655
rect 3015 14582 3061 14621
rect 3015 14548 3021 14582
rect 3055 14548 3061 14582
rect 3015 14509 3061 14548
rect 3015 14475 3021 14509
rect 3055 14475 3061 14509
rect 3015 14436 3061 14475
rect 3015 14402 3021 14436
rect 3055 14402 3061 14436
rect 3015 14363 3061 14402
rect 3015 14329 3021 14363
rect 3055 14329 3061 14363
rect 3015 14290 3061 14329
rect 3015 14256 3021 14290
rect 3055 14256 3061 14290
rect 3015 14217 3061 14256
rect 3015 14183 3021 14217
rect 3055 14183 3061 14217
rect 3015 14144 3061 14183
rect 3015 14110 3021 14144
rect 3055 14110 3061 14144
rect 3015 14071 3061 14110
rect 3015 14037 3021 14071
rect 3055 14037 3061 14071
rect 3015 13998 3061 14037
rect 3015 13964 3021 13998
rect 3055 13964 3061 13998
rect 3015 13925 3061 13964
rect 3015 13891 3021 13925
rect 3055 13891 3061 13925
rect 3015 13852 3061 13891
rect 3015 13818 3021 13852
rect 3055 13818 3061 13852
rect 3015 13779 3061 13818
rect 3015 13745 3021 13779
rect 3055 13745 3061 13779
rect 3015 13706 3061 13745
rect 3015 13672 3021 13706
rect 3055 13672 3061 13706
rect 3015 13633 3061 13672
rect 3015 13599 3021 13633
rect 3055 13599 3061 13633
rect 3015 13560 3061 13599
rect 3015 13526 3021 13560
rect 3055 13526 3061 13560
rect 3015 13487 3061 13526
rect 3015 13453 3021 13487
rect 3055 13453 3061 13487
rect 3015 13414 3061 13453
rect 3015 13380 3021 13414
rect 3055 13380 3061 13414
rect 3015 13341 3061 13380
rect 3015 13307 3021 13341
rect 3055 13307 3061 13341
rect 3015 13268 3061 13307
rect 3015 13234 3021 13268
rect 3055 13234 3061 13268
rect 3015 13195 3061 13234
rect 375 13144 381 13178
rect 415 13144 421 13178
rect 375 13105 421 13144
rect 375 13071 381 13105
rect 415 13071 421 13105
rect 375 13032 421 13071
rect 375 12998 381 13032
rect 415 12998 421 13032
rect 3015 13161 3021 13195
rect 3055 13161 3061 13195
rect 3015 13122 3061 13161
rect 3015 13088 3021 13122
rect 3055 13088 3061 13122
rect 3015 13048 3061 13088
rect 3015 13014 3021 13048
rect 3055 13014 3061 13048
rect 3015 13002 3061 13014
rect 375 12959 421 12998
rect 375 12925 381 12959
rect 415 12925 421 12959
rect 375 12886 421 12925
rect 375 12852 381 12886
rect 415 12852 421 12886
rect 375 12813 421 12852
rect 375 12779 381 12813
rect 415 12779 421 12813
rect 375 12740 421 12779
rect 375 12706 381 12740
rect 415 12706 421 12740
rect 375 12667 421 12706
rect 375 12633 381 12667
rect 415 12633 421 12667
rect 375 12594 421 12633
rect 375 12560 381 12594
rect 415 12560 421 12594
rect 375 12521 421 12560
rect 375 12487 381 12521
rect 415 12487 421 12521
rect 375 12448 421 12487
rect 375 12414 381 12448
rect 415 12414 421 12448
rect 375 12402 421 12414
tri 237 12260 301 12324 se
rect 301 12318 359 12324
rect 301 12266 304 12318
rect 356 12266 359 12318
rect 301 12260 359 12266
rect 0 12254 359 12260
rect 0 12202 304 12254
rect 356 12202 359 12254
rect 0 12196 359 12202
tri 1963 12196 1987 12220 se
rect 1987 12214 2045 12220
rect 1987 12196 1990 12214
tri 1923 12156 1963 12196 se
rect 1963 12162 1990 12196
rect 2042 12162 2045 12214
rect 1963 12156 2045 12162
rect 0 12150 2045 12156
rect 0 12098 1990 12150
rect 2042 12098 2045 12150
rect 0 12092 2045 12098
tri 84 11771 150 11837 se
rect 150 11791 421 11837
tri 421 11791 467 11837 sw
tri 150 11771 170 11791 nw
tri 401 11771 421 11791 ne
rect 421 11771 467 11791
tri 18 11705 84 11771 se
tri 84 11705 150 11771 nw
tri 421 11725 467 11771 ne
tri 467 11725 533 11791 sw
tri 1893 11725 1916 11748 se
rect 1916 11725 2316 11748
tri 467 11705 487 11725 ne
rect 487 11705 533 11725
tri -7 11680 18 11705 se
rect 18 11680 39 11705
rect -389 2938 -306 2984
tri -389 2927 -378 2938 ne
rect -378 2927 -306 2938
tri -378 2901 -352 2927 ne
rect -352 2901 -306 2927
rect -1262 2583 -772 2609
rect -1262 2558 -824 2583
tri -850 2532 -824 2558 ne
rect -824 2519 -772 2531
rect -824 2461 -772 2467
rect -7 216 39 11680
tri 39 11660 84 11705 nw
tri 487 11660 532 11705 ne
rect 532 11660 533 11705
tri 532 11659 533 11660 ne
tri 533 11659 599 11725 sw
tri 1850 11682 1893 11725 se
rect 1893 11702 2316 11725
rect 1893 11682 1916 11702
tri 1916 11682 1936 11702 nw
tri 1827 11659 1850 11682 se
tri 533 11596 596 11659 ne
rect 596 11596 599 11659
rect 375 11584 421 11596
tri 596 11593 599 11596 ne
tri 599 11593 665 11659 sw
tri 1784 11616 1827 11659 se
rect 1827 11616 1850 11659
tri 1850 11616 1916 11682 nw
tri 1761 11593 1784 11616 se
rect 1784 11593 1827 11616
tri 1827 11593 1850 11616 nw
rect 375 11550 381 11584
rect 415 11550 421 11584
rect 375 11512 421 11550
tri 599 11547 645 11593 ne
rect 645 11547 1781 11593
tri 1781 11547 1827 11593 nw
rect 375 11478 381 11512
rect 415 11478 421 11512
rect 375 11440 421 11478
rect 375 11406 381 11440
rect 415 11406 421 11440
rect 375 11368 421 11406
rect 375 11334 381 11368
rect 415 11334 421 11368
rect 375 11296 421 11334
rect 375 11262 381 11296
rect 415 11262 421 11296
rect 375 11224 421 11262
rect 375 11190 381 11224
rect 415 11190 421 11224
rect 375 11152 421 11190
rect 375 11118 381 11152
rect 415 11118 421 11152
rect 375 11080 421 11118
rect 375 11046 381 11080
rect 415 11046 421 11080
rect 375 11008 421 11046
rect 375 10974 381 11008
rect 415 10974 421 11008
rect 375 10936 421 10974
rect 375 10902 381 10936
rect 415 10902 421 10936
rect 375 10864 421 10902
rect 375 10830 381 10864
rect 415 10830 421 10864
rect 375 10792 421 10830
rect 375 10758 381 10792
rect 415 10758 421 10792
rect 375 10720 421 10758
rect 375 10686 381 10720
rect 415 10686 421 10720
rect 375 10648 421 10686
rect 375 10614 381 10648
rect 415 10614 421 10648
rect 375 10576 421 10614
rect 375 10542 381 10576
rect 415 10542 421 10576
rect 375 10504 421 10542
rect 375 10470 381 10504
rect 415 10470 421 10504
rect 375 10432 421 10470
rect 375 10398 381 10432
rect 415 10398 421 10432
rect 375 10360 421 10398
rect 375 10326 381 10360
rect 415 10326 421 10360
rect 375 10288 421 10326
rect 375 10254 381 10288
rect 415 10254 421 10288
rect 375 10216 421 10254
rect 375 10182 381 10216
rect 415 10182 421 10216
rect 375 10144 421 10182
rect 375 10110 381 10144
rect 415 10110 421 10144
rect 375 10072 421 10110
rect 375 10038 381 10072
rect 415 10038 421 10072
rect 375 10000 421 10038
rect 375 9966 381 10000
rect 415 9966 421 10000
rect 375 9928 421 9966
rect 375 9894 381 9928
rect 415 9894 421 9928
rect 375 9856 421 9894
rect 375 9822 381 9856
rect 415 9822 421 9856
rect 375 9784 421 9822
rect 375 9750 381 9784
rect 415 9750 421 9784
rect 375 9712 421 9750
rect 375 9678 381 9712
rect 415 9678 421 9712
rect 375 9640 421 9678
rect 375 9606 381 9640
rect 415 9606 421 9640
rect 375 9568 421 9606
rect 375 9534 381 9568
rect 415 9534 421 9568
rect 375 9496 421 9534
rect 375 9462 381 9496
rect 415 9462 421 9496
rect 375 9424 421 9462
rect 375 9390 381 9424
rect 415 9390 421 9424
rect 375 9352 421 9390
rect 375 9318 381 9352
rect 415 9318 421 9352
rect 375 9280 421 9318
rect 375 9246 381 9280
rect 415 9246 421 9280
rect 375 9208 421 9246
rect 375 9174 381 9208
rect 415 9174 421 9208
rect 375 9136 421 9174
rect 375 9102 381 9136
rect 415 9102 421 9136
rect 375 9064 421 9102
rect 375 9030 381 9064
rect 415 9030 421 9064
rect 375 8992 421 9030
rect 375 8958 381 8992
rect 415 8958 421 8992
rect 375 8920 421 8958
rect 375 8886 381 8920
rect 415 8886 421 8920
rect 375 8848 421 8886
rect 375 8814 381 8848
rect 415 8814 421 8848
rect 375 8776 421 8814
rect 375 8742 381 8776
rect 415 8742 421 8776
rect 375 8704 421 8742
rect 375 8670 381 8704
rect 415 8670 421 8704
rect 375 8632 421 8670
rect 375 8598 381 8632
rect 415 8598 421 8632
rect 375 8560 421 8598
rect 375 8526 381 8560
rect 415 8526 421 8560
rect 375 8488 421 8526
rect 375 8454 381 8488
rect 415 8454 421 8488
rect 375 8416 421 8454
rect 375 8382 381 8416
rect 415 8382 421 8416
rect 375 8344 421 8382
rect 375 8310 381 8344
rect 415 8310 421 8344
rect 375 8272 421 8310
rect 375 8238 381 8272
rect 415 8238 421 8272
rect 375 8200 421 8238
rect 375 8166 381 8200
rect 415 8166 421 8200
rect 375 8128 421 8166
rect 375 8094 381 8128
rect 415 8094 421 8128
rect 375 8056 421 8094
rect 375 8022 381 8056
rect 415 8022 421 8056
rect 375 7984 421 8022
rect 375 7950 381 7984
rect 415 7950 421 7984
rect 375 7912 421 7950
rect 375 7878 381 7912
rect 415 7878 421 7912
rect 375 7840 421 7878
rect 375 7806 381 7840
rect 415 7806 421 7840
rect 375 7768 421 7806
rect 375 7734 381 7768
rect 415 7734 421 7768
rect 375 7696 421 7734
rect 375 7662 381 7696
rect 415 7662 421 7696
rect 375 7624 421 7662
rect 375 7590 381 7624
rect 415 7590 421 7624
rect 375 7552 421 7590
rect 375 7518 381 7552
rect 415 7518 421 7552
rect 375 7480 421 7518
rect 375 7446 381 7480
rect 415 7446 421 7480
rect 375 7408 421 7446
rect 375 7374 381 7408
rect 415 7374 421 7408
rect 375 7336 421 7374
rect 375 7302 381 7336
rect 415 7302 421 7336
rect 375 7264 421 7302
rect 375 7230 381 7264
rect 415 7230 421 7264
rect 375 7192 421 7230
rect 375 7158 381 7192
rect 415 7158 421 7192
rect 375 7120 421 7158
rect 375 7086 381 7120
rect 415 7086 421 7120
rect 375 7048 421 7086
rect 375 7014 381 7048
rect 415 7014 421 7048
rect 375 6976 421 7014
rect 375 6942 381 6976
rect 415 6942 421 6976
rect 375 6904 421 6942
rect 375 6870 381 6904
rect 415 6870 421 6904
rect 375 6832 421 6870
rect 375 6798 381 6832
rect 415 6798 421 6832
rect 375 6760 421 6798
rect 375 6726 381 6760
rect 415 6726 421 6760
rect 375 6688 421 6726
rect 375 6654 381 6688
rect 415 6654 421 6688
rect 375 6616 421 6654
rect 375 6582 381 6616
rect 415 6582 421 6616
rect 375 6544 421 6582
rect 375 6510 381 6544
rect 415 6510 421 6544
rect 375 6472 421 6510
rect 375 6438 381 6472
rect 415 6438 421 6472
rect 375 6400 421 6438
rect 375 6366 381 6400
rect 415 6366 421 6400
rect 375 6328 421 6366
rect 375 6294 381 6328
rect 415 6294 421 6328
rect 375 6256 421 6294
rect 375 6222 381 6256
rect 415 6222 421 6256
rect 375 6184 421 6222
rect 375 6150 381 6184
rect 415 6150 421 6184
rect 375 6112 421 6150
rect 375 6078 381 6112
rect 415 6078 421 6112
rect 375 6040 421 6078
rect 375 6006 381 6040
rect 415 6006 421 6040
rect 375 5968 421 6006
rect 375 5934 381 5968
rect 415 5934 421 5968
rect 375 5896 421 5934
rect 375 5862 381 5896
rect 415 5862 421 5896
rect 375 5824 421 5862
rect 375 5790 381 5824
rect 415 5790 421 5824
rect 375 5752 421 5790
rect 375 5718 381 5752
rect 415 5718 421 5752
rect 375 5680 421 5718
rect 375 5646 381 5680
rect 415 5646 421 5680
rect 375 5608 421 5646
rect 375 5574 381 5608
rect 415 5574 421 5608
rect 375 5536 421 5574
rect 375 5502 381 5536
rect 415 5502 421 5536
rect 375 5464 421 5502
rect 375 5430 381 5464
rect 415 5430 421 5464
rect 375 5392 421 5430
rect 375 5358 381 5392
rect 415 5358 421 5392
rect 375 5320 421 5358
rect 375 5286 381 5320
rect 415 5286 421 5320
rect 375 5248 421 5286
rect 375 5214 381 5248
rect 415 5214 421 5248
rect 375 5176 421 5214
rect 375 5142 381 5176
rect 415 5142 421 5176
rect 375 5104 421 5142
rect 375 5070 381 5104
rect 415 5070 421 5104
rect 375 5032 421 5070
rect 375 4998 381 5032
rect 415 4998 421 5032
rect 375 4960 421 4998
rect 375 4926 381 4960
rect 415 4926 421 4960
rect 375 4888 421 4926
rect 375 4854 381 4888
rect 415 4854 421 4888
rect 375 4816 421 4854
rect 375 4782 381 4816
rect 415 4782 421 4816
rect 375 4744 421 4782
rect 375 4710 381 4744
rect 415 4710 421 4744
rect 375 4672 421 4710
rect 375 4638 381 4672
rect 415 4638 421 4672
rect 375 4600 421 4638
rect 375 4566 381 4600
rect 415 4566 421 4600
rect 375 4528 421 4566
rect 375 4494 381 4528
rect 415 4494 421 4528
rect 375 4456 421 4494
rect 375 4422 381 4456
rect 415 4422 421 4456
rect 375 4384 421 4422
rect 375 4350 381 4384
rect 415 4350 421 4384
rect 375 4312 421 4350
rect 375 4278 381 4312
rect 415 4278 421 4312
rect 375 4240 421 4278
rect 375 4206 381 4240
rect 415 4206 421 4240
rect 375 4168 421 4206
rect 3015 10350 3061 10362
rect 3015 10316 3021 10350
rect 3055 10316 3061 10350
rect 3015 10278 3061 10316
rect 3015 10244 3021 10278
rect 3055 10244 3061 10278
rect 3015 10206 3061 10244
rect 3015 10172 3021 10206
rect 3055 10172 3061 10206
rect 3015 10134 3061 10172
rect 3015 10100 3021 10134
rect 3055 10100 3061 10134
rect 3015 10062 3061 10100
rect 3015 10028 3021 10062
rect 3055 10028 3061 10062
rect 3015 9990 3061 10028
rect 3015 9956 3021 9990
rect 3055 9956 3061 9990
rect 3015 9918 3061 9956
rect 3015 9884 3021 9918
rect 3055 9884 3061 9918
rect 3015 9846 3061 9884
rect 3015 9812 3021 9846
rect 3055 9812 3061 9846
rect 3015 9774 3061 9812
rect 3015 9740 3021 9774
rect 3055 9740 3061 9774
rect 3015 9702 3061 9740
rect 3015 9668 3021 9702
rect 3055 9668 3061 9702
rect 3015 9630 3061 9668
rect 3015 9596 3021 9630
rect 3055 9596 3061 9630
rect 3015 9558 3061 9596
rect 3015 9524 3021 9558
rect 3055 9524 3061 9558
rect 3015 9486 3061 9524
rect 3015 9452 3021 9486
rect 3055 9452 3061 9486
rect 3015 9414 3061 9452
rect 3015 9380 3021 9414
rect 3055 9380 3061 9414
rect 3015 9342 3061 9380
rect 3015 9308 3021 9342
rect 3055 9308 3061 9342
rect 3015 9270 3061 9308
rect 3015 9236 3021 9270
rect 3055 9236 3061 9270
rect 3015 9198 3061 9236
rect 3015 9164 3021 9198
rect 3055 9164 3061 9198
rect 3015 9126 3061 9164
rect 3015 9092 3021 9126
rect 3055 9092 3061 9126
rect 3015 9054 3061 9092
rect 3015 9020 3021 9054
rect 3055 9020 3061 9054
rect 3015 8982 3061 9020
rect 3015 8948 3021 8982
rect 3055 8948 3061 8982
rect 3015 8910 3061 8948
rect 3015 8876 3021 8910
rect 3055 8876 3061 8910
rect 3015 8838 3061 8876
rect 3015 8804 3021 8838
rect 3055 8804 3061 8838
rect 3015 8766 3061 8804
rect 3015 8732 3021 8766
rect 3055 8732 3061 8766
rect 3015 8694 3061 8732
rect 3015 8660 3021 8694
rect 3055 8660 3061 8694
rect 3015 8622 3061 8660
rect 3015 8588 3021 8622
rect 3055 8588 3061 8622
rect 3015 8550 3061 8588
rect 3015 8516 3021 8550
rect 3055 8516 3061 8550
rect 3015 8478 3061 8516
rect 3015 8444 3021 8478
rect 3055 8444 3061 8478
rect 3015 8406 3061 8444
rect 3015 8372 3021 8406
rect 3055 8372 3061 8406
rect 3015 8334 3061 8372
rect 3015 8300 3021 8334
rect 3055 8300 3061 8334
rect 3015 8262 3061 8300
rect 3015 8228 3021 8262
rect 3055 8228 3061 8262
rect 3015 8190 3061 8228
rect 3015 8156 3021 8190
rect 3055 8156 3061 8190
rect 3015 8118 3061 8156
rect 3015 8084 3021 8118
rect 3055 8084 3061 8118
rect 3015 8046 3061 8084
rect 3015 8012 3021 8046
rect 3055 8012 3061 8046
rect 3015 7974 3061 8012
rect 3015 7940 3021 7974
rect 3055 7940 3061 7974
rect 3015 7902 3061 7940
rect 3015 7868 3021 7902
rect 3055 7868 3061 7902
rect 3015 7830 3061 7868
rect 3015 7796 3021 7830
rect 3055 7796 3061 7830
rect 3015 7758 3061 7796
rect 3015 7724 3021 7758
rect 3055 7724 3061 7758
rect 3015 7686 3061 7724
rect 3015 7652 3021 7686
rect 3055 7652 3061 7686
rect 3015 7614 3061 7652
rect 3015 7580 3021 7614
rect 3055 7580 3061 7614
rect 3015 7542 3061 7580
rect 3015 7508 3021 7542
rect 3055 7508 3061 7542
rect 3015 7470 3061 7508
rect 3015 7436 3021 7470
rect 3055 7436 3061 7470
rect 3015 7398 3061 7436
rect 3015 7364 3021 7398
rect 3055 7364 3061 7398
rect 3015 7326 3061 7364
rect 3015 7292 3021 7326
rect 3055 7292 3061 7326
rect 3015 7254 3061 7292
rect 3015 7220 3021 7254
rect 3055 7220 3061 7254
rect 3015 7182 3061 7220
rect 3015 7148 3021 7182
rect 3055 7148 3061 7182
rect 3015 7110 3061 7148
rect 3015 7076 3021 7110
rect 3055 7076 3061 7110
rect 3015 7038 3061 7076
rect 3015 7004 3021 7038
rect 3055 7004 3061 7038
rect 3015 6966 3061 7004
rect 3015 6932 3021 6966
rect 3055 6932 3061 6966
rect 3015 6894 3061 6932
rect 3015 6860 3021 6894
rect 3055 6860 3061 6894
rect 3015 6822 3061 6860
rect 3015 6788 3021 6822
rect 3055 6788 3061 6822
rect 3015 6750 3061 6788
rect 3015 6716 3021 6750
rect 3055 6716 3061 6750
rect 3015 6678 3061 6716
rect 3015 6644 3021 6678
rect 3055 6644 3061 6678
rect 3015 6606 3061 6644
rect 3015 6572 3021 6606
rect 3055 6572 3061 6606
rect 3015 6534 3061 6572
rect 3015 6500 3021 6534
rect 3055 6500 3061 6534
rect 3015 6462 3061 6500
rect 3015 6428 3021 6462
rect 3055 6428 3061 6462
rect 3015 6390 3061 6428
rect 3015 6356 3021 6390
rect 3055 6356 3061 6390
rect 3015 6318 3061 6356
rect 3015 6284 3021 6318
rect 3055 6284 3061 6318
rect 3015 6246 3061 6284
rect 3015 6212 3021 6246
rect 3055 6212 3061 6246
rect 3015 6174 3061 6212
rect 3015 6140 3021 6174
rect 3055 6140 3061 6174
rect 3015 6102 3061 6140
rect 3015 6068 3021 6102
rect 3055 6068 3061 6102
rect 3015 6030 3061 6068
rect 3015 5996 3021 6030
rect 3055 5996 3061 6030
rect 3015 5958 3061 5996
rect 3015 5924 3021 5958
rect 3055 5924 3061 5958
rect 3015 5886 3061 5924
rect 3015 5852 3021 5886
rect 3055 5852 3061 5886
rect 3015 5814 3061 5852
rect 3015 5780 3021 5814
rect 3055 5780 3061 5814
rect 3015 5742 3061 5780
rect 3015 5708 3021 5742
rect 3055 5708 3061 5742
rect 3015 5670 3061 5708
rect 3015 5636 3021 5670
rect 3055 5636 3061 5670
rect 3015 5598 3061 5636
rect 3015 5564 3021 5598
rect 3055 5564 3061 5598
rect 3015 5526 3061 5564
rect 3015 5492 3021 5526
rect 3055 5492 3061 5526
rect 3015 5454 3061 5492
rect 3015 5420 3021 5454
rect 3055 5420 3061 5454
rect 3015 5382 3061 5420
rect 3015 5348 3021 5382
rect 3055 5348 3061 5382
rect 3015 5309 3061 5348
rect 3015 5275 3021 5309
rect 3055 5275 3061 5309
rect 3015 5236 3061 5275
rect 3015 5202 3021 5236
rect 3055 5202 3061 5236
rect 3015 5163 3061 5202
rect 3015 5129 3021 5163
rect 3055 5129 3061 5163
rect 3015 5090 3061 5129
rect 3015 5056 3021 5090
rect 3055 5056 3061 5090
rect 3015 5017 3061 5056
rect 3015 4983 3021 5017
rect 3055 4983 3061 5017
rect 3015 4944 3061 4983
rect 3015 4910 3021 4944
rect 3055 4910 3061 4944
rect 3015 4871 3061 4910
rect 3015 4837 3021 4871
rect 3055 4837 3061 4871
rect 3015 4798 3061 4837
rect 3015 4764 3021 4798
rect 3055 4764 3061 4798
rect 3015 4725 3061 4764
rect 3015 4691 3021 4725
rect 3055 4691 3061 4725
rect 3015 4652 3061 4691
rect 3015 4618 3021 4652
rect 3055 4618 3061 4652
rect 3015 4579 3061 4618
rect 3015 4545 3021 4579
rect 3055 4545 3061 4579
rect 3015 4506 3061 4545
rect 3015 4472 3021 4506
rect 3055 4472 3061 4506
rect 3015 4433 3061 4472
rect 3015 4399 3021 4433
rect 3055 4399 3061 4433
rect 3015 4360 3061 4399
rect 3015 4326 3021 4360
rect 3055 4326 3061 4360
rect 3015 4287 3061 4326
rect 3015 4253 3021 4287
rect 3055 4253 3061 4287
rect 3015 4214 3061 4253
rect 3015 4180 3021 4214
rect 3055 4180 3061 4214
rect 3015 4168 3061 4180
rect 375 4134 381 4168
rect 415 4134 421 4168
rect 375 4095 421 4134
rect 375 4061 381 4095
rect 415 4061 421 4095
rect 375 4022 421 4061
rect 375 3988 381 4022
rect 415 3988 421 4022
rect 375 3949 421 3988
rect 375 3915 381 3949
rect 415 3915 421 3949
rect 375 3876 421 3915
rect 375 3842 381 3876
rect 415 3842 421 3876
rect 375 3803 421 3842
rect 375 3769 381 3803
rect 415 3769 421 3803
rect 375 3730 421 3769
rect 375 3696 381 3730
rect 415 3696 421 3730
rect 375 3657 421 3696
rect 375 3623 381 3657
rect 415 3623 421 3657
rect 375 3584 421 3623
rect 375 3550 381 3584
rect 415 3550 421 3584
rect 375 3511 421 3550
rect 375 3477 381 3511
rect 415 3477 421 3511
rect 375 3438 421 3477
rect 375 3404 381 3438
rect 415 3404 421 3438
rect 375 3365 421 3404
rect 375 3331 381 3365
rect 415 3331 421 3365
rect 375 3292 421 3331
rect 375 3258 381 3292
rect 415 3258 421 3292
rect 375 3219 421 3258
rect 375 3185 381 3219
rect 415 3185 421 3219
rect 375 3146 421 3185
rect 375 3112 381 3146
rect 415 3112 421 3146
rect 375 3073 421 3112
rect 375 3039 381 3073
rect 415 3039 421 3073
rect 375 3000 421 3039
rect 375 2966 381 3000
rect 415 2966 421 3000
rect 375 2927 421 2966
rect 375 2893 381 2927
rect 415 2893 421 2927
rect 375 2854 421 2893
rect 375 2820 381 2854
rect 415 2820 421 2854
rect 375 2781 421 2820
rect 375 2747 381 2781
rect 415 2747 421 2781
rect 375 2708 421 2747
rect 375 2674 381 2708
rect 415 2674 421 2708
rect 375 2635 421 2674
rect 375 2601 381 2635
rect 415 2601 421 2635
rect 375 2562 421 2601
rect 375 2528 381 2562
rect 415 2528 421 2562
rect 375 2489 421 2528
rect 375 2455 381 2489
rect 415 2455 421 2489
rect 375 2416 421 2455
rect 375 2382 381 2416
rect 415 2382 421 2416
rect 375 2343 421 2382
rect 375 2309 381 2343
rect 415 2309 421 2343
rect 375 2270 421 2309
rect 375 2236 381 2270
rect 415 2236 421 2270
rect 375 2197 421 2236
rect 375 2163 381 2197
rect 415 2163 421 2197
rect 375 2124 421 2163
rect 375 2090 381 2124
rect 415 2090 421 2124
rect 375 2051 421 2090
rect 375 2017 381 2051
rect 415 2017 421 2051
rect 375 1978 421 2017
rect 375 1944 381 1978
rect 415 1944 421 1978
rect 375 1905 421 1944
rect 375 1871 381 1905
rect 415 1871 421 1905
rect 375 1832 421 1871
rect 375 1798 381 1832
rect 415 1798 421 1832
rect 375 1759 421 1798
rect 375 1725 381 1759
rect 415 1725 421 1759
rect 375 1686 421 1725
rect 375 1652 381 1686
rect 415 1652 421 1686
rect 375 1613 421 1652
rect 375 1579 381 1613
rect 415 1579 421 1613
rect 375 1540 421 1579
rect 375 1506 381 1540
rect 415 1506 421 1540
rect 375 1467 421 1506
rect 375 1433 381 1467
rect 415 1433 421 1467
rect 375 1394 421 1433
rect 375 1360 381 1394
rect 415 1360 421 1394
rect 375 1321 421 1360
rect 375 1287 381 1321
rect 415 1287 421 1321
rect 375 1248 421 1287
rect 375 1214 381 1248
rect 415 1214 421 1248
rect 375 1175 421 1214
rect 375 1141 381 1175
rect 415 1141 421 1175
rect 375 1102 421 1141
rect 375 1068 381 1102
rect 415 1068 421 1102
rect 375 1029 421 1068
rect 375 995 381 1029
rect 415 995 421 1029
rect 375 956 421 995
rect 375 922 381 956
rect 415 922 421 956
rect 375 910 421 922
rect 1695 3642 1741 3674
rect 1695 3608 1701 3642
rect 1735 3608 1741 3642
rect 1695 3570 1741 3608
rect 1695 3536 1701 3570
rect 1735 3536 1741 3570
rect 1695 3498 1741 3536
rect 1695 3464 1701 3498
rect 1735 3464 1741 3498
rect 1695 3426 1741 3464
rect 1695 3392 1701 3426
rect 1735 3392 1741 3426
rect 1695 3354 1741 3392
rect 1695 3320 1701 3354
rect 1735 3320 1741 3354
rect 1695 3282 1741 3320
rect 1695 3248 1701 3282
rect 1735 3248 1741 3282
rect 1695 3210 1741 3248
rect 1695 3176 1701 3210
rect 1735 3176 1741 3210
rect 1695 3138 1741 3176
rect 1695 3104 1701 3138
rect 1735 3104 1741 3138
rect 1695 3066 1741 3104
rect 1695 3032 1701 3066
rect 1735 3032 1741 3066
rect 1695 2994 1741 3032
rect 1695 2960 1701 2994
rect 1735 2960 1741 2994
rect 1695 2922 1741 2960
rect 1695 2888 1701 2922
rect 1735 2888 1741 2922
rect 1695 2850 1741 2888
rect 1695 2816 1701 2850
rect 1735 2816 1741 2850
rect 1695 2778 1741 2816
rect 1695 2744 1701 2778
rect 1735 2744 1741 2778
rect 1695 2706 1741 2744
rect 1695 2672 1701 2706
rect 1735 2672 1741 2706
rect 1695 2634 1741 2672
rect 1695 2600 1701 2634
rect 1735 2600 1741 2634
rect 1695 2562 1741 2600
tri 2781 2576 2855 2650 se
rect 2855 2636 3898 2650
tri 3898 2636 3912 2650 sw
rect 2855 2598 3912 2636
tri 2855 2576 2877 2598 nw
tri 3876 2576 3898 2598 ne
rect 3898 2576 3912 2598
rect 1695 2528 1701 2562
rect 1735 2528 1741 2562
rect 1695 2490 1741 2528
rect 1695 2456 1701 2490
rect 1735 2456 1741 2490
rect 1695 2418 1741 2456
rect 1695 2384 1701 2418
rect 1735 2384 1741 2418
rect 1695 2346 1741 2384
tri 2739 2534 2781 2576 se
rect 2781 2534 2791 2576
rect 2739 2475 2791 2534
tri 2791 2512 2855 2576 nw
tri 3898 2562 3912 2576 ne
tri 3912 2562 3986 2636 sw
tri 3912 2534 3940 2562 ne
rect 2739 2411 2791 2423
rect 2739 2353 2791 2359
rect 1695 2312 1701 2346
rect 1735 2312 1741 2346
rect 1695 2274 1741 2312
rect 1695 2240 1701 2274
rect 1735 2240 1741 2274
rect 1695 2202 1741 2240
rect 1695 2168 1701 2202
rect 1735 2168 1741 2202
rect 1695 2130 1741 2168
rect 1695 2096 1701 2130
rect 1735 2096 1741 2130
rect 1695 2058 1741 2096
rect 1695 2024 1701 2058
rect 1735 2024 1741 2058
rect 3189 2336 3195 2388
rect 3247 2336 3259 2388
rect 3311 2336 3323 2388
rect 3375 2379 3414 2388
rect 3379 2345 3414 2379
rect 3375 2336 3414 2345
rect 3189 2305 3241 2336
rect 3189 2293 3198 2305
rect 3232 2293 3241 2305
rect 3189 2233 3241 2241
rect 3189 2229 3198 2233
rect 3232 2229 3241 2233
rect 3189 2165 3241 2177
rect 3189 2101 3241 2113
rect 3189 2043 3241 2049
rect 3338 2260 3684 2266
rect 3338 2226 3350 2260
rect 3384 2226 3422 2260
rect 3456 2226 3494 2260
rect 3528 2226 3566 2260
rect 3600 2226 3638 2260
rect 3672 2226 3684 2260
rect 3338 2220 3684 2226
rect 3940 2231 3986 2562
rect 3338 2197 3546 2220
tri 3546 2197 3569 2220 nw
rect 3940 2197 3946 2231
rect 3980 2197 3986 2231
rect 1695 1986 1741 2024
tri 3313 1989 3338 2014 se
rect 3338 1989 3544 2197
tri 3544 2195 3546 2197 nw
rect 3940 2159 3986 2197
rect 3940 2125 3946 2159
rect 3980 2125 3986 2159
rect 3940 2113 3986 2125
rect 3615 2104 3889 2110
rect 3615 2070 3627 2104
rect 3661 2070 3699 2104
rect 3733 2070 3771 2104
rect 3805 2070 3843 2104
rect 3877 2070 3889 2104
rect 3615 2064 3889 2070
tri 3687 2039 3712 2064 ne
rect 1695 1952 1701 1986
rect 1735 1952 1741 1986
rect 1695 1914 1741 1952
rect 1695 1880 1701 1914
rect 1735 1880 1741 1914
rect 1695 1842 1741 1880
rect 1695 1808 1701 1842
rect 1735 1808 1741 1842
rect 1695 1770 1741 1808
rect 1848 1983 3544 1989
rect 1848 1931 1865 1983
rect 1917 1931 2204 1983
rect 2256 1931 2328 1983
rect 2380 1931 2564 1983
rect 2616 1931 2638 1983
rect 2690 1931 2712 1983
rect 2764 1954 3544 1983
rect 3712 2015 3889 2064
tri 3889 2015 3918 2044 sw
tri 3544 1954 3569 1979 sw
rect 2764 1948 3684 1954
rect 2764 1931 3350 1948
rect 1848 1917 3350 1931
rect 1848 1865 1865 1917
rect 1917 1865 2204 1917
rect 2256 1865 2328 1917
rect 2380 1865 2564 1917
rect 2616 1865 2638 1917
rect 2690 1865 2712 1917
rect 2764 1914 3350 1917
rect 3384 1914 3422 1948
rect 3456 1914 3494 1948
rect 3528 1914 3566 1948
rect 3600 1914 3638 1948
rect 3672 1914 3684 1948
rect 2764 1908 3684 1914
rect 2764 1865 3544 1908
tri 3544 1883 3569 1908 nw
rect 1848 1850 3544 1865
rect 1848 1798 1865 1850
rect 1917 1798 2204 1850
rect 2256 1798 2328 1850
rect 2380 1798 2564 1850
rect 2616 1798 2638 1850
rect 2690 1798 2712 1850
rect 2764 1798 3544 1850
tri 3687 1798 3712 1823 se
rect 3712 1798 3918 2015
rect 1848 1792 3544 1798
rect 1695 1736 1701 1770
rect 1735 1736 1741 1770
tri 3313 1767 3338 1792 ne
rect 1695 1698 1741 1736
rect 1695 1664 1701 1698
rect 1735 1664 1741 1698
rect 1695 1626 1741 1664
rect 1695 1592 1701 1626
rect 1735 1592 1741 1626
rect 1695 1554 1741 1592
rect 1695 1520 1701 1554
rect 1735 1520 1741 1554
rect 1695 1482 1741 1520
rect 1695 1448 1701 1482
rect 1735 1448 1741 1482
rect 1695 1410 1741 1448
rect 1695 1376 1701 1410
rect 1735 1376 1741 1410
rect 1695 1338 1741 1376
rect 1695 1304 1701 1338
rect 1735 1304 1741 1338
rect 1695 1266 1741 1304
rect 1695 1232 1701 1266
rect 1735 1232 1741 1266
rect 1695 1194 1741 1232
rect 1695 1160 1701 1194
rect 1735 1160 1741 1194
rect 1695 1122 1741 1160
rect 1695 1088 1701 1122
rect 1735 1088 1741 1122
rect 1695 1050 1741 1088
rect 1695 1016 1701 1050
rect 1735 1016 1741 1050
rect 1695 978 1741 1016
rect 3189 1724 3241 1730
rect 3189 1660 3241 1672
rect 3189 1596 3241 1608
rect 3189 1540 3198 1544
rect 3232 1540 3241 1544
rect 3189 1532 3241 1540
rect 3189 1468 3198 1480
rect 3232 1468 3241 1480
rect 3189 1404 3198 1416
rect 3232 1404 3241 1416
rect 3189 1340 3198 1352
rect 3232 1340 3241 1352
rect 3189 1286 3241 1288
rect 3189 1276 3198 1286
rect 3232 1276 3241 1286
rect 3338 1642 3544 1792
rect 3572 1792 3918 1798
rect 3572 1758 3584 1792
rect 3618 1758 3656 1792
rect 3690 1758 3728 1792
rect 3762 1758 3800 1792
rect 3834 1758 3872 1792
rect 3906 1758 3918 1792
rect 3572 1752 3918 1758
tri 3687 1727 3712 1752 ne
tri 3544 1642 3569 1667 sw
rect 3338 1636 3684 1642
rect 3338 1602 3350 1636
rect 3384 1602 3422 1636
rect 3456 1602 3494 1636
rect 3528 1602 3566 1636
rect 3600 1602 3638 1636
rect 3672 1602 3684 1636
rect 3338 1596 3684 1602
rect 3338 1330 3544 1596
tri 3544 1571 3569 1596 nw
tri 3687 1486 3712 1511 se
rect 3712 1486 3918 1752
rect 3572 1480 3918 1486
rect 3572 1446 3584 1480
rect 3618 1446 3656 1480
rect 3690 1446 3728 1480
rect 3762 1446 3800 1480
rect 3834 1446 3872 1480
rect 3906 1446 3918 1480
rect 3572 1440 3918 1446
tri 3687 1415 3712 1440 ne
tri 3544 1330 3569 1355 sw
rect 3338 1324 3684 1330
rect 3338 1290 3350 1324
rect 3384 1290 3422 1324
rect 3456 1290 3494 1324
rect 3528 1290 3566 1324
rect 3600 1290 3638 1324
rect 3672 1290 3684 1324
rect 3338 1284 3684 1290
rect 3189 1214 3241 1224
rect 3189 1212 3198 1214
rect 3232 1212 3241 1214
tri 3687 1194 3712 1219 se
rect 3712 1194 3918 1440
rect 3189 1148 3241 1160
rect 3572 1188 3918 1194
rect 3572 1154 3584 1188
rect 3618 1154 3656 1188
rect 3690 1154 3728 1188
rect 3762 1154 3800 1188
rect 3834 1154 3872 1188
rect 3906 1154 3918 1188
rect 3572 1148 3918 1154
tri 3687 1123 3712 1148 ne
rect 3189 1059 3241 1096
rect 3189 1007 3195 1059
rect 3247 1007 3259 1059
rect 3311 1007 3323 1059
rect 3375 1050 3414 1059
rect 3379 1016 3414 1050
rect 3375 1007 3414 1016
tri 3674 1007 3712 1045 se
rect 3712 1007 3918 1148
tri 3645 978 3674 1007 se
rect 3674 978 3918 1007
rect 1695 944 1701 978
rect 1735 944 1741 978
rect 1695 906 1741 944
rect 1695 872 1701 906
rect 1735 872 1741 906
rect 1695 834 1741 872
rect 304 824 833 830
rect 356 802 833 824
tri 833 802 861 830 sw
rect 356 800 861 802
tri 861 800 863 802 sw
rect 1695 800 1701 834
rect 1735 800 1741 834
rect 356 772 863 800
rect 304 762 863 772
tri 863 762 901 800 sw
rect 1695 762 1741 800
tri 2855 799 3034 978 se
rect 3034 966 3918 978
rect 3034 848 3800 966
tri 3800 848 3918 966 nw
rect 3034 799 3039 848
tri 3039 799 3088 848 nw
rect 304 758 901 762
rect 356 728 901 758
tri 901 728 935 762 sw
rect 1695 728 1701 762
rect 1735 728 1741 762
rect 356 706 935 728
rect 304 700 935 706
tri 779 690 789 700 ne
rect 789 690 935 700
tri 935 690 973 728 sw
rect 1695 690 1741 728
tri 789 656 823 690 ne
rect 823 656 973 690
tri 973 656 1007 690 sw
rect 1695 656 1701 690
rect 1735 656 1741 690
tri 823 630 849 656 ne
rect 849 630 1007 656
rect 375 618 421 630
tri 849 618 861 630 ne
rect 861 618 1007 630
tri 1007 618 1045 656 sw
rect 375 584 381 618
rect 415 584 421 618
tri 861 617 862 618 ne
rect 862 617 1045 618
rect 375 530 421 584
tri 862 583 896 617 ne
rect 896 583 1045 617
tri 896 578 901 583 ne
rect 901 578 1045 583
rect 552 572 656 578
tri 537 553 552 568 se
rect 552 553 578 572
tri 528 544 537 553 se
rect 537 544 578 553
rect 375 496 381 530
rect 415 496 421 530
tri 494 510 528 544 se
rect 528 520 578 544
rect 630 520 656 572
tri 901 564 915 578 ne
rect 528 510 656 520
rect 375 442 421 496
tri 461 477 494 510 se
rect 494 506 656 510
rect 494 477 578 506
tri 455 471 461 477 se
rect 461 471 578 477
rect 375 408 381 442
rect 415 408 421 442
rect 375 353 421 408
rect 375 319 381 353
rect 415 319 421 353
tri 451 467 455 471 se
rect 455 467 578 471
rect 451 454 578 467
rect 630 454 656 506
rect 451 448 656 454
rect 451 437 605 448
tri 605 437 616 448 nw
rect 451 436 604 437
tri 604 436 605 437 nw
rect 915 436 1045 578
rect 1695 617 1741 656
rect 1990 761 2327 769
rect 2042 759 2327 761
tri 2327 759 2337 769 sw
rect 2042 709 2337 759
rect 1990 697 2337 709
rect 2042 645 2337 697
rect 1990 639 2337 645
rect 1695 583 1701 617
rect 1735 583 1741 617
tri 2273 587 2325 639 ne
rect 2325 587 2337 639
tri 2337 587 2509 759 sw
rect 1695 544 1741 583
tri 2325 575 2337 587 ne
rect 2337 575 2509 587
tri 2509 575 2521 587 sw
tri 2337 553 2359 575 ne
rect 2359 553 2521 575
rect 1695 510 1701 544
rect 1735 510 1741 544
tri 2359 521 2391 553 ne
rect 1695 471 1741 510
rect 1695 437 1701 471
rect 1735 437 1741 471
rect 451 352 581 436
tri 581 413 604 436 nw
rect 1695 398 1741 437
rect 2391 436 2521 553
rect 1695 364 1701 398
rect 1735 364 1741 398
rect 375 259 421 319
tri 421 259 443 281 sw
tri 39 216 41 218 sw
rect -7 211 41 216
tri 41 211 46 216 sw
rect -7 198 46 211
tri 46 198 59 211 sw
rect 228 207 234 259
rect 286 207 298 259
rect 350 207 362 259
rect 414 250 426 259
rect 478 256 496 259
tri 496 256 499 259 sw
tri 873 256 876 259 se
rect 876 256 882 259
rect 478 250 882 256
rect 934 250 946 259
rect 998 250 1010 259
rect 1062 250 1074 259
rect 1126 256 1144 259
tri 1144 256 1147 259 sw
tri 1197 256 1200 259 se
rect 1200 256 1206 259
rect 1126 250 1206 256
rect 1258 250 1270 259
rect 500 216 539 250
rect 573 216 612 250
rect 646 216 685 250
rect 719 216 758 250
rect 792 216 831 250
rect 865 216 882 250
rect 938 216 946 250
rect 1157 216 1196 250
rect 1258 216 1269 250
rect 414 207 426 216
rect 478 210 882 216
rect 478 207 496 210
tri 496 207 499 210 nw
tri 873 207 876 210 ne
rect 876 207 882 210
rect 934 207 946 216
rect 998 207 1010 216
rect 1062 207 1074 216
rect 1126 210 1206 216
rect 1126 207 1144 210
tri 1144 207 1147 210 nw
tri 1197 207 1200 210 ne
rect 1200 207 1206 210
rect 1258 207 1270 216
rect 1322 207 1334 259
rect 1386 207 1398 259
rect 1450 256 1468 259
tri 1468 256 1471 259 sw
rect 1695 256 1741 364
rect 2855 352 2985 799
tri 2985 745 3039 799 nw
rect 3564 593 3616 599
rect 3564 520 3616 541
rect 3564 447 3616 468
rect 3564 374 3616 395
rect 3564 301 3616 322
tri 1845 256 1848 259 se
rect 1848 256 1854 259
rect 1450 250 1854 256
rect 1450 216 1488 250
rect 1522 216 1561 250
rect 1595 216 1634 250
rect 1668 216 1707 250
rect 1741 216 1780 250
rect 1814 216 1853 250
rect 1450 210 1854 216
rect 1450 207 1468 210
tri 1468 207 1471 210 nw
tri 1845 207 1848 210 ne
rect 1848 207 1854 210
rect 1906 207 1918 259
rect 1970 207 1982 259
rect 2034 256 2081 259
tri 2081 256 2084 259 sw
tri 2201 256 2204 259 se
rect 2204 256 2210 259
rect 2034 250 2210 256
rect 2034 216 2072 250
rect 2106 216 2145 250
rect 2179 216 2210 250
rect 2034 210 2210 216
rect 2034 207 2081 210
tri 2081 207 2084 210 nw
tri 2201 207 2204 210 ne
rect 2204 207 2210 210
rect 2262 207 2274 259
rect 2326 256 2380 259
tri 2380 256 2383 259 sw
tri 2561 256 2564 259 se
rect 2564 256 2570 259
rect 2326 250 2570 256
rect 2326 216 2361 250
rect 2395 216 2433 250
rect 2467 216 2505 250
rect 2539 216 2570 250
rect 2326 210 2570 216
rect 2326 207 2380 210
tri 2380 207 2383 210 nw
tri 2561 207 2564 210 ne
rect 2564 207 2570 210
rect 2622 207 2634 259
rect 2686 207 2698 259
rect 2750 256 2764 259
tri 2764 256 2767 259 sw
rect 2750 250 3055 256
rect 2755 216 2793 250
rect 2827 216 2865 250
rect 2899 216 2937 250
rect 2971 216 3009 250
rect 3043 216 3055 250
rect 2750 210 3055 216
rect 3564 228 3616 249
rect 2750 207 2764 210
tri 2764 207 2767 210 nw
tri -7 177 14 198 ne
rect 14 177 59 198
tri 59 177 80 198 sw
tri 14 136 55 177 ne
rect 55 155 80 177
tri 80 155 102 177 sw
rect 2408 155 2414 161
rect 55 136 2414 155
tri 55 132 59 136 ne
rect 59 132 2414 136
tri 59 109 82 132 ne
rect 82 109 2414 132
rect 2466 109 2478 161
rect 2530 109 2536 161
rect 3564 156 3616 176
tri -377 67 -352 92 se
rect -352 67 -306 107
rect 3564 102 3576 104
rect 3610 102 3616 104
tri 3563 92 3564 93 se
rect 3564 92 3616 102
tri -306 67 -281 92 sw
tri 3538 67 3563 92 se
rect 3563 84 3616 92
rect 3563 67 3564 84
rect -1262 32 3564 67
rect -1262 27 3576 32
rect 3610 27 3616 32
rect -1262 0 3616 27
<< via1 >>
rect 2124 17544 2176 17596
rect 2124 17480 2176 17532
rect 304 12266 356 12318
rect 304 12202 356 12254
rect 1990 12162 2042 12214
rect 1990 12098 2042 12150
rect -824 2531 -772 2583
rect -824 2467 -772 2519
rect 2739 2423 2791 2475
rect 2739 2359 2791 2411
rect 3195 2379 3247 2388
rect 3195 2345 3201 2379
rect 3201 2345 3235 2379
rect 3235 2345 3247 2379
rect 3195 2336 3247 2345
rect 3259 2379 3311 2388
rect 3259 2345 3273 2379
rect 3273 2345 3307 2379
rect 3307 2345 3311 2379
rect 3259 2336 3311 2345
rect 3323 2379 3375 2388
rect 3323 2345 3345 2379
rect 3345 2345 3375 2379
rect 3323 2336 3375 2345
rect 3189 2271 3198 2293
rect 3198 2271 3232 2293
rect 3232 2271 3241 2293
rect 3189 2241 3241 2271
rect 3189 2199 3198 2229
rect 3198 2199 3232 2229
rect 3232 2199 3241 2229
rect 3189 2177 3241 2199
rect 3189 2161 3241 2165
rect 3189 2127 3198 2161
rect 3198 2127 3232 2161
rect 3232 2127 3241 2161
rect 3189 2113 3241 2127
rect 3189 2089 3241 2101
rect 3189 2055 3198 2089
rect 3198 2055 3232 2089
rect 3232 2055 3241 2089
rect 3189 2049 3241 2055
rect 1865 1931 1917 1983
rect 2204 1931 2256 1983
rect 2328 1931 2380 1983
rect 2564 1931 2616 1983
rect 2638 1931 2690 1983
rect 2712 1931 2764 1983
rect 1865 1865 1917 1917
rect 2204 1865 2256 1917
rect 2328 1865 2380 1917
rect 2564 1865 2616 1917
rect 2638 1865 2690 1917
rect 2712 1865 2764 1917
rect 1865 1798 1917 1850
rect 2204 1798 2256 1850
rect 2328 1798 2380 1850
rect 2564 1798 2616 1850
rect 2638 1798 2690 1850
rect 2712 1798 2764 1850
rect 3189 1718 3241 1724
rect 3189 1684 3198 1718
rect 3198 1684 3232 1718
rect 3232 1684 3241 1718
rect 3189 1672 3241 1684
rect 3189 1646 3241 1660
rect 3189 1612 3198 1646
rect 3198 1612 3232 1646
rect 3232 1612 3241 1646
rect 3189 1608 3241 1612
rect 3189 1574 3241 1596
rect 3189 1544 3198 1574
rect 3198 1544 3232 1574
rect 3232 1544 3241 1574
rect 3189 1502 3241 1532
rect 3189 1480 3198 1502
rect 3198 1480 3232 1502
rect 3232 1480 3241 1502
rect 3189 1430 3241 1468
rect 3189 1416 3198 1430
rect 3198 1416 3232 1430
rect 3232 1416 3241 1430
rect 3189 1396 3198 1404
rect 3198 1396 3232 1404
rect 3232 1396 3241 1404
rect 3189 1358 3241 1396
rect 3189 1352 3198 1358
rect 3198 1352 3232 1358
rect 3232 1352 3241 1358
rect 3189 1324 3198 1340
rect 3198 1324 3232 1340
rect 3232 1324 3241 1340
rect 3189 1288 3241 1324
rect 3189 1252 3198 1276
rect 3198 1252 3232 1276
rect 3232 1252 3241 1276
rect 3189 1224 3241 1252
rect 3189 1180 3198 1212
rect 3198 1180 3232 1212
rect 3232 1180 3241 1212
rect 3189 1160 3241 1180
rect 3189 1142 3241 1148
rect 3189 1108 3198 1142
rect 3198 1108 3232 1142
rect 3232 1108 3241 1142
rect 3189 1096 3241 1108
rect 3195 1050 3247 1059
rect 3195 1016 3201 1050
rect 3201 1016 3235 1050
rect 3235 1016 3247 1050
rect 3195 1007 3247 1016
rect 3259 1050 3311 1059
rect 3259 1016 3273 1050
rect 3273 1016 3307 1050
rect 3307 1016 3311 1050
rect 3259 1007 3311 1016
rect 3323 1050 3375 1059
rect 3323 1016 3345 1050
rect 3345 1016 3375 1050
rect 3323 1007 3375 1016
rect 304 772 356 824
rect 304 706 356 758
rect 578 520 630 572
rect 578 454 630 506
rect 1990 709 2042 761
rect 1990 645 2042 697
rect 234 207 286 259
rect 298 207 350 259
rect 362 250 414 259
rect 426 250 478 259
rect 882 250 934 259
rect 946 250 998 259
rect 1010 250 1062 259
rect 1074 250 1126 259
rect 1206 250 1258 259
rect 1270 250 1322 259
rect 362 216 393 250
rect 393 216 414 250
rect 426 216 427 250
rect 427 216 466 250
rect 466 216 478 250
rect 882 216 904 250
rect 904 216 934 250
rect 946 216 977 250
rect 977 216 998 250
rect 1010 216 1011 250
rect 1011 216 1050 250
rect 1050 216 1062 250
rect 1074 216 1084 250
rect 1084 216 1123 250
rect 1123 216 1126 250
rect 1206 216 1230 250
rect 1230 216 1258 250
rect 1270 216 1303 250
rect 1303 216 1322 250
rect 362 207 414 216
rect 426 207 478 216
rect 882 207 934 216
rect 946 207 998 216
rect 1010 207 1062 216
rect 1074 207 1126 216
rect 1206 207 1258 216
rect 1270 207 1322 216
rect 1334 250 1386 259
rect 1334 216 1342 250
rect 1342 216 1376 250
rect 1376 216 1386 250
rect 1334 207 1386 216
rect 1398 250 1450 259
rect 3564 587 3616 593
rect 3564 553 3576 587
rect 3576 553 3610 587
rect 3610 553 3616 587
rect 3564 541 3616 553
rect 3564 511 3616 520
rect 3564 477 3576 511
rect 3576 477 3610 511
rect 3610 477 3616 511
rect 3564 468 3616 477
rect 3564 436 3616 447
rect 3564 402 3576 436
rect 3576 402 3610 436
rect 3610 402 3616 436
rect 3564 395 3616 402
rect 3564 361 3616 374
rect 3564 327 3576 361
rect 3576 327 3610 361
rect 3610 327 3616 361
rect 3564 322 3616 327
rect 3564 286 3616 301
rect 1854 250 1906 259
rect 1398 216 1415 250
rect 1415 216 1449 250
rect 1449 216 1450 250
rect 1854 216 1887 250
rect 1887 216 1906 250
rect 1398 207 1450 216
rect 1854 207 1906 216
rect 1918 250 1970 259
rect 1918 216 1926 250
rect 1926 216 1960 250
rect 1960 216 1970 250
rect 1918 207 1970 216
rect 1982 250 2034 259
rect 2210 250 2262 259
rect 1982 216 1999 250
rect 1999 216 2033 250
rect 2033 216 2034 250
rect 2210 216 2217 250
rect 2217 216 2251 250
rect 2251 216 2262 250
rect 1982 207 2034 216
rect 2210 207 2262 216
rect 2274 250 2326 259
rect 2570 250 2622 259
rect 2274 216 2289 250
rect 2289 216 2323 250
rect 2323 216 2326 250
rect 2570 216 2577 250
rect 2577 216 2611 250
rect 2611 216 2622 250
rect 2274 207 2326 216
rect 2570 207 2622 216
rect 2634 250 2686 259
rect 2634 216 2649 250
rect 2649 216 2683 250
rect 2683 216 2686 250
rect 2634 207 2686 216
rect 2698 250 2750 259
rect 2698 216 2721 250
rect 2721 216 2750 250
rect 2698 207 2750 216
rect 3564 252 3576 286
rect 3576 252 3610 286
rect 3610 252 3616 286
rect 3564 249 3616 252
rect 3564 211 3616 228
rect 3564 177 3576 211
rect 3576 177 3610 211
rect 3610 177 3616 211
rect 3564 176 3616 177
rect 2414 109 2466 161
rect 2478 109 2530 161
rect 3564 136 3616 156
rect 3564 104 3576 136
rect 3576 104 3610 136
rect 3610 104 3616 136
rect 3564 61 3616 84
rect 3564 32 3576 61
rect 3576 32 3610 61
rect 3610 32 3616 61
<< metal2 >>
tri -1086 2423 -1048 2461 se
rect -1048 2423 -852 2917
tri -1098 2411 -1086 2423 se
rect -1086 2411 -852 2423
tri -1150 2359 -1098 2411 se
rect -1098 2359 -852 2411
tri -1173 2336 -1150 2359 se
rect -1150 2336 -852 2359
tri -1206 2303 -1173 2336 se
rect -1173 2303 -852 2336
rect -1206 0 -852 2303
rect -824 2583 -772 2589
rect -824 2519 -772 2531
rect -824 0 -772 2467
rect -744 0 -476 2917
rect -420 0 -152 2917
rect -96 0 49 2917
rect 120 0 172 17828
rect 228 16935 496 17855
rect 228 454 276 16935
tri 276 16903 308 16935 nw
tri 352 16903 384 16935 ne
rect 304 12318 356 16751
rect 304 12254 356 12266
rect 304 824 356 12202
rect 304 758 356 772
rect 304 624 356 706
tri 276 454 306 484 sw
tri 354 454 384 484 se
rect 384 454 496 16935
rect 228 452 306 454
tri 306 452 308 454 sw
tri 352 452 354 454 se
rect 354 452 496 454
rect 228 259 496 452
rect 228 207 234 259
rect 286 207 298 259
rect 350 207 362 259
rect 414 207 426 259
rect 478 207 496 259
rect 228 0 496 207
rect 552 16935 820 17855
rect 552 572 656 16935
tri 656 16903 688 16935 nw
rect 552 520 578 572
rect 630 520 656 572
rect 552 506 656 520
rect 552 454 578 506
rect 630 454 656 506
rect 552 0 656 454
rect 876 259 1144 17855
rect 876 207 882 259
rect 934 207 946 259
rect 998 207 1010 259
rect 1062 207 1074 259
rect 1126 207 1144 259
rect 876 85 1144 207
tri 876 84 877 85 ne
rect 877 84 1144 85
tri 877 32 929 84 ne
rect 929 32 1144 84
tri 929 0 961 32 ne
rect 961 0 1144 32
rect 1200 259 1468 17855
rect 1524 625 1792 17855
rect 1848 16935 2081 17964
rect 2204 17671 2440 17964
rect 2124 17596 2176 17602
rect 2124 17532 2176 17544
rect 1848 1983 1934 16935
tri 1934 16903 1966 16935 nw
rect 1848 1931 1865 1983
rect 1917 1931 1934 1983
rect 1848 1917 1934 1931
rect 1848 1865 1865 1917
rect 1917 1865 1934 1917
rect 1848 1850 1934 1865
rect 1848 1798 1865 1850
rect 1917 1798 1934 1850
rect 1200 207 1206 259
rect 1258 207 1270 259
rect 1322 207 1334 259
rect 1386 207 1398 259
rect 1450 207 1468 259
rect 1200 0 1468 207
rect 1500 0 1816 569
rect 1848 468 1934 1798
rect 1990 12214 2042 16751
rect 1990 12150 2042 12162
rect 1990 761 2042 12098
rect 1990 697 2042 709
rect 1990 639 2042 645
tri 1934 468 1950 484 sw
rect 1848 452 1950 468
tri 1950 452 1966 468 sw
rect 1848 259 2081 452
rect 1848 207 1854 259
rect 1906 207 1918 259
rect 1970 207 1982 259
rect 2034 207 2081 259
rect 1848 0 2081 207
rect 2124 0 2176 17480
rect 2204 1983 2380 17671
tri 2380 17611 2440 17671 nw
rect 2256 1931 2328 1983
rect 2204 1917 2380 1931
rect 2256 1865 2328 1917
rect 2204 1850 2380 1865
rect 2256 1798 2328 1850
rect 2204 259 2380 1798
rect 2204 207 2210 259
rect 2262 207 2274 259
rect 2326 207 2380 259
rect 2204 0 2380 207
rect 2564 3586 2764 17862
rect 2820 17675 3042 17964
tri 3042 17675 3136 17769 sw
tri 2820 17582 2913 17675 ne
rect 2564 2177 2711 3586
tri 2711 3533 2764 3586 nw
tri 2819 3402 2913 3496 se
rect 2913 3403 3136 17675
rect 2913 3402 3098 3403
rect 2819 3365 3098 3402
tri 3098 3365 3136 3403 nw
tri 3178 3365 3192 3379 se
rect 3192 3365 3414 17964
rect 2739 2475 2791 2481
rect 2739 2411 2791 2423
rect 2739 2299 2791 2359
rect 2819 2395 3042 3365
tri 3042 3309 3098 3365 nw
tri 3122 3309 3178 3365 se
rect 3178 3309 3414 3365
tri 3098 3285 3122 3309 se
rect 3122 3285 3414 3309
rect 3098 2475 3414 3285
tri 3098 2451 3122 2475 ne
rect 3122 2451 3414 2475
tri 3042 2395 3098 2451 sw
tri 3122 2395 3178 2451 ne
rect 3178 2395 3414 2451
rect 2819 2388 3098 2395
tri 3098 2388 3105 2395 sw
tri 3178 2388 3185 2395 ne
rect 3185 2388 3414 2395
rect 2819 2358 3105 2388
tri 2819 2336 2841 2358 ne
rect 2841 2357 3105 2358
tri 3105 2357 3136 2388 sw
tri 3185 2384 3189 2388 ne
rect 2841 2336 3136 2357
tri 2841 2306 2871 2336 ne
rect 2871 2306 3136 2336
tri 2791 2299 2798 2306 sw
tri 2871 2299 2878 2306 ne
rect 2878 2299 3136 2306
rect 2739 2293 2798 2299
tri 2798 2293 2804 2299 sw
tri 2878 2293 2884 2299 ne
rect 2884 2293 3136 2299
rect 2739 2284 2804 2293
tri 2739 2241 2782 2284 ne
rect 2782 2241 2804 2284
tri 2804 2241 2856 2293 sw
tri 2884 2264 2913 2293 ne
tri 2782 2229 2794 2241 ne
rect 2794 2229 2856 2241
tri 2856 2229 2868 2241 sw
tri 2794 2225 2798 2229 ne
rect 2798 2225 2868 2229
tri 2868 2225 2872 2229 sw
tri 2798 2203 2820 2225 ne
tri 2711 2177 2735 2201 sw
rect 2564 2165 2735 2177
tri 2735 2165 2747 2177 sw
rect 2564 2148 2747 2165
tri 2747 2148 2764 2165 sw
rect 2564 1983 2764 2148
rect 2616 1931 2638 1983
rect 2690 1931 2712 1983
rect 2564 1917 2764 1931
rect 2616 1865 2638 1917
rect 2690 1865 2712 1917
rect 2564 1850 2764 1865
rect 2616 1798 2638 1850
rect 2690 1798 2712 1850
rect 2564 259 2764 1798
rect 2564 207 2570 259
rect 2622 207 2634 259
rect 2686 207 2698 259
rect 2750 207 2764 259
rect 2408 109 2414 161
rect 2466 109 2478 161
rect 2530 109 2536 161
rect 2436 0 2488 109
rect 2564 32 2764 207
tri 2564 0 2596 32 ne
rect 2596 0 2764 32
rect 2820 0 2872 2225
rect 2913 0 3136 2293
rect 3189 2336 3195 2388
rect 3247 2336 3259 2388
rect 3311 2336 3323 2388
rect 3375 2336 3414 2388
rect 3189 2293 3414 2336
rect 3241 2241 3414 2293
rect 3189 2229 3414 2241
rect 3241 2177 3414 2229
rect 3189 2165 3414 2177
rect 3241 2113 3414 2165
rect 3189 2101 3414 2113
rect 3241 2049 3414 2101
rect 3189 2043 3414 2049
rect 3192 1730 3414 2043
rect 3189 1724 3414 1730
rect 3241 1672 3414 1724
rect 3189 1660 3414 1672
rect 3241 1608 3414 1660
rect 3189 1596 3414 1608
rect 3241 1544 3414 1596
rect 3189 1532 3414 1544
rect 3241 1480 3414 1532
rect 3189 1468 3414 1480
rect 3241 1416 3414 1468
rect 3189 1404 3414 1416
rect 3241 1352 3414 1404
rect 3189 1340 3414 1352
rect 3241 1288 3414 1340
rect 3189 1276 3414 1288
rect 3241 1224 3414 1276
rect 3189 1212 3414 1224
rect 3241 1160 3414 1212
rect 3189 1148 3414 1160
rect 3241 1096 3414 1148
rect 3189 1059 3414 1096
rect 3189 1007 3195 1059
rect 3247 1007 3259 1059
rect 3311 1007 3323 1059
rect 3375 1007 3414 1059
rect 3192 0 3414 1007
rect 3470 593 3781 18198
rect 3470 541 3564 593
rect 3616 541 3781 593
rect 3470 520 3781 541
rect 3470 468 3564 520
rect 3616 468 3781 520
rect 3470 447 3781 468
rect 3470 395 3564 447
rect 3616 395 3781 447
rect 3470 374 3781 395
rect 3470 322 3564 374
rect 3616 322 3781 374
rect 3470 301 3781 322
rect 3470 249 3564 301
rect 3616 249 3781 301
rect 3470 228 3781 249
rect 3470 176 3564 228
rect 3616 176 3781 228
rect 3470 156 3781 176
rect 3470 104 3564 156
rect 3616 104 3781 156
rect 3470 84 3781 104
rect 3470 32 3564 84
rect 3616 32 3781 84
rect 3470 0 3781 32
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform -1 0 3672 0 1 2226
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_1
timestamp 1704896540
transform -1 0 3672 0 1 1914
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_2
timestamp 1704896540
transform -1 0 3672 0 1 1602
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_3
timestamp 1704896540
transform -1 0 3672 0 1 1290
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_4
timestamp 1704896540
transform -1 0 3906 0 1 1154
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_5
timestamp 1704896540
transform -1 0 3906 0 1 1446
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_6
timestamp 1704896540
transform -1 0 3906 0 1 1758
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1704896540
transform -1 0 3877 0 1 2070
box 0 0 1 1
use L1M1_CDNS_52468879185940  L1M1_CDNS_52468879185940_0
timestamp 1704896540
transform 0 -1 -312 1 0 119
box -12 -6 2782 40
use L1M1_CDNS_524688791851140  L1M1_CDNS_524688791851140_0
timestamp 1704896540
transform -1 0 3533 0 1 27
box -12 -6 3718 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 2176 -1 0 17602
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 0 -1 356 1 0 12196
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 0 -1 2042 1 0 12092
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 0 -1 -772 1 0 2461
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1704896540
transform 0 1 1530 1 0 17663
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_1
timestamp 1704896540
transform 0 1 1207 1 0 17663
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_2
timestamp 1704896540
transform 0 1 888 1 0 17663
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_3
timestamp 1704896540
transform 0 1 563 1 0 17663
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_4
timestamp 1704896540
transform 0 1 238 1 0 17663
box 0 0 192 244
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1704896540
transform 0 1 2564 1 0 17663
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1704896540
transform 0 1 1875 1 0 17663
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1704896540
transform 0 -1 2428 1 0 17663
box 0 0 192 180
use nfet_CDNS_524688791851143  nfet_CDNS_524688791851143_0
timestamp 1704896540
transform 0 -1 3906 1 0 1179
box -79 -52 1118 652
use sky130_fd_io__refgen_res_ntwk_a  sky130_fd_io__refgen_res_ntwk_a_0
timestamp 1704896540
transform -1 0 2993 0 1 278
box -88 -88 1318 17258
use sky130_fd_io__refgen_res_ntwk_a  sky130_fd_io__refgen_res_ntwk_a_1
timestamp 1704896540
transform 1 0 443 0 1 278
box -88 -88 1318 17258
<< labels >>
flabel comment s 70 17571 70 17571 3 FreeSans 200 0 0 0 en_outop_h_n
flabel comment s 2144 13 2144 13 3 FreeSans 200 90 0 0 en_outop_h_n
flabel comment s -1233 2581 -1233 2581 3 FreeSans 200 0 0 0 en_inpop_h
flabel comment s -800 13 -800 13 3 FreeSans 200 90 0 0 en_inpop_h
flabel comment s 1656 53 1656 53 3 FreeSans 200 90 0 0 vpb
flabel comment s 143 13 143 13 3 FreeSans 200 90 0 0 biasen_n
flabel comment s 144 17708 144 17708 3 FreeSans 200 270 0 0 biasen_n
flabel comment s 3022 10 3022 10 3 FreeSans 200 90 0 0 vpwr
flabel comment s 2935 17959 2935 17959 3 FreeSans 200 270 0 0 vpwr
flabel metal1 s -1262 0 -1226 67 3 FreeSans 200 0 0 0 vcc
port 2 nsew
flabel metal1 s 0 12196 34 12260 3 FreeSans 200 0 0 0 fb_out
port 3 nsew
flabel metal1 s 1 12092 34 12156 3 FreeSans 200 0 0 0 res_stack
port 4 nsew
flabel metal2 s 876 17793 1144 17828 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s -744 2876 -476 2917 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s -1206 0 -852 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s -744 0 -476 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s -1003 11 -1003 11 3 FreeSans 200 90 0 0 vgnd
flabel metal2 s -1048 2876 -852 2917 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s -96 2896 49 2917 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 3470 18175 3616 18198 3 FreeSans 200 270 0 0 vcc
port 2 nsew
flabel metal2 s 3470 0 3616 21 3 FreeSans 200 90 0 0 vcc
port 2 nsew
flabel metal2 s -420 2896 -152 2917 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 2596 0 2764 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 2204 0 2380 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 1848 17921 2081 17964 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 1524 17793 1792 17828 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 1200 0 1468 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 961 0 1144 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 552 0 656 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 228 0 496 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s -420 0 -152 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 2436 0 2488 21 3 FreeSans 200 90 0 0 vohref_0p5
port 6 nsew
flabel metal2 s -96 0 49 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 3192 17921 3414 17964 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 2204 17921 2440 17964 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 1848 0 2081 21 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 1200 17793 1468 17828 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 3192 0 3414 43 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 2820 0 2872 21 3 FreeSans 200 90 0 0 sel_vohref_0p5
port 7 nsew
flabel metal2 s 228 17793 496 17828 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
flabel metal2 s 552 17793 820 17828 3 FreeSans 200 270 0 0 vgnd
port 5 nsew
<< properties >>
string GDS_END 79584798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79515280
string path 63.400 3.375 60.200 3.375 
<< end >>
