magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 98 157 800 203
rect 1 21 800 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 176 47 206 177
rect 260 47 290 177
rect 344 47 374 177
rect 428 47 458 177
rect 512 47 542 177
rect 596 47 626 177
rect 692 47 722 177
<< scpmoshvt >>
rect 79 360 109 444
rect 176 297 206 497
rect 260 297 290 497
rect 344 297 374 497
rect 428 297 458 497
rect 512 297 542 497
rect 596 297 626 497
rect 692 297 722 497
<< ndiff >>
rect 124 131 176 177
rect 27 108 79 131
rect 27 74 35 108
rect 69 74 79 108
rect 27 47 79 74
rect 109 97 176 131
rect 109 63 124 97
rect 158 63 176 97
rect 109 47 176 63
rect 206 164 260 177
rect 206 130 216 164
rect 250 130 260 164
rect 206 96 260 130
rect 206 62 216 96
rect 250 62 260 96
rect 206 47 260 62
rect 290 97 344 177
rect 290 63 300 97
rect 334 63 344 97
rect 290 47 344 63
rect 374 101 428 177
rect 374 67 384 101
rect 418 67 428 101
rect 374 47 428 67
rect 458 97 512 177
rect 458 63 468 97
rect 502 63 512 97
rect 458 47 512 63
rect 542 111 596 177
rect 542 77 552 111
rect 586 77 596 111
rect 542 47 596 77
rect 626 97 692 177
rect 626 63 636 97
rect 670 63 692 97
rect 626 47 692 63
rect 722 111 774 177
rect 722 77 732 111
rect 766 77 774 111
rect 722 47 774 77
<< pdiff >>
rect 124 476 176 497
rect 124 444 132 476
rect 27 412 79 444
rect 27 378 35 412
rect 69 378 79 412
rect 27 360 79 378
rect 109 442 132 444
rect 166 442 176 476
rect 109 360 176 442
rect 124 297 176 360
rect 206 340 260 497
rect 206 306 216 340
rect 250 306 260 340
rect 206 297 260 306
rect 290 476 344 497
rect 290 442 300 476
rect 334 442 344 476
rect 290 297 344 442
rect 374 340 428 497
rect 374 306 384 340
rect 418 306 428 340
rect 374 297 428 306
rect 458 476 512 497
rect 458 442 468 476
rect 502 442 512 476
rect 458 297 512 442
rect 542 297 596 497
rect 626 297 692 497
rect 722 476 774 497
rect 722 442 732 476
rect 766 442 774 476
rect 722 297 774 442
<< ndiffc >>
rect 35 74 69 108
rect 124 63 158 97
rect 216 130 250 164
rect 216 62 250 96
rect 300 63 334 97
rect 384 67 418 101
rect 468 63 502 97
rect 552 77 586 111
rect 636 63 670 97
rect 732 77 766 111
<< pdiffc >>
rect 35 378 69 412
rect 132 442 166 476
rect 216 306 250 340
rect 300 442 334 476
rect 384 306 418 340
rect 468 442 502 476
rect 732 442 766 476
<< poly >>
rect 176 497 206 523
rect 260 497 290 523
rect 344 497 374 523
rect 428 497 458 523
rect 512 497 542 523
rect 596 497 626 523
rect 692 497 722 523
rect 79 444 109 470
rect 79 265 109 360
rect 22 249 109 265
rect 22 215 35 249
rect 69 215 109 249
rect 22 199 109 215
rect 79 131 109 199
rect 176 265 206 297
rect 260 265 290 297
rect 344 265 374 297
rect 428 265 458 297
rect 512 265 542 297
rect 596 265 626 297
rect 692 265 722 297
rect 176 249 458 265
rect 176 215 271 249
rect 305 215 339 249
rect 373 215 407 249
rect 441 215 458 249
rect 176 199 458 215
rect 500 249 554 265
rect 500 215 510 249
rect 544 215 554 249
rect 500 199 554 215
rect 596 249 650 265
rect 596 215 606 249
rect 640 215 650 249
rect 596 199 650 215
rect 692 249 746 265
rect 692 215 702 249
rect 736 215 746 249
rect 692 199 746 215
rect 176 177 206 199
rect 260 177 290 199
rect 344 177 374 199
rect 428 177 458 199
rect 512 177 542 199
rect 596 177 626 199
rect 692 177 722 199
rect 79 21 109 47
rect 176 21 206 47
rect 260 21 290 47
rect 344 21 374 47
rect 428 21 458 47
rect 512 21 542 47
rect 596 21 626 47
rect 692 21 722 47
<< polycont >>
rect 35 215 69 249
rect 271 215 305 249
rect 339 215 373 249
rect 407 215 441 249
rect 510 215 544 249
rect 606 215 640 249
rect 702 215 736 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 110 476 182 527
rect 17 412 69 444
rect 110 442 132 476
rect 166 442 182 476
rect 284 476 350 527
rect 284 442 300 476
rect 334 442 350 476
rect 451 476 519 527
rect 451 442 468 476
rect 502 442 519 476
rect 704 476 811 485
rect 704 442 732 476
rect 766 442 811 476
rect 17 378 35 412
rect 69 378 724 408
rect 17 374 724 378
rect 17 362 153 374
rect 17 249 85 328
rect 17 215 35 249
rect 69 215 85 249
rect 119 181 153 362
rect 17 147 153 181
rect 187 306 216 340
rect 250 306 384 340
rect 418 306 444 340
rect 187 283 444 306
rect 480 283 544 340
rect 187 181 221 283
rect 507 249 544 283
rect 255 215 271 249
rect 305 215 339 249
rect 373 215 407 249
rect 441 215 473 249
rect 187 164 405 181
rect 187 147 216 164
rect 17 108 69 147
rect 200 130 216 147
rect 250 147 405 164
rect 250 130 266 147
rect 17 74 35 108
rect 17 58 69 74
rect 124 97 158 113
rect 124 17 158 63
rect 200 96 266 130
rect 371 117 405 147
rect 439 178 473 215
rect 507 215 510 249
rect 507 199 544 215
rect 578 249 640 340
rect 578 215 606 249
rect 578 199 640 215
rect 678 265 724 374
rect 678 249 736 265
rect 678 215 702 249
rect 678 199 736 215
rect 439 165 480 178
rect 770 165 811 442
rect 439 144 811 165
rect 450 131 811 144
rect 200 62 216 96
rect 250 62 266 96
rect 200 57 266 62
rect 300 97 334 113
rect 300 17 334 63
rect 371 101 418 117
rect 371 67 384 101
rect 552 111 586 131
rect 371 51 418 67
rect 452 63 468 97
rect 502 63 518 97
rect 452 17 518 63
rect 732 121 811 131
rect 732 111 783 121
rect 552 61 586 77
rect 620 63 636 97
rect 670 63 698 97
rect 620 17 698 63
rect 766 77 783 111
rect 732 61 783 77
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 490 289 524 323 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 200 180 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or3b_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1048222
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1041788
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
