magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 176 1426
<< mvnmos >>
rect 0 0 100 1400
<< mvndiff >>
rect -50 0 0 1400
rect 100 0 150 1400
<< poly >>
rect 0 1400 100 1432
rect 0 -32 100 0
<< metal1 >>
rect -51 -16 -5 1410
rect 105 -16 151 1410
use hvDFM1sd2_CDNS_52468879185610  hvDFM1sd2_CDNS_52468879185610_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 82 1426
use hvDFM1sd2_CDNS_52468879185610  hvDFM1sd2_CDNS_52468879185610_1
timestamp 1704896540
transform 1 0 100 0 1 0
box -26 -26 82 1426
<< labels >>
flabel comment s -28 697 -28 697 0 FreeSans 300 0 0 0 S
flabel comment s 128 697 128 697 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6693880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6692986
<< end >>
