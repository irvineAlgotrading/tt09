magic
tech sky130B
timestamp 1704896540
<< locali >>
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 108 17
rect 125 0 144 17
rect 161 0 180 17
rect 197 0 216 17
rect 233 0 252 17
rect 269 0 288 17
rect 305 0 324 17
rect 341 0 360 17
rect 377 0 396 17
rect 413 0 432 17
rect 449 0 468 17
rect 485 0 504 17
rect 521 0 540 17
rect 557 0 576 17
rect 593 0 612 17
rect 629 0 648 17
rect 665 0 684 17
rect 701 0 720 17
rect 737 0 756 17
rect 773 0 792 17
rect 809 0 828 17
rect 845 0 864 17
rect 881 0 900 17
rect 917 0 936 17
rect 953 0 972 17
rect 989 0 1008 17
rect 1025 0 1044 17
rect 1061 0 1080 17
rect 1097 0 1116 17
rect 1133 0 1152 17
rect 1169 0 1188 17
rect 1205 0 1224 17
rect 1241 0 1260 17
rect 1277 0 1296 17
rect 1313 0 1332 17
rect 1349 0 1368 17
rect 1385 0 1404 17
rect 1421 0 1440 17
rect 1457 0 1476 17
rect 1493 0 1512 17
rect 1529 0 1548 17
rect 1565 0 1584 17
rect 1601 0 1620 17
rect 1637 0 1656 17
rect 1673 0 1692 17
rect 1709 0 1728 17
rect 1745 0 1764 17
rect 1781 0 1800 17
rect 1817 0 1836 17
rect 1853 0 1872 17
rect 1889 0 1908 17
rect 1925 0 1944 17
rect 1961 0 1980 17
rect 1997 0 2016 17
rect 2033 0 2052 17
rect 2069 0 2088 17
rect 2105 0 2124 17
rect 2141 0 2160 17
rect 2177 0 2196 17
rect 2213 0 2232 17
rect 2249 0 2268 17
rect 2285 0 2304 17
rect 2321 0 2340 17
rect 2357 0 2376 17
rect 2393 0 2412 17
rect 2429 0 2448 17
rect 2465 0 2484 17
rect 2501 0 2520 17
rect 2537 0 2556 17
rect 2573 0 2592 17
rect 2609 0 2628 17
rect 2645 0 2664 17
rect 2681 0 2700 17
rect 2717 0 2736 17
rect 2753 0 2772 17
rect 2789 0 2808 17
rect 2825 0 2844 17
rect 2861 0 2880 17
rect 2897 0 2916 17
rect 2933 0 2952 17
rect 2969 0 2988 17
rect 3005 0 3024 17
<< viali >>
rect 0 0 17 17
rect 36 0 53 17
rect 72 0 89 17
rect 108 0 125 17
rect 144 0 161 17
rect 180 0 197 17
rect 216 0 233 17
rect 252 0 269 17
rect 288 0 305 17
rect 324 0 341 17
rect 360 0 377 17
rect 396 0 413 17
rect 432 0 449 17
rect 468 0 485 17
rect 504 0 521 17
rect 540 0 557 17
rect 576 0 593 17
rect 612 0 629 17
rect 648 0 665 17
rect 684 0 701 17
rect 720 0 737 17
rect 756 0 773 17
rect 792 0 809 17
rect 828 0 845 17
rect 864 0 881 17
rect 900 0 917 17
rect 936 0 953 17
rect 972 0 989 17
rect 1008 0 1025 17
rect 1044 0 1061 17
rect 1080 0 1097 17
rect 1116 0 1133 17
rect 1152 0 1169 17
rect 1188 0 1205 17
rect 1224 0 1241 17
rect 1260 0 1277 17
rect 1296 0 1313 17
rect 1332 0 1349 17
rect 1368 0 1385 17
rect 1404 0 1421 17
rect 1440 0 1457 17
rect 1476 0 1493 17
rect 1512 0 1529 17
rect 1548 0 1565 17
rect 1584 0 1601 17
rect 1620 0 1637 17
rect 1656 0 1673 17
rect 1692 0 1709 17
rect 1728 0 1745 17
rect 1764 0 1781 17
rect 1800 0 1817 17
rect 1836 0 1853 17
rect 1872 0 1889 17
rect 1908 0 1925 17
rect 1944 0 1961 17
rect 1980 0 1997 17
rect 2016 0 2033 17
rect 2052 0 2069 17
rect 2088 0 2105 17
rect 2124 0 2141 17
rect 2160 0 2177 17
rect 2196 0 2213 17
rect 2232 0 2249 17
rect 2268 0 2285 17
rect 2304 0 2321 17
rect 2340 0 2357 17
rect 2376 0 2393 17
rect 2412 0 2429 17
rect 2448 0 2465 17
rect 2484 0 2501 17
rect 2520 0 2537 17
rect 2556 0 2573 17
rect 2592 0 2609 17
rect 2628 0 2645 17
rect 2664 0 2681 17
rect 2700 0 2717 17
rect 2736 0 2753 17
rect 2772 0 2789 17
rect 2808 0 2825 17
rect 2844 0 2861 17
rect 2880 0 2897 17
rect 2916 0 2933 17
rect 2952 0 2969 17
rect 2988 0 3005 17
rect 3024 0 3041 17
<< metal1 >>
rect -6 17 3047 20
rect -6 0 0 17
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 108 17
rect 125 0 144 17
rect 161 0 180 17
rect 197 0 216 17
rect 233 0 252 17
rect 269 0 288 17
rect 305 0 324 17
rect 341 0 360 17
rect 377 0 396 17
rect 413 0 432 17
rect 449 0 468 17
rect 485 0 504 17
rect 521 0 540 17
rect 557 0 576 17
rect 593 0 612 17
rect 629 0 648 17
rect 665 0 684 17
rect 701 0 720 17
rect 737 0 756 17
rect 773 0 792 17
rect 809 0 828 17
rect 845 0 864 17
rect 881 0 900 17
rect 917 0 936 17
rect 953 0 972 17
rect 989 0 1008 17
rect 1025 0 1044 17
rect 1061 0 1080 17
rect 1097 0 1116 17
rect 1133 0 1152 17
rect 1169 0 1188 17
rect 1205 0 1224 17
rect 1241 0 1260 17
rect 1277 0 1296 17
rect 1313 0 1332 17
rect 1349 0 1368 17
rect 1385 0 1404 17
rect 1421 0 1440 17
rect 1457 0 1476 17
rect 1493 0 1512 17
rect 1529 0 1548 17
rect 1565 0 1584 17
rect 1601 0 1620 17
rect 1637 0 1656 17
rect 1673 0 1692 17
rect 1709 0 1728 17
rect 1745 0 1764 17
rect 1781 0 1800 17
rect 1817 0 1836 17
rect 1853 0 1872 17
rect 1889 0 1908 17
rect 1925 0 1944 17
rect 1961 0 1980 17
rect 1997 0 2016 17
rect 2033 0 2052 17
rect 2069 0 2088 17
rect 2105 0 2124 17
rect 2141 0 2160 17
rect 2177 0 2196 17
rect 2213 0 2232 17
rect 2249 0 2268 17
rect 2285 0 2304 17
rect 2321 0 2340 17
rect 2357 0 2376 17
rect 2393 0 2412 17
rect 2429 0 2448 17
rect 2465 0 2484 17
rect 2501 0 2520 17
rect 2537 0 2556 17
rect 2573 0 2592 17
rect 2609 0 2628 17
rect 2645 0 2664 17
rect 2681 0 2700 17
rect 2717 0 2736 17
rect 2753 0 2772 17
rect 2789 0 2808 17
rect 2825 0 2844 17
rect 2861 0 2880 17
rect 2897 0 2916 17
rect 2933 0 2952 17
rect 2969 0 2988 17
rect 3005 0 3024 17
rect 3041 0 3047 17
rect -6 -3 3047 0
<< properties >>
string GDS_END 80037614
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80032042
<< end >>
