magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 2754 897
<< pwell >>
rect 6 43 2605 317
rect -26 -43 2714 43
<< mvnmos >>
rect 85 141 185 291
rect 241 141 341 291
rect 397 141 497 291
rect 553 141 653 291
rect 709 141 809 291
rect 865 141 965 291
rect 1021 141 1121 291
rect 1177 141 1277 291
rect 1333 141 1433 291
rect 1489 141 1589 291
rect 1645 141 1745 291
rect 1801 141 1901 291
rect 1957 141 2057 291
rect 2113 141 2213 291
rect 2269 141 2369 291
rect 2425 141 2525 291
<< mvpmos >>
rect 86 443 186 743
rect 242 443 342 743
rect 398 443 498 743
rect 554 443 654 743
rect 710 443 810 743
rect 866 443 966 743
rect 1022 443 1122 743
rect 1178 443 1278 743
rect 1334 443 1434 743
rect 1490 443 1590 743
rect 1646 443 1746 743
rect 1802 443 1902 743
rect 1958 443 2058 743
rect 2114 443 2214 743
rect 2270 443 2370 743
rect 2426 443 2526 743
<< mvndiff >>
rect 32 279 85 291
rect 32 245 40 279
rect 74 245 85 279
rect 32 206 85 245
rect 32 172 40 206
rect 74 172 85 206
rect 32 141 85 172
rect 185 283 241 291
rect 185 249 196 283
rect 230 249 241 283
rect 185 209 241 249
rect 185 175 196 209
rect 230 175 241 209
rect 185 141 241 175
rect 341 279 397 291
rect 341 245 352 279
rect 386 245 397 279
rect 341 206 397 245
rect 341 172 352 206
rect 386 172 397 206
rect 341 141 397 172
rect 497 283 553 291
rect 497 249 508 283
rect 542 249 553 283
rect 497 209 553 249
rect 497 175 508 209
rect 542 175 553 209
rect 497 141 553 175
rect 653 279 709 291
rect 653 245 664 279
rect 698 245 709 279
rect 653 206 709 245
rect 653 172 664 206
rect 698 172 709 206
rect 653 141 709 172
rect 809 283 865 291
rect 809 249 820 283
rect 854 249 865 283
rect 809 209 865 249
rect 809 175 820 209
rect 854 175 865 209
rect 809 141 865 175
rect 965 279 1021 291
rect 965 245 976 279
rect 1010 245 1021 279
rect 965 206 1021 245
rect 965 172 976 206
rect 1010 172 1021 206
rect 965 141 1021 172
rect 1121 283 1177 291
rect 1121 249 1132 283
rect 1166 249 1177 283
rect 1121 209 1177 249
rect 1121 175 1132 209
rect 1166 175 1177 209
rect 1121 141 1177 175
rect 1277 279 1333 291
rect 1277 245 1288 279
rect 1322 245 1333 279
rect 1277 206 1333 245
rect 1277 172 1288 206
rect 1322 172 1333 206
rect 1277 141 1333 172
rect 1433 283 1489 291
rect 1433 249 1444 283
rect 1478 249 1489 283
rect 1433 209 1489 249
rect 1433 175 1444 209
rect 1478 175 1489 209
rect 1433 141 1489 175
rect 1589 279 1645 291
rect 1589 245 1600 279
rect 1634 245 1645 279
rect 1589 206 1645 245
rect 1589 172 1600 206
rect 1634 172 1645 206
rect 1589 141 1645 172
rect 1745 283 1801 291
rect 1745 249 1756 283
rect 1790 249 1801 283
rect 1745 209 1801 249
rect 1745 175 1756 209
rect 1790 175 1801 209
rect 1745 141 1801 175
rect 1901 279 1957 291
rect 1901 245 1912 279
rect 1946 245 1957 279
rect 1901 206 1957 245
rect 1901 172 1912 206
rect 1946 172 1957 206
rect 1901 141 1957 172
rect 2057 283 2113 291
rect 2057 249 2068 283
rect 2102 249 2113 283
rect 2057 209 2113 249
rect 2057 175 2068 209
rect 2102 175 2113 209
rect 2057 141 2113 175
rect 2213 279 2269 291
rect 2213 245 2224 279
rect 2258 245 2269 279
rect 2213 206 2269 245
rect 2213 172 2224 206
rect 2258 172 2269 206
rect 2213 141 2269 172
rect 2369 283 2425 291
rect 2369 249 2380 283
rect 2414 249 2425 283
rect 2369 209 2425 249
rect 2369 175 2380 209
rect 2414 175 2425 209
rect 2369 141 2425 175
rect 2525 279 2579 291
rect 2525 245 2536 279
rect 2570 245 2579 279
rect 2525 206 2579 245
rect 2525 172 2536 206
rect 2570 172 2579 206
rect 2525 141 2579 172
<< mvpdiff >>
rect 33 731 86 743
rect 33 697 41 731
rect 75 697 86 731
rect 33 663 86 697
rect 33 629 41 663
rect 75 629 86 663
rect 33 557 86 629
rect 33 523 41 557
rect 75 523 86 557
rect 33 489 86 523
rect 33 455 41 489
rect 75 455 86 489
rect 33 443 86 455
rect 186 735 242 743
rect 186 701 197 735
rect 231 701 242 735
rect 186 667 242 701
rect 186 633 197 667
rect 231 633 242 667
rect 186 553 242 633
rect 186 519 197 553
rect 231 519 242 553
rect 186 485 242 519
rect 186 451 197 485
rect 231 451 242 485
rect 186 443 242 451
rect 342 735 398 743
rect 342 701 353 735
rect 387 701 398 735
rect 342 667 398 701
rect 342 633 353 667
rect 387 633 398 667
rect 342 553 398 633
rect 342 519 353 553
rect 387 519 398 553
rect 342 485 398 519
rect 342 451 353 485
rect 387 451 398 485
rect 342 443 398 451
rect 498 735 554 743
rect 498 701 509 735
rect 543 701 554 735
rect 498 667 554 701
rect 498 633 509 667
rect 543 633 554 667
rect 498 553 554 633
rect 498 519 509 553
rect 543 519 554 553
rect 498 485 554 519
rect 498 451 509 485
rect 543 451 554 485
rect 498 443 554 451
rect 654 735 710 743
rect 654 701 665 735
rect 699 701 710 735
rect 654 667 710 701
rect 654 633 665 667
rect 699 633 710 667
rect 654 553 710 633
rect 654 519 665 553
rect 699 519 710 553
rect 654 485 710 519
rect 654 451 665 485
rect 699 451 710 485
rect 654 443 710 451
rect 810 735 866 743
rect 810 701 821 735
rect 855 701 866 735
rect 810 667 866 701
rect 810 633 821 667
rect 855 633 866 667
rect 810 553 866 633
rect 810 519 821 553
rect 855 519 866 553
rect 810 485 866 519
rect 810 451 821 485
rect 855 451 866 485
rect 810 443 866 451
rect 966 735 1022 743
rect 966 701 977 735
rect 1011 701 1022 735
rect 966 667 1022 701
rect 966 633 977 667
rect 1011 633 1022 667
rect 966 553 1022 633
rect 966 519 977 553
rect 1011 519 1022 553
rect 966 485 1022 519
rect 966 451 977 485
rect 1011 451 1022 485
rect 966 443 1022 451
rect 1122 735 1178 743
rect 1122 701 1133 735
rect 1167 701 1178 735
rect 1122 667 1178 701
rect 1122 633 1133 667
rect 1167 633 1178 667
rect 1122 553 1178 633
rect 1122 519 1133 553
rect 1167 519 1178 553
rect 1122 485 1178 519
rect 1122 451 1133 485
rect 1167 451 1178 485
rect 1122 443 1178 451
rect 1278 735 1334 743
rect 1278 701 1289 735
rect 1323 701 1334 735
rect 1278 667 1334 701
rect 1278 633 1289 667
rect 1323 633 1334 667
rect 1278 553 1334 633
rect 1278 519 1289 553
rect 1323 519 1334 553
rect 1278 485 1334 519
rect 1278 451 1289 485
rect 1323 451 1334 485
rect 1278 443 1334 451
rect 1434 735 1490 743
rect 1434 701 1445 735
rect 1479 701 1490 735
rect 1434 667 1490 701
rect 1434 633 1445 667
rect 1479 633 1490 667
rect 1434 553 1490 633
rect 1434 519 1445 553
rect 1479 519 1490 553
rect 1434 485 1490 519
rect 1434 451 1445 485
rect 1479 451 1490 485
rect 1434 443 1490 451
rect 1590 735 1646 743
rect 1590 701 1601 735
rect 1635 701 1646 735
rect 1590 667 1646 701
rect 1590 633 1601 667
rect 1635 633 1646 667
rect 1590 553 1646 633
rect 1590 519 1601 553
rect 1635 519 1646 553
rect 1590 485 1646 519
rect 1590 451 1601 485
rect 1635 451 1646 485
rect 1590 443 1646 451
rect 1746 735 1802 743
rect 1746 701 1757 735
rect 1791 701 1802 735
rect 1746 667 1802 701
rect 1746 633 1757 667
rect 1791 633 1802 667
rect 1746 553 1802 633
rect 1746 519 1757 553
rect 1791 519 1802 553
rect 1746 485 1802 519
rect 1746 451 1757 485
rect 1791 451 1802 485
rect 1746 443 1802 451
rect 1902 735 1958 743
rect 1902 701 1913 735
rect 1947 701 1958 735
rect 1902 667 1958 701
rect 1902 633 1913 667
rect 1947 633 1958 667
rect 1902 553 1958 633
rect 1902 519 1913 553
rect 1947 519 1958 553
rect 1902 485 1958 519
rect 1902 451 1913 485
rect 1947 451 1958 485
rect 1902 443 1958 451
rect 2058 735 2114 743
rect 2058 701 2069 735
rect 2103 701 2114 735
rect 2058 667 2114 701
rect 2058 633 2069 667
rect 2103 633 2114 667
rect 2058 553 2114 633
rect 2058 519 2069 553
rect 2103 519 2114 553
rect 2058 485 2114 519
rect 2058 451 2069 485
rect 2103 451 2114 485
rect 2058 443 2114 451
rect 2214 735 2270 743
rect 2214 701 2225 735
rect 2259 701 2270 735
rect 2214 667 2270 701
rect 2214 633 2225 667
rect 2259 633 2270 667
rect 2214 553 2270 633
rect 2214 519 2225 553
rect 2259 519 2270 553
rect 2214 485 2270 519
rect 2214 451 2225 485
rect 2259 451 2270 485
rect 2214 443 2270 451
rect 2370 735 2426 743
rect 2370 701 2381 735
rect 2415 701 2426 735
rect 2370 667 2426 701
rect 2370 633 2381 667
rect 2415 633 2426 667
rect 2370 553 2426 633
rect 2370 519 2381 553
rect 2415 519 2426 553
rect 2370 485 2426 519
rect 2370 451 2381 485
rect 2415 451 2426 485
rect 2370 443 2426 451
rect 2526 731 2579 743
rect 2526 697 2537 731
rect 2571 697 2579 731
rect 2526 663 2579 697
rect 2526 629 2537 663
rect 2571 629 2579 663
rect 2526 557 2579 629
rect 2526 523 2537 557
rect 2571 523 2579 557
rect 2526 489 2579 523
rect 2526 455 2537 489
rect 2571 455 2579 489
rect 2526 443 2579 455
<< mvndiffc >>
rect 40 245 74 279
rect 40 172 74 206
rect 196 249 230 283
rect 196 175 230 209
rect 352 245 386 279
rect 352 172 386 206
rect 508 249 542 283
rect 508 175 542 209
rect 664 245 698 279
rect 664 172 698 206
rect 820 249 854 283
rect 820 175 854 209
rect 976 245 1010 279
rect 976 172 1010 206
rect 1132 249 1166 283
rect 1132 175 1166 209
rect 1288 245 1322 279
rect 1288 172 1322 206
rect 1444 249 1478 283
rect 1444 175 1478 209
rect 1600 245 1634 279
rect 1600 172 1634 206
rect 1756 249 1790 283
rect 1756 175 1790 209
rect 1912 245 1946 279
rect 1912 172 1946 206
rect 2068 249 2102 283
rect 2068 175 2102 209
rect 2224 245 2258 279
rect 2224 172 2258 206
rect 2380 249 2414 283
rect 2380 175 2414 209
rect 2536 245 2570 279
rect 2536 172 2570 206
<< mvpdiffc >>
rect 41 697 75 731
rect 41 629 75 663
rect 41 523 75 557
rect 41 455 75 489
rect 197 701 231 735
rect 197 633 231 667
rect 197 519 231 553
rect 197 451 231 485
rect 353 701 387 735
rect 353 633 387 667
rect 353 519 387 553
rect 353 451 387 485
rect 509 701 543 735
rect 509 633 543 667
rect 509 519 543 553
rect 509 451 543 485
rect 665 701 699 735
rect 665 633 699 667
rect 665 519 699 553
rect 665 451 699 485
rect 821 701 855 735
rect 821 633 855 667
rect 821 519 855 553
rect 821 451 855 485
rect 977 701 1011 735
rect 977 633 1011 667
rect 977 519 1011 553
rect 977 451 1011 485
rect 1133 701 1167 735
rect 1133 633 1167 667
rect 1133 519 1167 553
rect 1133 451 1167 485
rect 1289 701 1323 735
rect 1289 633 1323 667
rect 1289 519 1323 553
rect 1289 451 1323 485
rect 1445 701 1479 735
rect 1445 633 1479 667
rect 1445 519 1479 553
rect 1445 451 1479 485
rect 1601 701 1635 735
rect 1601 633 1635 667
rect 1601 519 1635 553
rect 1601 451 1635 485
rect 1757 701 1791 735
rect 1757 633 1791 667
rect 1757 519 1791 553
rect 1757 451 1791 485
rect 1913 701 1947 735
rect 1913 633 1947 667
rect 1913 519 1947 553
rect 1913 451 1947 485
rect 2069 701 2103 735
rect 2069 633 2103 667
rect 2069 519 2103 553
rect 2069 451 2103 485
rect 2225 701 2259 735
rect 2225 633 2259 667
rect 2225 519 2259 553
rect 2225 451 2259 485
rect 2381 701 2415 735
rect 2381 633 2415 667
rect 2381 519 2415 553
rect 2381 451 2415 485
rect 2537 697 2571 731
rect 2537 629 2571 663
rect 2537 523 2571 557
rect 2537 455 2571 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2688 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
<< poly >>
rect 86 743 186 769
rect 242 743 342 769
rect 398 743 498 769
rect 554 743 654 769
rect 710 743 810 769
rect 866 743 966 769
rect 1022 743 1122 769
rect 1178 743 1278 769
rect 1334 743 1434 769
rect 1490 743 1590 769
rect 1646 743 1746 769
rect 1802 743 1902 769
rect 1958 743 2058 769
rect 2114 743 2214 769
rect 2270 743 2370 769
rect 2426 743 2526 769
rect 86 401 186 443
rect 242 401 342 443
rect 398 401 498 443
rect 554 401 654 443
rect 710 401 810 443
rect 866 401 966 443
rect 1022 401 1122 443
rect 1178 401 1278 443
rect 1334 401 1434 443
rect 1490 401 1590 443
rect 1646 401 1746 443
rect 1802 401 1902 443
rect 1958 401 2058 443
rect 2114 401 2214 443
rect 2270 401 2370 443
rect 2426 401 2526 443
rect 85 400 2526 401
rect 85 363 2525 400
rect 85 329 296 363
rect 330 329 409 363
rect 443 329 608 363
rect 642 329 721 363
rect 755 329 920 363
rect 954 329 1033 363
rect 1067 329 1232 363
rect 1266 329 1345 363
rect 1379 329 1544 363
rect 1578 329 1657 363
rect 1691 329 1856 363
rect 1890 329 1969 363
rect 2003 329 2168 363
rect 2202 329 2281 363
rect 2315 329 2525 363
rect 85 313 2525 329
rect 85 291 185 313
rect 241 291 341 313
rect 397 291 497 313
rect 553 291 653 313
rect 709 291 809 313
rect 865 291 965 313
rect 1021 291 1121 313
rect 1177 291 1277 313
rect 1333 291 1433 313
rect 1489 291 1589 313
rect 1645 291 1745 313
rect 1801 291 1901 313
rect 1957 291 2057 313
rect 2113 291 2213 313
rect 2269 291 2369 313
rect 2425 291 2525 313
rect 85 115 185 141
rect 241 115 341 141
rect 397 115 497 141
rect 553 115 653 141
rect 709 115 809 141
rect 865 115 965 141
rect 1021 115 1121 141
rect 1177 115 1277 141
rect 1333 115 1433 141
rect 1489 115 1589 141
rect 1645 115 1745 141
rect 1801 115 1901 141
rect 1957 115 2057 141
rect 2113 115 2213 141
rect 2269 115 2369 141
rect 2425 115 2525 141
<< polycont >>
rect 296 329 330 363
rect 409 329 443 363
rect 608 329 642 363
rect 721 329 755 363
rect 920 329 954 363
rect 1033 329 1067 363
rect 1232 329 1266 363
rect 1345 329 1379 363
rect 1544 329 1578 363
rect 1657 329 1691 363
rect 1856 329 1890 363
rect 1969 329 2003 363
rect 2168 329 2202 363
rect 2281 329 2315 363
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2688 831
rect 25 731 131 751
rect 25 729 41 731
rect 75 729 131 731
rect 75 697 97 729
rect 59 695 97 697
rect 25 663 131 695
rect 25 629 41 663
rect 75 629 131 663
rect 25 557 131 629
rect 25 523 41 557
rect 75 523 131 557
rect 25 489 131 523
rect 25 455 41 489
rect 75 455 131 489
rect 25 435 131 455
rect 180 735 246 751
rect 180 701 197 735
rect 231 701 246 735
rect 180 667 246 701
rect 180 633 197 667
rect 231 633 246 667
rect 180 553 246 633
rect 180 519 197 553
rect 231 519 246 553
rect 180 498 246 519
rect 180 451 197 498
rect 231 451 246 498
rect 19 279 126 295
rect 19 245 40 279
rect 74 245 126 279
rect 19 206 126 245
rect 19 172 40 206
rect 74 172 126 206
rect 19 119 126 172
rect 180 283 246 451
rect 280 735 458 751
rect 280 729 353 735
rect 387 729 458 735
rect 314 695 352 729
rect 387 701 424 729
rect 386 695 424 701
rect 280 667 458 695
rect 280 633 353 667
rect 387 633 458 667
rect 280 553 458 633
rect 280 519 353 553
rect 387 519 458 553
rect 280 485 458 519
rect 280 451 353 485
rect 387 451 458 485
rect 280 435 458 451
rect 492 735 558 751
rect 492 701 509 735
rect 543 701 558 735
rect 492 667 558 701
rect 492 633 509 667
rect 543 633 558 667
rect 492 553 558 633
rect 492 519 509 553
rect 543 519 558 553
rect 492 498 558 519
rect 492 451 509 498
rect 543 451 558 498
rect 280 363 458 379
rect 280 329 296 363
rect 330 350 409 363
rect 280 316 319 329
rect 353 316 391 350
rect 443 329 458 363
rect 425 316 458 329
rect 280 313 458 316
rect 180 249 196 283
rect 230 249 246 283
rect 492 283 558 451
rect 592 735 770 751
rect 592 729 665 735
rect 699 729 770 735
rect 626 695 664 729
rect 699 701 736 729
rect 698 695 736 701
rect 592 667 770 695
rect 592 633 665 667
rect 699 633 770 667
rect 592 553 770 633
rect 592 519 665 553
rect 699 519 770 553
rect 592 485 770 519
rect 592 451 665 485
rect 699 451 770 485
rect 592 435 770 451
rect 804 735 870 751
rect 804 701 821 735
rect 855 701 870 735
rect 804 667 870 701
rect 804 633 821 667
rect 855 633 870 667
rect 804 553 870 633
rect 804 519 821 553
rect 855 519 870 553
rect 804 498 870 519
rect 804 451 821 498
rect 855 451 870 498
rect 592 363 770 379
rect 592 329 608 363
rect 642 350 721 363
rect 592 316 629 329
rect 663 316 701 350
rect 755 329 770 363
rect 735 316 770 329
rect 592 313 770 316
rect 180 209 246 249
rect 180 175 196 209
rect 230 175 246 209
rect 180 159 246 175
rect 280 245 352 279
rect 386 245 458 279
rect 280 206 458 245
rect 280 172 352 206
rect 386 172 458 206
rect 53 85 91 119
rect 125 85 126 119
rect 19 75 126 85
rect 280 119 458 172
rect 492 249 508 283
rect 542 249 558 283
rect 804 283 870 451
rect 904 735 1082 751
rect 904 729 977 735
rect 1011 729 1082 735
rect 938 695 976 729
rect 1011 701 1048 729
rect 1010 695 1048 701
rect 904 667 1082 695
rect 904 633 977 667
rect 1011 633 1082 667
rect 904 553 1082 633
rect 904 519 977 553
rect 1011 519 1082 553
rect 904 485 1082 519
rect 904 451 977 485
rect 1011 451 1082 485
rect 904 435 1082 451
rect 1116 735 1182 751
rect 1116 701 1133 735
rect 1167 701 1182 735
rect 1116 667 1182 701
rect 1116 633 1133 667
rect 1167 633 1182 667
rect 1116 553 1182 633
rect 1116 519 1133 553
rect 1167 519 1182 553
rect 1116 498 1182 519
rect 1116 451 1133 498
rect 1167 451 1182 498
rect 904 363 1082 379
rect 904 329 920 363
rect 954 350 1033 363
rect 904 316 941 329
rect 975 316 1013 350
rect 1067 329 1082 363
rect 1047 316 1082 329
rect 904 313 1082 316
rect 492 209 558 249
rect 492 175 508 209
rect 542 175 558 209
rect 492 159 558 175
rect 592 245 664 279
rect 698 245 770 279
rect 592 206 770 245
rect 592 172 664 206
rect 698 172 770 206
rect 314 85 352 119
rect 386 85 424 119
rect 280 75 458 85
rect 592 119 770 172
rect 804 249 820 283
rect 854 249 870 283
rect 1116 283 1182 451
rect 1216 735 1394 751
rect 1216 729 1289 735
rect 1323 729 1394 735
rect 1250 695 1288 729
rect 1323 701 1360 729
rect 1322 695 1360 701
rect 1216 667 1394 695
rect 1216 633 1289 667
rect 1323 633 1394 667
rect 1216 553 1394 633
rect 1216 519 1289 553
rect 1323 519 1394 553
rect 1216 485 1394 519
rect 1216 451 1289 485
rect 1323 451 1394 485
rect 1216 435 1394 451
rect 1428 735 1494 751
rect 1428 701 1445 735
rect 1479 701 1494 735
rect 1428 667 1494 701
rect 1428 633 1445 667
rect 1479 633 1494 667
rect 1428 553 1494 633
rect 1428 519 1445 553
rect 1479 519 1494 553
rect 1428 498 1494 519
rect 1428 451 1445 498
rect 1479 451 1494 498
rect 1216 363 1394 379
rect 1216 329 1232 363
rect 1266 350 1345 363
rect 1216 316 1253 329
rect 1287 316 1325 350
rect 1379 329 1394 363
rect 1359 316 1394 329
rect 1216 313 1394 316
rect 804 209 870 249
rect 804 175 820 209
rect 854 175 870 209
rect 804 159 870 175
rect 904 245 976 279
rect 1010 245 1082 279
rect 904 206 1082 245
rect 904 172 976 206
rect 1010 172 1082 206
rect 626 85 664 119
rect 698 85 736 119
rect 592 75 770 85
rect 904 119 1082 172
rect 1116 249 1132 283
rect 1166 249 1182 283
rect 1428 283 1494 451
rect 1528 735 1706 751
rect 1528 729 1601 735
rect 1635 729 1706 735
rect 1562 695 1600 729
rect 1635 701 1672 729
rect 1634 695 1672 701
rect 1528 667 1706 695
rect 1528 633 1601 667
rect 1635 633 1706 667
rect 1528 553 1706 633
rect 1528 519 1601 553
rect 1635 519 1706 553
rect 1528 485 1706 519
rect 1528 451 1601 485
rect 1635 451 1706 485
rect 1528 435 1706 451
rect 1740 735 1806 751
rect 1740 701 1757 735
rect 1791 701 1806 735
rect 1740 667 1806 701
rect 1740 633 1757 667
rect 1791 633 1806 667
rect 1740 553 1806 633
rect 1740 519 1757 553
rect 1791 519 1806 553
rect 1740 498 1806 519
rect 1740 451 1757 498
rect 1791 451 1806 498
rect 1528 363 1706 379
rect 1528 329 1544 363
rect 1578 350 1657 363
rect 1528 316 1565 329
rect 1599 316 1637 350
rect 1691 329 1706 363
rect 1671 316 1706 329
rect 1528 313 1706 316
rect 1116 209 1182 249
rect 1116 175 1132 209
rect 1166 175 1182 209
rect 1116 159 1182 175
rect 1216 245 1288 279
rect 1322 245 1394 279
rect 1216 206 1394 245
rect 1216 172 1288 206
rect 1322 172 1394 206
rect 938 85 976 119
rect 1010 85 1048 119
rect 904 75 1082 85
rect 1216 119 1394 172
rect 1428 249 1444 283
rect 1478 249 1494 283
rect 1740 283 1806 451
rect 1840 735 2018 751
rect 1840 729 1913 735
rect 1947 729 2018 735
rect 1874 695 1912 729
rect 1947 701 1984 729
rect 1946 695 1984 701
rect 1840 667 2018 695
rect 1840 633 1913 667
rect 1947 633 2018 667
rect 1840 553 2018 633
rect 1840 519 1913 553
rect 1947 519 2018 553
rect 1840 485 2018 519
rect 1840 451 1913 485
rect 1947 451 2018 485
rect 1840 435 2018 451
rect 2052 735 2118 751
rect 2052 701 2069 735
rect 2103 701 2118 735
rect 2052 667 2118 701
rect 2052 633 2069 667
rect 2103 633 2118 667
rect 2052 553 2118 633
rect 2052 519 2069 553
rect 2103 519 2118 553
rect 2052 498 2118 519
rect 2052 451 2069 498
rect 2103 451 2118 498
rect 1840 363 2018 379
rect 1840 329 1856 363
rect 1890 350 1969 363
rect 1840 316 1877 329
rect 1911 316 1949 350
rect 2003 329 2018 363
rect 1983 316 2018 329
rect 1840 313 2018 316
rect 1428 209 1494 249
rect 1428 175 1444 209
rect 1478 175 1494 209
rect 1428 159 1494 175
rect 1528 245 1600 279
rect 1634 245 1706 279
rect 1528 206 1706 245
rect 1528 172 1600 206
rect 1634 172 1706 206
rect 1250 85 1288 119
rect 1322 85 1360 119
rect 1216 75 1394 85
rect 1528 119 1706 172
rect 1740 249 1756 283
rect 1790 249 1806 283
rect 2052 283 2118 451
rect 2152 735 2330 751
rect 2152 729 2225 735
rect 2259 729 2330 735
rect 2186 695 2224 729
rect 2259 701 2296 729
rect 2258 695 2296 701
rect 2152 667 2330 695
rect 2152 633 2225 667
rect 2259 633 2330 667
rect 2152 553 2330 633
rect 2152 519 2225 553
rect 2259 519 2330 553
rect 2152 485 2330 519
rect 2152 451 2225 485
rect 2259 451 2330 485
rect 2152 435 2330 451
rect 2364 735 2430 751
rect 2364 701 2381 735
rect 2415 701 2430 735
rect 2364 667 2430 701
rect 2364 633 2381 667
rect 2415 633 2430 667
rect 2364 553 2430 633
rect 2364 519 2381 553
rect 2415 519 2430 553
rect 2364 498 2430 519
rect 2364 451 2381 498
rect 2415 451 2430 498
rect 2152 363 2330 379
rect 2152 329 2168 363
rect 2202 350 2281 363
rect 2152 316 2189 329
rect 2223 316 2261 350
rect 2315 329 2330 363
rect 2295 316 2330 329
rect 2152 313 2330 316
rect 1740 209 1806 249
rect 1740 175 1756 209
rect 1790 175 1806 209
rect 1740 159 1806 175
rect 1840 245 1912 279
rect 1946 245 2018 279
rect 1840 206 2018 245
rect 1840 172 1912 206
rect 1946 172 2018 206
rect 1562 85 1600 119
rect 1634 85 1672 119
rect 1528 75 1706 85
rect 1840 119 2018 172
rect 2052 249 2068 283
rect 2102 249 2118 283
rect 2364 283 2430 451
rect 2464 731 2587 735
rect 2464 729 2537 731
rect 2571 729 2587 731
rect 2464 695 2473 729
rect 2507 697 2537 729
rect 2507 695 2545 697
rect 2579 695 2587 729
rect 2464 663 2587 695
rect 2464 629 2537 663
rect 2571 629 2587 663
rect 2464 557 2587 629
rect 2464 523 2537 557
rect 2571 523 2587 557
rect 2464 489 2587 523
rect 2464 455 2537 489
rect 2571 455 2587 489
rect 2464 435 2587 455
rect 2052 209 2118 249
rect 2052 175 2068 209
rect 2102 175 2118 209
rect 2052 159 2118 175
rect 2152 245 2224 279
rect 2258 245 2330 279
rect 2152 206 2330 245
rect 2152 172 2224 206
rect 2258 172 2330 206
rect 1874 85 1912 119
rect 1946 85 1984 119
rect 1840 75 2018 85
rect 2152 119 2330 172
rect 2364 249 2380 283
rect 2414 249 2430 283
rect 2364 209 2430 249
rect 2364 175 2380 209
rect 2414 175 2430 209
rect 2364 159 2430 175
rect 2464 245 2536 279
rect 2570 245 2587 279
rect 2464 206 2587 245
rect 2464 172 2536 206
rect 2570 172 2587 206
rect 2186 85 2224 119
rect 2258 85 2296 119
rect 2152 75 2330 85
rect 2464 119 2587 172
rect 2464 85 2473 119
rect 2507 85 2545 119
rect 2579 85 2587 119
rect 2464 75 2587 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 25 697 41 729
rect 41 697 59 729
rect 25 695 59 697
rect 97 695 131 729
rect 197 485 231 498
rect 197 464 231 485
rect 280 695 314 729
rect 352 701 353 729
rect 353 701 386 729
rect 352 695 386 701
rect 424 695 458 729
rect 509 485 543 498
rect 509 464 543 485
rect 319 329 330 350
rect 330 329 353 350
rect 319 316 353 329
rect 391 329 409 350
rect 409 329 425 350
rect 391 316 425 329
rect 592 695 626 729
rect 664 701 665 729
rect 665 701 698 729
rect 664 695 698 701
rect 736 695 770 729
rect 821 485 855 498
rect 821 464 855 485
rect 629 329 642 350
rect 642 329 663 350
rect 629 316 663 329
rect 701 329 721 350
rect 721 329 735 350
rect 701 316 735 329
rect 19 85 53 119
rect 91 85 125 119
rect 904 695 938 729
rect 976 701 977 729
rect 977 701 1010 729
rect 976 695 1010 701
rect 1048 695 1082 729
rect 1133 485 1167 498
rect 1133 464 1167 485
rect 941 329 954 350
rect 954 329 975 350
rect 941 316 975 329
rect 1013 329 1033 350
rect 1033 329 1047 350
rect 1013 316 1047 329
rect 280 85 314 119
rect 352 85 386 119
rect 424 85 458 119
rect 1216 695 1250 729
rect 1288 701 1289 729
rect 1289 701 1322 729
rect 1288 695 1322 701
rect 1360 695 1394 729
rect 1445 485 1479 498
rect 1445 464 1479 485
rect 1253 329 1266 350
rect 1266 329 1287 350
rect 1253 316 1287 329
rect 1325 329 1345 350
rect 1345 329 1359 350
rect 1325 316 1359 329
rect 592 85 626 119
rect 664 85 698 119
rect 736 85 770 119
rect 1528 695 1562 729
rect 1600 701 1601 729
rect 1601 701 1634 729
rect 1600 695 1634 701
rect 1672 695 1706 729
rect 1757 485 1791 498
rect 1757 464 1791 485
rect 1565 329 1578 350
rect 1578 329 1599 350
rect 1565 316 1599 329
rect 1637 329 1657 350
rect 1657 329 1671 350
rect 1637 316 1671 329
rect 904 85 938 119
rect 976 85 1010 119
rect 1048 85 1082 119
rect 1840 695 1874 729
rect 1912 701 1913 729
rect 1913 701 1946 729
rect 1912 695 1946 701
rect 1984 695 2018 729
rect 2069 485 2103 498
rect 2069 464 2103 485
rect 1877 329 1890 350
rect 1890 329 1911 350
rect 1877 316 1911 329
rect 1949 329 1969 350
rect 1969 329 1983 350
rect 1949 316 1983 329
rect 1216 85 1250 119
rect 1288 85 1322 119
rect 1360 85 1394 119
rect 2152 695 2186 729
rect 2224 701 2225 729
rect 2225 701 2258 729
rect 2224 695 2258 701
rect 2296 695 2330 729
rect 2381 485 2415 498
rect 2381 464 2415 485
rect 2189 329 2202 350
rect 2202 329 2223 350
rect 2189 316 2223 329
rect 2261 329 2281 350
rect 2281 329 2295 350
rect 2261 316 2295 329
rect 1528 85 1562 119
rect 1600 85 1634 119
rect 1672 85 1706 119
rect 2473 695 2507 729
rect 2545 697 2571 729
rect 2571 697 2579 729
rect 2545 695 2579 697
rect 1840 85 1874 119
rect 1912 85 1946 119
rect 1984 85 2018 119
rect 2152 85 2186 119
rect 2224 85 2258 119
rect 2296 85 2330 119
rect 2473 85 2507 119
rect 2545 85 2579 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
<< metal1 >>
rect 0 831 2688 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2688 831
rect 0 791 2688 797
rect 0 729 2688 763
rect 0 695 25 729
rect 59 695 97 729
rect 131 695 280 729
rect 314 695 352 729
rect 386 695 424 729
rect 458 695 592 729
rect 626 695 664 729
rect 698 695 736 729
rect 770 695 904 729
rect 938 695 976 729
rect 1010 695 1048 729
rect 1082 695 1216 729
rect 1250 695 1288 729
rect 1322 695 1360 729
rect 1394 695 1528 729
rect 1562 695 1600 729
rect 1634 695 1672 729
rect 1706 695 1840 729
rect 1874 695 1912 729
rect 1946 695 1984 729
rect 2018 695 2152 729
rect 2186 695 2224 729
rect 2258 695 2296 729
rect 2330 695 2473 729
rect 2507 695 2545 729
rect 2579 695 2688 729
rect 0 689 2688 695
rect 185 498 243 504
rect 497 498 555 504
rect 809 498 867 504
rect 1121 498 1179 504
rect 1433 498 1491 504
rect 1745 498 1803 504
rect 2057 498 2115 504
rect 2369 498 2427 504
rect 185 464 197 498
rect 231 464 509 498
rect 543 464 821 498
rect 855 464 1133 498
rect 1167 464 1445 498
rect 1479 464 1757 498
rect 1791 464 2069 498
rect 2103 464 2381 498
rect 2415 464 2427 498
rect 185 458 243 464
rect 497 458 555 464
rect 809 458 867 464
rect 1121 458 1179 464
rect 1433 458 1491 464
rect 1745 458 1803 464
rect 2057 458 2115 464
rect 2369 458 2427 464
rect 307 350 437 356
rect 617 350 747 356
rect 929 350 1059 356
rect 1241 350 1371 356
rect 1553 350 1683 356
rect 1865 350 1995 356
rect 2177 350 2307 356
rect 307 316 319 350
rect 353 316 391 350
rect 425 316 629 350
rect 663 316 701 350
rect 735 316 941 350
rect 975 316 1013 350
rect 1047 316 1253 350
rect 1287 316 1325 350
rect 1359 316 1565 350
rect 1599 316 1637 350
rect 1671 316 1877 350
rect 1911 316 1949 350
rect 1983 316 2189 350
rect 2223 316 2261 350
rect 2295 316 2307 350
rect 307 310 437 316
rect 617 310 747 316
rect 929 310 1059 316
rect 1241 310 1371 316
rect 1553 310 1683 316
rect 1865 310 1995 316
rect 2177 310 2307 316
rect 0 119 2688 125
rect 0 85 19 119
rect 53 85 91 119
rect 125 85 280 119
rect 314 85 352 119
rect 386 85 424 119
rect 458 85 592 119
rect 626 85 664 119
rect 698 85 736 119
rect 770 85 904 119
rect 938 85 976 119
rect 1010 85 1048 119
rect 1082 85 1216 119
rect 1250 85 1288 119
rect 1322 85 1360 119
rect 1394 85 1528 119
rect 1562 85 1600 119
rect 1634 85 1672 119
rect 1706 85 1840 119
rect 1874 85 1912 119
rect 1946 85 1984 119
rect 2018 85 2152 119
rect 2186 85 2224 119
rect 2258 85 2296 119
rect 2330 85 2473 119
rect 2507 85 2545 119
rect 2579 85 2688 119
rect 0 51 2688 85
rect 0 17 2688 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2688 17
rect 0 -23 2688 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_16
flabel metal1 s 185 464 2427 498 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel metal1 s 307 316 2307 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 0 0 2688 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 2688 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 2688 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 1344 802 1344 802 0 FreeSans 340 0 0 0 VPB
flabel metal1 s 0 51 2688 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 1344 11 1344 11 0 FreeSans 340 0 0 0 VNB
<< properties >>
string FIXED_BBOX 0 0 2688 814
string GDS_END 42530
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 12890
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
