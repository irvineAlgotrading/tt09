magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 250
rect 61 0 64 250
<< via1 >>
rect 3 0 61 250
<< metal2 >>
rect 0 0 3 250
rect 61 0 64 250
<< properties >>
string GDS_END 94935030
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94933874
<< end >>
