magic
tech sky130A
magscale 1 2
timestamp 1715166193
<< obsli1 >>
rect 1830 39689 14025 39939
rect 1830 34194 2080 39689
rect 2220 39367 13631 39545
rect 2220 34205 2398 39367
rect 2877 37032 3087 39037
rect 3121 36998 3339 39115
rect 3513 36998 3735 39115
rect 3797 37103 3975 39015
rect 4041 36998 4259 39115
rect 4433 36998 4655 39115
rect 4717 37103 4895 39006
rect 4961 36998 5179 39115
rect 5353 36998 5575 39115
rect 5637 37103 5815 39006
rect 5881 36998 6099 39115
rect 6273 36998 6495 39115
rect 6557 37103 6735 39006
rect 6801 36998 7019 39115
rect 7193 36998 7415 39115
rect 7477 37103 7655 39006
rect 7721 36998 7939 39115
rect 8113 36998 8335 39115
rect 8397 37103 8575 39006
rect 8641 36998 8859 39115
rect 9033 36998 9255 39115
rect 9317 37103 9495 39006
rect 9561 36998 9779 39115
rect 9953 36998 10175 39115
rect 10237 37103 10415 39006
rect 10481 36998 10699 39115
rect 10873 36998 11095 39115
rect 11157 37103 11335 39028
rect 11401 36998 11619 39115
rect 11793 36998 12015 39115
rect 12077 37103 12255 39028
rect 12321 36998 12539 39115
rect 12713 36998 12935 39115
rect 12969 37032 13175 39036
rect 2566 36514 13337 36998
rect 3121 36468 13337 36514
rect 1834 34144 2072 34194
rect 1702 26908 2072 34144
rect 2225 34103 2395 34205
rect 2154 27233 2395 34103
rect 2877 32432 3083 36386
rect 3121 32398 3339 36468
rect 3513 32398 3735 36468
rect 3797 32503 3975 36362
rect 4041 32398 4259 36468
rect 4433 32398 4655 36468
rect 4717 32503 4895 36353
rect 4961 32398 5179 36468
rect 5353 32398 5575 36468
rect 5637 32503 5815 36353
rect 5881 32398 6099 36468
rect 6273 32398 6495 36468
rect 6557 32503 6735 36353
rect 6801 32398 7019 36468
rect 7193 32398 7415 36468
rect 7477 32503 7655 36353
rect 7721 32398 7939 36468
rect 8113 32398 8335 36468
rect 8397 32503 8575 36353
rect 8641 32398 8859 36468
rect 9033 32398 9255 36468
rect 9317 32503 9495 36353
rect 9561 32398 9779 36468
rect 9953 32398 10175 36468
rect 10237 32503 10415 36353
rect 10481 32398 10699 36468
rect 10873 32398 11095 36468
rect 11157 32503 11335 36353
rect 11401 32398 11619 36468
rect 11793 32398 12015 36468
rect 12077 32503 12255 36353
rect 12321 32398 12539 36468
rect 12713 32398 12935 36468
rect 12969 32432 13175 36386
rect 13453 33198 13631 39367
rect 13458 33118 13628 33198
rect 2480 31911 12935 32398
rect 3121 31868 12935 31911
rect 2877 27832 3083 31786
rect 3121 27798 3339 31868
rect 3513 27798 3735 31868
rect 3797 27903 3975 31762
rect 4041 27798 4259 31868
rect 4433 27798 4655 31868
rect 4717 27903 4895 31753
rect 4961 27798 5179 31868
rect 5353 27798 5575 31868
rect 5637 27903 5815 31753
rect 5881 27798 6099 31868
rect 6273 27798 6495 31868
rect 6557 27903 6735 31753
rect 6801 27798 7019 31868
rect 7193 27798 7415 31868
rect 7477 27903 7655 31753
rect 7721 27798 7939 31868
rect 8113 27798 8335 31868
rect 8397 27903 8575 31753
rect 8641 27798 8859 31868
rect 9033 27798 9255 31868
rect 9317 27903 9495 31753
rect 9561 27798 9779 31868
rect 9953 27798 10175 31868
rect 10237 27903 10415 31753
rect 10481 27798 10699 31868
rect 10873 27798 11095 31868
rect 11157 27903 11335 31753
rect 11401 27798 11619 31868
rect 11793 27798 12015 31868
rect 12077 27903 12255 31753
rect 12321 27798 12539 31868
rect 12713 27798 12935 31868
rect 12969 27832 13175 31786
rect 3121 27308 12935 27798
rect 4961 27268 12935 27308
rect 2154 27105 4532 27233
rect 2225 27063 4532 27105
rect 1702 26670 4198 26908
rect 1702 26645 2738 26670
rect 3567 26629 4198 26670
rect 3913 19500 4198 26629
rect 3960 19379 4198 19500
rect 4362 19490 4532 27063
rect 4717 23232 4923 27186
rect 4961 23198 5179 27268
rect 5353 23198 5575 27268
rect 5637 23303 5815 27162
rect 5881 23198 6099 27268
rect 6273 23198 6495 27268
rect 6557 23303 6735 27153
rect 6801 23198 7019 27268
rect 7193 23198 7415 27268
rect 7477 23303 7655 27153
rect 7721 23198 7939 27268
rect 8113 23198 8335 27268
rect 8397 23303 8575 27153
rect 8641 23198 8859 27268
rect 9033 23198 9255 27268
rect 9317 23303 9495 27153
rect 9561 23198 9779 27268
rect 9953 23198 10175 27268
rect 10237 23303 10415 27153
rect 10481 23198 10699 27268
rect 10873 23198 11095 27268
rect 11157 23303 11335 27153
rect 11401 23198 11619 27268
rect 11793 23198 12015 27268
rect 12077 23303 12255 27153
rect 12321 23198 12539 27268
rect 12713 23198 12935 27268
rect 12969 26628 13175 27186
rect 12997 23790 13175 26628
rect 12969 23232 13175 23790
rect 4611 22668 12935 23198
rect 1861 14751 1997 14960
rect 3678 14745 3800 14918
rect 3960 14564 4217 19379
rect 1827 14314 4217 14564
rect 1827 8951 2077 14314
rect 4358 14173 4536 19490
rect 4717 18632 4923 22586
rect 4961 18598 5179 22668
rect 5353 18598 5575 22668
rect 5637 18703 5815 22571
rect 5881 18598 6099 22668
rect 6273 18598 6495 22668
rect 6557 18703 6735 22562
rect 6801 18598 7019 22668
rect 7193 18598 7415 22668
rect 7477 18703 7655 22562
rect 7721 18598 7939 22668
rect 8113 18598 8335 22668
rect 8397 18703 8575 22562
rect 8641 18598 8859 22668
rect 9033 18598 9255 22668
rect 9317 18703 9495 22562
rect 9561 18598 9779 22668
rect 9953 18598 10175 22668
rect 10237 18703 10415 22562
rect 10481 18598 10699 22668
rect 10873 18598 11095 22668
rect 11157 18703 11335 22562
rect 11401 18598 11619 22668
rect 11793 18598 12015 22668
rect 12077 18703 12255 22562
rect 12321 18598 12539 22668
rect 12713 18598 12935 22668
rect 12969 22029 13175 22587
rect 12997 19190 13175 22029
rect 13458 20342 13631 33118
rect 13458 20263 13628 20342
rect 12969 18632 13175 19190
rect 4605 18099 12935 18598
rect 4961 18068 12935 18099
rect 2221 13995 4536 14173
rect 4717 14032 4923 17986
rect 4961 13998 5179 18068
rect 5353 13998 5575 18068
rect 5637 14103 5815 17962
rect 5881 13998 6099 18068
rect 6273 13998 6495 18068
rect 6557 14103 6735 17953
rect 6801 13998 7019 18068
rect 7193 13998 7415 18068
rect 7477 14103 7655 17953
rect 7721 13998 7939 18068
rect 8113 13998 8335 18068
rect 8397 14103 8575 17953
rect 8641 13998 8859 18068
rect 9033 13998 9255 18068
rect 9317 14103 9495 17953
rect 9561 13998 9779 18068
rect 9953 13998 10175 18068
rect 10237 14103 10415 17953
rect 10481 13998 10699 18068
rect 10873 13998 11095 18068
rect 11157 14103 11335 17953
rect 11401 13998 11619 18068
rect 11793 13998 12015 18068
rect 12077 14103 12255 17953
rect 12321 13998 12539 18068
rect 12713 13998 12935 18068
rect 12969 17428 13175 17986
rect 12997 14590 13175 17428
rect 12969 14032 13175 14590
rect 2221 9270 2399 13995
rect 4702 13799 12935 13998
rect 2617 9398 2651 13593
rect 3121 13468 12935 13799
rect 2877 9432 3083 13386
rect 3121 9398 3339 13468
rect 3513 9398 3735 13468
rect 3797 9503 3975 13371
rect 4041 9398 4259 13468
rect 4433 9398 4655 13468
rect 4717 9503 4895 13362
rect 4961 9398 5179 13468
rect 5353 9398 5575 13468
rect 5637 9503 5815 13362
rect 5881 9398 6099 13468
rect 6273 9398 6495 13468
rect 6557 9503 6735 13362
rect 6801 9398 7019 13468
rect 7193 9398 7415 13468
rect 7477 9503 7655 13362
rect 7721 9398 7939 13468
rect 8113 9398 8335 13468
rect 8397 9503 8575 13362
rect 8641 9398 8859 13468
rect 9033 9398 9255 13468
rect 9317 9503 9495 13362
rect 9561 9398 9779 13468
rect 9953 9398 10175 13468
rect 10237 9503 10415 13362
rect 10481 9398 10699 13468
rect 10873 9398 11095 13468
rect 11157 9503 11335 13362
rect 11401 9398 11619 13468
rect 11793 9398 12015 13468
rect 12077 9503 12255 13362
rect 12321 9398 12539 13468
rect 12713 9398 12935 13468
rect 12969 9432 13175 13386
rect 2617 9363 12935 9398
rect 2618 9348 12935 9363
rect 13453 9270 13631 20263
rect 2221 9092 13631 9270
rect 13775 9237 14025 39689
rect 14449 39606 14555 39767
rect 13781 9199 14019 9237
rect 13775 8951 14025 9199
rect 214 8554 338 8720
rect 1591 8568 1743 8724
rect 1827 8701 14025 8951
rect 620 7683 10264 8533
rect 10473 8499 14019 8701
rect 620 5684 940 7683
rect 1107 7485 9191 7519
rect 1107 5886 1141 7485
rect 1268 7394 9012 7446
rect 1223 6668 1257 7298
rect 1535 6667 1569 7298
rect 1847 6668 1881 7298
rect 2159 6667 2193 7298
rect 2471 6668 2505 7298
rect 2783 6667 2817 7298
rect 3095 6668 3129 7298
rect 3407 6667 3441 7298
rect 3719 6668 3753 7298
rect 4031 6667 4065 7298
rect 4343 6668 4377 7298
rect 4655 6667 4689 7298
rect 4967 6668 5001 7298
rect 5279 6667 5313 7298
rect 5591 6668 5625 7298
rect 5903 6667 5937 7298
rect 6215 6668 6249 7298
rect 6527 6667 6561 7298
rect 6839 6668 6873 7298
rect 7151 6667 7185 7298
rect 7463 6668 7497 7298
rect 7775 6667 7809 7298
rect 8087 6667 8121 7298
rect 8399 6668 8433 7298
rect 8711 6667 8745 7298
rect 9023 6668 9057 7298
rect 1379 5955 1413 6572
rect 1691 5954 1725 6572
rect 2003 5955 2037 6572
rect 2315 5954 2349 6572
rect 2627 5955 2661 6572
rect 2939 5954 2973 6572
rect 3251 5954 3285 6572
rect 3563 5954 3597 6572
rect 3875 5955 3909 6572
rect 4187 5954 4221 6572
rect 4499 5955 4533 6572
rect 4811 5954 4845 6572
rect 5123 5955 5157 6572
rect 5435 5954 5469 6572
rect 5747 5955 5781 6572
rect 6059 5954 6093 6572
rect 6371 5955 6405 6572
rect 6683 5954 6717 6572
rect 6995 5955 7029 6572
rect 7307 5954 7341 6572
rect 7619 5955 7653 6572
rect 7931 5954 7965 6572
rect 8243 5954 8277 6572
rect 8555 5955 8589 6572
rect 8867 5954 8901 6572
rect 9151 5886 9191 7485
rect 1107 5846 9191 5886
rect 9354 5684 10264 7683
rect 620 4784 10264 5684
rect 10464 8291 14019 8499
rect 10464 6212 10642 8291
rect 13595 8263 14019 8291
rect 14106 8284 14229 8425
rect 10792 8082 13428 8116
rect 10792 6401 10826 8082
rect 10988 7954 13267 7988
rect 10939 7238 10973 7858
rect 11251 7238 11285 7858
rect 11563 7238 11597 7858
rect 11875 7238 11909 7858
rect 12187 7238 12221 7858
rect 12499 7238 12533 7858
rect 12811 7238 12845 7858
rect 13123 7238 13157 7858
rect 13387 7255 13428 8082
rect 13394 7213 13428 7255
rect 11093 6524 11127 7154
rect 11405 6524 11439 7154
rect 11717 6524 11751 7154
rect 12029 6524 12063 7154
rect 12341 6524 12375 7154
rect 12653 6524 12687 7154
rect 12965 6524 12999 7154
rect 13277 6524 13311 7154
rect 13387 6401 13428 7213
rect 10792 6367 13428 6401
rect 13600 6212 14019 8263
rect 10464 5865 14019 6212
rect 10464 5687 14126 5865
rect 620 213 2126 4784
rect 10464 4648 11199 5687
rect 11364 5497 12562 5543
rect 11364 4696 11410 5497
rect 11511 4696 11557 5286
rect 12370 4696 12416 5286
rect 12516 4696 12562 5497
rect 2330 4446 11199 4648
rect 2330 378 2508 4446
rect 10643 4445 11199 4446
rect 11370 4293 11404 4696
rect 11563 4347 12363 4393
rect 12522 4293 12556 4696
rect 13948 4504 14126 5687
rect 13956 4464 14126 4504
rect 13948 378 14126 4464
rect 2330 200 14126 378
<< metal1 >>
rect 621 7770 10263 8496
rect 621 7763 1123 7770
rect 9215 7769 10263 7770
rect 621 7749 1109 7763
rect 9229 7755 10263 7769
rect 621 7742 1095 7749
rect 621 7609 969 7742
rect 9243 7741 10263 7755
rect 9257 7727 10263 7741
rect 9271 7713 10263 7727
rect 9285 7699 10263 7713
rect 9299 7685 10263 7699
rect 9313 7671 10263 7685
rect 9327 7657 10263 7671
rect 9341 7643 10263 7657
rect 9355 7629 10263 7643
rect 9369 7615 10263 7629
rect 621 7595 955 7609
rect 9383 7601 10263 7615
rect 621 5831 941 7595
rect 9397 7587 10263 7601
rect 9411 7573 10263 7587
rect 9425 7559 10263 7573
rect 9439 7558 10263 7559
rect 9481 7503 10263 7558
rect 9495 7489 10263 7503
rect 9509 7475 10263 7489
rect 9523 7461 10263 7475
rect 9537 5826 10263 7461
rect 9523 5812 10263 5826
rect 9509 5798 10263 5812
rect 9495 5784 10263 5798
rect 9481 5770 10263 5784
rect 9467 5756 10263 5770
rect 9460 5546 10263 5756
rect 9243 5532 10263 5546
rect 9229 5518 10263 5532
rect 620 4792 10263 5518
rect 620 4781 2366 4792
rect 620 4767 2352 4781
rect 620 4764 2338 4767
rect 620 4109 1694 4764
rect 620 4095 1680 4109
rect 620 2 1666 4095
<< obsm1 >>
rect 0 8524 15000 40000
rect 0 5803 593 8524
rect 969 7698 9202 7742
rect 969 7684 9207 7698
rect 969 7670 9221 7684
rect 969 7656 9235 7670
rect 969 7642 9249 7656
rect 969 7628 9263 7642
rect 969 7614 9277 7628
rect 969 7600 9291 7614
rect 969 7586 9305 7600
rect 969 7572 9319 7586
rect 969 7569 9333 7572
rect 969 7558 9375 7569
rect 969 7435 9481 7558
rect 969 5803 9509 7435
rect 0 5775 9481 5803
rect 0 5546 9460 5775
rect 0 0 592 5546
rect 10291 4764 15000 8524
rect 1694 0 15000 4764
<< metal2 >>
rect 187 38112 13440 39015
rect 187 38099 3006 38112
rect 187 38085 2992 38099
rect 187 38071 2978 38085
rect 187 38057 2964 38071
rect 187 38043 2950 38057
rect 187 38031 2936 38043
rect 187 37973 2880 38031
rect 187 37959 2866 37973
rect 187 37945 2852 37959
rect 187 37931 2838 37945
rect 187 37005 2824 37931
rect 3361 37059 14858 38003
rect 11746 37052 14858 37059
rect 11760 37038 14858 37052
rect 11774 37024 14858 37038
rect 187 36991 2830 37005
rect 11788 37010 14858 37024
rect 11802 36996 14858 37010
rect 187 36977 2844 36991
rect 11816 36982 14858 36996
rect 187 36963 2858 36977
rect 11830 36968 14858 36982
rect 187 36949 2872 36963
rect 11844 36954 14858 36968
rect 187 36935 2886 36949
rect 11858 36940 14858 36954
rect 187 36921 2900 36935
rect 11872 36926 14858 36940
rect 187 36907 2914 36921
rect 11886 36912 14858 36926
rect 187 36893 2928 36907
rect 11900 36898 14858 36912
rect 187 36879 2942 36893
rect 11914 36884 14858 36898
rect 187 36865 2956 36879
rect 11928 36870 14858 36884
rect 187 36851 2970 36865
rect 11942 36856 14858 36870
rect 187 36837 2984 36851
rect 11956 36842 14858 36856
rect 187 36823 2998 36837
rect 187 36809 3012 36823
rect 187 36795 3026 36809
rect 187 36781 3040 36795
rect 11970 36828 14858 36842
rect 11984 36814 14858 36828
rect 11998 36800 14858 36814
rect 187 36758 3064 36781
rect 12012 36786 14858 36800
rect 12026 36772 14858 36786
rect 187 36744 3077 36758
rect 12040 36758 14858 36772
rect 187 36730 3091 36744
rect 12054 36744 14858 36758
rect 187 36716 3105 36730
rect 12068 36730 14858 36744
rect 187 36702 3119 36716
rect 12082 36716 14858 36730
rect 187 36688 3133 36702
rect 12096 36702 14858 36716
rect 187 36674 3147 36688
rect 12110 36688 14858 36702
rect 187 36660 3161 36674
rect 12124 36674 14858 36688
rect 187 36646 3175 36660
rect 12138 36660 14858 36674
rect 187 36632 3189 36646
rect 12152 36646 14858 36660
rect 187 36618 3203 36632
rect 12166 36632 14858 36646
rect 187 36604 3217 36618
rect 12180 36618 14858 36632
rect 187 36590 3231 36604
rect 12194 36604 14858 36618
rect 187 36576 3245 36590
rect 12208 36590 14858 36604
rect 187 36562 3259 36576
rect 187 36548 3273 36562
rect 187 36534 3287 36548
rect 187 36520 3301 36534
rect 187 36506 3315 36520
rect 187 36492 3329 36506
rect 187 36478 3343 36492
rect 187 36464 3357 36478
rect 187 36450 3371 36464
rect 187 36436 3385 36450
rect 187 36422 3399 36436
rect 187 36408 3413 36422
rect 187 36394 3427 36408
rect 187 36380 3441 36394
rect 187 36366 3455 36380
rect 187 36352 3469 36366
rect 187 36338 3483 36352
rect 187 36324 3497 36338
rect 187 36310 3511 36324
rect 187 36296 3525 36310
rect 187 34556 11592 36296
rect 187 34544 3524 34556
rect 187 34530 3510 34544
rect 187 34516 3496 34530
rect 187 34502 3482 34516
rect 187 34500 3468 34502
rect 12222 34931 14858 36590
rect 12213 34917 14858 34931
rect 12199 34903 14858 34917
rect 12194 34500 14858 34903
rect 187 34348 3318 34500
rect 187 34334 3314 34348
rect 187 34320 3300 34334
rect 187 34306 3286 34320
rect 187 34292 3272 34306
rect 187 34278 3258 34292
rect 187 34264 3244 34278
rect 187 34259 3230 34264
rect 11793 34497 14858 34500
rect 11779 34483 14858 34497
rect 11765 34469 14858 34483
rect 11751 34455 14858 34469
rect 11742 34259 14858 34455
rect 187 33900 2880 34259
rect 187 33886 2866 33900
rect 187 33872 2852 33886
rect 187 33858 2838 33872
rect 187 32410 2824 33858
rect 11541 34245 14858 34259
rect 11527 34231 14858 34245
rect 3361 32491 14858 34231
rect 11508 32488 14858 32491
rect 11522 32474 14858 32488
rect 11536 32460 14858 32474
rect 11550 32446 14858 32460
rect 11564 32432 14858 32446
rect 11578 32418 14858 32432
rect 187 32396 2830 32410
rect 11592 32404 14858 32418
rect 187 32382 2844 32396
rect 11606 32390 14858 32404
rect 187 32368 2858 32382
rect 11620 32376 14858 32390
rect 187 32354 2872 32368
rect 11634 32362 14858 32376
rect 187 32340 2886 32354
rect 11648 32348 14858 32362
rect 187 32326 2900 32340
rect 11662 32334 14858 32348
rect 187 32312 2914 32326
rect 11676 32320 14858 32334
rect 187 32298 2928 32312
rect 11690 32306 14858 32320
rect 187 32284 2942 32298
rect 11704 32292 14858 32306
rect 187 32270 2956 32284
rect 11718 32278 14858 32292
rect 187 32256 2970 32270
rect 11732 32264 14858 32278
rect 187 32242 2984 32256
rect 11746 32250 14858 32264
rect 187 32228 2998 32242
rect 11760 32236 14858 32250
rect 187 32214 3012 32228
rect 11774 32222 14858 32236
rect 187 32200 3026 32214
rect 11788 32208 14858 32222
rect 187 32186 3040 32200
rect 11802 32194 14858 32208
rect 187 32172 3054 32186
rect 11816 32180 14858 32194
rect 187 32158 3068 32172
rect 11830 32166 14858 32180
rect 187 32144 3082 32158
rect 11844 32152 14858 32166
rect 187 32130 3096 32144
rect 11858 32138 14858 32152
rect 187 32116 3110 32130
rect 11872 32124 14858 32138
rect 187 32102 3124 32116
rect 11886 32110 14858 32124
rect 187 32088 3138 32102
rect 11900 32096 14858 32110
rect 187 32074 3152 32088
rect 11914 32082 14858 32096
rect 187 32060 3166 32074
rect 11928 32068 14858 32082
rect 187 32046 3180 32060
rect 11942 32054 14858 32068
rect 187 32032 3194 32046
rect 11956 32040 14858 32054
rect 187 32018 3208 32032
rect 11970 32026 14858 32040
rect 187 32004 3222 32018
rect 11984 32012 14858 32026
rect 187 31990 3236 32004
rect 11998 31998 14858 32012
rect 187 31976 3250 31990
rect 12012 31984 14858 31998
rect 187 31962 3264 31976
rect 12026 31970 14858 31984
rect 187 31948 3278 31962
rect 12040 31956 14858 31970
rect 187 31934 3292 31948
rect 12054 31942 14858 31956
rect 187 31920 3306 31934
rect 12068 31928 14858 31942
rect 187 31906 3320 31920
rect 12082 31914 14858 31928
rect 187 31892 3334 31906
rect 12096 31900 14858 31914
rect 187 31878 3348 31892
rect 12110 31886 14858 31900
rect 187 31864 3362 31878
rect 12124 31872 14858 31886
rect 187 31850 3376 31864
rect 12138 31858 14858 31872
rect 187 31836 3390 31850
rect 12152 31844 14858 31858
rect 187 31822 3404 31836
rect 12166 31830 14858 31844
rect 187 31808 3418 31822
rect 12180 31816 14858 31830
rect 187 31794 3432 31808
rect 12194 31802 14858 31816
rect 187 31780 3446 31794
rect 12208 31788 14858 31802
rect 187 31766 3460 31780
rect 187 31752 3474 31766
rect 187 31738 3488 31752
rect 187 31724 3502 31738
rect 187 31710 3516 31724
rect 187 31696 3530 31710
rect 187 29956 11341 31696
rect 187 29943 3524 29956
rect 187 29929 3510 29943
rect 187 29915 3496 29929
rect 187 29901 3482 29915
rect 187 29900 3468 29901
rect 12222 30345 14858 31788
rect 12211 30331 14858 30345
rect 12197 30317 14858 30331
rect 12194 29900 14858 30317
rect 187 29747 3319 29900
rect 187 29733 3314 29747
rect 187 29719 3300 29733
rect 187 29705 3286 29719
rect 187 29691 3272 29705
rect 187 29677 3258 29691
rect 187 29663 3244 29677
rect 187 29659 3230 29663
rect 11777 29897 14858 29900
rect 11763 29883 14858 29897
rect 11749 29869 14858 29883
rect 11735 29855 14858 29869
rect 11726 29659 14858 29855
rect 187 29439 3014 29659
rect 187 29425 3006 29439
rect 187 29411 2992 29425
rect 187 29397 2978 29411
rect 187 29383 2964 29397
rect 187 29369 2950 29383
rect 187 29355 2936 29369
rect 187 29354 2922 29355
rect 11525 29645 14858 29659
rect 11511 29631 14858 29645
rect 3650 29622 14858 29631
rect 3641 29608 14858 29622
rect 3638 29354 14858 29608
rect 187 29299 2880 29354
rect 187 29285 2866 29299
rect 187 29271 2852 29285
rect 187 29257 2838 29271
rect 187 27824 2824 29257
rect 3375 29342 14858 29354
rect 3361 27891 14858 29342
rect 11508 27885 14858 27891
rect 11522 27871 14858 27885
rect 11536 27857 14858 27871
rect 11550 27843 14858 27857
rect 11564 27829 14858 27843
rect 187 27810 2834 27824
rect 11578 27815 14858 27829
rect 187 27796 2848 27810
rect 11592 27801 14858 27815
rect 187 27782 2862 27796
rect 11606 27787 14858 27801
rect 187 27768 2876 27782
rect 11620 27773 14858 27787
rect 187 27754 2890 27768
rect 11634 27759 14858 27773
rect 187 27740 2904 27754
rect 11648 27745 14858 27759
rect 187 27726 2918 27740
rect 11662 27731 14858 27745
rect 187 27712 2932 27726
rect 11676 27717 14858 27731
rect 187 27698 2946 27712
rect 11690 27703 14858 27717
rect 187 27684 2960 27698
rect 11704 27689 14858 27703
rect 187 27670 2974 27684
rect 11718 27675 14858 27689
rect 187 27656 2988 27670
rect 11732 27661 14858 27675
rect 187 27642 3002 27656
rect 11746 27647 14858 27661
rect 187 27628 3016 27642
rect 11760 27633 14858 27647
rect 187 27614 3030 27628
rect 11774 27619 14858 27633
rect 187 27600 3044 27614
rect 11788 27605 14858 27619
rect 187 27586 3058 27600
rect 11802 27591 14858 27605
rect 187 27572 3072 27586
rect 11816 27577 14858 27591
rect 187 27558 3086 27572
rect 11830 27563 14858 27577
rect 187 27544 3100 27558
rect 11844 27549 14858 27563
rect 187 27530 3114 27544
rect 11858 27535 14858 27549
rect 187 27516 3128 27530
rect 11872 27521 14858 27535
rect 187 27502 3142 27516
rect 11886 27507 14858 27521
rect 187 27488 3156 27502
rect 11900 27493 14858 27507
rect 187 27474 3170 27488
rect 11914 27479 14858 27493
rect 187 27460 3184 27474
rect 11928 27465 14858 27479
rect 187 27446 3198 27460
rect 11942 27451 14858 27465
rect 187 27432 3212 27446
rect 11956 27437 14858 27451
rect 187 27418 3226 27432
rect 11970 27423 14858 27437
rect 187 27404 3240 27418
rect 11984 27409 14858 27423
rect 187 27390 3254 27404
rect 11998 27395 14858 27409
rect 187 27376 3268 27390
rect 12012 27381 14858 27395
rect 187 27362 3282 27376
rect 12026 27367 14858 27381
rect 187 27348 3296 27362
rect 12040 27353 14858 27367
rect 187 27334 3310 27348
rect 12054 27339 14858 27353
rect 187 27320 3324 27334
rect 12068 27325 14858 27339
rect 187 27306 3338 27320
rect 12082 27311 14858 27325
rect 187 27292 3352 27306
rect 12096 27297 14858 27311
rect 187 27278 3366 27292
rect 12110 27283 14858 27297
rect 187 27264 3380 27278
rect 12124 27269 14858 27283
rect 187 27250 3394 27264
rect 12138 27255 14858 27269
rect 187 27236 3408 27250
rect 12152 27241 14858 27255
rect 187 27222 3422 27236
rect 12166 27227 14858 27241
rect 187 27208 3436 27222
rect 12180 27213 14858 27227
rect 187 27194 3450 27208
rect 12194 27199 14858 27213
rect 187 27180 3464 27194
rect 12208 27185 14858 27199
rect 187 27166 3478 27180
rect 187 27152 3492 27166
rect 187 27138 3506 27152
rect 187 27124 3520 27138
rect 187 27110 3534 27124
rect 187 27096 3548 27110
rect 187 25356 11341 27096
rect 187 25343 3538 25356
rect 187 25329 3524 25343
rect 187 25315 3510 25329
rect 187 25301 3496 25315
rect 187 25300 3482 25301
rect 12222 25731 14858 27185
rect 12211 25717 14858 25731
rect 12197 25703 14858 25717
rect 12194 25300 14858 25703
rect 187 25147 3333 25300
rect 187 25133 3328 25147
rect 187 25119 3314 25133
rect 187 25105 3300 25119
rect 187 25091 3286 25105
rect 187 25077 3272 25091
rect 187 25063 3258 25077
rect 187 25059 3244 25063
rect 11791 25297 14858 25300
rect 11777 25283 14858 25297
rect 11763 25269 14858 25283
rect 11749 25255 14858 25269
rect 11740 25059 14858 25255
rect 187 24685 2880 25059
rect 187 24671 2866 24685
rect 187 24657 2852 24671
rect 187 24643 2838 24657
rect 187 23210 2824 24643
rect 11539 25045 14858 25059
rect 11525 25031 14858 25045
rect 4964 23291 14858 25031
rect 11508 23278 14858 23291
rect 11522 23264 14858 23278
rect 11536 23250 14858 23264
rect 11550 23236 14858 23250
rect 11564 23222 14858 23236
rect 187 23196 2827 23210
rect 11578 23208 14858 23222
rect 187 23182 2841 23196
rect 11592 23194 14858 23208
rect 187 23168 2855 23182
rect 11606 23180 14858 23194
rect 187 23154 2869 23168
rect 11620 23166 14858 23180
rect 187 23140 2883 23154
rect 11634 23152 14858 23166
rect 187 23126 2897 23140
rect 11648 23138 14858 23152
rect 187 23112 2911 23126
rect 11662 23124 14858 23138
rect 187 23098 2925 23112
rect 11676 23110 14858 23124
rect 187 23084 2939 23098
rect 11690 23096 14858 23110
rect 187 23070 2953 23084
rect 11704 23082 14858 23096
rect 187 23056 2967 23070
rect 11718 23068 14858 23082
rect 187 23042 2981 23056
rect 11732 23054 14858 23068
rect 187 23028 2995 23042
rect 11746 23040 14858 23054
rect 187 23014 3009 23028
rect 11760 23026 14858 23040
rect 187 23000 3023 23014
rect 11774 23012 14858 23026
rect 187 22986 3037 23000
rect 11788 22998 14858 23012
rect 187 22972 3051 22986
rect 11802 22984 14858 22998
rect 187 22958 3065 22972
rect 11816 22970 14858 22984
rect 187 22944 3079 22958
rect 11830 22956 14858 22970
rect 187 22930 3093 22944
rect 11844 22942 14858 22956
rect 187 22916 3107 22930
rect 11858 22928 14858 22942
rect 187 22902 3121 22916
rect 11872 22914 14858 22928
rect 187 22888 3135 22902
rect 11886 22900 14858 22914
rect 187 22874 3149 22888
rect 11900 22886 14858 22900
rect 187 22860 3163 22874
rect 11914 22872 14858 22886
rect 187 22846 3177 22860
rect 11928 22858 14858 22872
rect 187 22832 3191 22846
rect 11942 22844 14858 22858
rect 187 22818 3205 22832
rect 11956 22830 14858 22844
rect 187 22804 3219 22818
rect 11970 22816 14858 22830
rect 187 22790 3233 22804
rect 11984 22802 14858 22816
rect 187 22776 3247 22790
rect 11998 22788 14858 22802
rect 187 22762 3261 22776
rect 12012 22774 14858 22788
rect 187 22748 3275 22762
rect 12026 22760 14858 22774
rect 187 22734 3289 22748
rect 12040 22746 14858 22760
rect 187 22720 3303 22734
rect 12054 22732 14858 22746
rect 187 22706 3317 22720
rect 12068 22718 14858 22732
rect 187 22692 3331 22706
rect 12082 22704 14858 22718
rect 187 22678 3345 22692
rect 12096 22690 14858 22704
rect 187 22664 3359 22678
rect 12110 22676 14858 22690
rect 187 22650 3373 22664
rect 12124 22662 14858 22676
rect 187 22636 3387 22650
rect 12138 22648 14858 22662
rect 187 22622 3401 22636
rect 12152 22634 14858 22648
rect 187 22608 3415 22622
rect 12166 22620 14858 22634
rect 187 22594 3429 22608
rect 12180 22606 14858 22620
rect 187 22580 3443 22594
rect 12194 22592 14858 22606
rect 187 22566 3457 22580
rect 12208 22578 14858 22592
rect 187 22552 3471 22566
rect 187 22538 3485 22552
rect 187 22524 3499 22538
rect 187 22510 3513 22524
rect 187 22496 3527 22510
rect 187 20756 11341 22496
rect 187 20748 3524 20756
rect 187 20734 3510 20748
rect 187 20720 3496 20734
rect 187 20706 3482 20720
rect 187 20700 3468 20706
rect 12222 21131 14858 22578
rect 12211 21117 14858 21131
rect 12197 21103 14858 21117
rect 12194 20700 14858 21103
rect 187 20538 3314 20700
rect 187 20524 3300 20538
rect 187 20510 3286 20524
rect 187 20496 3272 20510
rect 187 20482 3258 20496
rect 187 20468 3244 20482
rect 187 20459 3230 20468
rect 11791 20697 14858 20700
rect 11777 20683 14858 20697
rect 11763 20669 14858 20683
rect 11749 20655 14858 20669
rect 11740 20459 14858 20655
rect 187 20104 2880 20459
rect 187 20090 2866 20104
rect 187 20076 2852 20090
rect 187 20062 2838 20076
rect 187 18596 2824 20062
rect 11539 20445 14858 20459
rect 11525 20431 14858 20445
rect 4964 18691 14858 20431
rect 11522 18682 14858 18691
rect 11536 18668 14858 18682
rect 11550 18654 14858 18668
rect 11564 18640 14858 18654
rect 11578 18626 14858 18640
rect 11592 18612 14858 18626
rect 187 18582 2833 18596
rect 11606 18598 14858 18612
rect 187 18568 2847 18582
rect 11620 18584 14858 18598
rect 187 18554 2861 18568
rect 11634 18570 14858 18584
rect 187 18540 2875 18554
rect 11648 18556 14858 18570
rect 187 18526 2889 18540
rect 11662 18542 14858 18556
rect 187 18512 2903 18526
rect 11676 18528 14858 18542
rect 187 18498 2917 18512
rect 11690 18514 14858 18528
rect 187 18484 2931 18498
rect 11704 18500 14858 18514
rect 187 18470 2945 18484
rect 11718 18486 14858 18500
rect 187 18456 2959 18470
rect 11732 18472 14858 18486
rect 187 18442 2973 18456
rect 11746 18458 14858 18472
rect 187 18428 2987 18442
rect 11760 18444 14858 18458
rect 187 18414 3001 18428
rect 11774 18430 14858 18444
rect 187 18400 3015 18414
rect 11788 18416 14858 18430
rect 187 18386 3029 18400
rect 11802 18402 14858 18416
rect 187 18372 3043 18386
rect 11816 18388 14858 18402
rect 187 18358 3057 18372
rect 11830 18374 14858 18388
rect 187 18344 3071 18358
rect 11844 18360 14858 18374
rect 187 18330 3085 18344
rect 11858 18346 14858 18360
rect 187 18316 3099 18330
rect 11872 18332 14858 18346
rect 187 18302 3113 18316
rect 11886 18318 14858 18332
rect 187 18288 3127 18302
rect 11900 18304 14858 18318
rect 187 18274 3141 18288
rect 11914 18290 14858 18304
rect 187 18260 3155 18274
rect 11928 18276 14858 18290
rect 187 18246 3169 18260
rect 11942 18262 14858 18276
rect 187 18232 3183 18246
rect 11956 18248 14858 18262
rect 187 18218 3197 18232
rect 11970 18234 14858 18248
rect 187 18204 3211 18218
rect 11984 18220 14858 18234
rect 187 18190 3225 18204
rect 11998 18206 14858 18220
rect 187 18176 3239 18190
rect 12012 18192 14858 18206
rect 187 18162 3253 18176
rect 12026 18178 14858 18192
rect 187 18148 3267 18162
rect 12040 18164 14858 18178
rect 187 18134 3281 18148
rect 12054 18150 14858 18164
rect 187 18120 3295 18134
rect 12068 18136 14858 18150
rect 187 18106 3309 18120
rect 12082 18122 14858 18136
rect 187 18092 3323 18106
rect 12096 18108 14858 18122
rect 187 18078 3337 18092
rect 12110 18094 14858 18108
rect 187 18064 3351 18078
rect 12124 18080 14858 18094
rect 187 18050 3365 18064
rect 12138 18066 14858 18080
rect 187 18036 3379 18050
rect 12152 18052 14858 18066
rect 187 18022 3393 18036
rect 12166 18038 14858 18052
rect 187 18008 3407 18022
rect 12180 18024 14858 18038
rect 187 17994 3421 18008
rect 12194 18010 14858 18024
rect 187 17980 3435 17994
rect 12208 17996 14858 18010
rect 187 17966 3449 17980
rect 187 17952 3463 17966
rect 187 17938 3477 17952
rect 187 17924 3491 17938
rect 187 17910 3505 17924
rect 187 17896 3519 17910
rect 187 16156 11341 17896
rect 187 16148 3524 16156
rect 187 16134 3510 16148
rect 187 16120 3496 16134
rect 187 16106 3482 16120
rect 187 16100 3468 16106
rect 12222 16531 14858 17996
rect 12211 16517 14858 16531
rect 12197 16503 14858 16517
rect 12194 16100 14858 16503
rect 187 15938 3314 16100
rect 187 15924 3300 15938
rect 187 15910 3286 15924
rect 187 15896 3272 15910
rect 187 15882 3258 15896
rect 187 15868 3244 15882
rect 187 15859 3230 15868
rect 11791 16097 14858 16100
rect 11777 16083 14858 16097
rect 11763 16069 14858 16083
rect 11749 16055 14858 16069
rect 11740 15859 14858 16055
rect 187 15504 2880 15859
rect 187 15490 2866 15504
rect 187 15476 2852 15490
rect 187 15462 2838 15476
rect 187 13996 2824 15462
rect 11539 15845 14858 15859
rect 11525 15831 14858 15845
rect 4964 15112 14858 15831
rect 4953 15098 14858 15112
rect 4939 15084 14858 15098
rect 4936 14944 14858 15084
rect 4785 14930 14858 14944
rect 4771 14916 14858 14930
rect 3682 14798 14858 14916
rect 4768 14793 14858 14798
rect 4782 14779 14858 14793
rect 4796 14765 14858 14779
rect 4810 14751 14858 14765
rect 4824 14737 14858 14751
rect 4838 14723 14858 14737
rect 4852 14709 14858 14723
rect 4866 14695 14858 14709
rect 4880 14681 14858 14695
rect 4894 14667 14858 14681
rect 4908 14653 14858 14667
rect 4922 14639 14858 14653
rect 4936 14625 14858 14639
rect 4950 14611 14858 14625
rect 4964 14091 14858 14611
rect 11508 14084 14858 14091
rect 11522 14070 14858 14084
rect 11536 14056 14858 14070
rect 11550 14042 14858 14056
rect 11564 14028 14858 14042
rect 11578 14014 14858 14028
rect 11592 14000 14858 14014
rect 187 13982 2833 13996
rect 11606 13986 14858 14000
rect 187 13968 2847 13982
rect 11620 13972 14858 13986
rect 187 13954 2861 13968
rect 11634 13958 14858 13972
rect 187 13940 2875 13954
rect 11648 13944 14858 13958
rect 187 13926 2889 13940
rect 11662 13930 14858 13944
rect 187 13912 2903 13926
rect 11676 13916 14858 13930
rect 187 13898 2917 13912
rect 11690 13902 14858 13916
rect 187 13884 2931 13898
rect 11704 13888 14858 13902
rect 187 13870 2945 13884
rect 11718 13874 14858 13888
rect 187 13856 2959 13870
rect 11732 13860 14858 13874
rect 187 13842 2973 13856
rect 11746 13846 14858 13860
rect 187 13828 2987 13842
rect 11760 13832 14858 13846
rect 187 13814 3001 13828
rect 11774 13818 14858 13832
rect 187 13800 3015 13814
rect 11788 13804 14858 13818
rect 187 13786 3029 13800
rect 11802 13790 14858 13804
rect 187 13772 3043 13786
rect 11816 13776 14858 13790
rect 187 13758 3057 13772
rect 11830 13762 14858 13776
rect 187 13744 3071 13758
rect 11844 13748 14858 13762
rect 187 13730 3085 13744
rect 11858 13734 14858 13748
rect 187 13716 3099 13730
rect 11872 13720 14858 13734
rect 187 13702 3113 13716
rect 11886 13706 14858 13720
rect 187 13688 3127 13702
rect 11900 13692 14858 13706
rect 187 13674 3141 13688
rect 11914 13678 14858 13692
rect 187 13660 3155 13674
rect 11928 13664 14858 13678
rect 187 13646 3169 13660
rect 11942 13650 14858 13664
rect 187 13632 3183 13646
rect 11956 13636 14858 13650
rect 187 13618 3197 13632
rect 11970 13622 14858 13636
rect 187 13604 3211 13618
rect 11984 13608 14858 13622
rect 187 13590 3225 13604
rect 11998 13594 14858 13608
rect 187 13576 3239 13590
rect 12012 13580 14858 13594
rect 187 13562 3253 13576
rect 12026 13566 14858 13580
rect 187 13548 3267 13562
rect 12040 13552 14858 13566
rect 187 13534 3281 13548
rect 12054 13538 14858 13552
rect 187 13520 3295 13534
rect 12068 13524 14858 13538
rect 187 13506 3309 13520
rect 12082 13510 14858 13524
rect 187 13492 3323 13506
rect 12096 13496 14858 13510
rect 187 13478 3337 13492
rect 12110 13482 14858 13496
rect 187 13464 3351 13478
rect 12124 13468 14858 13482
rect 187 13450 3365 13464
rect 12138 13454 14858 13468
rect 187 13436 3379 13450
rect 12152 13440 14858 13454
rect 187 13422 3393 13436
rect 12166 13426 14858 13440
rect 187 13408 3407 13422
rect 12180 13412 14858 13426
rect 187 13394 3421 13408
rect 12194 13398 14858 13412
rect 187 13380 3435 13394
rect 12208 13384 14858 13398
rect 187 13366 3449 13380
rect 187 13352 3463 13366
rect 187 13338 3477 13352
rect 187 13324 3491 13338
rect 187 13310 3505 13324
rect 187 13296 3519 13310
rect 187 11556 11342 13296
rect 187 11543 3524 11556
rect 187 11529 3510 11543
rect 187 11515 3496 11529
rect 187 11501 3482 11515
rect 187 11500 3468 11501
rect 12222 11945 14858 13384
rect 12219 11931 14858 11945
rect 12205 11917 14858 11931
rect 12194 11500 14858 11917
rect 187 11347 3319 11500
rect 187 11333 3314 11347
rect 187 11319 3300 11333
rect 187 11305 3286 11319
rect 187 11291 3272 11305
rect 187 11277 3258 11291
rect 187 11263 3244 11277
rect 187 11259 3230 11263
rect 11785 11497 14858 11500
rect 11771 11483 14858 11497
rect 11757 11469 14858 11483
rect 11743 11455 14858 11469
rect 11734 11259 14858 11455
rect 187 11067 3041 11259
rect 187 11053 3034 11067
rect 187 11039 3020 11053
rect 187 11025 3006 11039
rect 187 11011 2992 11025
rect 187 10997 2978 11011
rect 187 10983 2964 10997
rect 187 10981 2950 10983
rect 11533 11245 14858 11259
rect 11519 11231 14858 11245
rect 3770 11219 14858 11231
rect 3758 10981 14858 11219
rect 187 10899 2880 10981
rect 187 10885 2866 10899
rect 187 10871 2852 10885
rect 187 10857 2838 10871
rect 187 8600 2824 10857
rect 3520 10967 14858 10981
rect 3506 10953 14858 10967
rect 3361 9491 14858 10953
rect 11508 9478 14858 9491
rect 11522 9464 14858 9478
rect 11536 9450 14858 9464
rect 11550 9436 14858 9450
rect 11564 9422 14858 9436
rect 11578 9408 14858 9422
rect 11592 9394 14858 9408
rect 11606 9380 14858 9394
rect 11620 9366 14858 9380
rect 11634 9352 14858 9366
rect 11648 9338 14858 9352
rect 11662 9324 14858 9338
rect 11676 9310 14858 9324
rect 11690 9296 14858 9310
rect 11704 9282 14858 9296
rect 11718 9268 14858 9282
rect 11732 9254 14858 9268
rect 11746 9240 14858 9254
rect 11760 9226 14858 9240
rect 11774 9212 14858 9226
rect 11788 9198 14858 9212
rect 11802 9184 14858 9198
rect 11816 9170 14858 9184
rect 11830 9156 14858 9170
rect 11844 9142 14858 9156
rect 11858 9128 14858 9142
rect 11872 9114 14858 9128
rect 11886 9100 14858 9114
rect 11900 9086 14858 9100
rect 11914 9072 14858 9086
rect 11928 9058 14858 9072
rect 11942 9044 14858 9058
rect 11956 9030 14858 9044
rect 11970 9016 14858 9030
rect 11984 9002 14858 9016
rect 11998 8988 14858 9002
rect 12012 8974 14858 8988
rect 12026 8960 14858 8974
rect 12040 8946 14858 8960
rect 12054 8932 14858 8946
rect 12068 8918 14858 8932
rect 12082 8904 14858 8918
rect 12096 8890 14858 8904
rect 12110 8876 14858 8890
rect 12124 8862 14858 8876
rect 12138 8848 14858 8862
rect 12152 8834 14858 8848
rect 12166 8820 14858 8834
rect 12180 8806 14858 8820
rect 12194 8792 14858 8806
rect 12208 8778 14858 8792
rect 187 8586 2837 8600
rect 187 8572 2851 8586
rect 187 8558 2865 8572
rect 187 8544 2879 8558
rect 187 8530 2893 8544
rect 187 8516 2907 8530
rect 187 8502 2921 8516
rect 187 8488 2935 8502
rect 187 8474 2949 8488
rect 187 8460 2963 8474
rect 187 8446 2977 8460
rect 187 8432 2991 8446
rect 187 8418 3005 8432
rect 187 8404 3019 8418
rect 187 8390 3033 8404
rect 187 8376 3047 8390
rect 187 8362 3061 8376
rect 187 8348 3075 8362
rect 187 8334 3089 8348
rect 187 8320 3103 8334
rect 187 8306 3117 8320
rect 187 8292 3131 8306
rect 187 8278 3145 8292
rect 187 8264 3159 8278
rect 187 8250 3173 8264
rect 187 8236 3187 8250
rect 187 8222 3201 8236
rect 187 8208 3215 8222
rect 187 8194 3229 8208
rect 187 8180 3243 8194
rect 187 8166 3257 8180
rect 187 8152 3271 8166
rect 187 8138 3285 8152
rect 187 8124 3299 8138
rect 187 8110 3313 8124
rect 187 8096 3327 8110
rect 187 8082 3341 8096
rect 187 8068 3355 8082
rect 187 8054 3369 8068
rect 187 8040 3383 8054
rect 187 8026 3397 8040
rect 187 8017 11290 8026
rect 187 8003 11299 8017
rect 187 7989 11313 8003
rect 187 7975 11327 7989
rect 187 7961 11341 7975
rect 187 7947 11355 7961
rect 187 7933 11369 7947
rect 187 7620 11383 7933
rect 187 7615 3545 7620
rect 187 7601 3531 7615
rect 10766 7610 11383 7620
rect 187 7587 3517 7601
rect 10780 7596 11383 7610
rect 187 7573 3503 7587
rect 187 7564 3489 7573
rect 10794 7582 11383 7596
rect 10808 7568 11383 7582
rect 187 7503 3428 7564
rect 10822 7554 11383 7568
rect 10836 7540 11383 7554
rect 10850 7526 11383 7540
rect 10864 7512 11383 7526
rect 187 7489 3419 7503
rect 10878 7498 11383 7512
rect 187 7475 3405 7489
rect 10892 7484 11383 7498
rect 187 7461 3391 7475
rect 10906 7470 11383 7484
rect 187 7447 3377 7461
rect 10920 7456 11383 7470
rect 187 7433 3363 7447
rect 187 7419 3349 7433
rect 187 7405 3335 7419
rect 187 7391 3321 7405
rect 187 7377 3307 7391
rect 187 7363 3293 7377
rect 187 7349 3279 7363
rect 187 7335 3265 7349
rect 187 7321 3251 7335
rect 187 7312 3237 7321
rect 187 7279 3204 7312
rect 187 7265 3195 7279
rect 187 7251 3181 7265
rect 187 7237 3167 7251
rect 187 7223 3153 7237
rect 187 7209 3139 7223
rect 187 7195 3125 7209
rect 10934 7223 11383 7456
rect 187 7181 3111 7195
rect 187 7167 3097 7181
rect 187 7153 3083 7167
rect 187 7139 3069 7153
rect 187 7125 3055 7139
rect 187 5854 3041 7125
rect 12222 6182 14858 8778
rect 12213 6168 14858 6182
rect 12199 6154 14858 6168
rect 12194 5886 14858 6154
rect 11919 5874 14858 5886
rect 11905 5860 14858 5874
rect 187 5840 3050 5854
rect 11891 5846 14858 5860
rect 187 5826 3064 5840
rect 187 5812 3078 5826
rect 187 5798 3092 5812
rect 187 5784 3106 5798
rect 187 5770 3120 5784
rect 187 5756 3134 5770
rect 187 5742 3148 5756
rect 187 5728 3162 5742
rect 187 5714 3176 5728
rect 187 5700 3190 5714
rect 187 5686 3204 5700
rect 187 5672 3218 5686
rect 187 5658 3232 5672
rect 187 5644 3246 5658
rect 187 5630 3260 5644
rect 187 5616 3274 5630
rect 187 5602 3288 5616
rect 187 5588 3302 5602
rect 187 5574 3316 5588
rect 187 5560 3330 5574
rect 187 5546 3344 5560
rect 187 5532 3358 5546
rect 187 5518 3372 5532
rect 187 5504 3386 5518
rect 187 5490 3400 5504
rect 187 5476 3414 5490
rect 187 5462 3428 5476
rect 187 5448 3442 5462
rect 187 5434 3456 5448
rect 187 5420 3470 5434
rect 187 5406 3484 5420
rect 187 5392 3498 5406
rect 187 5378 3512 5392
rect 187 5364 3526 5378
rect 187 5350 3540 5364
rect 187 5336 3554 5350
rect 187 5322 3568 5336
rect 187 5308 3582 5322
rect 187 5294 3596 5308
rect 187 5280 3610 5294
rect 187 5266 3624 5280
rect 187 5252 3638 5266
rect 187 5238 3652 5252
rect 187 5224 3666 5238
rect 187 5210 3680 5224
rect 187 5196 3694 5210
rect 11878 5196 14858 5846
rect 187 5182 3708 5196
rect 187 5168 3722 5182
rect 187 5154 3736 5168
rect 11233 5188 14858 5196
rect 11219 5174 14858 5188
rect 11205 5160 14858 5174
rect 187 5140 3750 5154
rect 187 2480 7379 5140
rect 187 2475 5635 2480
rect 187 2461 5621 2475
rect 187 2447 5607 2461
rect 187 2433 5593 2447
rect 187 2424 5579 2433
rect 11191 5146 14858 5160
rect 11177 5132 14858 5146
rect 7578 2459 14858 5132
rect 9350 2453 14858 2459
rect 9364 2439 14858 2453
rect 9378 2425 14858 2439
rect 187 1803 4953 2424
rect 9392 2411 14858 2425
rect 9406 2397 14858 2411
rect 9420 2383 14858 2397
rect 9434 2369 14858 2383
rect 9448 2355 14858 2369
rect 9462 2341 14858 2355
rect 9476 2327 14858 2341
rect 9490 2313 14858 2327
rect 9504 2299 14858 2313
rect 9518 2285 14858 2299
rect 9532 2271 14858 2285
rect 9546 2257 14858 2271
rect 9560 2243 14858 2257
rect 9574 2229 14858 2243
rect 9588 2215 14858 2229
rect 9602 2201 14858 2215
rect 9616 2187 14858 2201
rect 9630 2173 14858 2187
rect 9644 2159 14858 2173
rect 9658 2145 14858 2159
rect 9672 2131 14858 2145
rect 9686 2117 14858 2131
rect 9700 2103 14858 2117
rect 9714 2089 14858 2103
rect 9728 2075 14858 2089
rect 9742 2061 14858 2075
rect 9756 2047 14858 2061
rect 9770 2033 14858 2047
rect 9784 2019 14858 2033
rect 9798 2005 14858 2019
rect 9812 1991 14858 2005
rect 9826 1977 14858 1991
rect 9840 1963 14858 1977
rect 9854 1949 14858 1963
rect 9868 1935 14858 1949
rect 9882 1921 14858 1935
rect 9896 1907 14858 1921
rect 9910 1893 14858 1907
rect 9924 1879 14858 1893
rect 9938 1865 14858 1879
rect 9952 1851 14858 1865
rect 9966 1837 14858 1851
rect 9980 1823 14858 1837
rect 187 1789 4949 1803
rect 9994 1809 14858 1823
rect 187 1775 4935 1789
rect 10008 1795 14858 1809
rect 187 1761 4921 1775
rect 10022 1781 14858 1795
rect 187 1747 4907 1761
rect 10036 1767 14858 1781
rect 187 1733 4893 1747
rect 10050 1753 14858 1767
rect 187 495 4879 1733
rect 10064 1739 14858 1753
rect 183 481 4879 495
rect 169 467 4879 481
rect 155 453 4879 467
rect 141 439 4879 453
rect 131 434 4879 439
rect 127 425 4879 434
rect 113 411 4879 425
rect 99 0 4879 411
rect 5179 0 5579 384
rect 10078 0 14858 1739
<< obsm2 >>
rect 0 39071 15000 40000
rect 0 434 131 39071
rect 13496 38056 15000 39071
rect 3017 38031 15000 38056
rect 2880 37034 3333 38031
rect 2883 37031 3333 37034
rect 2897 37017 11727 37031
rect 2911 37003 11727 37017
rect 2923 36991 11727 37003
rect 2937 36977 11728 36991
rect 2951 36963 11742 36977
rect 2965 36949 11756 36963
rect 2979 36935 11770 36949
rect 2993 36921 11784 36935
rect 3007 36907 11798 36921
rect 3021 36893 11812 36907
rect 3035 36879 11826 36893
rect 3049 36865 11840 36879
rect 3063 36851 11854 36865
rect 3077 36837 11868 36851
rect 3120 36794 11921 36837
rect 3123 36791 11964 36794
rect 3137 36777 11964 36791
rect 3151 36763 11964 36777
rect 3165 36749 11964 36763
rect 3179 36735 11970 36749
rect 3193 36721 11984 36735
rect 3207 36707 11998 36721
rect 3221 36693 12012 36707
rect 3235 36679 12026 36693
rect 3249 36665 12040 36679
rect 3263 36651 12054 36665
rect 3277 36637 12068 36651
rect 3291 36623 12082 36637
rect 3305 36609 12096 36623
rect 3319 36595 12110 36609
rect 3333 36581 12124 36595
rect 3347 36567 12138 36581
rect 3350 36564 12152 36567
rect 3361 36553 12194 36564
rect 3366 36548 12194 36553
rect 3380 36534 12194 36548
rect 3394 36520 12194 36534
rect 3408 36506 12194 36520
rect 3422 36492 12194 36506
rect 3436 36478 12194 36492
rect 3450 36464 12194 36478
rect 3464 36450 12194 36464
rect 3478 36436 12194 36450
rect 3492 36422 12194 36436
rect 3506 36408 12194 36422
rect 3520 36394 12194 36408
rect 3534 36380 12194 36394
rect 3548 36366 12194 36380
rect 3562 36352 12194 36366
rect 11648 34500 12194 36352
rect 3318 34259 11742 34500
rect 2880 32463 3333 34259
rect 2880 32439 11493 32463
rect 2882 32437 3305 32439
rect 2884 32435 3305 32437
rect 3557 32435 11517 32439
rect 2895 32424 11517 32435
rect 2909 32410 11517 32424
rect 2923 32396 11517 32410
rect 2937 32382 11521 32396
rect 2951 32368 11535 32382
rect 2965 32354 11549 32368
rect 2979 32340 11563 32354
rect 2993 32326 11577 32340
rect 3007 32312 11591 32326
rect 3021 32298 11605 32312
rect 3035 32284 11619 32298
rect 3049 32270 11633 32284
rect 3063 32256 11647 32270
rect 3077 32242 11661 32256
rect 3091 32228 11675 32242
rect 3105 32214 11689 32228
rect 3119 32200 11703 32214
rect 3133 32186 11717 32200
rect 3147 32172 11731 32186
rect 3161 32158 11745 32172
rect 3175 32144 11759 32158
rect 3189 32130 11773 32144
rect 3203 32116 11787 32130
rect 3217 32102 11801 32116
rect 3231 32088 11815 32102
rect 3245 32074 11829 32088
rect 3259 32060 11843 32074
rect 3273 32046 11857 32060
rect 3287 32032 11871 32046
rect 3301 32018 11885 32032
rect 3315 32004 11899 32018
rect 3329 31990 11913 32004
rect 3343 31976 11927 31990
rect 3357 31962 11941 31976
rect 3371 31948 11955 31962
rect 3385 31934 11969 31948
rect 3399 31920 11983 31934
rect 3413 31906 11997 31920
rect 3427 31892 12011 31906
rect 3441 31878 12025 31892
rect 3455 31864 12039 31878
rect 3469 31850 12053 31864
rect 3483 31836 12067 31850
rect 3497 31822 12081 31836
rect 3511 31808 12095 31822
rect 3525 31794 12109 31808
rect 3539 31780 12123 31794
rect 3553 31766 12137 31780
rect 3557 31762 12151 31766
rect 3567 31752 12194 31762
rect 11397 29900 12194 31752
rect 3319 29659 11726 29900
rect 3014 29354 3638 29659
rect 2880 27863 3333 29354
rect 2880 27857 11490 27863
rect 2891 27846 3305 27857
rect 2902 27835 3305 27846
rect 3578 27835 11496 27857
rect 2913 27824 11496 27835
rect 2927 27810 11496 27824
rect 2941 27796 11504 27810
rect 2955 27782 11518 27796
rect 2969 27768 11532 27782
rect 2983 27754 11546 27768
rect 2997 27740 11560 27754
rect 3011 27726 11574 27740
rect 3025 27712 11588 27726
rect 3039 27698 11602 27712
rect 3053 27684 11616 27698
rect 3067 27670 11630 27684
rect 3081 27656 11644 27670
rect 3095 27642 11658 27656
rect 3109 27628 11672 27642
rect 3123 27614 11686 27628
rect 3137 27600 11700 27614
rect 3151 27586 11714 27600
rect 3165 27572 11728 27586
rect 3179 27558 11742 27572
rect 3193 27544 11756 27558
rect 3207 27530 11770 27544
rect 3221 27516 11784 27530
rect 3235 27502 11798 27516
rect 3249 27488 11812 27502
rect 3263 27474 11826 27488
rect 3277 27460 11840 27474
rect 3291 27446 11854 27460
rect 3305 27432 11868 27446
rect 3319 27418 11882 27432
rect 3333 27404 11896 27418
rect 3347 27390 11910 27404
rect 3361 27376 11924 27390
rect 3375 27362 11938 27376
rect 3389 27348 11952 27362
rect 3403 27334 11966 27348
rect 3417 27320 11980 27334
rect 3431 27306 11994 27320
rect 3445 27292 12008 27306
rect 3459 27278 12022 27292
rect 3473 27264 12036 27278
rect 3487 27250 12050 27264
rect 3501 27236 12064 27250
rect 3515 27222 12078 27236
rect 3529 27208 12092 27222
rect 3543 27194 12106 27208
rect 3557 27180 12120 27194
rect 3571 27166 12134 27180
rect 3578 27159 12148 27166
rect 3585 27152 12194 27159
rect 11397 25300 12194 27152
rect 3333 25059 11740 25300
rect 2880 23263 4936 25059
rect 2880 23236 11483 23263
rect 2881 23235 11510 23236
rect 2892 23224 11510 23235
rect 2906 23210 11510 23224
rect 2920 23196 11510 23210
rect 2934 23182 11511 23196
rect 2948 23168 11525 23182
rect 2962 23154 11539 23168
rect 2976 23140 11553 23154
rect 2990 23126 11567 23140
rect 3004 23112 11581 23126
rect 3018 23098 11595 23112
rect 3032 23084 11609 23098
rect 3046 23070 11623 23084
rect 3060 23056 11637 23070
rect 3074 23042 11651 23056
rect 3088 23028 11665 23042
rect 3102 23014 11679 23028
rect 3116 23000 11693 23014
rect 3130 22986 11707 23000
rect 3144 22972 11721 22986
rect 3158 22958 11735 22972
rect 3172 22944 11749 22958
rect 3186 22930 11763 22944
rect 3200 22916 11777 22930
rect 3214 22902 11791 22916
rect 3228 22888 11805 22902
rect 3242 22874 11819 22888
rect 3256 22860 11833 22874
rect 3270 22846 11847 22860
rect 3284 22832 11861 22846
rect 3298 22818 11875 22832
rect 3312 22804 11889 22818
rect 3326 22790 11903 22804
rect 3340 22776 11917 22790
rect 3354 22762 11931 22776
rect 3368 22748 11945 22762
rect 3382 22734 11959 22748
rect 3396 22720 11973 22734
rect 3410 22706 11987 22720
rect 3424 22692 12001 22706
rect 3438 22678 12015 22692
rect 3452 22664 12029 22678
rect 3466 22650 12043 22664
rect 3480 22636 12057 22650
rect 3494 22622 12071 22636
rect 3508 22608 12085 22622
rect 3522 22594 12099 22608
rect 3536 22580 12113 22594
rect 3550 22566 12127 22580
rect 3564 22552 12141 22566
rect 11397 20700 12194 22552
rect 3314 20459 11740 20700
rect 2880 18663 4936 20459
rect 2880 18628 11501 18663
rect 2891 18617 11536 18628
rect 2905 18603 11536 18617
rect 2919 18589 11536 18603
rect 2933 18575 11536 18589
rect 2947 18561 11550 18575
rect 2961 18547 11564 18561
rect 2975 18533 11578 18547
rect 2989 18519 11592 18533
rect 3003 18505 11606 18519
rect 3017 18491 11620 18505
rect 3031 18477 11634 18491
rect 3045 18463 11648 18477
rect 3059 18449 11662 18463
rect 3073 18435 11676 18449
rect 3087 18421 11690 18435
rect 3101 18407 11704 18421
rect 3115 18393 11718 18407
rect 3129 18379 11732 18393
rect 3143 18365 11746 18379
rect 3157 18351 11760 18365
rect 3171 18337 11774 18351
rect 3185 18323 11788 18337
rect 3199 18309 11802 18323
rect 3213 18295 11816 18309
rect 3227 18281 11830 18295
rect 3241 18267 11844 18281
rect 3255 18253 11858 18267
rect 3269 18239 11872 18253
rect 3283 18225 11886 18239
rect 3297 18211 11900 18225
rect 3311 18197 11914 18211
rect 3325 18183 11928 18197
rect 3339 18169 11942 18183
rect 3353 18155 11956 18169
rect 3367 18141 11970 18155
rect 3381 18127 11984 18141
rect 3395 18113 11998 18127
rect 3409 18099 12012 18113
rect 3423 18085 12026 18099
rect 3437 18071 12040 18085
rect 3451 18057 12054 18071
rect 3465 18043 12068 18057
rect 3479 18029 12082 18043
rect 3493 18015 12096 18029
rect 3507 18001 12110 18015
rect 3521 17987 12124 18001
rect 3535 17973 12138 17987
rect 3538 17970 12152 17973
rect 3549 17959 12194 17970
rect 3550 17958 12194 17959
rect 3553 17955 12194 17958
rect 3556 17952 12194 17955
rect 11397 16100 12194 17952
rect 3314 15859 11740 16100
rect 2880 14944 4936 15859
rect 2880 14770 3654 14944
rect 2880 14728 4751 14770
rect 2880 14714 4754 14728
rect 2880 14700 4768 14714
rect 2880 14686 4782 14700
rect 2880 14672 4796 14686
rect 2880 14658 4810 14672
rect 2880 14644 4824 14658
rect 2880 14630 4838 14644
rect 2880 14616 4852 14630
rect 2880 14602 4866 14616
rect 2880 14588 4880 14602
rect 2880 14585 4894 14588
rect 2880 14063 4936 14585
rect 2880 14028 11489 14063
rect 2884 14024 11524 14028
rect 2898 14010 11524 14024
rect 2912 13996 11524 14010
rect 2926 13982 11524 13996
rect 2940 13968 11531 13982
rect 2954 13954 11545 13968
rect 2968 13940 11559 13954
rect 2982 13926 11573 13940
rect 2996 13912 11587 13926
rect 3010 13898 11601 13912
rect 3024 13884 11615 13898
rect 3038 13870 11629 13884
rect 3052 13856 11643 13870
rect 3066 13842 11657 13856
rect 3080 13828 11671 13842
rect 3094 13814 11685 13828
rect 3108 13800 11699 13814
rect 3122 13786 11713 13800
rect 3136 13772 11727 13786
rect 3150 13758 11741 13772
rect 3164 13744 11755 13758
rect 3178 13730 11769 13744
rect 3192 13716 11783 13730
rect 3206 13702 11797 13716
rect 3220 13688 11811 13702
rect 3234 13674 11825 13688
rect 3248 13660 11839 13674
rect 3262 13646 11853 13660
rect 3276 13632 11867 13646
rect 3290 13618 11881 13632
rect 3304 13604 11895 13618
rect 3318 13590 11909 13604
rect 3332 13576 11923 13590
rect 3346 13562 11937 13576
rect 3360 13548 11951 13562
rect 3374 13534 11965 13548
rect 3388 13520 11979 13534
rect 3402 13506 11993 13520
rect 3416 13492 12007 13506
rect 3430 13478 12021 13492
rect 3444 13464 12035 13478
rect 3458 13450 12049 13464
rect 3472 13436 12063 13450
rect 3486 13422 12077 13436
rect 3500 13408 12091 13422
rect 3514 13394 12105 13408
rect 3528 13380 12119 13394
rect 3542 13366 12133 13380
rect 3550 13358 12147 13366
rect 3556 13352 12194 13358
rect 11398 11500 12194 13352
rect 3319 11259 11734 11500
rect 3041 10981 3758 11259
rect 2880 9463 3333 10981
rect 2880 9413 11483 9463
rect 2880 9399 11494 9413
rect 2880 9385 11508 9399
rect 2880 9371 11522 9385
rect 2880 9357 11536 9371
rect 2880 9343 11550 9357
rect 2880 9329 11564 9343
rect 2880 9315 11578 9329
rect 2880 9301 11592 9315
rect 2880 9287 11606 9301
rect 2880 9273 11620 9287
rect 2880 9259 11634 9273
rect 2880 9245 11648 9259
rect 2880 9231 11662 9245
rect 2880 9217 11676 9231
rect 2880 9203 11690 9217
rect 2880 9189 11704 9203
rect 2880 9175 11718 9189
rect 2880 9161 11732 9175
rect 2880 9147 11746 9161
rect 2880 9133 11760 9147
rect 2880 9119 11774 9133
rect 2880 9105 11788 9119
rect 2880 9091 11802 9105
rect 2880 9077 11816 9091
rect 2880 9063 11830 9077
rect 2880 9049 11844 9063
rect 2880 9035 11858 9049
rect 2880 9021 11872 9035
rect 2880 9007 11886 9021
rect 2880 8993 11900 9007
rect 2880 8979 11914 8993
rect 2880 8965 11928 8979
rect 2880 8951 11942 8965
rect 2880 8937 11956 8951
rect 2880 8923 11970 8937
rect 2880 8909 11984 8923
rect 2880 8895 11998 8909
rect 2880 8881 12012 8895
rect 2880 8867 12026 8881
rect 2880 8853 12040 8867
rect 2880 8839 12054 8853
rect 2880 8825 12068 8839
rect 2880 8811 12082 8825
rect 2880 8797 12096 8811
rect 2880 8783 12110 8797
rect 2880 8769 12124 8783
rect 2880 8755 12138 8769
rect 2880 8752 12152 8755
rect 2880 8636 12194 8752
rect 2888 8628 12194 8636
rect 2902 8614 12194 8628
rect 2916 8600 12194 8614
rect 2930 8586 12194 8600
rect 2944 8572 12194 8586
rect 2958 8558 12194 8572
rect 2972 8544 12194 8558
rect 2986 8530 12194 8544
rect 3000 8516 12194 8530
rect 3014 8502 12194 8516
rect 3028 8488 12194 8502
rect 3042 8474 12194 8488
rect 3056 8460 12194 8474
rect 3070 8446 12194 8460
rect 3084 8432 12194 8446
rect 3098 8418 12194 8432
rect 3112 8404 12194 8418
rect 3126 8390 12194 8404
rect 3140 8376 12194 8390
rect 3154 8362 12194 8376
rect 3168 8348 12194 8362
rect 3182 8334 12194 8348
rect 3196 8320 12194 8334
rect 3210 8306 12194 8320
rect 3224 8292 12194 8306
rect 3238 8278 12194 8292
rect 3252 8264 12194 8278
rect 3266 8250 12194 8264
rect 3280 8236 12194 8250
rect 3294 8222 12194 8236
rect 3308 8208 12194 8222
rect 3322 8194 12194 8208
rect 3336 8180 12194 8194
rect 3350 8166 12194 8180
rect 3364 8152 12194 8166
rect 3378 8138 12194 8152
rect 3392 8124 12194 8138
rect 3406 8110 12194 8124
rect 3420 8096 12194 8110
rect 3434 8082 12194 8096
rect 3541 8054 10136 8082
rect 11327 8068 12194 8082
rect 11341 8054 12194 8068
rect 11355 8040 12194 8054
rect 11369 8026 12194 8040
rect 11383 8012 12194 8026
rect 11397 7998 12194 8012
rect 11411 7984 12194 7998
rect 11425 7970 12194 7984
rect 3652 7564 10626 7592
rect 3428 7559 10733 7564
rect 3428 7545 10738 7559
rect 3428 7531 10752 7545
rect 3428 7517 10766 7531
rect 3428 7503 10780 7517
rect 3428 7489 10794 7503
rect 3428 7475 10808 7489
rect 3428 7461 10822 7475
rect 3428 7447 10836 7461
rect 3428 7433 10850 7447
rect 3428 7419 10864 7433
rect 3349 7340 10878 7419
rect 3321 7312 10878 7340
rect 3204 7195 10906 7312
rect 3176 7167 11023 7195
rect 11439 7167 12194 7970
rect 3097 5886 12194 7167
rect 3101 5882 11878 5886
rect 3115 5868 11878 5882
rect 3129 5854 11878 5868
rect 3143 5840 11878 5854
rect 3157 5826 11878 5840
rect 3171 5812 11878 5826
rect 3185 5798 11878 5812
rect 3199 5784 11878 5798
rect 3213 5770 11878 5784
rect 3227 5756 11878 5770
rect 3241 5742 11878 5756
rect 3255 5728 11878 5742
rect 3269 5714 11878 5728
rect 3283 5700 11878 5714
rect 3297 5686 11878 5700
rect 3311 5672 11878 5686
rect 3325 5658 11878 5672
rect 3339 5644 11878 5658
rect 3353 5630 11878 5644
rect 3367 5616 11878 5630
rect 3381 5602 11878 5616
rect 3395 5588 11878 5602
rect 3409 5574 11878 5588
rect 3423 5560 11878 5574
rect 3437 5546 11878 5560
rect 3451 5532 11878 5546
rect 3465 5518 11878 5532
rect 3479 5504 11878 5518
rect 3493 5490 11878 5504
rect 3507 5476 11878 5490
rect 3521 5462 11878 5476
rect 3535 5448 11878 5462
rect 3549 5434 11878 5448
rect 3563 5420 11878 5434
rect 3577 5406 11878 5420
rect 3591 5392 11878 5406
rect 3605 5378 11878 5392
rect 3619 5364 11878 5378
rect 3633 5350 11878 5364
rect 3647 5336 11878 5350
rect 3661 5322 11878 5336
rect 3675 5308 11878 5322
rect 3689 5294 11878 5308
rect 3703 5280 11878 5294
rect 3717 5266 11878 5280
rect 3731 5252 11878 5266
rect 3745 5238 11878 5252
rect 3759 5224 11878 5238
rect 3773 5210 11878 5224
rect 3787 5196 11878 5210
rect 7435 5160 11187 5196
rect 7435 2431 7550 5160
rect 7435 2424 9332 2431
rect 4953 2374 9339 2424
rect 4953 2360 9350 2374
rect 4953 2346 9364 2360
rect 4953 2332 9378 2346
rect 4953 2318 9392 2332
rect 4953 2304 9406 2318
rect 4953 2290 9420 2304
rect 4953 2276 9434 2290
rect 4953 2262 9448 2276
rect 4953 2248 9462 2262
rect 4953 2234 9476 2248
rect 4953 2220 9490 2234
rect 4953 2206 9504 2220
rect 4953 2192 9518 2206
rect 4953 2178 9532 2192
rect 4953 2164 9546 2178
rect 4953 2150 9560 2164
rect 4953 2136 9574 2150
rect 4953 2122 9588 2136
rect 4953 2108 9602 2122
rect 4953 2094 9616 2108
rect 4953 2080 9630 2094
rect 4953 2066 9644 2080
rect 4953 2052 9658 2066
rect 4953 2038 9672 2052
rect 4953 2024 9686 2038
rect 4953 2010 9700 2024
rect 4953 1996 9714 2010
rect 4953 1982 9728 1996
rect 4953 1968 9742 1982
rect 4953 1954 9756 1968
rect 4953 1940 9770 1954
rect 4953 1926 9784 1940
rect 4953 1912 9798 1926
rect 4953 1898 9812 1912
rect 4953 1884 9826 1898
rect 4953 1870 9840 1884
rect 4953 1856 9854 1870
rect 4953 1842 9868 1856
rect 4953 1828 9882 1842
rect 4953 1814 9896 1828
rect 4953 1800 9910 1814
rect 4953 1786 9924 1800
rect 4953 1772 9938 1786
rect 4953 1758 9952 1772
rect 4953 1744 9966 1758
rect 4953 1730 9980 1744
rect 4953 1716 9994 1730
rect 4953 1713 10008 1716
rect 0 0 43 434
rect 4935 412 10050 1713
rect 4935 0 5151 412
rect 5607 0 10050 412
rect 14886 0 15000 38031
<< metal3 >>
rect 2525 35179 5002 39015
rect 2530 35174 5002 35179
rect 2560 35144 5002 35174
rect 2590 35114 5002 35144
rect 2620 35084 5002 35114
rect 2650 35054 5002 35084
rect 2680 35024 5002 35054
rect 2710 34994 5002 35024
rect 2740 34964 5002 34994
rect 2770 34934 5002 34964
rect 2800 34904 5002 34934
rect 2830 34874 5002 34904
rect 2860 34844 5002 34874
rect 2890 34814 5002 34844
rect 2920 34784 5002 34814
rect 2950 34754 5002 34784
rect 2980 34724 5002 34754
rect 3010 34694 5002 34724
rect 3040 34664 5002 34694
rect 3070 34634 5002 34664
rect 3100 34528 5002 34634
rect 5186 35070 7364 39015
rect 7593 35070 9771 38004
rect 5186 35052 7346 35070
rect 7611 35052 9771 35070
rect 5186 35022 7316 35052
rect 7641 35022 9771 35052
rect 5186 34992 7286 35022
rect 7671 34992 9771 35022
rect 5186 34962 7256 34992
rect 7701 34962 9771 34992
rect 5186 34932 7226 34962
rect 7731 34932 9771 34962
rect 5186 34902 7196 34932
rect 7761 34902 9771 34932
rect 5186 34872 7166 34902
rect 7791 34872 9771 34902
rect 5186 34842 7136 34872
rect 7821 34842 9771 34872
rect 5186 34812 7106 34842
rect 7851 34812 9771 34842
rect 5186 34782 7076 34812
rect 7881 34782 9771 34812
rect 5186 34752 7046 34782
rect 7911 34752 9771 34782
rect 5186 34722 7016 34752
rect 7941 34722 9771 34752
rect 5186 34692 6986 34722
rect 7971 34692 9771 34722
rect 5186 34662 6956 34692
rect 8001 34662 9771 34692
rect 5186 34632 6926 34662
rect 8031 34632 9771 34662
rect 5186 34602 6896 34632
rect 8061 34602 9771 34632
rect 5186 34572 6866 34602
rect 8091 34572 9771 34602
rect 5186 34542 6836 34572
rect 8121 34542 9771 34572
rect 3100 34516 4990 34528
rect 3100 34486 4960 34516
rect 5186 34512 6806 34542
rect 8151 34512 9771 34542
rect 9955 35045 12298 38008
rect 9955 35024 12277 35045
rect 9955 34994 12247 35024
rect 9955 34964 12217 34994
rect 9955 34934 12187 34964
rect 9955 34904 12157 34934
rect 9955 34874 12127 34904
rect 9955 34844 12097 34874
rect 9955 34814 12067 34844
rect 9955 34784 12037 34814
rect 9955 34754 12007 34784
rect 9955 34724 11977 34754
rect 9955 34694 11947 34724
rect 9955 34664 11917 34694
rect 9955 34634 11887 34664
rect 9955 34529 11857 34634
rect 9967 34517 11857 34529
rect 3100 34456 4930 34486
rect 5186 34482 6776 34512
rect 8181 34482 9771 34512
rect 9997 34487 11857 34517
rect 3100 34426 4900 34456
rect 5186 34452 6746 34482
rect 8211 34452 9771 34482
rect 10027 34457 11857 34487
rect 3100 34396 4870 34426
rect 5186 34422 6716 34452
rect 8241 34422 9771 34452
rect 10057 34427 11857 34457
rect 3100 34366 4840 34396
rect 5186 34392 6686 34422
rect 8271 34392 9771 34422
rect 10087 34397 11857 34427
rect 3100 34336 4810 34366
rect 5186 34362 6656 34392
rect 8301 34362 9771 34392
rect 10117 34367 11857 34397
rect 3100 34306 4780 34336
rect 5186 34332 6626 34362
rect 8331 34332 9771 34362
rect 10147 34337 11857 34367
rect 3100 34276 4750 34306
rect 5186 34302 6596 34332
rect 8361 34302 9771 34332
rect 10177 34307 11857 34337
rect 3100 34246 4720 34276
rect 5186 34272 6566 34302
rect 8391 34272 9771 34302
rect 10207 34277 11857 34307
rect 3100 34216 4690 34246
rect 5186 34242 6536 34272
rect 8421 34242 9771 34272
rect 10237 34247 11857 34277
rect 3100 34186 4660 34216
rect 5186 34212 6506 34242
rect 8451 34212 9771 34242
rect 10267 34217 11857 34247
rect 3100 34156 4630 34186
rect 5186 34182 6476 34212
rect 8481 34182 9771 34212
rect 10297 34187 11857 34217
rect 3100 34126 4600 34156
rect 5186 34152 6446 34182
rect 8511 34152 9771 34182
rect 10327 34157 11857 34187
rect 3100 34096 4570 34126
rect 5186 34122 6416 34152
rect 8541 34122 9771 34152
rect 10357 34127 11857 34157
rect 3100 34066 4540 34096
rect 3100 34036 4510 34066
rect 3100 34006 4480 34036
rect 3100 33976 4450 34006
rect 3100 33946 4420 33976
rect 3100 33916 4390 33946
rect 3100 33886 4360 33916
rect 3100 33856 4330 33886
rect 3100 20920 4300 33856
rect 5186 20958 6386 34122
rect 8571 22110 9771 34122
rect 10387 34097 11857 34127
rect 10417 34067 11857 34097
rect 10447 34037 11857 34067
rect 10477 34007 11857 34037
rect 10507 33977 11857 34007
rect 10537 33947 11857 33977
rect 10567 33917 11857 33947
rect 10597 33887 11857 33917
rect 10627 33857 11857 33887
rect 8557 22080 9771 22110
rect 8527 22050 9771 22080
rect 10657 22072 11857 33857
rect 8497 22020 9771 22050
rect 10641 22042 11857 22072
rect 8467 21990 9771 22020
rect 10611 22012 11857 22042
rect 8437 21960 9771 21990
rect 10581 21982 11857 22012
rect 8407 21930 9771 21960
rect 10551 21952 11857 21982
rect 8377 21900 9771 21930
rect 10521 21922 11857 21952
rect 8347 21870 9771 21900
rect 10491 21892 11857 21922
rect 8317 21840 9771 21870
rect 10461 21862 11857 21892
rect 8287 21810 9771 21840
rect 10431 21832 11857 21862
rect 8257 21780 9771 21810
rect 10401 21802 11857 21832
rect 8227 21750 9771 21780
rect 10371 21772 11857 21802
rect 8197 21720 9771 21750
rect 10341 21742 11857 21772
rect 8167 21690 9771 21720
rect 10311 21712 11857 21742
rect 8137 21660 9771 21690
rect 10281 21682 11857 21712
rect 8107 21630 9771 21660
rect 10251 21652 11857 21682
rect 8077 21611 9752 21630
rect 10221 21622 11857 21652
rect 8058 21581 9722 21611
rect 10191 21592 11857 21622
rect 10161 21581 11846 21592
rect 8028 21551 9692 21581
rect 10150 21551 11816 21581
rect 7998 21521 9662 21551
rect 10120 21521 11786 21551
rect 7968 21491 9632 21521
rect 10090 21491 11756 21521
rect 7938 21461 9602 21491
rect 10060 21461 11726 21491
rect 7908 21431 9572 21461
rect 10030 21431 11696 21461
rect 7878 21401 9542 21431
rect 10000 21401 11666 21431
rect 7848 21371 9512 21401
rect 9970 21371 11636 21401
rect 7818 21341 9482 21371
rect 9940 21341 11606 21371
rect 7788 21311 9452 21341
rect 9910 21311 11576 21341
rect 7758 21281 9422 21311
rect 9880 21281 11546 21311
rect 7728 21251 9392 21281
rect 9850 21251 11516 21281
rect 7698 21221 9362 21251
rect 9820 21221 11486 21251
rect 7668 21191 9332 21221
rect 9790 21191 11456 21221
rect 7638 21161 9302 21191
rect 9760 21161 11426 21191
rect 7608 21131 9272 21161
rect 9730 21131 11396 21161
rect 7578 21117 9258 21131
rect 7578 21087 9228 21117
rect 9700 21101 11366 21131
rect 7578 21057 9198 21087
rect 9670 21071 11336 21101
rect 7578 21027 9168 21057
rect 9640 21041 11306 21071
rect 7578 20997 9138 21027
rect 9610 21011 11276 21041
rect 7578 20967 9108 20997
rect 9580 20981 11246 21011
rect 5186 20928 6400 20958
rect 7578 20937 9078 20967
rect 9550 20951 11216 20981
rect 3100 20890 4316 20920
rect 5186 20898 6430 20928
rect 7578 20907 9048 20937
rect 9520 20921 11186 20951
rect 3100 20860 4346 20890
rect 5186 20868 6460 20898
rect 7578 20877 9018 20907
rect 9490 20891 11156 20921
rect 3100 20830 4376 20860
rect 5186 20838 6490 20868
rect 7578 20847 8988 20877
rect 9460 20861 11126 20891
rect 3100 20800 4406 20830
rect 5186 20808 6520 20838
rect 7578 20817 8958 20847
rect 9430 20831 11096 20861
rect 3100 20770 4436 20800
rect 5186 20778 6550 20808
rect 7578 20787 8928 20817
rect 9400 20801 11066 20831
rect 3100 20740 4466 20770
rect 5186 20748 6580 20778
rect 7578 20757 8898 20787
rect 9370 20771 11036 20801
rect 3100 20710 4496 20740
rect 5186 20718 6610 20748
rect 7578 20727 8868 20757
rect 9340 20741 11006 20771
rect 3100 20680 4526 20710
rect 5186 20688 6640 20718
rect 7578 20697 8838 20727
rect 9310 20711 10976 20741
rect 3100 20650 4556 20680
rect 5186 20658 6670 20688
rect 7578 20667 8808 20697
rect 9280 20681 10946 20711
rect 3100 20620 4586 20650
rect 5186 20628 6700 20658
rect 7578 20637 8778 20667
rect 9250 20651 10916 20681
rect 3100 20590 4616 20620
rect 5186 20598 6730 20628
rect 7578 20607 8748 20637
rect 9220 20621 10886 20651
rect 3100 20560 4646 20590
rect 5186 20568 6760 20598
rect 7578 20577 8718 20607
rect 9190 20591 10856 20621
rect 3100 20530 4676 20560
rect 5186 20538 6790 20568
rect 7578 20547 8688 20577
rect 9160 20561 10826 20591
rect 3100 20500 4706 20530
rect 5186 20508 6820 20538
rect 7578 20517 8658 20547
rect 9130 20531 10796 20561
rect 3100 20470 4736 20500
rect 5186 20478 6850 20508
rect 7578 20487 8628 20517
rect 9100 20501 10766 20531
rect 9070 20496 10761 20501
rect 3100 20440 4766 20470
rect 5205 20459 6880 20478
rect 3129 20411 4796 20440
rect 5235 20429 6899 20459
rect 7578 20457 8598 20487
rect 9070 20466 10731 20496
rect 3159 20381 4825 20411
rect 5265 20399 6929 20429
rect 3189 20351 4855 20381
rect 5295 20369 6959 20399
rect 3219 20321 4885 20351
rect 5325 20339 6989 20369
rect 3249 20291 4915 20321
rect 5355 20309 7019 20339
rect 3279 20261 4945 20291
rect 5385 20279 7049 20309
rect 3309 20231 4975 20261
rect 5415 20249 7079 20279
rect 3339 20201 5005 20231
rect 5445 20219 7109 20249
rect 3369 20171 5035 20201
rect 5475 20189 7139 20219
rect 3399 20141 5065 20171
rect 5505 20159 7169 20189
rect 3429 20111 5095 20141
rect 5535 20129 7199 20159
rect 3459 20081 5125 20111
rect 5565 20099 7229 20129
rect 3489 20051 5155 20081
rect 5595 20069 7259 20099
rect 3519 20021 5185 20051
rect 5625 20039 7289 20069
rect 7578 20051 8568 20457
rect 9070 20436 10701 20466
rect 9070 20406 10671 20436
rect 9070 20376 10641 20406
rect 9070 20346 10611 20376
rect 9070 20316 10581 20346
rect 9070 20286 10551 20316
rect 9070 20256 10521 20286
rect 9070 20226 10491 20256
rect 9070 20196 10461 20226
rect 9070 20166 10431 20196
rect 9070 20136 10401 20166
rect 9070 20106 10371 20136
rect 9070 20076 10341 20106
rect 3549 19991 5215 20021
rect 5655 20009 7319 20039
rect 7578 20021 8574 20051
rect 9070 20046 10311 20076
rect 9070 20033 10298 20046
rect 3579 19961 5245 19991
rect 5685 19979 7349 20009
rect 7578 19991 8604 20021
rect 9057 20003 10268 20033
rect 5699 19965 7379 19979
rect 3609 19931 5275 19961
rect 5729 19935 7379 19965
rect 3639 19901 5305 19931
rect 5759 19905 7379 19935
rect 3669 19871 5335 19901
rect 5789 19875 7379 19905
rect 3699 19841 5365 19871
rect 5819 19845 7379 19875
rect 3729 19811 5395 19841
rect 5849 19815 7379 19845
rect 3759 19781 5425 19811
rect 5879 19785 7379 19815
rect 3789 19751 5455 19781
rect 5909 19755 7379 19785
rect 3819 19721 5485 19751
rect 5939 19725 7379 19755
rect 3849 19691 5515 19721
rect 5969 19695 7379 19725
rect 3879 19661 5545 19691
rect 5999 19665 7379 19695
rect 3909 19631 5575 19661
rect 6029 19635 7379 19665
rect 3939 19601 5605 19631
rect 6059 19605 7379 19635
rect 3969 19571 5635 19601
rect 6089 19575 7379 19605
rect 3999 19541 5665 19571
rect 6119 19545 7379 19575
rect 4029 19511 5695 19541
rect 6149 19515 7379 19545
rect 4059 19481 5725 19511
rect 6179 19485 7379 19515
rect 4089 19451 5755 19481
rect 6209 19455 7379 19485
rect 4119 19421 5785 19451
rect 6239 19425 7379 19455
rect 4149 19391 5815 19421
rect 6269 19395 7379 19425
rect 4179 19361 5845 19391
rect 6299 19365 7379 19395
rect 4209 19331 5875 19361
rect 6329 19335 7379 19365
rect 4239 19301 5905 19331
rect 6359 19305 7379 19335
rect 4269 19271 5905 19301
rect 4299 19241 5905 19271
rect 4329 19211 5905 19241
rect 4359 19181 5905 19211
rect 4389 19151 5905 19181
rect 4419 19121 5905 19151
rect 4449 19091 5905 19121
rect 4479 19061 5905 19091
rect 4509 19031 5905 19061
rect 4539 19001 5905 19031
rect 4569 18971 5905 19001
rect 4599 18941 5905 18971
rect 4629 18911 5905 18941
rect 4659 18881 5905 18911
rect 4689 18851 5905 18881
rect 4719 18821 5905 18851
rect 4749 18598 5905 18821
rect 6389 18598 7379 19305
rect 4749 18568 5927 18598
rect 6367 18568 7379 18598
rect 4749 18538 5957 18568
rect 6337 18538 7379 18568
rect 4749 18508 5987 18538
rect 6307 18508 7379 18538
rect 4764 18493 6017 18508
rect 4779 18478 6032 18493
rect 6277 18478 7379 18508
rect 4789 18468 7379 18478
rect 4819 18438 7379 18468
rect 4849 18408 7379 18438
rect 4879 18378 7379 18408
rect 4909 18348 7379 18378
rect 4939 18318 7379 18348
rect 4969 18288 7379 18318
rect 4999 18258 7379 18288
rect 5029 18228 7379 18258
rect 5059 18198 7379 18228
rect 5089 18168 7379 18198
rect 5119 18138 7379 18168
rect 5149 18108 7379 18138
rect 5179 0 7379 18108
rect 7578 19961 8634 19991
rect 9027 19973 10238 20003
rect 7578 19931 8664 19961
rect 8997 19943 10208 19973
rect 7578 19901 8694 19931
rect 8967 19922 10208 19943
rect 8946 19901 10208 19922
rect 7578 19660 10208 19901
rect 7578 19650 10198 19660
rect 7578 19620 10168 19650
rect 7578 19590 10138 19620
rect 7578 19560 10108 19590
rect 7578 19530 10078 19560
rect 7578 19500 10048 19530
rect 7578 19470 10018 19500
rect 7578 19440 9988 19470
rect 7578 19410 9958 19440
rect 7578 19380 9928 19410
rect 7578 19350 9898 19380
rect 7578 19320 9868 19350
rect 7578 19290 9838 19320
rect 7578 19260 9808 19290
rect 7578 0 9778 19260
<< labels >>
rlabel metal1 s 9537 5826 10263 5840 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9523 5812 10263 5826 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9509 5798 10263 5812 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9495 5784 10263 5798 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9481 5770 10263 5784 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9467 5756 10263 5770 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9453 5742 10263 5756 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9439 5728 10263 5742 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9425 5714 10263 5728 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9411 5700 10263 5714 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9397 5686 10263 5700 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9383 5672 10263 5686 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9369 5658 10263 5672 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9355 5644 10263 5658 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9341 5630 10263 5644 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9327 5616 10263 5630 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9313 5602 10263 5616 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9299 5588 10263 5602 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9285 5574 10263 5588 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9271 5560 10263 5574 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9257 5546 10263 5560 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9243 5532 10263 5546 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9229 5518 10263 5532 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9537 5840 10263 7447 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7763 1123 7770 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7749 1109 7763 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7735 1095 7749 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7721 1081 7735 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7707 1067 7721 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7693 1053 7707 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7679 1039 7693 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7665 1025 7679 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7651 1011 7665 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7637 997 7651 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7623 983 7637 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7609 969 7623 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7595 955 7609 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7581 941 7595 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 5831 941 7581 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7770 10263 8496 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9215 7769 10263 7770 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9229 7755 10263 7769 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9243 7741 10263 7755 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9257 7727 10263 7741 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9271 7713 10263 7727 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9285 7699 10263 7713 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9299 7685 10263 7699 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9313 7671 10263 7685 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9327 7657 10263 7671 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9341 7643 10263 7657 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9355 7629 10263 7643 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9369 7615 10263 7629 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9383 7601 10263 7615 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9397 7587 10263 7601 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9411 7573 10263 7587 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9425 7559 10263 7573 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9439 7545 10263 7559 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9453 7531 10263 7545 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9467 7517 10263 7531 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9481 7503 10263 7517 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9495 7489 10263 7503 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9509 7475 10263 7489 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9523 7461 10263 7475 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 9537 7447 10263 7461 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4781 2366 4792 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4767 2352 4781 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4753 2338 4767 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4739 2324 4753 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4725 2310 4739 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4711 2296 4725 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4697 2282 4711 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4683 2268 4697 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4669 2254 4683 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4655 2240 4669 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4641 2226 4655 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4627 2212 4641 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4613 2198 4627 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4599 2184 4613 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4585 2170 4599 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4571 2156 4585 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4557 2142 4571 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4543 2128 4557 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4529 2114 4543 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4515 2100 4529 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4501 2086 4515 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4487 2072 4501 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4473 2058 4487 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4459 2044 4473 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4445 2030 4459 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4431 2016 4445 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4417 2002 4431 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4403 1988 4417 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4389 1974 4403 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4375 1960 4389 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4361 1946 4375 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4347 1932 4361 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4333 1918 4347 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4319 1904 4333 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4305 1890 4319 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4291 1876 4305 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4277 1862 4291 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4263 1848 4277 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4249 1834 4263 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4235 1820 4249 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4221 1806 4235 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4207 1792 4221 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4193 1778 4207 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4179 1764 4193 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4165 1750 4179 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4151 1736 4165 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4137 1722 4151 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4123 1708 4137 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4109 1694 4123 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4095 1680 4109 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4081 1666 4095 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 2 1666 4081 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4792 10263 5518 6 vssd
port 1 nsew ground bidirectional
rlabel metal2 s 5179 0 5579 384 6 ogc_hvc
port 2 nsew power bidirectional
rlabel metal3 s 3100 34528 5002 34604 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2525 35179 5002 39015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2530 35174 5002 35179 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2560 35144 5002 35174 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2590 35114 5002 35144 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2620 35084 5002 35114 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2650 35054 5002 35084 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2680 35024 5002 35054 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2710 34994 5002 35024 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2740 34964 5002 34994 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2770 34934 5002 34964 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2800 34904 5002 34934 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2830 34874 5002 34904 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2860 34844 5002 34874 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2890 34814 5002 34844 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2920 34784 5002 34814 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2950 34754 5002 34784 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 2980 34724 5002 34754 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3010 34694 5002 34724 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3040 34664 5002 34694 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3070 34634 5002 34664 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34604 5002 34634 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34516 4990 34528 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34486 4960 34516 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34456 4930 34486 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34426 4900 34456 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34396 4870 34426 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34366 4840 34396 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34336 4810 34366 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34306 4780 34336 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34276 4750 34306 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34246 4720 34276 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34216 4690 34246 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34186 4660 34216 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34156 4630 34186 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34126 4600 34156 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34096 4570 34126 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34066 4540 34096 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34036 4510 34066 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34006 4480 34036 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33976 4450 34006 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33946 4420 33976 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33916 4390 33946 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33886 4360 33916 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33856 4330 33886 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33826 4300 33856 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 35070 7364 39015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20936 4300 33826 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 35052 7346 35070 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 35022 7316 35052 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34992 7286 35022 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34962 7256 34992 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34932 7226 34962 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34902 7196 34932 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34872 7166 34902 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34842 7136 34872 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34812 7106 34842 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34782 7076 34812 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34752 7046 34782 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34722 7016 34752 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34692 6986 34722 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34662 6956 34692 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34632 6926 34662 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34602 6896 34632 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34572 6866 34602 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34542 6836 34572 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34512 6806 34542 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34482 6776 34512 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34452 6746 34482 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34422 6716 34452 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34392 6686 34422 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34362 6656 34392 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34332 6626 34362 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34302 6596 34332 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34272 6566 34302 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34242 6536 34272 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34212 6506 34242 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34182 6476 34212 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34152 6446 34182 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34122 6416 34152 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34092 6386 34122 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20920 4300 20936 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20890 4316 20920 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20860 4346 20890 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20830 4376 20860 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20800 4406 20830 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20770 4436 20800 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20740 4466 20770 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20710 4496 20740 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20680 4526 20710 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20650 4556 20680 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20620 4586 20650 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20590 4616 20620 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20560 4646 20590 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20530 4676 20560 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20500 4706 20530 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20470 4736 20500 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20440 4766 20470 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20972 6386 34092 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3129 20411 4796 20440 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3159 20381 4825 20411 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3189 20351 4855 20381 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3219 20321 4885 20351 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3249 20291 4915 20321 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3279 20261 4945 20291 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3309 20231 4975 20261 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3339 20201 5005 20231 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3369 20171 5035 20201 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3399 20141 5065 20171 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3429 20111 5095 20141 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3459 20081 5125 20111 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3489 20051 5155 20081 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3519 20021 5185 20051 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3549 19991 5215 20021 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3579 19961 5245 19991 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3609 19931 5275 19961 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3639 19901 5305 19931 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3669 19871 5335 19901 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3699 19841 5365 19871 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3729 19811 5395 19841 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3759 19781 5425 19811 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3789 19751 5455 19781 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3819 19721 5485 19751 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3849 19691 5515 19721 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3879 19661 5545 19691 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3909 19631 5575 19661 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3939 19601 5605 19631 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3969 19571 5635 19601 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3999 19541 5665 19571 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4029 19511 5695 19541 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4059 19481 5725 19511 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4089 19451 5755 19481 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4119 19421 5785 19451 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4149 19391 5815 19421 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4179 19361 5845 19391 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4209 19331 5875 19361 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20958 6386 20972 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20928 6400 20958 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20898 6430 20928 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20868 6460 20898 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20838 6490 20868 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20808 6520 20838 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20778 6550 20808 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20748 6580 20778 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20718 6610 20748 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20688 6640 20718 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20658 6670 20688 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20628 6700 20658 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20598 6730 20628 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20568 6760 20598 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20538 6790 20568 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20508 6820 20538 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20478 6850 20508 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4239 19301 5905 19331 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4269 19271 5905 19301 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4299 19241 5905 19271 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4329 19211 5905 19241 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4359 19181 5905 19211 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4389 19151 5905 19181 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4419 19121 5905 19151 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4449 19091 5905 19121 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4479 19061 5905 19091 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4509 19031 5905 19061 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4539 19001 5905 19031 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4569 18971 5905 19001 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4599 18941 5905 18971 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4629 18911 5905 18941 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4659 18881 5905 18911 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4689 18851 5905 18881 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4719 18821 5905 18851 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18791 5905 18821 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5205 20459 6880 20478 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5235 20429 6899 20459 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5265 20399 6929 20429 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5295 20369 6959 20399 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5325 20339 6989 20369 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5355 20309 7019 20339 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5385 20279 7049 20309 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5415 20249 7079 20279 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5445 20219 7109 20249 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5475 20189 7139 20219 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5505 20159 7169 20189 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5535 20129 7199 20159 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5565 20099 7229 20129 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5595 20069 7259 20099 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5625 20039 7289 20069 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5655 20009 7319 20039 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5685 19979 7349 20009 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18620 5905 18791 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5699 19965 7379 19979 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5729 19935 7379 19965 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5759 19905 7379 19935 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5789 19875 7379 19905 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5819 19845 7379 19875 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5849 19815 7379 19845 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5879 19785 7379 19815 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5909 19755 7379 19785 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5939 19725 7379 19755 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5969 19695 7379 19725 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5999 19665 7379 19695 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6029 19635 7379 19665 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6059 19605 7379 19635 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6089 19575 7379 19605 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6119 19545 7379 19575 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6149 19515 7379 19545 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6179 19485 7379 19515 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6209 19455 7379 19485 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6239 19425 7379 19455 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6269 19395 7379 19425 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6299 19365 7379 19395 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6329 19335 7379 19365 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6359 19305 7379 19335 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6389 19275 7379 19305 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18598 5905 18620 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18568 5927 18598 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18538 5957 18568 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18508 5987 18538 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6389 18620 7379 19275 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4764 18493 6017 18508 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4779 18478 6032 18493 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6389 18598 7379 18620 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6367 18568 7379 18598 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6337 18538 7379 18568 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6307 18508 7379 18538 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6277 18478 7379 18508 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4789 18468 7379 18478 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4819 18438 7379 18468 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4849 18408 7379 18438 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4879 18378 7379 18408 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4909 18348 7379 18378 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4939 18318 7379 18348 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4969 18288 7379 18318 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4999 18258 7379 18288 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5029 18228 7379 18258 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5059 18198 7379 18228 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5089 18168 7379 18198 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5119 18138 7379 18168 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5149 18108 7379 18138 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5179 18078 7379 18108 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5179 0 7379 18078 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 99 0 4879 411 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 495 4879 499 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 183 481 4879 495 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 169 467 4879 481 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 155 453 4879 467 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 141 439 4879 453 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 127 425 4879 439 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 113 411 4879 425 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 499 4879 1719 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2475 5635 2480 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2461 5621 2475 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2447 5607 2461 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2433 5593 2447 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2419 5579 2433 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2405 5565 2419 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2391 5551 2405 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2377 5537 2391 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2363 5523 2377 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2349 5509 2363 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2335 5495 2349 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2321 5481 2335 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2307 5467 2321 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2293 5453 2307 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2279 5439 2293 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2265 5425 2279 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2251 5411 2265 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2237 5397 2251 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2223 5383 2237 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2209 5369 2223 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2195 5355 2209 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2181 5341 2195 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2167 5327 2181 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2153 5313 2167 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2139 5299 2153 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2125 5285 2139 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2111 5271 2125 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2097 5257 2111 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2083 5243 2097 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2069 5229 2083 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2055 5215 2069 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2041 5201 2055 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2027 5187 2041 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2013 5173 2027 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1999 5159 2013 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1985 5145 1999 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1971 5131 1985 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1957 5117 1971 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1943 5103 1957 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1929 5089 1943 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1915 5075 1929 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1901 5061 1915 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1887 5047 1901 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1873 5033 1887 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1859 5019 1873 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1845 5005 1859 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1831 4991 1845 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1817 4977 1831 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1803 4963 1817 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1789 4949 1803 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1775 4935 1789 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1761 4921 1775 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1747 4907 1761 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1733 4893 1747 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 1719 4879 1733 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 2480 7379 5140 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5854 3041 5863 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5840 3050 5854 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5826 3064 5840 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5812 3078 5826 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5798 3092 5812 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5784 3106 5798 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5770 3120 5784 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5756 3134 5770 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5742 3148 5756 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5728 3162 5742 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5714 3176 5728 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5700 3190 5714 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5686 3204 5700 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5672 3218 5686 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5658 3232 5672 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5644 3246 5658 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5630 3260 5644 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5616 3274 5630 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5602 3288 5616 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5588 3302 5602 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5574 3316 5588 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5560 3330 5574 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5546 3344 5560 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5532 3358 5546 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5518 3372 5532 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5504 3386 5518 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5490 3400 5504 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5476 3414 5490 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5462 3428 5476 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5448 3442 5462 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5434 3456 5448 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5420 3470 5434 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5406 3484 5420 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5392 3498 5406 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5378 3512 5392 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5364 3526 5378 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5350 3540 5364 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5336 3554 5350 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5322 3568 5336 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5308 3582 5322 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5294 3596 5308 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5280 3610 5294 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5266 3624 5280 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5252 3638 5266 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5238 3652 5252 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5224 3666 5238 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5210 3680 5224 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5196 3694 5210 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5182 3708 5196 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5168 3722 5182 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5154 3736 5168 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5140 3750 5154 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 5863 3041 7111 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7615 3545 7620 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7601 3531 7615 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7587 3517 7601 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7573 3503 7587 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7559 3489 7573 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7545 3475 7559 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7531 3461 7545 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7517 3447 7531 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7503 3433 7517 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7489 3419 7503 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7475 3405 7489 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7461 3391 7475 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7447 3377 7461 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7433 3363 7447 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7419 3349 7433 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7405 3335 7419 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7391 3321 7405 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7377 3307 7391 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7363 3293 7377 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7349 3279 7363 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7335 3265 7349 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7321 3251 7335 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7307 3237 7321 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7293 3223 7307 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7279 3209 7293 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7265 3195 7279 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7251 3181 7265 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7237 3167 7251 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7223 3153 7237 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7209 3139 7223 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7195 3125 7209 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7181 3111 7195 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7167 3097 7181 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7153 3083 7167 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7139 3069 7153 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7125 3055 7139 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7111 3041 7125 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10934 7223 11383 7442 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10766 7610 11383 7620 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10780 7596 11383 7610 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10794 7582 11383 7596 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10808 7568 11383 7582 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10822 7554 11383 7568 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10836 7540 11383 7554 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10850 7526 11383 7540 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10864 7512 11383 7526 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10878 7498 11383 7512 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10892 7484 11383 7498 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10906 7470 11383 7484 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10920 7456 11383 7470 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10934 7442 11383 7456 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7620 11383 7933 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8017 11290 8026 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8003 11299 8017 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7989 11313 8003 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7975 11327 7989 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7961 11341 7975 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7947 11355 7961 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 7933 11369 7947 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8600 2824 8613 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8586 2837 8600 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8572 2851 8586 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8558 2865 8572 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8544 2879 8558 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8530 2893 8544 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8516 2907 8530 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8502 2921 8516 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8488 2935 8502 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8474 2949 8488 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8460 2963 8474 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8446 2977 8460 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8432 2991 8446 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8418 3005 8432 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8404 3019 8418 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8390 3033 8404 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8376 3047 8390 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8362 3061 8376 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8348 3075 8362 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8334 3089 8348 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8320 3103 8334 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8306 3117 8320 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8292 3131 8306 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8278 3145 8292 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8264 3159 8278 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8250 3173 8264 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8236 3187 8250 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8222 3201 8236 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8208 3215 8222 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8194 3229 8208 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8180 3243 8194 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8166 3257 8180 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8152 3271 8166 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8138 3285 8152 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8124 3299 8138 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8110 3313 8124 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8096 3327 8110 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8082 3341 8096 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8068 3355 8082 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8054 3369 8068 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8040 3383 8054 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8026 3397 8040 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8613 2824 10843 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11543 3524 11556 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11529 3510 11543 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11515 3496 11529 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11501 3482 11515 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11487 3468 11501 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11473 3454 11487 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11459 3440 11473 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11445 3426 11459 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11431 3412 11445 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11417 3398 11431 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11403 3384 11417 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11389 3370 11403 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11375 3356 11389 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11361 3342 11375 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11347 3328 11361 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11333 3314 11347 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11319 3300 11333 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11305 3286 11319 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11291 3272 11305 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11277 3258 11291 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11263 3244 11277 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11249 3230 11263 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11235 3216 11249 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11221 3202 11235 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11207 3188 11221 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11193 3174 11207 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11179 3160 11193 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11165 3146 11179 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11151 3132 11165 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11137 3118 11151 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11123 3104 11137 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11109 3090 11123 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11095 3076 11109 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11081 3062 11095 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11067 3048 11081 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11053 3034 11067 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11039 3020 11053 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11025 3006 11039 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11011 2992 11025 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10997 2978 11011 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10983 2964 10997 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10969 2950 10983 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10955 2936 10969 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10941 2922 10955 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10927 2908 10941 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10913 2894 10927 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10899 2880 10913 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10885 2866 10899 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10871 2852 10885 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10857 2838 10871 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 10843 2824 10857 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 11556 11342 13296 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13996 2824 14005 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13982 2833 13996 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13968 2847 13982 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13954 2861 13968 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13940 2875 13954 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13926 2889 13940 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13912 2903 13926 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13898 2917 13912 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13884 2931 13898 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13870 2945 13884 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13856 2959 13870 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13842 2973 13856 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13828 2987 13842 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13814 3001 13828 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13800 3015 13814 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13786 3029 13800 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13772 3043 13786 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13758 3057 13772 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13744 3071 13758 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13730 3085 13744 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13716 3099 13730 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13702 3113 13716 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13688 3127 13702 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13674 3141 13688 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13660 3155 13674 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13646 3169 13660 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13632 3183 13646 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13618 3197 13632 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13604 3211 13618 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13590 3225 13604 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13576 3239 13590 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13562 3253 13576 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13548 3267 13562 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13534 3281 13548 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13520 3295 13534 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13506 3309 13520 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13492 3323 13506 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13478 3337 13492 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13464 3351 13478 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13450 3365 13464 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13436 3379 13450 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13422 3393 13436 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13408 3407 13422 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13394 3421 13408 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13380 3435 13394 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13366 3449 13380 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13352 3463 13366 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13338 3477 13352 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13324 3491 13338 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13310 3505 13324 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 13296 3519 13310 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 14005 2824 15448 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16148 3524 16156 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16134 3510 16148 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16120 3496 16134 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16106 3482 16120 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16092 3468 16106 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16078 3454 16092 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16064 3440 16078 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16050 3426 16064 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16036 3412 16050 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16022 3398 16036 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16008 3384 16022 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15994 3370 16008 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15980 3356 15994 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15966 3342 15980 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15952 3328 15966 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15938 3314 15952 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15924 3300 15938 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15910 3286 15924 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15896 3272 15910 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15882 3258 15896 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15868 3244 15882 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15854 3230 15868 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15840 3216 15854 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15826 3202 15840 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15812 3188 15826 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15798 3174 15812 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15784 3160 15798 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15770 3146 15784 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15756 3132 15770 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15742 3118 15756 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15728 3104 15742 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15714 3090 15728 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15700 3076 15714 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15686 3062 15700 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15672 3048 15686 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15658 3034 15672 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15644 3020 15658 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15630 3006 15644 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15616 2992 15630 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15602 2978 15616 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15588 2964 15602 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15574 2950 15588 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15560 2936 15574 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15546 2922 15560 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15532 2908 15546 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15518 2894 15532 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15504 2880 15518 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15490 2866 15504 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15476 2852 15490 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15462 2838 15476 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 15448 2824 15462 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 16156 11341 17896 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18596 2824 18605 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18582 2833 18596 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18568 2847 18582 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18554 2861 18568 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18540 2875 18554 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18526 2889 18540 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18512 2903 18526 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18498 2917 18512 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18484 2931 18498 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18470 2945 18484 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18456 2959 18470 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18442 2973 18456 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18428 2987 18442 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18414 3001 18428 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18400 3015 18414 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18386 3029 18400 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18372 3043 18386 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18358 3057 18372 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18344 3071 18358 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18330 3085 18344 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18316 3099 18330 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18302 3113 18316 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18288 3127 18302 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18274 3141 18288 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18260 3155 18274 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18246 3169 18260 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18232 3183 18246 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18218 3197 18232 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18204 3211 18218 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18190 3225 18204 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18176 3239 18190 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18162 3253 18176 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18148 3267 18162 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18134 3281 18148 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18120 3295 18134 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18106 3309 18120 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18092 3323 18106 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18078 3337 18092 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18064 3351 18078 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18050 3365 18064 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18036 3379 18050 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18022 3393 18036 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18008 3407 18022 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17994 3421 18008 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17980 3435 17994 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17966 3449 17980 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17952 3463 17966 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17938 3477 17952 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17924 3491 17938 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17910 3505 17924 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 17896 3519 17910 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 18605 2824 20048 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20748 3524 20756 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20734 3510 20748 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20720 3496 20734 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20706 3482 20720 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20692 3468 20706 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20678 3454 20692 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20664 3440 20678 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20650 3426 20664 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20636 3412 20650 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20622 3398 20636 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20608 3384 20622 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20594 3370 20608 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20580 3356 20594 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20566 3342 20580 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20552 3328 20566 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20538 3314 20552 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20524 3300 20538 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20510 3286 20524 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20496 3272 20510 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20482 3258 20496 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20468 3244 20482 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20454 3230 20468 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20440 3216 20454 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20426 3202 20440 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20412 3188 20426 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20398 3174 20412 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20384 3160 20398 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20370 3146 20384 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20356 3132 20370 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20342 3118 20356 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20328 3104 20342 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20314 3090 20328 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20300 3076 20314 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20286 3062 20300 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20272 3048 20286 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20258 3034 20272 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20244 3020 20258 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20230 3006 20244 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20216 2992 20230 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20202 2978 20216 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20188 2964 20202 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20174 2950 20188 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20160 2936 20174 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20146 2922 20160 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20132 2908 20146 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20118 2894 20132 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20104 2880 20118 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20090 2866 20104 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20076 2852 20090 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20062 2838 20076 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20048 2824 20062 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 20756 11341 22496 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23210 2824 23213 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23196 2827 23210 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23182 2841 23196 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23168 2855 23182 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23154 2869 23168 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23140 2883 23154 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23126 2897 23140 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23112 2911 23126 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23098 2925 23112 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23084 2939 23098 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23070 2953 23084 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23056 2967 23070 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23042 2981 23056 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23028 2995 23042 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23014 3009 23028 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23000 3023 23014 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22986 3037 23000 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22972 3051 22986 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22958 3065 22972 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22944 3079 22958 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22930 3093 22944 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22916 3107 22930 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22902 3121 22916 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22888 3135 22902 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22874 3149 22888 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22860 3163 22874 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22846 3177 22860 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22832 3191 22846 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22818 3205 22832 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22804 3219 22818 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22790 3233 22804 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22776 3247 22790 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22762 3261 22776 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22748 3275 22762 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22734 3289 22748 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22720 3303 22734 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22706 3317 22720 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22692 3331 22706 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22678 3345 22692 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22664 3359 22678 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22650 3373 22664 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22636 3387 22650 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22622 3401 22636 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22608 3415 22622 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22594 3429 22608 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22580 3443 22594 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22566 3457 22580 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22552 3471 22566 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22538 3485 22552 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22524 3499 22538 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22510 3513 22524 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 22496 3527 22510 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 23213 2824 24629 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25343 3538 25356 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25329 3524 25343 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25315 3510 25329 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25301 3496 25315 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25287 3482 25301 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25273 3468 25287 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25259 3454 25273 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25245 3440 25259 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25231 3426 25245 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25217 3412 25231 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25203 3398 25217 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25189 3384 25203 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25175 3370 25189 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25161 3356 25175 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25147 3342 25161 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25133 3328 25147 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25119 3314 25133 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25105 3300 25119 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25091 3286 25105 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25077 3272 25091 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25063 3258 25077 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25049 3244 25063 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25035 3230 25049 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25021 3216 25035 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25007 3202 25021 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24993 3188 25007 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24979 3174 24993 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24965 3160 24979 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24951 3146 24965 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24937 3132 24951 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24923 3118 24937 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24909 3104 24923 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24895 3090 24909 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24881 3076 24895 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24867 3062 24881 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24853 3048 24867 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24839 3034 24853 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24825 3020 24839 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24811 3006 24825 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24797 2992 24811 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24783 2978 24797 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24769 2964 24783 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24755 2950 24769 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24741 2936 24755 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24727 2922 24741 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24713 2908 24727 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24699 2894 24713 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24685 2880 24699 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24671 2866 24685 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24657 2852 24671 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24643 2838 24657 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 24629 2824 24643 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 25356 11341 27096 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27824 2824 27834 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27810 2834 27824 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27796 2848 27810 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27782 2862 27796 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27768 2876 27782 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27754 2890 27768 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27740 2904 27754 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27726 2918 27740 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27712 2932 27726 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27698 2946 27712 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27684 2960 27698 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27670 2974 27684 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27656 2988 27670 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27642 3002 27656 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27628 3016 27642 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27614 3030 27628 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27600 3044 27614 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27586 3058 27600 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27572 3072 27586 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27558 3086 27572 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27544 3100 27558 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27530 3114 27544 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27516 3128 27530 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27502 3142 27516 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27488 3156 27502 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27474 3170 27488 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27460 3184 27474 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27446 3198 27460 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27432 3212 27446 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27418 3226 27432 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27404 3240 27418 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27390 3254 27404 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27376 3268 27390 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27362 3282 27376 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27348 3296 27362 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27334 3310 27348 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27320 3324 27334 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27306 3338 27320 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27292 3352 27306 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27278 3366 27292 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27264 3380 27278 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27250 3394 27264 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27236 3408 27250 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27222 3422 27236 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27208 3436 27222 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27194 3450 27208 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27180 3464 27194 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27166 3478 27180 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27152 3492 27166 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27138 3506 27152 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27124 3520 27138 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27110 3534 27124 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27096 3548 27110 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 27834 2824 29243 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29943 3524 29956 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29929 3510 29943 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29915 3496 29929 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29901 3482 29915 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29887 3468 29901 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29873 3454 29887 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29859 3440 29873 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29845 3426 29859 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29831 3412 29845 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29817 3398 29831 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29803 3384 29817 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29789 3370 29803 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29775 3356 29789 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29761 3342 29775 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29747 3328 29761 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29733 3314 29747 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29719 3300 29733 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29705 3286 29719 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29691 3272 29705 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29677 3258 29691 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29663 3244 29677 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29649 3230 29663 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29635 3216 29649 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29621 3202 29635 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29607 3188 29621 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29593 3174 29607 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29579 3160 29593 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29565 3146 29579 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29551 3132 29565 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29537 3118 29551 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29523 3104 29537 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29509 3090 29523 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29495 3076 29509 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29481 3062 29495 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29467 3048 29481 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29453 3034 29467 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29439 3020 29453 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29425 3006 29439 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29411 2992 29425 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29397 2978 29411 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29383 2964 29397 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29369 2950 29383 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29355 2936 29369 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29341 2922 29355 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29327 2908 29341 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29313 2894 29327 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29299 2880 29313 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29285 2866 29299 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29271 2852 29285 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29257 2838 29271 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29243 2824 29257 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 29956 11341 31696 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32410 2824 32416 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32396 2830 32410 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32382 2844 32396 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32368 2858 32382 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32354 2872 32368 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32340 2886 32354 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32326 2900 32340 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32312 2914 32326 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32298 2928 32312 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32284 2942 32298 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32270 2956 32284 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32256 2970 32270 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32242 2984 32256 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32228 2998 32242 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32214 3012 32228 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32200 3026 32214 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32186 3040 32200 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32172 3054 32186 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32158 3068 32172 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32144 3082 32158 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32130 3096 32144 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32116 3110 32130 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32102 3124 32116 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32088 3138 32102 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32074 3152 32088 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32060 3166 32074 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32046 3180 32060 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32032 3194 32046 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32018 3208 32032 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32004 3222 32018 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31990 3236 32004 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31976 3250 31990 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31962 3264 31976 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31948 3278 31962 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31934 3292 31948 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31920 3306 31934 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31906 3320 31920 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31892 3334 31906 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31878 3348 31892 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31864 3362 31878 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31850 3376 31864 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31836 3390 31850 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31822 3404 31836 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31808 3418 31822 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31794 3432 31808 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31780 3446 31794 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31766 3460 31780 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31752 3474 31766 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31738 3488 31752 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31724 3502 31738 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31710 3516 31724 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 31696 3530 31710 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 32416 2824 33844 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34544 3524 34556 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34530 3510 34544 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34516 3496 34530 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34502 3482 34516 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34488 3468 34502 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34474 3454 34488 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34460 3440 34474 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34446 3426 34460 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34432 3412 34446 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34418 3398 34432 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34404 3384 34418 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34390 3370 34404 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34376 3356 34390 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34362 3342 34376 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34348 3328 34362 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34334 3314 34348 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34320 3300 34334 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34306 3286 34320 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34292 3272 34306 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34278 3258 34292 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34264 3244 34278 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34250 3230 34264 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34236 3216 34250 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34222 3202 34236 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34208 3188 34222 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34194 3174 34208 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34180 3160 34194 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34166 3146 34180 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34152 3132 34166 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34138 3118 34152 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34124 3104 34138 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34110 3090 34124 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34096 3076 34110 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34082 3062 34096 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34068 3048 34082 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34054 3034 34068 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34040 3020 34054 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34026 3006 34040 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34012 2992 34026 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33998 2978 34012 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33984 2964 33998 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33970 2950 33984 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33956 2936 33970 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33942 2922 33956 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33928 2908 33942 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33914 2894 33928 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33900 2880 33914 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33886 2866 33900 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33872 2852 33886 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33858 2838 33872 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 33844 2824 33858 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 34556 11592 36296 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36758 3064 36771 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36744 3077 36758 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36730 3091 36744 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36716 3105 36730 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36702 3119 36716 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36688 3133 36702 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36674 3147 36688 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36660 3161 36674 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36646 3175 36660 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36632 3189 36646 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36618 3203 36632 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36604 3217 36618 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36590 3231 36604 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36576 3245 36590 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36562 3259 36576 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36548 3273 36562 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36534 3287 36548 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36520 3301 36534 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36506 3315 36520 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36492 3329 36506 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36478 3343 36492 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36464 3357 36478 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36450 3371 36464 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36436 3385 36450 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36422 3399 36436 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36408 3413 36422 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36394 3427 36408 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36380 3441 36394 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36366 3455 36380 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36352 3469 36366 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36338 3483 36352 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36324 3497 36338 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36310 3511 36324 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36296 3525 36310 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36771 3064 36781 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37005 2824 37011 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36991 2830 37005 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36977 2844 36991 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36963 2858 36977 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36949 2872 36963 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36935 2886 36949 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36921 2900 36935 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36907 2914 36921 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36893 2928 36907 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36879 2942 36893 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36865 2956 36879 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36851 2970 36865 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36837 2984 36851 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36823 2998 36837 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36809 3012 36823 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36795 3026 36809 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 36781 3040 36795 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37011 2824 37917 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38099 3006 38112 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38085 2992 38099 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38071 2978 38085 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38057 2964 38071 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38043 2950 38057 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38029 2936 38043 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38015 2922 38029 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38001 2908 38015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37987 2894 38001 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37973 2880 37987 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37959 2866 37973 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37945 2852 37959 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37931 2838 37945 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 37917 2824 37931 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 38112 13440 39015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 8571 22124 9771 34092 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10657 22088 11857 33827 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 35045 12298 38008 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 35024 12277 35045 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34994 12247 35024 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34964 12217 34994 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34934 12187 34964 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34904 12157 34934 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34874 12127 34904 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34844 12097 34874 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34814 12067 34844 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34784 12037 34814 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34754 12007 34784 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34724 11977 34754 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34694 11947 34724 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34664 11917 34694 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34634 11887 34664 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34604 11857 34634 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7593 35070 9771 38004 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9955 34529 11857 34604 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7611 35052 9771 35070 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7641 35022 9771 35052 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7671 34992 9771 35022 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7701 34962 9771 34992 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7731 34932 9771 34962 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7761 34902 9771 34932 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7791 34872 9771 34902 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7821 34842 9771 34872 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7851 34812 9771 34842 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7881 34782 9771 34812 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7911 34752 9771 34782 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7941 34722 9771 34752 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7971 34692 9771 34722 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8001 34662 9771 34692 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8031 34632 9771 34662 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8061 34602 9771 34632 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8091 34572 9771 34602 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8121 34542 9771 34572 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8151 34512 9771 34542 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8181 34482 9771 34512 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8211 34452 9771 34482 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8241 34422 9771 34452 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8271 34392 9771 34422 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8301 34362 9771 34392 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8331 34332 9771 34362 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8361 34302 9771 34332 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8391 34272 9771 34302 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8421 34242 9771 34272 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8451 34212 9771 34242 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8481 34182 9771 34212 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8511 34152 9771 34182 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8541 34122 9771 34152 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8571 34092 9771 34122 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9967 34517 11857 34529 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9997 34487 11857 34517 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10027 34457 11857 34487 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10057 34427 11857 34457 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10087 34397 11857 34427 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10117 34367 11857 34397 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10147 34337 11857 34367 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10177 34307 11857 34337 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10207 34277 11857 34307 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10237 34247 11857 34277 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10267 34217 11857 34247 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10297 34187 11857 34217 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10327 34157 11857 34187 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10357 34127 11857 34157 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10387 34097 11857 34127 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10417 34067 11857 34097 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10447 34037 11857 34067 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10477 34007 11857 34037 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10507 33977 11857 34007 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10537 33947 11857 33977 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10567 33917 11857 33947 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10597 33887 11857 33917 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10627 33857 11857 33887 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10657 33827 11857 33857 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8571 22110 9771 22124 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8557 22080 9771 22110 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8527 22050 9771 22080 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8497 22020 9771 22050 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8467 21990 9771 22020 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8437 21960 9771 21990 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8407 21930 9771 21960 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8377 21900 9771 21930 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8347 21870 9771 21900 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8317 21840 9771 21870 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8287 21810 9771 21840 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8257 21780 9771 21810 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8227 21750 9771 21780 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8197 21720 9771 21750 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8167 21690 9771 21720 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8137 21660 9771 21690 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8107 21630 9771 21660 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10657 22072 11857 22088 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10641 22042 11857 22072 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10611 22012 11857 22042 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10581 21982 11857 22012 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10551 21952 11857 21982 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10521 21922 11857 21952 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10491 21892 11857 21922 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10461 21862 11857 21892 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10431 21832 11857 21862 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10401 21802 11857 21832 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10371 21772 11857 21802 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10341 21742 11857 21772 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10311 21712 11857 21742 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10281 21682 11857 21712 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10251 21652 11857 21682 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10221 21622 11857 21652 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10191 21592 11857 21622 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8077 21611 9752 21630 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8058 21581 9722 21611 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8028 21551 9692 21581 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7998 21521 9662 21551 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7968 21491 9632 21521 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7938 21461 9602 21491 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7908 21431 9572 21461 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7878 21401 9542 21431 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7848 21371 9512 21401 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7818 21341 9482 21371 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7788 21311 9452 21341 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7758 21281 9422 21311 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7728 21251 9392 21281 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7698 21221 9362 21251 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7668 21191 9332 21221 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7638 21161 9302 21191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7608 21131 9272 21161 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10161 21581 11846 21592 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10150 21551 11816 21581 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10120 21521 11786 21551 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10090 21491 11756 21521 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10060 21461 11726 21491 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10030 21431 11696 21461 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10000 21401 11666 21431 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9970 21371 11636 21401 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9940 21341 11606 21371 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9910 21311 11576 21341 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9880 21281 11546 21311 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9850 21251 11516 21281 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9820 21221 11486 21251 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9790 21191 11456 21221 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9760 21161 11426 21191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9730 21131 11396 21161 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9700 21101 11366 21131 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9670 21071 11336 21101 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9640 21041 11306 21071 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9610 21011 11276 21041 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9580 20981 11246 21011 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9550 20951 11216 20981 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9520 20921 11186 20951 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9490 20891 11156 20921 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9460 20861 11126 20891 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9430 20831 11096 20861 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9400 20801 11066 20831 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9370 20771 11036 20801 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9340 20741 11006 20771 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9310 20711 10976 20741 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9280 20681 10946 20711 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9250 20651 10916 20681 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9220 20621 10886 20651 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9190 20591 10856 20621 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9160 20561 10826 20591 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9130 20531 10796 20561 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9100 20501 10766 20531 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21117 9258 21131 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21087 9228 21117 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21057 9198 21087 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21027 9168 21057 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20997 9138 21027 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20967 9108 20997 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20937 9078 20967 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20907 9048 20937 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20877 9018 20907 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20847 8988 20877 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20817 8958 20847 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20787 8928 20817 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20757 8898 20787 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20727 8868 20757 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20697 8838 20727 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20667 8808 20697 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20637 8778 20667 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20607 8748 20637 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20577 8718 20607 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20547 8688 20577 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20517 8658 20547 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20487 8628 20517 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20457 8598 20487 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20427 8568 20457 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20057 8568 20427 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20051 8568 20057 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20021 8574 20051 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19991 8604 20021 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19961 8634 19991 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19931 8664 19961 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19901 8694 19931 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19660 10208 19901 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8967 19922 10208 19943 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8946 19901 10208 19922 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20033 10298 20046 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9057 20003 10268 20033 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9027 19973 10238 20003 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8997 19943 10208 19973 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20496 10761 20501 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20466 10731 20496 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20436 10701 20466 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20406 10671 20436 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20376 10641 20406 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20346 10611 20376 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20316 10581 20346 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20286 10551 20316 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20256 10521 20286 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20226 10491 20256 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20196 10461 20226 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20166 10431 20196 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20136 10401 20166 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20106 10371 20136 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20076 10341 20106 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20046 10311 20076 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19650 10198 19660 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19620 10168 19650 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19590 10138 19620 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19560 10108 19590 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19530 10078 19560 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19500 10048 19530 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19470 10018 19500 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19440 9988 19470 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19410 9958 19440 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19380 9928 19410 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19350 9898 19380 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19320 9868 19350 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19290 9838 19320 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19260 9808 19290 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 19230 9778 19260 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 0 9778 19230 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10078 0 14858 1725 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9350 2453 14858 2459 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9364 2439 14858 2453 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9378 2425 14858 2439 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9392 2411 14858 2425 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9406 2397 14858 2411 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9420 2383 14858 2397 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9434 2369 14858 2383 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9448 2355 14858 2369 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9462 2341 14858 2355 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9476 2327 14858 2341 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9490 2313 14858 2327 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9504 2299 14858 2313 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9518 2285 14858 2299 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9532 2271 14858 2285 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9546 2257 14858 2271 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9560 2243 14858 2257 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9574 2229 14858 2243 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9588 2215 14858 2229 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9602 2201 14858 2215 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9616 2187 14858 2201 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9630 2173 14858 2187 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9644 2159 14858 2173 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9658 2145 14858 2159 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9672 2131 14858 2145 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9686 2117 14858 2131 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9700 2103 14858 2117 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9714 2089 14858 2103 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9728 2075 14858 2089 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9742 2061 14858 2075 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9756 2047 14858 2061 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9770 2033 14858 2047 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9784 2019 14858 2033 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9798 2005 14858 2019 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9812 1991 14858 2005 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9826 1977 14858 1991 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9840 1963 14858 1977 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9854 1949 14858 1963 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9868 1935 14858 1949 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9882 1921 14858 1935 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9896 1907 14858 1921 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9910 1893 14858 1907 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9924 1879 14858 1893 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9938 1865 14858 1879 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9952 1851 14858 1865 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9966 1837 14858 1851 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9980 1823 14858 1837 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 9994 1809 14858 1823 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10008 1795 14858 1809 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10022 1781 14858 1795 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10036 1767 14858 1781 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10050 1753 14858 1767 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10064 1739 14858 1753 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10078 1725 14858 1739 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 7578 2459 14858 5132 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11177 5132 14858 5146 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11191 5146 14858 5160 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11205 5160 14858 5174 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11219 5174 14858 5188 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11233 5188 14858 5202 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11247 5202 14858 5216 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11261 5216 14858 5230 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11275 5230 14858 5244 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11289 5244 14858 5258 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11303 5258 14858 5272 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11317 5272 14858 5286 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11331 5286 14858 5300 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11345 5300 14858 5314 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11359 5314 14858 5328 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11373 5328 14858 5342 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11387 5342 14858 5356 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11401 5356 14858 5370 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11415 5370 14858 5384 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11429 5384 14858 5398 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11443 5398 14858 5412 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11457 5412 14858 5426 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11471 5426 14858 5440 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11485 5440 14858 5454 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11499 5454 14858 5468 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11513 5468 14858 5482 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11527 5482 14858 5496 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11541 5496 14858 5510 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11555 5510 14858 5524 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11569 5524 14858 5538 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11583 5538 14858 5552 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11597 5552 14858 5566 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11611 5566 14858 5580 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11625 5580 14858 5594 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11639 5594 14858 5608 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11653 5608 14858 5622 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11667 5622 14858 5636 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11681 5636 14858 5650 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11695 5650 14858 5664 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11709 5664 14858 5678 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11723 5678 14858 5692 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11737 5692 14858 5706 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11751 5706 14858 5720 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11765 5720 14858 5734 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11779 5734 14858 5748 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11793 5748 14858 5762 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11807 5762 14858 5776 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11821 5776 14858 5790 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11835 5790 14858 5804 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11849 5804 14858 5818 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11863 5818 14858 5832 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11877 5832 14858 5846 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11891 5846 14858 5860 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11905 5860 14858 5874 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11919 5874 14858 5888 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11933 5888 14858 5902 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11947 5902 14858 5916 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11961 5916 14858 5930 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11975 5930 14858 5944 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11989 5944 14858 5958 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12003 5958 14858 5972 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12017 5972 14858 5986 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12031 5986 14858 6000 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12045 6000 14858 6014 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12059 6014 14858 6028 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12073 6028 14858 6042 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12087 6042 14858 6056 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12101 6056 14858 6070 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12115 6070 14858 6084 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12129 6084 14858 6098 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12143 6098 14858 6112 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12157 6112 14858 6126 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12171 6126 14858 6140 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12185 6140 14858 6154 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12199 6154 14858 6168 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12213 6168 14858 6182 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 6182 14858 6191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 6191 14858 8764 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11508 9478 14858 9491 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11522 9464 14858 9478 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11536 9450 14858 9464 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11550 9436 14858 9450 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11564 9422 14858 9436 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11578 9408 14858 9422 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11592 9394 14858 9408 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11606 9380 14858 9394 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11620 9366 14858 9380 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11634 9352 14858 9366 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11648 9338 14858 9352 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11662 9324 14858 9338 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11676 9310 14858 9324 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11690 9296 14858 9310 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11704 9282 14858 9296 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11718 9268 14858 9282 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11732 9254 14858 9268 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 9240 14858 9254 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 9226 14858 9240 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 9212 14858 9226 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 9198 14858 9212 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 9184 14858 9198 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 9170 14858 9184 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 9156 14858 9170 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 9142 14858 9156 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 9128 14858 9142 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 9114 14858 9128 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 9100 14858 9114 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 9086 14858 9100 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 9072 14858 9086 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 9058 14858 9072 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 9044 14858 9058 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 9030 14858 9044 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 9016 14858 9030 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 9002 14858 9016 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 8988 14858 9002 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 8974 14858 8988 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 8960 14858 8974 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 8946 14858 8960 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 8932 14858 8946 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 8918 14858 8932 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 8904 14858 8918 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 8890 14858 8904 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 8876 14858 8890 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 8862 14858 8876 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 8848 14858 8862 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 8834 14858 8848 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 8820 14858 8834 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 8806 14858 8820 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 8792 14858 8806 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 8778 14858 8792 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 8764 14858 8778 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3361 9491 14858 10953 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3770 11219 14858 11231 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3758 11205 14858 11219 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3744 11191 14858 11205 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3730 11177 14858 11191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3716 11163 14858 11177 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3702 11149 14858 11163 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3688 11135 14858 11149 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3674 11121 14858 11135 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3660 11107 14858 11121 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3646 11093 14858 11107 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3632 11079 14858 11093 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3618 11065 14858 11079 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3604 11051 14858 11065 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3590 11037 14858 11051 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3576 11023 14858 11037 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3562 11009 14858 11023 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3548 10995 14858 11009 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3534 10981 14858 10995 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3520 10967 14858 10981 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3506 10953 14858 10967 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 11945 14858 11948 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12219 11931 14858 11945 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12205 11917 14858 11931 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12191 11903 14858 11917 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12177 11889 14858 11903 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12163 11875 14858 11889 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12149 11861 14858 11875 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12135 11847 14858 11861 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12121 11833 14858 11847 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12107 11819 14858 11833 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12093 11805 14858 11819 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12079 11791 14858 11805 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12065 11777 14858 11791 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12051 11763 14858 11777 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12037 11749 14858 11763 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12023 11735 14858 11749 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12009 11721 14858 11735 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11995 11707 14858 11721 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11981 11693 14858 11707 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11967 11679 14858 11693 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11953 11665 14858 11679 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11939 11651 14858 11665 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11925 11637 14858 11651 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11911 11623 14858 11637 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11897 11609 14858 11623 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11883 11595 14858 11609 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11869 11581 14858 11595 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11855 11567 14858 11581 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11841 11553 14858 11567 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11827 11539 14858 11553 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11813 11525 14858 11539 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11799 11511 14858 11525 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11785 11497 14858 11511 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11771 11483 14858 11497 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11757 11469 14858 11483 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11743 11455 14858 11469 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11729 11441 14858 11455 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11715 11427 14858 11441 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11701 11413 14858 11427 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11687 11399 14858 11413 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11673 11385 14858 11399 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11659 11371 14858 11385 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11645 11357 14858 11371 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11631 11343 14858 11357 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11617 11329 14858 11343 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11603 11315 14858 11329 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11589 11301 14858 11315 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11575 11287 14858 11301 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11561 11273 14858 11287 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11547 11259 14858 11273 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11533 11245 14858 11259 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11519 11231 14858 11245 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 11948 14858 13370 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11508 14084 14858 14091 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11522 14070 14858 14084 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11536 14056 14858 14070 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11550 14042 14858 14056 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11564 14028 14858 14042 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11578 14014 14858 14028 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11592 14000 14858 14014 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11606 13986 14858 14000 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11620 13972 14858 13986 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11634 13958 14858 13972 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11648 13944 14858 13958 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11662 13930 14858 13944 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11676 13916 14858 13930 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11690 13902 14858 13916 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11704 13888 14858 13902 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11718 13874 14858 13888 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11732 13860 14858 13874 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 13846 14858 13860 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 13832 14858 13846 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 13818 14858 13832 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 13804 14858 13818 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 13790 14858 13804 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 13776 14858 13790 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 13762 14858 13776 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 13748 14858 13762 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 13734 14858 13748 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 13720 14858 13734 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 13706 14858 13720 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 13692 14858 13706 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 13678 14858 13692 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 13664 14858 13678 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 13650 14858 13664 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 13636 14858 13650 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 13622 14858 13636 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 13608 14858 13622 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 13594 14858 13608 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 13580 14858 13594 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 13566 14858 13580 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 13552 14858 13566 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 13538 14858 13552 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 13524 14858 13538 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 13510 14858 13524 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 13496 14858 13510 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 13482 14858 13496 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 13468 14858 13482 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 13454 14858 13468 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 13440 14858 13454 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 13426 14858 13440 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 13412 14858 13426 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 13398 14858 13412 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 13384 14858 13398 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 13370 14858 13384 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4964 14091 14858 14597 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4768 14793 14858 14798 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4782 14779 14858 14793 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4796 14765 14858 14779 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4810 14751 14858 14765 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4824 14737 14858 14751 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4838 14723 14858 14737 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4852 14709 14858 14723 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4866 14695 14858 14709 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4880 14681 14858 14695 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4894 14667 14858 14681 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4908 14653 14858 14667 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4922 14639 14858 14653 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4936 14625 14858 14639 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4950 14611 14858 14625 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4964 14597 14858 14611 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3682 14798 14858 14916 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4964 15112 14858 15123 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4953 15098 14858 15112 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4939 15084 14858 15098 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4925 15070 14858 15084 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4911 15056 14858 15070 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4897 15042 14858 15056 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4883 15028 14858 15042 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4869 15014 14858 15028 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4855 15000 14858 15014 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4841 14986 14858 15000 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4827 14972 14858 14986 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4813 14958 14858 14972 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4799 14944 14858 14958 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4785 14930 14858 14944 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4771 14916 14858 14930 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4964 15123 14858 15831 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 16531 14858 16542 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12211 16517 14858 16531 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12197 16503 14858 16517 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12183 16489 14858 16503 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12169 16475 14858 16489 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12155 16461 14858 16475 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12141 16447 14858 16461 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12127 16433 14858 16447 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12113 16419 14858 16433 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12099 16405 14858 16419 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12085 16391 14858 16405 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12071 16377 14858 16391 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12057 16363 14858 16377 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12043 16349 14858 16363 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12029 16335 14858 16349 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12015 16321 14858 16335 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12001 16307 14858 16321 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11987 16293 14858 16307 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11973 16279 14858 16293 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11959 16265 14858 16279 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11945 16251 14858 16265 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11931 16237 14858 16251 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11917 16223 14858 16237 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11903 16209 14858 16223 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11889 16195 14858 16209 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11875 16181 14858 16195 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11861 16167 14858 16181 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11847 16153 14858 16167 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11833 16139 14858 16153 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11819 16125 14858 16139 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11805 16111 14858 16125 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11791 16097 14858 16111 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11777 16083 14858 16097 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11763 16069 14858 16083 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11749 16055 14858 16069 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11735 16041 14858 16055 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11721 16027 14858 16041 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11707 16013 14858 16027 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11693 15999 14858 16013 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11679 15985 14858 15999 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11665 15971 14858 15985 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11651 15957 14858 15971 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11637 15943 14858 15957 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11623 15929 14858 15943 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11609 15915 14858 15929 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11595 15901 14858 15915 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11581 15887 14858 15901 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11567 15873 14858 15887 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11553 15859 14858 15873 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11539 15845 14858 15859 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11525 15831 14858 15845 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 16542 14858 17982 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11522 18682 14858 18691 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11536 18668 14858 18682 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11550 18654 14858 18668 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11564 18640 14858 18654 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11578 18626 14858 18640 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11592 18612 14858 18626 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11606 18598 14858 18612 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11620 18584 14858 18598 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11634 18570 14858 18584 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11648 18556 14858 18570 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11662 18542 14858 18556 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11676 18528 14858 18542 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11690 18514 14858 18528 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11704 18500 14858 18514 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11718 18486 14858 18500 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11732 18472 14858 18486 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 18458 14858 18472 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 18444 14858 18458 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 18430 14858 18444 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 18416 14858 18430 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 18402 14858 18416 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 18388 14858 18402 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 18374 14858 18388 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 18360 14858 18374 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 18346 14858 18360 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 18332 14858 18346 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 18318 14858 18332 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 18304 14858 18318 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 18290 14858 18304 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 18276 14858 18290 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 18262 14858 18276 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 18248 14858 18262 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 18234 14858 18248 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 18220 14858 18234 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 18206 14858 18220 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 18192 14858 18206 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 18178 14858 18192 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 18164 14858 18178 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 18150 14858 18164 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 18136 14858 18150 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 18122 14858 18136 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 18108 14858 18122 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 18094 14858 18108 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 18080 14858 18094 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 18066 14858 18080 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 18052 14858 18066 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 18038 14858 18052 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 18024 14858 18038 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 18010 14858 18024 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 17996 14858 18010 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 17982 14858 17996 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4964 18691 14858 20431 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 21131 14858 21142 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12211 21117 14858 21131 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12197 21103 14858 21117 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12183 21089 14858 21103 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12169 21075 14858 21089 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12155 21061 14858 21075 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12141 21047 14858 21061 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12127 21033 14858 21047 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12113 21019 14858 21033 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12099 21005 14858 21019 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12085 20991 14858 21005 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12071 20977 14858 20991 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12057 20963 14858 20977 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12043 20949 14858 20963 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12029 20935 14858 20949 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12015 20921 14858 20935 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12001 20907 14858 20921 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11987 20893 14858 20907 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11973 20879 14858 20893 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11959 20865 14858 20879 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11945 20851 14858 20865 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11931 20837 14858 20851 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11917 20823 14858 20837 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11903 20809 14858 20823 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11889 20795 14858 20809 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11875 20781 14858 20795 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11861 20767 14858 20781 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11847 20753 14858 20767 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11833 20739 14858 20753 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11819 20725 14858 20739 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11805 20711 14858 20725 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11791 20697 14858 20711 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11777 20683 14858 20697 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11763 20669 14858 20683 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11749 20655 14858 20669 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11735 20641 14858 20655 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11721 20627 14858 20641 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11707 20613 14858 20627 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11693 20599 14858 20613 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11679 20585 14858 20599 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11665 20571 14858 20585 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11651 20557 14858 20571 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11637 20543 14858 20557 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11623 20529 14858 20543 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11609 20515 14858 20529 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11595 20501 14858 20515 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11581 20487 14858 20501 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11567 20473 14858 20487 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11553 20459 14858 20473 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11539 20445 14858 20459 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11525 20431 14858 20445 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 21142 14858 22564 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11508 23278 14858 23291 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11522 23264 14858 23278 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11536 23250 14858 23264 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11550 23236 14858 23250 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11564 23222 14858 23236 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11578 23208 14858 23222 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11592 23194 14858 23208 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11606 23180 14858 23194 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11620 23166 14858 23180 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11634 23152 14858 23166 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11648 23138 14858 23152 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11662 23124 14858 23138 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11676 23110 14858 23124 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11690 23096 14858 23110 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11704 23082 14858 23096 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11718 23068 14858 23082 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11732 23054 14858 23068 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 23040 14858 23054 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 23026 14858 23040 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 23012 14858 23026 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 22998 14858 23012 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 22984 14858 22998 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 22970 14858 22984 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 22956 14858 22970 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 22942 14858 22956 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 22928 14858 22942 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 22914 14858 22928 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 22900 14858 22914 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 22886 14858 22900 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 22872 14858 22886 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 22858 14858 22872 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 22844 14858 22858 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 22830 14858 22844 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 22816 14858 22830 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 22802 14858 22816 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 22788 14858 22802 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 22774 14858 22788 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 22760 14858 22774 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 22746 14858 22760 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 22732 14858 22746 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 22718 14858 22732 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 22704 14858 22718 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 22690 14858 22704 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 22676 14858 22690 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 22662 14858 22676 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 22648 14858 22662 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 22634 14858 22648 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 22620 14858 22634 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 22606 14858 22620 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 22592 14858 22606 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 22578 14858 22592 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 22564 14858 22578 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 4964 23291 14858 25031 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 25731 14858 25742 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12211 25717 14858 25731 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12197 25703 14858 25717 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12183 25689 14858 25703 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12169 25675 14858 25689 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12155 25661 14858 25675 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12141 25647 14858 25661 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12127 25633 14858 25647 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12113 25619 14858 25633 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12099 25605 14858 25619 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12085 25591 14858 25605 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12071 25577 14858 25591 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12057 25563 14858 25577 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12043 25549 14858 25563 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12029 25535 14858 25549 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12015 25521 14858 25535 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12001 25507 14858 25521 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11987 25493 14858 25507 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11973 25479 14858 25493 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11959 25465 14858 25479 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11945 25451 14858 25465 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11931 25437 14858 25451 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11917 25423 14858 25437 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11903 25409 14858 25423 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11889 25395 14858 25409 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11875 25381 14858 25395 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11861 25367 14858 25381 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11847 25353 14858 25367 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11833 25339 14858 25353 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11819 25325 14858 25339 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11805 25311 14858 25325 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11791 25297 14858 25311 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11777 25283 14858 25297 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11763 25269 14858 25283 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11749 25255 14858 25269 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11735 25241 14858 25255 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11721 25227 14858 25241 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11707 25213 14858 25227 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11693 25199 14858 25213 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11679 25185 14858 25199 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11665 25171 14858 25185 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11651 25157 14858 25171 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11637 25143 14858 25157 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11623 25129 14858 25143 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11609 25115 14858 25129 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11595 25101 14858 25115 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11581 25087 14858 25101 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11567 25073 14858 25087 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11553 25059 14858 25073 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11539 25045 14858 25059 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11525 25031 14858 25045 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 25742 14858 27171 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11508 27885 14858 27891 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11522 27871 14858 27885 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11536 27857 14858 27871 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11550 27843 14858 27857 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11564 27829 14858 27843 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11578 27815 14858 27829 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11592 27801 14858 27815 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11606 27787 14858 27801 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11620 27773 14858 27787 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11634 27759 14858 27773 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11648 27745 14858 27759 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11662 27731 14858 27745 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11676 27717 14858 27731 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11690 27703 14858 27717 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11704 27689 14858 27703 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11718 27675 14858 27689 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11732 27661 14858 27675 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 27647 14858 27661 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 27633 14858 27647 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 27619 14858 27633 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 27605 14858 27619 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 27591 14858 27605 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 27577 14858 27591 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 27563 14858 27577 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 27549 14858 27563 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 27535 14858 27549 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 27521 14858 27535 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 27507 14858 27521 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 27493 14858 27507 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 27479 14858 27493 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 27465 14858 27479 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 27451 14858 27465 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 27437 14858 27451 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 27423 14858 27437 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 27409 14858 27423 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 27395 14858 27409 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 27381 14858 27395 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 27367 14858 27381 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 27353 14858 27367 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 27339 14858 27353 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 27325 14858 27339 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 27311 14858 27325 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 27297 14858 27311 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 27283 14858 27297 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 27269 14858 27283 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 27255 14858 27269 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 27241 14858 27255 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 27227 14858 27241 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 27213 14858 27227 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 27199 14858 27213 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 27185 14858 27199 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 27171 14858 27185 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3361 27891 14858 29342 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3650 29622 14858 29631 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3641 29608 14858 29622 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3627 29594 14858 29608 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3613 29580 14858 29594 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3599 29566 14858 29580 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3585 29552 14858 29566 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3571 29538 14858 29552 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3557 29524 14858 29538 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3543 29510 14858 29524 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3529 29496 14858 29510 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3515 29482 14858 29496 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3501 29468 14858 29482 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3487 29454 14858 29468 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3473 29440 14858 29454 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3459 29426 14858 29440 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3445 29412 14858 29426 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3431 29398 14858 29412 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3417 29384 14858 29398 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3403 29370 14858 29384 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3389 29356 14858 29370 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3375 29342 14858 29356 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 30345 14858 30356 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12211 30331 14858 30345 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12197 30317 14858 30331 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12183 30303 14858 30317 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12169 30289 14858 30303 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12155 30275 14858 30289 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12141 30261 14858 30275 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12127 30247 14858 30261 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12113 30233 14858 30247 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12099 30219 14858 30233 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12085 30205 14858 30219 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12071 30191 14858 30205 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12057 30177 14858 30191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12043 30163 14858 30177 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12029 30149 14858 30163 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12015 30135 14858 30149 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12001 30121 14858 30135 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11987 30107 14858 30121 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11973 30093 14858 30107 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11959 30079 14858 30093 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11945 30065 14858 30079 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11931 30051 14858 30065 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11917 30037 14858 30051 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11903 30023 14858 30037 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11889 30009 14858 30023 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11875 29995 14858 30009 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11861 29981 14858 29995 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11847 29967 14858 29981 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11833 29953 14858 29967 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11819 29939 14858 29953 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11805 29925 14858 29939 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11791 29911 14858 29925 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11777 29897 14858 29911 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11763 29883 14858 29897 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11749 29869 14858 29883 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11735 29855 14858 29869 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11721 29841 14858 29855 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11707 29827 14858 29841 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11693 29813 14858 29827 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11679 29799 14858 29813 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11665 29785 14858 29799 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11651 29771 14858 29785 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11637 29757 14858 29771 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11623 29743 14858 29757 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11609 29729 14858 29743 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11595 29715 14858 29729 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11581 29701 14858 29715 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11567 29687 14858 29701 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11553 29673 14858 29687 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11539 29659 14858 29673 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11525 29645 14858 29659 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11511 29631 14858 29645 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 30356 14858 31774 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11508 32488 14858 32491 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11522 32474 14858 32488 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11536 32460 14858 32474 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11550 32446 14858 32460 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11564 32432 14858 32446 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11578 32418 14858 32432 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11592 32404 14858 32418 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11606 32390 14858 32404 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11620 32376 14858 32390 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11634 32362 14858 32376 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11648 32348 14858 32362 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11662 32334 14858 32348 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11676 32320 14858 32334 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11690 32306 14858 32320 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11704 32292 14858 32306 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11718 32278 14858 32292 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11732 32264 14858 32278 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 32250 14858 32264 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 32236 14858 32250 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 32222 14858 32236 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 32208 14858 32222 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 32194 14858 32208 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 32180 14858 32194 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 32166 14858 32180 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 32152 14858 32166 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 32138 14858 32152 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 32124 14858 32138 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 32110 14858 32124 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 32096 14858 32110 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 32082 14858 32096 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 32068 14858 32082 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 32054 14858 32068 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 32040 14858 32054 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 32026 14858 32040 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 32012 14858 32026 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 31998 14858 32012 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 31984 14858 31998 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 31970 14858 31984 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 31956 14858 31970 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 31942 14858 31956 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 31928 14858 31942 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 31914 14858 31928 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 31900 14858 31914 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 31886 14858 31900 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 31872 14858 31886 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 31858 14858 31872 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 31844 14858 31858 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 31830 14858 31844 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 31816 14858 31830 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 31802 14858 31816 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 31788 14858 31802 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 31774 14858 31788 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3361 32491 14858 34231 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 34931 14858 34940 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12213 34917 14858 34931 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12199 34903 14858 34917 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12185 34889 14858 34903 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12171 34875 14858 34889 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12157 34861 14858 34875 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12143 34847 14858 34861 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12129 34833 14858 34847 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12115 34819 14858 34833 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12101 34805 14858 34819 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12087 34791 14858 34805 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12073 34777 14858 34791 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12059 34763 14858 34777 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12045 34749 14858 34763 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12031 34735 14858 34749 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12017 34721 14858 34735 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12003 34707 14858 34721 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11989 34693 14858 34707 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11975 34679 14858 34693 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11961 34665 14858 34679 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11947 34651 14858 34665 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11933 34637 14858 34651 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11919 34623 14858 34637 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11905 34609 14858 34623 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11891 34595 14858 34609 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11877 34581 14858 34595 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11863 34567 14858 34581 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11849 34553 14858 34567 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11835 34539 14858 34553 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11821 34525 14858 34539 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11807 34511 14858 34525 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11793 34497 14858 34511 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11779 34483 14858 34497 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11765 34469 14858 34483 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11751 34455 14858 34469 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11737 34441 14858 34455 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11723 34427 14858 34441 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11709 34413 14858 34427 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11695 34399 14858 34413 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11681 34385 14858 34399 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11667 34371 14858 34385 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11653 34357 14858 34371 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11639 34343 14858 34357 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11625 34329 14858 34343 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11611 34315 14858 34329 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11597 34301 14858 34315 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11583 34287 14858 34301 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11569 34273 14858 34287 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11555 34259 14858 34273 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11541 34245 14858 34259 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11527 34231 14858 34245 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 34940 14858 36576 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11746 37052 14858 37059 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11760 37038 14858 37052 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11774 37024 14858 37038 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11788 37010 14858 37024 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11802 36996 14858 37010 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11816 36982 14858 36996 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11830 36968 14858 36982 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11844 36954 14858 36968 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11858 36940 14858 36954 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11872 36926 14858 36940 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11886 36912 14858 36926 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11900 36898 14858 36912 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11914 36884 14858 36898 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11928 36870 14858 36884 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11942 36856 14858 36870 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11956 36842 14858 36856 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11970 36828 14858 36842 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11984 36814 14858 36828 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11998 36800 14858 36814 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12012 36786 14858 36800 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12026 36772 14858 36786 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12040 36758 14858 36772 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12054 36744 14858 36758 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12068 36730 14858 36744 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12082 36716 14858 36730 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12096 36702 14858 36716 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12110 36688 14858 36702 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12124 36674 14858 36688 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12138 36660 14858 36674 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12152 36646 14858 36660 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12166 36632 14858 36646 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12180 36618 14858 36632 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12194 36604 14858 36618 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12208 36590 14858 36604 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 36576 14858 36590 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 3361 37059 14858 38003 6 drn_hvc
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
<< end >>
