magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< metal1 >>
rect -32 51671 -26 51723
rect 26 51671 32 51723
rect -32 637 -26 689
rect 26 637 32 689
rect 972 0 1008 52140
rect 1044 0 1080 52140
rect 1116 51429 1152 51770
rect 1116 50639 1152 51271
rect 1116 49849 1152 50481
rect 1116 49059 1152 49691
rect 1116 48269 1152 48901
rect 1116 47479 1152 48111
rect 1116 46689 1152 47321
rect 1116 45899 1152 46531
rect 1116 45109 1152 45741
rect 1116 44319 1152 44951
rect 1116 43529 1152 44161
rect 1116 42739 1152 43371
rect 1116 41949 1152 42581
rect 1116 41159 1152 41791
rect 1116 40369 1152 41001
rect 1116 39579 1152 40211
rect 1116 38789 1152 39421
rect 1116 37999 1152 38631
rect 1116 37209 1152 37841
rect 1116 36419 1152 37051
rect 1116 35629 1152 36261
rect 1116 34839 1152 35471
rect 1116 34049 1152 34681
rect 1116 33259 1152 33891
rect 1116 32469 1152 33101
rect 1116 31679 1152 32311
rect 1116 30889 1152 31521
rect 1116 30099 1152 30731
rect 1116 29309 1152 29941
rect 1116 28519 1152 29151
rect 1116 27729 1152 28361
rect 1116 26939 1152 27571
rect 1116 26149 1152 26781
rect 1116 25359 1152 25991
rect 1116 24569 1152 25201
rect 1116 23779 1152 24411
rect 1116 22989 1152 23621
rect 1116 22199 1152 22831
rect 1116 21409 1152 22041
rect 1116 20619 1152 21251
rect 1116 19829 1152 20461
rect 1116 19039 1152 19671
rect 1116 18249 1152 18881
rect 1116 17459 1152 18091
rect 1116 16669 1152 17301
rect 1116 15879 1152 16511
rect 1116 15089 1152 15721
rect 1116 14299 1152 14931
rect 1116 13509 1152 14141
rect 1116 12719 1152 13351
rect 1116 11929 1152 12561
rect 1116 11139 1152 11771
rect 1116 10349 1152 10981
rect 1116 9559 1152 10191
rect 1116 8769 1152 9401
rect 1116 7979 1152 8611
rect 1116 7189 1152 7821
rect 1116 6399 1152 7031
rect 1116 5609 1152 6241
rect 1116 4819 1152 5451
rect 1116 4029 1152 4661
rect 1116 3239 1152 3871
rect 1116 2449 1152 3081
rect 1116 1659 1152 2291
rect 1116 869 1152 1501
rect 1116 370 1152 711
rect 1188 0 1224 52140
rect 1260 0 1296 52140
rect 1452 0 1488 52140
rect 1524 0 1560 52140
rect 1668 0 1704 52140
rect 1740 0 1776 52140
rect 2220 0 2256 52140
rect 2292 0 2328 52140
rect 2436 0 2472 52140
rect 2508 0 2544 52140
rect 2700 0 2736 52140
rect 2772 0 2808 52140
rect 2916 0 2952 52140
rect 2988 0 3024 52140
rect 3468 0 3504 52140
rect 3540 0 3576 52140
rect 3684 0 3720 52140
rect 3756 0 3792 52140
rect 3948 0 3984 52140
rect 4020 0 4056 52140
rect 4164 0 4200 52140
rect 4236 0 4272 52140
rect 4716 0 4752 52140
rect 4788 0 4824 52140
rect 4932 0 4968 52140
rect 5004 0 5040 52140
rect 5196 0 5232 52140
rect 5268 0 5304 52140
rect 5412 0 5448 52140
rect 5484 0 5520 52140
rect 5964 0 6000 52140
rect 6036 0 6072 52140
rect 6180 0 6216 52140
rect 6252 0 6288 52140
rect 6444 0 6480 52140
rect 6516 0 6552 52140
rect 6660 0 6696 52140
rect 6732 0 6768 52140
rect 7212 0 7248 52140
rect 7284 0 7320 52140
rect 7428 0 7464 52140
rect 7500 0 7536 52140
rect 7692 0 7728 52140
rect 7764 0 7800 52140
rect 7908 0 7944 52140
rect 7980 0 8016 52140
rect 8460 0 8496 52140
rect 8532 0 8568 52140
rect 8676 0 8712 52140
rect 8748 0 8784 52140
rect 8940 0 8976 52140
rect 9012 0 9048 52140
rect 9156 0 9192 52140
rect 9228 0 9264 52140
rect 9708 0 9744 52140
rect 9780 0 9816 52140
rect 9924 0 9960 52140
rect 9996 0 10032 52140
rect 10188 0 10224 52140
rect 10260 0 10296 52140
rect 10404 0 10440 52140
rect 10476 0 10512 52140
rect 10956 0 10992 52140
rect 11028 0 11064 52140
rect 11172 0 11208 52140
rect 11244 0 11280 52140
rect 11436 0 11472 52140
rect 11508 0 11544 52140
rect 11652 0 11688 52140
rect 11724 0 11760 52140
rect 12204 0 12240 52140
rect 12276 0 12312 52140
rect 12420 0 12456 52140
rect 12492 0 12528 52140
rect 12684 0 12720 52140
rect 12756 0 12792 52140
rect 12900 0 12936 52140
rect 12972 0 13008 52140
rect 13452 0 13488 52140
rect 13524 0 13560 52140
rect 13668 0 13704 52140
rect 13740 0 13776 52140
rect 13932 0 13968 52140
rect 14004 0 14040 52140
rect 14148 0 14184 52140
rect 14220 0 14256 52140
rect 14700 0 14736 52140
rect 14772 0 14808 52140
rect 14916 0 14952 52140
rect 14988 0 15024 52140
rect 15180 0 15216 52140
rect 15252 0 15288 52140
rect 15396 0 15432 52140
rect 15468 0 15504 52140
rect 15948 0 15984 52140
rect 16020 0 16056 52140
rect 16164 0 16200 52140
rect 16236 0 16272 52140
rect 16428 0 16464 52140
rect 16500 0 16536 52140
rect 16644 0 16680 52140
rect 16716 0 16752 52140
rect 17196 0 17232 52140
rect 17268 0 17304 52140
rect 17412 0 17448 52140
rect 17484 0 17520 52140
rect 17676 0 17712 52140
rect 17748 0 17784 52140
rect 17892 0 17928 52140
rect 17964 0 18000 52140
rect 18444 0 18480 52140
rect 18516 0 18552 52140
rect 18660 0 18696 52140
rect 18732 0 18768 52140
rect 18924 0 18960 52140
rect 18996 0 19032 52140
rect 19140 0 19176 52140
rect 19212 0 19248 52140
rect 19692 0 19728 52140
rect 19764 0 19800 52140
rect 19908 0 19944 52140
rect 19980 0 20016 52140
rect 20172 0 20208 52140
rect 20244 0 20280 52140
rect 20388 0 20424 52140
rect 20460 0 20496 52140
rect 20940 0 20976 52140
rect 21012 0 21048 52140
rect 21156 0 21192 52140
rect 21228 0 21264 52140
rect 21420 0 21456 52140
rect 21492 0 21528 52140
rect 21636 0 21672 52140
rect 21708 0 21744 52140
rect 22188 0 22224 52140
rect 22260 0 22296 52140
rect 22404 0 22440 52140
rect 22476 0 22512 52140
rect 22668 0 22704 52140
rect 22740 0 22776 52140
rect 22884 0 22920 52140
rect 22956 0 22992 52140
rect 23436 0 23472 52140
rect 23508 0 23544 52140
rect 23652 0 23688 52140
rect 23724 0 23760 52140
rect 23916 0 23952 52140
rect 23988 0 24024 52140
rect 24132 0 24168 52140
rect 24204 0 24240 52140
rect 24684 0 24720 52140
rect 24756 0 24792 52140
rect 24900 0 24936 52140
rect 24972 0 25008 52140
rect 25164 0 25200 52140
rect 25236 0 25272 52140
rect 25380 0 25416 52140
rect 25452 0 25488 52140
rect 25932 0 25968 52140
rect 26004 0 26040 52140
rect 26148 0 26184 52140
rect 26220 0 26256 52140
rect 26412 0 26448 52140
rect 26484 0 26520 52140
rect 26628 0 26664 52140
rect 26700 0 26736 52140
rect 27180 0 27216 52140
rect 27252 0 27288 52140
rect 27396 0 27432 52140
rect 27468 0 27504 52140
rect 27660 0 27696 52140
rect 27732 0 27768 52140
rect 27876 0 27912 52140
rect 27948 0 27984 52140
rect 28428 0 28464 52140
rect 28500 0 28536 52140
rect 28644 0 28680 52140
rect 28716 0 28752 52140
rect 28908 0 28944 52140
rect 28980 0 29016 52140
rect 29124 0 29160 52140
rect 29196 0 29232 52140
rect 29676 0 29712 52140
rect 29748 0 29784 52140
rect 29892 0 29928 52140
rect 29964 0 30000 52140
rect 30156 0 30192 52140
rect 30228 0 30264 52140
rect 30372 0 30408 52140
rect 30444 0 30480 52140
rect 30924 0 30960 52140
rect 30996 0 31032 52140
rect 31140 0 31176 52140
rect 31212 0 31248 52140
rect 31404 0 31440 52140
rect 31476 0 31512 52140
rect 31620 0 31656 52140
rect 31692 0 31728 52140
rect 32172 0 32208 52140
rect 32244 0 32280 52140
rect 32388 0 32424 52140
rect 32460 0 32496 52140
rect 32652 0 32688 52140
rect 32724 0 32760 52140
rect 32868 0 32904 52140
rect 32940 0 32976 52140
rect 33420 0 33456 52140
rect 33492 0 33528 52140
rect 33636 0 33672 52140
rect 33708 0 33744 52140
rect 33900 0 33936 52140
rect 33972 0 34008 52140
rect 34116 0 34152 52140
rect 34188 0 34224 52140
rect 34668 0 34704 52140
rect 34740 0 34776 52140
rect 34884 0 34920 52140
rect 34956 0 34992 52140
rect 35148 0 35184 52140
rect 35220 0 35256 52140
rect 35364 0 35400 52140
rect 35436 0 35472 52140
rect 35916 0 35952 52140
rect 35988 0 36024 52140
rect 36132 0 36168 52140
rect 36204 0 36240 52140
rect 36396 0 36432 52140
rect 36468 0 36504 52140
rect 36612 0 36648 52140
rect 36684 0 36720 52140
rect 37164 0 37200 52140
rect 37236 0 37272 52140
rect 37380 0 37416 52140
rect 37452 0 37488 52140
rect 37644 0 37680 52140
rect 37716 0 37752 52140
rect 37860 0 37896 52140
rect 37932 0 37968 52140
rect 38412 0 38448 52140
rect 38484 0 38520 52140
rect 38628 0 38664 52140
rect 38700 0 38736 52140
rect 38892 0 38928 52140
rect 38964 0 39000 52140
rect 39108 0 39144 52140
rect 39180 0 39216 52140
rect 39660 0 39696 52140
rect 39732 0 39768 52140
rect 39876 0 39912 52140
rect 39948 0 39984 52140
rect 40140 0 40176 52140
rect 40212 0 40248 52140
rect 40356 0 40392 52140
rect 40428 0 40464 52140
rect 40908 0 40944 52140
rect 40980 0 41016 52140
rect 41124 0 41160 52140
rect 41196 0 41232 52140
rect 41388 0 41424 52140
rect 41460 0 41496 52140
rect 41532 51429 41568 51770
rect 41532 50639 41568 51271
rect 41532 49849 41568 50481
rect 41532 49059 41568 49691
rect 41532 48269 41568 48901
rect 41532 47479 41568 48111
rect 41532 46689 41568 47321
rect 41532 45899 41568 46531
rect 41532 45109 41568 45741
rect 41532 44319 41568 44951
rect 41532 43529 41568 44161
rect 41532 42739 41568 43371
rect 41532 41949 41568 42581
rect 41532 41159 41568 41791
rect 41532 40369 41568 41001
rect 41532 39579 41568 40211
rect 41532 38789 41568 39421
rect 41532 37999 41568 38631
rect 41532 37209 41568 37841
rect 41532 36419 41568 37051
rect 41532 35629 41568 36261
rect 41532 34839 41568 35471
rect 41532 34049 41568 34681
rect 41532 33259 41568 33891
rect 41532 32469 41568 33101
rect 41532 31679 41568 32311
rect 41532 30889 41568 31521
rect 41532 30099 41568 30731
rect 41532 29309 41568 29941
rect 41532 28519 41568 29151
rect 41532 27729 41568 28361
rect 41532 26939 41568 27571
rect 41532 26149 41568 26781
rect 41532 25359 41568 25991
rect 41532 24569 41568 25201
rect 41532 23779 41568 24411
rect 41532 22989 41568 23621
rect 41532 22199 41568 22831
rect 41532 21409 41568 22041
rect 41532 20619 41568 21251
rect 41532 19829 41568 20461
rect 41532 19039 41568 19671
rect 41532 18249 41568 18881
rect 41532 17459 41568 18091
rect 41532 16669 41568 17301
rect 41532 15879 41568 16511
rect 41532 15089 41568 15721
rect 41532 14299 41568 14931
rect 41532 13509 41568 14141
rect 41532 12719 41568 13351
rect 41532 11929 41568 12561
rect 41532 11139 41568 11771
rect 41532 10349 41568 10981
rect 41532 9559 41568 10191
rect 41532 8769 41568 9401
rect 41532 7979 41568 8611
rect 41532 7189 41568 7821
rect 41532 6399 41568 7031
rect 41532 5609 41568 6241
rect 41532 4819 41568 5451
rect 41532 4029 41568 4661
rect 41532 3239 41568 3871
rect 41532 2449 41568 3081
rect 41532 1659 41568 2291
rect 41532 869 41568 1501
rect 41532 370 41568 711
rect 41604 0 41640 52140
rect 41676 0 41712 52140
rect 42652 51671 42658 51723
rect 42710 51671 42716 51723
rect 42652 637 42658 689
rect 42710 637 42716 689
<< via1 >>
rect -26 51671 26 51723
rect -26 637 26 689
rect 42658 51671 42710 51723
rect 42658 637 42710 689
<< metal2 >>
rect -37 51669 -28 51725
rect 28 51721 37 51725
rect 42647 51721 42656 51725
rect 28 51673 42656 51721
rect 28 51669 37 51673
rect 42647 51669 42656 51673
rect 42712 51669 42721 51725
rect 1080 51549 1188 51625
rect 41496 51549 41604 51625
rect 0 51453 42684 51501
rect 1080 51295 1188 51405
rect 41496 51295 41604 51405
rect 0 51199 42684 51247
rect 1080 51075 1188 51151
rect 41496 51075 41604 51151
rect 0 50979 42684 51027
rect 0 50883 42684 50931
rect 1080 50759 1188 50835
rect 41496 50759 41604 50835
rect 0 50663 42684 50711
rect 1080 50505 1188 50615
rect 41496 50505 41604 50615
rect 0 50409 42684 50457
rect 1080 50285 1188 50361
rect 41496 50285 41604 50361
rect 0 50189 42684 50237
rect 0 50093 42684 50141
rect 1080 49969 1188 50045
rect 41496 49969 41604 50045
rect 0 49873 42684 49921
rect 1080 49715 1188 49825
rect 41496 49715 41604 49825
rect 0 49619 42684 49667
rect 1080 49495 1188 49571
rect 41496 49495 41604 49571
rect 0 49399 42684 49447
rect 0 49303 42684 49351
rect 1080 49179 1188 49255
rect 41496 49179 41604 49255
rect 0 49083 42684 49131
rect 1080 48925 1188 49035
rect 41496 48925 41604 49035
rect 0 48829 42684 48877
rect 1080 48705 1188 48781
rect 41496 48705 41604 48781
rect 0 48609 42684 48657
rect 0 48513 42684 48561
rect 1080 48389 1188 48465
rect 41496 48389 41604 48465
rect 0 48293 42684 48341
rect 1080 48135 1188 48245
rect 41496 48135 41604 48245
rect 0 48039 42684 48087
rect 1080 47915 1188 47991
rect 41496 47915 41604 47991
rect 0 47819 42684 47867
rect 0 47723 42684 47771
rect 1080 47599 1188 47675
rect 41496 47599 41604 47675
rect 0 47503 42684 47551
rect 1080 47345 1188 47455
rect 41496 47345 41604 47455
rect 0 47249 42684 47297
rect 1080 47125 1188 47201
rect 41496 47125 41604 47201
rect 0 47029 42684 47077
rect 0 46933 42684 46981
rect 1080 46809 1188 46885
rect 41496 46809 41604 46885
rect 0 46713 42684 46761
rect 1080 46555 1188 46665
rect 41496 46555 41604 46665
rect 0 46459 42684 46507
rect 1080 46335 1188 46411
rect 41496 46335 41604 46411
rect 0 46239 42684 46287
rect 0 46143 42684 46191
rect 1080 46019 1188 46095
rect 41496 46019 41604 46095
rect 0 45923 42684 45971
rect 1080 45765 1188 45875
rect 41496 45765 41604 45875
rect 0 45669 42684 45717
rect 1080 45545 1188 45621
rect 41496 45545 41604 45621
rect 0 45449 42684 45497
rect 0 45353 42684 45401
rect 1080 45229 1188 45305
rect 41496 45229 41604 45305
rect 0 45133 42684 45181
rect 1080 44975 1188 45085
rect 41496 44975 41604 45085
rect 0 44879 42684 44927
rect 1080 44755 1188 44831
rect 41496 44755 41604 44831
rect 0 44659 42684 44707
rect 0 44563 42684 44611
rect 1080 44439 1188 44515
rect 41496 44439 41604 44515
rect 0 44343 42684 44391
rect 1080 44185 1188 44295
rect 41496 44185 41604 44295
rect 0 44089 42684 44137
rect 1080 43965 1188 44041
rect 41496 43965 41604 44041
rect 0 43869 42684 43917
rect 0 43773 42684 43821
rect 1080 43649 1188 43725
rect 41496 43649 41604 43725
rect 0 43553 42684 43601
rect 1080 43395 1188 43505
rect 41496 43395 41604 43505
rect 0 43299 42684 43347
rect 1080 43175 1188 43251
rect 41496 43175 41604 43251
rect 0 43079 42684 43127
rect 0 42983 42684 43031
rect 1080 42859 1188 42935
rect 41496 42859 41604 42935
rect 0 42763 42684 42811
rect 1080 42605 1188 42715
rect 41496 42605 41604 42715
rect 0 42509 42684 42557
rect 1080 42385 1188 42461
rect 41496 42385 41604 42461
rect 0 42289 42684 42337
rect 0 42193 42684 42241
rect 1080 42069 1188 42145
rect 41496 42069 41604 42145
rect 0 41973 42684 42021
rect 1080 41815 1188 41925
rect 41496 41815 41604 41925
rect 0 41719 42684 41767
rect 1080 41595 1188 41671
rect 41496 41595 41604 41671
rect 0 41499 42684 41547
rect 0 41403 42684 41451
rect 1080 41279 1188 41355
rect 41496 41279 41604 41355
rect 0 41183 42684 41231
rect 1080 41025 1188 41135
rect 41496 41025 41604 41135
rect 0 40929 42684 40977
rect 1080 40805 1188 40881
rect 41496 40805 41604 40881
rect 0 40709 42684 40757
rect 0 40613 42684 40661
rect 1080 40489 1188 40565
rect 41496 40489 41604 40565
rect 0 40393 42684 40441
rect 1080 40235 1188 40345
rect 41496 40235 41604 40345
rect 0 40139 42684 40187
rect 1080 40015 1188 40091
rect 41496 40015 41604 40091
rect 0 39919 42684 39967
rect 0 39823 42684 39871
rect 1080 39699 1188 39775
rect 41496 39699 41604 39775
rect 0 39603 42684 39651
rect 1080 39445 1188 39555
rect 41496 39445 41604 39555
rect 0 39349 42684 39397
rect 1080 39225 1188 39301
rect 41496 39225 41604 39301
rect 0 39129 42684 39177
rect 0 39033 42684 39081
rect 1080 38909 1188 38985
rect 41496 38909 41604 38985
rect 0 38813 42684 38861
rect 1080 38655 1188 38765
rect 41496 38655 41604 38765
rect 0 38559 42684 38607
rect 1080 38435 1188 38511
rect 41496 38435 41604 38511
rect 0 38339 42684 38387
rect 0 38243 42684 38291
rect 1080 38119 1188 38195
rect 41496 38119 41604 38195
rect 0 38023 42684 38071
rect 1080 37865 1188 37975
rect 41496 37865 41604 37975
rect 0 37769 42684 37817
rect 1080 37645 1188 37721
rect 41496 37645 41604 37721
rect 0 37549 42684 37597
rect 0 37453 42684 37501
rect 1080 37329 1188 37405
rect 41496 37329 41604 37405
rect 0 37233 42684 37281
rect 1080 37075 1188 37185
rect 41496 37075 41604 37185
rect 0 36979 42684 37027
rect 1080 36855 1188 36931
rect 41496 36855 41604 36931
rect 0 36759 42684 36807
rect 0 36663 42684 36711
rect 1080 36539 1188 36615
rect 41496 36539 41604 36615
rect 0 36443 42684 36491
rect 1080 36285 1188 36395
rect 41496 36285 41604 36395
rect 0 36189 42684 36237
rect 1080 36065 1188 36141
rect 41496 36065 41604 36141
rect 0 35969 42684 36017
rect 0 35873 42684 35921
rect 1080 35749 1188 35825
rect 41496 35749 41604 35825
rect 0 35653 42684 35701
rect 1080 35495 1188 35605
rect 41496 35495 41604 35605
rect 0 35399 42684 35447
rect 1080 35275 1188 35351
rect 41496 35275 41604 35351
rect 0 35179 42684 35227
rect 0 35083 42684 35131
rect 1080 34959 1188 35035
rect 41496 34959 41604 35035
rect 0 34863 42684 34911
rect 1080 34705 1188 34815
rect 41496 34705 41604 34815
rect 0 34609 42684 34657
rect 1080 34485 1188 34561
rect 41496 34485 41604 34561
rect 0 34389 42684 34437
rect 0 34293 42684 34341
rect 1080 34169 1188 34245
rect 41496 34169 41604 34245
rect 0 34073 42684 34121
rect 1080 33915 1188 34025
rect 41496 33915 41604 34025
rect 0 33819 42684 33867
rect 1080 33695 1188 33771
rect 41496 33695 41604 33771
rect 0 33599 42684 33647
rect 0 33503 42684 33551
rect 1080 33379 1188 33455
rect 41496 33379 41604 33455
rect 0 33283 42684 33331
rect 1080 33125 1188 33235
rect 41496 33125 41604 33235
rect 0 33029 42684 33077
rect 1080 32905 1188 32981
rect 41496 32905 41604 32981
rect 0 32809 42684 32857
rect 0 32713 42684 32761
rect 1080 32589 1188 32665
rect 41496 32589 41604 32665
rect 0 32493 42684 32541
rect 1080 32335 1188 32445
rect 41496 32335 41604 32445
rect 0 32239 42684 32287
rect 1080 32115 1188 32191
rect 41496 32115 41604 32191
rect 0 32019 42684 32067
rect 0 31923 42684 31971
rect 1080 31799 1188 31875
rect 41496 31799 41604 31875
rect 0 31703 42684 31751
rect 1080 31545 1188 31655
rect 41496 31545 41604 31655
rect 0 31449 42684 31497
rect 1080 31325 1188 31401
rect 41496 31325 41604 31401
rect 0 31229 42684 31277
rect 0 31133 42684 31181
rect 1080 31009 1188 31085
rect 41496 31009 41604 31085
rect 0 30913 42684 30961
rect 1080 30755 1188 30865
rect 41496 30755 41604 30865
rect 0 30659 42684 30707
rect 1080 30535 1188 30611
rect 41496 30535 41604 30611
rect 0 30439 42684 30487
rect 0 30343 42684 30391
rect 1080 30219 1188 30295
rect 41496 30219 41604 30295
rect 0 30123 42684 30171
rect 1080 29965 1188 30075
rect 41496 29965 41604 30075
rect 0 29869 42684 29917
rect 1080 29745 1188 29821
rect 41496 29745 41604 29821
rect 0 29649 42684 29697
rect 0 29553 42684 29601
rect 1080 29429 1188 29505
rect 41496 29429 41604 29505
rect 0 29333 42684 29381
rect 1080 29175 1188 29285
rect 41496 29175 41604 29285
rect 0 29079 42684 29127
rect 1080 28955 1188 29031
rect 41496 28955 41604 29031
rect 0 28859 42684 28907
rect 0 28763 42684 28811
rect 1080 28639 1188 28715
rect 41496 28639 41604 28715
rect 0 28543 42684 28591
rect 1080 28385 1188 28495
rect 41496 28385 41604 28495
rect 0 28289 42684 28337
rect 1080 28165 1188 28241
rect 41496 28165 41604 28241
rect 0 28069 42684 28117
rect 0 27973 42684 28021
rect 1080 27849 1188 27925
rect 41496 27849 41604 27925
rect 0 27753 42684 27801
rect 1080 27595 1188 27705
rect 41496 27595 41604 27705
rect 0 27499 42684 27547
rect 1080 27375 1188 27451
rect 41496 27375 41604 27451
rect 0 27279 42684 27327
rect 0 27183 42684 27231
rect 1080 27059 1188 27135
rect 41496 27059 41604 27135
rect 0 26963 42684 27011
rect 1080 26805 1188 26915
rect 41496 26805 41604 26915
rect 0 26709 42684 26757
rect 1080 26585 1188 26661
rect 41496 26585 41604 26661
rect 0 26489 42684 26537
rect 0 26393 42684 26441
rect 1080 26269 1188 26345
rect 41496 26269 41604 26345
rect 0 26173 42684 26221
rect 1080 26015 1188 26125
rect 41496 26015 41604 26125
rect 0 25919 42684 25967
rect 1080 25795 1188 25871
rect 41496 25795 41604 25871
rect 0 25699 42684 25747
rect 0 25603 42684 25651
rect 1080 25479 1188 25555
rect 41496 25479 41604 25555
rect 0 25383 42684 25431
rect 1080 25225 1188 25335
rect 41496 25225 41604 25335
rect 0 25129 42684 25177
rect 1080 25005 1188 25081
rect 41496 25005 41604 25081
rect 0 24909 42684 24957
rect 0 24813 42684 24861
rect 1080 24689 1188 24765
rect 41496 24689 41604 24765
rect 0 24593 42684 24641
rect 1080 24435 1188 24545
rect 41496 24435 41604 24545
rect 0 24339 42684 24387
rect 1080 24215 1188 24291
rect 41496 24215 41604 24291
rect 0 24119 42684 24167
rect 0 24023 42684 24071
rect 1080 23899 1188 23975
rect 41496 23899 41604 23975
rect 0 23803 42684 23851
rect 1080 23645 1188 23755
rect 41496 23645 41604 23755
rect 0 23549 42684 23597
rect 1080 23425 1188 23501
rect 41496 23425 41604 23501
rect 0 23329 42684 23377
rect 0 23233 42684 23281
rect 1080 23109 1188 23185
rect 41496 23109 41604 23185
rect 0 23013 42684 23061
rect 1080 22855 1188 22965
rect 41496 22855 41604 22965
rect 0 22759 42684 22807
rect 1080 22635 1188 22711
rect 41496 22635 41604 22711
rect 0 22539 42684 22587
rect 0 22443 42684 22491
rect 1080 22319 1188 22395
rect 41496 22319 41604 22395
rect 0 22223 42684 22271
rect 1080 22065 1188 22175
rect 41496 22065 41604 22175
rect 0 21969 42684 22017
rect 1080 21845 1188 21921
rect 41496 21845 41604 21921
rect 0 21749 42684 21797
rect 0 21653 42684 21701
rect 1080 21529 1188 21605
rect 41496 21529 41604 21605
rect 0 21433 42684 21481
rect 1080 21275 1188 21385
rect 41496 21275 41604 21385
rect 0 21179 42684 21227
rect 1080 21055 1188 21131
rect 41496 21055 41604 21131
rect 0 20959 42684 21007
rect 0 20863 42684 20911
rect 1080 20739 1188 20815
rect 41496 20739 41604 20815
rect 0 20643 42684 20691
rect 1080 20485 1188 20595
rect 41496 20485 41604 20595
rect 0 20389 42684 20437
rect 1080 20265 1188 20341
rect 41496 20265 41604 20341
rect 0 20169 42684 20217
rect 0 20073 42684 20121
rect 1080 19949 1188 20025
rect 41496 19949 41604 20025
rect 0 19853 42684 19901
rect 1080 19695 1188 19805
rect 41496 19695 41604 19805
rect 0 19599 42684 19647
rect 1080 19475 1188 19551
rect 41496 19475 41604 19551
rect 0 19379 42684 19427
rect 0 19283 42684 19331
rect 1080 19159 1188 19235
rect 41496 19159 41604 19235
rect 0 19063 42684 19111
rect 1080 18905 1188 19015
rect 41496 18905 41604 19015
rect 0 18809 42684 18857
rect 1080 18685 1188 18761
rect 41496 18685 41604 18761
rect 0 18589 42684 18637
rect 0 18493 42684 18541
rect 1080 18369 1188 18445
rect 41496 18369 41604 18445
rect 0 18273 42684 18321
rect 1080 18115 1188 18225
rect 41496 18115 41604 18225
rect 0 18019 42684 18067
rect 1080 17895 1188 17971
rect 41496 17895 41604 17971
rect 0 17799 42684 17847
rect 0 17703 42684 17751
rect 1080 17579 1188 17655
rect 41496 17579 41604 17655
rect 0 17483 42684 17531
rect 1080 17325 1188 17435
rect 41496 17325 41604 17435
rect 0 17229 42684 17277
rect 1080 17105 1188 17181
rect 41496 17105 41604 17181
rect 0 17009 42684 17057
rect 0 16913 42684 16961
rect 1080 16789 1188 16865
rect 41496 16789 41604 16865
rect 0 16693 42684 16741
rect 1080 16535 1188 16645
rect 41496 16535 41604 16645
rect 0 16439 42684 16487
rect 1080 16315 1188 16391
rect 41496 16315 41604 16391
rect 0 16219 42684 16267
rect 0 16123 42684 16171
rect 1080 15999 1188 16075
rect 41496 15999 41604 16075
rect 0 15903 42684 15951
rect 1080 15745 1188 15855
rect 41496 15745 41604 15855
rect 0 15649 42684 15697
rect 1080 15525 1188 15601
rect 41496 15525 41604 15601
rect 0 15429 42684 15477
rect 0 15333 42684 15381
rect 1080 15209 1188 15285
rect 41496 15209 41604 15285
rect 0 15113 42684 15161
rect 1080 14955 1188 15065
rect 41496 14955 41604 15065
rect 0 14859 42684 14907
rect 1080 14735 1188 14811
rect 41496 14735 41604 14811
rect 0 14639 42684 14687
rect 0 14543 42684 14591
rect 1080 14419 1188 14495
rect 41496 14419 41604 14495
rect 0 14323 42684 14371
rect 1080 14165 1188 14275
rect 41496 14165 41604 14275
rect 0 14069 42684 14117
rect 1080 13945 1188 14021
rect 41496 13945 41604 14021
rect 0 13849 42684 13897
rect 0 13753 42684 13801
rect 1080 13629 1188 13705
rect 41496 13629 41604 13705
rect 0 13533 42684 13581
rect 1080 13375 1188 13485
rect 41496 13375 41604 13485
rect 0 13279 42684 13327
rect 1080 13155 1188 13231
rect 41496 13155 41604 13231
rect 0 13059 42684 13107
rect 0 12963 42684 13011
rect 1080 12839 1188 12915
rect 41496 12839 41604 12915
rect 0 12743 42684 12791
rect 1080 12585 1188 12695
rect 41496 12585 41604 12695
rect 0 12489 42684 12537
rect 1080 12365 1188 12441
rect 41496 12365 41604 12441
rect 0 12269 42684 12317
rect 0 12173 42684 12221
rect 1080 12049 1188 12125
rect 41496 12049 41604 12125
rect 0 11953 42684 12001
rect 1080 11795 1188 11905
rect 41496 11795 41604 11905
rect 0 11699 42684 11747
rect 1080 11575 1188 11651
rect 41496 11575 41604 11651
rect 0 11479 42684 11527
rect 0 11383 42684 11431
rect 1080 11259 1188 11335
rect 41496 11259 41604 11335
rect 0 11163 42684 11211
rect 1080 11005 1188 11115
rect 41496 11005 41604 11115
rect 0 10909 42684 10957
rect 1080 10785 1188 10861
rect 41496 10785 41604 10861
rect 0 10689 42684 10737
rect 0 10593 42684 10641
rect 1080 10469 1188 10545
rect 41496 10469 41604 10545
rect 0 10373 42684 10421
rect 1080 10215 1188 10325
rect 41496 10215 41604 10325
rect 0 10119 42684 10167
rect 1080 9995 1188 10071
rect 41496 9995 41604 10071
rect 0 9899 42684 9947
rect 0 9803 42684 9851
rect 1080 9679 1188 9755
rect 41496 9679 41604 9755
rect 0 9583 42684 9631
rect 1080 9425 1188 9535
rect 41496 9425 41604 9535
rect 0 9329 42684 9377
rect 1080 9205 1188 9281
rect 41496 9205 41604 9281
rect 0 9109 42684 9157
rect 0 9013 42684 9061
rect 1080 8889 1188 8965
rect 41496 8889 41604 8965
rect 0 8793 42684 8841
rect 1080 8635 1188 8745
rect 41496 8635 41604 8745
rect 0 8539 42684 8587
rect 1080 8415 1188 8491
rect 41496 8415 41604 8491
rect 0 8319 42684 8367
rect 0 8223 42684 8271
rect 1080 8099 1188 8175
rect 41496 8099 41604 8175
rect 0 8003 42684 8051
rect 1080 7845 1188 7955
rect 41496 7845 41604 7955
rect 0 7749 42684 7797
rect 1080 7625 1188 7701
rect 41496 7625 41604 7701
rect 0 7529 42684 7577
rect 0 7433 42684 7481
rect 1080 7309 1188 7385
rect 41496 7309 41604 7385
rect 0 7213 42684 7261
rect 1080 7055 1188 7165
rect 41496 7055 41604 7165
rect 0 6959 42684 7007
rect 1080 6835 1188 6911
rect 41496 6835 41604 6911
rect 0 6739 42684 6787
rect 0 6643 42684 6691
rect 1080 6519 1188 6595
rect 41496 6519 41604 6595
rect 0 6423 42684 6471
rect 1080 6265 1188 6375
rect 41496 6265 41604 6375
rect 0 6169 42684 6217
rect 1080 6045 1188 6121
rect 41496 6045 41604 6121
rect 0 5949 42684 5997
rect 0 5853 42684 5901
rect 1080 5729 1188 5805
rect 41496 5729 41604 5805
rect 0 5633 42684 5681
rect 1080 5475 1188 5585
rect 41496 5475 41604 5585
rect 0 5379 42684 5427
rect 1080 5255 1188 5331
rect 41496 5255 41604 5331
rect 0 5159 42684 5207
rect 0 5063 42684 5111
rect 1080 4939 1188 5015
rect 41496 4939 41604 5015
rect 0 4843 42684 4891
rect 1080 4685 1188 4795
rect 41496 4685 41604 4795
rect 0 4589 42684 4637
rect 1080 4465 1188 4541
rect 41496 4465 41604 4541
rect 0 4369 42684 4417
rect 0 4273 42684 4321
rect 1080 4149 1188 4225
rect 41496 4149 41604 4225
rect 0 4053 42684 4101
rect 1080 3895 1188 4005
rect 41496 3895 41604 4005
rect 0 3799 42684 3847
rect 1080 3675 1188 3751
rect 41496 3675 41604 3751
rect 0 3579 42684 3627
rect 0 3483 42684 3531
rect 1080 3359 1188 3435
rect 41496 3359 41604 3435
rect 0 3263 42684 3311
rect 1080 3105 1188 3215
rect 41496 3105 41604 3215
rect 0 3009 42684 3057
rect 1080 2885 1188 2961
rect 41496 2885 41604 2961
rect 0 2789 42684 2837
rect 0 2693 42684 2741
rect 1080 2569 1188 2645
rect 41496 2569 41604 2645
rect 0 2473 42684 2521
rect 1080 2315 1188 2425
rect 41496 2315 41604 2425
rect 0 2219 42684 2267
rect 1080 2095 1188 2171
rect 41496 2095 41604 2171
rect 0 1999 42684 2047
rect 0 1903 42684 1951
rect 1080 1779 1188 1855
rect 41496 1779 41604 1855
rect 0 1683 42684 1731
rect 1080 1525 1188 1635
rect 41496 1525 41604 1635
rect 0 1429 42684 1477
rect 1080 1305 1188 1381
rect 41496 1305 41604 1381
rect 0 1209 42684 1257
rect 0 1113 42684 1161
rect 1080 989 1188 1065
rect 41496 989 41604 1065
rect 0 893 42684 941
rect 1080 735 1188 845
rect 41496 735 41604 845
rect -37 635 -28 691
rect 28 687 37 691
rect 42647 687 42656 691
rect 28 639 42656 687
rect 28 635 37 639
rect 42647 635 42656 639
rect 42712 635 42721 691
rect 1080 515 1188 591
rect 41496 515 41604 591
rect 0 419 42684 467
<< via2 >>
rect -28 51723 28 51725
rect -28 51671 -26 51723
rect -26 51671 26 51723
rect 26 51671 28 51723
rect 42656 51723 42712 51725
rect -28 51669 28 51671
rect 42656 51671 42658 51723
rect 42658 51671 42710 51723
rect 42710 51671 42712 51723
rect 42656 51669 42712 51671
rect -28 689 28 691
rect -28 637 -26 689
rect -26 637 26 689
rect 26 637 28 689
rect 42656 689 42712 691
rect -28 635 28 637
rect 42656 637 42658 689
rect 42658 637 42710 689
rect 42710 637 42712 689
rect 42656 635 42712 637
<< metal3 >>
rect 1013 51862 1111 51960
rect 1637 51862 1735 51960
rect 2261 51862 2359 51960
rect 2885 51862 2983 51960
rect 3509 51862 3607 51960
rect 4133 51862 4231 51960
rect 4757 51862 4855 51960
rect 5381 51862 5479 51960
rect 6005 51862 6103 51960
rect 6629 51862 6727 51960
rect 7253 51862 7351 51960
rect 7877 51862 7975 51960
rect 8501 51862 8599 51960
rect 9125 51862 9223 51960
rect 9749 51862 9847 51960
rect 10373 51862 10471 51960
rect 10997 51862 11095 51960
rect 11621 51862 11719 51960
rect 12245 51862 12343 51960
rect 12869 51862 12967 51960
rect 13493 51862 13591 51960
rect 14117 51862 14215 51960
rect 14741 51862 14839 51960
rect 15365 51862 15463 51960
rect 15989 51862 16087 51960
rect 16613 51862 16711 51960
rect 17237 51862 17335 51960
rect 17861 51862 17959 51960
rect 18485 51862 18583 51960
rect 19109 51862 19207 51960
rect 19733 51862 19831 51960
rect 20357 51862 20455 51960
rect 20981 51862 21079 51960
rect 21605 51862 21703 51960
rect 22229 51862 22327 51960
rect 22853 51862 22951 51960
rect 23477 51862 23575 51960
rect 24101 51862 24199 51960
rect 24725 51862 24823 51960
rect 25349 51862 25447 51960
rect 25973 51862 26071 51960
rect 26597 51862 26695 51960
rect 27221 51862 27319 51960
rect 27845 51862 27943 51960
rect 28469 51862 28567 51960
rect 29093 51862 29191 51960
rect 29717 51862 29815 51960
rect 30341 51862 30439 51960
rect 30965 51862 31063 51960
rect 31589 51862 31687 51960
rect 32213 51862 32311 51960
rect 32837 51862 32935 51960
rect 33461 51862 33559 51960
rect 34085 51862 34183 51960
rect 34709 51862 34807 51960
rect 35333 51862 35431 51960
rect 35957 51862 36055 51960
rect 36581 51862 36679 51960
rect 37205 51862 37303 51960
rect 37829 51862 37927 51960
rect 38453 51862 38551 51960
rect 39077 51862 39175 51960
rect 39701 51862 39799 51960
rect 40325 51862 40423 51960
rect 40949 51862 41047 51960
rect 41573 51862 41671 51960
rect -49 51725 49 51746
rect -49 51669 -28 51725
rect 28 51669 49 51725
rect -49 51648 49 51669
rect 42635 51725 42733 51746
rect 42635 51669 42656 51725
rect 42712 51669 42733 51725
rect 42635 51648 42733 51669
rect 317 51301 415 51399
rect 42269 51301 42367 51399
rect 317 51064 415 51162
rect 42269 51064 42367 51162
rect 317 50748 415 50846
rect 42269 50748 42367 50846
rect 317 50511 415 50609
rect 42269 50511 42367 50609
rect 317 50274 415 50372
rect 42269 50274 42367 50372
rect 317 49958 415 50056
rect 42269 49958 42367 50056
rect 317 49721 415 49819
rect 42269 49721 42367 49819
rect 317 49484 415 49582
rect 42269 49484 42367 49582
rect 317 49168 415 49266
rect 42269 49168 42367 49266
rect 317 48931 415 49029
rect 42269 48931 42367 49029
rect 317 48694 415 48792
rect 42269 48694 42367 48792
rect 317 48378 415 48476
rect 42269 48378 42367 48476
rect 317 48141 415 48239
rect 42269 48141 42367 48239
rect 317 47904 415 48002
rect 42269 47904 42367 48002
rect 317 47588 415 47686
rect 42269 47588 42367 47686
rect 317 47351 415 47449
rect 42269 47351 42367 47449
rect 317 47114 415 47212
rect 42269 47114 42367 47212
rect 317 46798 415 46896
rect 42269 46798 42367 46896
rect 317 46561 415 46659
rect 42269 46561 42367 46659
rect 317 46324 415 46422
rect 42269 46324 42367 46422
rect 317 46008 415 46106
rect 42269 46008 42367 46106
rect 317 45771 415 45869
rect 42269 45771 42367 45869
rect 317 45534 415 45632
rect 42269 45534 42367 45632
rect 317 45218 415 45316
rect 42269 45218 42367 45316
rect 317 44981 415 45079
rect 42269 44981 42367 45079
rect 317 44744 415 44842
rect 42269 44744 42367 44842
rect 317 44428 415 44526
rect 42269 44428 42367 44526
rect 317 44191 415 44289
rect 42269 44191 42367 44289
rect 317 43954 415 44052
rect 42269 43954 42367 44052
rect 317 43638 415 43736
rect 42269 43638 42367 43736
rect 317 43401 415 43499
rect 42269 43401 42367 43499
rect 317 43164 415 43262
rect 42269 43164 42367 43262
rect 317 42848 415 42946
rect 42269 42848 42367 42946
rect 317 42611 415 42709
rect 42269 42611 42367 42709
rect 317 42374 415 42472
rect 42269 42374 42367 42472
rect 317 42058 415 42156
rect 42269 42058 42367 42156
rect 317 41821 415 41919
rect 42269 41821 42367 41919
rect 317 41584 415 41682
rect 42269 41584 42367 41682
rect 317 41268 415 41366
rect 42269 41268 42367 41366
rect 317 41031 415 41129
rect 42269 41031 42367 41129
rect 317 40794 415 40892
rect 42269 40794 42367 40892
rect 317 40478 415 40576
rect 42269 40478 42367 40576
rect 317 40241 415 40339
rect 42269 40241 42367 40339
rect 317 40004 415 40102
rect 42269 40004 42367 40102
rect 317 39688 415 39786
rect 42269 39688 42367 39786
rect 317 39451 415 39549
rect 42269 39451 42367 39549
rect 317 39214 415 39312
rect 42269 39214 42367 39312
rect 317 38898 415 38996
rect 42269 38898 42367 38996
rect 317 38661 415 38759
rect 42269 38661 42367 38759
rect 317 38424 415 38522
rect 42269 38424 42367 38522
rect 317 38108 415 38206
rect 42269 38108 42367 38206
rect 317 37871 415 37969
rect 42269 37871 42367 37969
rect 317 37634 415 37732
rect 42269 37634 42367 37732
rect 317 37318 415 37416
rect 42269 37318 42367 37416
rect 317 37081 415 37179
rect 42269 37081 42367 37179
rect 317 36844 415 36942
rect 42269 36844 42367 36942
rect 317 36528 415 36626
rect 42269 36528 42367 36626
rect 317 36291 415 36389
rect 42269 36291 42367 36389
rect 317 36054 415 36152
rect 42269 36054 42367 36152
rect 317 35738 415 35836
rect 42269 35738 42367 35836
rect 317 35501 415 35599
rect 42269 35501 42367 35599
rect 317 35264 415 35362
rect 42269 35264 42367 35362
rect 317 34948 415 35046
rect 42269 34948 42367 35046
rect 317 34711 415 34809
rect 42269 34711 42367 34809
rect 317 34474 415 34572
rect 42269 34474 42367 34572
rect 317 34158 415 34256
rect 42269 34158 42367 34256
rect 317 33921 415 34019
rect 42269 33921 42367 34019
rect 317 33684 415 33782
rect 42269 33684 42367 33782
rect 317 33368 415 33466
rect 42269 33368 42367 33466
rect 317 33131 415 33229
rect 42269 33131 42367 33229
rect 317 32894 415 32992
rect 42269 32894 42367 32992
rect 317 32578 415 32676
rect 42269 32578 42367 32676
rect 317 32341 415 32439
rect 42269 32341 42367 32439
rect 317 32104 415 32202
rect 42269 32104 42367 32202
rect 317 31788 415 31886
rect 42269 31788 42367 31886
rect 317 31551 415 31649
rect 42269 31551 42367 31649
rect 317 31314 415 31412
rect 42269 31314 42367 31412
rect 317 30998 415 31096
rect 42269 30998 42367 31096
rect 317 30761 415 30859
rect 42269 30761 42367 30859
rect 317 30524 415 30622
rect 42269 30524 42367 30622
rect 317 30208 415 30306
rect 42269 30208 42367 30306
rect 317 29971 415 30069
rect 42269 29971 42367 30069
rect 317 29734 415 29832
rect 42269 29734 42367 29832
rect 317 29418 415 29516
rect 42269 29418 42367 29516
rect 317 29181 415 29279
rect 42269 29181 42367 29279
rect 317 28944 415 29042
rect 42269 28944 42367 29042
rect 317 28628 415 28726
rect 42269 28628 42367 28726
rect 317 28391 415 28489
rect 42269 28391 42367 28489
rect 317 28154 415 28252
rect 42269 28154 42367 28252
rect 317 27838 415 27936
rect 42269 27838 42367 27936
rect 317 27601 415 27699
rect 42269 27601 42367 27699
rect 317 27364 415 27462
rect 42269 27364 42367 27462
rect 317 27048 415 27146
rect 42269 27048 42367 27146
rect 317 26811 415 26909
rect 42269 26811 42367 26909
rect 317 26574 415 26672
rect 42269 26574 42367 26672
rect 317 26258 415 26356
rect 42269 26258 42367 26356
rect 317 26021 415 26119
rect 42269 26021 42367 26119
rect 317 25784 415 25882
rect 42269 25784 42367 25882
rect 317 25468 415 25566
rect 42269 25468 42367 25566
rect 317 25231 415 25329
rect 42269 25231 42367 25329
rect 317 24994 415 25092
rect 42269 24994 42367 25092
rect 317 24678 415 24776
rect 42269 24678 42367 24776
rect 317 24441 415 24539
rect 42269 24441 42367 24539
rect 317 24204 415 24302
rect 42269 24204 42367 24302
rect 317 23888 415 23986
rect 42269 23888 42367 23986
rect 317 23651 415 23749
rect 42269 23651 42367 23749
rect 317 23414 415 23512
rect 42269 23414 42367 23512
rect 317 23098 415 23196
rect 42269 23098 42367 23196
rect 317 22861 415 22959
rect 42269 22861 42367 22959
rect 317 22624 415 22722
rect 42269 22624 42367 22722
rect 317 22308 415 22406
rect 42269 22308 42367 22406
rect 317 22071 415 22169
rect 42269 22071 42367 22169
rect 317 21834 415 21932
rect 42269 21834 42367 21932
rect 317 21518 415 21616
rect 42269 21518 42367 21616
rect 317 21281 415 21379
rect 42269 21281 42367 21379
rect 317 21044 415 21142
rect 42269 21044 42367 21142
rect 317 20728 415 20826
rect 42269 20728 42367 20826
rect 317 20491 415 20589
rect 42269 20491 42367 20589
rect 317 20254 415 20352
rect 42269 20254 42367 20352
rect 317 19938 415 20036
rect 42269 19938 42367 20036
rect 317 19701 415 19799
rect 42269 19701 42367 19799
rect 317 19464 415 19562
rect 42269 19464 42367 19562
rect 317 19148 415 19246
rect 42269 19148 42367 19246
rect 317 18911 415 19009
rect 42269 18911 42367 19009
rect 317 18674 415 18772
rect 42269 18674 42367 18772
rect 317 18358 415 18456
rect 42269 18358 42367 18456
rect 317 18121 415 18219
rect 42269 18121 42367 18219
rect 317 17884 415 17982
rect 42269 17884 42367 17982
rect 317 17568 415 17666
rect 42269 17568 42367 17666
rect 317 17331 415 17429
rect 42269 17331 42367 17429
rect 317 17094 415 17192
rect 42269 17094 42367 17192
rect 317 16778 415 16876
rect 42269 16778 42367 16876
rect 317 16541 415 16639
rect 42269 16541 42367 16639
rect 317 16304 415 16402
rect 42269 16304 42367 16402
rect 317 15988 415 16086
rect 42269 15988 42367 16086
rect 317 15751 415 15849
rect 42269 15751 42367 15849
rect 317 15514 415 15612
rect 42269 15514 42367 15612
rect 317 15198 415 15296
rect 42269 15198 42367 15296
rect 317 14961 415 15059
rect 42269 14961 42367 15059
rect 317 14724 415 14822
rect 42269 14724 42367 14822
rect 317 14408 415 14506
rect 42269 14408 42367 14506
rect 317 14171 415 14269
rect 42269 14171 42367 14269
rect 317 13934 415 14032
rect 42269 13934 42367 14032
rect 317 13618 415 13716
rect 42269 13618 42367 13716
rect 317 13381 415 13479
rect 42269 13381 42367 13479
rect 317 13144 415 13242
rect 42269 13144 42367 13242
rect 317 12828 415 12926
rect 42269 12828 42367 12926
rect 317 12591 415 12689
rect 42269 12591 42367 12689
rect 317 12354 415 12452
rect 42269 12354 42367 12452
rect 317 12038 415 12136
rect 42269 12038 42367 12136
rect 317 11801 415 11899
rect 42269 11801 42367 11899
rect 317 11564 415 11662
rect 42269 11564 42367 11662
rect 317 11248 415 11346
rect 42269 11248 42367 11346
rect 317 11011 415 11109
rect 42269 11011 42367 11109
rect 317 10774 415 10872
rect 42269 10774 42367 10872
rect 317 10458 415 10556
rect 42269 10458 42367 10556
rect 317 10221 415 10319
rect 42269 10221 42367 10319
rect 317 9984 415 10082
rect 42269 9984 42367 10082
rect 317 9668 415 9766
rect 42269 9668 42367 9766
rect 317 9431 415 9529
rect 42269 9431 42367 9529
rect 317 9194 415 9292
rect 42269 9194 42367 9292
rect 317 8878 415 8976
rect 42269 8878 42367 8976
rect 317 8641 415 8739
rect 42269 8641 42367 8739
rect 317 8404 415 8502
rect 42269 8404 42367 8502
rect 317 8088 415 8186
rect 42269 8088 42367 8186
rect 317 7851 415 7949
rect 42269 7851 42367 7949
rect 317 7614 415 7712
rect 42269 7614 42367 7712
rect 317 7298 415 7396
rect 42269 7298 42367 7396
rect 317 7061 415 7159
rect 42269 7061 42367 7159
rect 317 6824 415 6922
rect 42269 6824 42367 6922
rect 317 6508 415 6606
rect 42269 6508 42367 6606
rect 317 6271 415 6369
rect 42269 6271 42367 6369
rect 317 6034 415 6132
rect 42269 6034 42367 6132
rect 317 5718 415 5816
rect 42269 5718 42367 5816
rect 317 5481 415 5579
rect 42269 5481 42367 5579
rect 317 5244 415 5342
rect 42269 5244 42367 5342
rect 317 4928 415 5026
rect 42269 4928 42367 5026
rect 317 4691 415 4789
rect 42269 4691 42367 4789
rect 317 4454 415 4552
rect 42269 4454 42367 4552
rect 317 4138 415 4236
rect 42269 4138 42367 4236
rect 317 3901 415 3999
rect 42269 3901 42367 3999
rect 317 3664 415 3762
rect 42269 3664 42367 3762
rect 317 3348 415 3446
rect 42269 3348 42367 3446
rect 317 3111 415 3209
rect 42269 3111 42367 3209
rect 317 2874 415 2972
rect 42269 2874 42367 2972
rect 317 2558 415 2656
rect 42269 2558 42367 2656
rect 317 2321 415 2419
rect 42269 2321 42367 2419
rect 317 2084 415 2182
rect 42269 2084 42367 2182
rect 317 1768 415 1866
rect 42269 1768 42367 1866
rect 317 1531 415 1629
rect 42269 1531 42367 1629
rect 317 1294 415 1392
rect 42269 1294 42367 1392
rect 317 978 415 1076
rect 42269 978 42367 1076
rect 317 741 415 839
rect 42269 741 42367 839
rect -49 691 49 712
rect -49 635 -28 691
rect 28 635 49 691
rect -49 614 49 635
rect 42635 691 42733 712
rect 42635 635 42656 691
rect 42712 635 42733 691
rect 42635 614 42733 635
rect 1013 180 1111 278
rect 1637 180 1735 278
rect 2261 180 2359 278
rect 2885 180 2983 278
rect 3509 180 3607 278
rect 4133 180 4231 278
rect 4757 180 4855 278
rect 5381 180 5479 278
rect 6005 180 6103 278
rect 6629 180 6727 278
rect 7253 180 7351 278
rect 7877 180 7975 278
rect 8501 180 8599 278
rect 9125 180 9223 278
rect 9749 180 9847 278
rect 10373 180 10471 278
rect 10997 180 11095 278
rect 11621 180 11719 278
rect 12245 180 12343 278
rect 12869 180 12967 278
rect 13493 180 13591 278
rect 14117 180 14215 278
rect 14741 180 14839 278
rect 15365 180 15463 278
rect 15989 180 16087 278
rect 16613 180 16711 278
rect 17237 180 17335 278
rect 17861 180 17959 278
rect 18485 180 18583 278
rect 19109 180 19207 278
rect 19733 180 19831 278
rect 20357 180 20455 278
rect 20981 180 21079 278
rect 21605 180 21703 278
rect 22229 180 22327 278
rect 22853 180 22951 278
rect 23477 180 23575 278
rect 24101 180 24199 278
rect 24725 180 24823 278
rect 25349 180 25447 278
rect 25973 180 26071 278
rect 26597 180 26695 278
rect 27221 180 27319 278
rect 27845 180 27943 278
rect 28469 180 28567 278
rect 29093 180 29191 278
rect 29717 180 29815 278
rect 30341 180 30439 278
rect 30965 180 31063 278
rect 31589 180 31687 278
rect 32213 180 32311 278
rect 32837 180 32935 278
rect 33461 180 33559 278
rect 34085 180 34183 278
rect 34709 180 34807 278
rect 35333 180 35431 278
rect 35957 180 36055 278
rect 36581 180 36679 278
rect 37205 180 37303 278
rect 37829 180 37927 278
rect 38453 180 38551 278
rect 39077 180 39175 278
rect 39701 180 39799 278
rect 40325 180 40423 278
rect 40949 180 41047 278
rect 41573 180 41671 278
use sky130_sram_1kbyte_1rw1r_8x1024_8_bitcell_array  sky130_sram_1kbyte_1rw1r_8x1024_8_bitcell_array_0
timestamp 1704896540
transform 1 0 1374 0 1 790
box -42 -105 39978 50665
use sky130_sram_1kbyte_1rw1r_8x1024_8_col_cap_array  sky130_sram_1kbyte_1rw1r_8x1024_8_col_cap_array_0
timestamp 1704896540
transform 1 0 1374 0 -1 52140
box 0 0 39936 474
use sky130_sram_1kbyte_1rw1r_8x1024_8_col_cap_array_0  sky130_sram_1kbyte_1rw1r_8x1024_8_col_cap_array_0_0
timestamp 1704896540
transform 1 0 1374 0 1 0
box 0 0 39936 474
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8_0
timestamp 1704896540
transform 1 0 42652 0 1 51671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8_1
timestamp 1704896540
transform 1 0 -32 0 1 51671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8_2
timestamp 1704896540
transform 1 0 42652 0 1 637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_8_3
timestamp 1704896540
transform 1 0 -32 0 1 637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9_0
timestamp 1704896540
transform 1 0 42647 0 1 51664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9_1
timestamp 1704896540
transform 1 0 -37 0 1 51664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9_2
timestamp 1704896540
transform 1 0 42647 0 1 630
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_9_3
timestamp 1704896540
transform 1 0 -37 0 1 630
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_dummy_array  sky130_sram_1kbyte_1rw1r_8x1024_8_dummy_array_0
timestamp 1704896540
transform 1 0 1374 0 1 51350
box -42 -105 39978 421
use sky130_sram_1kbyte_1rw1r_8x1024_8_dummy_array  sky130_sram_1kbyte_1rw1r_8x1024_8_dummy_array_1
timestamp 1704896540
transform 1 0 1374 0 -1 790
box -42 -105 39978 421
use sky130_sram_1kbyte_1rw1r_8x1024_8_replica_column  sky130_sram_1kbyte_1rw1r_8x1024_8_replica_column_0
timestamp 1704896540
transform 1 0 750 0 1 0
box -26 0 666 52140
use sky130_sram_1kbyte_1rw1r_8x1024_8_replica_column_0  sky130_sram_1kbyte_1rw1r_8x1024_8_replica_column_0_0
timestamp 1704896540
transform 1 0 41310 0 1 0
box -42 0 650 52140
use sky130_sram_1kbyte_1rw1r_8x1024_8_row_cap_array  sky130_sram_1kbyte_1rw1r_8x1024_8_row_cap_array_0
timestamp 1704896540
transform 1 0 126 0 1 0
box -42 419 624 51721
use sky130_sram_1kbyte_1rw1r_8x1024_8_row_cap_array_0  sky130_sram_1kbyte_1rw1r_8x1024_8_row_cap_array_0_0
timestamp 1704896540
transform 1 0 41934 0 1 0
box 0 419 666 51721
<< labels >>
rlabel metal3 s 40949 51862 41047 51960 4 vdd
port 1 nsew
rlabel metal3 s 38453 51862 38551 51960 4 vdd
port 1 nsew
rlabel metal3 s 32837 51862 32935 51960 4 vdd
port 1 nsew
rlabel metal3 s 39701 51862 39799 51960 4 vdd
port 1 nsew
rlabel metal3 s 34085 51862 34183 51960 4 vdd
port 1 nsew
rlabel metal3 s 35333 51862 35431 51960 4 vdd
port 1 nsew
rlabel metal3 s 32213 51862 32311 51960 4 vdd
port 1 nsew
rlabel metal3 s 37829 51862 37927 51960 4 vdd
port 1 nsew
rlabel metal3 s 37205 51862 37303 51960 4 vdd
port 1 nsew
rlabel metal3 s 35957 51862 36055 51960 4 vdd
port 1 nsew
rlabel metal3 s 39077 51862 39175 51960 4 vdd
port 1 nsew
rlabel metal3 s 36581 51862 36679 51960 4 vdd
port 1 nsew
rlabel metal3 s 41573 51862 41671 51960 4 vdd
port 1 nsew
rlabel metal3 s 40325 51862 40423 51960 4 vdd
port 1 nsew
rlabel metal3 s 33461 51862 33559 51960 4 vdd
port 1 nsew
rlabel metal3 s 34709 51862 34807 51960 4 vdd
port 1 nsew
rlabel metal3 s 42269 46561 42367 46659 4 gnd
port 2 nsew
rlabel metal3 s 42269 50748 42367 50846 4 gnd
port 2 nsew
rlabel metal3 s 42269 44191 42367 44289 4 gnd
port 2 nsew
rlabel metal3 s 42269 40004 42367 40102 4 gnd
port 2 nsew
rlabel metal3 s 42635 51648 42733 51746 4 gnd
port 2 nsew
rlabel metal3 s 42269 47904 42367 48002 4 gnd
port 2 nsew
rlabel metal3 s 42269 47351 42367 47449 4 gnd
port 2 nsew
rlabel metal3 s 42269 40478 42367 40576 4 gnd
port 2 nsew
rlabel metal3 s 42269 48378 42367 48476 4 gnd
port 2 nsew
rlabel metal3 s 42269 43401 42367 43499 4 gnd
port 2 nsew
rlabel metal3 s 42269 49484 42367 49582 4 gnd
port 2 nsew
rlabel metal3 s 42269 41268 42367 41366 4 gnd
port 2 nsew
rlabel metal3 s 42269 48931 42367 49029 4 gnd
port 2 nsew
rlabel metal3 s 42269 49721 42367 49819 4 gnd
port 2 nsew
rlabel metal3 s 42269 43164 42367 43262 4 gnd
port 2 nsew
rlabel metal3 s 42269 44428 42367 44526 4 gnd
port 2 nsew
rlabel metal3 s 42269 46008 42367 46106 4 gnd
port 2 nsew
rlabel metal3 s 42269 50511 42367 50609 4 gnd
port 2 nsew
rlabel metal3 s 42269 48694 42367 48792 4 gnd
port 2 nsew
rlabel metal3 s 42269 44981 42367 45079 4 gnd
port 2 nsew
rlabel metal3 s 42269 49958 42367 50056 4 gnd
port 2 nsew
rlabel metal3 s 42269 47588 42367 47686 4 gnd
port 2 nsew
rlabel metal3 s 42269 43954 42367 44052 4 gnd
port 2 nsew
rlabel metal3 s 42269 42058 42367 42156 4 gnd
port 2 nsew
rlabel metal3 s 42269 41821 42367 41919 4 gnd
port 2 nsew
rlabel metal3 s 42269 41584 42367 41682 4 gnd
port 2 nsew
rlabel metal3 s 42269 40241 42367 40339 4 gnd
port 2 nsew
rlabel metal3 s 42269 41031 42367 41129 4 gnd
port 2 nsew
rlabel metal3 s 42269 48141 42367 48239 4 gnd
port 2 nsew
rlabel metal3 s 42269 43638 42367 43736 4 gnd
port 2 nsew
rlabel metal3 s 42269 42848 42367 42946 4 gnd
port 2 nsew
rlabel metal3 s 42269 49168 42367 49266 4 gnd
port 2 nsew
rlabel metal3 s 42269 51301 42367 51399 4 gnd
port 2 nsew
rlabel metal3 s 42269 45534 42367 45632 4 gnd
port 2 nsew
rlabel metal3 s 42269 39451 42367 39549 4 gnd
port 2 nsew
rlabel metal3 s 42269 50274 42367 50372 4 gnd
port 2 nsew
rlabel metal3 s 42269 45771 42367 45869 4 gnd
port 2 nsew
rlabel metal3 s 42269 47114 42367 47212 4 gnd
port 2 nsew
rlabel metal3 s 42269 42374 42367 42472 4 gnd
port 2 nsew
rlabel metal3 s 42269 45218 42367 45316 4 gnd
port 2 nsew
rlabel metal3 s 42269 46798 42367 46896 4 gnd
port 2 nsew
rlabel metal3 s 42269 44744 42367 44842 4 gnd
port 2 nsew
rlabel metal3 s 42269 40794 42367 40892 4 gnd
port 2 nsew
rlabel metal3 s 42269 39688 42367 39786 4 gnd
port 2 nsew
rlabel metal3 s 42269 46324 42367 46422 4 gnd
port 2 nsew
rlabel metal3 s 42269 42611 42367 42709 4 gnd
port 2 nsew
rlabel metal3 s 42269 51064 42367 51162 4 gnd
port 2 nsew
rlabel metal3 s 42269 39214 42367 39312 4 gnd
port 2 nsew
rlabel metal3 s 25973 51862 26071 51960 4 vdd
port 1 nsew
rlabel metal3 s 24725 51862 24823 51960 4 vdd
port 1 nsew
rlabel metal3 s 30965 51862 31063 51960 4 vdd
port 1 nsew
rlabel metal3 s 21605 51862 21703 51960 4 vdd
port 1 nsew
rlabel metal3 s 25349 51862 25447 51960 4 vdd
port 1 nsew
rlabel metal3 s 29093 51862 29191 51960 4 vdd
port 1 nsew
rlabel metal3 s 29717 51862 29815 51960 4 vdd
port 1 nsew
rlabel metal3 s 27221 51862 27319 51960 4 vdd
port 1 nsew
rlabel metal3 s 24101 51862 24199 51960 4 vdd
port 1 nsew
rlabel metal3 s 26597 51862 26695 51960 4 vdd
port 1 nsew
rlabel metal3 s 31589 51862 31687 51960 4 vdd
port 1 nsew
rlabel metal3 s 22853 51862 22951 51960 4 vdd
port 1 nsew
rlabel metal3 s 23477 51862 23575 51960 4 vdd
port 1 nsew
rlabel metal3 s 28469 51862 28567 51960 4 vdd
port 1 nsew
rlabel metal3 s 30341 51862 30439 51960 4 vdd
port 1 nsew
rlabel metal3 s 22229 51862 22327 51960 4 vdd
port 1 nsew
rlabel metal3 s 27845 51862 27943 51960 4 vdd
port 1 nsew
rlabel metal3 s 42269 27048 42367 27146 4 gnd
port 2 nsew
rlabel metal3 s 42269 36528 42367 36626 4 gnd
port 2 nsew
rlabel metal3 s 42269 30761 42367 30859 4 gnd
port 2 nsew
rlabel metal3 s 42269 32578 42367 32676 4 gnd
port 2 nsew
rlabel metal3 s 42269 31788 42367 31886 4 gnd
port 2 nsew
rlabel metal3 s 42269 34948 42367 35046 4 gnd
port 2 nsew
rlabel metal3 s 42269 37081 42367 37179 4 gnd
port 2 nsew
rlabel metal3 s 42269 37318 42367 37416 4 gnd
port 2 nsew
rlabel metal3 s 42269 30524 42367 30622 4 gnd
port 2 nsew
rlabel metal3 s 42269 29734 42367 29832 4 gnd
port 2 nsew
rlabel metal3 s 42269 38661 42367 38759 4 gnd
port 2 nsew
rlabel metal3 s 42269 34158 42367 34256 4 gnd
port 2 nsew
rlabel metal3 s 42269 36291 42367 36389 4 gnd
port 2 nsew
rlabel metal3 s 42269 31551 42367 31649 4 gnd
port 2 nsew
rlabel metal3 s 42269 30208 42367 30306 4 gnd
port 2 nsew
rlabel metal3 s 42269 34474 42367 34572 4 gnd
port 2 nsew
rlabel metal3 s 42269 36054 42367 36152 4 gnd
port 2 nsew
rlabel metal3 s 42269 38424 42367 38522 4 gnd
port 2 nsew
rlabel metal3 s 42269 37871 42367 37969 4 gnd
port 2 nsew
rlabel metal3 s 42269 28628 42367 28726 4 gnd
port 2 nsew
rlabel metal3 s 42269 32341 42367 32439 4 gnd
port 2 nsew
rlabel metal3 s 42269 35738 42367 35836 4 gnd
port 2 nsew
rlabel metal3 s 42269 33684 42367 33782 4 gnd
port 2 nsew
rlabel metal3 s 42269 36844 42367 36942 4 gnd
port 2 nsew
rlabel metal3 s 42269 30998 42367 31096 4 gnd
port 2 nsew
rlabel metal3 s 42269 32104 42367 32202 4 gnd
port 2 nsew
rlabel metal3 s 42269 29971 42367 30069 4 gnd
port 2 nsew
rlabel metal3 s 42269 28391 42367 28489 4 gnd
port 2 nsew
rlabel metal3 s 42269 38108 42367 38206 4 gnd
port 2 nsew
rlabel metal3 s 42269 26574 42367 26672 4 gnd
port 2 nsew
rlabel metal3 s 42269 35501 42367 35599 4 gnd
port 2 nsew
rlabel metal3 s 42269 33131 42367 33229 4 gnd
port 2 nsew
rlabel metal3 s 42269 35264 42367 35362 4 gnd
port 2 nsew
rlabel metal3 s 42269 33368 42367 33466 4 gnd
port 2 nsew
rlabel metal3 s 42269 28944 42367 29042 4 gnd
port 2 nsew
rlabel metal3 s 42269 27601 42367 27699 4 gnd
port 2 nsew
rlabel metal3 s 42269 32894 42367 32992 4 gnd
port 2 nsew
rlabel metal3 s 42269 27838 42367 27936 4 gnd
port 2 nsew
rlabel metal3 s 42269 26811 42367 26909 4 gnd
port 2 nsew
rlabel metal3 s 42269 27364 42367 27462 4 gnd
port 2 nsew
rlabel metal3 s 42269 29418 42367 29516 4 gnd
port 2 nsew
rlabel metal3 s 42269 33921 42367 34019 4 gnd
port 2 nsew
rlabel metal3 s 42269 37634 42367 37732 4 gnd
port 2 nsew
rlabel metal3 s 42269 26258 42367 26356 4 gnd
port 2 nsew
rlabel metal3 s 42269 29181 42367 29279 4 gnd
port 2 nsew
rlabel metal3 s 42269 38898 42367 38996 4 gnd
port 2 nsew
rlabel metal3 s 42269 34711 42367 34809 4 gnd
port 2 nsew
rlabel metal3 s 42269 28154 42367 28252 4 gnd
port 2 nsew
rlabel metal3 s 42269 31314 42367 31412 4 gnd
port 2 nsew
rlabel metal3 s 14741 51862 14839 51960 4 vdd
port 1 nsew
rlabel metal3 s 13493 51862 13591 51960 4 vdd
port 1 nsew
rlabel metal3 s 17861 51862 17959 51960 4 vdd
port 1 nsew
rlabel metal3 s 19733 51862 19831 51960 4 vdd
port 1 nsew
rlabel metal3 s 14117 51862 14215 51960 4 vdd
port 1 nsew
rlabel metal3 s 20981 51862 21079 51960 4 vdd
port 1 nsew
rlabel metal3 s 18485 51862 18583 51960 4 vdd
port 1 nsew
rlabel metal3 s 15365 51862 15463 51960 4 vdd
port 1 nsew
rlabel metal3 s 12245 51862 12343 51960 4 vdd
port 1 nsew
rlabel metal3 s 12869 51862 12967 51960 4 vdd
port 1 nsew
rlabel metal3 s 16613 51862 16711 51960 4 vdd
port 1 nsew
rlabel metal3 s 20357 51862 20455 51960 4 vdd
port 1 nsew
rlabel metal3 s 15989 51862 16087 51960 4 vdd
port 1 nsew
rlabel metal3 s 19109 51862 19207 51960 4 vdd
port 1 nsew
rlabel metal3 s 10997 51862 11095 51960 4 vdd
port 1 nsew
rlabel metal3 s 17237 51862 17335 51960 4 vdd
port 1 nsew
rlabel metal3 s 11621 51862 11719 51960 4 vdd
port 1 nsew
rlabel metal3 s -49 51648 49 51746 4 gnd
port 2 nsew
rlabel metal3 s 5381 51862 5479 51960 4 vdd
port 1 nsew
rlabel metal3 s 10373 51862 10471 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 42848 415 42946 4 gnd
port 2 nsew
rlabel metal3 s 317 49721 415 49819 4 gnd
port 2 nsew
rlabel metal3 s 317 46798 415 46896 4 gnd
port 2 nsew
rlabel metal3 s 317 43954 415 44052 4 gnd
port 2 nsew
rlabel metal3 s 317 44428 415 44526 4 gnd
port 2 nsew
rlabel metal3 s 317 50511 415 50609 4 gnd
port 2 nsew
rlabel metal3 s 317 39451 415 39549 4 gnd
port 2 nsew
rlabel metal3 s 317 39214 415 39312 4 gnd
port 2 nsew
rlabel metal3 s 7877 51862 7975 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 40241 415 40339 4 gnd
port 2 nsew
rlabel metal3 s 317 42374 415 42472 4 gnd
port 2 nsew
rlabel metal3 s 317 47114 415 47212 4 gnd
port 2 nsew
rlabel metal3 s 317 50274 415 50372 4 gnd
port 2 nsew
rlabel metal3 s 1013 51862 1111 51960 4 vdd
port 1 nsew
rlabel metal3 s 4757 51862 4855 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 48931 415 49029 4 gnd
port 2 nsew
rlabel metal3 s 317 41268 415 41366 4 gnd
port 2 nsew
rlabel metal3 s 317 44744 415 44842 4 gnd
port 2 nsew
rlabel metal3 s 317 45534 415 45632 4 gnd
port 2 nsew
rlabel metal3 s 317 49484 415 49582 4 gnd
port 2 nsew
rlabel metal3 s 8501 51862 8599 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 46008 415 46106 4 gnd
port 2 nsew
rlabel metal3 s 317 49168 415 49266 4 gnd
port 2 nsew
rlabel metal3 s 317 44981 415 45079 4 gnd
port 2 nsew
rlabel metal3 s 317 39688 415 39786 4 gnd
port 2 nsew
rlabel metal3 s 317 42058 415 42156 4 gnd
port 2 nsew
rlabel metal3 s 3509 51862 3607 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 43401 415 43499 4 gnd
port 2 nsew
rlabel metal3 s 317 47904 415 48002 4 gnd
port 2 nsew
rlabel metal3 s 317 43638 415 43736 4 gnd
port 2 nsew
rlabel metal3 s 9749 51862 9847 51960 4 vdd
port 1 nsew
rlabel metal3 s 9125 51862 9223 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 47588 415 47686 4 gnd
port 2 nsew
rlabel metal3 s 2261 51862 2359 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 40004 415 40102 4 gnd
port 2 nsew
rlabel metal3 s 317 49958 415 50056 4 gnd
port 2 nsew
rlabel metal3 s 317 46324 415 46422 4 gnd
port 2 nsew
rlabel metal3 s 317 43164 415 43262 4 gnd
port 2 nsew
rlabel metal3 s 317 41031 415 41129 4 gnd
port 2 nsew
rlabel metal3 s 317 47351 415 47449 4 gnd
port 2 nsew
rlabel metal3 s 6629 51862 6727 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 50748 415 50846 4 gnd
port 2 nsew
rlabel metal3 s 317 46561 415 46659 4 gnd
port 2 nsew
rlabel metal3 s 7253 51862 7351 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 51064 415 51162 4 gnd
port 2 nsew
rlabel metal3 s 317 41821 415 41919 4 gnd
port 2 nsew
rlabel metal3 s 1637 51862 1735 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 44191 415 44289 4 gnd
port 2 nsew
rlabel metal3 s 317 51301 415 51399 4 gnd
port 2 nsew
rlabel metal3 s 317 41584 415 41682 4 gnd
port 2 nsew
rlabel metal3 s 317 42611 415 42709 4 gnd
port 2 nsew
rlabel metal3 s 317 45771 415 45869 4 gnd
port 2 nsew
rlabel metal3 s 4133 51862 4231 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 45218 415 45316 4 gnd
port 2 nsew
rlabel metal3 s 317 48141 415 48239 4 gnd
port 2 nsew
rlabel metal3 s 6005 51862 6103 51960 4 vdd
port 1 nsew
rlabel metal3 s 2885 51862 2983 51960 4 vdd
port 1 nsew
rlabel metal3 s 317 48378 415 48476 4 gnd
port 2 nsew
rlabel metal3 s 317 40478 415 40576 4 gnd
port 2 nsew
rlabel metal3 s 317 48694 415 48792 4 gnd
port 2 nsew
rlabel metal3 s 317 40794 415 40892 4 gnd
port 2 nsew
rlabel metal3 s 317 38898 415 38996 4 gnd
port 2 nsew
rlabel metal3 s 317 28154 415 28252 4 gnd
port 2 nsew
rlabel metal3 s 317 38661 415 38759 4 gnd
port 2 nsew
rlabel metal3 s 317 28391 415 28489 4 gnd
port 2 nsew
rlabel metal3 s 317 34158 415 34256 4 gnd
port 2 nsew
rlabel metal3 s 317 27048 415 27146 4 gnd
port 2 nsew
rlabel metal3 s 317 30761 415 30859 4 gnd
port 2 nsew
rlabel metal3 s 317 30524 415 30622 4 gnd
port 2 nsew
rlabel metal3 s 317 33921 415 34019 4 gnd
port 2 nsew
rlabel metal3 s 317 37081 415 37179 4 gnd
port 2 nsew
rlabel metal3 s 317 26811 415 26909 4 gnd
port 2 nsew
rlabel metal3 s 317 36291 415 36389 4 gnd
port 2 nsew
rlabel metal3 s 317 37871 415 37969 4 gnd
port 2 nsew
rlabel metal3 s 317 32894 415 32992 4 gnd
port 2 nsew
rlabel metal3 s 317 32578 415 32676 4 gnd
port 2 nsew
rlabel metal3 s 317 31314 415 31412 4 gnd
port 2 nsew
rlabel metal3 s 317 26258 415 26356 4 gnd
port 2 nsew
rlabel metal3 s 317 34474 415 34572 4 gnd
port 2 nsew
rlabel metal3 s 317 37318 415 37416 4 gnd
port 2 nsew
rlabel metal3 s 317 33684 415 33782 4 gnd
port 2 nsew
rlabel metal3 s 317 29734 415 29832 4 gnd
port 2 nsew
rlabel metal3 s 317 36528 415 36626 4 gnd
port 2 nsew
rlabel metal3 s 317 28628 415 28726 4 gnd
port 2 nsew
rlabel metal3 s 317 36844 415 36942 4 gnd
port 2 nsew
rlabel metal3 s 317 33131 415 33229 4 gnd
port 2 nsew
rlabel metal3 s 317 38108 415 38206 4 gnd
port 2 nsew
rlabel metal3 s 317 36054 415 36152 4 gnd
port 2 nsew
rlabel metal3 s 317 26574 415 26672 4 gnd
port 2 nsew
rlabel metal3 s 317 30998 415 31096 4 gnd
port 2 nsew
rlabel metal3 s 317 29181 415 29279 4 gnd
port 2 nsew
rlabel metal3 s 317 32341 415 32439 4 gnd
port 2 nsew
rlabel metal3 s 317 28944 415 29042 4 gnd
port 2 nsew
rlabel metal3 s 317 35501 415 35599 4 gnd
port 2 nsew
rlabel metal3 s 317 27838 415 27936 4 gnd
port 2 nsew
rlabel metal3 s 317 32104 415 32202 4 gnd
port 2 nsew
rlabel metal3 s 317 31551 415 31649 4 gnd
port 2 nsew
rlabel metal3 s 317 30208 415 30306 4 gnd
port 2 nsew
rlabel metal3 s 317 35264 415 35362 4 gnd
port 2 nsew
rlabel metal3 s 317 27601 415 27699 4 gnd
port 2 nsew
rlabel metal3 s 317 35738 415 35836 4 gnd
port 2 nsew
rlabel metal3 s 317 29971 415 30069 4 gnd
port 2 nsew
rlabel metal3 s 317 38424 415 38522 4 gnd
port 2 nsew
rlabel metal3 s 317 37634 415 37732 4 gnd
port 2 nsew
rlabel metal3 s 317 33368 415 33466 4 gnd
port 2 nsew
rlabel metal3 s 317 34948 415 35046 4 gnd
port 2 nsew
rlabel metal3 s 317 34711 415 34809 4 gnd
port 2 nsew
rlabel metal3 s 317 27364 415 27462 4 gnd
port 2 nsew
rlabel metal3 s 317 31788 415 31886 4 gnd
port 2 nsew
rlabel metal3 s 317 29418 415 29516 4 gnd
port 2 nsew
rlabel metal3 s 317 13618 415 13716 4 gnd
port 2 nsew
rlabel metal3 s 317 14171 415 14269 4 gnd
port 2 nsew
rlabel metal3 s 317 14408 415 14506 4 gnd
port 2 nsew
rlabel metal3 s 317 14724 415 14822 4 gnd
port 2 nsew
rlabel metal3 s 317 16778 415 16876 4 gnd
port 2 nsew
rlabel metal3 s 317 25784 415 25882 4 gnd
port 2 nsew
rlabel metal3 s 317 17568 415 17666 4 gnd
port 2 nsew
rlabel metal3 s 317 22861 415 22959 4 gnd
port 2 nsew
rlabel metal3 s 317 20728 415 20826 4 gnd
port 2 nsew
rlabel metal3 s 317 19701 415 19799 4 gnd
port 2 nsew
rlabel metal3 s 317 15514 415 15612 4 gnd
port 2 nsew
rlabel metal3 s 317 15198 415 15296 4 gnd
port 2 nsew
rlabel metal3 s 317 23414 415 23512 4 gnd
port 2 nsew
rlabel metal3 s 317 26021 415 26119 4 gnd
port 2 nsew
rlabel metal3 s 317 18121 415 18219 4 gnd
port 2 nsew
rlabel metal3 s 317 22308 415 22406 4 gnd
port 2 nsew
rlabel metal3 s 317 13144 415 13242 4 gnd
port 2 nsew
rlabel metal3 s 317 25231 415 25329 4 gnd
port 2 nsew
rlabel metal3 s 317 22624 415 22722 4 gnd
port 2 nsew
rlabel metal3 s 317 24441 415 24539 4 gnd
port 2 nsew
rlabel metal3 s 317 20254 415 20352 4 gnd
port 2 nsew
rlabel metal3 s 317 23651 415 23749 4 gnd
port 2 nsew
rlabel metal3 s 317 16304 415 16402 4 gnd
port 2 nsew
rlabel metal3 s 317 24994 415 25092 4 gnd
port 2 nsew
rlabel metal3 s 317 18674 415 18772 4 gnd
port 2 nsew
rlabel metal3 s 317 15751 415 15849 4 gnd
port 2 nsew
rlabel metal3 s 317 21281 415 21379 4 gnd
port 2 nsew
rlabel metal3 s 317 18911 415 19009 4 gnd
port 2 nsew
rlabel metal3 s 317 17094 415 17192 4 gnd
port 2 nsew
rlabel metal3 s 317 17884 415 17982 4 gnd
port 2 nsew
rlabel metal3 s 317 19464 415 19562 4 gnd
port 2 nsew
rlabel metal3 s 317 13934 415 14032 4 gnd
port 2 nsew
rlabel metal3 s 317 21044 415 21142 4 gnd
port 2 nsew
rlabel metal3 s 317 14961 415 15059 4 gnd
port 2 nsew
rlabel metal3 s 317 21518 415 21616 4 gnd
port 2 nsew
rlabel metal3 s 317 19938 415 20036 4 gnd
port 2 nsew
rlabel metal3 s 317 18358 415 18456 4 gnd
port 2 nsew
rlabel metal3 s 317 21834 415 21932 4 gnd
port 2 nsew
rlabel metal3 s 317 23098 415 23196 4 gnd
port 2 nsew
rlabel metal3 s 317 16541 415 16639 4 gnd
port 2 nsew
rlabel metal3 s 317 24678 415 24776 4 gnd
port 2 nsew
rlabel metal3 s 317 23888 415 23986 4 gnd
port 2 nsew
rlabel metal3 s 317 17331 415 17429 4 gnd
port 2 nsew
rlabel metal3 s 317 24204 415 24302 4 gnd
port 2 nsew
rlabel metal3 s 317 20491 415 20589 4 gnd
port 2 nsew
rlabel metal3 s 317 13381 415 13479 4 gnd
port 2 nsew
rlabel metal3 s 317 25468 415 25566 4 gnd
port 2 nsew
rlabel metal3 s 317 15988 415 16086 4 gnd
port 2 nsew
rlabel metal3 s 317 22071 415 22169 4 gnd
port 2 nsew
rlabel metal3 s 317 19148 415 19246 4 gnd
port 2 nsew
rlabel metal3 s 317 9431 415 9529 4 gnd
port 2 nsew
rlabel metal3 s 6629 180 6727 278 4 vdd
port 1 nsew
rlabel metal3 s 6005 180 6103 278 4 vdd
port 1 nsew
rlabel metal3 s 317 2321 415 2419 4 gnd
port 2 nsew
rlabel metal3 s 317 4138 415 4236 4 gnd
port 2 nsew
rlabel metal3 s 317 9984 415 10082 4 gnd
port 2 nsew
rlabel metal3 s 317 10221 415 10319 4 gnd
port 2 nsew
rlabel metal3 s 317 11011 415 11109 4 gnd
port 2 nsew
rlabel metal3 s 317 11248 415 11346 4 gnd
port 2 nsew
rlabel metal3 s 317 11564 415 11662 4 gnd
port 2 nsew
rlabel metal3 s 317 11801 415 11899 4 gnd
port 2 nsew
rlabel metal3 s 4757 180 4855 278 4 vdd
port 1 nsew
rlabel metal3 s 317 2084 415 2182 4 gnd
port 2 nsew
rlabel metal3 s 317 6508 415 6606 4 gnd
port 2 nsew
rlabel metal3 s 317 10774 415 10872 4 gnd
port 2 nsew
rlabel metal3 s 317 6034 415 6132 4 gnd
port 2 nsew
rlabel metal3 s 9749 180 9847 278 4 vdd
port 1 nsew
rlabel metal3 s 317 8088 415 8186 4 gnd
port 2 nsew
rlabel metal3 s 1637 180 1735 278 4 vdd
port 1 nsew
rlabel metal3 s -49 614 49 712 4 gnd
port 2 nsew
rlabel metal3 s 317 8641 415 8739 4 gnd
port 2 nsew
rlabel metal3 s 317 8878 415 8976 4 gnd
port 2 nsew
rlabel metal3 s 10373 180 10471 278 4 vdd
port 1 nsew
rlabel metal3 s 4133 180 4231 278 4 vdd
port 1 nsew
rlabel metal3 s 317 5481 415 5579 4 gnd
port 2 nsew
rlabel metal3 s 317 9194 415 9292 4 gnd
port 2 nsew
rlabel metal3 s 8501 180 8599 278 4 vdd
port 1 nsew
rlabel metal3 s 317 5718 415 5816 4 gnd
port 2 nsew
rlabel metal3 s 317 5244 415 5342 4 gnd
port 2 nsew
rlabel metal3 s 317 12038 415 12136 4 gnd
port 2 nsew
rlabel metal3 s 317 1768 415 1866 4 gnd
port 2 nsew
rlabel metal3 s 317 10458 415 10556 4 gnd
port 2 nsew
rlabel metal3 s 317 9668 415 9766 4 gnd
port 2 nsew
rlabel metal3 s 7877 180 7975 278 4 vdd
port 1 nsew
rlabel metal3 s 317 978 415 1076 4 gnd
port 2 nsew
rlabel metal3 s 2885 180 2983 278 4 vdd
port 1 nsew
rlabel metal3 s 317 7851 415 7949 4 gnd
port 2 nsew
rlabel metal3 s 2261 180 2359 278 4 vdd
port 1 nsew
rlabel metal3 s 9125 180 9223 278 4 vdd
port 1 nsew
rlabel metal3 s 317 7614 415 7712 4 gnd
port 2 nsew
rlabel metal3 s 317 4928 415 5026 4 gnd
port 2 nsew
rlabel metal3 s 317 2558 415 2656 4 gnd
port 2 nsew
rlabel metal3 s 317 8404 415 8502 4 gnd
port 2 nsew
rlabel metal3 s 317 2874 415 2972 4 gnd
port 2 nsew
rlabel metal3 s 317 12354 415 12452 4 gnd
port 2 nsew
rlabel metal3 s 317 1531 415 1629 4 gnd
port 2 nsew
rlabel metal3 s 317 6824 415 6922 4 gnd
port 2 nsew
rlabel metal3 s 5381 180 5479 278 4 vdd
port 1 nsew
rlabel metal3 s 317 4454 415 4552 4 gnd
port 2 nsew
rlabel metal3 s 317 1294 415 1392 4 gnd
port 2 nsew
rlabel metal3 s 317 4691 415 4789 4 gnd
port 2 nsew
rlabel metal3 s 317 3348 415 3446 4 gnd
port 2 nsew
rlabel metal3 s 317 6271 415 6369 4 gnd
port 2 nsew
rlabel metal3 s 317 7061 415 7159 4 gnd
port 2 nsew
rlabel metal3 s 7253 180 7351 278 4 vdd
port 1 nsew
rlabel metal3 s 317 3901 415 3999 4 gnd
port 2 nsew
rlabel metal3 s 1013 180 1111 278 4 vdd
port 1 nsew
rlabel metal3 s 317 12828 415 12926 4 gnd
port 2 nsew
rlabel metal3 s 317 741 415 839 4 gnd
port 2 nsew
rlabel metal3 s 317 12591 415 12689 4 gnd
port 2 nsew
rlabel metal3 s 317 3111 415 3209 4 gnd
port 2 nsew
rlabel metal3 s 317 3664 415 3762 4 gnd
port 2 nsew
rlabel metal3 s 3509 180 3607 278 4 vdd
port 1 nsew
rlabel metal3 s 317 7298 415 7396 4 gnd
port 2 nsew
rlabel metal3 s 20981 180 21079 278 4 vdd
port 1 nsew
rlabel metal3 s 19109 180 19207 278 4 vdd
port 1 nsew
rlabel metal3 s 15989 180 16087 278 4 vdd
port 1 nsew
rlabel metal3 s 17237 180 17335 278 4 vdd
port 1 nsew
rlabel metal3 s 19733 180 19831 278 4 vdd
port 1 nsew
rlabel metal3 s 10997 180 11095 278 4 vdd
port 1 nsew
rlabel metal3 s 12245 180 12343 278 4 vdd
port 1 nsew
rlabel metal3 s 20357 180 20455 278 4 vdd
port 1 nsew
rlabel metal3 s 13493 180 13591 278 4 vdd
port 1 nsew
rlabel metal3 s 16613 180 16711 278 4 vdd
port 1 nsew
rlabel metal3 s 12869 180 12967 278 4 vdd
port 1 nsew
rlabel metal3 s 14741 180 14839 278 4 vdd
port 1 nsew
rlabel metal3 s 14117 180 14215 278 4 vdd
port 1 nsew
rlabel metal3 s 11621 180 11719 278 4 vdd
port 1 nsew
rlabel metal3 s 17861 180 17959 278 4 vdd
port 1 nsew
rlabel metal3 s 15365 180 15463 278 4 vdd
port 1 nsew
rlabel metal3 s 18485 180 18583 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 15988 42367 16086 4 gnd
port 2 nsew
rlabel metal3 s 42269 23414 42367 23512 4 gnd
port 2 nsew
rlabel metal3 s 42269 19938 42367 20036 4 gnd
port 2 nsew
rlabel metal3 s 42269 23651 42367 23749 4 gnd
port 2 nsew
rlabel metal3 s 42269 14408 42367 14506 4 gnd
port 2 nsew
rlabel metal3 s 42269 14171 42367 14269 4 gnd
port 2 nsew
rlabel metal3 s 42269 24204 42367 24302 4 gnd
port 2 nsew
rlabel metal3 s 42269 13144 42367 13242 4 gnd
port 2 nsew
rlabel metal3 s 42269 22624 42367 22722 4 gnd
port 2 nsew
rlabel metal3 s 42269 18121 42367 18219 4 gnd
port 2 nsew
rlabel metal3 s 42269 14961 42367 15059 4 gnd
port 2 nsew
rlabel metal3 s 42269 21281 42367 21379 4 gnd
port 2 nsew
rlabel metal3 s 42269 20491 42367 20589 4 gnd
port 2 nsew
rlabel metal3 s 42269 17331 42367 17429 4 gnd
port 2 nsew
rlabel metal3 s 42269 23098 42367 23196 4 gnd
port 2 nsew
rlabel metal3 s 42269 19701 42367 19799 4 gnd
port 2 nsew
rlabel metal3 s 42269 17568 42367 17666 4 gnd
port 2 nsew
rlabel metal3 s 42269 24441 42367 24539 4 gnd
port 2 nsew
rlabel metal3 s 42269 17094 42367 17192 4 gnd
port 2 nsew
rlabel metal3 s 42269 18911 42367 19009 4 gnd
port 2 nsew
rlabel metal3 s 42269 13381 42367 13479 4 gnd
port 2 nsew
rlabel metal3 s 42269 22861 42367 22959 4 gnd
port 2 nsew
rlabel metal3 s 42269 25468 42367 25566 4 gnd
port 2 nsew
rlabel metal3 s 42269 22071 42367 22169 4 gnd
port 2 nsew
rlabel metal3 s 42269 26021 42367 26119 4 gnd
port 2 nsew
rlabel metal3 s 42269 18358 42367 18456 4 gnd
port 2 nsew
rlabel metal3 s 42269 16541 42367 16639 4 gnd
port 2 nsew
rlabel metal3 s 42269 15751 42367 15849 4 gnd
port 2 nsew
rlabel metal3 s 42269 21834 42367 21932 4 gnd
port 2 nsew
rlabel metal3 s 42269 25231 42367 25329 4 gnd
port 2 nsew
rlabel metal3 s 42269 25784 42367 25882 4 gnd
port 2 nsew
rlabel metal3 s 42269 18674 42367 18772 4 gnd
port 2 nsew
rlabel metal3 s 42269 17884 42367 17982 4 gnd
port 2 nsew
rlabel metal3 s 42269 20728 42367 20826 4 gnd
port 2 nsew
rlabel metal3 s 42269 24994 42367 25092 4 gnd
port 2 nsew
rlabel metal3 s 42269 21044 42367 21142 4 gnd
port 2 nsew
rlabel metal3 s 42269 24678 42367 24776 4 gnd
port 2 nsew
rlabel metal3 s 42269 21518 42367 21616 4 gnd
port 2 nsew
rlabel metal3 s 42269 19148 42367 19246 4 gnd
port 2 nsew
rlabel metal3 s 42269 16304 42367 16402 4 gnd
port 2 nsew
rlabel metal3 s 42269 13618 42367 13716 4 gnd
port 2 nsew
rlabel metal3 s 42269 13934 42367 14032 4 gnd
port 2 nsew
rlabel metal3 s 42269 15514 42367 15612 4 gnd
port 2 nsew
rlabel metal3 s 42269 16778 42367 16876 4 gnd
port 2 nsew
rlabel metal3 s 42269 20254 42367 20352 4 gnd
port 2 nsew
rlabel metal3 s 42269 14724 42367 14822 4 gnd
port 2 nsew
rlabel metal3 s 42269 15198 42367 15296 4 gnd
port 2 nsew
rlabel metal3 s 42269 23888 42367 23986 4 gnd
port 2 nsew
rlabel metal3 s 42269 19464 42367 19562 4 gnd
port 2 nsew
rlabel metal3 s 42269 22308 42367 22406 4 gnd
port 2 nsew
rlabel metal3 s 24725 180 24823 278 4 vdd
port 1 nsew
rlabel metal3 s 29093 180 29191 278 4 vdd
port 1 nsew
rlabel metal3 s 30341 180 30439 278 4 vdd
port 1 nsew
rlabel metal3 s 26597 180 26695 278 4 vdd
port 1 nsew
rlabel metal3 s 25973 180 26071 278 4 vdd
port 1 nsew
rlabel metal3 s 22853 180 22951 278 4 vdd
port 1 nsew
rlabel metal3 s 27845 180 27943 278 4 vdd
port 1 nsew
rlabel metal3 s 21605 180 21703 278 4 vdd
port 1 nsew
rlabel metal3 s 27221 180 27319 278 4 vdd
port 1 nsew
rlabel metal3 s 22229 180 22327 278 4 vdd
port 1 nsew
rlabel metal3 s 24101 180 24199 278 4 vdd
port 1 nsew
rlabel metal3 s 29717 180 29815 278 4 vdd
port 1 nsew
rlabel metal3 s 23477 180 23575 278 4 vdd
port 1 nsew
rlabel metal3 s 30965 180 31063 278 4 vdd
port 1 nsew
rlabel metal3 s 31589 180 31687 278 4 vdd
port 1 nsew
rlabel metal3 s 25349 180 25447 278 4 vdd
port 1 nsew
rlabel metal3 s 28469 180 28567 278 4 vdd
port 1 nsew
rlabel metal3 s 35957 180 36055 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 6824 42367 6922 4 gnd
port 2 nsew
rlabel metal3 s 42269 12591 42367 12689 4 gnd
port 2 nsew
rlabel metal3 s 41573 180 41671 278 4 vdd
port 1 nsew
rlabel metal3 s 35333 180 35431 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 4691 42367 4789 4 gnd
port 2 nsew
rlabel metal3 s 42269 11011 42367 11109 4 gnd
port 2 nsew
rlabel metal3 s 42269 5481 42367 5579 4 gnd
port 2 nsew
rlabel metal3 s 42269 11248 42367 11346 4 gnd
port 2 nsew
rlabel metal3 s 42269 12354 42367 12452 4 gnd
port 2 nsew
rlabel metal3 s 42269 4454 42367 4552 4 gnd
port 2 nsew
rlabel metal3 s 42269 6508 42367 6606 4 gnd
port 2 nsew
rlabel metal3 s 42269 9194 42367 9292 4 gnd
port 2 nsew
rlabel metal3 s 37829 180 37927 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 2874 42367 2972 4 gnd
port 2 nsew
rlabel metal3 s 42269 2321 42367 2419 4 gnd
port 2 nsew
rlabel metal3 s 42269 7851 42367 7949 4 gnd
port 2 nsew
rlabel metal3 s 32213 180 32311 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 7061 42367 7159 4 gnd
port 2 nsew
rlabel metal3 s 42269 12828 42367 12926 4 gnd
port 2 nsew
rlabel metal3 s 42269 1294 42367 1392 4 gnd
port 2 nsew
rlabel metal3 s 42269 3348 42367 3446 4 gnd
port 2 nsew
rlabel metal3 s 42269 5718 42367 5816 4 gnd
port 2 nsew
rlabel metal3 s 40325 180 40423 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 978 42367 1076 4 gnd
port 2 nsew
rlabel metal3 s 42269 8404 42367 8502 4 gnd
port 2 nsew
rlabel metal3 s 32837 180 32935 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 9668 42367 9766 4 gnd
port 2 nsew
rlabel metal3 s 42269 9984 42367 10082 4 gnd
port 2 nsew
rlabel metal3 s 42269 11801 42367 11899 4 gnd
port 2 nsew
rlabel metal3 s 42635 614 42733 712 4 gnd
port 2 nsew
rlabel metal3 s 42269 8878 42367 8976 4 gnd
port 2 nsew
rlabel metal3 s 42269 9431 42367 9529 4 gnd
port 2 nsew
rlabel metal3 s 42269 10221 42367 10319 4 gnd
port 2 nsew
rlabel metal3 s 42269 6271 42367 6369 4 gnd
port 2 nsew
rlabel metal3 s 42269 10774 42367 10872 4 gnd
port 2 nsew
rlabel metal3 s 36581 180 36679 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 3901 42367 3999 4 gnd
port 2 nsew
rlabel metal3 s 34085 180 34183 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 1531 42367 1629 4 gnd
port 2 nsew
rlabel metal3 s 39701 180 39799 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 4928 42367 5026 4 gnd
port 2 nsew
rlabel metal3 s 42269 10458 42367 10556 4 gnd
port 2 nsew
rlabel metal3 s 42269 8088 42367 8186 4 gnd
port 2 nsew
rlabel metal3 s 42269 4138 42367 4236 4 gnd
port 2 nsew
rlabel metal3 s 42269 6034 42367 6132 4 gnd
port 2 nsew
rlabel metal3 s 42269 11564 42367 11662 4 gnd
port 2 nsew
rlabel metal3 s 39077 180 39175 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 7614 42367 7712 4 gnd
port 2 nsew
rlabel metal3 s 42269 741 42367 839 4 gnd
port 2 nsew
rlabel metal3 s 42269 2558 42367 2656 4 gnd
port 2 nsew
rlabel metal3 s 42269 2084 42367 2182 4 gnd
port 2 nsew
rlabel metal3 s 42269 5244 42367 5342 4 gnd
port 2 nsew
rlabel metal3 s 42269 3111 42367 3209 4 gnd
port 2 nsew
rlabel metal3 s 42269 8641 42367 8739 4 gnd
port 2 nsew
rlabel metal3 s 42269 7298 42367 7396 4 gnd
port 2 nsew
rlabel metal3 s 40949 180 41047 278 4 vdd
port 1 nsew
rlabel metal3 s 38453 180 38551 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 1768 42367 1866 4 gnd
port 2 nsew
rlabel metal3 s 42269 3664 42367 3762 4 gnd
port 2 nsew
rlabel metal3 s 34709 180 34807 278 4 vdd
port 1 nsew
rlabel metal3 s 37205 180 37303 278 4 vdd
port 1 nsew
rlabel metal3 s 42269 12038 42367 12136 4 gnd
port 2 nsew
rlabel metal3 s 33461 180 33559 278 4 vdd
port 1 nsew
rlabel metal2 s 41496 30219 41604 30295 4 gnd
port 2 nsew
rlabel metal2 s 41496 43175 41604 43251 4 gnd
port 2 nsew
rlabel metal2 s 41496 33379 41604 33455 4 gnd
port 2 nsew
rlabel metal2 s 41496 34959 41604 35035 4 gnd
port 2 nsew
rlabel metal2 s 41496 31799 41604 31875 4 gnd
port 2 nsew
rlabel metal2 s 41496 50285 41604 50361 4 gnd
port 2 nsew
rlabel metal2 s 41496 46335 41604 46411 4 gnd
port 2 nsew
rlabel metal2 s 41496 26015 41604 26125 4 gnd
port 2 nsew
rlabel metal2 s 41496 35495 41604 35605 4 gnd
port 2 nsew
rlabel metal2 s 41496 26805 41604 26915 4 gnd
port 2 nsew
rlabel metal2 s 41496 28165 41604 28241 4 gnd
port 2 nsew
rlabel metal2 s 41496 41279 41604 41355 4 gnd
port 2 nsew
rlabel metal2 s 41496 42859 41604 42935 4 gnd
port 2 nsew
rlabel metal2 s 41496 49179 41604 49255 4 gnd
port 2 nsew
rlabel metal2 s 41496 48389 41604 48465 4 gnd
port 2 nsew
rlabel metal2 s 41496 48705 41604 48781 4 gnd
port 2 nsew
rlabel metal2 s 41496 51549 41604 51625 4 gnd
port 2 nsew
rlabel metal2 s 41496 45545 41604 45621 4 gnd
port 2 nsew
rlabel metal2 s 41496 34705 41604 34815 4 gnd
port 2 nsew
rlabel metal2 s 41496 26585 41604 26661 4 gnd
port 2 nsew
rlabel metal2 s 41496 47125 41604 47201 4 gnd
port 2 nsew
rlabel metal2 s 41496 51295 41604 51405 4 gnd
port 2 nsew
rlabel metal2 s 41496 27595 41604 27705 4 gnd
port 2 nsew
rlabel metal2 s 41496 41815 41604 41925 4 gnd
port 2 nsew
rlabel metal2 s 41496 50505 41604 50615 4 gnd
port 2 nsew
rlabel metal2 s 41496 32589 41604 32665 4 gnd
port 2 nsew
rlabel metal2 s 41496 51075 41604 51151 4 gnd
port 2 nsew
rlabel metal2 s 41496 38909 41604 38985 4 gnd
port 2 nsew
rlabel metal2 s 41496 44975 41604 45085 4 gnd
port 2 nsew
rlabel metal2 s 41496 37865 41604 37975 4 gnd
port 2 nsew
rlabel metal2 s 41496 34485 41604 34561 4 gnd
port 2 nsew
rlabel metal2 s 41496 45229 41604 45305 4 gnd
port 2 nsew
rlabel metal2 s 41496 48135 41604 48245 4 gnd
port 2 nsew
rlabel metal2 s 41496 46555 41604 46665 4 gnd
port 2 nsew
rlabel metal2 s 41496 33695 41604 33771 4 gnd
port 2 nsew
rlabel metal2 s 41496 33915 41604 34025 4 gnd
port 2 nsew
rlabel metal2 s 41496 30755 41604 30865 4 gnd
port 2 nsew
rlabel metal2 s 41496 32905 41604 32981 4 gnd
port 2 nsew
rlabel metal2 s 41496 35749 41604 35825 4 gnd
port 2 nsew
rlabel metal2 s 41496 36065 41604 36141 4 gnd
port 2 nsew
rlabel metal2 s 41496 32115 41604 32191 4 gnd
port 2 nsew
rlabel metal2 s 41496 41025 41604 41135 4 gnd
port 2 nsew
rlabel metal2 s 41496 46019 41604 46095 4 gnd
port 2 nsew
rlabel metal2 s 41496 31325 41604 31401 4 gnd
port 2 nsew
rlabel metal2 s 41496 49715 41604 49825 4 gnd
port 2 nsew
rlabel metal2 s 41496 38435 41604 38511 4 gnd
port 2 nsew
rlabel metal2 s 41496 44439 41604 44515 4 gnd
port 2 nsew
rlabel metal2 s 41496 28955 41604 29031 4 gnd
port 2 nsew
rlabel metal2 s 41496 49969 41604 50045 4 gnd
port 2 nsew
rlabel metal2 s 41496 29965 41604 30075 4 gnd
port 2 nsew
rlabel metal2 s 41496 26269 41604 26345 4 gnd
port 2 nsew
rlabel metal2 s 41496 50759 41604 50835 4 gnd
port 2 nsew
rlabel metal2 s 41496 47599 41604 47675 4 gnd
port 2 nsew
rlabel metal2 s 41496 37645 41604 37721 4 gnd
port 2 nsew
rlabel metal2 s 41496 29745 41604 29821 4 gnd
port 2 nsew
rlabel metal2 s 41496 45765 41604 45875 4 gnd
port 2 nsew
rlabel metal2 s 41496 42385 41604 42461 4 gnd
port 2 nsew
rlabel metal2 s 41496 27849 41604 27925 4 gnd
port 2 nsew
rlabel metal2 s 41496 43395 41604 43505 4 gnd
port 2 nsew
rlabel metal2 s 41496 31545 41604 31655 4 gnd
port 2 nsew
rlabel metal2 s 41496 37075 41604 37185 4 gnd
port 2 nsew
rlabel metal2 s 41496 36855 41604 36931 4 gnd
port 2 nsew
rlabel metal2 s 41496 30535 41604 30611 4 gnd
port 2 nsew
rlabel metal2 s 41496 34169 41604 34245 4 gnd
port 2 nsew
rlabel metal2 s 41496 29175 41604 29285 4 gnd
port 2 nsew
rlabel metal2 s 41496 39699 41604 39775 4 gnd
port 2 nsew
rlabel metal2 s 41496 39225 41604 39301 4 gnd
port 2 nsew
rlabel metal2 s 41496 48925 41604 49035 4 gnd
port 2 nsew
rlabel metal2 s 41496 28385 41604 28495 4 gnd
port 2 nsew
rlabel metal2 s 41496 41595 41604 41671 4 gnd
port 2 nsew
rlabel metal2 s 41496 38119 41604 38195 4 gnd
port 2 nsew
rlabel metal2 s 41496 28639 41604 28715 4 gnd
port 2 nsew
rlabel metal2 s 41496 39445 41604 39555 4 gnd
port 2 nsew
rlabel metal2 s 41496 42605 41604 42715 4 gnd
port 2 nsew
rlabel metal2 s 41496 36539 41604 36615 4 gnd
port 2 nsew
rlabel metal2 s 41496 32335 41604 32445 4 gnd
port 2 nsew
rlabel metal2 s 41496 40489 41604 40565 4 gnd
port 2 nsew
rlabel metal2 s 41496 38655 41604 38765 4 gnd
port 2 nsew
rlabel metal2 s 41496 44185 41604 44295 4 gnd
port 2 nsew
rlabel metal2 s 41496 49495 41604 49571 4 gnd
port 2 nsew
rlabel metal2 s 41496 40015 41604 40091 4 gnd
port 2 nsew
rlabel metal2 s 41496 43649 41604 43725 4 gnd
port 2 nsew
rlabel metal2 s 41496 43965 41604 44041 4 gnd
port 2 nsew
rlabel metal2 s 41496 27375 41604 27451 4 gnd
port 2 nsew
rlabel metal2 s 41496 47915 41604 47991 4 gnd
port 2 nsew
rlabel metal2 s 41496 31009 41604 31085 4 gnd
port 2 nsew
rlabel metal2 s 41496 46809 41604 46885 4 gnd
port 2 nsew
rlabel metal2 s 41496 29429 41604 29505 4 gnd
port 2 nsew
rlabel metal2 s 41496 40235 41604 40345 4 gnd
port 2 nsew
rlabel metal2 s 41496 47345 41604 47455 4 gnd
port 2 nsew
rlabel metal2 s 41496 36285 41604 36395 4 gnd
port 2 nsew
rlabel metal2 s 41496 42069 41604 42145 4 gnd
port 2 nsew
rlabel metal2 s 41496 27059 41604 27135 4 gnd
port 2 nsew
rlabel metal2 s 41496 44755 41604 44831 4 gnd
port 2 nsew
rlabel metal2 s 41496 37329 41604 37405 4 gnd
port 2 nsew
rlabel metal2 s 41496 40805 41604 40881 4 gnd
port 2 nsew
rlabel metal2 s 41496 35275 41604 35351 4 gnd
port 2 nsew
rlabel metal2 s 41496 33125 41604 33235 4 gnd
port 2 nsew
rlabel metal2 s 0 45449 42684 45497 4 wl_0_113
port 3 nsew
rlabel metal2 s 0 45669 42684 45717 4 wl_1_113
port 4 nsew
rlabel metal2 s 0 46143 42684 46191 4 wl_0_114
port 5 nsew
rlabel metal2 s 0 45923 42684 45971 4 wl_1_114
port 6 nsew
rlabel metal2 s 0 46239 42684 46287 4 wl_0_115
port 7 nsew
rlabel metal2 s 0 46459 42684 46507 4 wl_1_115
port 8 nsew
rlabel metal2 s 0 46933 42684 46981 4 wl_0_116
port 9 nsew
rlabel metal2 s 0 46713 42684 46761 4 wl_1_116
port 10 nsew
rlabel metal2 s 0 47029 42684 47077 4 wl_0_117
port 11 nsew
rlabel metal2 s 0 47249 42684 47297 4 wl_1_117
port 12 nsew
rlabel metal2 s 0 47723 42684 47771 4 wl_0_118
port 13 nsew
rlabel metal2 s 0 47503 42684 47551 4 wl_1_118
port 14 nsew
rlabel metal2 s 0 47819 42684 47867 4 wl_0_119
port 15 nsew
rlabel metal2 s 0 48039 42684 48087 4 wl_1_119
port 16 nsew
rlabel metal2 s 0 48513 42684 48561 4 wl_0_120
port 17 nsew
rlabel metal2 s 0 48293 42684 48341 4 wl_1_120
port 18 nsew
rlabel metal2 s 0 48609 42684 48657 4 wl_0_121
port 19 nsew
rlabel metal2 s 0 48829 42684 48877 4 wl_1_121
port 20 nsew
rlabel metal2 s 0 49303 42684 49351 4 wl_0_122
port 21 nsew
rlabel metal2 s 0 49083 42684 49131 4 wl_1_122
port 22 nsew
rlabel metal2 s 0 49399 42684 49447 4 wl_0_123
port 23 nsew
rlabel metal2 s 0 49619 42684 49667 4 wl_1_123
port 24 nsew
rlabel metal2 s 0 50093 42684 50141 4 wl_0_124
port 25 nsew
rlabel metal2 s 0 49873 42684 49921 4 wl_1_124
port 26 nsew
rlabel metal2 s 0 50189 42684 50237 4 wl_0_125
port 27 nsew
rlabel metal2 s 0 50409 42684 50457 4 wl_1_125
port 28 nsew
rlabel metal2 s 0 50883 42684 50931 4 wl_0_126
port 29 nsew
rlabel metal2 s 0 50663 42684 50711 4 wl_1_126
port 30 nsew
rlabel metal2 s 0 50979 42684 51027 4 wl_0_127
port 31 nsew
rlabel metal2 s 0 51199 42684 51247 4 wl_1_127
port 32 nsew
rlabel metal2 s 0 51453 42684 51501 4 rbl_wl_1_1
port 33 nsew
rlabel metal2 s 0 39033 42684 39081 4 wl_0_96
port 34 nsew
rlabel metal2 s 0 38813 42684 38861 4 wl_1_96
port 35 nsew
rlabel metal2 s 0 39129 42684 39177 4 wl_0_97
port 36 nsew
rlabel metal2 s 0 39349 42684 39397 4 wl_1_97
port 37 nsew
rlabel metal2 s 0 39823 42684 39871 4 wl_0_98
port 38 nsew
rlabel metal2 s 0 39603 42684 39651 4 wl_1_98
port 39 nsew
rlabel metal2 s 0 39919 42684 39967 4 wl_0_99
port 40 nsew
rlabel metal2 s 0 40139 42684 40187 4 wl_1_99
port 41 nsew
rlabel metal2 s 0 40613 42684 40661 4 wl_0_100
port 42 nsew
rlabel metal2 s 0 40393 42684 40441 4 wl_1_100
port 43 nsew
rlabel metal2 s 0 40709 42684 40757 4 wl_0_101
port 44 nsew
rlabel metal2 s 0 40929 42684 40977 4 wl_1_101
port 45 nsew
rlabel metal2 s 0 41403 42684 41451 4 wl_0_102
port 46 nsew
rlabel metal2 s 0 41183 42684 41231 4 wl_1_102
port 47 nsew
rlabel metal2 s 0 41499 42684 41547 4 wl_0_103
port 48 nsew
rlabel metal2 s 0 41719 42684 41767 4 wl_1_103
port 49 nsew
rlabel metal2 s 0 42193 42684 42241 4 wl_0_104
port 50 nsew
rlabel metal2 s 0 41973 42684 42021 4 wl_1_104
port 51 nsew
rlabel metal2 s 0 42289 42684 42337 4 wl_0_105
port 52 nsew
rlabel metal2 s 0 42509 42684 42557 4 wl_1_105
port 53 nsew
rlabel metal2 s 0 42983 42684 43031 4 wl_0_106
port 54 nsew
rlabel metal2 s 0 42763 42684 42811 4 wl_1_106
port 55 nsew
rlabel metal2 s 0 43079 42684 43127 4 wl_0_107
port 56 nsew
rlabel metal2 s 0 43299 42684 43347 4 wl_1_107
port 57 nsew
rlabel metal2 s 0 43773 42684 43821 4 wl_0_108
port 58 nsew
rlabel metal2 s 0 43553 42684 43601 4 wl_1_108
port 59 nsew
rlabel metal2 s 0 43869 42684 43917 4 wl_0_109
port 60 nsew
rlabel metal2 s 0 44089 42684 44137 4 wl_1_109
port 61 nsew
rlabel metal2 s 0 44563 42684 44611 4 wl_0_110
port 62 nsew
rlabel metal2 s 0 44343 42684 44391 4 wl_1_110
port 63 nsew
rlabel metal2 s 0 44659 42684 44707 4 wl_0_111
port 64 nsew
rlabel metal2 s 0 44879 42684 44927 4 wl_1_111
port 65 nsew
rlabel metal2 s 0 45353 42684 45401 4 wl_0_112
port 66 nsew
rlabel metal2 s 0 45133 42684 45181 4 wl_1_112
port 67 nsew
rlabel metal2 s 1080 43395 1188 43505 4 gnd
port 2 nsew
rlabel metal2 s 1080 49969 1188 50045 4 gnd
port 2 nsew
rlabel metal2 s 1080 51075 1188 51151 4 gnd
port 2 nsew
rlabel metal2 s 1080 49495 1188 49571 4 gnd
port 2 nsew
rlabel metal2 s 1080 40015 1188 40091 4 gnd
port 2 nsew
rlabel metal2 s 1080 48135 1188 48245 4 gnd
port 2 nsew
rlabel metal2 s 1080 45765 1188 45875 4 gnd
port 2 nsew
rlabel metal2 s 1080 50759 1188 50835 4 gnd
port 2 nsew
rlabel metal2 s 1080 49715 1188 49825 4 gnd
port 2 nsew
rlabel metal2 s 1080 51295 1188 51405 4 gnd
port 2 nsew
rlabel metal2 s 1080 42069 1188 42145 4 gnd
port 2 nsew
rlabel metal2 s 1080 41025 1188 41135 4 gnd
port 2 nsew
rlabel metal2 s 1080 46809 1188 46885 4 gnd
port 2 nsew
rlabel metal2 s 1080 43965 1188 44041 4 gnd
port 2 nsew
rlabel metal2 s 1080 42385 1188 42461 4 gnd
port 2 nsew
rlabel metal2 s 1080 51549 1188 51625 4 gnd
port 2 nsew
rlabel metal2 s 1080 41595 1188 41671 4 gnd
port 2 nsew
rlabel metal2 s 1080 41279 1188 41355 4 gnd
port 2 nsew
rlabel metal2 s 1080 48705 1188 48781 4 gnd
port 2 nsew
rlabel metal2 s 1080 42859 1188 42935 4 gnd
port 2 nsew
rlabel metal2 s 1080 46555 1188 46665 4 gnd
port 2 nsew
rlabel metal2 s 1080 40489 1188 40565 4 gnd
port 2 nsew
rlabel metal2 s 1080 45229 1188 45305 4 gnd
port 2 nsew
rlabel metal2 s 1080 46335 1188 46411 4 gnd
port 2 nsew
rlabel metal2 s 1080 38909 1188 38985 4 gnd
port 2 nsew
rlabel metal2 s 1080 44975 1188 45085 4 gnd
port 2 nsew
rlabel metal2 s 1080 44439 1188 44515 4 gnd
port 2 nsew
rlabel metal2 s 1080 47915 1188 47991 4 gnd
port 2 nsew
rlabel metal2 s 1080 49179 1188 49255 4 gnd
port 2 nsew
rlabel metal2 s 1080 44185 1188 44295 4 gnd
port 2 nsew
rlabel metal2 s 1080 47599 1188 47675 4 gnd
port 2 nsew
rlabel metal2 s 1080 47125 1188 47201 4 gnd
port 2 nsew
rlabel metal2 s 1080 48925 1188 49035 4 gnd
port 2 nsew
rlabel metal2 s 1080 48389 1188 48465 4 gnd
port 2 nsew
rlabel metal2 s 1080 40235 1188 40345 4 gnd
port 2 nsew
rlabel metal2 s 1080 39445 1188 39555 4 gnd
port 2 nsew
rlabel metal2 s 1080 42605 1188 42715 4 gnd
port 2 nsew
rlabel metal2 s 1080 47345 1188 47455 4 gnd
port 2 nsew
rlabel metal2 s 1080 44755 1188 44831 4 gnd
port 2 nsew
rlabel metal2 s 1080 43649 1188 43725 4 gnd
port 2 nsew
rlabel metal2 s 1080 46019 1188 46095 4 gnd
port 2 nsew
rlabel metal2 s 1080 41815 1188 41925 4 gnd
port 2 nsew
rlabel metal2 s 1080 39699 1188 39775 4 gnd
port 2 nsew
rlabel metal2 s 1080 50285 1188 50361 4 gnd
port 2 nsew
rlabel metal2 s 1080 43175 1188 43251 4 gnd
port 2 nsew
rlabel metal2 s 1080 39225 1188 39301 4 gnd
port 2 nsew
rlabel metal2 s 1080 40805 1188 40881 4 gnd
port 2 nsew
rlabel metal2 s 1080 45545 1188 45621 4 gnd
port 2 nsew
rlabel metal2 s 1080 50505 1188 50615 4 gnd
port 2 nsew
rlabel metal2 s 1080 38119 1188 38195 4 gnd
port 2 nsew
rlabel metal2 s 1080 27059 1188 27135 4 gnd
port 2 nsew
rlabel metal2 s 1080 32335 1188 32445 4 gnd
port 2 nsew
rlabel metal2 s 1080 36539 1188 36615 4 gnd
port 2 nsew
rlabel metal2 s 1080 29965 1188 30075 4 gnd
port 2 nsew
rlabel metal2 s 1080 37865 1188 37975 4 gnd
port 2 nsew
rlabel metal2 s 1080 28639 1188 28715 4 gnd
port 2 nsew
rlabel metal2 s 1080 37329 1188 37405 4 gnd
port 2 nsew
rlabel metal2 s 1080 31325 1188 31401 4 gnd
port 2 nsew
rlabel metal2 s 1080 26805 1188 26915 4 gnd
port 2 nsew
rlabel metal2 s 1080 29175 1188 29285 4 gnd
port 2 nsew
rlabel metal2 s 1080 32115 1188 32191 4 gnd
port 2 nsew
rlabel metal2 s 1080 26269 1188 26345 4 gnd
port 2 nsew
rlabel metal2 s 1080 26585 1188 26661 4 gnd
port 2 nsew
rlabel metal2 s 1080 35275 1188 35351 4 gnd
port 2 nsew
rlabel metal2 s 1080 36285 1188 36395 4 gnd
port 2 nsew
rlabel metal2 s 1080 28385 1188 28495 4 gnd
port 2 nsew
rlabel metal2 s 1080 32589 1188 32665 4 gnd
port 2 nsew
rlabel metal2 s 1080 28165 1188 28241 4 gnd
port 2 nsew
rlabel metal2 s 1080 29745 1188 29821 4 gnd
port 2 nsew
rlabel metal2 s 1080 34485 1188 34561 4 gnd
port 2 nsew
rlabel metal2 s 1080 26015 1188 26125 4 gnd
port 2 nsew
rlabel metal2 s 1080 38435 1188 38511 4 gnd
port 2 nsew
rlabel metal2 s 1080 36065 1188 36141 4 gnd
port 2 nsew
rlabel metal2 s 1080 30755 1188 30865 4 gnd
port 2 nsew
rlabel metal2 s 1080 28955 1188 29031 4 gnd
port 2 nsew
rlabel metal2 s 1080 27849 1188 27925 4 gnd
port 2 nsew
rlabel metal2 s 1080 31009 1188 31085 4 gnd
port 2 nsew
rlabel metal2 s 1080 35749 1188 35825 4 gnd
port 2 nsew
rlabel metal2 s 1080 27595 1188 27705 4 gnd
port 2 nsew
rlabel metal2 s 1080 30535 1188 30611 4 gnd
port 2 nsew
rlabel metal2 s 1080 32905 1188 32981 4 gnd
port 2 nsew
rlabel metal2 s 1080 29429 1188 29505 4 gnd
port 2 nsew
rlabel metal2 s 1080 30219 1188 30295 4 gnd
port 2 nsew
rlabel metal2 s 1080 34705 1188 34815 4 gnd
port 2 nsew
rlabel metal2 s 1080 38655 1188 38765 4 gnd
port 2 nsew
rlabel metal2 s 1080 37075 1188 37185 4 gnd
port 2 nsew
rlabel metal2 s 1080 31799 1188 31875 4 gnd
port 2 nsew
rlabel metal2 s 1080 37645 1188 37721 4 gnd
port 2 nsew
rlabel metal2 s 1080 27375 1188 27451 4 gnd
port 2 nsew
rlabel metal2 s 1080 33379 1188 33455 4 gnd
port 2 nsew
rlabel metal2 s 1080 34959 1188 35035 4 gnd
port 2 nsew
rlabel metal2 s 1080 33125 1188 33235 4 gnd
port 2 nsew
rlabel metal2 s 1080 33695 1188 33771 4 gnd
port 2 nsew
rlabel metal2 s 1080 33915 1188 34025 4 gnd
port 2 nsew
rlabel metal2 s 1080 36855 1188 36931 4 gnd
port 2 nsew
rlabel metal2 s 1080 35495 1188 35605 4 gnd
port 2 nsew
rlabel metal2 s 1080 31545 1188 31655 4 gnd
port 2 nsew
rlabel metal2 s 1080 34169 1188 34245 4 gnd
port 2 nsew
rlabel metal2 s 0 32239 42684 32287 4 wl_1_79
port 68 nsew
rlabel metal2 s 0 32713 42684 32761 4 wl_0_80
port 69 nsew
rlabel metal2 s 0 28859 42684 28907 4 wl_0_71
port 70 nsew
rlabel metal2 s 0 32493 42684 32541 4 wl_1_80
port 71 nsew
rlabel metal2 s 0 29079 42684 29127 4 wl_1_71
port 72 nsew
rlabel metal2 s 0 32809 42684 32857 4 wl_0_81
port 73 nsew
rlabel metal2 s 0 29553 42684 29601 4 wl_0_72
port 74 nsew
rlabel metal2 s 0 27753 42684 27801 4 wl_1_68
port 75 nsew
rlabel metal2 s 0 33029 42684 33077 4 wl_1_81
port 76 nsew
rlabel metal2 s 0 33503 42684 33551 4 wl_0_82
port 77 nsew
rlabel metal2 s 0 33283 42684 33331 4 wl_1_82
port 78 nsew
rlabel metal2 s 0 28069 42684 28117 4 wl_0_69
port 79 nsew
rlabel metal2 s 0 33599 42684 33647 4 wl_0_83
port 80 nsew
rlabel metal2 s 0 33819 42684 33867 4 wl_1_83
port 81 nsew
rlabel metal2 s 0 29333 42684 29381 4 wl_1_72
port 82 nsew
rlabel metal2 s 0 34293 42684 34341 4 wl_0_84
port 83 nsew
rlabel metal2 s 0 34073 42684 34121 4 wl_1_84
port 84 nsew
rlabel metal2 s 0 27279 42684 27327 4 wl_0_67
port 85 nsew
rlabel metal2 s 0 34389 42684 34437 4 wl_0_85
port 86 nsew
rlabel metal2 s 0 34609 42684 34657 4 wl_1_85
port 87 nsew
rlabel metal2 s 0 35083 42684 35131 4 wl_0_86
port 88 nsew
rlabel metal2 s 0 26709 42684 26757 4 wl_1_65
port 89 nsew
rlabel metal2 s 0 34863 42684 34911 4 wl_1_86
port 90 nsew
rlabel metal2 s 0 35179 42684 35227 4 wl_0_87
port 91 nsew
rlabel metal2 s 0 35399 42684 35447 4 wl_1_87
port 92 nsew
rlabel metal2 s 0 26173 42684 26221 4 wl_1_64
port 93 nsew
rlabel metal2 s 0 26393 42684 26441 4 wl_0_64
port 94 nsew
rlabel metal2 s 0 35873 42684 35921 4 wl_0_88
port 95 nsew
rlabel metal2 s 0 35653 42684 35701 4 wl_1_88
port 96 nsew
rlabel metal2 s 0 35969 42684 36017 4 wl_0_89
port 97 nsew
rlabel metal2 s 0 29649 42684 29697 4 wl_0_73
port 98 nsew
rlabel metal2 s 0 29869 42684 29917 4 wl_1_73
port 99 nsew
rlabel metal2 s 0 30343 42684 30391 4 wl_0_74
port 100 nsew
rlabel metal2 s 0 27499 42684 27547 4 wl_1_67
port 101 nsew
rlabel metal2 s 0 36189 42684 36237 4 wl_1_89
port 102 nsew
rlabel metal2 s 0 36663 42684 36711 4 wl_0_90
port 103 nsew
rlabel metal2 s 0 36443 42684 36491 4 wl_1_90
port 104 nsew
rlabel metal2 s 0 36759 42684 36807 4 wl_0_91
port 105 nsew
rlabel metal2 s 0 36979 42684 37027 4 wl_1_91
port 106 nsew
rlabel metal2 s 0 27183 42684 27231 4 wl_0_66
port 107 nsew
rlabel metal2 s 0 30123 42684 30171 4 wl_1_74
port 108 nsew
rlabel metal2 s 0 37453 42684 37501 4 wl_0_92
port 109 nsew
rlabel metal2 s 0 37233 42684 37281 4 wl_1_92
port 110 nsew
rlabel metal2 s 0 37549 42684 37597 4 wl_0_93
port 111 nsew
rlabel metal2 s 0 37769 42684 37817 4 wl_1_93
port 112 nsew
rlabel metal2 s 0 30439 42684 30487 4 wl_0_75
port 113 nsew
rlabel metal2 s 0 30659 42684 30707 4 wl_1_75
port 114 nsew
rlabel metal2 s 0 31133 42684 31181 4 wl_0_76
port 115 nsew
rlabel metal2 s 0 38243 42684 38291 4 wl_0_94
port 116 nsew
rlabel metal2 s 0 30913 42684 30961 4 wl_1_76
port 117 nsew
rlabel metal2 s 0 27973 42684 28021 4 wl_0_68
port 118 nsew
rlabel metal2 s 0 31229 42684 31277 4 wl_0_77
port 119 nsew
rlabel metal2 s 0 38023 42684 38071 4 wl_1_94
port 120 nsew
rlabel metal2 s 0 38339 42684 38387 4 wl_0_95
port 121 nsew
rlabel metal2 s 0 31449 42684 31497 4 wl_1_77
port 122 nsew
rlabel metal2 s 0 38559 42684 38607 4 wl_1_95
port 123 nsew
rlabel metal2 s 0 28289 42684 28337 4 wl_1_69
port 124 nsew
rlabel metal2 s 0 28763 42684 28811 4 wl_0_70
port 125 nsew
rlabel metal2 s 0 26489 42684 26537 4 wl_0_65
port 126 nsew
rlabel metal2 s 0 31923 42684 31971 4 wl_0_78
port 127 nsew
rlabel metal2 s 0 31703 42684 31751 4 wl_1_78
port 128 nsew
rlabel metal2 s 0 28543 42684 28591 4 wl_1_70
port 129 nsew
rlabel metal2 s 0 26963 42684 27011 4 wl_1_66
port 130 nsew
rlabel metal2 s 0 32019 42684 32067 4 wl_0_79
port 131 nsew
rlabel metal2 s 0 13279 42684 13327 4 wl_1_31
port 132 nsew
rlabel metal2 s 0 13753 42684 13801 4 wl_0_32
port 133 nsew
rlabel metal2 s 0 13533 42684 13581 4 wl_1_32
port 134 nsew
rlabel metal2 s 0 13849 42684 13897 4 wl_0_33
port 135 nsew
rlabel metal2 s 0 14069 42684 14117 4 wl_1_33
port 136 nsew
rlabel metal2 s 0 14543 42684 14591 4 wl_0_34
port 137 nsew
rlabel metal2 s 0 14323 42684 14371 4 wl_1_34
port 138 nsew
rlabel metal2 s 0 14639 42684 14687 4 wl_0_35
port 139 nsew
rlabel metal2 s 0 14859 42684 14907 4 wl_1_35
port 140 nsew
rlabel metal2 s 0 15333 42684 15381 4 wl_0_36
port 141 nsew
rlabel metal2 s 0 15113 42684 15161 4 wl_1_36
port 142 nsew
rlabel metal2 s 0 15429 42684 15477 4 wl_0_37
port 143 nsew
rlabel metal2 s 0 15649 42684 15697 4 wl_1_37
port 144 nsew
rlabel metal2 s 0 16123 42684 16171 4 wl_0_38
port 145 nsew
rlabel metal2 s 0 15903 42684 15951 4 wl_1_38
port 146 nsew
rlabel metal2 s 0 16219 42684 16267 4 wl_0_39
port 147 nsew
rlabel metal2 s 0 16439 42684 16487 4 wl_1_39
port 148 nsew
rlabel metal2 s 0 16913 42684 16961 4 wl_0_40
port 149 nsew
rlabel metal2 s 0 16693 42684 16741 4 wl_1_40
port 150 nsew
rlabel metal2 s 0 17009 42684 17057 4 wl_0_41
port 151 nsew
rlabel metal2 s 0 17229 42684 17277 4 wl_1_41
port 152 nsew
rlabel metal2 s 0 17703 42684 17751 4 wl_0_42
port 153 nsew
rlabel metal2 s 0 17483 42684 17531 4 wl_1_42
port 154 nsew
rlabel metal2 s 0 17799 42684 17847 4 wl_0_43
port 155 nsew
rlabel metal2 s 0 18019 42684 18067 4 wl_1_43
port 156 nsew
rlabel metal2 s 0 18493 42684 18541 4 wl_0_44
port 157 nsew
rlabel metal2 s 0 18273 42684 18321 4 wl_1_44
port 158 nsew
rlabel metal2 s 0 18589 42684 18637 4 wl_0_45
port 159 nsew
rlabel metal2 s 0 18809 42684 18857 4 wl_1_45
port 160 nsew
rlabel metal2 s 0 19283 42684 19331 4 wl_0_46
port 161 nsew
rlabel metal2 s 0 19063 42684 19111 4 wl_1_46
port 162 nsew
rlabel metal2 s 0 19379 42684 19427 4 wl_0_47
port 163 nsew
rlabel metal2 s 0 19599 42684 19647 4 wl_1_47
port 164 nsew
rlabel metal2 s 0 20073 42684 20121 4 wl_0_48
port 165 nsew
rlabel metal2 s 0 19853 42684 19901 4 wl_1_48
port 166 nsew
rlabel metal2 s 0 20169 42684 20217 4 wl_0_49
port 167 nsew
rlabel metal2 s 0 20389 42684 20437 4 wl_1_49
port 168 nsew
rlabel metal2 s 0 20863 42684 20911 4 wl_0_50
port 169 nsew
rlabel metal2 s 0 20643 42684 20691 4 wl_1_50
port 170 nsew
rlabel metal2 s 0 20959 42684 21007 4 wl_0_51
port 171 nsew
rlabel metal2 s 0 21179 42684 21227 4 wl_1_51
port 172 nsew
rlabel metal2 s 0 21653 42684 21701 4 wl_0_52
port 173 nsew
rlabel metal2 s 0 21433 42684 21481 4 wl_1_52
port 174 nsew
rlabel metal2 s 0 21749 42684 21797 4 wl_0_53
port 175 nsew
rlabel metal2 s 0 21969 42684 22017 4 wl_1_53
port 176 nsew
rlabel metal2 s 0 22443 42684 22491 4 wl_0_54
port 177 nsew
rlabel metal2 s 0 22223 42684 22271 4 wl_1_54
port 178 nsew
rlabel metal2 s 0 22539 42684 22587 4 wl_0_55
port 179 nsew
rlabel metal2 s 0 22759 42684 22807 4 wl_1_55
port 180 nsew
rlabel metal2 s 0 23233 42684 23281 4 wl_0_56
port 181 nsew
rlabel metal2 s 0 23013 42684 23061 4 wl_1_56
port 182 nsew
rlabel metal2 s 0 23329 42684 23377 4 wl_0_57
port 183 nsew
rlabel metal2 s 0 23549 42684 23597 4 wl_1_57
port 184 nsew
rlabel metal2 s 0 24023 42684 24071 4 wl_0_58
port 185 nsew
rlabel metal2 s 0 23803 42684 23851 4 wl_1_58
port 186 nsew
rlabel metal2 s 0 24119 42684 24167 4 wl_0_59
port 187 nsew
rlabel metal2 s 0 24339 42684 24387 4 wl_1_59
port 188 nsew
rlabel metal2 s 0 24813 42684 24861 4 wl_0_60
port 189 nsew
rlabel metal2 s 0 24593 42684 24641 4 wl_1_60
port 190 nsew
rlabel metal2 s 0 24909 42684 24957 4 wl_0_61
port 191 nsew
rlabel metal2 s 0 25129 42684 25177 4 wl_1_61
port 192 nsew
rlabel metal2 s 0 25603 42684 25651 4 wl_0_62
port 193 nsew
rlabel metal2 s 0 25383 42684 25431 4 wl_1_62
port 194 nsew
rlabel metal2 s 0 25699 42684 25747 4 wl_0_63
port 195 nsew
rlabel metal2 s 0 25919 42684 25967 4 wl_1_63
port 196 nsew
rlabel metal2 s 1080 14419 1188 14495 4 gnd
port 2 nsew
rlabel metal2 s 1080 13945 1188 14021 4 gnd
port 2 nsew
rlabel metal2 s 1080 19695 1188 19805 4 gnd
port 2 nsew
rlabel metal2 s 1080 17895 1188 17971 4 gnd
port 2 nsew
rlabel metal2 s 1080 21055 1188 21131 4 gnd
port 2 nsew
rlabel metal2 s 1080 15525 1188 15601 4 gnd
port 2 nsew
rlabel metal2 s 1080 17325 1188 17435 4 gnd
port 2 nsew
rlabel metal2 s 1080 20265 1188 20341 4 gnd
port 2 nsew
rlabel metal2 s 1080 13375 1188 13485 4 gnd
port 2 nsew
rlabel metal2 s 1080 16789 1188 16865 4 gnd
port 2 nsew
rlabel metal2 s 1080 15209 1188 15285 4 gnd
port 2 nsew
rlabel metal2 s 1080 23109 1188 23185 4 gnd
port 2 nsew
rlabel metal2 s 1080 17105 1188 17181 4 gnd
port 2 nsew
rlabel metal2 s 1080 16315 1188 16391 4 gnd
port 2 nsew
rlabel metal2 s 1080 23645 1188 23755 4 gnd
port 2 nsew
rlabel metal2 s 1080 21845 1188 21921 4 gnd
port 2 nsew
rlabel metal2 s 1080 19159 1188 19235 4 gnd
port 2 nsew
rlabel metal2 s 1080 19475 1188 19551 4 gnd
port 2 nsew
rlabel metal2 s 1080 25479 1188 25555 4 gnd
port 2 nsew
rlabel metal2 s 1080 25005 1188 25081 4 gnd
port 2 nsew
rlabel metal2 s 1080 25795 1188 25871 4 gnd
port 2 nsew
rlabel metal2 s 1080 24215 1188 24291 4 gnd
port 2 nsew
rlabel metal2 s 1080 21529 1188 21605 4 gnd
port 2 nsew
rlabel metal2 s 1080 24435 1188 24545 4 gnd
port 2 nsew
rlabel metal2 s 1080 22065 1188 22175 4 gnd
port 2 nsew
rlabel metal2 s 1080 18115 1188 18225 4 gnd
port 2 nsew
rlabel metal2 s 1080 18369 1188 18445 4 gnd
port 2 nsew
rlabel metal2 s 1080 20739 1188 20815 4 gnd
port 2 nsew
rlabel metal2 s 1080 23899 1188 23975 4 gnd
port 2 nsew
rlabel metal2 s 1080 17579 1188 17655 4 gnd
port 2 nsew
rlabel metal2 s 1080 18685 1188 18761 4 gnd
port 2 nsew
rlabel metal2 s 1080 16535 1188 16645 4 gnd
port 2 nsew
rlabel metal2 s 1080 19949 1188 20025 4 gnd
port 2 nsew
rlabel metal2 s 1080 15999 1188 16075 4 gnd
port 2 nsew
rlabel metal2 s 1080 14955 1188 15065 4 gnd
port 2 nsew
rlabel metal2 s 1080 18905 1188 19015 4 gnd
port 2 nsew
rlabel metal2 s 1080 20485 1188 20595 4 gnd
port 2 nsew
rlabel metal2 s 1080 13629 1188 13705 4 gnd
port 2 nsew
rlabel metal2 s 1080 14165 1188 14275 4 gnd
port 2 nsew
rlabel metal2 s 1080 22855 1188 22965 4 gnd
port 2 nsew
rlabel metal2 s 1080 23425 1188 23501 4 gnd
port 2 nsew
rlabel metal2 s 1080 25225 1188 25335 4 gnd
port 2 nsew
rlabel metal2 s 1080 15745 1188 15855 4 gnd
port 2 nsew
rlabel metal2 s 1080 24689 1188 24765 4 gnd
port 2 nsew
rlabel metal2 s 1080 22635 1188 22711 4 gnd
port 2 nsew
rlabel metal2 s 1080 22319 1188 22395 4 gnd
port 2 nsew
rlabel metal2 s 1080 14735 1188 14811 4 gnd
port 2 nsew
rlabel metal2 s 1080 21275 1188 21385 4 gnd
port 2 nsew
rlabel metal2 s 1080 4939 1188 5015 4 gnd
port 2 nsew
rlabel metal2 s 1080 5255 1188 5331 4 gnd
port 2 nsew
rlabel metal2 s 1080 735 1188 845 4 gnd
port 2 nsew
rlabel metal2 s 1080 11259 1188 11335 4 gnd
port 2 nsew
rlabel metal2 s 1080 12839 1188 12915 4 gnd
port 2 nsew
rlabel metal2 s 1080 2885 1188 2961 4 gnd
port 2 nsew
rlabel metal2 s 1080 5729 1188 5805 4 gnd
port 2 nsew
rlabel metal2 s 1080 11005 1188 11115 4 gnd
port 2 nsew
rlabel metal2 s 1080 6045 1188 6121 4 gnd
port 2 nsew
rlabel metal2 s 1080 3359 1188 3435 4 gnd
port 2 nsew
rlabel metal2 s 1080 7055 1188 7165 4 gnd
port 2 nsew
rlabel metal2 s 1080 3675 1188 3751 4 gnd
port 2 nsew
rlabel metal2 s 1080 4149 1188 4225 4 gnd
port 2 nsew
rlabel metal2 s 1080 3895 1188 4005 4 gnd
port 2 nsew
rlabel metal2 s 1080 515 1188 591 4 gnd
port 2 nsew
rlabel metal2 s 1080 11795 1188 11905 4 gnd
port 2 nsew
rlabel metal2 s 1080 989 1188 1065 4 gnd
port 2 nsew
rlabel metal2 s 1080 13155 1188 13231 4 gnd
port 2 nsew
rlabel metal2 s 1080 6835 1188 6911 4 gnd
port 2 nsew
rlabel metal2 s 1080 9205 1188 9281 4 gnd
port 2 nsew
rlabel metal2 s 1080 7309 1188 7385 4 gnd
port 2 nsew
rlabel metal2 s 1080 4685 1188 4795 4 gnd
port 2 nsew
rlabel metal2 s 1080 9679 1188 9755 4 gnd
port 2 nsew
rlabel metal2 s 1080 1305 1188 1381 4 gnd
port 2 nsew
rlabel metal2 s 1080 2315 1188 2425 4 gnd
port 2 nsew
rlabel metal2 s 1080 5475 1188 5585 4 gnd
port 2 nsew
rlabel metal2 s 1080 7845 1188 7955 4 gnd
port 2 nsew
rlabel metal2 s 1080 2569 1188 2645 4 gnd
port 2 nsew
rlabel metal2 s 1080 3105 1188 3215 4 gnd
port 2 nsew
rlabel metal2 s 1080 12365 1188 12441 4 gnd
port 2 nsew
rlabel metal2 s 1080 8635 1188 8745 4 gnd
port 2 nsew
rlabel metal2 s 1080 10215 1188 10325 4 gnd
port 2 nsew
rlabel metal2 s 1080 9425 1188 9535 4 gnd
port 2 nsew
rlabel metal2 s 1080 1779 1188 1855 4 gnd
port 2 nsew
rlabel metal2 s 1080 4465 1188 4541 4 gnd
port 2 nsew
rlabel metal2 s 1080 11575 1188 11651 4 gnd
port 2 nsew
rlabel metal2 s 1080 7625 1188 7701 4 gnd
port 2 nsew
rlabel metal2 s 1080 8889 1188 8965 4 gnd
port 2 nsew
rlabel metal2 s 1080 12049 1188 12125 4 gnd
port 2 nsew
rlabel metal2 s 1080 9995 1188 10071 4 gnd
port 2 nsew
rlabel metal2 s 1080 10785 1188 10861 4 gnd
port 2 nsew
rlabel metal2 s 1080 10469 1188 10545 4 gnd
port 2 nsew
rlabel metal2 s 1080 8099 1188 8175 4 gnd
port 2 nsew
rlabel metal2 s 1080 12585 1188 12695 4 gnd
port 2 nsew
rlabel metal2 s 1080 2095 1188 2171 4 gnd
port 2 nsew
rlabel metal2 s 1080 8415 1188 8491 4 gnd
port 2 nsew
rlabel metal2 s 1080 1525 1188 1635 4 gnd
port 2 nsew
rlabel metal2 s 1080 6265 1188 6375 4 gnd
port 2 nsew
rlabel metal2 s 1080 6519 1188 6595 4 gnd
port 2 nsew
rlabel metal2 s 0 3799 42684 3847 4 wl_1_7
port 197 nsew
rlabel metal2 s 0 419 42684 467 4 rbl_wl_0_0
port 198 nsew
rlabel metal2 s 0 1113 42684 1161 4 wl_0_0
port 199 nsew
rlabel metal2 s 0 4273 42684 4321 4 wl_0_8
port 200 nsew
rlabel metal2 s 0 4053 42684 4101 4 wl_1_8
port 201 nsew
rlabel metal2 s 0 4369 42684 4417 4 wl_0_9
port 202 nsew
rlabel metal2 s 0 12269 42684 12317 4 wl_0_29
port 203 nsew
rlabel metal2 s 0 893 42684 941 4 wl_1_0
port 204 nsew
rlabel metal2 s 0 1209 42684 1257 4 wl_0_1
port 205 nsew
rlabel metal2 s 0 10593 42684 10641 4 wl_0_24
port 206 nsew
rlabel metal2 s 0 4589 42684 4637 4 wl_1_9
port 207 nsew
rlabel metal2 s 0 10689 42684 10737 4 wl_0_25
port 208 nsew
rlabel metal2 s 0 12489 42684 12537 4 wl_1_29
port 209 nsew
rlabel metal2 s 0 5063 42684 5111 4 wl_0_10
port 210 nsew
rlabel metal2 s 0 1429 42684 1477 4 wl_1_1
port 211 nsew
rlabel metal2 s 0 12963 42684 13011 4 wl_0_30
port 212 nsew
rlabel metal2 s 0 4843 42684 4891 4 wl_1_10
port 213 nsew
rlabel metal2 s 0 5159 42684 5207 4 wl_0_11
port 214 nsew
rlabel metal2 s 0 10119 42684 10167 4 wl_1_23
port 215 nsew
rlabel metal2 s 0 10909 42684 10957 4 wl_1_25
port 216 nsew
rlabel metal2 s 0 1903 42684 1951 4 wl_0_2
port 217 nsew
rlabel metal2 s 0 5379 42684 5427 4 wl_1_11
port 218 nsew
rlabel metal2 s 0 12743 42684 12791 4 wl_1_30
port 219 nsew
rlabel metal2 s 0 1683 42684 1731 4 wl_1_2
port 220 nsew
rlabel metal2 s 0 5853 42684 5901 4 wl_0_12
port 221 nsew
rlabel metal2 s 0 11383 42684 11431 4 wl_0_26
port 222 nsew
rlabel metal2 s 0 13059 42684 13107 4 wl_0_31
port 223 nsew
rlabel metal2 s 0 5633 42684 5681 4 wl_1_12
port 224 nsew
rlabel metal2 s 0 5949 42684 5997 4 wl_0_13
port 225 nsew
rlabel metal2 s 0 11163 42684 11211 4 wl_1_26
port 226 nsew
rlabel metal2 s 0 6169 42684 6217 4 wl_1_13
port 227 nsew
rlabel metal2 s 0 6643 42684 6691 4 wl_0_14
port 228 nsew
rlabel metal2 s 0 6423 42684 6471 4 wl_1_14
port 229 nsew
rlabel metal2 s 0 11479 42684 11527 4 wl_0_27
port 230 nsew
rlabel metal2 s 0 6739 42684 6787 4 wl_0_15
port 231 nsew
rlabel metal2 s 0 10373 42684 10421 4 wl_1_24
port 232 nsew
rlabel metal2 s 0 6959 42684 7007 4 wl_1_15
port 233 nsew
rlabel metal2 s 0 7433 42684 7481 4 wl_0_16
port 234 nsew
rlabel metal2 s 0 7213 42684 7261 4 wl_1_16
port 235 nsew
rlabel metal2 s 0 7529 42684 7577 4 wl_0_17
port 236 nsew
rlabel metal2 s 0 7749 42684 7797 4 wl_1_17
port 237 nsew
rlabel metal2 s 0 8223 42684 8271 4 wl_0_18
port 238 nsew
rlabel metal2 s 0 8003 42684 8051 4 wl_1_18
port 239 nsew
rlabel metal2 s 0 11699 42684 11747 4 wl_1_27
port 240 nsew
rlabel metal2 s 0 8319 42684 8367 4 wl_0_19
port 241 nsew
rlabel metal2 s 0 12173 42684 12221 4 wl_0_28
port 242 nsew
rlabel metal2 s 0 1999 42684 2047 4 wl_0_3
port 243 nsew
rlabel metal2 s 0 2219 42684 2267 4 wl_1_3
port 244 nsew
rlabel metal2 s 0 2693 42684 2741 4 wl_0_4
port 245 nsew
rlabel metal2 s 0 2473 42684 2521 4 wl_1_4
port 246 nsew
rlabel metal2 s 0 2789 42684 2837 4 wl_0_5
port 247 nsew
rlabel metal2 s 0 8539 42684 8587 4 wl_1_19
port 248 nsew
rlabel metal2 s 0 3009 42684 3057 4 wl_1_5
port 249 nsew
rlabel metal2 s 0 9013 42684 9061 4 wl_0_20
port 250 nsew
rlabel metal2 s 0 8793 42684 8841 4 wl_1_20
port 251 nsew
rlabel metal2 s 0 9109 42684 9157 4 wl_0_21
port 252 nsew
rlabel metal2 s 0 11953 42684 12001 4 wl_1_28
port 253 nsew
rlabel metal2 s 0 9329 42684 9377 4 wl_1_21
port 254 nsew
rlabel metal2 s 0 9803 42684 9851 4 wl_0_22
port 255 nsew
rlabel metal2 s 0 9583 42684 9631 4 wl_1_22
port 256 nsew
rlabel metal2 s 0 3483 42684 3531 4 wl_0_6
port 257 nsew
rlabel metal2 s 0 3263 42684 3311 4 wl_1_6
port 258 nsew
rlabel metal2 s 0 9899 42684 9947 4 wl_0_23
port 259 nsew
rlabel metal2 s 0 3579 42684 3627 4 wl_0_7
port 260 nsew
rlabel metal2 s 41496 19475 41604 19551 4 gnd
port 2 nsew
rlabel metal2 s 41496 1525 41604 1635 4 gnd
port 2 nsew
rlabel metal2 s 41496 13375 41604 13485 4 gnd
port 2 nsew
rlabel metal2 s 41496 9205 41604 9281 4 gnd
port 2 nsew
rlabel metal2 s 41496 515 41604 591 4 gnd
port 2 nsew
rlabel metal2 s 41496 13629 41604 13705 4 gnd
port 2 nsew
rlabel metal2 s 41496 10785 41604 10861 4 gnd
port 2 nsew
rlabel metal2 s 41496 20265 41604 20341 4 gnd
port 2 nsew
rlabel metal2 s 41496 5475 41604 5585 4 gnd
port 2 nsew
rlabel metal2 s 41496 22855 41604 22965 4 gnd
port 2 nsew
rlabel metal2 s 41496 735 41604 845 4 gnd
port 2 nsew
rlabel metal2 s 41496 4149 41604 4225 4 gnd
port 2 nsew
rlabel metal2 s 41496 14955 41604 15065 4 gnd
port 2 nsew
rlabel metal2 s 41496 19949 41604 20025 4 gnd
port 2 nsew
rlabel metal2 s 41496 14735 41604 14811 4 gnd
port 2 nsew
rlabel metal2 s 41496 3675 41604 3751 4 gnd
port 2 nsew
rlabel metal2 s 41496 25005 41604 25081 4 gnd
port 2 nsew
rlabel metal2 s 41496 22635 41604 22711 4 gnd
port 2 nsew
rlabel metal2 s 41496 2569 41604 2645 4 gnd
port 2 nsew
rlabel metal2 s 41496 5729 41604 5805 4 gnd
port 2 nsew
rlabel metal2 s 41496 17579 41604 17655 4 gnd
port 2 nsew
rlabel metal2 s 41496 11005 41604 11115 4 gnd
port 2 nsew
rlabel metal2 s 41496 989 41604 1065 4 gnd
port 2 nsew
rlabel metal2 s 41496 2095 41604 2171 4 gnd
port 2 nsew
rlabel metal2 s 41496 11259 41604 11335 4 gnd
port 2 nsew
rlabel metal2 s 41496 8889 41604 8965 4 gnd
port 2 nsew
rlabel metal2 s 41496 6045 41604 6121 4 gnd
port 2 nsew
rlabel metal2 s 41496 15745 41604 15855 4 gnd
port 2 nsew
rlabel metal2 s 41496 23425 41604 23501 4 gnd
port 2 nsew
rlabel metal2 s 41496 3359 41604 3435 4 gnd
port 2 nsew
rlabel metal2 s 41496 3105 41604 3215 4 gnd
port 2 nsew
rlabel metal2 s 41496 5255 41604 5331 4 gnd
port 2 nsew
rlabel metal2 s 41496 12049 41604 12125 4 gnd
port 2 nsew
rlabel metal2 s 41496 1779 41604 1855 4 gnd
port 2 nsew
rlabel metal2 s 41496 7055 41604 7165 4 gnd
port 2 nsew
rlabel metal2 s 41496 4465 41604 4541 4 gnd
port 2 nsew
rlabel metal2 s 41496 3895 41604 4005 4 gnd
port 2 nsew
rlabel metal2 s 41496 12365 41604 12441 4 gnd
port 2 nsew
rlabel metal2 s 41496 12839 41604 12915 4 gnd
port 2 nsew
rlabel metal2 s 41496 11575 41604 11651 4 gnd
port 2 nsew
rlabel metal2 s 41496 21055 41604 21131 4 gnd
port 2 nsew
rlabel metal2 s 41496 4939 41604 5015 4 gnd
port 2 nsew
rlabel metal2 s 41496 10469 41604 10545 4 gnd
port 2 nsew
rlabel metal2 s 41496 6265 41604 6375 4 gnd
port 2 nsew
rlabel metal2 s 41496 15999 41604 16075 4 gnd
port 2 nsew
rlabel metal2 s 41496 21275 41604 21385 4 gnd
port 2 nsew
rlabel metal2 s 41496 18905 41604 19015 4 gnd
port 2 nsew
rlabel metal2 s 41496 24435 41604 24545 4 gnd
port 2 nsew
rlabel metal2 s 41496 23109 41604 23185 4 gnd
port 2 nsew
rlabel metal2 s 41496 1305 41604 1381 4 gnd
port 2 nsew
rlabel metal2 s 41496 2315 41604 2425 4 gnd
port 2 nsew
rlabel metal2 s 41496 18115 41604 18225 4 gnd
port 2 nsew
rlabel metal2 s 41496 21845 41604 21921 4 gnd
port 2 nsew
rlabel metal2 s 41496 16535 41604 16645 4 gnd
port 2 nsew
rlabel metal2 s 41496 25795 41604 25871 4 gnd
port 2 nsew
rlabel metal2 s 41496 2885 41604 2961 4 gnd
port 2 nsew
rlabel metal2 s 41496 14419 41604 14495 4 gnd
port 2 nsew
rlabel metal2 s 41496 22319 41604 22395 4 gnd
port 2 nsew
rlabel metal2 s 41496 18369 41604 18445 4 gnd
port 2 nsew
rlabel metal2 s 41496 15525 41604 15601 4 gnd
port 2 nsew
rlabel metal2 s 41496 13155 41604 13231 4 gnd
port 2 nsew
rlabel metal2 s 41496 8415 41604 8491 4 gnd
port 2 nsew
rlabel metal2 s 41496 20485 41604 20595 4 gnd
port 2 nsew
rlabel metal2 s 41496 25225 41604 25335 4 gnd
port 2 nsew
rlabel metal2 s 41496 9425 41604 9535 4 gnd
port 2 nsew
rlabel metal2 s 41496 4685 41604 4795 4 gnd
port 2 nsew
rlabel metal2 s 41496 21529 41604 21605 4 gnd
port 2 nsew
rlabel metal2 s 41496 15209 41604 15285 4 gnd
port 2 nsew
rlabel metal2 s 41496 7625 41604 7701 4 gnd
port 2 nsew
rlabel metal2 s 41496 7845 41604 7955 4 gnd
port 2 nsew
rlabel metal2 s 41496 9995 41604 10071 4 gnd
port 2 nsew
rlabel metal2 s 41496 24215 41604 24291 4 gnd
port 2 nsew
rlabel metal2 s 41496 24689 41604 24765 4 gnd
port 2 nsew
rlabel metal2 s 41496 17325 41604 17435 4 gnd
port 2 nsew
rlabel metal2 s 41496 8099 41604 8175 4 gnd
port 2 nsew
rlabel metal2 s 41496 8635 41604 8745 4 gnd
port 2 nsew
rlabel metal2 s 41496 6835 41604 6911 4 gnd
port 2 nsew
rlabel metal2 s 41496 11795 41604 11905 4 gnd
port 2 nsew
rlabel metal2 s 41496 25479 41604 25555 4 gnd
port 2 nsew
rlabel metal2 s 41496 20739 41604 20815 4 gnd
port 2 nsew
rlabel metal2 s 41496 9679 41604 9755 4 gnd
port 2 nsew
rlabel metal2 s 41496 7309 41604 7385 4 gnd
port 2 nsew
rlabel metal2 s 41496 16789 41604 16865 4 gnd
port 2 nsew
rlabel metal2 s 41496 22065 41604 22175 4 gnd
port 2 nsew
rlabel metal2 s 41496 19159 41604 19235 4 gnd
port 2 nsew
rlabel metal2 s 41496 6519 41604 6595 4 gnd
port 2 nsew
rlabel metal2 s 41496 23645 41604 23755 4 gnd
port 2 nsew
rlabel metal2 s 41496 14165 41604 14275 4 gnd
port 2 nsew
rlabel metal2 s 41496 12585 41604 12695 4 gnd
port 2 nsew
rlabel metal2 s 41496 17895 41604 17971 4 gnd
port 2 nsew
rlabel metal2 s 41496 19695 41604 19805 4 gnd
port 2 nsew
rlabel metal2 s 41496 13945 41604 14021 4 gnd
port 2 nsew
rlabel metal2 s 41496 16315 41604 16391 4 gnd
port 2 nsew
rlabel metal2 s 41496 17105 41604 17181 4 gnd
port 2 nsew
rlabel metal2 s 41496 10215 41604 10325 4 gnd
port 2 nsew
rlabel metal2 s 41496 18685 41604 18761 4 gnd
port 2 nsew
rlabel metal2 s 41496 23899 41604 23975 4 gnd
port 2 nsew
rlabel metal1 s 41532 41159 41568 41500 4 vdd
port 1 nsew
rlabel metal1 s 41532 40369 41568 40710 4 vdd
port 1 nsew
rlabel metal1 s 41532 37500 41568 37841 4 vdd
port 1 nsew
rlabel metal1 s 41532 32469 41568 32810 4 vdd
port 1 nsew
rlabel metal1 s 41532 36710 41568 37051 4 vdd
port 1 nsew
rlabel metal1 s 41532 47770 41568 48111 4 vdd
port 1 nsew
rlabel metal1 s 41532 45109 41568 45450 4 vdd
port 1 nsew
rlabel metal1 s 41532 30099 41568 30440 4 vdd
port 1 nsew
rlabel metal1 s 41532 50930 41568 51271 4 vdd
port 1 nsew
rlabel metal1 s 41532 43529 41568 43870 4 vdd
port 1 nsew
rlabel metal1 s 41532 50639 41568 50980 4 vdd
port 1 nsew
rlabel metal1 s 41532 42240 41568 42581 4 vdd
port 1 nsew
rlabel metal1 s 41532 32760 41568 33101 4 vdd
port 1 nsew
rlabel metal1 s 41532 28810 41568 29151 4 vdd
port 1 nsew
rlabel metal1 s 41532 41450 41568 41791 4 vdd
port 1 nsew
rlabel metal1 s 41532 48560 41568 48901 4 vdd
port 1 nsew
rlabel metal1 s 41532 38290 41568 38631 4 vdd
port 1 nsew
rlabel metal1 s 41532 45400 41568 45741 4 vdd
port 1 nsew
rlabel metal1 s 41532 49849 41568 50190 4 vdd
port 1 nsew
rlabel metal1 s 41532 29600 41568 29941 4 vdd
port 1 nsew
rlabel metal1 s 41532 35130 41568 35471 4 vdd
port 1 nsew
rlabel metal1 s 41532 26939 41568 27280 4 vdd
port 1 nsew
rlabel metal1 s 41532 46689 41568 47030 4 vdd
port 1 nsew
rlabel metal1 s 41532 40660 41568 41001 4 vdd
port 1 nsew
rlabel metal1 s 41532 36419 41568 36760 4 vdd
port 1 nsew
rlabel metal1 s 41532 39579 41568 39920 4 vdd
port 1 nsew
rlabel metal1 s 41532 43030 41568 43371 4 vdd
port 1 nsew
rlabel metal1 s 41532 33550 41568 33891 4 vdd
port 1 nsew
rlabel metal1 s 41532 51429 41568 51770 4 vdd
port 1 nsew
rlabel metal1 s 41532 47479 41568 47820 4 vdd
port 1 nsew
rlabel metal1 s 41532 26440 41568 26781 4 vdd
port 1 nsew
rlabel metal1 s 41532 48269 41568 48610 4 vdd
port 1 nsew
rlabel metal1 s 41532 33259 41568 33600 4 vdd
port 1 nsew
rlabel metal1 s 41532 39080 41568 39421 4 vdd
port 1 nsew
rlabel metal1 s 41532 28020 41568 28361 4 vdd
port 1 nsew
rlabel metal1 s 41532 39870 41568 40211 4 vdd
port 1 nsew
rlabel metal1 s 41532 34340 41568 34681 4 vdd
port 1 nsew
rlabel metal1 s 41532 50140 41568 50481 4 vdd
port 1 nsew
rlabel metal1 s 41532 49350 41568 49691 4 vdd
port 1 nsew
rlabel metal1 s 41532 43820 41568 44161 4 vdd
port 1 nsew
rlabel metal1 s 41532 41949 41568 42290 4 vdd
port 1 nsew
rlabel metal1 s 41532 46980 41568 47321 4 vdd
port 1 nsew
rlabel metal1 s 41532 30889 41568 31230 4 vdd
port 1 nsew
rlabel metal1 s 41532 29309 41568 29650 4 vdd
port 1 nsew
rlabel metal1 s 41532 37209 41568 37550 4 vdd
port 1 nsew
rlabel metal1 s 41532 49059 41568 49400 4 vdd
port 1 nsew
rlabel metal1 s 41532 27230 41568 27571 4 vdd
port 1 nsew
rlabel metal1 s 41532 28519 41568 28860 4 vdd
port 1 nsew
rlabel metal1 s 41532 34049 41568 34390 4 vdd
port 1 nsew
rlabel metal1 s 41532 46190 41568 46531 4 vdd
port 1 nsew
rlabel metal1 s 41532 30390 41568 30731 4 vdd
port 1 nsew
rlabel metal1 s 41532 34839 41568 35180 4 vdd
port 1 nsew
rlabel metal1 s 41532 42739 41568 43080 4 vdd
port 1 nsew
rlabel metal1 s 41532 37999 41568 38340 4 vdd
port 1 nsew
rlabel metal1 s 41532 38789 41568 39130 4 vdd
port 1 nsew
rlabel metal1 s 41532 44319 41568 44660 4 vdd
port 1 nsew
rlabel metal1 s 41532 44610 41568 44951 4 vdd
port 1 nsew
rlabel metal1 s 41532 27729 41568 28070 4 vdd
port 1 nsew
rlabel metal1 s 41532 31180 41568 31521 4 vdd
port 1 nsew
rlabel metal1 s 41532 35629 41568 35970 4 vdd
port 1 nsew
rlabel metal1 s 41532 35920 41568 36261 4 vdd
port 1 nsew
rlabel metal1 s 41532 31970 41568 32311 4 vdd
port 1 nsew
rlabel metal1 s 41532 31679 41568 32020 4 vdd
port 1 nsew
rlabel metal1 s 41532 45899 41568 46240 4 vdd
port 1 nsew
rlabel metal1 s 41532 26149 41568 26490 4 vdd
port 1 nsew
rlabel metal1 s 1116 38290 1152 38631 4 vdd
port 1 nsew
rlabel metal1 s 1116 39579 1152 39920 4 vdd
port 1 nsew
rlabel metal1 s 1116 41450 1152 41791 4 vdd
port 1 nsew
rlabel metal1 s 1116 50140 1152 50481 4 vdd
port 1 nsew
rlabel metal1 s 1116 45400 1152 45741 4 vdd
port 1 nsew
rlabel metal1 s 1116 26440 1152 26781 4 vdd
port 1 nsew
rlabel metal1 s 1116 50639 1152 50980 4 vdd
port 1 nsew
rlabel metal1 s 1116 34340 1152 34681 4 vdd
port 1 nsew
rlabel metal1 s 1116 44319 1152 44660 4 vdd
port 1 nsew
rlabel metal1 s 1116 33550 1152 33891 4 vdd
port 1 nsew
rlabel metal1 s 1116 31970 1152 32311 4 vdd
port 1 nsew
rlabel metal1 s 1116 48560 1152 48901 4 vdd
port 1 nsew
rlabel metal1 s 1116 37209 1152 37550 4 vdd
port 1 nsew
rlabel metal1 s 1116 45109 1152 45450 4 vdd
port 1 nsew
rlabel metal1 s 1116 33259 1152 33600 4 vdd
port 1 nsew
rlabel metal1 s 1116 47770 1152 48111 4 vdd
port 1 nsew
rlabel metal1 s 1116 43820 1152 44161 4 vdd
port 1 nsew
rlabel metal1 s 1116 42739 1152 43080 4 vdd
port 1 nsew
rlabel metal1 s 1116 30390 1152 30731 4 vdd
port 1 nsew
rlabel metal1 s 1116 35920 1152 36261 4 vdd
port 1 nsew
rlabel metal1 s 1116 36710 1152 37051 4 vdd
port 1 nsew
rlabel metal1 s 1116 49059 1152 49400 4 vdd
port 1 nsew
rlabel metal1 s 1116 35130 1152 35471 4 vdd
port 1 nsew
rlabel metal1 s 1116 48269 1152 48610 4 vdd
port 1 nsew
rlabel metal1 s 1116 47479 1152 47820 4 vdd
port 1 nsew
rlabel metal1 s 1116 27230 1152 27571 4 vdd
port 1 nsew
rlabel metal1 s 1116 49350 1152 49691 4 vdd
port 1 nsew
rlabel metal1 s 1116 40660 1152 41001 4 vdd
port 1 nsew
rlabel metal1 s 1116 28519 1152 28860 4 vdd
port 1 nsew
rlabel metal1 s 1116 28020 1152 28361 4 vdd
port 1 nsew
rlabel metal1 s 1116 31679 1152 32020 4 vdd
port 1 nsew
rlabel metal1 s 1116 46190 1152 46531 4 vdd
port 1 nsew
rlabel metal1 s 1116 38789 1152 39130 4 vdd
port 1 nsew
rlabel metal1 s 1116 26149 1152 26490 4 vdd
port 1 nsew
rlabel metal1 s 1116 36419 1152 36760 4 vdd
port 1 nsew
rlabel metal1 s 1116 30889 1152 31230 4 vdd
port 1 nsew
rlabel metal1 s 1116 30099 1152 30440 4 vdd
port 1 nsew
rlabel metal1 s 1116 27729 1152 28070 4 vdd
port 1 nsew
rlabel metal1 s 1116 43030 1152 43371 4 vdd
port 1 nsew
rlabel metal1 s 1116 32760 1152 33101 4 vdd
port 1 nsew
rlabel metal1 s 1116 49849 1152 50190 4 vdd
port 1 nsew
rlabel metal1 s 1116 42240 1152 42581 4 vdd
port 1 nsew
rlabel metal1 s 1116 37500 1152 37841 4 vdd
port 1 nsew
rlabel metal1 s 1116 34839 1152 35180 4 vdd
port 1 nsew
rlabel metal1 s 1116 41949 1152 42290 4 vdd
port 1 nsew
rlabel metal1 s 1116 45899 1152 46240 4 vdd
port 1 nsew
rlabel metal1 s 1116 41159 1152 41500 4 vdd
port 1 nsew
rlabel metal1 s 1116 39080 1152 39421 4 vdd
port 1 nsew
rlabel metal1 s 1116 26939 1152 27280 4 vdd
port 1 nsew
rlabel metal1 s 1116 29600 1152 29941 4 vdd
port 1 nsew
rlabel metal1 s 1116 31180 1152 31521 4 vdd
port 1 nsew
rlabel metal1 s 1116 51429 1152 51770 4 vdd
port 1 nsew
rlabel metal1 s 1116 50930 1152 51271 4 vdd
port 1 nsew
rlabel metal1 s 1116 35629 1152 35970 4 vdd
port 1 nsew
rlabel metal1 s 1116 40369 1152 40710 4 vdd
port 1 nsew
rlabel metal1 s 1116 44610 1152 44951 4 vdd
port 1 nsew
rlabel metal1 s 1116 39870 1152 40211 4 vdd
port 1 nsew
rlabel metal1 s 1116 43529 1152 43870 4 vdd
port 1 nsew
rlabel metal1 s 1116 34049 1152 34390 4 vdd
port 1 nsew
rlabel metal1 s 1116 46689 1152 47030 4 vdd
port 1 nsew
rlabel metal1 s 1116 37999 1152 38340 4 vdd
port 1 nsew
rlabel metal1 s 1116 29309 1152 29650 4 vdd
port 1 nsew
rlabel metal1 s 1116 32469 1152 32810 4 vdd
port 1 nsew
rlabel metal1 s 1116 28810 1152 29151 4 vdd
port 1 nsew
rlabel metal1 s 1116 46980 1152 47321 4 vdd
port 1 nsew
rlabel metal1 s 11244 0 11280 52140 4 bl_0_15
port 261 nsew
rlabel metal1 s 11172 0 11208 52140 4 br_0_15
port 262 nsew
rlabel metal1 s 11436 0 11472 52140 4 bl_0_16
port 263 nsew
rlabel metal1 s 11652 0 11688 52140 4 bl_1_16
port 264 nsew
rlabel metal1 s 11508 0 11544 52140 4 br_0_16
port 265 nsew
rlabel metal1 s 11724 0 11760 52140 4 br_1_16
port 266 nsew
rlabel metal1 s 12492 0 12528 52140 4 bl_0_17
port 267 nsew
rlabel metal1 s 12276 0 12312 52140 4 bl_1_17
port 268 nsew
rlabel metal1 s 12420 0 12456 52140 4 br_0_17
port 269 nsew
rlabel metal1 s 12204 0 12240 52140 4 br_1_17
port 270 nsew
rlabel metal1 s 12684 0 12720 52140 4 bl_0_18
port 271 nsew
rlabel metal1 s 12900 0 12936 52140 4 bl_1_18
port 272 nsew
rlabel metal1 s 12756 0 12792 52140 4 br_0_18
port 273 nsew
rlabel metal1 s 12972 0 13008 52140 4 br_1_18
port 274 nsew
rlabel metal1 s 13740 0 13776 52140 4 bl_0_19
port 275 nsew
rlabel metal1 s 13524 0 13560 52140 4 bl_1_19
port 276 nsew
rlabel metal1 s 13668 0 13704 52140 4 br_0_19
port 277 nsew
rlabel metal1 s 13452 0 13488 52140 4 br_1_19
port 278 nsew
rlabel metal1 s 13932 0 13968 52140 4 bl_0_20
port 279 nsew
rlabel metal1 s 14148 0 14184 52140 4 bl_1_20
port 280 nsew
rlabel metal1 s 14004 0 14040 52140 4 br_0_20
port 281 nsew
rlabel metal1 s 14220 0 14256 52140 4 br_1_20
port 282 nsew
rlabel metal1 s 14988 0 15024 52140 4 bl_0_21
port 283 nsew
rlabel metal1 s 14772 0 14808 52140 4 bl_1_21
port 284 nsew
rlabel metal1 s 14916 0 14952 52140 4 br_0_21
port 285 nsew
rlabel metal1 s 14700 0 14736 52140 4 br_1_21
port 286 nsew
rlabel metal1 s 15180 0 15216 52140 4 bl_0_22
port 287 nsew
rlabel metal1 s 15396 0 15432 52140 4 bl_1_22
port 288 nsew
rlabel metal1 s 15252 0 15288 52140 4 br_0_22
port 289 nsew
rlabel metal1 s 15468 0 15504 52140 4 br_1_22
port 290 nsew
rlabel metal1 s 16236 0 16272 52140 4 bl_0_23
port 291 nsew
rlabel metal1 s 16020 0 16056 52140 4 bl_1_23
port 292 nsew
rlabel metal1 s 16164 0 16200 52140 4 br_0_23
port 293 nsew
rlabel metal1 s 15948 0 15984 52140 4 br_1_23
port 294 nsew
rlabel metal1 s 16428 0 16464 52140 4 bl_0_24
port 295 nsew
rlabel metal1 s 16644 0 16680 52140 4 bl_1_24
port 296 nsew
rlabel metal1 s 16500 0 16536 52140 4 br_0_24
port 297 nsew
rlabel metal1 s 16716 0 16752 52140 4 br_1_24
port 298 nsew
rlabel metal1 s 17484 0 17520 52140 4 bl_0_25
port 299 nsew
rlabel metal1 s 17268 0 17304 52140 4 bl_1_25
port 300 nsew
rlabel metal1 s 17412 0 17448 52140 4 br_0_25
port 301 nsew
rlabel metal1 s 17196 0 17232 52140 4 br_1_25
port 302 nsew
rlabel metal1 s 17676 0 17712 52140 4 bl_0_26
port 303 nsew
rlabel metal1 s 17892 0 17928 52140 4 bl_1_26
port 304 nsew
rlabel metal1 s 17748 0 17784 52140 4 br_0_26
port 305 nsew
rlabel metal1 s 17964 0 18000 52140 4 br_1_26
port 306 nsew
rlabel metal1 s 18732 0 18768 52140 4 bl_0_27
port 307 nsew
rlabel metal1 s 18516 0 18552 52140 4 bl_1_27
port 308 nsew
rlabel metal1 s 18660 0 18696 52140 4 br_0_27
port 309 nsew
rlabel metal1 s 18444 0 18480 52140 4 br_1_27
port 310 nsew
rlabel metal1 s 18924 0 18960 52140 4 bl_0_28
port 311 nsew
rlabel metal1 s 19140 0 19176 52140 4 bl_1_28
port 312 nsew
rlabel metal1 s 18996 0 19032 52140 4 br_0_28
port 313 nsew
rlabel metal1 s 19212 0 19248 52140 4 br_1_28
port 314 nsew
rlabel metal1 s 19980 0 20016 52140 4 bl_0_29
port 315 nsew
rlabel metal1 s 19764 0 19800 52140 4 bl_1_29
port 316 nsew
rlabel metal1 s 19908 0 19944 52140 4 br_0_29
port 317 nsew
rlabel metal1 s 19692 0 19728 52140 4 br_1_29
port 318 nsew
rlabel metal1 s 20172 0 20208 52140 4 bl_0_30
port 319 nsew
rlabel metal1 s 20388 0 20424 52140 4 bl_1_30
port 320 nsew
rlabel metal1 s 20244 0 20280 52140 4 br_0_30
port 321 nsew
rlabel metal1 s 20460 0 20496 52140 4 br_1_30
port 322 nsew
rlabel metal1 s 21228 0 21264 52140 4 bl_0_31
port 323 nsew
rlabel metal1 s 21012 0 21048 52140 4 bl_1_31
port 324 nsew
rlabel metal1 s 21156 0 21192 52140 4 br_0_31
port 325 nsew
rlabel metal1 s 20940 0 20976 52140 4 br_1_31
port 326 nsew
rlabel metal1 s 9156 0 9192 52140 4 bl_1_12
port 327 nsew
rlabel metal1 s 9012 0 9048 52140 4 br_0_12
port 328 nsew
rlabel metal1 s 9228 0 9264 52140 4 br_1_12
port 329 nsew
rlabel metal1 s 9996 0 10032 52140 4 bl_0_13
port 330 nsew
rlabel metal1 s 9780 0 9816 52140 4 bl_1_13
port 331 nsew
rlabel metal1 s 9924 0 9960 52140 4 br_0_13
port 332 nsew
rlabel metal1 s 9708 0 9744 52140 4 br_1_13
port 333 nsew
rlabel metal1 s 10188 0 10224 52140 4 bl_0_14
port 334 nsew
rlabel metal1 s 10404 0 10440 52140 4 bl_1_14
port 335 nsew
rlabel metal1 s 10260 0 10296 52140 4 br_0_14
port 336 nsew
rlabel metal1 s 10476 0 10512 52140 4 br_1_14
port 337 nsew
rlabel metal1 s 1188 0 1224 52140 4 rbl_br_0_0
port 338 nsew
rlabel metal1 s 11028 0 11064 52140 4 bl_1_15
port 339 nsew
rlabel metal1 s 972 0 1008 52140 4 rbl_br_1_0
port 340 nsew
rlabel metal1 s 10956 0 10992 52140 4 br_1_15
port 341 nsew
rlabel metal1 s 1116 22989 1152 23330 4 vdd
port 1 nsew
rlabel metal1 s 1116 19829 1152 20170 4 vdd
port 1 nsew
rlabel metal1 s 1452 0 1488 52140 4 bl_0_0
port 342 nsew
rlabel metal1 s 1668 0 1704 52140 4 bl_1_0
port 343 nsew
rlabel metal1 s 1524 0 1560 52140 4 br_0_0
port 344 nsew
rlabel metal1 s 1740 0 1776 52140 4 br_1_0
port 345 nsew
rlabel metal1 s 2508 0 2544 52140 4 bl_0_1
port 346 nsew
rlabel metal1 s 2292 0 2328 52140 4 bl_1_1
port 347 nsew
rlabel metal1 s 2436 0 2472 52140 4 br_0_1
port 348 nsew
rlabel metal1 s 2220 0 2256 52140 4 br_1_1
port 349 nsew
rlabel metal1 s 2700 0 2736 52140 4 bl_0_2
port 350 nsew
rlabel metal1 s 2916 0 2952 52140 4 bl_1_2
port 351 nsew
rlabel metal1 s 1116 24860 1152 25201 4 vdd
port 1 nsew
rlabel metal1 s 1116 15879 1152 16220 4 vdd
port 1 nsew
rlabel metal1 s 1116 25650 1152 25991 4 vdd
port 1 nsew
rlabel metal1 s 1116 20120 1152 20461 4 vdd
port 1 nsew
rlabel metal1 s 2772 0 2808 52140 4 br_0_2
port 352 nsew
rlabel metal1 s 2988 0 3024 52140 4 br_1_2
port 353 nsew
rlabel metal1 s 3756 0 3792 52140 4 bl_0_3
port 354 nsew
rlabel metal1 s 3540 0 3576 52140 4 bl_1_3
port 355 nsew
rlabel metal1 s 1116 24569 1152 24910 4 vdd
port 1 nsew
rlabel metal1 s 1116 18249 1152 18590 4 vdd
port 1 nsew
rlabel metal1 s 3684 0 3720 52140 4 br_0_3
port 356 nsew
rlabel metal1 s 3468 0 3504 52140 4 br_1_3
port 357 nsew
rlabel metal1 s 1116 14299 1152 14640 4 vdd
port 1 nsew
rlabel metal1 s 3948 0 3984 52140 4 bl_0_4
port 358 nsew
rlabel metal1 s 4164 0 4200 52140 4 bl_1_4
port 359 nsew
rlabel metal1 s 4020 0 4056 52140 4 br_0_4
port 360 nsew
rlabel metal1 s 4236 0 4272 52140 4 br_1_4
port 361 nsew
rlabel metal1 s 5004 0 5040 52140 4 bl_0_5
port 362 nsew
rlabel metal1 s 1116 17750 1152 18091 4 vdd
port 1 nsew
rlabel metal1 s 4788 0 4824 52140 4 bl_1_5
port 363 nsew
rlabel metal1 s 4932 0 4968 52140 4 br_0_5
port 364 nsew
rlabel metal1 s 4716 0 4752 52140 4 br_1_5
port 365 nsew
rlabel metal1 s 5196 0 5232 52140 4 bl_0_6
port 366 nsew
rlabel metal1 s 1116 21700 1152 22041 4 vdd
port 1 nsew
rlabel metal1 s 1116 20619 1152 20960 4 vdd
port 1 nsew
rlabel metal1 s 1116 17459 1152 17800 4 vdd
port 1 nsew
rlabel metal1 s 5412 0 5448 52140 4 bl_1_6
port 367 nsew
rlabel metal1 s 1116 23280 1152 23621 4 vdd
port 1 nsew
rlabel metal1 s 5268 0 5304 52140 4 br_0_6
port 368 nsew
rlabel metal1 s 1116 15089 1152 15430 4 vdd
port 1 nsew
rlabel metal1 s 1116 13509 1152 13850 4 vdd
port 1 nsew
rlabel metal1 s 1116 23779 1152 24120 4 vdd
port 1 nsew
rlabel metal1 s 5484 0 5520 52140 4 br_1_6
port 369 nsew
rlabel metal1 s 1116 13800 1152 14141 4 vdd
port 1 nsew
rlabel metal1 s 6252 0 6288 52140 4 bl_0_7
port 370 nsew
rlabel metal1 s 6036 0 6072 52140 4 bl_1_7
port 371 nsew
rlabel metal1 s 1116 25359 1152 25700 4 vdd
port 1 nsew
rlabel metal1 s 6180 0 6216 52140 4 br_0_7
port 372 nsew
rlabel metal1 s 1116 21409 1152 21750 4 vdd
port 1 nsew
rlabel metal1 s 5964 0 6000 52140 4 br_1_7
port 373 nsew
rlabel metal1 s 6444 0 6480 52140 4 bl_0_8
port 374 nsew
rlabel metal1 s 6660 0 6696 52140 4 bl_1_8
port 375 nsew
rlabel metal1 s 6516 0 6552 52140 4 br_0_8
port 376 nsew
rlabel metal1 s 1116 15380 1152 15721 4 vdd
port 1 nsew
rlabel metal1 s 1116 18540 1152 18881 4 vdd
port 1 nsew
rlabel metal1 s 6732 0 6768 52140 4 br_1_8
port 377 nsew
rlabel metal1 s 7500 0 7536 52140 4 bl_0_9
port 378 nsew
rlabel metal1 s 7284 0 7320 52140 4 bl_1_9
port 379 nsew
rlabel metal1 s 7428 0 7464 52140 4 br_0_9
port 380 nsew
rlabel metal1 s 1116 16170 1152 16511 4 vdd
port 1 nsew
rlabel metal1 s 1116 22490 1152 22831 4 vdd
port 1 nsew
rlabel metal1 s 1116 20910 1152 21251 4 vdd
port 1 nsew
rlabel metal1 s 7212 0 7248 52140 4 br_1_9
port 381 nsew
rlabel metal1 s 7692 0 7728 52140 4 bl_0_10
port 382 nsew
rlabel metal1 s 1116 24070 1152 24411 4 vdd
port 1 nsew
rlabel metal1 s 1116 19330 1152 19671 4 vdd
port 1 nsew
rlabel metal1 s 7908 0 7944 52140 4 bl_1_10
port 383 nsew
rlabel metal1 s 7764 0 7800 52140 4 br_0_10
port 384 nsew
rlabel metal1 s 1116 16669 1152 17010 4 vdd
port 1 nsew
rlabel metal1 s 7980 0 8016 52140 4 br_1_10
port 385 nsew
rlabel metal1 s 8748 0 8784 52140 4 bl_0_11
port 386 nsew
rlabel metal1 s 1116 16960 1152 17301 4 vdd
port 1 nsew
rlabel metal1 s 8532 0 8568 52140 4 bl_1_11
port 387 nsew
rlabel metal1 s 1116 22199 1152 22540 4 vdd
port 1 nsew
rlabel metal1 s 1116 14590 1152 14931 4 vdd
port 1 nsew
rlabel metal1 s 1116 19039 1152 19380 4 vdd
port 1 nsew
rlabel metal1 s 8676 0 8712 52140 4 br_0_11
port 388 nsew
rlabel metal1 s 8460 0 8496 52140 4 br_1_11
port 389 nsew
rlabel metal1 s 8940 0 8976 52140 4 bl_0_12
port 390 nsew
rlabel metal1 s 1260 0 1296 52140 4 rbl_bl_0_0
port 391 nsew
rlabel metal1 s 1044 0 1080 52140 4 rbl_bl_1_0
port 392 nsew
rlabel metal1 s 1116 370 1152 711 4 vdd
port 1 nsew
rlabel metal1 s 1116 12719 1152 13060 4 vdd
port 1 nsew
rlabel metal1 s 1116 7189 1152 7530 4 vdd
port 1 nsew
rlabel metal1 s 1116 2449 1152 2790 4 vdd
port 1 nsew
rlabel metal1 s 1116 9850 1152 10191 4 vdd
port 1 nsew
rlabel metal1 s 1116 7979 1152 8320 4 vdd
port 1 nsew
rlabel metal1 s 1116 13010 1152 13351 4 vdd
port 1 nsew
rlabel metal1 s 1116 7480 1152 7821 4 vdd
port 1 nsew
rlabel metal1 s 1116 8270 1152 8611 4 vdd
port 1 nsew
rlabel metal1 s 1116 1160 1152 1501 4 vdd
port 1 nsew
rlabel metal1 s 1116 4819 1152 5160 4 vdd
port 1 nsew
rlabel metal1 s 1116 6690 1152 7031 4 vdd
port 1 nsew
rlabel metal1 s 1116 11929 1152 12270 4 vdd
port 1 nsew
rlabel metal1 s 1116 4320 1152 4661 4 vdd
port 1 nsew
rlabel metal1 s 1116 2740 1152 3081 4 vdd
port 1 nsew
rlabel metal1 s 1116 3239 1152 3580 4 vdd
port 1 nsew
rlabel metal1 s 1116 10349 1152 10690 4 vdd
port 1 nsew
rlabel metal1 s 1116 1659 1152 2000 4 vdd
port 1 nsew
rlabel metal1 s 1116 869 1152 1210 4 vdd
port 1 nsew
rlabel metal1 s 1116 6399 1152 6740 4 vdd
port 1 nsew
rlabel metal1 s 1116 10640 1152 10981 4 vdd
port 1 nsew
rlabel metal1 s 1116 4029 1152 4370 4 vdd
port 1 nsew
rlabel metal1 s 1116 1950 1152 2291 4 vdd
port 1 nsew
rlabel metal1 s 1116 11430 1152 11771 4 vdd
port 1 nsew
rlabel metal1 s 1116 12220 1152 12561 4 vdd
port 1 nsew
rlabel metal1 s 1116 5110 1152 5451 4 vdd
port 1 nsew
rlabel metal1 s 1116 3530 1152 3871 4 vdd
port 1 nsew
rlabel metal1 s 1116 5900 1152 6241 4 vdd
port 1 nsew
rlabel metal1 s 1116 8769 1152 9110 4 vdd
port 1 nsew
rlabel metal1 s 1116 9559 1152 9900 4 vdd
port 1 nsew
rlabel metal1 s 1116 11139 1152 11480 4 vdd
port 1 nsew
rlabel metal1 s 1116 9060 1152 9401 4 vdd
port 1 nsew
rlabel metal1 s 1116 5609 1152 5950 4 vdd
port 1 nsew
rlabel metal1 s 41532 16960 41568 17301 4 vdd
port 1 nsew
rlabel metal1 s 41532 24070 41568 24411 4 vdd
port 1 nsew
rlabel metal1 s 41532 20910 41568 21251 4 vdd
port 1 nsew
rlabel metal1 s 41532 19330 41568 19671 4 vdd
port 1 nsew
rlabel metal1 s 31620 0 31656 52140 4 bl_1_48
port 393 nsew
rlabel metal1 s 41532 21409 41568 21750 4 vdd
port 1 nsew
rlabel metal1 s 31692 0 31728 52140 4 br_1_48
port 394 nsew
rlabel metal1 s 32460 0 32496 52140 4 bl_0_49
port 395 nsew
rlabel metal1 s 32244 0 32280 52140 4 bl_1_49
port 396 nsew
rlabel metal1 s 32388 0 32424 52140 4 br_0_49
port 397 nsew
rlabel metal1 s 32172 0 32208 52140 4 br_1_49
port 398 nsew
rlabel metal1 s 32652 0 32688 52140 4 bl_0_50
port 399 nsew
rlabel metal1 s 32868 0 32904 52140 4 bl_1_50
port 400 nsew
rlabel metal1 s 32724 0 32760 52140 4 br_0_50
port 401 nsew
rlabel metal1 s 32940 0 32976 52140 4 br_1_50
port 402 nsew
rlabel metal1 s 33708 0 33744 52140 4 bl_0_51
port 403 nsew
rlabel metal1 s 33492 0 33528 52140 4 bl_1_51
port 404 nsew
rlabel metal1 s 33636 0 33672 52140 4 br_0_51
port 405 nsew
rlabel metal1 s 33420 0 33456 52140 4 br_1_51
port 406 nsew
rlabel metal1 s 33900 0 33936 52140 4 bl_0_52
port 407 nsew
rlabel metal1 s 34116 0 34152 52140 4 bl_1_52
port 408 nsew
rlabel metal1 s 33972 0 34008 52140 4 br_0_52
port 409 nsew
rlabel metal1 s 34188 0 34224 52140 4 br_1_52
port 410 nsew
rlabel metal1 s 34956 0 34992 52140 4 bl_0_53
port 411 nsew
rlabel metal1 s 34740 0 34776 52140 4 bl_1_53
port 412 nsew
rlabel metal1 s 41532 18249 41568 18590 4 vdd
port 1 nsew
rlabel metal1 s 34884 0 34920 52140 4 br_0_53
port 413 nsew
rlabel metal1 s 34668 0 34704 52140 4 br_1_53
port 414 nsew
rlabel metal1 s 35148 0 35184 52140 4 bl_0_54
port 415 nsew
rlabel metal1 s 35364 0 35400 52140 4 bl_1_54
port 416 nsew
rlabel metal1 s 35220 0 35256 52140 4 br_0_54
port 417 nsew
rlabel metal1 s 35436 0 35472 52140 4 br_1_54
port 418 nsew
rlabel metal1 s 41532 21700 41568 22041 4 vdd
port 1 nsew
rlabel metal1 s 36204 0 36240 52140 4 bl_0_55
port 419 nsew
rlabel metal1 s 35988 0 36024 52140 4 bl_1_55
port 420 nsew
rlabel metal1 s 36132 0 36168 52140 4 br_0_55
port 421 nsew
rlabel metal1 s 35916 0 35952 52140 4 br_1_55
port 422 nsew
rlabel metal1 s 36396 0 36432 52140 4 bl_0_56
port 423 nsew
rlabel metal1 s 41532 22490 41568 22831 4 vdd
port 1 nsew
rlabel metal1 s 36612 0 36648 52140 4 bl_1_56
port 424 nsew
rlabel metal1 s 36468 0 36504 52140 4 br_0_56
port 425 nsew
rlabel metal1 s 41532 15879 41568 16220 4 vdd
port 1 nsew
rlabel metal1 s 41532 25650 41568 25991 4 vdd
port 1 nsew
rlabel metal1 s 36684 0 36720 52140 4 br_1_56
port 426 nsew
rlabel metal1 s 37452 0 37488 52140 4 bl_0_57
port 427 nsew
rlabel metal1 s 37236 0 37272 52140 4 bl_1_57
port 428 nsew
rlabel metal1 s 37380 0 37416 52140 4 br_0_57
port 429 nsew
rlabel metal1 s 41532 22199 41568 22540 4 vdd
port 1 nsew
rlabel metal1 s 41532 24569 41568 24910 4 vdd
port 1 nsew
rlabel metal1 s 37164 0 37200 52140 4 br_1_57
port 430 nsew
rlabel metal1 s 37644 0 37680 52140 4 bl_0_58
port 431 nsew
rlabel metal1 s 37860 0 37896 52140 4 bl_1_58
port 432 nsew
rlabel metal1 s 37716 0 37752 52140 4 br_0_58
port 433 nsew
rlabel metal1 s 41532 13800 41568 14141 4 vdd
port 1 nsew
rlabel metal1 s 37932 0 37968 52140 4 br_1_58
port 434 nsew
rlabel metal1 s 38700 0 38736 52140 4 bl_0_59
port 435 nsew
rlabel metal1 s 38484 0 38520 52140 4 bl_1_59
port 436 nsew
rlabel metal1 s 38628 0 38664 52140 4 br_0_59
port 437 nsew
rlabel metal1 s 38412 0 38448 52140 4 br_1_59
port 438 nsew
rlabel metal1 s 38892 0 38928 52140 4 bl_0_60
port 439 nsew
rlabel metal1 s 39108 0 39144 52140 4 bl_1_60
port 440 nsew
rlabel metal1 s 38964 0 39000 52140 4 br_0_60
port 441 nsew
rlabel metal1 s 39180 0 39216 52140 4 br_1_60
port 442 nsew
rlabel metal1 s 39948 0 39984 52140 4 bl_0_61
port 443 nsew
rlabel metal1 s 39732 0 39768 52140 4 bl_1_61
port 444 nsew
rlabel metal1 s 39876 0 39912 52140 4 br_0_61
port 445 nsew
rlabel metal1 s 39660 0 39696 52140 4 br_1_61
port 446 nsew
rlabel metal1 s 40140 0 40176 52140 4 bl_0_62
port 447 nsew
rlabel metal1 s 40356 0 40392 52140 4 bl_1_62
port 448 nsew
rlabel metal1 s 40212 0 40248 52140 4 br_0_62
port 449 nsew
rlabel metal1 s 40428 0 40464 52140 4 br_1_62
port 450 nsew
rlabel metal1 s 41196 0 41232 52140 4 bl_0_63
port 451 nsew
rlabel metal1 s 41532 15380 41568 15721 4 vdd
port 1 nsew
rlabel metal1 s 40980 0 41016 52140 4 bl_1_63
port 452 nsew
rlabel metal1 s 41124 0 41160 52140 4 br_0_63
port 453 nsew
rlabel metal1 s 40908 0 40944 52140 4 br_1_63
port 454 nsew
rlabel metal1 s 41532 17459 41568 17800 4 vdd
port 1 nsew
rlabel metal1 s 41388 0 41424 52140 4 rbl_bl_0_1
port 455 nsew
rlabel metal1 s 41532 16170 41568 16511 4 vdd
port 1 nsew
rlabel metal1 s 41604 0 41640 52140 4 rbl_bl_1_1
port 456 nsew
rlabel metal1 s 41460 0 41496 52140 4 rbl_br_0_1
port 457 nsew
rlabel metal1 s 41676 0 41712 52140 4 rbl_br_1_1
port 458 nsew
rlabel metal1 s 41532 14299 41568 14640 4 vdd
port 1 nsew
rlabel metal1 s 41532 19829 41568 20170 4 vdd
port 1 nsew
rlabel metal1 s 41532 14590 41568 14931 4 vdd
port 1 nsew
rlabel metal1 s 41532 24860 41568 25201 4 vdd
port 1 nsew
rlabel metal1 s 41532 22989 41568 23330 4 vdd
port 1 nsew
rlabel metal1 s 41532 23779 41568 24120 4 vdd
port 1 nsew
rlabel metal1 s 41532 17750 41568 18091 4 vdd
port 1 nsew
rlabel metal1 s 41532 15089 41568 15430 4 vdd
port 1 nsew
rlabel metal1 s 41532 25359 41568 25700 4 vdd
port 1 nsew
rlabel metal1 s 41532 19039 41568 19380 4 vdd
port 1 nsew
rlabel metal1 s 41532 20120 41568 20461 4 vdd
port 1 nsew
rlabel metal1 s 41532 13509 41568 13850 4 vdd
port 1 nsew
rlabel metal1 s 41532 18540 41568 18881 4 vdd
port 1 nsew
rlabel metal1 s 41532 23280 41568 23621 4 vdd
port 1 nsew
rlabel metal1 s 41532 16669 41568 17010 4 vdd
port 1 nsew
rlabel metal1 s 41532 20619 41568 20960 4 vdd
port 1 nsew
rlabel metal1 s 29676 0 29712 52140 4 br_1_45
port 459 nsew
rlabel metal1 s 31476 0 31512 52140 4 br_0_48
port 460 nsew
rlabel metal1 s 30156 0 30192 52140 4 bl_0_46
port 461 nsew
rlabel metal1 s 30372 0 30408 52140 4 bl_1_46
port 462 nsew
rlabel metal1 s 22476 0 22512 52140 4 bl_0_33
port 463 nsew
rlabel metal1 s 30228 0 30264 52140 4 br_0_46
port 464 nsew
rlabel metal1 s 22260 0 22296 52140 4 bl_1_33
port 465 nsew
rlabel metal1 s 22404 0 22440 52140 4 br_0_33
port 466 nsew
rlabel metal1 s 22188 0 22224 52140 4 br_1_33
port 467 nsew
rlabel metal1 s 22668 0 22704 52140 4 bl_0_34
port 468 nsew
rlabel metal1 s 22884 0 22920 52140 4 bl_1_34
port 469 nsew
rlabel metal1 s 22740 0 22776 52140 4 br_0_34
port 470 nsew
rlabel metal1 s 22956 0 22992 52140 4 br_1_34
port 471 nsew
rlabel metal1 s 23724 0 23760 52140 4 bl_0_35
port 472 nsew
rlabel metal1 s 30444 0 30480 52140 4 br_1_46
port 473 nsew
rlabel metal1 s 23508 0 23544 52140 4 bl_1_35
port 474 nsew
rlabel metal1 s 29196 0 29232 52140 4 br_1_44
port 475 nsew
rlabel metal1 s 23652 0 23688 52140 4 br_0_35
port 476 nsew
rlabel metal1 s 23436 0 23472 52140 4 br_1_35
port 477 nsew
rlabel metal1 s 23916 0 23952 52140 4 bl_0_36
port 478 nsew
rlabel metal1 s 31212 0 31248 52140 4 bl_0_47
port 479 nsew
rlabel metal1 s 24132 0 24168 52140 4 bl_1_36
port 480 nsew
rlabel metal1 s 23988 0 24024 52140 4 br_0_36
port 481 nsew
rlabel metal1 s 30996 0 31032 52140 4 bl_1_47
port 482 nsew
rlabel metal1 s 29964 0 30000 52140 4 bl_0_45
port 483 nsew
rlabel metal1 s 24204 0 24240 52140 4 br_1_36
port 484 nsew
rlabel metal1 s 31140 0 31176 52140 4 br_0_47
port 485 nsew
rlabel metal1 s 30924 0 30960 52140 4 br_1_47
port 486 nsew
rlabel metal1 s 24972 0 25008 52140 4 bl_0_37
port 487 nsew
rlabel metal1 s 24756 0 24792 52140 4 bl_1_37
port 488 nsew
rlabel metal1 s 24900 0 24936 52140 4 br_0_37
port 489 nsew
rlabel metal1 s 24684 0 24720 52140 4 br_1_37
port 490 nsew
rlabel metal1 s 25164 0 25200 52140 4 bl_0_38
port 491 nsew
rlabel metal1 s 25380 0 25416 52140 4 bl_1_38
port 492 nsew
rlabel metal1 s 25236 0 25272 52140 4 br_0_38
port 493 nsew
rlabel metal1 s 21420 0 21456 52140 4 bl_0_32
port 494 nsew
rlabel metal1 s 25452 0 25488 52140 4 br_1_38
port 495 nsew
rlabel metal1 s 26220 0 26256 52140 4 bl_0_39
port 496 nsew
rlabel metal1 s 26004 0 26040 52140 4 bl_1_39
port 497 nsew
rlabel metal1 s 26148 0 26184 52140 4 br_0_39
port 498 nsew
rlabel metal1 s 25932 0 25968 52140 4 br_1_39
port 499 nsew
rlabel metal1 s 26412 0 26448 52140 4 bl_0_40
port 500 nsew
rlabel metal1 s 21636 0 21672 52140 4 bl_1_32
port 501 nsew
rlabel metal1 s 26628 0 26664 52140 4 bl_1_40
port 502 nsew
rlabel metal1 s 26484 0 26520 52140 4 br_0_40
port 503 nsew
rlabel metal1 s 21492 0 21528 52140 4 br_0_32
port 504 nsew
rlabel metal1 s 26700 0 26736 52140 4 br_1_40
port 505 nsew
rlabel metal1 s 27468 0 27504 52140 4 bl_0_41
port 506 nsew
rlabel metal1 s 27252 0 27288 52140 4 bl_1_41
port 507 nsew
rlabel metal1 s 29748 0 29784 52140 4 bl_1_45
port 508 nsew
rlabel metal1 s 27396 0 27432 52140 4 br_0_41
port 509 nsew
rlabel metal1 s 27180 0 27216 52140 4 br_1_41
port 510 nsew
rlabel metal1 s 21708 0 21744 52140 4 br_1_32
port 511 nsew
rlabel metal1 s 27660 0 27696 52140 4 bl_0_42
port 512 nsew
rlabel metal1 s 27876 0 27912 52140 4 bl_1_42
port 513 nsew
rlabel metal1 s 31404 0 31440 52140 4 bl_0_48
port 514 nsew
rlabel metal1 s 27732 0 27768 52140 4 br_0_42
port 515 nsew
rlabel metal1 s 27948 0 27984 52140 4 br_1_42
port 516 nsew
rlabel metal1 s 28716 0 28752 52140 4 bl_0_43
port 517 nsew
rlabel metal1 s 28500 0 28536 52140 4 bl_1_43
port 518 nsew
rlabel metal1 s 28644 0 28680 52140 4 br_0_43
port 519 nsew
rlabel metal1 s 28428 0 28464 52140 4 br_1_43
port 520 nsew
rlabel metal1 s 28908 0 28944 52140 4 bl_0_44
port 521 nsew
rlabel metal1 s 29124 0 29160 52140 4 bl_1_44
port 522 nsew
rlabel metal1 s 29892 0 29928 52140 4 br_0_45
port 523 nsew
rlabel metal1 s 28980 0 29016 52140 4 br_0_44
port 524 nsew
rlabel metal1 s 41532 13010 41568 13351 4 vdd
port 1 nsew
rlabel metal1 s 41532 6690 41568 7031 4 vdd
port 1 nsew
rlabel metal1 s 41532 8270 41568 8611 4 vdd
port 1 nsew
rlabel metal1 s 41532 370 41568 711 4 vdd
port 1 nsew
rlabel metal1 s 41532 5609 41568 5950 4 vdd
port 1 nsew
rlabel metal1 s 41532 10640 41568 10981 4 vdd
port 1 nsew
rlabel metal1 s 41532 9060 41568 9401 4 vdd
port 1 nsew
rlabel metal1 s 41532 11929 41568 12270 4 vdd
port 1 nsew
rlabel metal1 s 41532 1659 41568 2000 4 vdd
port 1 nsew
rlabel metal1 s 41532 3530 41568 3871 4 vdd
port 1 nsew
rlabel metal1 s 41532 3239 41568 3580 4 vdd
port 1 nsew
rlabel metal1 s 41532 1950 41568 2291 4 vdd
port 1 nsew
rlabel metal1 s 41532 4819 41568 5160 4 vdd
port 1 nsew
rlabel metal1 s 41532 1160 41568 1501 4 vdd
port 1 nsew
rlabel metal1 s 41532 7979 41568 8320 4 vdd
port 1 nsew
rlabel metal1 s 41532 7480 41568 7821 4 vdd
port 1 nsew
rlabel metal1 s 41532 2449 41568 2790 4 vdd
port 1 nsew
rlabel metal1 s 41532 11139 41568 11480 4 vdd
port 1 nsew
rlabel metal1 s 41532 869 41568 1210 4 vdd
port 1 nsew
rlabel metal1 s 41532 12220 41568 12561 4 vdd
port 1 nsew
rlabel metal1 s 41532 4029 41568 4370 4 vdd
port 1 nsew
rlabel metal1 s 41532 6399 41568 6740 4 vdd
port 1 nsew
rlabel metal1 s 41532 2740 41568 3081 4 vdd
port 1 nsew
rlabel metal1 s 41532 9850 41568 10191 4 vdd
port 1 nsew
rlabel metal1 s 41532 4320 41568 4661 4 vdd
port 1 nsew
rlabel metal1 s 41532 10349 41568 10690 4 vdd
port 1 nsew
rlabel metal1 s 41532 9559 41568 9900 4 vdd
port 1 nsew
rlabel metal1 s 41532 12719 41568 13060 4 vdd
port 1 nsew
rlabel metal1 s 41532 8769 41568 9110 4 vdd
port 1 nsew
rlabel metal1 s 41532 7189 41568 7530 4 vdd
port 1 nsew
rlabel metal1 s 41532 5900 41568 6241 4 vdd
port 1 nsew
rlabel metal1 s 41532 5110 41568 5451 4 vdd
port 1 nsew
rlabel metal1 s 41532 11430 41568 11771 4 vdd
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 42684 630
string GDS_END 7019604
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 6721048
<< end >>
