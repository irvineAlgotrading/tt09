magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 17745 20216 17979 23522
<< pwell >>
rect 28615 7182 31021 7966
rect 28615 6758 29005 7182
rect 28615 6175 28837 6758
rect 30066 5796 32083 6028
rect 30066 5566 30256 5796
rect 19929 4159 20508 5449
rect 22786 5090 30256 5566
rect 20139 2663 20508 4159
rect 26641 4691 30256 5090
rect 26641 4143 28740 4691
rect 22497 2663 22815 3099
rect 20139 2611 22815 2663
rect 18122 2541 22815 2611
rect 16497 2420 22815 2541
rect 22249 1712 22815 2420
rect 26696 1669 28418 2374
rect 26696 805 27005 1669
<< psubdiff >>
rect 28641 7906 28665 7940
rect 28699 7906 28734 7940
rect 28768 7906 28803 7940
rect 28837 7906 28872 7940
rect 28906 7906 28941 7940
rect 28975 7906 29010 7940
rect 29044 7906 29079 7940
rect 29113 7906 29148 7940
rect 29182 7906 29217 7940
rect 29251 7906 29286 7940
rect 29320 7906 29355 7940
rect 29389 7906 29424 7940
rect 29458 7906 29493 7940
rect 29527 7906 29562 7940
rect 29596 7906 29631 7940
rect 29665 7906 29700 7940
rect 29734 7906 29769 7940
rect 29803 7906 29838 7940
rect 29872 7906 29907 7940
rect 29941 7906 29976 7940
rect 30010 7906 30045 7940
rect 30079 7906 30114 7940
rect 30148 7906 30183 7940
rect 30217 7906 30252 7940
rect 30286 7906 30321 7940
rect 30355 7906 30390 7940
rect 30424 7906 30459 7940
rect 30493 7906 30528 7940
rect 30562 7906 30597 7940
rect 28641 7872 30597 7906
rect 28641 7838 28665 7872
rect 28699 7838 28734 7872
rect 28768 7838 28803 7872
rect 28837 7838 28872 7872
rect 28906 7838 28941 7872
rect 28975 7838 29010 7872
rect 29044 7838 29079 7872
rect 29113 7838 29148 7872
rect 29182 7838 29217 7872
rect 29251 7838 29286 7872
rect 29320 7838 29355 7872
rect 29389 7838 29424 7872
rect 29458 7838 29493 7872
rect 29527 7838 29562 7872
rect 29596 7838 29631 7872
rect 29665 7838 29700 7872
rect 29734 7838 29769 7872
rect 29803 7838 29838 7872
rect 29872 7838 29907 7872
rect 29941 7838 29976 7872
rect 30010 7838 30045 7872
rect 30079 7838 30114 7872
rect 30148 7838 30183 7872
rect 30217 7838 30252 7872
rect 30286 7838 30321 7872
rect 30355 7838 30390 7872
rect 30424 7838 30459 7872
rect 30493 7838 30528 7872
rect 30562 7838 30597 7872
rect 28641 7804 30597 7838
rect 28641 7770 28665 7804
rect 28699 7770 28734 7804
rect 28768 7770 28803 7804
rect 28837 7770 28872 7804
rect 28906 7770 28941 7804
rect 28975 7770 29010 7804
rect 29044 7770 29079 7804
rect 29113 7770 29148 7804
rect 29182 7770 29217 7804
rect 29251 7770 29286 7804
rect 29320 7770 29355 7804
rect 29389 7770 29424 7804
rect 29458 7770 29493 7804
rect 29527 7770 29562 7804
rect 29596 7770 29631 7804
rect 29665 7770 29700 7804
rect 29734 7770 29769 7804
rect 29803 7770 29838 7804
rect 29872 7770 29907 7804
rect 29941 7770 29976 7804
rect 30010 7770 30045 7804
rect 30079 7770 30114 7804
rect 30148 7770 30183 7804
rect 30217 7770 30252 7804
rect 30286 7770 30321 7804
rect 30355 7770 30390 7804
rect 30424 7770 30459 7804
rect 30493 7770 30528 7804
rect 30562 7770 30597 7804
rect 28641 7736 30597 7770
rect 28641 7702 28665 7736
rect 28699 7702 28734 7736
rect 28768 7702 28803 7736
rect 28837 7702 28872 7736
rect 28906 7702 28941 7736
rect 28975 7702 29010 7736
rect 29044 7702 29079 7736
rect 29113 7702 29148 7736
rect 29182 7702 29217 7736
rect 29251 7702 29286 7736
rect 29320 7702 29355 7736
rect 29389 7702 29424 7736
rect 29458 7702 29493 7736
rect 29527 7702 29562 7736
rect 29596 7702 29631 7736
rect 29665 7702 29700 7736
rect 29734 7702 29769 7736
rect 29803 7702 29838 7736
rect 29872 7702 29907 7736
rect 29941 7702 29976 7736
rect 30010 7702 30045 7736
rect 30079 7702 30114 7736
rect 30148 7702 30183 7736
rect 30217 7702 30252 7736
rect 30286 7702 30321 7736
rect 30355 7702 30390 7736
rect 30424 7702 30459 7736
rect 30493 7702 30528 7736
rect 30562 7702 30597 7736
rect 28641 7668 30597 7702
rect 28641 7634 28665 7668
rect 28699 7634 28734 7668
rect 28768 7634 28803 7668
rect 28837 7634 28872 7668
rect 28906 7634 28941 7668
rect 28975 7634 29010 7668
rect 29044 7634 29079 7668
rect 29113 7634 29148 7668
rect 29182 7634 29217 7668
rect 29251 7634 29286 7668
rect 29320 7634 29355 7668
rect 29389 7634 29424 7668
rect 29458 7634 29493 7668
rect 29527 7634 29562 7668
rect 29596 7634 29631 7668
rect 29665 7634 29700 7668
rect 29734 7634 29769 7668
rect 29803 7634 29838 7668
rect 29872 7634 29907 7668
rect 29941 7634 29976 7668
rect 30010 7634 30045 7668
rect 30079 7634 30114 7668
rect 30148 7634 30183 7668
rect 30217 7634 30252 7668
rect 30286 7634 30321 7668
rect 30355 7634 30390 7668
rect 30424 7634 30459 7668
rect 30493 7634 30528 7668
rect 30562 7634 30597 7668
rect 28641 7600 30597 7634
rect 28641 7566 28665 7600
rect 28699 7566 28734 7600
rect 28768 7566 28803 7600
rect 28837 7566 28872 7600
rect 28906 7566 28941 7600
rect 28975 7566 29010 7600
rect 29044 7566 29079 7600
rect 29113 7566 29148 7600
rect 29182 7566 29217 7600
rect 29251 7566 29286 7600
rect 29320 7566 29355 7600
rect 29389 7566 29424 7600
rect 29458 7566 29493 7600
rect 29527 7566 29562 7600
rect 29596 7566 29631 7600
rect 29665 7566 29700 7600
rect 29734 7566 29769 7600
rect 29803 7566 29838 7600
rect 29872 7566 29907 7600
rect 29941 7566 29976 7600
rect 30010 7566 30045 7600
rect 30079 7566 30114 7600
rect 30148 7566 30183 7600
rect 30217 7566 30252 7600
rect 30286 7566 30321 7600
rect 30355 7566 30390 7600
rect 30424 7566 30459 7600
rect 30493 7566 30528 7600
rect 30562 7566 30597 7600
rect 28641 7532 30597 7566
rect 28641 7498 28665 7532
rect 28699 7498 28734 7532
rect 28768 7498 28803 7532
rect 28837 7498 28872 7532
rect 28906 7498 28941 7532
rect 28975 7498 29010 7532
rect 29044 7498 29079 7532
rect 29113 7498 29148 7532
rect 29182 7498 29217 7532
rect 29251 7498 29286 7532
rect 29320 7498 29355 7532
rect 29389 7498 29424 7532
rect 29458 7498 29493 7532
rect 29527 7498 29562 7532
rect 29596 7498 29631 7532
rect 29665 7498 29700 7532
rect 29734 7498 29769 7532
rect 29803 7498 29838 7532
rect 29872 7498 29907 7532
rect 29941 7498 29976 7532
rect 30010 7498 30045 7532
rect 30079 7498 30114 7532
rect 30148 7498 30183 7532
rect 30217 7498 30252 7532
rect 30286 7498 30321 7532
rect 30355 7498 30390 7532
rect 30424 7498 30459 7532
rect 30493 7498 30528 7532
rect 30562 7498 30597 7532
rect 28641 7464 30597 7498
rect 28641 7430 28665 7464
rect 28699 7430 28734 7464
rect 28768 7430 28803 7464
rect 28837 7430 28872 7464
rect 28906 7430 28941 7464
rect 28975 7430 29010 7464
rect 29044 7430 29079 7464
rect 29113 7430 29148 7464
rect 29182 7430 29217 7464
rect 29251 7430 29286 7464
rect 29320 7430 29355 7464
rect 29389 7430 29424 7464
rect 29458 7430 29493 7464
rect 29527 7430 29562 7464
rect 29596 7430 29631 7464
rect 29665 7430 29700 7464
rect 29734 7430 29769 7464
rect 29803 7430 29838 7464
rect 29872 7430 29907 7464
rect 29941 7430 29976 7464
rect 30010 7430 30045 7464
rect 30079 7430 30114 7464
rect 30148 7430 30183 7464
rect 30217 7430 30252 7464
rect 30286 7430 30321 7464
rect 30355 7430 30390 7464
rect 30424 7430 30459 7464
rect 30493 7430 30528 7464
rect 30562 7430 30597 7464
rect 28641 7396 30597 7430
rect 28641 7362 28665 7396
rect 28699 7362 28734 7396
rect 28768 7362 28803 7396
rect 28837 7362 28872 7396
rect 28906 7362 28941 7396
rect 28975 7362 29010 7396
rect 29044 7362 29079 7396
rect 29113 7362 29148 7396
rect 29182 7362 29217 7396
rect 29251 7362 29286 7396
rect 29320 7362 29355 7396
rect 29389 7362 29424 7396
rect 29458 7362 29493 7396
rect 29527 7362 29562 7396
rect 29596 7362 29631 7396
rect 29665 7362 29700 7396
rect 29734 7362 29769 7396
rect 29803 7362 29838 7396
rect 29872 7362 29907 7396
rect 29941 7362 29976 7396
rect 30010 7362 30045 7396
rect 30079 7362 30114 7396
rect 30148 7362 30183 7396
rect 30217 7362 30252 7396
rect 30286 7362 30321 7396
rect 30355 7362 30390 7396
rect 30424 7362 30459 7396
rect 30493 7362 30528 7396
rect 30562 7362 30597 7396
rect 28641 7328 30597 7362
rect 28641 7294 28665 7328
rect 28699 7294 28734 7328
rect 28768 7294 28803 7328
rect 28837 7294 28872 7328
rect 28906 7294 28941 7328
rect 28975 7294 29010 7328
rect 29044 7294 29079 7328
rect 29113 7294 29148 7328
rect 29182 7294 29217 7328
rect 29251 7294 29286 7328
rect 29320 7294 29355 7328
rect 29389 7294 29424 7328
rect 29458 7294 29493 7328
rect 29527 7294 29562 7328
rect 29596 7294 29631 7328
rect 29665 7294 29700 7328
rect 29734 7294 29769 7328
rect 29803 7294 29838 7328
rect 29872 7294 29907 7328
rect 29941 7294 29976 7328
rect 30010 7294 30045 7328
rect 30079 7294 30114 7328
rect 30148 7294 30183 7328
rect 30217 7294 30252 7328
rect 30286 7294 30321 7328
rect 30355 7294 30390 7328
rect 30424 7294 30459 7328
rect 30493 7294 30528 7328
rect 30562 7294 30597 7328
rect 30971 7294 30995 7940
rect 28641 7221 30995 7294
rect 28811 7208 30995 7221
rect 28811 6915 28979 7208
rect 28641 6880 28979 6915
rect 28675 6846 28709 6880
rect 28743 6846 28777 6880
rect 28811 6846 28979 6880
rect 28641 6811 28979 6846
rect 28675 6777 28709 6811
rect 28743 6777 28777 6811
rect 28811 6784 28979 6811
rect 28641 6742 28811 6777
rect 28675 6708 28709 6742
rect 28743 6708 28777 6742
rect 28641 6673 28811 6708
rect 28675 6639 28709 6673
rect 28743 6639 28777 6673
rect 28641 6604 28811 6639
rect 28675 6570 28709 6604
rect 28743 6570 28777 6604
rect 28641 6535 28811 6570
rect 28675 6501 28709 6535
rect 28743 6501 28777 6535
rect 28641 6466 28811 6501
rect 28675 6432 28709 6466
rect 28743 6432 28777 6466
rect 28641 6397 28811 6432
rect 28675 6363 28709 6397
rect 28743 6363 28777 6397
rect 28641 6328 28811 6363
rect 28675 6294 28709 6328
rect 28743 6294 28777 6328
rect 28641 6259 28811 6294
rect 28675 6225 28709 6259
rect 28743 6225 28777 6259
rect 28641 6201 28811 6225
rect 26667 4169 26708 5042
rect 26722 831 26979 860
<< mvpsubdiff >>
rect 30092 6001 32057 6002
rect 30092 5967 30214 6001
rect 30248 5967 30283 6001
rect 30317 5967 30352 6001
rect 30386 5967 30421 6001
rect 30455 5967 30490 6001
rect 30524 5967 30559 6001
rect 30593 5967 30628 6001
rect 30662 5967 30697 6001
rect 30731 5967 30766 6001
rect 30800 5967 30835 6001
rect 30869 5967 30904 6001
rect 30938 5967 30973 6001
rect 31007 5967 31042 6001
rect 31076 5967 31111 6001
rect 31145 5967 31180 6001
rect 31214 5967 31249 6001
rect 31283 5967 31318 6001
rect 31352 5967 31387 6001
rect 31421 5967 31455 6001
rect 31489 5967 31523 6001
rect 31557 5967 31591 6001
rect 31625 5967 31659 6001
rect 31693 5967 31727 6001
rect 31761 5967 31795 6001
rect 31829 5967 31863 6001
rect 31897 5967 31931 6001
rect 31965 5967 31999 6001
rect 32033 5967 32057 6001
rect 30092 5929 32057 5967
rect 30092 5895 30214 5929
rect 30248 5895 30283 5929
rect 30317 5895 30352 5929
rect 30386 5895 30421 5929
rect 30455 5895 30490 5929
rect 30524 5895 30559 5929
rect 30593 5895 30628 5929
rect 30662 5895 30697 5929
rect 30731 5895 30766 5929
rect 30800 5895 30835 5929
rect 30869 5895 30904 5929
rect 30938 5895 30973 5929
rect 31007 5895 31042 5929
rect 31076 5895 31111 5929
rect 31145 5895 31180 5929
rect 31214 5895 31249 5929
rect 31283 5895 31318 5929
rect 31352 5895 31387 5929
rect 31421 5895 31455 5929
rect 31489 5895 31523 5929
rect 31557 5895 31591 5929
rect 31625 5895 31659 5929
rect 31693 5895 31727 5929
rect 31761 5895 31795 5929
rect 31829 5895 31863 5929
rect 31897 5895 31931 5929
rect 31965 5895 31999 5929
rect 32033 5895 32057 5929
rect 30092 5857 32057 5895
rect 30092 5823 30214 5857
rect 30248 5823 30283 5857
rect 30317 5823 30352 5857
rect 30386 5823 30421 5857
rect 30455 5823 30490 5857
rect 30524 5823 30559 5857
rect 30593 5823 30628 5857
rect 30662 5823 30697 5857
rect 30731 5823 30766 5857
rect 30800 5823 30835 5857
rect 30869 5823 30904 5857
rect 30938 5823 30973 5857
rect 31007 5823 31042 5857
rect 31076 5823 31111 5857
rect 31145 5823 31180 5857
rect 31214 5823 31249 5857
rect 31283 5823 31318 5857
rect 31352 5823 31387 5857
rect 31421 5823 31455 5857
rect 31489 5823 31523 5857
rect 31557 5823 31591 5857
rect 31625 5823 31659 5857
rect 31693 5823 31727 5857
rect 31761 5823 31795 5857
rect 31829 5823 31863 5857
rect 31897 5823 31931 5857
rect 31965 5823 31999 5857
rect 32033 5823 32057 5857
rect 30092 5822 32057 5823
rect 30092 5540 30230 5822
rect 22812 5499 30230 5540
rect 22812 5465 22836 5499
rect 22870 5465 22905 5499
rect 22939 5465 22974 5499
rect 23008 5465 23043 5499
rect 23077 5465 23112 5499
rect 23146 5465 23181 5499
rect 23215 5465 23250 5499
rect 23284 5465 23319 5499
rect 23353 5465 23388 5499
rect 23422 5465 23457 5499
rect 23491 5465 23526 5499
rect 23560 5465 23595 5499
rect 23629 5465 23664 5499
rect 23698 5465 23733 5499
rect 23767 5465 23802 5499
rect 23836 5465 23871 5499
rect 23905 5465 23940 5499
rect 23974 5465 24009 5499
rect 24043 5465 24078 5499
rect 24112 5465 24147 5499
rect 24181 5465 24216 5499
rect 24250 5465 24285 5499
rect 24319 5465 24354 5499
rect 24388 5465 24423 5499
rect 24457 5465 24492 5499
rect 24526 5465 24561 5499
rect 24595 5465 24630 5499
rect 24664 5465 24699 5499
rect 24733 5465 24768 5499
rect 24802 5465 24837 5499
rect 24871 5465 24906 5499
rect 24940 5465 24975 5499
rect 25009 5465 25044 5499
rect 25078 5465 25113 5499
rect 25147 5465 25181 5499
rect 25215 5465 25249 5499
rect 25283 5465 25317 5499
rect 25351 5465 25385 5499
rect 25419 5465 25453 5499
rect 25487 5465 25521 5499
rect 25555 5465 25589 5499
rect 25623 5465 25657 5499
rect 25691 5465 25725 5499
rect 25759 5465 25793 5499
rect 25827 5465 25861 5499
rect 25895 5465 25929 5499
rect 25963 5465 25997 5499
rect 26031 5465 26065 5499
rect 26099 5465 26133 5499
rect 26167 5465 26201 5499
rect 26235 5465 26269 5499
rect 26303 5465 26337 5499
rect 26371 5465 26405 5499
rect 26439 5465 26473 5499
rect 26507 5465 26541 5499
rect 26575 5465 26609 5499
rect 26643 5465 26740 5499
rect 26774 5465 26809 5499
rect 26843 5465 26878 5499
rect 26912 5465 26947 5499
rect 26981 5465 27016 5499
rect 27050 5465 27085 5499
rect 27119 5465 27154 5499
rect 27188 5465 27223 5499
rect 27257 5465 27292 5499
rect 27326 5465 27361 5499
rect 27395 5465 27430 5499
rect 27464 5465 27499 5499
rect 27533 5465 27568 5499
rect 22812 5431 27568 5465
rect 19955 5399 20482 5423
rect 20125 5365 20167 5399
rect 20201 5365 20247 5399
rect 20281 5365 20327 5399
rect 20361 5365 20407 5399
rect 20441 5365 20482 5399
rect 20125 5331 20482 5365
rect 20125 5297 20167 5331
rect 20201 5297 20247 5331
rect 20281 5297 20327 5331
rect 20361 5297 20407 5331
rect 20441 5297 20482 5331
rect 20125 5263 20482 5297
rect 20125 5229 20167 5263
rect 20201 5229 20247 5263
rect 20281 5229 20327 5263
rect 20361 5229 20407 5263
rect 20441 5229 20482 5263
rect 20125 5195 20482 5229
rect 20125 5161 20167 5195
rect 20201 5161 20247 5195
rect 20281 5161 20327 5195
rect 20361 5161 20407 5195
rect 20441 5161 20482 5195
rect 20125 5127 20482 5161
rect 20125 5093 20167 5127
rect 20201 5093 20247 5127
rect 20281 5093 20327 5127
rect 20361 5093 20407 5127
rect 20441 5093 20482 5127
rect 22812 5421 26740 5431
rect 22812 5387 22836 5421
rect 22870 5387 22905 5421
rect 22939 5387 22974 5421
rect 23008 5387 23043 5421
rect 23077 5387 23112 5421
rect 23146 5387 23181 5421
rect 23215 5387 23250 5421
rect 23284 5387 23319 5421
rect 23353 5387 23388 5421
rect 23422 5387 23457 5421
rect 23491 5387 23526 5421
rect 23560 5387 23595 5421
rect 23629 5387 23664 5421
rect 23698 5387 23733 5421
rect 23767 5387 23802 5421
rect 23836 5387 23871 5421
rect 23905 5387 23940 5421
rect 23974 5387 24009 5421
rect 24043 5387 24078 5421
rect 24112 5387 24147 5421
rect 24181 5387 24216 5421
rect 24250 5387 24285 5421
rect 24319 5387 24354 5421
rect 24388 5387 24423 5421
rect 24457 5387 24492 5421
rect 24526 5387 24561 5421
rect 24595 5387 24630 5421
rect 24664 5387 24699 5421
rect 24733 5387 24768 5421
rect 24802 5387 24837 5421
rect 24871 5387 24906 5421
rect 24940 5387 24975 5421
rect 25009 5387 25044 5421
rect 25078 5387 25113 5421
rect 25147 5387 25181 5421
rect 25215 5387 25249 5421
rect 25283 5387 25317 5421
rect 25351 5387 25385 5421
rect 25419 5387 25453 5421
rect 25487 5387 25521 5421
rect 25555 5387 25589 5421
rect 25623 5387 25657 5421
rect 25691 5387 25725 5421
rect 25759 5387 25793 5421
rect 25827 5387 25861 5421
rect 25895 5387 25929 5421
rect 25963 5387 25997 5421
rect 26031 5387 26065 5421
rect 26099 5387 26133 5421
rect 26167 5387 26201 5421
rect 26235 5387 26269 5421
rect 26303 5387 26337 5421
rect 26371 5387 26405 5421
rect 26439 5387 26473 5421
rect 26507 5387 26541 5421
rect 26575 5387 26609 5421
rect 26643 5397 26740 5421
rect 26774 5397 26809 5431
rect 26843 5397 26878 5431
rect 26912 5397 26947 5431
rect 26981 5397 27016 5431
rect 27050 5397 27085 5431
rect 27119 5397 27154 5431
rect 27188 5397 27223 5431
rect 27257 5397 27292 5431
rect 27326 5397 27361 5431
rect 27395 5397 27430 5431
rect 27464 5397 27499 5431
rect 27533 5397 27568 5431
rect 26643 5387 27568 5397
rect 22812 5363 27568 5387
rect 22812 5343 26740 5363
rect 22812 5309 22836 5343
rect 22870 5309 22905 5343
rect 22939 5309 22974 5343
rect 23008 5309 23043 5343
rect 23077 5309 23112 5343
rect 23146 5309 23181 5343
rect 23215 5309 23250 5343
rect 23284 5309 23319 5343
rect 23353 5309 23388 5343
rect 23422 5309 23457 5343
rect 23491 5309 23526 5343
rect 23560 5309 23595 5343
rect 23629 5309 23664 5343
rect 23698 5309 23733 5343
rect 23767 5309 23802 5343
rect 23836 5309 23871 5343
rect 23905 5309 23940 5343
rect 23974 5309 24009 5343
rect 24043 5309 24078 5343
rect 24112 5309 24147 5343
rect 24181 5309 24216 5343
rect 24250 5309 24285 5343
rect 24319 5309 24354 5343
rect 24388 5309 24423 5343
rect 24457 5309 24492 5343
rect 24526 5309 24561 5343
rect 24595 5309 24630 5343
rect 24664 5309 24699 5343
rect 24733 5309 24768 5343
rect 24802 5309 24837 5343
rect 24871 5309 24906 5343
rect 24940 5309 24975 5343
rect 25009 5309 25044 5343
rect 25078 5309 25113 5343
rect 25147 5309 25181 5343
rect 25215 5309 25249 5343
rect 25283 5309 25317 5343
rect 25351 5309 25385 5343
rect 25419 5309 25453 5343
rect 25487 5309 25521 5343
rect 25555 5309 25589 5343
rect 25623 5309 25657 5343
rect 25691 5309 25725 5343
rect 25759 5309 25793 5343
rect 25827 5309 25861 5343
rect 25895 5309 25929 5343
rect 25963 5309 25997 5343
rect 26031 5309 26065 5343
rect 26099 5309 26133 5343
rect 26167 5309 26201 5343
rect 26235 5309 26269 5343
rect 26303 5309 26337 5343
rect 26371 5309 26405 5343
rect 26439 5309 26473 5343
rect 26507 5309 26541 5343
rect 26575 5309 26609 5343
rect 26643 5329 26740 5343
rect 26774 5329 26809 5363
rect 26843 5329 26878 5363
rect 26912 5329 26947 5363
rect 26981 5329 27016 5363
rect 27050 5329 27085 5363
rect 27119 5329 27154 5363
rect 27188 5329 27223 5363
rect 27257 5329 27292 5363
rect 27326 5329 27361 5363
rect 27395 5329 27430 5363
rect 27464 5329 27499 5363
rect 27533 5329 27568 5363
rect 26643 5309 27568 5329
rect 22812 5295 27568 5309
rect 22812 5265 26740 5295
rect 22812 5231 22836 5265
rect 22870 5231 22905 5265
rect 22939 5231 22974 5265
rect 23008 5231 23043 5265
rect 23077 5231 23112 5265
rect 23146 5231 23181 5265
rect 23215 5231 23250 5265
rect 23284 5231 23319 5265
rect 23353 5231 23388 5265
rect 23422 5231 23457 5265
rect 23491 5231 23526 5265
rect 23560 5231 23595 5265
rect 23629 5231 23664 5265
rect 23698 5231 23733 5265
rect 23767 5231 23802 5265
rect 23836 5231 23871 5265
rect 23905 5231 23940 5265
rect 23974 5231 24009 5265
rect 24043 5231 24078 5265
rect 24112 5231 24147 5265
rect 24181 5231 24216 5265
rect 24250 5231 24285 5265
rect 24319 5231 24354 5265
rect 24388 5231 24423 5265
rect 24457 5231 24492 5265
rect 24526 5231 24561 5265
rect 24595 5231 24630 5265
rect 24664 5231 24699 5265
rect 24733 5231 24768 5265
rect 24802 5231 24837 5265
rect 24871 5231 24906 5265
rect 24940 5231 24975 5265
rect 25009 5231 25044 5265
rect 25078 5231 25113 5265
rect 25147 5231 25181 5265
rect 25215 5231 25249 5265
rect 25283 5231 25317 5265
rect 25351 5231 25385 5265
rect 25419 5231 25453 5265
rect 25487 5231 25521 5265
rect 25555 5231 25589 5265
rect 25623 5231 25657 5265
rect 25691 5231 25725 5265
rect 25759 5231 25793 5265
rect 25827 5231 25861 5265
rect 25895 5231 25929 5265
rect 25963 5231 25997 5265
rect 26031 5231 26065 5265
rect 26099 5231 26133 5265
rect 26167 5231 26201 5265
rect 26235 5231 26269 5265
rect 26303 5231 26337 5265
rect 26371 5231 26405 5265
rect 26439 5231 26473 5265
rect 26507 5231 26541 5265
rect 26575 5231 26609 5265
rect 26643 5261 26740 5265
rect 26774 5261 26809 5295
rect 26843 5261 26878 5295
rect 26912 5261 26947 5295
rect 26981 5261 27016 5295
rect 27050 5261 27085 5295
rect 27119 5261 27154 5295
rect 27188 5261 27223 5295
rect 27257 5261 27292 5295
rect 27326 5261 27361 5295
rect 27395 5261 27430 5295
rect 27464 5261 27499 5295
rect 27533 5261 27568 5295
rect 26643 5231 27568 5261
rect 22812 5227 27568 5231
rect 22812 5193 26740 5227
rect 26774 5193 26809 5227
rect 26843 5193 26878 5227
rect 26912 5193 26947 5227
rect 26981 5193 27016 5227
rect 27050 5193 27085 5227
rect 27119 5193 27154 5227
rect 27188 5193 27223 5227
rect 27257 5193 27292 5227
rect 27326 5193 27361 5227
rect 27395 5193 27430 5227
rect 27464 5193 27499 5227
rect 27533 5193 27568 5227
rect 22812 5187 27568 5193
rect 22812 5153 22836 5187
rect 22870 5153 22905 5187
rect 22939 5153 22974 5187
rect 23008 5153 23043 5187
rect 23077 5153 23112 5187
rect 23146 5153 23181 5187
rect 23215 5153 23250 5187
rect 23284 5153 23319 5187
rect 23353 5153 23388 5187
rect 23422 5153 23457 5187
rect 23491 5153 23526 5187
rect 23560 5153 23595 5187
rect 23629 5153 23664 5187
rect 23698 5153 23733 5187
rect 23767 5153 23802 5187
rect 23836 5153 23871 5187
rect 23905 5153 23940 5187
rect 23974 5153 24009 5187
rect 24043 5153 24078 5187
rect 24112 5153 24147 5187
rect 24181 5153 24216 5187
rect 24250 5153 24285 5187
rect 24319 5153 24354 5187
rect 24388 5153 24423 5187
rect 24457 5153 24492 5187
rect 24526 5153 24561 5187
rect 24595 5153 24630 5187
rect 24664 5153 24699 5187
rect 24733 5153 24768 5187
rect 24802 5153 24837 5187
rect 24871 5153 24906 5187
rect 24940 5153 24975 5187
rect 25009 5153 25044 5187
rect 25078 5153 25113 5187
rect 25147 5153 25181 5187
rect 25215 5153 25249 5187
rect 25283 5153 25317 5187
rect 25351 5153 25385 5187
rect 25419 5153 25453 5187
rect 25487 5153 25521 5187
rect 25555 5153 25589 5187
rect 25623 5153 25657 5187
rect 25691 5153 25725 5187
rect 25759 5153 25793 5187
rect 25827 5153 25861 5187
rect 25895 5153 25929 5187
rect 25963 5153 25997 5187
rect 26031 5153 26065 5187
rect 26099 5153 26133 5187
rect 26167 5153 26201 5187
rect 26235 5153 26269 5187
rect 26303 5153 26337 5187
rect 26371 5153 26405 5187
rect 26439 5153 26473 5187
rect 26507 5153 26541 5187
rect 26575 5153 26609 5187
rect 26643 5159 27568 5187
rect 26643 5153 26740 5159
rect 22812 5125 26740 5153
rect 26774 5125 26809 5159
rect 26843 5125 26878 5159
rect 26912 5125 26947 5159
rect 26981 5125 27016 5159
rect 27050 5125 27085 5159
rect 27119 5125 27154 5159
rect 27188 5125 27223 5159
rect 27257 5125 27292 5159
rect 27326 5125 27361 5159
rect 27395 5125 27430 5159
rect 27464 5125 27499 5159
rect 27533 5125 27568 5159
rect 22812 5116 27568 5125
rect 20125 5059 20482 5093
rect 20125 5025 20167 5059
rect 20201 5025 20247 5059
rect 20281 5025 20327 5059
rect 20361 5025 20407 5059
rect 20441 5025 20482 5059
rect 20125 4991 20482 5025
rect 20125 4957 20167 4991
rect 20201 4957 20247 4991
rect 20281 4957 20327 4991
rect 20361 4957 20407 4991
rect 20441 4957 20482 4991
rect 20125 4923 20482 4957
rect 20125 4889 20167 4923
rect 20201 4889 20247 4923
rect 20281 4889 20327 4923
rect 20361 4889 20407 4923
rect 20441 4889 20482 4923
rect 20125 4855 20482 4889
rect 20125 4821 20167 4855
rect 20201 4821 20247 4855
rect 20281 4821 20327 4855
rect 20361 4821 20407 4855
rect 20441 4821 20482 4855
rect 20125 4787 20482 4821
rect 20125 4753 20167 4787
rect 20201 4753 20247 4787
rect 20281 4753 20327 4787
rect 20361 4753 20407 4787
rect 20441 4753 20482 4787
rect 20125 4719 20482 4753
rect 20125 4685 20167 4719
rect 20201 4685 20247 4719
rect 20281 4685 20327 4719
rect 20361 4685 20407 4719
rect 20441 4685 20482 4719
rect 20125 4651 20482 4685
rect 20125 4617 20167 4651
rect 20201 4617 20247 4651
rect 20281 4617 20327 4651
rect 20361 4617 20407 4651
rect 20441 4617 20482 4651
rect 20125 4583 20482 4617
rect 20125 4549 20167 4583
rect 20201 4549 20247 4583
rect 20281 4549 20327 4583
rect 20361 4549 20407 4583
rect 20441 4549 20482 4583
rect 20125 4515 20482 4549
rect 20125 4481 20167 4515
rect 20201 4481 20247 4515
rect 20281 4481 20327 4515
rect 20361 4481 20407 4515
rect 20441 4481 20482 4515
rect 20125 4447 20482 4481
rect 20125 4413 20167 4447
rect 20201 4413 20247 4447
rect 20281 4413 20327 4447
rect 20361 4413 20407 4447
rect 20441 4413 20482 4447
rect 20125 4379 20482 4413
rect 20125 4345 20167 4379
rect 20201 4345 20247 4379
rect 20281 4345 20327 4379
rect 20361 4345 20407 4379
rect 20441 4345 20482 4379
rect 20125 4311 20482 4345
rect 20125 4277 20167 4311
rect 20201 4277 20247 4311
rect 20281 4277 20327 4311
rect 20361 4277 20407 4311
rect 20441 4277 20482 4311
rect 20125 4243 20482 4277
rect 20125 4209 20167 4243
rect 20201 4209 20247 4243
rect 20281 4209 20327 4243
rect 20361 4209 20407 4243
rect 20441 4209 20482 4243
rect 19955 4185 20482 4209
rect 20165 4175 20482 4185
rect 20165 4141 20167 4175
rect 20201 4141 20247 4175
rect 20281 4141 20327 4175
rect 20361 4141 20407 4175
rect 20441 4141 20482 4175
rect 26667 5091 27568 5116
rect 26667 5057 26740 5091
rect 26774 5057 26809 5091
rect 26843 5057 26878 5091
rect 26912 5057 26947 5091
rect 26981 5057 27016 5091
rect 27050 5057 27085 5091
rect 27119 5057 27154 5091
rect 27188 5057 27223 5091
rect 27257 5057 27292 5091
rect 27326 5057 27361 5091
rect 27395 5057 27430 5091
rect 27464 5057 27499 5091
rect 27533 5057 27568 5091
rect 26667 5042 27568 5057
rect 26708 5023 27568 5042
rect 26708 4989 26740 5023
rect 26774 4989 26809 5023
rect 26843 4989 26878 5023
rect 26912 4989 26947 5023
rect 26981 4989 27016 5023
rect 27050 4989 27085 5023
rect 27119 4989 27154 5023
rect 27188 4989 27223 5023
rect 27257 4989 27292 5023
rect 27326 4989 27361 5023
rect 27395 4989 27430 5023
rect 27464 4989 27499 5023
rect 27533 4989 27568 5023
rect 26708 4955 27568 4989
rect 26708 4921 26740 4955
rect 26774 4921 26809 4955
rect 26843 4921 26878 4955
rect 26912 4921 26947 4955
rect 26981 4921 27016 4955
rect 27050 4921 27085 4955
rect 27119 4921 27154 4955
rect 27188 4921 27223 4955
rect 27257 4921 27292 4955
rect 27326 4921 27361 4955
rect 27395 4921 27430 4955
rect 27464 4921 27499 4955
rect 27533 4921 27568 4955
rect 26708 4887 27568 4921
rect 26708 4853 26740 4887
rect 26774 4853 26809 4887
rect 26843 4853 26878 4887
rect 26912 4853 26947 4887
rect 26981 4853 27016 4887
rect 27050 4853 27085 4887
rect 27119 4853 27154 4887
rect 27188 4853 27223 4887
rect 27257 4853 27292 4887
rect 27326 4853 27361 4887
rect 27395 4853 27430 4887
rect 27464 4853 27499 4887
rect 27533 4853 27568 4887
rect 26708 4819 27568 4853
rect 26708 4785 26740 4819
rect 26774 4785 26809 4819
rect 26843 4785 26878 4819
rect 26912 4785 26947 4819
rect 26981 4785 27016 4819
rect 27050 4785 27085 4819
rect 27119 4785 27154 4819
rect 27188 4785 27223 4819
rect 27257 4785 27292 4819
rect 27326 4785 27361 4819
rect 27395 4785 27430 4819
rect 27464 4785 27499 4819
rect 27533 4785 27568 4819
rect 26708 4751 27568 4785
rect 26708 4717 26740 4751
rect 26774 4717 26809 4751
rect 26843 4717 26878 4751
rect 26912 4717 26947 4751
rect 26981 4717 27016 4751
rect 27050 4717 27085 4751
rect 27119 4717 27154 4751
rect 27188 4717 27223 4751
rect 27257 4717 27292 4751
rect 27326 4717 27361 4751
rect 27395 4717 27430 4751
rect 27464 4717 27499 4751
rect 27533 4717 27568 4751
rect 26708 4683 27568 4717
rect 26708 4649 26740 4683
rect 26774 4649 26809 4683
rect 26843 4649 26878 4683
rect 26912 4649 26947 4683
rect 26981 4649 27016 4683
rect 27050 4649 27085 4683
rect 27119 4649 27154 4683
rect 27188 4649 27223 4683
rect 27257 4649 27292 4683
rect 27326 4649 27361 4683
rect 27395 4649 27430 4683
rect 27464 4649 27499 4683
rect 27533 4649 27568 4683
rect 26708 4615 27568 4649
rect 26708 4581 26740 4615
rect 26774 4581 26809 4615
rect 26843 4581 26878 4615
rect 26912 4581 26947 4615
rect 26981 4581 27016 4615
rect 27050 4581 27085 4615
rect 27119 4581 27154 4615
rect 27188 4581 27223 4615
rect 27257 4581 27292 4615
rect 27326 4581 27361 4615
rect 27395 4581 27430 4615
rect 27464 4581 27499 4615
rect 27533 4581 27568 4615
rect 26708 4547 27568 4581
rect 26708 4513 26740 4547
rect 26774 4513 26809 4547
rect 26843 4513 26878 4547
rect 26912 4513 26947 4547
rect 26981 4513 27016 4547
rect 27050 4513 27085 4547
rect 27119 4513 27154 4547
rect 27188 4513 27223 4547
rect 27257 4513 27292 4547
rect 27326 4513 27361 4547
rect 27395 4513 27430 4547
rect 27464 4513 27499 4547
rect 27533 4513 27568 4547
rect 26708 4479 27568 4513
rect 26708 4445 26740 4479
rect 26774 4445 26809 4479
rect 26843 4445 26878 4479
rect 26912 4445 26947 4479
rect 26981 4445 27016 4479
rect 27050 4445 27085 4479
rect 27119 4445 27154 4479
rect 27188 4445 27223 4479
rect 27257 4445 27292 4479
rect 27326 4445 27361 4479
rect 27395 4445 27430 4479
rect 27464 4445 27499 4479
rect 27533 4445 27568 4479
rect 26708 4411 27568 4445
rect 26708 4377 26740 4411
rect 26774 4377 26809 4411
rect 26843 4377 26878 4411
rect 26912 4377 26947 4411
rect 26981 4377 27016 4411
rect 27050 4377 27085 4411
rect 27119 4377 27154 4411
rect 27188 4377 27223 4411
rect 27257 4377 27292 4411
rect 27326 4377 27361 4411
rect 27395 4377 27430 4411
rect 27464 4377 27499 4411
rect 27533 4377 27568 4411
rect 26708 4343 27568 4377
rect 26708 4309 26740 4343
rect 26774 4309 26809 4343
rect 26843 4309 26878 4343
rect 26912 4309 26947 4343
rect 26981 4309 27016 4343
rect 27050 4309 27085 4343
rect 27119 4309 27154 4343
rect 27188 4309 27223 4343
rect 27257 4309 27292 4343
rect 27326 4309 27361 4343
rect 27395 4309 27430 4343
rect 27464 4309 27499 4343
rect 27533 4309 27568 4343
rect 26708 4275 27568 4309
rect 26708 4241 26740 4275
rect 26774 4241 26809 4275
rect 26843 4241 26878 4275
rect 26912 4241 26947 4275
rect 26981 4241 27016 4275
rect 27050 4241 27085 4275
rect 27119 4241 27154 4275
rect 27188 4241 27223 4275
rect 27257 4241 27292 4275
rect 27326 4241 27361 4275
rect 27395 4241 27430 4275
rect 27464 4241 27499 4275
rect 27533 4241 27568 4275
rect 28690 5465 28777 5499
rect 28811 5465 28847 5499
rect 28881 5465 28917 5499
rect 28951 5465 28987 5499
rect 29021 5465 29057 5499
rect 29091 5465 29127 5499
rect 29161 5465 29197 5499
rect 29231 5465 29267 5499
rect 29301 5465 29337 5499
rect 29371 5465 29407 5499
rect 29441 5465 29477 5499
rect 29511 5465 29547 5499
rect 29581 5465 29617 5499
rect 29651 5465 29687 5499
rect 29721 5465 29757 5499
rect 29791 5465 29827 5499
rect 29861 5465 29896 5499
rect 29930 5465 29965 5499
rect 29999 5465 30034 5499
rect 30068 5465 30103 5499
rect 30137 5465 30172 5499
rect 30206 5465 30230 5499
rect 28690 5431 30230 5465
rect 28690 5397 28777 5431
rect 28811 5397 28847 5431
rect 28881 5397 28917 5431
rect 28951 5397 28987 5431
rect 29021 5397 29057 5431
rect 29091 5397 29127 5431
rect 29161 5397 29197 5431
rect 29231 5397 29267 5431
rect 29301 5397 29337 5431
rect 29371 5397 29407 5431
rect 29441 5397 29477 5431
rect 29511 5397 29547 5431
rect 29581 5397 29617 5431
rect 29651 5397 29687 5431
rect 29721 5397 29757 5431
rect 29791 5397 29827 5431
rect 29861 5397 29896 5431
rect 29930 5397 29965 5431
rect 29999 5397 30034 5431
rect 30068 5397 30103 5431
rect 30137 5397 30172 5431
rect 30206 5397 30230 5431
rect 28690 5363 30230 5397
rect 28690 5329 28777 5363
rect 28811 5329 28847 5363
rect 28881 5329 28917 5363
rect 28951 5329 28987 5363
rect 29021 5329 29057 5363
rect 29091 5329 29127 5363
rect 29161 5329 29197 5363
rect 29231 5329 29267 5363
rect 29301 5329 29337 5363
rect 29371 5329 29407 5363
rect 29441 5329 29477 5363
rect 29511 5329 29547 5363
rect 29581 5329 29617 5363
rect 29651 5329 29687 5363
rect 29721 5329 29757 5363
rect 29791 5329 29827 5363
rect 29861 5329 29896 5363
rect 29930 5329 29965 5363
rect 29999 5329 30034 5363
rect 30068 5329 30103 5363
rect 30137 5329 30172 5363
rect 30206 5329 30230 5363
rect 28690 5295 30230 5329
rect 28690 5261 28777 5295
rect 28811 5261 28847 5295
rect 28881 5261 28917 5295
rect 28951 5261 28987 5295
rect 29021 5261 29057 5295
rect 29091 5261 29127 5295
rect 29161 5261 29197 5295
rect 29231 5261 29267 5295
rect 29301 5261 29337 5295
rect 29371 5261 29407 5295
rect 29441 5261 29477 5295
rect 29511 5261 29547 5295
rect 29581 5261 29617 5295
rect 29651 5261 29687 5295
rect 29721 5261 29757 5295
rect 29791 5261 29827 5295
rect 29861 5261 29896 5295
rect 29930 5261 29965 5295
rect 29999 5261 30034 5295
rect 30068 5261 30103 5295
rect 30137 5261 30172 5295
rect 30206 5261 30230 5295
rect 28690 5227 30230 5261
rect 28690 5193 28777 5227
rect 28811 5193 28847 5227
rect 28881 5193 28917 5227
rect 28951 5193 28987 5227
rect 29021 5193 29057 5227
rect 29091 5193 29127 5227
rect 29161 5193 29197 5227
rect 29231 5193 29267 5227
rect 29301 5193 29337 5227
rect 29371 5193 29407 5227
rect 29441 5193 29477 5227
rect 29511 5193 29547 5227
rect 29581 5193 29617 5227
rect 29651 5193 29687 5227
rect 29721 5193 29757 5227
rect 29791 5193 29827 5227
rect 29861 5193 29896 5227
rect 29930 5193 29965 5227
rect 29999 5193 30034 5227
rect 30068 5193 30103 5227
rect 30137 5193 30172 5227
rect 30206 5193 30230 5227
rect 28690 5159 30230 5193
rect 28690 5125 28777 5159
rect 28811 5125 28847 5159
rect 28881 5125 28917 5159
rect 28951 5125 28987 5159
rect 29021 5125 29057 5159
rect 29091 5125 29127 5159
rect 29161 5125 29197 5159
rect 29231 5125 29267 5159
rect 29301 5125 29337 5159
rect 29371 5125 29407 5159
rect 29441 5125 29477 5159
rect 29511 5125 29547 5159
rect 29581 5125 29617 5159
rect 29651 5125 29687 5159
rect 29721 5125 29757 5159
rect 29791 5125 29827 5159
rect 29861 5125 29896 5159
rect 29930 5125 29965 5159
rect 29999 5125 30034 5159
rect 30068 5125 30103 5159
rect 30137 5125 30172 5159
rect 30206 5125 30230 5159
rect 28690 5091 30230 5125
rect 28690 5057 28777 5091
rect 28811 5057 28847 5091
rect 28881 5057 28917 5091
rect 28951 5057 28987 5091
rect 29021 5057 29057 5091
rect 29091 5057 29127 5091
rect 29161 5057 29197 5091
rect 29231 5057 29267 5091
rect 29301 5057 29337 5091
rect 29371 5057 29407 5091
rect 29441 5057 29477 5091
rect 29511 5057 29547 5091
rect 29581 5057 29617 5091
rect 29651 5057 29687 5091
rect 29721 5057 29757 5091
rect 29791 5057 29827 5091
rect 29861 5057 29896 5091
rect 29930 5057 29965 5091
rect 29999 5057 30034 5091
rect 30068 5057 30103 5091
rect 30137 5057 30172 5091
rect 30206 5057 30230 5091
rect 28690 5023 30230 5057
rect 28690 4989 28777 5023
rect 28811 4989 28847 5023
rect 28881 4989 28917 5023
rect 28951 4989 28987 5023
rect 29021 4989 29057 5023
rect 29091 4989 29127 5023
rect 29161 4989 29197 5023
rect 29231 4989 29267 5023
rect 29301 4989 29337 5023
rect 29371 4989 29407 5023
rect 29441 4989 29477 5023
rect 29511 4989 29547 5023
rect 29581 4989 29617 5023
rect 29651 4989 29687 5023
rect 29721 4989 29757 5023
rect 29791 4989 29827 5023
rect 29861 4989 29896 5023
rect 29930 4989 29965 5023
rect 29999 4989 30034 5023
rect 30068 4989 30103 5023
rect 30137 4989 30172 5023
rect 30206 4989 30230 5023
rect 28690 4955 30230 4989
rect 28690 4921 28777 4955
rect 28811 4921 28847 4955
rect 28881 4921 28917 4955
rect 28951 4921 28987 4955
rect 29021 4921 29057 4955
rect 29091 4921 29127 4955
rect 29161 4921 29197 4955
rect 29231 4921 29267 4955
rect 29301 4921 29337 4955
rect 29371 4921 29407 4955
rect 29441 4921 29477 4955
rect 29511 4921 29547 4955
rect 29581 4921 29617 4955
rect 29651 4921 29687 4955
rect 29721 4921 29757 4955
rect 29791 4921 29827 4955
rect 29861 4921 29896 4955
rect 29930 4921 29965 4955
rect 29999 4921 30034 4955
rect 30068 4921 30103 4955
rect 30137 4921 30172 4955
rect 30206 4921 30230 4955
rect 28690 4887 30230 4921
rect 28690 4853 28777 4887
rect 28811 4853 28847 4887
rect 28881 4853 28917 4887
rect 28951 4853 28987 4887
rect 29021 4853 29057 4887
rect 29091 4853 29127 4887
rect 29161 4853 29197 4887
rect 29231 4853 29267 4887
rect 29301 4853 29337 4887
rect 29371 4853 29407 4887
rect 29441 4853 29477 4887
rect 29511 4853 29547 4887
rect 29581 4853 29617 4887
rect 29651 4853 29687 4887
rect 29721 4853 29757 4887
rect 29791 4853 29827 4887
rect 29861 4853 29896 4887
rect 29930 4853 29965 4887
rect 29999 4853 30034 4887
rect 30068 4853 30103 4887
rect 30137 4853 30172 4887
rect 30206 4853 30230 4887
rect 28690 4819 30230 4853
rect 28690 4785 28777 4819
rect 28811 4785 28847 4819
rect 28881 4785 28917 4819
rect 28951 4785 28987 4819
rect 29021 4785 29057 4819
rect 29091 4785 29127 4819
rect 29161 4785 29197 4819
rect 29231 4785 29267 4819
rect 29301 4785 29337 4819
rect 29371 4785 29407 4819
rect 29441 4785 29477 4819
rect 29511 4785 29547 4819
rect 29581 4785 29617 4819
rect 29651 4785 29687 4819
rect 29721 4785 29757 4819
rect 29791 4785 29827 4819
rect 29861 4785 29896 4819
rect 29930 4785 29965 4819
rect 29999 4785 30034 4819
rect 30068 4785 30103 4819
rect 30137 4785 30172 4819
rect 30206 4785 30230 4819
rect 28690 4751 30230 4785
rect 28690 4717 28777 4751
rect 28811 4717 28847 4751
rect 28881 4717 28917 4751
rect 28951 4717 28987 4751
rect 29021 4717 29057 4751
rect 29091 4717 29127 4751
rect 29161 4717 29197 4751
rect 29231 4717 29267 4751
rect 29301 4717 29337 4751
rect 29371 4717 29407 4751
rect 29441 4717 29477 4751
rect 29511 4717 29547 4751
rect 29581 4717 29617 4751
rect 29651 4717 29687 4751
rect 29721 4717 29757 4751
rect 29791 4717 29827 4751
rect 29861 4717 29896 4751
rect 29930 4717 29965 4751
rect 29999 4717 30034 4751
rect 30068 4717 30103 4751
rect 30137 4717 30172 4751
rect 30206 4717 30230 4751
rect 28690 4241 28714 4717
rect 26708 4169 28714 4241
rect 20165 4107 20482 4141
rect 20165 4073 20167 4107
rect 20201 4073 20247 4107
rect 20281 4073 20327 4107
rect 20361 4073 20407 4107
rect 20441 4073 20482 4107
rect 20165 4039 20482 4073
rect 20165 4005 20167 4039
rect 20201 4005 20247 4039
rect 20281 4005 20327 4039
rect 20361 4005 20407 4039
rect 20441 4005 20482 4039
rect 20165 3971 20482 4005
rect 20165 3937 20167 3971
rect 20201 3937 20247 3971
rect 20281 3937 20327 3971
rect 20361 3937 20407 3971
rect 20441 3937 20482 3971
rect 20165 3903 20482 3937
rect 20165 3869 20167 3903
rect 20201 3869 20247 3903
rect 20281 3869 20327 3903
rect 20361 3869 20407 3903
rect 20441 3869 20482 3903
rect 20165 3835 20482 3869
rect 20165 3801 20167 3835
rect 20201 3801 20247 3835
rect 20281 3801 20327 3835
rect 20361 3801 20407 3835
rect 20441 3801 20482 3835
rect 20165 3767 20482 3801
rect 20165 3733 20167 3767
rect 20201 3733 20247 3767
rect 20281 3733 20327 3767
rect 20361 3733 20407 3767
rect 20441 3733 20482 3767
rect 20165 3699 20482 3733
rect 20165 3665 20167 3699
rect 20201 3665 20247 3699
rect 20281 3665 20327 3699
rect 20361 3665 20407 3699
rect 20441 3665 20482 3699
rect 20165 3631 20482 3665
rect 20165 3597 20167 3631
rect 20201 3597 20247 3631
rect 20281 3597 20327 3631
rect 20361 3597 20407 3631
rect 20441 3597 20482 3631
rect 20165 3563 20482 3597
rect 20165 3529 20167 3563
rect 20201 3529 20247 3563
rect 20281 3529 20327 3563
rect 20361 3529 20407 3563
rect 20441 3529 20482 3563
rect 20165 3495 20482 3529
rect 20165 3461 20167 3495
rect 20201 3461 20247 3495
rect 20281 3461 20327 3495
rect 20361 3461 20407 3495
rect 20441 3461 20482 3495
rect 20165 3427 20482 3461
rect 20165 3393 20167 3427
rect 20201 3393 20247 3427
rect 20281 3393 20327 3427
rect 20361 3393 20407 3427
rect 20441 3393 20482 3427
rect 20165 3359 20482 3393
rect 20165 3325 20167 3359
rect 20201 3325 20247 3359
rect 20281 3325 20327 3359
rect 20361 3325 20407 3359
rect 20441 3325 20482 3359
rect 20165 3291 20482 3325
rect 20165 3257 20167 3291
rect 20201 3257 20247 3291
rect 20281 3257 20327 3291
rect 20361 3257 20407 3291
rect 20441 3257 20482 3291
rect 20165 3223 20482 3257
rect 20165 3189 20167 3223
rect 20201 3189 20247 3223
rect 20281 3189 20327 3223
rect 20361 3189 20407 3223
rect 20441 3189 20482 3223
rect 20165 3155 20482 3189
rect 20165 3121 20167 3155
rect 20201 3121 20247 3155
rect 20281 3121 20327 3155
rect 20361 3121 20407 3155
rect 20441 3121 20482 3155
rect 20165 3087 20482 3121
rect 20165 3053 20167 3087
rect 20201 3053 20247 3087
rect 20281 3053 20327 3087
rect 20361 3053 20407 3087
rect 20441 3053 20482 3087
rect 20165 3019 20482 3053
rect 20165 2985 20167 3019
rect 20201 2985 20247 3019
rect 20281 2985 20327 3019
rect 20361 2985 20407 3019
rect 20441 2985 20482 3019
rect 20165 2951 20482 2985
rect 20165 2917 20167 2951
rect 20201 2917 20247 2951
rect 20281 2917 20327 2951
rect 20361 2917 20407 2951
rect 20441 2917 20482 2951
rect 20165 2883 20482 2917
rect 20165 2849 20167 2883
rect 20201 2849 20247 2883
rect 20281 2849 20327 2883
rect 20361 2849 20407 2883
rect 20441 2849 20482 2883
rect 20165 2815 20482 2849
rect 20165 2781 20167 2815
rect 20201 2781 20247 2815
rect 20281 2781 20327 2815
rect 20361 2781 20407 2815
rect 20441 2781 20482 2815
rect 20165 2747 20482 2781
rect 20165 2713 20167 2747
rect 20201 2713 20247 2747
rect 20281 2713 20327 2747
rect 20361 2713 20407 2747
rect 20441 2713 20482 2747
rect 20165 2678 20482 2713
rect 20165 2644 20167 2678
rect 20201 2644 20247 2678
rect 20281 2644 20327 2678
rect 20361 2644 20407 2678
rect 20441 2644 20482 2678
rect 20165 2637 20482 2644
rect 22523 3049 22789 3073
rect 22523 3015 22559 3049
rect 22593 3015 22657 3049
rect 22691 3015 22755 3049
rect 22523 2977 22789 3015
rect 22523 2943 22559 2977
rect 22593 2943 22657 2977
rect 22691 2943 22755 2977
rect 22523 2904 22789 2943
rect 22523 2870 22559 2904
rect 22593 2870 22657 2904
rect 22691 2870 22755 2904
rect 22523 2831 22789 2870
rect 22523 2797 22559 2831
rect 22593 2797 22657 2831
rect 22691 2797 22755 2831
rect 22523 2758 22789 2797
rect 22523 2724 22559 2758
rect 22593 2724 22657 2758
rect 22691 2724 22755 2758
rect 22523 2685 22789 2724
rect 22523 2651 22559 2685
rect 22593 2651 22657 2685
rect 22691 2651 22755 2685
rect 22523 2637 22789 2651
rect 20165 2612 22789 2637
rect 20165 2585 22559 2612
rect 18148 2551 18172 2585
rect 18206 2551 18241 2585
rect 18275 2551 18310 2585
rect 18344 2551 18379 2585
rect 18413 2551 18448 2585
rect 18482 2551 18517 2585
rect 18551 2551 18586 2585
rect 18620 2551 18655 2585
rect 18689 2551 18724 2585
rect 18758 2551 18793 2585
rect 18827 2551 18861 2585
rect 18895 2551 18929 2585
rect 18963 2551 18997 2585
rect 19031 2551 19065 2585
rect 19099 2551 19133 2585
rect 19167 2551 19201 2585
rect 19235 2551 19269 2585
rect 19303 2551 19337 2585
rect 19371 2551 19405 2585
rect 19439 2551 19473 2585
rect 19507 2551 19541 2585
rect 19575 2551 19609 2585
rect 19643 2551 19677 2585
rect 19711 2551 19745 2585
rect 19779 2551 19813 2585
rect 19847 2551 19881 2585
rect 19915 2551 19949 2585
rect 19983 2551 20017 2585
rect 20051 2551 20085 2585
rect 20119 2551 20153 2585
rect 20187 2551 20221 2585
rect 20255 2551 20289 2585
rect 20323 2551 20357 2585
rect 20391 2551 20425 2585
rect 20459 2551 20493 2585
rect 20527 2551 20561 2585
rect 20595 2551 20629 2585
rect 20663 2551 20697 2585
rect 20731 2551 20765 2585
rect 20799 2551 20833 2585
rect 20867 2551 20901 2585
rect 20935 2551 20969 2585
rect 21003 2551 21037 2585
rect 21071 2551 21105 2585
rect 21139 2551 21173 2585
rect 21207 2551 21241 2585
rect 21275 2551 21309 2585
rect 21343 2551 21377 2585
rect 21411 2551 21445 2585
rect 21479 2551 21513 2585
rect 21547 2551 21581 2585
rect 21615 2551 21649 2585
rect 21683 2551 21717 2585
rect 21751 2551 21785 2585
rect 21819 2551 21853 2585
rect 21887 2551 21921 2585
rect 21955 2551 21989 2585
rect 22023 2551 22057 2585
rect 22091 2551 22125 2585
rect 22159 2551 22193 2585
rect 22227 2551 22261 2585
rect 22295 2551 22329 2585
rect 22363 2551 22397 2585
rect 22431 2551 22465 2585
rect 22499 2578 22559 2585
rect 22593 2578 22657 2612
rect 22691 2578 22755 2612
rect 22499 2551 22789 2578
rect 18148 2539 22789 2551
rect 18148 2515 22559 2539
rect 16523 2481 16579 2515
rect 16613 2481 16650 2515
rect 16684 2481 16721 2515
rect 16755 2481 16792 2515
rect 16826 2481 16863 2515
rect 16897 2481 16933 2515
rect 16967 2481 17003 2515
rect 17037 2481 17073 2515
rect 17107 2481 17143 2515
rect 17177 2481 17213 2515
rect 17247 2481 17283 2515
rect 17317 2481 17353 2515
rect 17387 2481 17423 2515
rect 17457 2481 17493 2515
rect 17527 2481 17563 2515
rect 17597 2481 17633 2515
rect 17667 2481 17703 2515
rect 17737 2481 17773 2515
rect 17807 2481 17843 2515
rect 17877 2481 17913 2515
rect 17947 2481 17983 2515
rect 18017 2481 18053 2515
rect 18087 2481 18172 2515
rect 18206 2481 18241 2515
rect 18275 2481 18310 2515
rect 18344 2481 18379 2515
rect 18413 2481 18448 2515
rect 18482 2481 18517 2515
rect 18551 2481 18586 2515
rect 18620 2481 18655 2515
rect 18689 2481 18724 2515
rect 18758 2481 18793 2515
rect 18827 2481 18861 2515
rect 18895 2481 18929 2515
rect 18963 2481 18997 2515
rect 19031 2481 19065 2515
rect 19099 2481 19133 2515
rect 19167 2481 19201 2515
rect 19235 2481 19269 2515
rect 19303 2481 19337 2515
rect 19371 2481 19405 2515
rect 19439 2481 19473 2515
rect 19507 2481 19541 2515
rect 19575 2481 19609 2515
rect 19643 2481 19677 2515
rect 19711 2481 19745 2515
rect 19779 2481 19813 2515
rect 19847 2481 19881 2515
rect 19915 2481 19949 2515
rect 19983 2481 20017 2515
rect 20051 2481 20085 2515
rect 20119 2481 20153 2515
rect 20187 2481 20221 2515
rect 20255 2481 20289 2515
rect 20323 2481 20357 2515
rect 20391 2481 20425 2515
rect 20459 2481 20493 2515
rect 20527 2481 20561 2515
rect 20595 2481 20629 2515
rect 20663 2481 20697 2515
rect 20731 2481 20765 2515
rect 20799 2481 20833 2515
rect 20867 2481 20901 2515
rect 20935 2481 20969 2515
rect 21003 2481 21037 2515
rect 21071 2481 21105 2515
rect 21139 2481 21173 2515
rect 21207 2481 21241 2515
rect 21275 2481 21309 2515
rect 21343 2481 21377 2515
rect 21411 2481 21445 2515
rect 21479 2481 21513 2515
rect 21547 2481 21581 2515
rect 21615 2481 21649 2515
rect 21683 2481 21717 2515
rect 21751 2481 21785 2515
rect 21819 2481 21853 2515
rect 21887 2481 21921 2515
rect 21955 2481 21989 2515
rect 22023 2481 22057 2515
rect 22091 2481 22125 2515
rect 22159 2481 22193 2515
rect 22227 2481 22261 2515
rect 22295 2481 22329 2515
rect 22363 2481 22397 2515
rect 22431 2481 22465 2515
rect 22499 2505 22559 2515
rect 22593 2505 22657 2539
rect 22691 2505 22755 2539
rect 22499 2481 22789 2505
rect 16523 2446 22789 2481
rect 22275 2403 22789 2446
rect 22275 2369 22347 2403
rect 22381 2369 22415 2403
rect 22449 2369 22483 2403
rect 22517 2369 22551 2403
rect 22585 2369 22619 2403
rect 22653 2369 22687 2403
rect 22721 2369 22755 2403
rect 22275 2328 22789 2369
rect 22275 2294 22347 2328
rect 22381 2294 22415 2328
rect 22449 2294 22483 2328
rect 22517 2294 22551 2328
rect 22585 2294 22619 2328
rect 22653 2294 22687 2328
rect 22721 2294 22755 2328
rect 22275 2252 22789 2294
rect 22275 2218 22347 2252
rect 22381 2218 22415 2252
rect 22449 2218 22483 2252
rect 22517 2218 22551 2252
rect 22585 2218 22619 2252
rect 22653 2218 22687 2252
rect 22721 2218 22755 2252
rect 22275 2176 22789 2218
rect 22275 2142 22347 2176
rect 22381 2142 22415 2176
rect 22449 2142 22483 2176
rect 22517 2142 22551 2176
rect 22585 2142 22619 2176
rect 22653 2142 22687 2176
rect 22721 2142 22755 2176
rect 22275 2100 22789 2142
rect 22275 2066 22347 2100
rect 22381 2066 22415 2100
rect 22449 2066 22483 2100
rect 22517 2066 22551 2100
rect 22585 2066 22619 2100
rect 22653 2066 22687 2100
rect 22721 2066 22755 2100
rect 22275 2024 22789 2066
rect 22275 1990 22347 2024
rect 22381 1990 22415 2024
rect 22449 1990 22483 2024
rect 22517 1990 22551 2024
rect 22585 1990 22619 2024
rect 22653 1990 22687 2024
rect 22721 1990 22755 2024
rect 22275 1948 22789 1990
rect 22275 1914 22347 1948
rect 22381 1914 22415 1948
rect 22449 1914 22483 1948
rect 22517 1914 22551 1948
rect 22585 1914 22619 1948
rect 22653 1914 22687 1948
rect 22721 1914 22755 1948
rect 22275 1872 22789 1914
rect 22275 1838 22347 1872
rect 22381 1838 22415 1872
rect 22449 1838 22483 1872
rect 22517 1838 22551 1872
rect 22585 1838 22619 1872
rect 22653 1838 22687 1872
rect 22721 1838 22755 1872
rect 22275 1796 22789 1838
rect 22275 1762 22347 1796
rect 22381 1762 22415 1796
rect 22449 1762 22483 1796
rect 22517 1762 22551 1796
rect 22585 1762 22619 1796
rect 22653 1762 22687 1796
rect 22721 1762 22755 1796
rect 22275 1738 22789 1762
rect 26722 2273 28392 2348
rect 26722 2239 26787 2273
rect 26821 2239 26858 2273
rect 26892 2239 26929 2273
rect 26963 2239 27000 2273
rect 27034 2239 27071 2273
rect 27105 2239 27142 2273
rect 27176 2239 27213 2273
rect 27247 2239 27284 2273
rect 27318 2239 27354 2273
rect 27388 2239 27424 2273
rect 27458 2239 27494 2273
rect 27528 2239 27564 2273
rect 27598 2239 27634 2273
rect 27668 2239 27704 2273
rect 27738 2239 27774 2273
rect 27808 2239 27844 2273
rect 27878 2239 27914 2273
rect 27948 2239 27984 2273
rect 28018 2239 28054 2273
rect 28088 2239 28124 2273
rect 28158 2239 28194 2273
rect 28228 2239 28264 2273
rect 28298 2239 28334 2273
rect 28368 2239 28392 2273
rect 26722 2205 28392 2239
rect 26722 2171 26787 2205
rect 26821 2171 26858 2205
rect 26892 2171 26929 2205
rect 26963 2171 27000 2205
rect 27034 2171 27071 2205
rect 27105 2171 27142 2205
rect 27176 2171 27213 2205
rect 27247 2171 27284 2205
rect 27318 2171 27354 2205
rect 27388 2171 27424 2205
rect 27458 2171 27494 2205
rect 27528 2171 27564 2205
rect 27598 2171 27634 2205
rect 27668 2171 27704 2205
rect 27738 2171 27774 2205
rect 27808 2171 27844 2205
rect 27878 2171 27914 2205
rect 27948 2171 27984 2205
rect 28018 2171 28054 2205
rect 28088 2171 28124 2205
rect 28158 2171 28194 2205
rect 28228 2171 28264 2205
rect 28298 2171 28334 2205
rect 28368 2171 28392 2205
rect 26722 2137 28392 2171
rect 26722 2103 26787 2137
rect 26821 2103 26858 2137
rect 26892 2103 26929 2137
rect 26963 2103 27000 2137
rect 27034 2103 27071 2137
rect 27105 2103 27142 2137
rect 27176 2103 27213 2137
rect 27247 2103 27284 2137
rect 27318 2103 27354 2137
rect 27388 2103 27424 2137
rect 27458 2103 27494 2137
rect 27528 2103 27564 2137
rect 27598 2103 27634 2137
rect 27668 2103 27704 2137
rect 27738 2103 27774 2137
rect 27808 2103 27844 2137
rect 27878 2103 27914 2137
rect 27948 2103 27984 2137
rect 28018 2103 28054 2137
rect 28088 2103 28124 2137
rect 28158 2103 28194 2137
rect 28228 2103 28264 2137
rect 28298 2103 28334 2137
rect 28368 2103 28392 2137
rect 26722 2069 28392 2103
rect 26722 2035 26787 2069
rect 26821 2035 26858 2069
rect 26892 2035 26929 2069
rect 26963 2035 27000 2069
rect 27034 2035 27071 2069
rect 27105 2035 27142 2069
rect 27176 2035 27213 2069
rect 27247 2035 27284 2069
rect 27318 2035 27354 2069
rect 27388 2035 27424 2069
rect 27458 2035 27494 2069
rect 27528 2035 27564 2069
rect 27598 2035 27634 2069
rect 27668 2035 27704 2069
rect 27738 2035 27774 2069
rect 27808 2035 27844 2069
rect 27878 2035 27914 2069
rect 27948 2035 27984 2069
rect 28018 2035 28054 2069
rect 28088 2035 28124 2069
rect 28158 2035 28194 2069
rect 28228 2035 28264 2069
rect 28298 2035 28334 2069
rect 28368 2035 28392 2069
rect 26722 2001 28392 2035
rect 26722 1967 26787 2001
rect 26821 1967 26858 2001
rect 26892 1967 26929 2001
rect 26963 1967 27000 2001
rect 27034 1967 27071 2001
rect 27105 1967 27142 2001
rect 27176 1967 27213 2001
rect 27247 1967 27284 2001
rect 27318 1967 27354 2001
rect 27388 1967 27424 2001
rect 27458 1967 27494 2001
rect 27528 1967 27564 2001
rect 27598 1967 27634 2001
rect 27668 1967 27704 2001
rect 27738 1967 27774 2001
rect 27808 1967 27844 2001
rect 27878 1967 27914 2001
rect 27948 1967 27984 2001
rect 28018 1967 28054 2001
rect 28088 1967 28124 2001
rect 28158 1967 28194 2001
rect 28228 1967 28264 2001
rect 28298 1967 28334 2001
rect 28368 1967 28392 2001
rect 26722 1933 28392 1967
rect 26722 1899 26787 1933
rect 26821 1899 26858 1933
rect 26892 1899 26929 1933
rect 26963 1899 27000 1933
rect 27034 1899 27071 1933
rect 27105 1899 27142 1933
rect 27176 1899 27213 1933
rect 27247 1899 27284 1933
rect 27318 1899 27354 1933
rect 27388 1899 27424 1933
rect 27458 1899 27494 1933
rect 27528 1899 27564 1933
rect 27598 1899 27634 1933
rect 27668 1899 27704 1933
rect 27738 1899 27774 1933
rect 27808 1899 27844 1933
rect 27878 1899 27914 1933
rect 27948 1899 27984 1933
rect 28018 1899 28054 1933
rect 28088 1899 28124 1933
rect 28158 1899 28194 1933
rect 28228 1899 28264 1933
rect 28298 1899 28334 1933
rect 28368 1899 28392 1933
rect 26722 1865 28392 1899
rect 26722 1831 26787 1865
rect 26821 1831 26858 1865
rect 26892 1831 26929 1865
rect 26963 1831 27000 1865
rect 27034 1831 27071 1865
rect 27105 1831 27142 1865
rect 27176 1831 27213 1865
rect 27247 1831 27284 1865
rect 27318 1831 27354 1865
rect 27388 1831 27424 1865
rect 27458 1831 27494 1865
rect 27528 1831 27564 1865
rect 27598 1831 27634 1865
rect 27668 1831 27704 1865
rect 27738 1831 27774 1865
rect 27808 1831 27844 1865
rect 27878 1831 27914 1865
rect 27948 1831 27984 1865
rect 28018 1831 28054 1865
rect 28088 1831 28124 1865
rect 28158 1831 28194 1865
rect 28228 1831 28264 1865
rect 28298 1831 28334 1865
rect 28368 1831 28392 1865
rect 26722 1797 28392 1831
rect 26722 1763 26787 1797
rect 26821 1763 26858 1797
rect 26892 1763 26929 1797
rect 26963 1763 27000 1797
rect 27034 1763 27071 1797
rect 27105 1763 27142 1797
rect 27176 1763 27213 1797
rect 27247 1763 27284 1797
rect 27318 1763 27354 1797
rect 27388 1763 27424 1797
rect 27458 1763 27494 1797
rect 27528 1763 27564 1797
rect 27598 1763 27634 1797
rect 27668 1763 27704 1797
rect 27738 1763 27774 1797
rect 27808 1763 27844 1797
rect 27878 1763 27914 1797
rect 27948 1763 27984 1797
rect 28018 1763 28054 1797
rect 28088 1763 28124 1797
rect 28158 1763 28194 1797
rect 28228 1763 28264 1797
rect 28298 1763 28334 1797
rect 28368 1763 28392 1797
rect 26722 1729 28392 1763
rect 26722 1695 26787 1729
rect 26821 1695 26858 1729
rect 26892 1695 26929 1729
rect 26963 1695 27000 1729
rect 27034 1695 27071 1729
rect 27105 1695 27142 1729
rect 27176 1695 27213 1729
rect 27247 1695 27284 1729
rect 27318 1695 27354 1729
rect 27388 1695 27424 1729
rect 27458 1695 27494 1729
rect 27528 1695 27564 1729
rect 27598 1695 27634 1729
rect 27668 1695 27704 1729
rect 27738 1695 27774 1729
rect 27808 1695 27844 1729
rect 27878 1695 27914 1729
rect 27948 1695 27984 1729
rect 28018 1695 28054 1729
rect 28088 1695 28124 1729
rect 28158 1695 28194 1729
rect 28228 1695 28264 1729
rect 28298 1695 28334 1729
rect 28368 1695 28392 1729
rect 26722 1643 26979 1695
rect 26722 1609 26753 1643
rect 26787 1609 26849 1643
rect 26883 1609 26945 1643
rect 26722 1571 26979 1609
rect 26722 1537 26753 1571
rect 26787 1537 26849 1571
rect 26883 1537 26945 1571
rect 26722 1499 26979 1537
rect 26722 1465 26753 1499
rect 26787 1465 26849 1499
rect 26883 1465 26945 1499
rect 26722 1426 26979 1465
rect 26722 1392 26753 1426
rect 26787 1392 26849 1426
rect 26883 1392 26945 1426
rect 26722 1353 26979 1392
rect 26722 1319 26753 1353
rect 26787 1319 26849 1353
rect 26883 1319 26945 1353
rect 26722 1280 26979 1319
rect 26722 1246 26753 1280
rect 26787 1246 26849 1280
rect 26883 1246 26945 1280
rect 26722 1207 26979 1246
rect 26722 1173 26753 1207
rect 26787 1173 26849 1207
rect 26883 1173 26945 1207
rect 26722 1134 26979 1173
rect 26722 1100 26753 1134
rect 26787 1100 26849 1134
rect 26883 1100 26945 1134
rect 26722 1061 26979 1100
rect 26722 1027 26753 1061
rect 26787 1027 26849 1061
rect 26883 1027 26945 1061
rect 26722 988 26979 1027
rect 26722 954 26753 988
rect 26787 954 26849 988
rect 26883 954 26945 988
rect 26722 915 26979 954
rect 26722 881 26753 915
rect 26787 881 26849 915
rect 26883 881 26945 915
rect 26722 860 26979 881
<< mvnsubdiff >>
rect 17811 23432 17913 23456
rect 17811 22479 17913 22514
rect 17845 22445 17879 22479
rect 17811 22410 17913 22445
rect 17845 22376 17879 22410
rect 17811 22341 17913 22376
rect 17845 22307 17879 22341
rect 17811 22272 17913 22307
rect 17845 22238 17879 22272
rect 17811 22203 17913 22238
rect 17845 22169 17879 22203
rect 17811 22134 17913 22169
rect 17845 22100 17879 22134
rect 17811 22065 17913 22100
rect 17845 22031 17879 22065
rect 17811 21996 17913 22031
rect 17845 21962 17879 21996
rect 17811 21927 17913 21962
rect 17845 21893 17879 21927
rect 17811 21858 17913 21893
rect 17845 21824 17879 21858
rect 17811 21789 17913 21824
rect 17845 21755 17879 21789
rect 17811 21720 17913 21755
rect 17845 21686 17879 21720
rect 17811 21651 17913 21686
rect 17845 21617 17879 21651
rect 17811 21582 17913 21617
rect 17845 21548 17879 21582
rect 17811 21513 17913 21548
rect 17845 21479 17879 21513
rect 17811 21444 17913 21479
rect 17845 21410 17879 21444
rect 17811 21375 17913 21410
rect 17845 21341 17879 21375
rect 17811 21306 17913 21341
rect 17845 21272 17879 21306
rect 17811 21237 17913 21272
rect 17845 21203 17879 21237
rect 17811 21168 17913 21203
rect 17845 21134 17879 21168
rect 17811 21099 17913 21134
rect 17845 21065 17879 21099
rect 17811 21030 17913 21065
rect 17845 20996 17879 21030
rect 17811 20961 17913 20996
rect 17845 20927 17879 20961
rect 17811 20892 17913 20927
rect 17845 20858 17879 20892
rect 17811 20823 17913 20858
rect 17845 20789 17879 20823
rect 17811 20754 17913 20789
rect 17845 20720 17879 20754
rect 17811 20685 17913 20720
rect 17845 20651 17879 20685
rect 17811 20616 17913 20651
rect 17845 20582 17879 20616
rect 17811 20547 17913 20582
rect 17845 20513 17879 20547
rect 17811 20478 17913 20513
rect 17845 20444 17879 20478
rect 17811 20409 17913 20444
rect 17845 20375 17879 20409
rect 17811 20340 17913 20375
rect 17845 20306 17879 20340
rect 17811 20282 17913 20306
<< psubdiffcont >>
rect 28665 7906 28699 7940
rect 28734 7906 28768 7940
rect 28803 7906 28837 7940
rect 28872 7906 28906 7940
rect 28941 7906 28975 7940
rect 29010 7906 29044 7940
rect 29079 7906 29113 7940
rect 29148 7906 29182 7940
rect 29217 7906 29251 7940
rect 29286 7906 29320 7940
rect 29355 7906 29389 7940
rect 29424 7906 29458 7940
rect 29493 7906 29527 7940
rect 29562 7906 29596 7940
rect 29631 7906 29665 7940
rect 29700 7906 29734 7940
rect 29769 7906 29803 7940
rect 29838 7906 29872 7940
rect 29907 7906 29941 7940
rect 29976 7906 30010 7940
rect 30045 7906 30079 7940
rect 30114 7906 30148 7940
rect 30183 7906 30217 7940
rect 30252 7906 30286 7940
rect 30321 7906 30355 7940
rect 30390 7906 30424 7940
rect 30459 7906 30493 7940
rect 30528 7906 30562 7940
rect 28665 7838 28699 7872
rect 28734 7838 28768 7872
rect 28803 7838 28837 7872
rect 28872 7838 28906 7872
rect 28941 7838 28975 7872
rect 29010 7838 29044 7872
rect 29079 7838 29113 7872
rect 29148 7838 29182 7872
rect 29217 7838 29251 7872
rect 29286 7838 29320 7872
rect 29355 7838 29389 7872
rect 29424 7838 29458 7872
rect 29493 7838 29527 7872
rect 29562 7838 29596 7872
rect 29631 7838 29665 7872
rect 29700 7838 29734 7872
rect 29769 7838 29803 7872
rect 29838 7838 29872 7872
rect 29907 7838 29941 7872
rect 29976 7838 30010 7872
rect 30045 7838 30079 7872
rect 30114 7838 30148 7872
rect 30183 7838 30217 7872
rect 30252 7838 30286 7872
rect 30321 7838 30355 7872
rect 30390 7838 30424 7872
rect 30459 7838 30493 7872
rect 30528 7838 30562 7872
rect 28665 7770 28699 7804
rect 28734 7770 28768 7804
rect 28803 7770 28837 7804
rect 28872 7770 28906 7804
rect 28941 7770 28975 7804
rect 29010 7770 29044 7804
rect 29079 7770 29113 7804
rect 29148 7770 29182 7804
rect 29217 7770 29251 7804
rect 29286 7770 29320 7804
rect 29355 7770 29389 7804
rect 29424 7770 29458 7804
rect 29493 7770 29527 7804
rect 29562 7770 29596 7804
rect 29631 7770 29665 7804
rect 29700 7770 29734 7804
rect 29769 7770 29803 7804
rect 29838 7770 29872 7804
rect 29907 7770 29941 7804
rect 29976 7770 30010 7804
rect 30045 7770 30079 7804
rect 30114 7770 30148 7804
rect 30183 7770 30217 7804
rect 30252 7770 30286 7804
rect 30321 7770 30355 7804
rect 30390 7770 30424 7804
rect 30459 7770 30493 7804
rect 30528 7770 30562 7804
rect 28665 7702 28699 7736
rect 28734 7702 28768 7736
rect 28803 7702 28837 7736
rect 28872 7702 28906 7736
rect 28941 7702 28975 7736
rect 29010 7702 29044 7736
rect 29079 7702 29113 7736
rect 29148 7702 29182 7736
rect 29217 7702 29251 7736
rect 29286 7702 29320 7736
rect 29355 7702 29389 7736
rect 29424 7702 29458 7736
rect 29493 7702 29527 7736
rect 29562 7702 29596 7736
rect 29631 7702 29665 7736
rect 29700 7702 29734 7736
rect 29769 7702 29803 7736
rect 29838 7702 29872 7736
rect 29907 7702 29941 7736
rect 29976 7702 30010 7736
rect 30045 7702 30079 7736
rect 30114 7702 30148 7736
rect 30183 7702 30217 7736
rect 30252 7702 30286 7736
rect 30321 7702 30355 7736
rect 30390 7702 30424 7736
rect 30459 7702 30493 7736
rect 30528 7702 30562 7736
rect 28665 7634 28699 7668
rect 28734 7634 28768 7668
rect 28803 7634 28837 7668
rect 28872 7634 28906 7668
rect 28941 7634 28975 7668
rect 29010 7634 29044 7668
rect 29079 7634 29113 7668
rect 29148 7634 29182 7668
rect 29217 7634 29251 7668
rect 29286 7634 29320 7668
rect 29355 7634 29389 7668
rect 29424 7634 29458 7668
rect 29493 7634 29527 7668
rect 29562 7634 29596 7668
rect 29631 7634 29665 7668
rect 29700 7634 29734 7668
rect 29769 7634 29803 7668
rect 29838 7634 29872 7668
rect 29907 7634 29941 7668
rect 29976 7634 30010 7668
rect 30045 7634 30079 7668
rect 30114 7634 30148 7668
rect 30183 7634 30217 7668
rect 30252 7634 30286 7668
rect 30321 7634 30355 7668
rect 30390 7634 30424 7668
rect 30459 7634 30493 7668
rect 30528 7634 30562 7668
rect 28665 7566 28699 7600
rect 28734 7566 28768 7600
rect 28803 7566 28837 7600
rect 28872 7566 28906 7600
rect 28941 7566 28975 7600
rect 29010 7566 29044 7600
rect 29079 7566 29113 7600
rect 29148 7566 29182 7600
rect 29217 7566 29251 7600
rect 29286 7566 29320 7600
rect 29355 7566 29389 7600
rect 29424 7566 29458 7600
rect 29493 7566 29527 7600
rect 29562 7566 29596 7600
rect 29631 7566 29665 7600
rect 29700 7566 29734 7600
rect 29769 7566 29803 7600
rect 29838 7566 29872 7600
rect 29907 7566 29941 7600
rect 29976 7566 30010 7600
rect 30045 7566 30079 7600
rect 30114 7566 30148 7600
rect 30183 7566 30217 7600
rect 30252 7566 30286 7600
rect 30321 7566 30355 7600
rect 30390 7566 30424 7600
rect 30459 7566 30493 7600
rect 30528 7566 30562 7600
rect 28665 7498 28699 7532
rect 28734 7498 28768 7532
rect 28803 7498 28837 7532
rect 28872 7498 28906 7532
rect 28941 7498 28975 7532
rect 29010 7498 29044 7532
rect 29079 7498 29113 7532
rect 29148 7498 29182 7532
rect 29217 7498 29251 7532
rect 29286 7498 29320 7532
rect 29355 7498 29389 7532
rect 29424 7498 29458 7532
rect 29493 7498 29527 7532
rect 29562 7498 29596 7532
rect 29631 7498 29665 7532
rect 29700 7498 29734 7532
rect 29769 7498 29803 7532
rect 29838 7498 29872 7532
rect 29907 7498 29941 7532
rect 29976 7498 30010 7532
rect 30045 7498 30079 7532
rect 30114 7498 30148 7532
rect 30183 7498 30217 7532
rect 30252 7498 30286 7532
rect 30321 7498 30355 7532
rect 30390 7498 30424 7532
rect 30459 7498 30493 7532
rect 30528 7498 30562 7532
rect 28665 7430 28699 7464
rect 28734 7430 28768 7464
rect 28803 7430 28837 7464
rect 28872 7430 28906 7464
rect 28941 7430 28975 7464
rect 29010 7430 29044 7464
rect 29079 7430 29113 7464
rect 29148 7430 29182 7464
rect 29217 7430 29251 7464
rect 29286 7430 29320 7464
rect 29355 7430 29389 7464
rect 29424 7430 29458 7464
rect 29493 7430 29527 7464
rect 29562 7430 29596 7464
rect 29631 7430 29665 7464
rect 29700 7430 29734 7464
rect 29769 7430 29803 7464
rect 29838 7430 29872 7464
rect 29907 7430 29941 7464
rect 29976 7430 30010 7464
rect 30045 7430 30079 7464
rect 30114 7430 30148 7464
rect 30183 7430 30217 7464
rect 30252 7430 30286 7464
rect 30321 7430 30355 7464
rect 30390 7430 30424 7464
rect 30459 7430 30493 7464
rect 30528 7430 30562 7464
rect 28665 7362 28699 7396
rect 28734 7362 28768 7396
rect 28803 7362 28837 7396
rect 28872 7362 28906 7396
rect 28941 7362 28975 7396
rect 29010 7362 29044 7396
rect 29079 7362 29113 7396
rect 29148 7362 29182 7396
rect 29217 7362 29251 7396
rect 29286 7362 29320 7396
rect 29355 7362 29389 7396
rect 29424 7362 29458 7396
rect 29493 7362 29527 7396
rect 29562 7362 29596 7396
rect 29631 7362 29665 7396
rect 29700 7362 29734 7396
rect 29769 7362 29803 7396
rect 29838 7362 29872 7396
rect 29907 7362 29941 7396
rect 29976 7362 30010 7396
rect 30045 7362 30079 7396
rect 30114 7362 30148 7396
rect 30183 7362 30217 7396
rect 30252 7362 30286 7396
rect 30321 7362 30355 7396
rect 30390 7362 30424 7396
rect 30459 7362 30493 7396
rect 30528 7362 30562 7396
rect 28665 7294 28699 7328
rect 28734 7294 28768 7328
rect 28803 7294 28837 7328
rect 28872 7294 28906 7328
rect 28941 7294 28975 7328
rect 29010 7294 29044 7328
rect 29079 7294 29113 7328
rect 29148 7294 29182 7328
rect 29217 7294 29251 7328
rect 29286 7294 29320 7328
rect 29355 7294 29389 7328
rect 29424 7294 29458 7328
rect 29493 7294 29527 7328
rect 29562 7294 29596 7328
rect 29631 7294 29665 7328
rect 29700 7294 29734 7328
rect 29769 7294 29803 7328
rect 29838 7294 29872 7328
rect 29907 7294 29941 7328
rect 29976 7294 30010 7328
rect 30045 7294 30079 7328
rect 30114 7294 30148 7328
rect 30183 7294 30217 7328
rect 30252 7294 30286 7328
rect 30321 7294 30355 7328
rect 30390 7294 30424 7328
rect 30459 7294 30493 7328
rect 30528 7294 30562 7328
rect 30597 7294 30971 7940
rect 28641 6915 28811 7221
rect 28641 6846 28675 6880
rect 28709 6846 28743 6880
rect 28777 6846 28811 6880
rect 28641 6777 28675 6811
rect 28709 6777 28743 6811
rect 28777 6777 28811 6811
rect 28641 6708 28675 6742
rect 28709 6708 28743 6742
rect 28777 6708 28811 6742
rect 28641 6639 28675 6673
rect 28709 6639 28743 6673
rect 28777 6639 28811 6673
rect 28641 6570 28675 6604
rect 28709 6570 28743 6604
rect 28777 6570 28811 6604
rect 28641 6501 28675 6535
rect 28709 6501 28743 6535
rect 28777 6501 28811 6535
rect 28641 6432 28675 6466
rect 28709 6432 28743 6466
rect 28777 6432 28811 6466
rect 28641 6363 28675 6397
rect 28709 6363 28743 6397
rect 28777 6363 28811 6397
rect 28641 6294 28675 6328
rect 28709 6294 28743 6328
rect 28777 6294 28811 6328
rect 28641 6225 28675 6259
rect 28709 6225 28743 6259
rect 28777 6225 28811 6259
<< mvpsubdiffcont >>
rect 30214 5967 30248 6001
rect 30283 5967 30317 6001
rect 30352 5967 30386 6001
rect 30421 5967 30455 6001
rect 30490 5967 30524 6001
rect 30559 5967 30593 6001
rect 30628 5967 30662 6001
rect 30697 5967 30731 6001
rect 30766 5967 30800 6001
rect 30835 5967 30869 6001
rect 30904 5967 30938 6001
rect 30973 5967 31007 6001
rect 31042 5967 31076 6001
rect 31111 5967 31145 6001
rect 31180 5967 31214 6001
rect 31249 5967 31283 6001
rect 31318 5967 31352 6001
rect 31387 5967 31421 6001
rect 31455 5967 31489 6001
rect 31523 5967 31557 6001
rect 31591 5967 31625 6001
rect 31659 5967 31693 6001
rect 31727 5967 31761 6001
rect 31795 5967 31829 6001
rect 31863 5967 31897 6001
rect 31931 5967 31965 6001
rect 31999 5967 32033 6001
rect 30214 5895 30248 5929
rect 30283 5895 30317 5929
rect 30352 5895 30386 5929
rect 30421 5895 30455 5929
rect 30490 5895 30524 5929
rect 30559 5895 30593 5929
rect 30628 5895 30662 5929
rect 30697 5895 30731 5929
rect 30766 5895 30800 5929
rect 30835 5895 30869 5929
rect 30904 5895 30938 5929
rect 30973 5895 31007 5929
rect 31042 5895 31076 5929
rect 31111 5895 31145 5929
rect 31180 5895 31214 5929
rect 31249 5895 31283 5929
rect 31318 5895 31352 5929
rect 31387 5895 31421 5929
rect 31455 5895 31489 5929
rect 31523 5895 31557 5929
rect 31591 5895 31625 5929
rect 31659 5895 31693 5929
rect 31727 5895 31761 5929
rect 31795 5895 31829 5929
rect 31863 5895 31897 5929
rect 31931 5895 31965 5929
rect 31999 5895 32033 5929
rect 30214 5823 30248 5857
rect 30283 5823 30317 5857
rect 30352 5823 30386 5857
rect 30421 5823 30455 5857
rect 30490 5823 30524 5857
rect 30559 5823 30593 5857
rect 30628 5823 30662 5857
rect 30697 5823 30731 5857
rect 30766 5823 30800 5857
rect 30835 5823 30869 5857
rect 30904 5823 30938 5857
rect 30973 5823 31007 5857
rect 31042 5823 31076 5857
rect 31111 5823 31145 5857
rect 31180 5823 31214 5857
rect 31249 5823 31283 5857
rect 31318 5823 31352 5857
rect 31387 5823 31421 5857
rect 31455 5823 31489 5857
rect 31523 5823 31557 5857
rect 31591 5823 31625 5857
rect 31659 5823 31693 5857
rect 31727 5823 31761 5857
rect 31795 5823 31829 5857
rect 31863 5823 31897 5857
rect 31931 5823 31965 5857
rect 31999 5823 32033 5857
rect 22836 5465 22870 5499
rect 22905 5465 22939 5499
rect 22974 5465 23008 5499
rect 23043 5465 23077 5499
rect 23112 5465 23146 5499
rect 23181 5465 23215 5499
rect 23250 5465 23284 5499
rect 23319 5465 23353 5499
rect 23388 5465 23422 5499
rect 23457 5465 23491 5499
rect 23526 5465 23560 5499
rect 23595 5465 23629 5499
rect 23664 5465 23698 5499
rect 23733 5465 23767 5499
rect 23802 5465 23836 5499
rect 23871 5465 23905 5499
rect 23940 5465 23974 5499
rect 24009 5465 24043 5499
rect 24078 5465 24112 5499
rect 24147 5465 24181 5499
rect 24216 5465 24250 5499
rect 24285 5465 24319 5499
rect 24354 5465 24388 5499
rect 24423 5465 24457 5499
rect 24492 5465 24526 5499
rect 24561 5465 24595 5499
rect 24630 5465 24664 5499
rect 24699 5465 24733 5499
rect 24768 5465 24802 5499
rect 24837 5465 24871 5499
rect 24906 5465 24940 5499
rect 24975 5465 25009 5499
rect 25044 5465 25078 5499
rect 25113 5465 25147 5499
rect 25181 5465 25215 5499
rect 25249 5465 25283 5499
rect 25317 5465 25351 5499
rect 25385 5465 25419 5499
rect 25453 5465 25487 5499
rect 25521 5465 25555 5499
rect 25589 5465 25623 5499
rect 25657 5465 25691 5499
rect 25725 5465 25759 5499
rect 25793 5465 25827 5499
rect 25861 5465 25895 5499
rect 25929 5465 25963 5499
rect 25997 5465 26031 5499
rect 26065 5465 26099 5499
rect 26133 5465 26167 5499
rect 26201 5465 26235 5499
rect 26269 5465 26303 5499
rect 26337 5465 26371 5499
rect 26405 5465 26439 5499
rect 26473 5465 26507 5499
rect 26541 5465 26575 5499
rect 26609 5465 26643 5499
rect 26740 5465 26774 5499
rect 26809 5465 26843 5499
rect 26878 5465 26912 5499
rect 26947 5465 26981 5499
rect 27016 5465 27050 5499
rect 27085 5465 27119 5499
rect 27154 5465 27188 5499
rect 27223 5465 27257 5499
rect 27292 5465 27326 5499
rect 27361 5465 27395 5499
rect 27430 5465 27464 5499
rect 27499 5465 27533 5499
rect 19955 4209 20125 5399
rect 20167 5365 20201 5399
rect 20247 5365 20281 5399
rect 20327 5365 20361 5399
rect 20407 5365 20441 5399
rect 20167 5297 20201 5331
rect 20247 5297 20281 5331
rect 20327 5297 20361 5331
rect 20407 5297 20441 5331
rect 20167 5229 20201 5263
rect 20247 5229 20281 5263
rect 20327 5229 20361 5263
rect 20407 5229 20441 5263
rect 20167 5161 20201 5195
rect 20247 5161 20281 5195
rect 20327 5161 20361 5195
rect 20407 5161 20441 5195
rect 20167 5093 20201 5127
rect 20247 5093 20281 5127
rect 20327 5093 20361 5127
rect 20407 5093 20441 5127
rect 22836 5387 22870 5421
rect 22905 5387 22939 5421
rect 22974 5387 23008 5421
rect 23043 5387 23077 5421
rect 23112 5387 23146 5421
rect 23181 5387 23215 5421
rect 23250 5387 23284 5421
rect 23319 5387 23353 5421
rect 23388 5387 23422 5421
rect 23457 5387 23491 5421
rect 23526 5387 23560 5421
rect 23595 5387 23629 5421
rect 23664 5387 23698 5421
rect 23733 5387 23767 5421
rect 23802 5387 23836 5421
rect 23871 5387 23905 5421
rect 23940 5387 23974 5421
rect 24009 5387 24043 5421
rect 24078 5387 24112 5421
rect 24147 5387 24181 5421
rect 24216 5387 24250 5421
rect 24285 5387 24319 5421
rect 24354 5387 24388 5421
rect 24423 5387 24457 5421
rect 24492 5387 24526 5421
rect 24561 5387 24595 5421
rect 24630 5387 24664 5421
rect 24699 5387 24733 5421
rect 24768 5387 24802 5421
rect 24837 5387 24871 5421
rect 24906 5387 24940 5421
rect 24975 5387 25009 5421
rect 25044 5387 25078 5421
rect 25113 5387 25147 5421
rect 25181 5387 25215 5421
rect 25249 5387 25283 5421
rect 25317 5387 25351 5421
rect 25385 5387 25419 5421
rect 25453 5387 25487 5421
rect 25521 5387 25555 5421
rect 25589 5387 25623 5421
rect 25657 5387 25691 5421
rect 25725 5387 25759 5421
rect 25793 5387 25827 5421
rect 25861 5387 25895 5421
rect 25929 5387 25963 5421
rect 25997 5387 26031 5421
rect 26065 5387 26099 5421
rect 26133 5387 26167 5421
rect 26201 5387 26235 5421
rect 26269 5387 26303 5421
rect 26337 5387 26371 5421
rect 26405 5387 26439 5421
rect 26473 5387 26507 5421
rect 26541 5387 26575 5421
rect 26609 5387 26643 5421
rect 26740 5397 26774 5431
rect 26809 5397 26843 5431
rect 26878 5397 26912 5431
rect 26947 5397 26981 5431
rect 27016 5397 27050 5431
rect 27085 5397 27119 5431
rect 27154 5397 27188 5431
rect 27223 5397 27257 5431
rect 27292 5397 27326 5431
rect 27361 5397 27395 5431
rect 27430 5397 27464 5431
rect 27499 5397 27533 5431
rect 22836 5309 22870 5343
rect 22905 5309 22939 5343
rect 22974 5309 23008 5343
rect 23043 5309 23077 5343
rect 23112 5309 23146 5343
rect 23181 5309 23215 5343
rect 23250 5309 23284 5343
rect 23319 5309 23353 5343
rect 23388 5309 23422 5343
rect 23457 5309 23491 5343
rect 23526 5309 23560 5343
rect 23595 5309 23629 5343
rect 23664 5309 23698 5343
rect 23733 5309 23767 5343
rect 23802 5309 23836 5343
rect 23871 5309 23905 5343
rect 23940 5309 23974 5343
rect 24009 5309 24043 5343
rect 24078 5309 24112 5343
rect 24147 5309 24181 5343
rect 24216 5309 24250 5343
rect 24285 5309 24319 5343
rect 24354 5309 24388 5343
rect 24423 5309 24457 5343
rect 24492 5309 24526 5343
rect 24561 5309 24595 5343
rect 24630 5309 24664 5343
rect 24699 5309 24733 5343
rect 24768 5309 24802 5343
rect 24837 5309 24871 5343
rect 24906 5309 24940 5343
rect 24975 5309 25009 5343
rect 25044 5309 25078 5343
rect 25113 5309 25147 5343
rect 25181 5309 25215 5343
rect 25249 5309 25283 5343
rect 25317 5309 25351 5343
rect 25385 5309 25419 5343
rect 25453 5309 25487 5343
rect 25521 5309 25555 5343
rect 25589 5309 25623 5343
rect 25657 5309 25691 5343
rect 25725 5309 25759 5343
rect 25793 5309 25827 5343
rect 25861 5309 25895 5343
rect 25929 5309 25963 5343
rect 25997 5309 26031 5343
rect 26065 5309 26099 5343
rect 26133 5309 26167 5343
rect 26201 5309 26235 5343
rect 26269 5309 26303 5343
rect 26337 5309 26371 5343
rect 26405 5309 26439 5343
rect 26473 5309 26507 5343
rect 26541 5309 26575 5343
rect 26609 5309 26643 5343
rect 26740 5329 26774 5363
rect 26809 5329 26843 5363
rect 26878 5329 26912 5363
rect 26947 5329 26981 5363
rect 27016 5329 27050 5363
rect 27085 5329 27119 5363
rect 27154 5329 27188 5363
rect 27223 5329 27257 5363
rect 27292 5329 27326 5363
rect 27361 5329 27395 5363
rect 27430 5329 27464 5363
rect 27499 5329 27533 5363
rect 22836 5231 22870 5265
rect 22905 5231 22939 5265
rect 22974 5231 23008 5265
rect 23043 5231 23077 5265
rect 23112 5231 23146 5265
rect 23181 5231 23215 5265
rect 23250 5231 23284 5265
rect 23319 5231 23353 5265
rect 23388 5231 23422 5265
rect 23457 5231 23491 5265
rect 23526 5231 23560 5265
rect 23595 5231 23629 5265
rect 23664 5231 23698 5265
rect 23733 5231 23767 5265
rect 23802 5231 23836 5265
rect 23871 5231 23905 5265
rect 23940 5231 23974 5265
rect 24009 5231 24043 5265
rect 24078 5231 24112 5265
rect 24147 5231 24181 5265
rect 24216 5231 24250 5265
rect 24285 5231 24319 5265
rect 24354 5231 24388 5265
rect 24423 5231 24457 5265
rect 24492 5231 24526 5265
rect 24561 5231 24595 5265
rect 24630 5231 24664 5265
rect 24699 5231 24733 5265
rect 24768 5231 24802 5265
rect 24837 5231 24871 5265
rect 24906 5231 24940 5265
rect 24975 5231 25009 5265
rect 25044 5231 25078 5265
rect 25113 5231 25147 5265
rect 25181 5231 25215 5265
rect 25249 5231 25283 5265
rect 25317 5231 25351 5265
rect 25385 5231 25419 5265
rect 25453 5231 25487 5265
rect 25521 5231 25555 5265
rect 25589 5231 25623 5265
rect 25657 5231 25691 5265
rect 25725 5231 25759 5265
rect 25793 5231 25827 5265
rect 25861 5231 25895 5265
rect 25929 5231 25963 5265
rect 25997 5231 26031 5265
rect 26065 5231 26099 5265
rect 26133 5231 26167 5265
rect 26201 5231 26235 5265
rect 26269 5231 26303 5265
rect 26337 5231 26371 5265
rect 26405 5231 26439 5265
rect 26473 5231 26507 5265
rect 26541 5231 26575 5265
rect 26609 5231 26643 5265
rect 26740 5261 26774 5295
rect 26809 5261 26843 5295
rect 26878 5261 26912 5295
rect 26947 5261 26981 5295
rect 27016 5261 27050 5295
rect 27085 5261 27119 5295
rect 27154 5261 27188 5295
rect 27223 5261 27257 5295
rect 27292 5261 27326 5295
rect 27361 5261 27395 5295
rect 27430 5261 27464 5295
rect 27499 5261 27533 5295
rect 26740 5193 26774 5227
rect 26809 5193 26843 5227
rect 26878 5193 26912 5227
rect 26947 5193 26981 5227
rect 27016 5193 27050 5227
rect 27085 5193 27119 5227
rect 27154 5193 27188 5227
rect 27223 5193 27257 5227
rect 27292 5193 27326 5227
rect 27361 5193 27395 5227
rect 27430 5193 27464 5227
rect 27499 5193 27533 5227
rect 22836 5153 22870 5187
rect 22905 5153 22939 5187
rect 22974 5153 23008 5187
rect 23043 5153 23077 5187
rect 23112 5153 23146 5187
rect 23181 5153 23215 5187
rect 23250 5153 23284 5187
rect 23319 5153 23353 5187
rect 23388 5153 23422 5187
rect 23457 5153 23491 5187
rect 23526 5153 23560 5187
rect 23595 5153 23629 5187
rect 23664 5153 23698 5187
rect 23733 5153 23767 5187
rect 23802 5153 23836 5187
rect 23871 5153 23905 5187
rect 23940 5153 23974 5187
rect 24009 5153 24043 5187
rect 24078 5153 24112 5187
rect 24147 5153 24181 5187
rect 24216 5153 24250 5187
rect 24285 5153 24319 5187
rect 24354 5153 24388 5187
rect 24423 5153 24457 5187
rect 24492 5153 24526 5187
rect 24561 5153 24595 5187
rect 24630 5153 24664 5187
rect 24699 5153 24733 5187
rect 24768 5153 24802 5187
rect 24837 5153 24871 5187
rect 24906 5153 24940 5187
rect 24975 5153 25009 5187
rect 25044 5153 25078 5187
rect 25113 5153 25147 5187
rect 25181 5153 25215 5187
rect 25249 5153 25283 5187
rect 25317 5153 25351 5187
rect 25385 5153 25419 5187
rect 25453 5153 25487 5187
rect 25521 5153 25555 5187
rect 25589 5153 25623 5187
rect 25657 5153 25691 5187
rect 25725 5153 25759 5187
rect 25793 5153 25827 5187
rect 25861 5153 25895 5187
rect 25929 5153 25963 5187
rect 25997 5153 26031 5187
rect 26065 5153 26099 5187
rect 26133 5153 26167 5187
rect 26201 5153 26235 5187
rect 26269 5153 26303 5187
rect 26337 5153 26371 5187
rect 26405 5153 26439 5187
rect 26473 5153 26507 5187
rect 26541 5153 26575 5187
rect 26609 5153 26643 5187
rect 26740 5125 26774 5159
rect 26809 5125 26843 5159
rect 26878 5125 26912 5159
rect 26947 5125 26981 5159
rect 27016 5125 27050 5159
rect 27085 5125 27119 5159
rect 27154 5125 27188 5159
rect 27223 5125 27257 5159
rect 27292 5125 27326 5159
rect 27361 5125 27395 5159
rect 27430 5125 27464 5159
rect 27499 5125 27533 5159
rect 20167 5025 20201 5059
rect 20247 5025 20281 5059
rect 20327 5025 20361 5059
rect 20407 5025 20441 5059
rect 20167 4957 20201 4991
rect 20247 4957 20281 4991
rect 20327 4957 20361 4991
rect 20407 4957 20441 4991
rect 20167 4889 20201 4923
rect 20247 4889 20281 4923
rect 20327 4889 20361 4923
rect 20407 4889 20441 4923
rect 20167 4821 20201 4855
rect 20247 4821 20281 4855
rect 20327 4821 20361 4855
rect 20407 4821 20441 4855
rect 20167 4753 20201 4787
rect 20247 4753 20281 4787
rect 20327 4753 20361 4787
rect 20407 4753 20441 4787
rect 20167 4685 20201 4719
rect 20247 4685 20281 4719
rect 20327 4685 20361 4719
rect 20407 4685 20441 4719
rect 20167 4617 20201 4651
rect 20247 4617 20281 4651
rect 20327 4617 20361 4651
rect 20407 4617 20441 4651
rect 20167 4549 20201 4583
rect 20247 4549 20281 4583
rect 20327 4549 20361 4583
rect 20407 4549 20441 4583
rect 20167 4481 20201 4515
rect 20247 4481 20281 4515
rect 20327 4481 20361 4515
rect 20407 4481 20441 4515
rect 20167 4413 20201 4447
rect 20247 4413 20281 4447
rect 20327 4413 20361 4447
rect 20407 4413 20441 4447
rect 20167 4345 20201 4379
rect 20247 4345 20281 4379
rect 20327 4345 20361 4379
rect 20407 4345 20441 4379
rect 20167 4277 20201 4311
rect 20247 4277 20281 4311
rect 20327 4277 20361 4311
rect 20407 4277 20441 4311
rect 20167 4209 20201 4243
rect 20247 4209 20281 4243
rect 20327 4209 20361 4243
rect 20407 4209 20441 4243
rect 20167 4141 20201 4175
rect 20247 4141 20281 4175
rect 20327 4141 20361 4175
rect 20407 4141 20441 4175
rect 26740 5057 26774 5091
rect 26809 5057 26843 5091
rect 26878 5057 26912 5091
rect 26947 5057 26981 5091
rect 27016 5057 27050 5091
rect 27085 5057 27119 5091
rect 27154 5057 27188 5091
rect 27223 5057 27257 5091
rect 27292 5057 27326 5091
rect 27361 5057 27395 5091
rect 27430 5057 27464 5091
rect 27499 5057 27533 5091
rect 26740 4989 26774 5023
rect 26809 4989 26843 5023
rect 26878 4989 26912 5023
rect 26947 4989 26981 5023
rect 27016 4989 27050 5023
rect 27085 4989 27119 5023
rect 27154 4989 27188 5023
rect 27223 4989 27257 5023
rect 27292 4989 27326 5023
rect 27361 4989 27395 5023
rect 27430 4989 27464 5023
rect 27499 4989 27533 5023
rect 26740 4921 26774 4955
rect 26809 4921 26843 4955
rect 26878 4921 26912 4955
rect 26947 4921 26981 4955
rect 27016 4921 27050 4955
rect 27085 4921 27119 4955
rect 27154 4921 27188 4955
rect 27223 4921 27257 4955
rect 27292 4921 27326 4955
rect 27361 4921 27395 4955
rect 27430 4921 27464 4955
rect 27499 4921 27533 4955
rect 26740 4853 26774 4887
rect 26809 4853 26843 4887
rect 26878 4853 26912 4887
rect 26947 4853 26981 4887
rect 27016 4853 27050 4887
rect 27085 4853 27119 4887
rect 27154 4853 27188 4887
rect 27223 4853 27257 4887
rect 27292 4853 27326 4887
rect 27361 4853 27395 4887
rect 27430 4853 27464 4887
rect 27499 4853 27533 4887
rect 26740 4785 26774 4819
rect 26809 4785 26843 4819
rect 26878 4785 26912 4819
rect 26947 4785 26981 4819
rect 27016 4785 27050 4819
rect 27085 4785 27119 4819
rect 27154 4785 27188 4819
rect 27223 4785 27257 4819
rect 27292 4785 27326 4819
rect 27361 4785 27395 4819
rect 27430 4785 27464 4819
rect 27499 4785 27533 4819
rect 26740 4717 26774 4751
rect 26809 4717 26843 4751
rect 26878 4717 26912 4751
rect 26947 4717 26981 4751
rect 27016 4717 27050 4751
rect 27085 4717 27119 4751
rect 27154 4717 27188 4751
rect 27223 4717 27257 4751
rect 27292 4717 27326 4751
rect 27361 4717 27395 4751
rect 27430 4717 27464 4751
rect 27499 4717 27533 4751
rect 26740 4649 26774 4683
rect 26809 4649 26843 4683
rect 26878 4649 26912 4683
rect 26947 4649 26981 4683
rect 27016 4649 27050 4683
rect 27085 4649 27119 4683
rect 27154 4649 27188 4683
rect 27223 4649 27257 4683
rect 27292 4649 27326 4683
rect 27361 4649 27395 4683
rect 27430 4649 27464 4683
rect 27499 4649 27533 4683
rect 26740 4581 26774 4615
rect 26809 4581 26843 4615
rect 26878 4581 26912 4615
rect 26947 4581 26981 4615
rect 27016 4581 27050 4615
rect 27085 4581 27119 4615
rect 27154 4581 27188 4615
rect 27223 4581 27257 4615
rect 27292 4581 27326 4615
rect 27361 4581 27395 4615
rect 27430 4581 27464 4615
rect 27499 4581 27533 4615
rect 26740 4513 26774 4547
rect 26809 4513 26843 4547
rect 26878 4513 26912 4547
rect 26947 4513 26981 4547
rect 27016 4513 27050 4547
rect 27085 4513 27119 4547
rect 27154 4513 27188 4547
rect 27223 4513 27257 4547
rect 27292 4513 27326 4547
rect 27361 4513 27395 4547
rect 27430 4513 27464 4547
rect 27499 4513 27533 4547
rect 26740 4445 26774 4479
rect 26809 4445 26843 4479
rect 26878 4445 26912 4479
rect 26947 4445 26981 4479
rect 27016 4445 27050 4479
rect 27085 4445 27119 4479
rect 27154 4445 27188 4479
rect 27223 4445 27257 4479
rect 27292 4445 27326 4479
rect 27361 4445 27395 4479
rect 27430 4445 27464 4479
rect 27499 4445 27533 4479
rect 26740 4377 26774 4411
rect 26809 4377 26843 4411
rect 26878 4377 26912 4411
rect 26947 4377 26981 4411
rect 27016 4377 27050 4411
rect 27085 4377 27119 4411
rect 27154 4377 27188 4411
rect 27223 4377 27257 4411
rect 27292 4377 27326 4411
rect 27361 4377 27395 4411
rect 27430 4377 27464 4411
rect 27499 4377 27533 4411
rect 26740 4309 26774 4343
rect 26809 4309 26843 4343
rect 26878 4309 26912 4343
rect 26947 4309 26981 4343
rect 27016 4309 27050 4343
rect 27085 4309 27119 4343
rect 27154 4309 27188 4343
rect 27223 4309 27257 4343
rect 27292 4309 27326 4343
rect 27361 4309 27395 4343
rect 27430 4309 27464 4343
rect 27499 4309 27533 4343
rect 26740 4241 26774 4275
rect 26809 4241 26843 4275
rect 26878 4241 26912 4275
rect 26947 4241 26981 4275
rect 27016 4241 27050 4275
rect 27085 4241 27119 4275
rect 27154 4241 27188 4275
rect 27223 4241 27257 4275
rect 27292 4241 27326 4275
rect 27361 4241 27395 4275
rect 27430 4241 27464 4275
rect 27499 4241 27533 4275
rect 27568 4241 28690 5499
rect 28777 5465 28811 5499
rect 28847 5465 28881 5499
rect 28917 5465 28951 5499
rect 28987 5465 29021 5499
rect 29057 5465 29091 5499
rect 29127 5465 29161 5499
rect 29197 5465 29231 5499
rect 29267 5465 29301 5499
rect 29337 5465 29371 5499
rect 29407 5465 29441 5499
rect 29477 5465 29511 5499
rect 29547 5465 29581 5499
rect 29617 5465 29651 5499
rect 29687 5465 29721 5499
rect 29757 5465 29791 5499
rect 29827 5465 29861 5499
rect 29896 5465 29930 5499
rect 29965 5465 29999 5499
rect 30034 5465 30068 5499
rect 30103 5465 30137 5499
rect 30172 5465 30206 5499
rect 28777 5397 28811 5431
rect 28847 5397 28881 5431
rect 28917 5397 28951 5431
rect 28987 5397 29021 5431
rect 29057 5397 29091 5431
rect 29127 5397 29161 5431
rect 29197 5397 29231 5431
rect 29267 5397 29301 5431
rect 29337 5397 29371 5431
rect 29407 5397 29441 5431
rect 29477 5397 29511 5431
rect 29547 5397 29581 5431
rect 29617 5397 29651 5431
rect 29687 5397 29721 5431
rect 29757 5397 29791 5431
rect 29827 5397 29861 5431
rect 29896 5397 29930 5431
rect 29965 5397 29999 5431
rect 30034 5397 30068 5431
rect 30103 5397 30137 5431
rect 30172 5397 30206 5431
rect 28777 5329 28811 5363
rect 28847 5329 28881 5363
rect 28917 5329 28951 5363
rect 28987 5329 29021 5363
rect 29057 5329 29091 5363
rect 29127 5329 29161 5363
rect 29197 5329 29231 5363
rect 29267 5329 29301 5363
rect 29337 5329 29371 5363
rect 29407 5329 29441 5363
rect 29477 5329 29511 5363
rect 29547 5329 29581 5363
rect 29617 5329 29651 5363
rect 29687 5329 29721 5363
rect 29757 5329 29791 5363
rect 29827 5329 29861 5363
rect 29896 5329 29930 5363
rect 29965 5329 29999 5363
rect 30034 5329 30068 5363
rect 30103 5329 30137 5363
rect 30172 5329 30206 5363
rect 28777 5261 28811 5295
rect 28847 5261 28881 5295
rect 28917 5261 28951 5295
rect 28987 5261 29021 5295
rect 29057 5261 29091 5295
rect 29127 5261 29161 5295
rect 29197 5261 29231 5295
rect 29267 5261 29301 5295
rect 29337 5261 29371 5295
rect 29407 5261 29441 5295
rect 29477 5261 29511 5295
rect 29547 5261 29581 5295
rect 29617 5261 29651 5295
rect 29687 5261 29721 5295
rect 29757 5261 29791 5295
rect 29827 5261 29861 5295
rect 29896 5261 29930 5295
rect 29965 5261 29999 5295
rect 30034 5261 30068 5295
rect 30103 5261 30137 5295
rect 30172 5261 30206 5295
rect 28777 5193 28811 5227
rect 28847 5193 28881 5227
rect 28917 5193 28951 5227
rect 28987 5193 29021 5227
rect 29057 5193 29091 5227
rect 29127 5193 29161 5227
rect 29197 5193 29231 5227
rect 29267 5193 29301 5227
rect 29337 5193 29371 5227
rect 29407 5193 29441 5227
rect 29477 5193 29511 5227
rect 29547 5193 29581 5227
rect 29617 5193 29651 5227
rect 29687 5193 29721 5227
rect 29757 5193 29791 5227
rect 29827 5193 29861 5227
rect 29896 5193 29930 5227
rect 29965 5193 29999 5227
rect 30034 5193 30068 5227
rect 30103 5193 30137 5227
rect 30172 5193 30206 5227
rect 28777 5125 28811 5159
rect 28847 5125 28881 5159
rect 28917 5125 28951 5159
rect 28987 5125 29021 5159
rect 29057 5125 29091 5159
rect 29127 5125 29161 5159
rect 29197 5125 29231 5159
rect 29267 5125 29301 5159
rect 29337 5125 29371 5159
rect 29407 5125 29441 5159
rect 29477 5125 29511 5159
rect 29547 5125 29581 5159
rect 29617 5125 29651 5159
rect 29687 5125 29721 5159
rect 29757 5125 29791 5159
rect 29827 5125 29861 5159
rect 29896 5125 29930 5159
rect 29965 5125 29999 5159
rect 30034 5125 30068 5159
rect 30103 5125 30137 5159
rect 30172 5125 30206 5159
rect 28777 5057 28811 5091
rect 28847 5057 28881 5091
rect 28917 5057 28951 5091
rect 28987 5057 29021 5091
rect 29057 5057 29091 5091
rect 29127 5057 29161 5091
rect 29197 5057 29231 5091
rect 29267 5057 29301 5091
rect 29337 5057 29371 5091
rect 29407 5057 29441 5091
rect 29477 5057 29511 5091
rect 29547 5057 29581 5091
rect 29617 5057 29651 5091
rect 29687 5057 29721 5091
rect 29757 5057 29791 5091
rect 29827 5057 29861 5091
rect 29896 5057 29930 5091
rect 29965 5057 29999 5091
rect 30034 5057 30068 5091
rect 30103 5057 30137 5091
rect 30172 5057 30206 5091
rect 28777 4989 28811 5023
rect 28847 4989 28881 5023
rect 28917 4989 28951 5023
rect 28987 4989 29021 5023
rect 29057 4989 29091 5023
rect 29127 4989 29161 5023
rect 29197 4989 29231 5023
rect 29267 4989 29301 5023
rect 29337 4989 29371 5023
rect 29407 4989 29441 5023
rect 29477 4989 29511 5023
rect 29547 4989 29581 5023
rect 29617 4989 29651 5023
rect 29687 4989 29721 5023
rect 29757 4989 29791 5023
rect 29827 4989 29861 5023
rect 29896 4989 29930 5023
rect 29965 4989 29999 5023
rect 30034 4989 30068 5023
rect 30103 4989 30137 5023
rect 30172 4989 30206 5023
rect 28777 4921 28811 4955
rect 28847 4921 28881 4955
rect 28917 4921 28951 4955
rect 28987 4921 29021 4955
rect 29057 4921 29091 4955
rect 29127 4921 29161 4955
rect 29197 4921 29231 4955
rect 29267 4921 29301 4955
rect 29337 4921 29371 4955
rect 29407 4921 29441 4955
rect 29477 4921 29511 4955
rect 29547 4921 29581 4955
rect 29617 4921 29651 4955
rect 29687 4921 29721 4955
rect 29757 4921 29791 4955
rect 29827 4921 29861 4955
rect 29896 4921 29930 4955
rect 29965 4921 29999 4955
rect 30034 4921 30068 4955
rect 30103 4921 30137 4955
rect 30172 4921 30206 4955
rect 28777 4853 28811 4887
rect 28847 4853 28881 4887
rect 28917 4853 28951 4887
rect 28987 4853 29021 4887
rect 29057 4853 29091 4887
rect 29127 4853 29161 4887
rect 29197 4853 29231 4887
rect 29267 4853 29301 4887
rect 29337 4853 29371 4887
rect 29407 4853 29441 4887
rect 29477 4853 29511 4887
rect 29547 4853 29581 4887
rect 29617 4853 29651 4887
rect 29687 4853 29721 4887
rect 29757 4853 29791 4887
rect 29827 4853 29861 4887
rect 29896 4853 29930 4887
rect 29965 4853 29999 4887
rect 30034 4853 30068 4887
rect 30103 4853 30137 4887
rect 30172 4853 30206 4887
rect 28777 4785 28811 4819
rect 28847 4785 28881 4819
rect 28917 4785 28951 4819
rect 28987 4785 29021 4819
rect 29057 4785 29091 4819
rect 29127 4785 29161 4819
rect 29197 4785 29231 4819
rect 29267 4785 29301 4819
rect 29337 4785 29371 4819
rect 29407 4785 29441 4819
rect 29477 4785 29511 4819
rect 29547 4785 29581 4819
rect 29617 4785 29651 4819
rect 29687 4785 29721 4819
rect 29757 4785 29791 4819
rect 29827 4785 29861 4819
rect 29896 4785 29930 4819
rect 29965 4785 29999 4819
rect 30034 4785 30068 4819
rect 30103 4785 30137 4819
rect 30172 4785 30206 4819
rect 28777 4717 28811 4751
rect 28847 4717 28881 4751
rect 28917 4717 28951 4751
rect 28987 4717 29021 4751
rect 29057 4717 29091 4751
rect 29127 4717 29161 4751
rect 29197 4717 29231 4751
rect 29267 4717 29301 4751
rect 29337 4717 29371 4751
rect 29407 4717 29441 4751
rect 29477 4717 29511 4751
rect 29547 4717 29581 4751
rect 29617 4717 29651 4751
rect 29687 4717 29721 4751
rect 29757 4717 29791 4751
rect 29827 4717 29861 4751
rect 29896 4717 29930 4751
rect 29965 4717 29999 4751
rect 30034 4717 30068 4751
rect 30103 4717 30137 4751
rect 30172 4717 30206 4751
rect 20167 4073 20201 4107
rect 20247 4073 20281 4107
rect 20327 4073 20361 4107
rect 20407 4073 20441 4107
rect 20167 4005 20201 4039
rect 20247 4005 20281 4039
rect 20327 4005 20361 4039
rect 20407 4005 20441 4039
rect 20167 3937 20201 3971
rect 20247 3937 20281 3971
rect 20327 3937 20361 3971
rect 20407 3937 20441 3971
rect 20167 3869 20201 3903
rect 20247 3869 20281 3903
rect 20327 3869 20361 3903
rect 20407 3869 20441 3903
rect 20167 3801 20201 3835
rect 20247 3801 20281 3835
rect 20327 3801 20361 3835
rect 20407 3801 20441 3835
rect 20167 3733 20201 3767
rect 20247 3733 20281 3767
rect 20327 3733 20361 3767
rect 20407 3733 20441 3767
rect 20167 3665 20201 3699
rect 20247 3665 20281 3699
rect 20327 3665 20361 3699
rect 20407 3665 20441 3699
rect 20167 3597 20201 3631
rect 20247 3597 20281 3631
rect 20327 3597 20361 3631
rect 20407 3597 20441 3631
rect 20167 3529 20201 3563
rect 20247 3529 20281 3563
rect 20327 3529 20361 3563
rect 20407 3529 20441 3563
rect 20167 3461 20201 3495
rect 20247 3461 20281 3495
rect 20327 3461 20361 3495
rect 20407 3461 20441 3495
rect 20167 3393 20201 3427
rect 20247 3393 20281 3427
rect 20327 3393 20361 3427
rect 20407 3393 20441 3427
rect 20167 3325 20201 3359
rect 20247 3325 20281 3359
rect 20327 3325 20361 3359
rect 20407 3325 20441 3359
rect 20167 3257 20201 3291
rect 20247 3257 20281 3291
rect 20327 3257 20361 3291
rect 20407 3257 20441 3291
rect 20167 3189 20201 3223
rect 20247 3189 20281 3223
rect 20327 3189 20361 3223
rect 20407 3189 20441 3223
rect 20167 3121 20201 3155
rect 20247 3121 20281 3155
rect 20327 3121 20361 3155
rect 20407 3121 20441 3155
rect 20167 3053 20201 3087
rect 20247 3053 20281 3087
rect 20327 3053 20361 3087
rect 20407 3053 20441 3087
rect 20167 2985 20201 3019
rect 20247 2985 20281 3019
rect 20327 2985 20361 3019
rect 20407 2985 20441 3019
rect 20167 2917 20201 2951
rect 20247 2917 20281 2951
rect 20327 2917 20361 2951
rect 20407 2917 20441 2951
rect 20167 2849 20201 2883
rect 20247 2849 20281 2883
rect 20327 2849 20361 2883
rect 20407 2849 20441 2883
rect 20167 2781 20201 2815
rect 20247 2781 20281 2815
rect 20327 2781 20361 2815
rect 20407 2781 20441 2815
rect 20167 2713 20201 2747
rect 20247 2713 20281 2747
rect 20327 2713 20361 2747
rect 20407 2713 20441 2747
rect 20167 2644 20201 2678
rect 20247 2644 20281 2678
rect 20327 2644 20361 2678
rect 20407 2644 20441 2678
rect 22559 3015 22593 3049
rect 22657 3015 22691 3049
rect 22755 3015 22789 3049
rect 22559 2943 22593 2977
rect 22657 2943 22691 2977
rect 22755 2943 22789 2977
rect 22559 2870 22593 2904
rect 22657 2870 22691 2904
rect 22755 2870 22789 2904
rect 22559 2797 22593 2831
rect 22657 2797 22691 2831
rect 22755 2797 22789 2831
rect 22559 2724 22593 2758
rect 22657 2724 22691 2758
rect 22755 2724 22789 2758
rect 22559 2651 22593 2685
rect 22657 2651 22691 2685
rect 22755 2651 22789 2685
rect 18172 2551 18206 2585
rect 18241 2551 18275 2585
rect 18310 2551 18344 2585
rect 18379 2551 18413 2585
rect 18448 2551 18482 2585
rect 18517 2551 18551 2585
rect 18586 2551 18620 2585
rect 18655 2551 18689 2585
rect 18724 2551 18758 2585
rect 18793 2551 18827 2585
rect 18861 2551 18895 2585
rect 18929 2551 18963 2585
rect 18997 2551 19031 2585
rect 19065 2551 19099 2585
rect 19133 2551 19167 2585
rect 19201 2551 19235 2585
rect 19269 2551 19303 2585
rect 19337 2551 19371 2585
rect 19405 2551 19439 2585
rect 19473 2551 19507 2585
rect 19541 2551 19575 2585
rect 19609 2551 19643 2585
rect 19677 2551 19711 2585
rect 19745 2551 19779 2585
rect 19813 2551 19847 2585
rect 19881 2551 19915 2585
rect 19949 2551 19983 2585
rect 20017 2551 20051 2585
rect 20085 2551 20119 2585
rect 20153 2551 20187 2585
rect 20221 2551 20255 2585
rect 20289 2551 20323 2585
rect 20357 2551 20391 2585
rect 20425 2551 20459 2585
rect 20493 2551 20527 2585
rect 20561 2551 20595 2585
rect 20629 2551 20663 2585
rect 20697 2551 20731 2585
rect 20765 2551 20799 2585
rect 20833 2551 20867 2585
rect 20901 2551 20935 2585
rect 20969 2551 21003 2585
rect 21037 2551 21071 2585
rect 21105 2551 21139 2585
rect 21173 2551 21207 2585
rect 21241 2551 21275 2585
rect 21309 2551 21343 2585
rect 21377 2551 21411 2585
rect 21445 2551 21479 2585
rect 21513 2551 21547 2585
rect 21581 2551 21615 2585
rect 21649 2551 21683 2585
rect 21717 2551 21751 2585
rect 21785 2551 21819 2585
rect 21853 2551 21887 2585
rect 21921 2551 21955 2585
rect 21989 2551 22023 2585
rect 22057 2551 22091 2585
rect 22125 2551 22159 2585
rect 22193 2551 22227 2585
rect 22261 2551 22295 2585
rect 22329 2551 22363 2585
rect 22397 2551 22431 2585
rect 22465 2551 22499 2585
rect 22559 2578 22593 2612
rect 22657 2578 22691 2612
rect 22755 2578 22789 2612
rect 16579 2481 16613 2515
rect 16650 2481 16684 2515
rect 16721 2481 16755 2515
rect 16792 2481 16826 2515
rect 16863 2481 16897 2515
rect 16933 2481 16967 2515
rect 17003 2481 17037 2515
rect 17073 2481 17107 2515
rect 17143 2481 17177 2515
rect 17213 2481 17247 2515
rect 17283 2481 17317 2515
rect 17353 2481 17387 2515
rect 17423 2481 17457 2515
rect 17493 2481 17527 2515
rect 17563 2481 17597 2515
rect 17633 2481 17667 2515
rect 17703 2481 17737 2515
rect 17773 2481 17807 2515
rect 17843 2481 17877 2515
rect 17913 2481 17947 2515
rect 17983 2481 18017 2515
rect 18053 2481 18087 2515
rect 18172 2481 18206 2515
rect 18241 2481 18275 2515
rect 18310 2481 18344 2515
rect 18379 2481 18413 2515
rect 18448 2481 18482 2515
rect 18517 2481 18551 2515
rect 18586 2481 18620 2515
rect 18655 2481 18689 2515
rect 18724 2481 18758 2515
rect 18793 2481 18827 2515
rect 18861 2481 18895 2515
rect 18929 2481 18963 2515
rect 18997 2481 19031 2515
rect 19065 2481 19099 2515
rect 19133 2481 19167 2515
rect 19201 2481 19235 2515
rect 19269 2481 19303 2515
rect 19337 2481 19371 2515
rect 19405 2481 19439 2515
rect 19473 2481 19507 2515
rect 19541 2481 19575 2515
rect 19609 2481 19643 2515
rect 19677 2481 19711 2515
rect 19745 2481 19779 2515
rect 19813 2481 19847 2515
rect 19881 2481 19915 2515
rect 19949 2481 19983 2515
rect 20017 2481 20051 2515
rect 20085 2481 20119 2515
rect 20153 2481 20187 2515
rect 20221 2481 20255 2515
rect 20289 2481 20323 2515
rect 20357 2481 20391 2515
rect 20425 2481 20459 2515
rect 20493 2481 20527 2515
rect 20561 2481 20595 2515
rect 20629 2481 20663 2515
rect 20697 2481 20731 2515
rect 20765 2481 20799 2515
rect 20833 2481 20867 2515
rect 20901 2481 20935 2515
rect 20969 2481 21003 2515
rect 21037 2481 21071 2515
rect 21105 2481 21139 2515
rect 21173 2481 21207 2515
rect 21241 2481 21275 2515
rect 21309 2481 21343 2515
rect 21377 2481 21411 2515
rect 21445 2481 21479 2515
rect 21513 2481 21547 2515
rect 21581 2481 21615 2515
rect 21649 2481 21683 2515
rect 21717 2481 21751 2515
rect 21785 2481 21819 2515
rect 21853 2481 21887 2515
rect 21921 2481 21955 2515
rect 21989 2481 22023 2515
rect 22057 2481 22091 2515
rect 22125 2481 22159 2515
rect 22193 2481 22227 2515
rect 22261 2481 22295 2515
rect 22329 2481 22363 2515
rect 22397 2481 22431 2515
rect 22465 2481 22499 2515
rect 22559 2505 22593 2539
rect 22657 2505 22691 2539
rect 22755 2505 22789 2539
rect 22347 2369 22381 2403
rect 22415 2369 22449 2403
rect 22483 2369 22517 2403
rect 22551 2369 22585 2403
rect 22619 2369 22653 2403
rect 22687 2369 22721 2403
rect 22755 2369 22789 2403
rect 22347 2294 22381 2328
rect 22415 2294 22449 2328
rect 22483 2294 22517 2328
rect 22551 2294 22585 2328
rect 22619 2294 22653 2328
rect 22687 2294 22721 2328
rect 22755 2294 22789 2328
rect 22347 2218 22381 2252
rect 22415 2218 22449 2252
rect 22483 2218 22517 2252
rect 22551 2218 22585 2252
rect 22619 2218 22653 2252
rect 22687 2218 22721 2252
rect 22755 2218 22789 2252
rect 22347 2142 22381 2176
rect 22415 2142 22449 2176
rect 22483 2142 22517 2176
rect 22551 2142 22585 2176
rect 22619 2142 22653 2176
rect 22687 2142 22721 2176
rect 22755 2142 22789 2176
rect 22347 2066 22381 2100
rect 22415 2066 22449 2100
rect 22483 2066 22517 2100
rect 22551 2066 22585 2100
rect 22619 2066 22653 2100
rect 22687 2066 22721 2100
rect 22755 2066 22789 2100
rect 22347 1990 22381 2024
rect 22415 1990 22449 2024
rect 22483 1990 22517 2024
rect 22551 1990 22585 2024
rect 22619 1990 22653 2024
rect 22687 1990 22721 2024
rect 22755 1990 22789 2024
rect 22347 1914 22381 1948
rect 22415 1914 22449 1948
rect 22483 1914 22517 1948
rect 22551 1914 22585 1948
rect 22619 1914 22653 1948
rect 22687 1914 22721 1948
rect 22755 1914 22789 1948
rect 22347 1838 22381 1872
rect 22415 1838 22449 1872
rect 22483 1838 22517 1872
rect 22551 1838 22585 1872
rect 22619 1838 22653 1872
rect 22687 1838 22721 1872
rect 22755 1838 22789 1872
rect 22347 1762 22381 1796
rect 22415 1762 22449 1796
rect 22483 1762 22517 1796
rect 22551 1762 22585 1796
rect 22619 1762 22653 1796
rect 22687 1762 22721 1796
rect 22755 1762 22789 1796
rect 26787 2239 26821 2273
rect 26858 2239 26892 2273
rect 26929 2239 26963 2273
rect 27000 2239 27034 2273
rect 27071 2239 27105 2273
rect 27142 2239 27176 2273
rect 27213 2239 27247 2273
rect 27284 2239 27318 2273
rect 27354 2239 27388 2273
rect 27424 2239 27458 2273
rect 27494 2239 27528 2273
rect 27564 2239 27598 2273
rect 27634 2239 27668 2273
rect 27704 2239 27738 2273
rect 27774 2239 27808 2273
rect 27844 2239 27878 2273
rect 27914 2239 27948 2273
rect 27984 2239 28018 2273
rect 28054 2239 28088 2273
rect 28124 2239 28158 2273
rect 28194 2239 28228 2273
rect 28264 2239 28298 2273
rect 28334 2239 28368 2273
rect 26787 2171 26821 2205
rect 26858 2171 26892 2205
rect 26929 2171 26963 2205
rect 27000 2171 27034 2205
rect 27071 2171 27105 2205
rect 27142 2171 27176 2205
rect 27213 2171 27247 2205
rect 27284 2171 27318 2205
rect 27354 2171 27388 2205
rect 27424 2171 27458 2205
rect 27494 2171 27528 2205
rect 27564 2171 27598 2205
rect 27634 2171 27668 2205
rect 27704 2171 27738 2205
rect 27774 2171 27808 2205
rect 27844 2171 27878 2205
rect 27914 2171 27948 2205
rect 27984 2171 28018 2205
rect 28054 2171 28088 2205
rect 28124 2171 28158 2205
rect 28194 2171 28228 2205
rect 28264 2171 28298 2205
rect 28334 2171 28368 2205
rect 26787 2103 26821 2137
rect 26858 2103 26892 2137
rect 26929 2103 26963 2137
rect 27000 2103 27034 2137
rect 27071 2103 27105 2137
rect 27142 2103 27176 2137
rect 27213 2103 27247 2137
rect 27284 2103 27318 2137
rect 27354 2103 27388 2137
rect 27424 2103 27458 2137
rect 27494 2103 27528 2137
rect 27564 2103 27598 2137
rect 27634 2103 27668 2137
rect 27704 2103 27738 2137
rect 27774 2103 27808 2137
rect 27844 2103 27878 2137
rect 27914 2103 27948 2137
rect 27984 2103 28018 2137
rect 28054 2103 28088 2137
rect 28124 2103 28158 2137
rect 28194 2103 28228 2137
rect 28264 2103 28298 2137
rect 28334 2103 28368 2137
rect 26787 2035 26821 2069
rect 26858 2035 26892 2069
rect 26929 2035 26963 2069
rect 27000 2035 27034 2069
rect 27071 2035 27105 2069
rect 27142 2035 27176 2069
rect 27213 2035 27247 2069
rect 27284 2035 27318 2069
rect 27354 2035 27388 2069
rect 27424 2035 27458 2069
rect 27494 2035 27528 2069
rect 27564 2035 27598 2069
rect 27634 2035 27668 2069
rect 27704 2035 27738 2069
rect 27774 2035 27808 2069
rect 27844 2035 27878 2069
rect 27914 2035 27948 2069
rect 27984 2035 28018 2069
rect 28054 2035 28088 2069
rect 28124 2035 28158 2069
rect 28194 2035 28228 2069
rect 28264 2035 28298 2069
rect 28334 2035 28368 2069
rect 26787 1967 26821 2001
rect 26858 1967 26892 2001
rect 26929 1967 26963 2001
rect 27000 1967 27034 2001
rect 27071 1967 27105 2001
rect 27142 1967 27176 2001
rect 27213 1967 27247 2001
rect 27284 1967 27318 2001
rect 27354 1967 27388 2001
rect 27424 1967 27458 2001
rect 27494 1967 27528 2001
rect 27564 1967 27598 2001
rect 27634 1967 27668 2001
rect 27704 1967 27738 2001
rect 27774 1967 27808 2001
rect 27844 1967 27878 2001
rect 27914 1967 27948 2001
rect 27984 1967 28018 2001
rect 28054 1967 28088 2001
rect 28124 1967 28158 2001
rect 28194 1967 28228 2001
rect 28264 1967 28298 2001
rect 28334 1967 28368 2001
rect 26787 1899 26821 1933
rect 26858 1899 26892 1933
rect 26929 1899 26963 1933
rect 27000 1899 27034 1933
rect 27071 1899 27105 1933
rect 27142 1899 27176 1933
rect 27213 1899 27247 1933
rect 27284 1899 27318 1933
rect 27354 1899 27388 1933
rect 27424 1899 27458 1933
rect 27494 1899 27528 1933
rect 27564 1899 27598 1933
rect 27634 1899 27668 1933
rect 27704 1899 27738 1933
rect 27774 1899 27808 1933
rect 27844 1899 27878 1933
rect 27914 1899 27948 1933
rect 27984 1899 28018 1933
rect 28054 1899 28088 1933
rect 28124 1899 28158 1933
rect 28194 1899 28228 1933
rect 28264 1899 28298 1933
rect 28334 1899 28368 1933
rect 26787 1831 26821 1865
rect 26858 1831 26892 1865
rect 26929 1831 26963 1865
rect 27000 1831 27034 1865
rect 27071 1831 27105 1865
rect 27142 1831 27176 1865
rect 27213 1831 27247 1865
rect 27284 1831 27318 1865
rect 27354 1831 27388 1865
rect 27424 1831 27458 1865
rect 27494 1831 27528 1865
rect 27564 1831 27598 1865
rect 27634 1831 27668 1865
rect 27704 1831 27738 1865
rect 27774 1831 27808 1865
rect 27844 1831 27878 1865
rect 27914 1831 27948 1865
rect 27984 1831 28018 1865
rect 28054 1831 28088 1865
rect 28124 1831 28158 1865
rect 28194 1831 28228 1865
rect 28264 1831 28298 1865
rect 28334 1831 28368 1865
rect 26787 1763 26821 1797
rect 26858 1763 26892 1797
rect 26929 1763 26963 1797
rect 27000 1763 27034 1797
rect 27071 1763 27105 1797
rect 27142 1763 27176 1797
rect 27213 1763 27247 1797
rect 27284 1763 27318 1797
rect 27354 1763 27388 1797
rect 27424 1763 27458 1797
rect 27494 1763 27528 1797
rect 27564 1763 27598 1797
rect 27634 1763 27668 1797
rect 27704 1763 27738 1797
rect 27774 1763 27808 1797
rect 27844 1763 27878 1797
rect 27914 1763 27948 1797
rect 27984 1763 28018 1797
rect 28054 1763 28088 1797
rect 28124 1763 28158 1797
rect 28194 1763 28228 1797
rect 28264 1763 28298 1797
rect 28334 1763 28368 1797
rect 26787 1695 26821 1729
rect 26858 1695 26892 1729
rect 26929 1695 26963 1729
rect 27000 1695 27034 1729
rect 27071 1695 27105 1729
rect 27142 1695 27176 1729
rect 27213 1695 27247 1729
rect 27284 1695 27318 1729
rect 27354 1695 27388 1729
rect 27424 1695 27458 1729
rect 27494 1695 27528 1729
rect 27564 1695 27598 1729
rect 27634 1695 27668 1729
rect 27704 1695 27738 1729
rect 27774 1695 27808 1729
rect 27844 1695 27878 1729
rect 27914 1695 27948 1729
rect 27984 1695 28018 1729
rect 28054 1695 28088 1729
rect 28124 1695 28158 1729
rect 28194 1695 28228 1729
rect 28264 1695 28298 1729
rect 28334 1695 28368 1729
rect 26753 1609 26787 1643
rect 26849 1609 26883 1643
rect 26945 1609 26979 1643
rect 26753 1537 26787 1571
rect 26849 1537 26883 1571
rect 26945 1537 26979 1571
rect 26753 1465 26787 1499
rect 26849 1465 26883 1499
rect 26945 1465 26979 1499
rect 26753 1392 26787 1426
rect 26849 1392 26883 1426
rect 26945 1392 26979 1426
rect 26753 1319 26787 1353
rect 26849 1319 26883 1353
rect 26945 1319 26979 1353
rect 26753 1246 26787 1280
rect 26849 1246 26883 1280
rect 26945 1246 26979 1280
rect 26753 1173 26787 1207
rect 26849 1173 26883 1207
rect 26945 1173 26979 1207
rect 26753 1100 26787 1134
rect 26849 1100 26883 1134
rect 26945 1100 26979 1134
rect 26753 1027 26787 1061
rect 26849 1027 26883 1061
rect 26945 1027 26979 1061
rect 26753 954 26787 988
rect 26849 954 26883 988
rect 26945 954 26979 988
rect 26753 881 26787 915
rect 26849 881 26883 915
rect 26945 881 26979 915
<< mvnsubdiffcont >>
rect 17811 22514 17913 23432
rect 17811 22445 17845 22479
rect 17879 22445 17913 22479
rect 17811 22376 17845 22410
rect 17879 22376 17913 22410
rect 17811 22307 17845 22341
rect 17879 22307 17913 22341
rect 17811 22238 17845 22272
rect 17879 22238 17913 22272
rect 17811 22169 17845 22203
rect 17879 22169 17913 22203
rect 17811 22100 17845 22134
rect 17879 22100 17913 22134
rect 17811 22031 17845 22065
rect 17879 22031 17913 22065
rect 17811 21962 17845 21996
rect 17879 21962 17913 21996
rect 17811 21893 17845 21927
rect 17879 21893 17913 21927
rect 17811 21824 17845 21858
rect 17879 21824 17913 21858
rect 17811 21755 17845 21789
rect 17879 21755 17913 21789
rect 17811 21686 17845 21720
rect 17879 21686 17913 21720
rect 17811 21617 17845 21651
rect 17879 21617 17913 21651
rect 17811 21548 17845 21582
rect 17879 21548 17913 21582
rect 17811 21479 17845 21513
rect 17879 21479 17913 21513
rect 17811 21410 17845 21444
rect 17879 21410 17913 21444
rect 17811 21341 17845 21375
rect 17879 21341 17913 21375
rect 17811 21272 17845 21306
rect 17879 21272 17913 21306
rect 17811 21203 17845 21237
rect 17879 21203 17913 21237
rect 17811 21134 17845 21168
rect 17879 21134 17913 21168
rect 17811 21065 17845 21099
rect 17879 21065 17913 21099
rect 17811 20996 17845 21030
rect 17879 20996 17913 21030
rect 17811 20927 17845 20961
rect 17879 20927 17913 20961
rect 17811 20858 17845 20892
rect 17879 20858 17913 20892
rect 17811 20789 17845 20823
rect 17879 20789 17913 20823
rect 17811 20720 17845 20754
rect 17879 20720 17913 20754
rect 17811 20651 17845 20685
rect 17879 20651 17913 20685
rect 17811 20582 17845 20616
rect 17879 20582 17913 20616
rect 17811 20513 17845 20547
rect 17879 20513 17913 20547
rect 17811 20444 17845 20478
rect 17879 20444 17913 20478
rect 17811 20375 17845 20409
rect 17879 20375 17913 20409
rect 17811 20306 17845 20340
rect 17879 20306 17913 20340
<< locali >>
rect 447 33062 448 41880
rect 626 33062 627 41880
rect 447 33023 627 33062
rect 447 32989 448 33023
rect 482 32989 520 33023
rect 554 32989 592 33023
rect 626 32989 627 33023
rect 447 32950 627 32989
rect 447 32916 448 32950
rect 482 32916 520 32950
rect 554 32916 592 32950
rect 626 32916 627 32950
rect 447 32877 627 32916
rect 447 32843 448 32877
rect 482 32843 520 32877
rect 554 32843 592 32877
rect 626 32843 627 32877
rect 447 32804 627 32843
rect 447 32770 448 32804
rect 482 32770 520 32804
rect 554 32770 592 32804
rect 626 32770 627 32804
rect 447 32731 627 32770
rect 447 32697 448 32731
rect 482 32697 520 32731
rect 554 32697 592 32731
rect 626 32697 627 32731
rect 447 32658 627 32697
rect 447 32624 448 32658
rect 482 32624 520 32658
rect 554 32624 592 32658
rect 626 32624 627 32658
rect 447 32585 627 32624
rect 447 32551 448 32585
rect 482 32551 520 32585
rect 554 32551 592 32585
rect 626 32551 627 32585
rect 447 32512 627 32551
rect 447 32478 448 32512
rect 482 32478 520 32512
rect 554 32478 592 32512
rect 626 32478 627 32512
rect 447 32439 627 32478
rect 447 32405 448 32439
rect 482 32405 520 32439
rect 554 32405 592 32439
rect 626 32405 627 32439
rect 447 32366 627 32405
rect 447 32332 448 32366
rect 482 32332 520 32366
rect 554 32332 592 32366
rect 626 32332 627 32366
rect 447 32293 627 32332
rect 447 32259 448 32293
rect 482 32259 520 32293
rect 554 32259 592 32293
rect 626 32259 627 32293
rect 447 32220 627 32259
rect 447 32186 448 32220
rect 482 32186 520 32220
rect 554 32186 592 32220
rect 626 32186 627 32220
rect 447 32147 627 32186
rect 447 32113 448 32147
rect 482 32113 520 32147
rect 554 32113 592 32147
rect 626 32113 627 32147
rect 447 32074 627 32113
rect 447 32040 448 32074
rect 482 32040 520 32074
rect 554 32040 592 32074
rect 626 32040 627 32074
rect 447 32001 627 32040
rect 447 31967 448 32001
rect 482 31967 520 32001
rect 554 31967 592 32001
rect 626 31967 627 32001
rect 447 31928 627 31967
rect 447 31894 448 31928
rect 482 31894 520 31928
rect 554 31894 592 31928
rect 626 31894 627 31928
rect 447 31855 627 31894
rect 447 31821 448 31855
rect 482 31821 520 31855
rect 554 31821 592 31855
rect 626 31821 627 31855
rect 447 31782 627 31821
rect 447 31748 448 31782
rect 482 31748 520 31782
rect 554 31748 592 31782
rect 626 31748 627 31782
rect 447 31709 627 31748
rect 447 31675 448 31709
rect 482 31675 520 31709
rect 554 31675 592 31709
rect 626 31675 627 31709
rect 447 31636 627 31675
rect 447 31602 448 31636
rect 482 31602 520 31636
rect 554 31602 592 31636
rect 626 31602 627 31636
rect 447 31563 627 31602
rect 447 31529 448 31563
rect 482 31529 520 31563
rect 554 31529 592 31563
rect 626 31529 627 31563
rect 447 31490 627 31529
rect 447 31456 448 31490
rect 482 31456 520 31490
rect 554 31456 592 31490
rect 626 31456 627 31490
rect 447 31417 627 31456
rect 447 31383 448 31417
rect 482 31383 520 31417
rect 554 31383 592 31417
rect 626 31383 627 31417
rect 447 31344 627 31383
rect 447 31310 448 31344
rect 482 31310 520 31344
rect 554 31310 592 31344
rect 626 31310 627 31344
rect 447 31271 627 31310
rect 447 31237 448 31271
rect 482 31237 520 31271
rect 554 31237 592 31271
rect 626 31237 627 31271
rect 447 31198 627 31237
rect 447 31164 448 31198
rect 482 31164 520 31198
rect 554 31164 592 31198
rect 626 31164 627 31198
rect 447 31125 627 31164
rect 447 31091 448 31125
rect 482 31091 520 31125
rect 554 31091 592 31125
rect 626 31091 627 31125
rect 447 31052 627 31091
rect 447 31018 448 31052
rect 482 31018 520 31052
rect 554 31018 592 31052
rect 626 31018 627 31052
rect 447 30979 627 31018
rect 447 30945 448 30979
rect 482 30945 520 30979
rect 554 30945 592 30979
rect 626 30945 627 30979
rect 447 30906 627 30945
rect 447 30872 448 30906
rect 482 30872 520 30906
rect 554 30872 592 30906
rect 626 30872 627 30906
rect 447 30833 627 30872
rect 447 30799 448 30833
rect 482 30799 520 30833
rect 554 30799 592 30833
rect 626 30799 627 30833
rect 447 30760 627 30799
rect 447 30726 448 30760
rect 482 30726 520 30760
rect 554 30726 592 30760
rect 626 30726 627 30760
rect 447 30687 627 30726
rect 447 30653 448 30687
rect 482 30653 520 30687
rect 554 30653 592 30687
rect 626 30653 627 30687
rect 447 30614 627 30653
rect 447 30580 448 30614
rect 482 30580 520 30614
rect 554 30580 592 30614
rect 626 30580 627 30614
rect 447 30541 627 30580
rect 447 30507 448 30541
rect 482 30507 520 30541
rect 554 30507 592 30541
rect 626 30507 627 30541
rect 447 30468 627 30507
rect 447 30434 448 30468
rect 482 30434 520 30468
rect 554 30434 592 30468
rect 626 30434 627 30468
rect 447 30395 627 30434
rect 447 30361 448 30395
rect 482 30361 520 30395
rect 554 30361 592 30395
rect 626 30361 627 30395
rect 26913 31540 26916 31574
rect 26950 31540 26996 31574
rect 27030 31540 27076 31574
rect 27110 31540 27156 31574
rect 27190 31540 27236 31574
rect 27270 31540 27273 31574
rect 26913 31501 27273 31540
rect 26913 31467 26916 31501
rect 26950 31467 26996 31501
rect 27030 31467 27076 31501
rect 27110 31467 27156 31501
rect 27190 31467 27236 31501
rect 27270 31467 27273 31501
rect 26913 31428 27273 31467
rect 26913 31394 26916 31428
rect 26950 31394 26996 31428
rect 27030 31394 27076 31428
rect 27110 31394 27156 31428
rect 27190 31394 27236 31428
rect 27270 31394 27273 31428
rect 26913 31355 27273 31394
rect 26913 31321 26916 31355
rect 26950 31321 26996 31355
rect 27030 31321 27076 31355
rect 27110 31321 27156 31355
rect 27190 31321 27236 31355
rect 27270 31321 27273 31355
rect 26913 31282 27273 31321
rect 26913 31248 26916 31282
rect 26950 31248 26996 31282
rect 27030 31248 27076 31282
rect 27110 31248 27156 31282
rect 27190 31248 27236 31282
rect 27270 31248 27273 31282
rect 26913 31209 27273 31248
rect 26913 31175 26916 31209
rect 26950 31175 26996 31209
rect 27030 31175 27076 31209
rect 27110 31175 27156 31209
rect 27190 31175 27236 31209
rect 27270 31175 27273 31209
rect 26913 31136 27273 31175
rect 26913 31102 26916 31136
rect 26950 31102 26996 31136
rect 27030 31102 27076 31136
rect 27110 31102 27156 31136
rect 27190 31102 27236 31136
rect 27270 31102 27273 31136
rect 26913 31063 27273 31102
rect 26913 31029 26916 31063
rect 26950 31029 26996 31063
rect 27030 31029 27076 31063
rect 27110 31029 27156 31063
rect 27190 31029 27236 31063
rect 27270 31029 27273 31063
rect 26913 30990 27273 31029
rect 26913 30956 26916 30990
rect 26950 30956 26996 30990
rect 27030 30956 27076 30990
rect 27110 30956 27156 30990
rect 27190 30956 27236 30990
rect 27270 30956 27273 30990
rect 26913 30917 27273 30956
rect 26913 30883 26916 30917
rect 26950 30883 26996 30917
rect 27030 30883 27076 30917
rect 27110 30883 27156 30917
rect 27190 30883 27236 30917
rect 27270 30883 27273 30917
rect 26913 30844 27273 30883
rect 26913 30810 26916 30844
rect 26950 30810 26996 30844
rect 27030 30810 27076 30844
rect 27110 30810 27156 30844
rect 27190 30810 27236 30844
rect 27270 30810 27273 30844
rect 26913 30771 27273 30810
rect 26913 30737 26916 30771
rect 26950 30737 26996 30771
rect 27030 30737 27076 30771
rect 27110 30737 27156 30771
rect 27190 30737 27236 30771
rect 27270 30737 27273 30771
rect 26913 30698 27273 30737
rect 26913 30664 26916 30698
rect 26950 30664 26996 30698
rect 27030 30664 27076 30698
rect 27110 30664 27156 30698
rect 27190 30664 27236 30698
rect 27270 30664 27273 30698
rect 26913 30625 27273 30664
rect 26913 30591 26916 30625
rect 26950 30591 26996 30625
rect 27030 30591 27076 30625
rect 27110 30591 27156 30625
rect 27190 30591 27236 30625
rect 27270 30591 27273 30625
rect 26913 30551 27273 30591
rect 26913 30517 26916 30551
rect 26950 30517 26996 30551
rect 27030 30517 27076 30551
rect 27110 30517 27156 30551
rect 27190 30517 27236 30551
rect 27270 30517 27273 30551
rect 26913 30477 27273 30517
rect 26913 30443 26916 30477
rect 26950 30443 26996 30477
rect 27030 30443 27076 30477
rect 27110 30443 27156 30477
rect 27190 30443 27236 30477
rect 27270 30443 27273 30477
rect 26913 30403 27273 30443
rect 26913 30369 26916 30403
rect 26950 30369 26996 30403
rect 27030 30369 27076 30403
rect 27110 30369 27156 30403
rect 27190 30369 27236 30403
rect 27270 30369 27273 30403
rect 26913 30329 27273 30369
rect 26913 30295 26916 30329
rect 26950 30295 26996 30329
rect 27030 30295 27076 30329
rect 27110 30295 27156 30329
rect 27190 30295 27236 30329
rect 27270 30295 27273 30329
rect 473 30241 579 30275
rect 439 30203 613 30241
rect 473 30169 579 30203
rect 439 30131 613 30169
rect 473 30097 579 30131
rect 439 30059 613 30097
rect 473 30025 579 30059
rect 439 29987 613 30025
rect 473 29953 579 29987
rect 439 29915 613 29953
rect 473 29881 579 29915
rect 439 29843 613 29881
rect 473 29809 579 29843
rect 439 29771 613 29809
rect 473 29737 579 29771
rect 439 29699 613 29737
rect 473 29665 579 29699
rect 439 29627 613 29665
rect 473 29593 579 29627
rect 439 29555 613 29593
rect 473 29521 579 29555
rect 439 29483 613 29521
rect 473 29449 579 29483
rect 439 29411 613 29449
rect 473 29377 579 29411
rect 439 29339 613 29377
rect 473 29305 579 29339
rect 439 29267 613 29305
rect 473 29233 579 29267
rect 439 29195 613 29233
rect 473 29161 579 29195
rect 439 29123 613 29161
rect 473 29089 579 29123
rect 439 29051 613 29089
rect 473 29017 579 29051
rect 439 28979 613 29017
rect 473 28945 579 28979
rect 439 28907 613 28945
rect 473 28873 579 28907
rect 439 28835 613 28873
rect 473 28801 579 28835
rect 439 28763 613 28801
rect 473 28729 579 28763
rect 439 28691 613 28729
rect 473 28657 579 28691
rect 439 28619 613 28657
rect 473 28585 579 28619
rect 439 28547 613 28585
rect 473 28513 579 28547
rect 26913 30255 27273 30295
rect 26913 30221 26916 30255
rect 26950 30221 26996 30255
rect 27030 30221 27076 30255
rect 27110 30221 27156 30255
rect 27190 30221 27236 30255
rect 27270 30221 27273 30255
rect 26913 30181 27273 30221
rect 26913 30147 26916 30181
rect 26950 30147 26996 30181
rect 27030 30147 27076 30181
rect 27110 30147 27156 30181
rect 27190 30147 27236 30181
rect 27270 30147 27273 30181
rect 26913 30107 27273 30147
rect 26913 30073 26916 30107
rect 26950 30073 26996 30107
rect 27030 30073 27076 30107
rect 27110 30073 27156 30107
rect 27190 30073 27236 30107
rect 27270 30073 27273 30107
rect 26913 30033 27273 30073
rect 26913 29999 26916 30033
rect 26950 29999 26996 30033
rect 27030 29999 27076 30033
rect 27110 29999 27156 30033
rect 27190 29999 27236 30033
rect 27270 29999 27273 30033
rect 26913 29959 27273 29999
rect 26913 29925 26916 29959
rect 26950 29925 26996 29959
rect 27030 29925 27076 29959
rect 27110 29925 27156 29959
rect 27190 29925 27236 29959
rect 27270 29925 27273 29959
rect 26913 29885 27273 29925
rect 26913 29851 26916 29885
rect 26950 29851 26996 29885
rect 27030 29851 27076 29885
rect 27110 29851 27156 29885
rect 27190 29851 27236 29885
rect 27270 29851 27273 29885
rect 26913 29811 27273 29851
rect 26913 29777 26916 29811
rect 26950 29777 26996 29811
rect 27030 29777 27076 29811
rect 27110 29777 27156 29811
rect 27190 29777 27236 29811
rect 27270 29777 27273 29811
rect 26913 29737 27273 29777
rect 26913 29703 26916 29737
rect 26950 29703 26996 29737
rect 27030 29703 27076 29737
rect 27110 29703 27156 29737
rect 27190 29703 27236 29737
rect 27270 29703 27273 29737
rect 26913 29663 27273 29703
rect 26913 29629 26916 29663
rect 26950 29629 26996 29663
rect 27030 29629 27076 29663
rect 27110 29629 27156 29663
rect 27190 29629 27236 29663
rect 27270 29629 27273 29663
rect 26913 29589 27273 29629
rect 26913 29555 26916 29589
rect 26950 29555 26996 29589
rect 27030 29555 27076 29589
rect 27110 29555 27156 29589
rect 27190 29555 27236 29589
rect 27270 29555 27273 29589
rect 26913 29515 27273 29555
rect 26913 29481 26916 29515
rect 26950 29481 26996 29515
rect 27030 29481 27076 29515
rect 27110 29481 27156 29515
rect 27190 29481 27236 29515
rect 27270 29481 27273 29515
rect 26913 29441 27273 29481
rect 26913 29407 26916 29441
rect 26950 29407 26996 29441
rect 27030 29407 27076 29441
rect 27110 29407 27156 29441
rect 27190 29407 27236 29441
rect 27270 29407 27273 29441
rect 26913 29367 27273 29407
rect 26913 29333 26916 29367
rect 26950 29333 26996 29367
rect 27030 29333 27076 29367
rect 27110 29333 27156 29367
rect 27190 29333 27236 29367
rect 27270 29333 27273 29367
rect 26913 29293 27273 29333
rect 26913 29259 26916 29293
rect 26950 29259 26996 29293
rect 27030 29259 27076 29293
rect 27110 29259 27156 29293
rect 27190 29259 27236 29293
rect 27270 29259 27273 29293
rect 26913 29219 27273 29259
rect 26913 29185 26916 29219
rect 26950 29185 26996 29219
rect 27030 29185 27076 29219
rect 27110 29185 27156 29219
rect 27190 29185 27236 29219
rect 27270 29185 27273 29219
rect 26913 29145 27273 29185
rect 26913 29111 26916 29145
rect 26950 29111 26996 29145
rect 27030 29111 27076 29145
rect 27110 29111 27156 29145
rect 27190 29111 27236 29145
rect 27270 29111 27273 29145
rect 26913 29071 27273 29111
rect 26913 29037 26916 29071
rect 26950 29037 26996 29071
rect 27030 29037 27076 29071
rect 27110 29037 27156 29071
rect 27190 29037 27236 29071
rect 27270 29037 27273 29071
rect 26913 28997 27273 29037
rect 26913 28963 26916 28997
rect 26950 28963 26996 28997
rect 27030 28963 27076 28997
rect 27110 28963 27156 28997
rect 27190 28963 27236 28997
rect 27270 28963 27273 28997
rect 26913 28923 27273 28963
rect 26913 28889 26916 28923
rect 26950 28889 26996 28923
rect 27030 28889 27076 28923
rect 27110 28889 27156 28923
rect 27190 28889 27236 28923
rect 27270 28889 27273 28923
rect 26913 28849 27273 28889
rect 26913 28815 26916 28849
rect 26950 28815 26996 28849
rect 27030 28815 27076 28849
rect 27110 28815 27156 28849
rect 27190 28815 27236 28849
rect 27270 28815 27273 28849
rect 26913 28775 27273 28815
rect 26913 28741 26916 28775
rect 26950 28741 26996 28775
rect 27030 28741 27076 28775
rect 27110 28741 27156 28775
rect 27190 28741 27236 28775
rect 27270 28741 27273 28775
rect 26913 28701 27273 28741
rect 26913 28667 26916 28701
rect 26950 28667 26996 28701
rect 27030 28667 27076 28701
rect 27110 28667 27156 28701
rect 27190 28667 27236 28701
rect 27270 28667 27273 28701
rect 26913 28627 27273 28667
rect 26913 28593 26916 28627
rect 26950 28593 26996 28627
rect 27030 28593 27076 28627
rect 27110 28593 27156 28627
rect 27190 28593 27236 28627
rect 27270 28593 27273 28627
rect 26913 28553 27273 28593
rect 26913 28519 26916 28553
rect 26950 28519 26996 28553
rect 27030 28519 27076 28553
rect 27110 28519 27156 28553
rect 27190 28519 27236 28553
rect 27270 28519 27273 28553
rect 439 28475 613 28513
rect 473 28441 579 28475
rect 439 28403 613 28441
rect 473 28369 579 28403
rect 439 28331 613 28369
rect 473 28297 579 28331
rect 439 28259 613 28297
rect 473 28225 579 28259
rect 439 28187 613 28225
rect 473 28153 579 28187
rect 439 28115 613 28153
rect 473 28081 579 28115
rect 439 28043 613 28081
rect 473 28009 579 28043
rect 439 27971 613 28009
rect 473 27937 579 27971
rect 439 27899 613 27937
rect 473 27865 579 27899
rect 439 27827 613 27865
rect 473 27793 579 27827
rect 439 27755 613 27793
rect 473 27721 579 27755
rect 439 27683 613 27721
rect 473 27649 579 27683
rect 439 27611 613 27649
rect 473 27577 579 27611
rect 439 27539 613 27577
rect 473 27505 579 27539
rect 439 27467 613 27505
rect 473 27433 579 27467
rect 439 27395 613 27433
rect 473 27361 579 27395
rect 439 27323 613 27361
rect 473 27289 579 27323
rect 439 27251 613 27289
rect 473 27217 579 27251
rect 439 27179 613 27217
rect 473 27145 579 27179
rect 439 27107 613 27145
rect 473 27073 579 27107
rect 439 27035 613 27073
rect 473 27001 579 27035
rect 439 26963 613 27001
rect 473 26929 579 26963
rect 439 26891 613 26929
rect 473 26857 579 26891
rect 439 26819 613 26857
rect 473 26785 579 26819
rect 439 26747 613 26785
rect 473 26713 579 26747
rect 439 26675 613 26713
rect 473 26641 579 26675
rect 439 26603 613 26641
rect 473 26569 579 26603
rect 439 26530 613 26569
rect 473 26496 579 26530
rect 439 26457 613 26496
rect 473 26423 579 26457
rect 439 26384 613 26423
rect 473 26350 579 26384
rect 439 26311 613 26350
rect 473 26277 579 26311
rect 439 26238 613 26277
rect 473 26204 579 26238
rect 439 26165 613 26204
rect 473 26131 579 26165
rect -2255 26071 -1419 26073
rect -2221 26037 -2182 26071
rect -2148 26037 -2109 26071
rect -2075 26037 -2036 26071
rect -2002 26037 -1963 26071
rect -1929 26037 -1890 26071
rect -1856 26037 -1817 26071
rect -1783 26037 -1744 26071
rect -1710 26037 -1671 26071
rect -1637 26037 -1598 26071
rect -1564 26037 -1525 26071
rect -1491 26037 -1453 26071
rect -2255 25997 -1419 26037
rect -2221 25963 -2182 25997
rect -2148 25963 -2109 25997
rect -2075 25963 -2036 25997
rect -2002 25963 -1963 25997
rect -1929 25963 -1890 25997
rect -1856 25963 -1817 25997
rect -1783 25963 -1744 25997
rect -1710 25963 -1671 25997
rect -1637 25963 -1598 25997
rect -1564 25963 -1525 25997
rect -1491 25963 -1453 25997
rect -2255 25923 -1419 25963
rect -2221 25889 -2182 25923
rect -2148 25889 -2109 25923
rect -2075 25889 -2036 25923
rect -2002 25889 -1963 25923
rect -1929 25889 -1890 25923
rect -1856 25889 -1817 25923
rect -1783 25889 -1744 25923
rect -1710 25889 -1671 25923
rect -1637 25889 -1598 25923
rect -1564 25889 -1525 25923
rect -1491 25889 -1453 25923
rect -2255 25849 -1419 25889
rect -2221 25815 -2182 25849
rect -2148 25815 -2109 25849
rect -2075 25815 -2036 25849
rect -2002 25815 -1963 25849
rect -1929 25815 -1890 25849
rect -1856 25815 -1817 25849
rect -1783 25815 -1744 25849
rect -1710 25815 -1671 25849
rect -1637 25815 -1598 25849
rect -1564 25815 -1525 25849
rect -1491 25815 -1453 25849
rect -2255 25775 -1419 25815
rect -2221 25741 -2182 25775
rect -2148 25741 -2109 25775
rect -2075 25741 -2036 25775
rect -2002 25741 -1963 25775
rect -1929 25741 -1890 25775
rect -1856 25741 -1817 25775
rect -1783 25741 -1744 25775
rect -1710 25741 -1671 25775
rect -1637 25741 -1598 25775
rect -1564 25741 -1525 25775
rect -1491 25741 -1453 25775
rect -2255 25701 -1419 25741
rect -2221 25667 -2182 25701
rect -2148 25667 -2109 25701
rect -2075 25667 -2036 25701
rect -2002 25667 -1963 25701
rect -1929 25667 -1890 25701
rect -1856 25667 -1817 25701
rect -1783 25667 -1744 25701
rect -1710 25667 -1671 25701
rect -1637 25667 -1598 25701
rect -1564 25667 -1525 25701
rect -1491 25667 -1453 25701
rect -2255 25627 -1419 25667
rect -2221 25593 -2182 25627
rect -2148 25593 -2109 25627
rect -2075 25593 -2036 25627
rect -2002 25593 -1963 25627
rect -1929 25593 -1890 25627
rect -1856 25593 -1817 25627
rect -1783 25593 -1744 25627
rect -1710 25593 -1671 25627
rect -1637 25593 -1598 25627
rect -1564 25593 -1525 25627
rect -1491 25593 -1453 25627
rect -2255 25591 -1419 25593
rect -1181 25915 2679 25917
rect -1147 25881 -1108 25915
rect -1074 25881 -1035 25915
rect -1001 25881 -962 25915
rect -928 25881 -889 25915
rect -855 25881 -816 25915
rect -782 25881 -743 25915
rect -709 25881 -670 25915
rect -636 25881 -597 25915
rect -563 25881 -524 25915
rect -490 25881 -451 25915
rect -1181 25843 -451 25881
rect -1147 25809 -1108 25843
rect -1074 25809 -1035 25843
rect -1001 25809 -962 25843
rect -928 25809 -889 25843
rect -855 25809 -816 25843
rect -782 25809 -743 25843
rect -709 25809 -670 25843
rect -636 25809 -597 25843
rect -563 25809 -524 25843
rect -490 25809 -451 25843
rect -1181 25771 -451 25809
rect -1147 25737 -1108 25771
rect -1074 25737 -1035 25771
rect -1001 25737 -962 25771
rect -928 25737 -889 25771
rect -855 25737 -816 25771
rect -782 25737 -743 25771
rect -709 25737 -670 25771
rect -636 25737 -597 25771
rect -563 25737 -524 25771
rect -490 25737 -451 25771
rect -1181 25699 -451 25737
rect -1147 25665 -1108 25699
rect -1074 25665 -1035 25699
rect -1001 25665 -962 25699
rect -928 25665 -889 25699
rect -855 25665 -816 25699
rect -782 25665 -743 25699
rect -709 25665 -670 25699
rect -636 25665 -597 25699
rect -563 25665 -524 25699
rect -490 25665 -451 25699
rect -1181 25627 -451 25665
rect -1147 25593 -1108 25627
rect -1074 25593 -1035 25627
rect -1001 25593 -962 25627
rect -928 25593 -889 25627
rect -855 25593 -816 25627
rect -782 25593 -743 25627
rect -709 25593 -670 25627
rect -636 25593 -597 25627
rect -563 25593 -524 25627
rect -490 25593 -451 25627
rect -1181 25591 2679 25593
rect 31966 23611 32020 23645
rect 31932 23570 32054 23611
rect 31966 23536 32020 23570
rect 31932 23495 32054 23536
rect 31966 23461 32020 23495
rect 17811 23432 17913 23456
rect 17777 23395 17778 23429
rect 17913 23395 17978 23429
rect 18012 23395 18013 23429
rect 17777 23356 17811 23395
rect 17913 23356 18013 23395
rect 17777 23322 17778 23356
rect 17913 23322 17978 23356
rect 18012 23322 18013 23356
rect 17777 23283 17811 23322
rect 17913 23283 18013 23322
rect 17777 23249 17778 23283
rect 17913 23249 17978 23283
rect 18012 23249 18013 23283
rect 17777 23210 17811 23249
rect 17913 23210 18013 23249
rect 31932 23420 32054 23461
rect 31966 23386 32020 23420
rect 31932 23345 32054 23386
rect 31966 23311 32020 23345
rect 31932 23270 32054 23311
rect 31966 23236 32020 23270
rect 17777 23176 17778 23210
rect 17913 23176 17978 23210
rect 18012 23176 18013 23210
rect 17777 23137 17811 23176
rect 17913 23137 18013 23176
rect 17777 23103 17778 23137
rect 17913 23103 17978 23137
rect 18012 23103 18013 23137
rect 17777 23064 17811 23103
rect 17913 23064 18013 23103
rect 17777 23030 17778 23064
rect 17913 23030 17978 23064
rect 18012 23030 18013 23064
rect 17777 22991 17811 23030
rect 17913 22991 18013 23030
rect 17777 22957 17778 22991
rect 17913 22957 17978 22991
rect 18012 22957 18013 22991
rect 17777 22918 17811 22957
rect 17913 22918 18013 22957
rect 17777 22884 17778 22918
rect 17913 22884 17978 22918
rect 18012 22884 18013 22918
rect 17777 22845 17811 22884
rect 17913 22845 18013 22884
rect 17777 22811 17778 22845
rect 17913 22811 17978 22845
rect 18012 22811 18013 22845
rect 17777 22772 17811 22811
rect 17913 22772 18013 22811
rect 17777 22738 17778 22772
rect 17913 22738 17978 22772
rect 18012 22738 18013 22772
rect 17777 22699 17811 22738
rect 17913 22699 18013 22738
rect 17777 22665 17778 22699
rect 17913 22665 17978 22699
rect 18012 22665 18013 22699
rect 17777 22626 17811 22665
rect 17913 22626 18013 22665
rect 17777 22592 17778 22626
rect 17913 22592 17978 22626
rect 18012 22592 18013 22626
rect 17777 22553 17811 22592
rect 17913 22553 18013 22592
rect 17777 22519 17778 22553
rect 17913 22519 17978 22553
rect 18012 22519 18013 22553
rect 17777 22514 17811 22519
rect 17913 22514 18013 22519
rect 17777 22480 18013 22514
rect 17777 22446 17778 22480
rect 17812 22479 17878 22480
rect 17912 22479 17978 22480
rect 17845 22446 17878 22479
rect 17913 22446 17978 22479
rect 18012 22446 18013 22480
rect 17777 22445 17811 22446
rect 17845 22445 17879 22446
rect 17913 22445 18013 22446
rect 17777 22410 18013 22445
rect 17777 22407 17811 22410
rect 17845 22407 17879 22410
rect 17913 22407 18013 22410
rect 17777 22373 17778 22407
rect 17845 22376 17878 22407
rect 17913 22376 17978 22407
rect 17812 22373 17878 22376
rect 17912 22373 17978 22376
rect 18012 22373 18013 22407
rect 17777 22341 18013 22373
rect 17777 22334 17811 22341
rect 17845 22334 17879 22341
rect 17913 22334 18013 22341
rect 17777 22300 17778 22334
rect 17845 22307 17878 22334
rect 17913 22307 17978 22334
rect 17812 22300 17878 22307
rect 17912 22300 17978 22307
rect 18012 22300 18013 22334
rect 17777 22272 18013 22300
rect 17777 22261 17811 22272
rect 17845 22261 17879 22272
rect 17913 22261 18013 22272
rect 17777 22227 17778 22261
rect 17845 22238 17878 22261
rect 17913 22238 17978 22261
rect 17812 22227 17878 22238
rect 17912 22227 17978 22238
rect 18012 22227 18013 22261
rect 17777 22203 18013 22227
rect 17777 22188 17811 22203
rect 17845 22188 17879 22203
rect 17913 22188 18013 22203
rect 17777 22154 17778 22188
rect 17845 22169 17878 22188
rect 17913 22169 17978 22188
rect 17812 22154 17878 22169
rect 17912 22154 17978 22169
rect 18012 22154 18013 22188
rect 17777 22134 18013 22154
rect 17777 22115 17811 22134
rect 17845 22115 17879 22134
rect 17913 22115 18013 22134
rect 17777 22081 17778 22115
rect 17845 22100 17878 22115
rect 17913 22100 17978 22115
rect 17812 22081 17878 22100
rect 17912 22081 17978 22100
rect 18012 22081 18013 22115
rect 17777 22065 18013 22081
rect 17777 22042 17811 22065
rect 17845 22042 17879 22065
rect 17913 22042 18013 22065
rect 17777 22008 17778 22042
rect 17845 22031 17878 22042
rect 17913 22031 17978 22042
rect 17812 22008 17878 22031
rect 17912 22008 17978 22031
rect 18012 22008 18013 22042
rect 17777 21996 18013 22008
rect 17777 21968 17811 21996
rect 17845 21968 17879 21996
rect 17913 21968 18013 21996
rect 17777 21934 17778 21968
rect 17845 21962 17878 21968
rect 17913 21962 17978 21968
rect 17812 21934 17878 21962
rect 17912 21934 17978 21962
rect 18012 21934 18013 21968
rect 17777 21927 18013 21934
rect 17777 21894 17811 21927
rect 17845 21894 17879 21927
rect 17913 21894 18013 21927
rect 17777 21860 17778 21894
rect 17845 21893 17878 21894
rect 17913 21893 17978 21894
rect 17812 21860 17878 21893
rect 17912 21860 17978 21893
rect 18012 21860 18013 21894
rect 17777 21858 18013 21860
rect 17777 21824 17811 21858
rect 17845 21824 17879 21858
rect 17913 21824 18013 21858
rect 17777 21820 18013 21824
rect 17777 21786 17778 21820
rect 17812 21789 17878 21820
rect 17912 21789 17978 21820
rect 17845 21786 17878 21789
rect 17913 21786 17978 21789
rect 18012 21786 18013 21820
rect 17777 21755 17811 21786
rect 17845 21755 17879 21786
rect 17913 21755 18013 21786
rect 17777 21746 18013 21755
rect 17777 21712 17778 21746
rect 17812 21720 17878 21746
rect 17912 21720 17978 21746
rect 17845 21712 17878 21720
rect 17913 21712 17978 21720
rect 18012 21712 18013 21746
rect 17777 21686 17811 21712
rect 17845 21686 17879 21712
rect 17913 21686 18013 21712
rect 17777 21672 18013 21686
rect 17777 21638 17778 21672
rect 17812 21651 17878 21672
rect 17912 21651 17978 21672
rect 17845 21638 17878 21651
rect 17913 21638 17978 21651
rect 18012 21638 18013 21672
rect 17777 21617 17811 21638
rect 17845 21617 17879 21638
rect 17913 21617 18013 21638
rect 17777 21598 18013 21617
rect 17777 21564 17778 21598
rect 17812 21582 17878 21598
rect 17912 21582 17978 21598
rect 17845 21564 17878 21582
rect 17913 21564 17978 21582
rect 18012 21564 18013 21598
rect 17777 21548 17811 21564
rect 17845 21548 17879 21564
rect 17913 21548 18013 21564
rect 17777 21524 18013 21548
rect 17777 21490 17778 21524
rect 17812 21513 17878 21524
rect 17912 21513 17978 21524
rect 17845 21490 17878 21513
rect 17913 21490 17978 21513
rect 18012 21490 18013 21524
rect 17777 21479 17811 21490
rect 17845 21479 17879 21490
rect 17913 21479 18013 21490
rect 17777 21450 18013 21479
rect 17777 21416 17778 21450
rect 17812 21444 17878 21450
rect 17912 21444 17978 21450
rect 17845 21416 17878 21444
rect 17913 21416 17978 21444
rect 18012 21416 18013 21450
rect 17777 21410 17811 21416
rect 17845 21410 17879 21416
rect 17913 21410 18013 21416
rect 17777 21376 18013 21410
rect 17777 21342 17778 21376
rect 17812 21375 17878 21376
rect 17912 21375 17978 21376
rect 17845 21342 17878 21375
rect 17913 21342 17978 21375
rect 18012 21342 18013 21376
rect 17777 21341 17811 21342
rect 17845 21341 17879 21342
rect 17913 21341 18013 21342
rect 17777 21306 18013 21341
rect 17777 21302 17811 21306
rect 17845 21302 17879 21306
rect 17913 21302 18013 21306
rect 17777 21268 17778 21302
rect 17845 21272 17878 21302
rect 17913 21272 17978 21302
rect 17812 21268 17878 21272
rect 17912 21268 17978 21272
rect 18012 21268 18013 21302
rect 17777 21237 18013 21268
rect 17777 21228 17811 21237
rect 17845 21228 17879 21237
rect 17913 21228 18013 21237
rect 17777 21194 17778 21228
rect 17845 21203 17878 21228
rect 17913 21203 17978 21228
rect 17812 21194 17878 21203
rect 17912 21194 17978 21203
rect 18012 21194 18013 21228
rect 17777 21168 18013 21194
rect 17777 21154 17811 21168
rect 17845 21154 17879 21168
rect 17913 21154 18013 21168
rect 17777 21120 17778 21154
rect 17845 21134 17878 21154
rect 17913 21134 17978 21154
rect 17812 21120 17878 21134
rect 17912 21120 17978 21134
rect 18012 21120 18013 21154
rect 17777 21099 18013 21120
rect 17777 21080 17811 21099
rect 17845 21080 17879 21099
rect 17913 21080 18013 21099
rect 17777 21046 17778 21080
rect 17845 21065 17878 21080
rect 17913 21065 17978 21080
rect 17812 21046 17878 21065
rect 17912 21046 17978 21065
rect 18012 21046 18013 21080
rect 17777 21030 18013 21046
rect 17777 21006 17811 21030
rect 17845 21006 17879 21030
rect 17913 21006 18013 21030
rect 17777 20972 17778 21006
rect 17845 20996 17878 21006
rect 17913 20996 17978 21006
rect 17812 20972 17878 20996
rect 17912 20972 17978 20996
rect 18012 20972 18013 21006
rect 17777 20961 18013 20972
rect 31758 23121 31802 23155
rect 31836 23121 31880 23155
rect 31914 23121 31958 23155
rect 31992 23121 32036 23155
rect 31724 23081 32070 23121
rect 31758 23047 31802 23081
rect 31836 23047 31880 23081
rect 31914 23047 31958 23081
rect 31992 23047 32036 23081
rect 31724 23007 32070 23047
rect 31758 22973 31802 23007
rect 31836 22973 31880 23007
rect 31914 22973 31958 23007
rect 31992 22973 32036 23007
rect 31724 22933 32070 22973
rect 31758 22899 31802 22933
rect 31836 22899 31880 22933
rect 31914 22899 31958 22933
rect 31992 22899 32036 22933
rect 31724 22859 32070 22899
rect 31758 22825 31802 22859
rect 31836 22825 31880 22859
rect 31914 22825 31958 22859
rect 31992 22825 32036 22859
rect 31724 22785 32070 22825
rect 31758 22751 31802 22785
rect 31836 22751 31880 22785
rect 31914 22751 31958 22785
rect 31992 22751 32036 22785
rect 31724 22711 32070 22751
rect 31758 22677 31802 22711
rect 31836 22677 31880 22711
rect 31914 22677 31958 22711
rect 31992 22677 32036 22711
rect 31724 22637 32070 22677
rect 31758 22603 31802 22637
rect 31836 22603 31880 22637
rect 31914 22603 31958 22637
rect 31992 22603 32036 22637
rect 31724 22563 32070 22603
rect 31758 22529 31802 22563
rect 31836 22529 31880 22563
rect 31914 22529 31958 22563
rect 31992 22529 32036 22563
rect 31724 22489 32070 22529
rect 31758 22455 31802 22489
rect 31836 22455 31880 22489
rect 31914 22455 31958 22489
rect 31992 22455 32036 22489
rect 31724 22415 32070 22455
rect 31758 22381 31802 22415
rect 31836 22381 31880 22415
rect 31914 22381 31958 22415
rect 31992 22381 32036 22415
rect 31724 22341 32070 22381
rect 31758 22307 31802 22341
rect 31836 22307 31880 22341
rect 31914 22307 31958 22341
rect 31992 22307 32036 22341
rect 31724 22267 32070 22307
rect 31758 22233 31802 22267
rect 31836 22233 31880 22267
rect 31914 22233 31958 22267
rect 31992 22233 32036 22267
rect 31724 22193 32070 22233
rect 31758 22159 31802 22193
rect 31836 22159 31880 22193
rect 31914 22159 31958 22193
rect 31992 22159 32036 22193
rect 31724 22119 32070 22159
rect 31758 22085 31802 22119
rect 31836 22085 31880 22119
rect 31914 22085 31958 22119
rect 31992 22085 32036 22119
rect 31724 22045 32070 22085
rect 31758 22011 31802 22045
rect 31836 22011 31880 22045
rect 31914 22011 31958 22045
rect 31992 22011 32036 22045
rect 31724 21971 32070 22011
rect 31758 21937 31802 21971
rect 31836 21937 31880 21971
rect 31914 21937 31958 21971
rect 31992 21937 32036 21971
rect 31724 21897 32070 21937
rect 31758 21863 31802 21897
rect 31836 21863 31880 21897
rect 31914 21863 31958 21897
rect 31992 21863 32036 21897
rect 31724 21823 32070 21863
rect 31758 21789 31802 21823
rect 31836 21789 31880 21823
rect 31914 21789 31958 21823
rect 31992 21789 32036 21823
rect 31724 21749 32070 21789
rect 31758 21715 31802 21749
rect 31836 21715 31880 21749
rect 31914 21715 31958 21749
rect 31992 21715 32036 21749
rect 31724 21675 32070 21715
rect 31758 21641 31802 21675
rect 31836 21641 31880 21675
rect 31914 21641 31958 21675
rect 31992 21641 32036 21675
rect 31724 21601 32070 21641
rect 31758 21567 31802 21601
rect 31836 21567 31880 21601
rect 31914 21567 31958 21601
rect 31992 21567 32036 21601
rect 31724 21527 32070 21567
rect 31758 21493 31802 21527
rect 31836 21493 31880 21527
rect 31914 21493 31958 21527
rect 31992 21493 32036 21527
rect 31724 21452 32070 21493
rect 31758 21418 31802 21452
rect 31836 21418 31880 21452
rect 31914 21418 31958 21452
rect 31992 21418 32036 21452
rect 31724 21377 32070 21418
rect 31758 21343 31802 21377
rect 31836 21343 31880 21377
rect 31914 21343 31958 21377
rect 31992 21343 32036 21377
rect 31724 21302 32070 21343
rect 31758 21268 31802 21302
rect 31836 21268 31880 21302
rect 31914 21268 31958 21302
rect 31992 21268 32036 21302
rect 31724 21227 32070 21268
rect 31758 21193 31802 21227
rect 31836 21193 31880 21227
rect 31914 21193 31958 21227
rect 31992 21193 32036 21227
rect 31724 21152 32070 21193
rect 31758 21118 31802 21152
rect 31836 21118 31880 21152
rect 31914 21118 31958 21152
rect 31992 21118 32036 21152
rect 31724 21077 32070 21118
rect 31758 21043 31802 21077
rect 31836 21043 31880 21077
rect 31914 21043 31958 21077
rect 31992 21043 32036 21077
rect 31724 21002 32070 21043
rect 31758 20968 31802 21002
rect 31836 20968 31880 21002
rect 31914 20968 31958 21002
rect 31992 20968 32036 21002
rect 17777 20932 17811 20961
rect 17845 20932 17879 20961
rect 17913 20932 18013 20961
rect 17777 20898 17778 20932
rect 17845 20927 17878 20932
rect 17913 20927 17978 20932
rect 17812 20898 17878 20927
rect 17912 20898 17978 20927
rect 18012 20898 18013 20932
rect 17777 20892 18013 20898
rect 17777 20858 17811 20892
rect 17845 20858 17879 20892
rect 17913 20858 18013 20892
rect 17777 20824 17778 20858
rect 17812 20824 17878 20858
rect 17912 20824 17978 20858
rect 18012 20824 18013 20858
rect 17777 20823 18013 20824
rect 17777 20789 17811 20823
rect 17845 20789 17879 20823
rect 17913 20789 18013 20823
rect 17777 20784 18013 20789
rect 17777 20750 17778 20784
rect 17812 20754 17878 20784
rect 17912 20754 17978 20784
rect 17845 20750 17878 20754
rect 17913 20750 17978 20754
rect 18012 20750 18013 20784
rect 17777 20720 17811 20750
rect 17845 20720 17879 20750
rect 17913 20720 18013 20750
rect 17777 20710 18013 20720
rect 17777 20676 17778 20710
rect 17812 20685 17878 20710
rect 17912 20685 17978 20710
rect 17845 20676 17878 20685
rect 17913 20676 17978 20685
rect 18012 20676 18013 20710
rect 17777 20651 17811 20676
rect 17845 20651 17879 20676
rect 17913 20651 18013 20676
rect 17777 20636 18013 20651
rect 17777 20602 17778 20636
rect 17812 20616 17878 20636
rect 17912 20616 17978 20636
rect 17845 20602 17878 20616
rect 17913 20602 17978 20616
rect 18012 20602 18013 20636
rect 17777 20582 17811 20602
rect 17845 20582 17879 20602
rect 17913 20582 18013 20602
rect 17777 20562 18013 20582
rect 17777 20528 17778 20562
rect 17812 20547 17878 20562
rect 17912 20547 17978 20562
rect 17845 20528 17878 20547
rect 17913 20528 17978 20547
rect 18012 20528 18013 20562
rect 17777 20513 17811 20528
rect 17845 20513 17879 20528
rect 17913 20513 18013 20528
rect 17777 20488 18013 20513
rect 17777 20454 17778 20488
rect 17812 20478 17878 20488
rect 17912 20478 17978 20488
rect 17845 20454 17878 20478
rect 17913 20454 17978 20478
rect 18012 20454 18013 20488
rect 17777 20444 17811 20454
rect 17845 20444 17879 20454
rect 17913 20444 18013 20454
rect 17777 20414 18013 20444
rect 17777 20380 17778 20414
rect 17812 20409 17878 20414
rect 17912 20409 17978 20414
rect 17845 20380 17878 20409
rect 17913 20380 17978 20409
rect 18012 20380 18013 20414
rect 17777 20375 17811 20380
rect 17845 20375 17879 20380
rect 17913 20375 18013 20380
rect 17777 20340 18013 20375
rect 17777 20306 17778 20340
rect 17845 20306 17878 20340
rect 17913 20306 17978 20340
rect 18012 20306 18013 20340
rect 17811 20282 17913 20306
rect -2255 13313 -2215 13347
rect -2181 13313 -2141 13347
rect -2107 13313 -2067 13347
rect -2033 13313 -1993 13347
rect -1959 13313 -1919 13347
rect -1885 13313 -1845 13347
rect -1811 13313 -1771 13347
rect -1737 13313 -1698 13347
rect -1664 13313 -1625 13347
rect -1591 13313 -1552 13347
rect -2289 13263 -1518 13313
rect -2255 13229 -2215 13263
rect -2181 13229 -2141 13263
rect -2107 13229 -2067 13263
rect -2033 13229 -1993 13263
rect -1959 13229 -1919 13263
rect -1885 13229 -1845 13263
rect -1811 13229 -1771 13263
rect -1737 13229 -1698 13263
rect -1664 13229 -1625 13263
rect -1591 13229 -1552 13263
rect 28641 7906 28665 7940
rect 28699 7906 28734 7940
rect 28768 7906 28803 7940
rect 28837 7906 28872 7940
rect 28906 7906 28941 7940
rect 28975 7906 29010 7940
rect 29044 7906 29079 7940
rect 29113 7906 29148 7940
rect 29182 7906 29217 7940
rect 29251 7906 29286 7940
rect 29320 7906 29355 7940
rect 29389 7906 29424 7940
rect 29458 7906 29493 7940
rect 29527 7906 29562 7940
rect 29596 7906 29631 7940
rect 29665 7906 29700 7940
rect 29734 7906 29769 7940
rect 29803 7906 29838 7940
rect 29872 7906 29907 7940
rect 29941 7906 29976 7940
rect 30010 7906 30045 7940
rect 30079 7906 30114 7940
rect 30148 7906 30183 7940
rect 30217 7906 30252 7940
rect 30286 7906 30321 7940
rect 30355 7906 30390 7940
rect 30424 7906 30459 7940
rect 30493 7906 30528 7940
rect 30562 7906 30597 7940
rect 28641 7872 30597 7906
rect 28641 7838 28665 7872
rect 28699 7838 28734 7872
rect 28768 7838 28803 7872
rect 28837 7838 28872 7872
rect 28906 7838 28941 7872
rect 28975 7838 29010 7872
rect 29044 7838 29079 7872
rect 29113 7838 29148 7872
rect 29182 7838 29217 7872
rect 29251 7838 29286 7872
rect 29320 7838 29355 7872
rect 29389 7838 29424 7872
rect 29458 7838 29493 7872
rect 29527 7838 29562 7872
rect 29596 7838 29631 7872
rect 29665 7838 29700 7872
rect 29734 7838 29769 7872
rect 29803 7838 29838 7872
rect 29872 7838 29907 7872
rect 29941 7838 29976 7872
rect 30010 7838 30045 7872
rect 30079 7838 30114 7872
rect 30148 7838 30183 7872
rect 30217 7838 30252 7872
rect 30286 7838 30321 7872
rect 30355 7838 30390 7872
rect 30424 7838 30459 7872
rect 30493 7838 30528 7872
rect 30562 7838 30597 7872
rect 28641 7804 30597 7838
rect 28641 7770 28665 7804
rect 28699 7770 28734 7804
rect 28768 7770 28803 7804
rect 28837 7770 28872 7804
rect 28906 7770 28941 7804
rect 28975 7770 29010 7804
rect 29044 7770 29079 7804
rect 29113 7770 29148 7804
rect 29182 7770 29217 7804
rect 29251 7770 29286 7804
rect 29320 7770 29355 7804
rect 29389 7770 29424 7804
rect 29458 7770 29493 7804
rect 29527 7770 29562 7804
rect 29596 7770 29631 7804
rect 29665 7770 29700 7804
rect 29734 7770 29769 7804
rect 29803 7770 29838 7804
rect 29872 7770 29907 7804
rect 29941 7770 29976 7804
rect 30010 7770 30045 7804
rect 30079 7770 30114 7804
rect 30148 7770 30183 7804
rect 30217 7770 30252 7804
rect 30286 7770 30321 7804
rect 30355 7770 30390 7804
rect 30424 7770 30459 7804
rect 30493 7770 30528 7804
rect 30562 7770 30597 7804
rect 28641 7736 30597 7770
rect 28641 7702 28665 7736
rect 28699 7702 28734 7736
rect 28768 7702 28803 7736
rect 28837 7702 28872 7736
rect 28906 7702 28941 7736
rect 28975 7702 29010 7736
rect 29044 7702 29079 7736
rect 29113 7702 29148 7736
rect 29182 7702 29217 7736
rect 29251 7702 29286 7736
rect 29320 7702 29355 7736
rect 29389 7702 29424 7736
rect 29458 7702 29493 7736
rect 29527 7702 29562 7736
rect 29596 7702 29631 7736
rect 29665 7702 29700 7736
rect 29734 7702 29769 7736
rect 29803 7702 29838 7736
rect 29872 7702 29907 7736
rect 29941 7702 29976 7736
rect 30010 7702 30045 7736
rect 30079 7702 30114 7736
rect 30148 7702 30183 7736
rect 30217 7702 30252 7736
rect 30286 7702 30321 7736
rect 30355 7702 30390 7736
rect 30424 7702 30459 7736
rect 30493 7702 30528 7736
rect 30562 7702 30597 7736
rect 28641 7668 30597 7702
rect 28641 7634 28665 7668
rect 28699 7634 28734 7668
rect 28768 7634 28803 7668
rect 28837 7634 28872 7668
rect 28906 7634 28941 7668
rect 28975 7634 29010 7668
rect 29044 7634 29079 7668
rect 29113 7634 29148 7668
rect 29182 7634 29217 7668
rect 29251 7634 29286 7668
rect 29320 7634 29355 7668
rect 29389 7634 29424 7668
rect 29458 7634 29493 7668
rect 29527 7634 29562 7668
rect 29596 7634 29631 7668
rect 29665 7634 29700 7668
rect 29734 7634 29769 7668
rect 29803 7634 29838 7668
rect 29872 7634 29907 7668
rect 29941 7634 29976 7668
rect 30010 7634 30045 7668
rect 30079 7634 30114 7668
rect 30148 7634 30183 7668
rect 30217 7634 30252 7668
rect 30286 7634 30321 7668
rect 30355 7634 30390 7668
rect 30424 7634 30459 7668
rect 30493 7634 30528 7668
rect 30562 7634 30597 7668
rect 28641 7600 30597 7634
rect 28641 7566 28665 7600
rect 28699 7566 28734 7600
rect 28768 7566 28803 7600
rect 28837 7566 28872 7600
rect 28906 7566 28941 7600
rect 28975 7566 29010 7600
rect 29044 7566 29079 7600
rect 29113 7566 29148 7600
rect 29182 7566 29217 7600
rect 29251 7566 29286 7600
rect 29320 7566 29355 7600
rect 29389 7566 29424 7600
rect 29458 7566 29493 7600
rect 29527 7566 29562 7600
rect 29596 7566 29631 7600
rect 29665 7566 29700 7600
rect 29734 7566 29769 7600
rect 29803 7566 29838 7600
rect 29872 7566 29907 7600
rect 29941 7566 29976 7600
rect 30010 7566 30045 7600
rect 30079 7566 30114 7600
rect 30148 7566 30183 7600
rect 30217 7566 30252 7600
rect 30286 7566 30321 7600
rect 30355 7566 30390 7600
rect 30424 7566 30459 7600
rect 30493 7566 30528 7600
rect 30562 7566 30597 7600
rect 28641 7532 30597 7566
rect 28641 7498 28665 7532
rect 28699 7498 28734 7532
rect 28768 7498 28803 7532
rect 28837 7498 28872 7532
rect 28906 7498 28941 7532
rect 28975 7498 29010 7532
rect 29044 7498 29079 7532
rect 29113 7498 29148 7532
rect 29182 7498 29217 7532
rect 29251 7498 29286 7532
rect 29320 7498 29355 7532
rect 29389 7498 29424 7532
rect 29458 7498 29493 7532
rect 29527 7498 29562 7532
rect 29596 7498 29631 7532
rect 29665 7498 29700 7532
rect 29734 7498 29769 7532
rect 29803 7498 29838 7532
rect 29872 7498 29907 7532
rect 29941 7498 29976 7532
rect 30010 7498 30045 7532
rect 30079 7498 30114 7532
rect 30148 7498 30183 7532
rect 30217 7498 30252 7532
rect 30286 7498 30321 7532
rect 30355 7498 30390 7532
rect 30424 7498 30459 7532
rect 30493 7498 30528 7532
rect 30562 7498 30597 7532
rect 28641 7464 30597 7498
rect 28641 7430 28665 7464
rect 28699 7430 28734 7464
rect 28768 7430 28803 7464
rect 28837 7439 28872 7464
rect 28906 7439 28941 7464
rect 28975 7439 29010 7464
rect 28860 7430 28872 7439
rect 28933 7430 28941 7439
rect 29006 7430 29010 7439
rect 29044 7439 29079 7464
rect 29044 7430 29045 7439
rect 28641 7405 28826 7430
rect 28860 7405 28899 7430
rect 28933 7405 28972 7430
rect 29006 7405 29045 7430
rect 29113 7439 29148 7464
rect 29182 7439 29217 7464
rect 29251 7439 29286 7464
rect 29320 7439 29355 7464
rect 29389 7439 29424 7464
rect 29458 7439 29493 7464
rect 29527 7439 29562 7464
rect 29596 7439 29631 7464
rect 29665 7439 29700 7464
rect 29734 7439 29769 7464
rect 29803 7439 29838 7464
rect 29113 7430 29117 7439
rect 29182 7430 29189 7439
rect 29251 7430 29261 7439
rect 29320 7430 29333 7439
rect 29389 7430 29405 7439
rect 29458 7430 29477 7439
rect 29527 7430 29549 7439
rect 29596 7430 29621 7439
rect 29665 7430 29693 7439
rect 29734 7430 29765 7439
rect 29803 7430 29837 7439
rect 29872 7430 29907 7464
rect 29941 7439 29976 7464
rect 30010 7439 30045 7464
rect 30079 7439 30114 7464
rect 30148 7439 30183 7464
rect 30217 7439 30252 7464
rect 30286 7439 30321 7464
rect 30355 7439 30390 7464
rect 30424 7439 30459 7464
rect 30493 7439 30528 7464
rect 30562 7439 30597 7464
rect 29943 7430 29976 7439
rect 30015 7430 30045 7439
rect 30087 7430 30114 7439
rect 30159 7430 30183 7439
rect 30231 7430 30252 7439
rect 30303 7430 30321 7439
rect 30375 7430 30390 7439
rect 30447 7430 30459 7439
rect 30519 7430 30528 7439
rect 29079 7405 29117 7430
rect 29151 7405 29189 7430
rect 29223 7405 29261 7430
rect 29295 7405 29333 7430
rect 29367 7405 29405 7430
rect 29439 7405 29477 7430
rect 29511 7405 29549 7430
rect 29583 7405 29621 7430
rect 29655 7405 29693 7430
rect 29727 7405 29765 7430
rect 29799 7405 29837 7430
rect 29871 7405 29909 7430
rect 29943 7405 29981 7430
rect 30015 7405 30053 7430
rect 30087 7405 30125 7430
rect 30159 7405 30197 7430
rect 30231 7405 30269 7430
rect 30303 7405 30341 7430
rect 30375 7405 30413 7430
rect 30447 7405 30485 7430
rect 30519 7405 30557 7430
rect 30591 7405 30597 7439
rect 28641 7396 30597 7405
rect 28641 7375 28665 7396
rect 28555 7362 28665 7375
rect 28699 7362 28734 7396
rect 28768 7364 28803 7396
rect 28788 7362 28803 7364
rect 28837 7362 28872 7396
rect 28906 7362 28941 7396
rect 28975 7362 29010 7396
rect 29044 7362 29079 7396
rect 29113 7362 29148 7396
rect 29182 7362 29217 7396
rect 29251 7362 29286 7396
rect 29320 7362 29355 7396
rect 29389 7362 29424 7396
rect 29458 7362 29493 7396
rect 29527 7362 29562 7396
rect 29596 7362 29631 7396
rect 29665 7362 29700 7396
rect 29734 7362 29769 7396
rect 29803 7362 29838 7396
rect 29872 7362 29907 7396
rect 29941 7362 29976 7396
rect 30010 7362 30045 7396
rect 30079 7362 30114 7396
rect 30148 7362 30183 7396
rect 30217 7362 30252 7396
rect 30286 7362 30321 7396
rect 30355 7362 30390 7396
rect 30424 7362 30459 7396
rect 30493 7362 30528 7396
rect 30562 7362 30597 7396
rect 28555 7330 28754 7362
rect 28788 7330 30597 7362
rect 28555 7328 30597 7330
rect 28555 7294 28665 7328
rect 28699 7294 28734 7328
rect 28768 7294 28803 7328
rect 28837 7327 28872 7328
rect 28906 7327 28941 7328
rect 28837 7294 28866 7327
rect 28906 7294 28940 7327
rect 28975 7294 29010 7328
rect 29044 7327 29079 7328
rect 29113 7327 29148 7328
rect 29182 7327 29217 7328
rect 29251 7327 29286 7328
rect 29320 7327 29355 7328
rect 29389 7327 29424 7328
rect 29458 7327 29493 7328
rect 29048 7294 29079 7327
rect 29122 7294 29148 7327
rect 29196 7294 29217 7327
rect 29270 7294 29286 7327
rect 29344 7294 29355 7327
rect 29418 7294 29424 7327
rect 29491 7294 29493 7327
rect 29527 7327 29562 7328
rect 29596 7327 29631 7328
rect 29665 7327 29700 7328
rect 29734 7327 29769 7328
rect 29803 7327 29838 7328
rect 29872 7327 29907 7328
rect 29941 7327 29976 7328
rect 30010 7327 30045 7328
rect 29527 7294 29530 7327
rect 29596 7294 29603 7327
rect 29665 7294 29676 7327
rect 29734 7294 29749 7327
rect 29803 7294 29822 7327
rect 29872 7294 29895 7327
rect 29941 7294 29968 7327
rect 30010 7294 30041 7327
rect 30079 7294 30114 7328
rect 30148 7294 30183 7328
rect 30217 7327 30252 7328
rect 30286 7327 30321 7328
rect 30355 7327 30390 7328
rect 30424 7327 30459 7328
rect 30493 7327 30528 7328
rect 30562 7327 30597 7328
rect 30221 7294 30252 7327
rect 30294 7294 30321 7327
rect 30367 7294 30390 7327
rect 30440 7294 30459 7327
rect 30513 7294 30528 7327
rect 30586 7294 30597 7327
rect 30971 7294 30995 7940
rect 28555 7293 28866 7294
rect 28900 7293 28940 7294
rect 28974 7293 29014 7294
rect 29048 7293 29088 7294
rect 29122 7293 29162 7294
rect 29196 7293 29236 7294
rect 29270 7293 29310 7294
rect 29344 7293 29384 7294
rect 29418 7293 29457 7294
rect 29491 7293 29530 7294
rect 29564 7293 29603 7294
rect 29637 7293 29676 7294
rect 29710 7293 29749 7294
rect 29783 7293 29822 7294
rect 29856 7293 29895 7294
rect 29929 7293 29968 7294
rect 30002 7293 30041 7294
rect 30075 7293 30114 7294
rect 30148 7293 30187 7294
rect 30221 7293 30260 7294
rect 30294 7293 30333 7294
rect 30367 7293 30406 7294
rect 30440 7293 30479 7294
rect 30513 7293 30552 7294
rect 30586 7293 30625 7294
rect 30659 7293 30698 7294
rect 30732 7293 30771 7294
rect 30805 7293 30844 7294
rect 30878 7293 30917 7294
rect 30951 7293 30983 7294
rect 28555 7289 30983 7293
rect 28555 7255 28754 7289
rect 28788 7255 30983 7289
rect 28555 7246 30983 7255
rect 28555 7221 28866 7246
rect 28555 6915 28641 7221
rect 28811 7212 28866 7221
rect 28900 7212 30983 7246
rect 28811 7208 30983 7212
rect 28811 7165 28979 7208
rect 28811 7131 28866 7165
rect 28900 7131 28979 7165
rect 28811 7083 28979 7131
rect 28811 7049 28866 7083
rect 28900 7049 28979 7083
rect 28811 7001 28979 7049
rect 28811 6967 28866 7001
rect 28900 6967 28979 7001
rect 28811 6919 28979 6967
rect 28811 6915 28866 6919
rect 28555 6913 28866 6915
rect 28555 6880 28754 6913
rect 28788 6885 28866 6913
rect 28900 6885 28979 6919
rect 28788 6880 28979 6885
rect 28555 6846 28641 6880
rect 28675 6846 28709 6880
rect 28743 6879 28754 6880
rect 28743 6846 28777 6879
rect 28811 6846 28979 6880
rect 28555 6837 28979 6846
rect 28555 6811 28754 6837
rect 28788 6811 28866 6837
rect 28555 6777 28641 6811
rect 28675 6777 28709 6811
rect 28743 6803 28754 6811
rect 28811 6803 28866 6811
rect 28900 6803 28979 6837
rect 28743 6777 28777 6803
rect 28811 6784 28979 6803
rect 28555 6742 28811 6777
rect 28555 6708 28641 6742
rect 28675 6708 28709 6742
rect 28743 6708 28777 6742
rect 28555 6673 28811 6708
rect 28555 6639 28641 6673
rect 28675 6639 28709 6673
rect 28743 6639 28777 6673
rect 28555 6604 28811 6639
rect 28555 6570 28641 6604
rect 28675 6570 28709 6604
rect 28743 6570 28777 6604
rect 28555 6535 28811 6570
rect 28555 6501 28641 6535
rect 28675 6501 28709 6535
rect 28743 6501 28777 6535
rect 28555 6466 28811 6501
rect 28555 6432 28641 6466
rect 28675 6432 28709 6466
rect 28743 6432 28777 6466
rect 28555 6397 28811 6432
rect 28555 6363 28641 6397
rect 28675 6363 28709 6397
rect 28743 6363 28777 6397
rect 28555 6328 28811 6363
rect 28555 6294 28641 6328
rect 28675 6294 28709 6328
rect 28743 6294 28777 6328
rect 28555 6259 28811 6294
rect 28555 6225 28641 6259
rect 28675 6225 28709 6259
rect 28743 6225 28777 6259
rect 28555 6201 28811 6225
rect 30092 6001 32057 6002
rect 30092 5967 30214 6001
rect 30248 5967 30283 6001
rect 30317 5967 30352 6001
rect 30386 5967 30421 6001
rect 30455 5967 30490 6001
rect 30524 5967 30559 6001
rect 30593 5967 30628 6001
rect 30662 5967 30697 6001
rect 30731 5967 30766 6001
rect 30800 5967 30835 6001
rect 30869 5967 30904 6001
rect 30938 5967 30973 6001
rect 31007 5967 31042 6001
rect 31076 5967 31111 6001
rect 31145 5967 31180 6001
rect 31214 5967 31249 6001
rect 31283 5967 31318 6001
rect 31352 5967 31387 6001
rect 31421 5967 31455 6001
rect 31489 5967 31523 6001
rect 31557 5967 31591 6001
rect 31625 5967 31659 6001
rect 31693 5967 31727 6001
rect 31761 5967 31795 6001
rect 31829 5967 31863 6001
rect 31897 5967 31931 6001
rect 31965 5967 31999 6001
rect 32033 5967 32057 6001
rect 30092 5929 32057 5967
rect 30092 5895 30214 5929
rect 30248 5895 30283 5929
rect 30317 5895 30352 5929
rect 30386 5895 30421 5929
rect 30455 5895 30490 5929
rect 30524 5895 30559 5929
rect 30593 5895 30628 5929
rect 30662 5895 30697 5929
rect 30731 5895 30766 5929
rect 30800 5895 30835 5929
rect 30869 5895 30904 5929
rect 30938 5895 30973 5929
rect 31007 5895 31042 5929
rect 31076 5895 31111 5929
rect 31145 5895 31180 5929
rect 31214 5895 31249 5929
rect 31283 5895 31318 5929
rect 31352 5895 31387 5929
rect 31421 5895 31455 5929
rect 31489 5895 31523 5929
rect 31557 5895 31591 5929
rect 31625 5895 31659 5929
rect 31693 5895 31727 5929
rect 31761 5895 31795 5929
rect 31829 5895 31863 5929
rect 31897 5895 31931 5929
rect 31965 5895 31999 5929
rect 32033 5895 32057 5929
rect 30092 5857 32057 5895
rect 30092 5823 30214 5857
rect 30248 5835 30283 5857
rect 30317 5835 30352 5857
rect 30386 5835 30421 5857
rect 30455 5835 30490 5857
rect 30524 5835 30559 5857
rect 30593 5835 30628 5857
rect 30250 5823 30283 5835
rect 30325 5823 30352 5835
rect 30400 5823 30421 5835
rect 30475 5823 30490 5835
rect 30550 5823 30559 5835
rect 30625 5823 30628 5835
rect 30662 5835 30697 5857
rect 30731 5835 30766 5857
rect 30800 5835 30835 5857
rect 30869 5835 30904 5857
rect 30938 5835 30973 5857
rect 31007 5835 31042 5857
rect 30662 5823 30666 5835
rect 30731 5823 30741 5835
rect 30800 5823 30816 5835
rect 30869 5823 30891 5835
rect 30938 5823 30966 5835
rect 31007 5823 31041 5835
rect 31076 5823 31111 5857
rect 31145 5835 31180 5857
rect 31214 5835 31249 5857
rect 31283 5835 31318 5857
rect 31352 5835 31387 5857
rect 31421 5835 31455 5857
rect 31150 5823 31180 5835
rect 31225 5823 31249 5835
rect 31300 5823 31318 5835
rect 31375 5823 31387 5835
rect 31450 5823 31455 5835
rect 31489 5835 31523 5857
rect 31557 5835 31591 5857
rect 31625 5835 31659 5857
rect 31693 5835 31727 5857
rect 31761 5835 31795 5857
rect 31829 5835 31863 5857
rect 31489 5823 31491 5835
rect 31557 5823 31566 5835
rect 31625 5823 31640 5835
rect 31693 5823 31714 5835
rect 31761 5823 31788 5835
rect 31829 5823 31862 5835
rect 31897 5823 31931 5857
rect 31965 5835 31999 5857
rect 32033 5835 32057 5857
rect 31970 5823 31999 5835
rect 30092 5801 30216 5823
rect 30250 5801 30291 5823
rect 30325 5801 30366 5823
rect 30400 5801 30441 5823
rect 30475 5801 30516 5823
rect 30550 5801 30591 5823
rect 30625 5801 30666 5823
rect 30700 5801 30741 5823
rect 30775 5801 30816 5823
rect 30850 5801 30891 5823
rect 30925 5801 30966 5823
rect 31000 5801 31041 5823
rect 31075 5801 31116 5823
rect 31150 5801 31191 5823
rect 31225 5801 31266 5823
rect 31300 5801 31341 5823
rect 31375 5801 31416 5823
rect 31450 5801 31491 5823
rect 31525 5801 31566 5823
rect 31600 5801 31640 5823
rect 31674 5801 31714 5823
rect 31748 5801 31788 5823
rect 31822 5801 31862 5823
rect 31896 5801 31936 5823
rect 31970 5801 32010 5823
rect 32044 5822 32057 5835
rect 30092 5768 32044 5801
rect 16808 5545 18955 5546
rect 16842 5511 16881 5545
rect 16915 5511 16954 5545
rect 16988 5511 17027 5545
rect 17061 5511 17100 5545
rect 17134 5511 17173 5545
rect 17207 5511 17246 5545
rect 17280 5511 17319 5545
rect 17353 5511 17392 5545
rect 17426 5511 17465 5545
rect 17499 5511 17538 5545
rect 17572 5511 17611 5545
rect 17645 5511 17684 5545
rect 17718 5511 17757 5545
rect 17791 5511 17830 5545
rect 17864 5511 17903 5545
rect 17937 5511 17976 5545
rect 18010 5511 18049 5545
rect 18083 5511 18122 5545
rect 18156 5511 18195 5545
rect 18229 5511 18268 5545
rect 18302 5511 18341 5545
rect 18375 5511 18414 5545
rect 18448 5511 18487 5545
rect 18521 5511 18560 5545
rect 18594 5511 18633 5545
rect 18667 5511 18705 5545
rect 18739 5511 18777 5545
rect 18811 5511 18849 5545
rect 18883 5511 18921 5545
rect 30092 5540 30230 5768
rect 16808 5467 18955 5511
rect 16842 5433 16881 5467
rect 16915 5433 16954 5467
rect 16988 5433 17027 5467
rect 17061 5433 17100 5467
rect 17134 5433 17173 5467
rect 17207 5433 17246 5467
rect 17280 5433 17319 5467
rect 17353 5433 17392 5467
rect 17426 5433 17465 5467
rect 17499 5433 17538 5467
rect 17572 5433 17611 5467
rect 17645 5433 17684 5467
rect 17718 5433 17757 5467
rect 17791 5433 17830 5467
rect 17864 5433 17903 5467
rect 17937 5433 17976 5467
rect 18010 5433 18049 5467
rect 18083 5433 18122 5467
rect 18156 5433 18195 5467
rect 18229 5433 18268 5467
rect 18302 5433 18341 5467
rect 18375 5433 18414 5467
rect 18448 5433 18487 5467
rect 18521 5433 18560 5467
rect 18594 5433 18633 5467
rect 18667 5433 18705 5467
rect 18739 5433 18777 5467
rect 18811 5433 18849 5467
rect 18883 5433 18921 5467
rect 16808 5389 18955 5433
rect 22812 5499 30230 5540
rect 22812 5465 22836 5499
rect 22870 5465 22905 5499
rect 22939 5465 22974 5499
rect 23008 5465 23043 5499
rect 23077 5465 23112 5499
rect 23146 5465 23181 5499
rect 23215 5465 23250 5499
rect 23284 5465 23319 5499
rect 23353 5465 23388 5499
rect 23422 5465 23457 5499
rect 23491 5465 23526 5499
rect 23560 5465 23595 5499
rect 23629 5465 23664 5499
rect 23698 5465 23733 5499
rect 23767 5465 23802 5499
rect 23836 5465 23871 5499
rect 23905 5465 23940 5499
rect 23974 5465 24009 5499
rect 24043 5465 24078 5499
rect 24112 5465 24147 5499
rect 24181 5465 24216 5499
rect 24250 5465 24285 5499
rect 24319 5465 24354 5499
rect 24388 5465 24423 5499
rect 24457 5465 24492 5499
rect 24526 5465 24561 5499
rect 24595 5465 24630 5499
rect 24664 5465 24699 5499
rect 24733 5465 24768 5499
rect 24802 5465 24837 5499
rect 24871 5465 24906 5499
rect 24940 5465 24975 5499
rect 25009 5465 25044 5499
rect 25078 5465 25113 5499
rect 25147 5465 25181 5499
rect 25215 5465 25249 5499
rect 25283 5465 25317 5499
rect 25351 5465 25385 5499
rect 25419 5465 25453 5499
rect 25487 5465 25521 5499
rect 25555 5465 25589 5499
rect 25623 5465 25657 5499
rect 25691 5465 25725 5499
rect 25759 5465 25793 5499
rect 25827 5465 25861 5499
rect 25895 5465 25929 5499
rect 25963 5465 25997 5499
rect 26031 5465 26065 5499
rect 26099 5465 26133 5499
rect 26167 5465 26201 5499
rect 26235 5465 26269 5499
rect 26303 5465 26337 5499
rect 26371 5465 26405 5499
rect 26439 5465 26473 5499
rect 26507 5465 26541 5499
rect 26575 5465 26609 5499
rect 26643 5465 26740 5499
rect 26774 5465 26809 5499
rect 26843 5465 26878 5499
rect 26912 5465 26947 5499
rect 26981 5465 27016 5499
rect 27050 5465 27085 5499
rect 27119 5465 27154 5499
rect 27188 5465 27223 5499
rect 27257 5465 27292 5499
rect 27326 5465 27361 5499
rect 27395 5465 27430 5499
rect 27464 5465 27499 5499
rect 27533 5465 27568 5499
rect 22812 5431 27568 5465
rect 16842 5355 16881 5389
rect 16915 5355 16954 5389
rect 16988 5355 17027 5389
rect 17061 5355 17100 5389
rect 17134 5355 17173 5389
rect 17207 5355 17246 5389
rect 17280 5355 17319 5389
rect 17353 5355 17392 5389
rect 17426 5355 17465 5389
rect 17499 5355 17538 5389
rect 17572 5355 17611 5389
rect 17645 5355 17684 5389
rect 17718 5355 17757 5389
rect 17791 5355 17830 5389
rect 17864 5355 17903 5389
rect 17937 5355 17976 5389
rect 18010 5355 18049 5389
rect 18083 5355 18122 5389
rect 18156 5355 18195 5389
rect 18229 5355 18268 5389
rect 18302 5355 18341 5389
rect 18375 5355 18414 5389
rect 18448 5355 18487 5389
rect 18521 5355 18560 5389
rect 18594 5355 18633 5389
rect 18667 5355 18705 5389
rect 18739 5355 18777 5389
rect 18811 5355 18849 5389
rect 18883 5355 18921 5389
rect 16808 5311 18955 5355
rect 16842 5277 16881 5311
rect 16915 5277 16954 5311
rect 16988 5277 17027 5311
rect 17061 5277 17100 5311
rect 17134 5277 17173 5311
rect 17207 5277 17246 5311
rect 17280 5277 17319 5311
rect 17353 5277 17392 5311
rect 17426 5277 17465 5311
rect 17499 5277 17538 5311
rect 17572 5277 17611 5311
rect 17645 5277 17684 5311
rect 17718 5277 17757 5311
rect 17791 5277 17830 5311
rect 17864 5277 17903 5311
rect 17937 5277 17976 5311
rect 18010 5277 18049 5311
rect 18083 5277 18122 5311
rect 18156 5277 18195 5311
rect 18229 5277 18268 5311
rect 18302 5277 18341 5311
rect 18375 5277 18414 5311
rect 18448 5277 18487 5311
rect 18521 5277 18560 5311
rect 18594 5277 18633 5311
rect 18667 5277 18705 5311
rect 18739 5277 18777 5311
rect 18811 5277 18849 5311
rect 18883 5277 18921 5311
rect 16808 5276 18955 5277
rect 19955 5399 20482 5423
rect 20125 5365 20167 5399
rect 20201 5365 20247 5399
rect 20281 5365 20327 5399
rect 20361 5365 20407 5399
rect 20441 5365 20482 5399
rect 20125 5331 20482 5365
rect 20125 5297 20167 5331
rect 20201 5297 20247 5331
rect 20281 5297 20327 5331
rect 20361 5297 20407 5331
rect 20441 5297 20482 5331
rect 20125 5263 20482 5297
rect 20125 5229 20167 5263
rect 20201 5229 20247 5263
rect 20281 5229 20327 5263
rect 20361 5229 20407 5263
rect 20441 5229 20482 5263
rect 20125 5195 20482 5229
rect 20125 5161 20167 5195
rect 20201 5161 20247 5195
rect 20281 5161 20327 5195
rect 20361 5161 20407 5195
rect 20441 5161 20482 5195
rect 20125 5127 20482 5161
rect 20125 5093 20167 5127
rect 20201 5093 20247 5127
rect 20281 5093 20327 5127
rect 20361 5093 20407 5127
rect 20441 5093 20482 5127
rect 22812 5421 26740 5431
rect 22812 5387 22836 5421
rect 22870 5387 22905 5421
rect 22939 5387 22974 5421
rect 23008 5387 23043 5421
rect 23077 5387 23112 5421
rect 23146 5387 23181 5421
rect 23215 5387 23250 5421
rect 23284 5387 23319 5421
rect 23353 5387 23388 5421
rect 23422 5387 23457 5421
rect 23491 5387 23526 5421
rect 23560 5387 23595 5421
rect 23629 5387 23664 5421
rect 23698 5387 23733 5421
rect 23767 5387 23802 5421
rect 23836 5387 23871 5421
rect 23905 5387 23940 5421
rect 23974 5387 24009 5421
rect 24043 5387 24078 5421
rect 24112 5387 24147 5421
rect 24181 5387 24216 5421
rect 24250 5387 24285 5421
rect 24319 5387 24354 5421
rect 24388 5387 24423 5421
rect 24457 5387 24492 5421
rect 24526 5387 24561 5421
rect 24595 5387 24630 5421
rect 24664 5387 24699 5421
rect 24733 5387 24768 5421
rect 24802 5387 24837 5421
rect 24871 5387 24906 5421
rect 24940 5387 24975 5421
rect 25009 5387 25044 5421
rect 25078 5387 25113 5421
rect 25147 5387 25181 5421
rect 25215 5387 25249 5421
rect 25283 5387 25317 5421
rect 25351 5387 25385 5421
rect 25419 5387 25453 5421
rect 25487 5387 25521 5421
rect 25555 5387 25589 5421
rect 25623 5387 25657 5421
rect 25691 5387 25725 5421
rect 25759 5387 25793 5421
rect 25827 5387 25861 5421
rect 25895 5387 25929 5421
rect 25963 5387 25997 5421
rect 26031 5387 26065 5421
rect 26099 5387 26133 5421
rect 26167 5387 26201 5421
rect 26235 5387 26269 5421
rect 26303 5387 26337 5421
rect 26371 5387 26405 5421
rect 26439 5387 26473 5421
rect 26507 5387 26541 5421
rect 26575 5387 26609 5421
rect 26643 5397 26740 5421
rect 26774 5397 26809 5431
rect 26843 5397 26878 5431
rect 26912 5397 26947 5431
rect 26981 5397 27016 5431
rect 27050 5397 27085 5431
rect 27119 5397 27154 5431
rect 27188 5397 27223 5431
rect 27257 5397 27292 5431
rect 27326 5397 27361 5431
rect 27395 5397 27430 5431
rect 27464 5397 27499 5431
rect 27533 5397 27568 5431
rect 26643 5387 27568 5397
rect 22812 5363 27568 5387
rect 22812 5343 26740 5363
rect 22812 5309 22836 5343
rect 22870 5309 22905 5343
rect 22939 5309 22974 5343
rect 23008 5309 23043 5343
rect 23077 5309 23112 5343
rect 23146 5309 23181 5343
rect 23215 5309 23250 5343
rect 23284 5309 23319 5343
rect 23353 5309 23388 5343
rect 23422 5309 23457 5343
rect 23491 5309 23526 5343
rect 23560 5309 23595 5343
rect 23629 5309 23664 5343
rect 23698 5309 23733 5343
rect 23767 5309 23802 5343
rect 23836 5309 23871 5343
rect 23905 5309 23940 5343
rect 23974 5309 24009 5343
rect 24043 5309 24078 5343
rect 24112 5309 24147 5343
rect 24181 5309 24216 5343
rect 24250 5309 24285 5343
rect 24319 5309 24354 5343
rect 24388 5309 24423 5343
rect 24457 5309 24492 5343
rect 24526 5309 24561 5343
rect 24595 5309 24630 5343
rect 24664 5309 24699 5343
rect 24733 5309 24768 5343
rect 24802 5309 24837 5343
rect 24871 5309 24906 5343
rect 24940 5309 24975 5343
rect 25009 5309 25044 5343
rect 25078 5309 25113 5343
rect 25147 5309 25181 5343
rect 25215 5309 25249 5343
rect 25283 5309 25317 5343
rect 25351 5309 25385 5343
rect 25419 5309 25453 5343
rect 25487 5309 25521 5343
rect 25555 5309 25589 5343
rect 25623 5309 25657 5343
rect 25691 5309 25725 5343
rect 25759 5309 25793 5343
rect 25827 5309 25861 5343
rect 25895 5309 25929 5343
rect 25963 5309 25997 5343
rect 26031 5309 26065 5343
rect 26099 5309 26133 5343
rect 26167 5309 26201 5343
rect 26235 5309 26269 5343
rect 26303 5309 26337 5343
rect 26371 5309 26405 5343
rect 26439 5309 26473 5343
rect 26507 5309 26541 5343
rect 26575 5309 26609 5343
rect 26643 5329 26740 5343
rect 26774 5329 26809 5363
rect 26843 5329 26878 5363
rect 26912 5329 26947 5363
rect 26981 5329 27016 5363
rect 27050 5329 27085 5363
rect 27119 5329 27154 5363
rect 27188 5329 27223 5363
rect 27257 5329 27292 5363
rect 27326 5329 27361 5363
rect 27395 5329 27430 5363
rect 27464 5329 27499 5363
rect 27533 5329 27568 5363
rect 26643 5309 27568 5329
rect 22812 5295 27568 5309
rect 22812 5265 26740 5295
rect 22812 5231 22836 5265
rect 22870 5231 22905 5265
rect 22939 5231 22974 5265
rect 23008 5231 23043 5265
rect 23077 5231 23112 5265
rect 23146 5231 23181 5265
rect 23215 5231 23250 5265
rect 23284 5231 23319 5265
rect 23353 5231 23388 5265
rect 23422 5231 23457 5265
rect 23491 5231 23526 5265
rect 23560 5231 23595 5265
rect 23629 5231 23664 5265
rect 23698 5231 23733 5265
rect 23767 5231 23802 5265
rect 23836 5231 23871 5265
rect 23905 5231 23940 5265
rect 23974 5231 24009 5265
rect 24043 5231 24078 5265
rect 24112 5231 24147 5265
rect 24181 5231 24216 5265
rect 24250 5231 24285 5265
rect 24319 5231 24354 5265
rect 24388 5231 24423 5265
rect 24457 5231 24492 5265
rect 24526 5231 24561 5265
rect 24595 5231 24630 5265
rect 24664 5231 24699 5265
rect 24733 5231 24768 5265
rect 24802 5231 24837 5265
rect 24871 5231 24906 5265
rect 24940 5231 24975 5265
rect 25009 5231 25044 5265
rect 25078 5231 25113 5265
rect 25147 5231 25181 5265
rect 25215 5231 25249 5265
rect 25283 5231 25317 5265
rect 25351 5231 25385 5265
rect 25419 5231 25453 5265
rect 25487 5231 25521 5265
rect 25555 5231 25589 5265
rect 25623 5231 25657 5265
rect 25691 5231 25725 5265
rect 25759 5231 25793 5265
rect 25827 5231 25861 5265
rect 25895 5231 25929 5265
rect 25963 5231 25997 5265
rect 26031 5231 26065 5265
rect 26099 5231 26133 5265
rect 26167 5231 26201 5265
rect 26235 5231 26269 5265
rect 26303 5231 26337 5265
rect 26371 5231 26405 5265
rect 26439 5231 26473 5265
rect 26507 5231 26541 5265
rect 26575 5231 26609 5265
rect 26643 5261 26740 5265
rect 26774 5261 26809 5295
rect 26843 5261 26878 5295
rect 26912 5261 26947 5295
rect 26981 5261 27016 5295
rect 27050 5261 27085 5295
rect 27119 5261 27154 5295
rect 27188 5261 27223 5295
rect 27257 5261 27292 5295
rect 27326 5261 27361 5295
rect 27395 5261 27430 5295
rect 27464 5261 27499 5295
rect 27533 5261 27568 5295
rect 26643 5231 27568 5261
rect 22812 5227 27568 5231
rect 22812 5193 26740 5227
rect 26774 5193 26809 5227
rect 26843 5193 26878 5227
rect 26912 5193 26947 5227
rect 26981 5193 27016 5227
rect 27050 5193 27085 5227
rect 27119 5193 27154 5227
rect 27188 5193 27223 5227
rect 27257 5193 27292 5227
rect 27326 5193 27361 5227
rect 27395 5193 27430 5227
rect 27464 5193 27499 5227
rect 27533 5193 27568 5227
rect 22812 5187 27568 5193
rect 22812 5153 22836 5187
rect 22870 5153 22905 5187
rect 22939 5153 22974 5187
rect 23008 5153 23043 5187
rect 23077 5153 23112 5187
rect 23146 5153 23181 5187
rect 23215 5153 23250 5187
rect 23284 5153 23319 5187
rect 23353 5153 23388 5187
rect 23422 5153 23457 5187
rect 23491 5153 23526 5187
rect 23560 5153 23595 5187
rect 23629 5153 23664 5187
rect 23698 5153 23733 5187
rect 23767 5153 23802 5187
rect 23836 5153 23871 5187
rect 23905 5153 23940 5187
rect 23974 5153 24009 5187
rect 24043 5153 24078 5187
rect 24112 5153 24147 5187
rect 24181 5153 24216 5187
rect 24250 5153 24285 5187
rect 24319 5153 24354 5187
rect 24388 5153 24423 5187
rect 24457 5153 24492 5187
rect 24526 5153 24561 5187
rect 24595 5153 24630 5187
rect 24664 5153 24699 5187
rect 24733 5153 24768 5187
rect 24802 5153 24837 5187
rect 24871 5153 24906 5187
rect 24940 5153 24975 5187
rect 25009 5153 25044 5187
rect 25078 5153 25113 5187
rect 25147 5153 25181 5187
rect 25215 5153 25249 5187
rect 25283 5153 25317 5187
rect 25351 5153 25385 5187
rect 25419 5153 25453 5187
rect 25487 5153 25521 5187
rect 25555 5153 25589 5187
rect 25623 5153 25657 5187
rect 25691 5153 25725 5187
rect 25759 5153 25793 5187
rect 25827 5153 25861 5187
rect 25895 5153 25929 5187
rect 25963 5153 25997 5187
rect 26031 5153 26065 5187
rect 26099 5153 26133 5187
rect 26167 5153 26201 5187
rect 26235 5153 26269 5187
rect 26303 5153 26337 5187
rect 26371 5153 26405 5187
rect 26439 5153 26473 5187
rect 26507 5153 26541 5187
rect 26575 5153 26609 5187
rect 26643 5159 27568 5187
rect 26643 5153 26740 5159
rect 22812 5125 26740 5153
rect 26774 5125 26809 5159
rect 26843 5125 26878 5159
rect 26912 5125 26947 5159
rect 26981 5125 27016 5159
rect 27050 5125 27085 5159
rect 27119 5125 27154 5159
rect 27188 5125 27223 5159
rect 27257 5125 27292 5159
rect 27326 5125 27361 5159
rect 27395 5125 27430 5159
rect 27464 5125 27499 5159
rect 27533 5125 27568 5159
rect 28690 5465 28777 5499
rect 28811 5465 28847 5499
rect 28881 5465 28917 5499
rect 28951 5465 28987 5499
rect 29021 5465 29057 5499
rect 29091 5465 29127 5499
rect 29161 5465 29197 5499
rect 29231 5465 29267 5499
rect 29301 5465 29337 5499
rect 29371 5465 29407 5499
rect 29441 5465 29477 5499
rect 29511 5465 29547 5499
rect 29581 5465 29617 5499
rect 29651 5465 29687 5499
rect 29721 5465 29757 5499
rect 29791 5465 29827 5499
rect 29861 5465 29896 5499
rect 29930 5465 29965 5499
rect 29999 5465 30034 5499
rect 30068 5465 30103 5499
rect 30137 5465 30172 5499
rect 30206 5465 30230 5499
rect 28690 5431 30230 5465
rect 28690 5397 28777 5431
rect 28811 5397 28847 5431
rect 28881 5397 28917 5431
rect 28951 5397 28987 5431
rect 29021 5397 29057 5431
rect 29091 5397 29127 5431
rect 29161 5397 29197 5431
rect 29231 5397 29267 5431
rect 29301 5397 29337 5431
rect 29371 5397 29407 5431
rect 29441 5397 29477 5431
rect 29511 5397 29547 5431
rect 29581 5397 29617 5431
rect 29651 5397 29687 5431
rect 29721 5397 29757 5431
rect 29791 5397 29827 5431
rect 29861 5397 29896 5431
rect 29930 5397 29965 5431
rect 29999 5397 30034 5431
rect 30068 5397 30103 5431
rect 30137 5397 30172 5431
rect 30206 5397 30230 5431
rect 28690 5363 30230 5397
rect 28690 5329 28777 5363
rect 28811 5329 28847 5363
rect 28881 5329 28917 5363
rect 28951 5329 28987 5363
rect 29021 5329 29057 5363
rect 29091 5329 29127 5363
rect 29161 5329 29197 5363
rect 29231 5329 29267 5363
rect 29301 5329 29337 5363
rect 29371 5329 29407 5363
rect 29441 5329 29477 5363
rect 29511 5329 29547 5363
rect 29581 5329 29617 5363
rect 29651 5329 29687 5363
rect 29721 5329 29757 5363
rect 29791 5329 29827 5363
rect 29861 5329 29896 5363
rect 29930 5329 29965 5363
rect 29999 5329 30034 5363
rect 30068 5329 30103 5363
rect 30137 5329 30172 5363
rect 30206 5329 30230 5363
rect 28690 5295 30230 5329
rect 28690 5261 28777 5295
rect 28811 5261 28847 5295
rect 28881 5261 28917 5295
rect 28951 5261 28987 5295
rect 29021 5261 29057 5295
rect 29091 5261 29127 5295
rect 29161 5261 29197 5295
rect 29231 5261 29267 5295
rect 29301 5261 29337 5295
rect 29371 5261 29407 5295
rect 29441 5261 29477 5295
rect 29511 5261 29547 5295
rect 29581 5261 29617 5295
rect 29651 5261 29687 5295
rect 29721 5261 29757 5295
rect 29791 5261 29827 5295
rect 29861 5261 29896 5295
rect 29930 5261 29965 5295
rect 29999 5261 30034 5295
rect 30068 5261 30103 5295
rect 30137 5261 30172 5295
rect 30206 5261 30230 5295
rect 28690 5227 30230 5261
rect 28690 5193 28777 5227
rect 28811 5193 28847 5227
rect 28881 5193 28917 5227
rect 28951 5193 28987 5227
rect 29021 5193 29057 5227
rect 29091 5193 29127 5227
rect 29161 5193 29197 5227
rect 29231 5193 29267 5227
rect 29301 5193 29337 5227
rect 29371 5193 29407 5227
rect 29441 5193 29477 5227
rect 29511 5193 29547 5227
rect 29581 5193 29617 5227
rect 29651 5193 29687 5227
rect 29721 5193 29757 5227
rect 29791 5193 29827 5227
rect 29861 5193 29896 5227
rect 29930 5193 29965 5227
rect 29999 5193 30034 5227
rect 30068 5193 30103 5227
rect 30137 5193 30172 5227
rect 30206 5193 30230 5227
rect 28690 5159 30230 5193
rect 22812 5116 27568 5125
rect 20125 5059 20482 5093
rect 20125 5025 20167 5059
rect 20201 5025 20247 5059
rect 20281 5025 20327 5059
rect 20361 5025 20407 5059
rect 20441 5025 20482 5059
rect 20125 4991 20482 5025
rect 20125 4957 20167 4991
rect 20201 4957 20247 4991
rect 20281 4957 20327 4991
rect 20361 4957 20407 4991
rect 20441 4957 20482 4991
rect 20125 4923 20482 4957
rect 20125 4889 20167 4923
rect 20201 4889 20247 4923
rect 20281 4889 20327 4923
rect 20361 4889 20407 4923
rect 20441 4889 20482 4923
rect 20125 4855 20482 4889
rect 20125 4821 20167 4855
rect 20201 4821 20247 4855
rect 20281 4821 20327 4855
rect 20361 4821 20407 4855
rect 20441 4821 20482 4855
rect 20125 4787 20482 4821
rect 20125 4753 20167 4787
rect 20201 4753 20247 4787
rect 20281 4753 20327 4787
rect 20361 4753 20407 4787
rect 20441 4753 20482 4787
rect 20125 4719 20482 4753
rect 20125 4685 20167 4719
rect 20201 4685 20247 4719
rect 20281 4685 20327 4719
rect 20361 4685 20407 4719
rect 20441 4685 20482 4719
rect 20125 4651 20482 4685
rect 20125 4617 20167 4651
rect 20201 4617 20247 4651
rect 20281 4617 20327 4651
rect 20361 4617 20407 4651
rect 20441 4617 20482 4651
rect 20125 4583 20482 4617
rect 20125 4549 20167 4583
rect 20201 4549 20247 4583
rect 20281 4549 20327 4583
rect 20361 4549 20407 4583
rect 20441 4549 20482 4583
rect 20125 4515 20482 4549
rect 20125 4481 20167 4515
rect 20201 4481 20247 4515
rect 20281 4481 20327 4515
rect 20361 4481 20407 4515
rect 20441 4481 20482 4515
rect 20125 4447 20482 4481
rect 20125 4413 20167 4447
rect 20201 4413 20247 4447
rect 20281 4413 20327 4447
rect 20361 4413 20407 4447
rect 20441 4413 20482 4447
rect 20125 4379 20482 4413
rect 20125 4345 20167 4379
rect 20201 4345 20247 4379
rect 20281 4345 20327 4379
rect 20361 4345 20407 4379
rect 20441 4345 20482 4379
rect 20125 4311 20482 4345
rect 20125 4277 20167 4311
rect 20201 4277 20247 4311
rect 20281 4277 20327 4311
rect 20361 4277 20407 4311
rect 20441 4277 20482 4311
rect 20125 4243 20482 4277
rect 20125 4209 20167 4243
rect 20201 4209 20247 4243
rect 20281 4209 20327 4243
rect 20361 4209 20407 4243
rect 20441 4209 20482 4243
rect 19955 4185 20482 4209
rect 20165 4175 20482 4185
rect 20165 4141 20167 4175
rect 20201 4141 20247 4175
rect 20281 4141 20327 4175
rect 20361 4141 20407 4175
rect 20441 4141 20482 4175
rect 26667 5091 27568 5116
rect 28690 5125 28777 5159
rect 28811 5125 28847 5159
rect 28881 5125 28917 5159
rect 28951 5125 28987 5159
rect 29021 5125 29057 5159
rect 29091 5125 29127 5159
rect 29161 5125 29197 5159
rect 29231 5125 29267 5159
rect 29301 5125 29337 5159
rect 29371 5125 29407 5159
rect 29441 5125 29477 5159
rect 29511 5125 29547 5159
rect 29581 5125 29617 5159
rect 29651 5125 29687 5159
rect 29721 5125 29757 5159
rect 29791 5125 29827 5159
rect 29861 5125 29896 5159
rect 29930 5125 29965 5159
rect 29999 5125 30034 5159
rect 30068 5125 30103 5159
rect 30137 5125 30172 5159
rect 30206 5125 30230 5159
rect 26667 5057 26740 5091
rect 26774 5057 26809 5091
rect 26843 5057 26878 5091
rect 26912 5057 26947 5091
rect 26981 5057 27016 5091
rect 27050 5057 27085 5091
rect 27119 5057 27154 5091
rect 27188 5057 27223 5091
rect 27257 5057 27292 5091
rect 27326 5057 27361 5091
rect 27395 5057 27430 5091
rect 27464 5057 27499 5091
rect 27533 5057 27568 5091
rect 28690 5091 30230 5125
rect 26667 5023 27568 5057
rect 28690 5057 28777 5091
rect 28811 5057 28847 5091
rect 28881 5057 28917 5091
rect 28951 5057 28987 5091
rect 29021 5057 29057 5091
rect 29091 5057 29127 5091
rect 29161 5057 29197 5091
rect 29231 5057 29267 5091
rect 29301 5057 29337 5091
rect 29371 5057 29407 5091
rect 29441 5057 29477 5091
rect 29511 5057 29547 5091
rect 29581 5057 29617 5091
rect 29651 5057 29687 5091
rect 29721 5057 29757 5091
rect 29791 5057 29827 5091
rect 29861 5057 29896 5091
rect 29930 5057 29965 5091
rect 29999 5057 30034 5091
rect 30068 5057 30103 5091
rect 30137 5057 30172 5091
rect 30206 5057 30230 5091
rect 26667 4989 26740 5023
rect 26774 4989 26809 5023
rect 26843 4989 26878 5023
rect 26912 4989 26947 5023
rect 26981 4989 27016 5023
rect 27050 4989 27085 5023
rect 27119 4989 27154 5023
rect 27188 4989 27223 5023
rect 27257 4989 27292 5023
rect 27326 4989 27361 5023
rect 27395 4989 27430 5023
rect 27464 4989 27499 5023
rect 27533 4989 27568 5023
rect 26667 4955 27568 4989
rect 28690 5023 30230 5057
rect 28690 4989 28777 5023
rect 28811 4989 28847 5023
rect 28881 4989 28917 5023
rect 28951 4989 28987 5023
rect 29021 4989 29057 5023
rect 29091 4989 29127 5023
rect 29161 4989 29197 5023
rect 29231 4989 29267 5023
rect 29301 4989 29337 5023
rect 29371 4989 29407 5023
rect 29441 4989 29477 5023
rect 29511 4989 29547 5023
rect 29581 4989 29617 5023
rect 29651 4989 29687 5023
rect 29721 4989 29757 5023
rect 29791 4989 29827 5023
rect 29861 4989 29896 5023
rect 29930 4989 29965 5023
rect 29999 4989 30034 5023
rect 30068 4989 30103 5023
rect 30137 4989 30172 5023
rect 30206 4989 30230 5023
rect 26667 4921 26740 4955
rect 26774 4921 26809 4955
rect 26843 4921 26878 4955
rect 26912 4921 26947 4955
rect 26981 4921 27016 4955
rect 27050 4921 27085 4955
rect 27119 4921 27154 4955
rect 27188 4921 27223 4955
rect 27257 4921 27292 4955
rect 27326 4921 27361 4955
rect 27395 4921 27430 4955
rect 27464 4921 27499 4955
rect 27533 4921 27568 4955
rect 28690 4955 30230 4989
rect 26667 4887 27568 4921
rect 28690 4921 28777 4955
rect 28811 4921 28847 4955
rect 28881 4921 28917 4955
rect 28951 4921 28987 4955
rect 29021 4921 29057 4955
rect 29091 4921 29127 4955
rect 29161 4921 29197 4955
rect 29231 4921 29267 4955
rect 29301 4921 29337 4955
rect 29371 4921 29407 4955
rect 29441 4921 29477 4955
rect 29511 4921 29547 4955
rect 29581 4921 29617 4955
rect 29651 4921 29687 4955
rect 29721 4921 29757 4955
rect 29791 4921 29827 4955
rect 29861 4921 29896 4955
rect 29930 4921 29965 4955
rect 29999 4921 30034 4955
rect 30068 4921 30103 4955
rect 30137 4921 30172 4955
rect 30206 4921 30230 4955
rect 26667 4853 26740 4887
rect 26774 4853 26809 4887
rect 26843 4853 26878 4887
rect 26912 4853 26947 4887
rect 26981 4853 27016 4887
rect 27050 4853 27085 4887
rect 27119 4853 27154 4887
rect 27188 4853 27223 4887
rect 27257 4853 27292 4887
rect 27326 4853 27361 4887
rect 27395 4853 27430 4887
rect 27464 4853 27499 4887
rect 27533 4853 27568 4887
rect 28690 4887 30230 4921
rect 26667 4819 27568 4853
rect 28690 4853 28777 4887
rect 28811 4853 28847 4887
rect 28881 4853 28917 4887
rect 28951 4853 28987 4887
rect 29021 4853 29057 4887
rect 29091 4853 29127 4887
rect 29161 4853 29197 4887
rect 29231 4853 29267 4887
rect 29301 4853 29337 4887
rect 29371 4853 29407 4887
rect 29441 4853 29477 4887
rect 29511 4853 29547 4887
rect 29581 4853 29617 4887
rect 29651 4853 29687 4887
rect 29721 4853 29757 4887
rect 29791 4853 29827 4887
rect 29861 4853 29896 4887
rect 29930 4853 29965 4887
rect 29999 4853 30034 4887
rect 30068 4853 30103 4887
rect 30137 4853 30172 4887
rect 30206 4853 30230 4887
rect 26667 4785 26740 4819
rect 26774 4785 26809 4819
rect 26843 4785 26878 4819
rect 26912 4785 26947 4819
rect 26981 4785 27016 4819
rect 27050 4785 27085 4819
rect 27119 4785 27154 4819
rect 27188 4785 27223 4819
rect 27257 4785 27292 4819
rect 27326 4785 27361 4819
rect 27395 4785 27430 4819
rect 27464 4785 27499 4819
rect 27533 4785 27568 4819
rect 28690 4819 30230 4853
rect 26667 4751 27568 4785
rect 26667 4717 26740 4751
rect 26774 4717 26809 4751
rect 26843 4717 26878 4751
rect 26912 4717 26947 4751
rect 26981 4717 27016 4751
rect 27050 4717 27085 4751
rect 27119 4717 27154 4751
rect 27188 4717 27223 4751
rect 27257 4717 27292 4751
rect 27326 4717 27361 4751
rect 27395 4717 27430 4751
rect 27464 4717 27499 4751
rect 27533 4717 27568 4751
rect 28690 4785 28777 4819
rect 28811 4785 28847 4819
rect 28881 4785 28917 4819
rect 28951 4785 28987 4819
rect 29021 4785 29057 4819
rect 29091 4785 29127 4819
rect 29161 4785 29197 4819
rect 29231 4785 29267 4819
rect 29301 4785 29337 4819
rect 29371 4785 29407 4819
rect 29441 4785 29477 4819
rect 29511 4785 29547 4819
rect 29581 4785 29617 4819
rect 29651 4785 29687 4819
rect 29721 4785 29757 4819
rect 29791 4785 29827 4819
rect 29861 4785 29896 4819
rect 29930 4785 29965 4819
rect 29999 4785 30034 4819
rect 30068 4785 30103 4819
rect 30137 4785 30172 4819
rect 30206 4785 30230 4819
rect 28690 4751 30230 4785
rect 26667 4683 27568 4717
rect 28690 4717 28777 4751
rect 28811 4717 28847 4751
rect 28881 4717 28917 4751
rect 28951 4717 28987 4751
rect 29021 4717 29057 4751
rect 29091 4717 29127 4751
rect 29161 4717 29197 4751
rect 29231 4717 29267 4751
rect 29301 4717 29337 4751
rect 29371 4717 29407 4751
rect 29441 4717 29477 4751
rect 29511 4717 29547 4751
rect 29581 4717 29617 4751
rect 29651 4717 29687 4751
rect 29721 4717 29757 4751
rect 29791 4717 29827 4751
rect 29861 4717 29896 4751
rect 29930 4717 29965 4751
rect 29999 4717 30034 4751
rect 30068 4717 30103 4751
rect 30137 4717 30172 4751
rect 30206 4717 30230 4751
rect 26667 4649 26740 4683
rect 26774 4649 26809 4683
rect 26843 4649 26878 4683
rect 26912 4649 26947 4683
rect 26981 4649 27016 4683
rect 27050 4649 27085 4683
rect 27119 4649 27154 4683
rect 27188 4649 27223 4683
rect 27257 4649 27292 4683
rect 27326 4649 27361 4683
rect 27395 4649 27430 4683
rect 27464 4649 27499 4683
rect 27533 4649 27568 4683
rect 26667 4615 27568 4649
rect 26667 4581 26713 4615
rect 26774 4581 26788 4615
rect 26843 4581 26863 4615
rect 26912 4581 26938 4615
rect 26981 4581 27013 4615
rect 27050 4581 27085 4615
rect 27122 4581 27154 4615
rect 27197 4581 27223 4615
rect 27272 4581 27292 4615
rect 27346 4581 27361 4615
rect 27420 4581 27430 4615
rect 27494 4581 27499 4615
rect 27533 4581 27534 4615
rect 26667 4547 27568 4581
rect 26667 4535 26740 4547
rect 26774 4535 26809 4547
rect 26843 4535 26878 4547
rect 26912 4535 26947 4547
rect 26981 4535 27016 4547
rect 26667 4501 26713 4535
rect 26774 4513 26788 4535
rect 26843 4513 26863 4535
rect 26912 4513 26938 4535
rect 26981 4513 27013 4535
rect 27050 4513 27085 4547
rect 27119 4535 27154 4547
rect 27188 4535 27223 4547
rect 27257 4535 27292 4547
rect 27326 4535 27361 4547
rect 27395 4535 27430 4547
rect 27464 4535 27499 4547
rect 27122 4513 27154 4535
rect 27197 4513 27223 4535
rect 27272 4513 27292 4535
rect 27346 4513 27361 4535
rect 27420 4513 27430 4535
rect 27494 4513 27499 4535
rect 27533 4535 27568 4547
rect 27533 4513 27534 4535
rect 26747 4501 26788 4513
rect 26822 4501 26863 4513
rect 26897 4501 26938 4513
rect 26972 4501 27013 4513
rect 27047 4501 27088 4513
rect 27122 4501 27163 4513
rect 27197 4501 27238 4513
rect 27272 4501 27312 4513
rect 27346 4501 27386 4513
rect 27420 4501 27460 4513
rect 27494 4501 27534 4513
rect 26667 4479 27568 4501
rect 26667 4455 26740 4479
rect 26774 4455 26809 4479
rect 26843 4455 26878 4479
rect 26912 4455 26947 4479
rect 26981 4455 27016 4479
rect 26667 4421 26713 4455
rect 26774 4445 26788 4455
rect 26843 4445 26863 4455
rect 26912 4445 26938 4455
rect 26981 4445 27013 4455
rect 27050 4445 27085 4479
rect 27119 4455 27154 4479
rect 27188 4455 27223 4479
rect 27257 4455 27292 4479
rect 27326 4455 27361 4479
rect 27395 4455 27430 4479
rect 27464 4455 27499 4479
rect 27122 4445 27154 4455
rect 27197 4445 27223 4455
rect 27272 4445 27292 4455
rect 27346 4445 27361 4455
rect 27420 4445 27430 4455
rect 27494 4445 27499 4455
rect 27533 4455 27568 4479
rect 27533 4445 27534 4455
rect 26747 4421 26788 4445
rect 26822 4421 26863 4445
rect 26897 4421 26938 4445
rect 26972 4421 27013 4445
rect 27047 4421 27088 4445
rect 27122 4421 27163 4445
rect 27197 4421 27238 4445
rect 27272 4421 27312 4445
rect 27346 4421 27386 4445
rect 27420 4421 27460 4445
rect 27494 4421 27534 4445
rect 26667 4411 27568 4421
rect 26667 4377 26740 4411
rect 26774 4377 26809 4411
rect 26843 4377 26878 4411
rect 26912 4377 26947 4411
rect 26981 4377 27016 4411
rect 27050 4377 27085 4411
rect 27119 4377 27154 4411
rect 27188 4377 27223 4411
rect 27257 4377 27292 4411
rect 27326 4377 27361 4411
rect 27395 4377 27430 4411
rect 27464 4377 27499 4411
rect 27533 4377 27568 4411
rect 26667 4375 27568 4377
rect 26667 4341 26713 4375
rect 26747 4343 26788 4375
rect 26822 4343 26863 4375
rect 26897 4343 26938 4375
rect 26972 4343 27013 4375
rect 27047 4343 27088 4375
rect 27122 4343 27163 4375
rect 27197 4343 27238 4375
rect 27272 4343 27312 4375
rect 27346 4343 27386 4375
rect 27420 4343 27460 4375
rect 27494 4343 27534 4375
rect 26774 4341 26788 4343
rect 26843 4341 26863 4343
rect 26912 4341 26938 4343
rect 26981 4341 27013 4343
rect 26667 4309 26740 4341
rect 26774 4309 26809 4341
rect 26843 4309 26878 4341
rect 26912 4309 26947 4341
rect 26981 4309 27016 4341
rect 27050 4309 27085 4343
rect 27122 4341 27154 4343
rect 27197 4341 27223 4343
rect 27272 4341 27292 4343
rect 27346 4341 27361 4343
rect 27420 4341 27430 4343
rect 27494 4341 27499 4343
rect 27119 4309 27154 4341
rect 27188 4309 27223 4341
rect 27257 4309 27292 4341
rect 27326 4309 27361 4341
rect 27395 4309 27430 4341
rect 27464 4309 27499 4341
rect 27533 4341 27534 4343
rect 27533 4309 27568 4341
rect 26667 4295 27568 4309
rect 26667 4261 26713 4295
rect 26747 4275 26788 4295
rect 26822 4275 26863 4295
rect 26897 4275 26938 4295
rect 26972 4275 27013 4295
rect 27047 4275 27088 4295
rect 27122 4275 27163 4295
rect 27197 4275 27238 4295
rect 27272 4275 27312 4295
rect 27346 4275 27386 4295
rect 27420 4275 27460 4295
rect 27494 4275 27534 4295
rect 26774 4261 26788 4275
rect 26843 4261 26863 4275
rect 26912 4261 26938 4275
rect 26981 4261 27013 4275
rect 26667 4241 26740 4261
rect 26774 4241 26809 4261
rect 26843 4241 26878 4261
rect 26912 4241 26947 4261
rect 26981 4241 27016 4261
rect 27050 4241 27085 4275
rect 27122 4261 27154 4275
rect 27197 4261 27223 4275
rect 27272 4261 27292 4275
rect 27346 4261 27361 4275
rect 27420 4261 27430 4275
rect 27494 4261 27499 4275
rect 27119 4241 27154 4261
rect 27188 4241 27223 4261
rect 27257 4241 27292 4261
rect 27326 4241 27361 4261
rect 27395 4241 27430 4261
rect 27464 4241 27499 4261
rect 27533 4261 27534 4275
rect 27533 4241 27568 4261
rect 28690 4241 28714 4717
rect 26667 4215 28714 4241
rect 26667 4181 26713 4215
rect 26747 4181 26788 4215
rect 26822 4181 26863 4215
rect 26897 4181 26938 4215
rect 26972 4181 27013 4215
rect 27047 4181 27088 4215
rect 27122 4181 27163 4215
rect 27197 4181 27238 4215
rect 27272 4181 27312 4215
rect 27346 4181 27386 4215
rect 27420 4181 27460 4215
rect 27494 4181 27534 4215
rect 27568 4181 27608 4215
rect 27642 4181 27682 4215
rect 27716 4181 27756 4215
rect 27790 4200 28714 4215
rect 27790 4181 27910 4200
rect 26667 4169 27910 4181
rect 27872 4166 27910 4169
rect 27944 4166 27988 4200
rect 28022 4166 28066 4200
rect 28100 4166 28144 4200
rect 28178 4166 28222 4200
rect 28256 4166 28300 4200
rect 28334 4166 28378 4200
rect 28412 4166 28456 4200
rect 28490 4166 28534 4200
rect 28568 4166 28612 4200
rect 28646 4169 28714 4200
rect 28646 4166 28684 4169
rect 20165 4107 20482 4141
rect 20165 4073 20167 4107
rect 20201 4073 20247 4107
rect 20281 4073 20327 4107
rect 20361 4073 20407 4107
rect 20441 4073 20482 4107
rect 20165 4039 20482 4073
rect 20165 4005 20167 4039
rect 20201 4005 20247 4039
rect 20281 4005 20327 4039
rect 20361 4005 20407 4039
rect 20441 4005 20482 4039
rect 20165 3971 20482 4005
rect 20165 3937 20167 3971
rect 20201 3937 20247 3971
rect 20281 3937 20327 3971
rect 20361 3937 20407 3971
rect 20441 3937 20482 3971
rect 20165 3903 20482 3937
rect 20165 3869 20167 3903
rect 20201 3869 20247 3903
rect 20281 3869 20327 3903
rect 20361 3869 20407 3903
rect 20441 3869 20482 3903
rect 20165 3835 20482 3869
rect 20165 3801 20167 3835
rect 20201 3801 20247 3835
rect 20281 3801 20327 3835
rect 20361 3801 20407 3835
rect 20441 3801 20482 3835
rect 20165 3767 20482 3801
rect 20165 3733 20167 3767
rect 20201 3733 20247 3767
rect 20281 3733 20327 3767
rect 20361 3733 20407 3767
rect 20441 3733 20482 3767
rect 20165 3699 20482 3733
rect 20165 3665 20167 3699
rect 20201 3665 20247 3699
rect 20281 3665 20327 3699
rect 20361 3665 20407 3699
rect 20441 3665 20482 3699
rect 20165 3631 20482 3665
rect 20165 3597 20167 3631
rect 20201 3597 20247 3631
rect 20281 3597 20327 3631
rect 20361 3597 20407 3631
rect 20441 3597 20482 3631
rect 20165 3563 20482 3597
rect 20165 3529 20167 3563
rect 20201 3529 20247 3563
rect 20281 3529 20327 3563
rect 20361 3529 20407 3563
rect 20441 3529 20482 3563
rect 9055 3273 9109 3529
rect 9055 3235 9143 3273
rect 9055 1453 9109 3235
rect 9315 3273 9397 3529
rect 9281 3235 9397 3273
rect 9315 1453 9397 3235
rect 10687 3273 10769 3529
rect 10687 3235 10803 3273
rect 10687 1453 10769 3235
rect 10975 3273 11029 3529
rect 10941 3235 11029 3273
rect 10975 1453 11029 3235
rect 20165 3495 20482 3529
rect 20165 3461 20167 3495
rect 20201 3461 20247 3495
rect 20281 3461 20327 3495
rect 20361 3461 20407 3495
rect 20441 3461 20482 3495
rect 20165 3427 20482 3461
rect 20165 3393 20167 3427
rect 20201 3393 20247 3427
rect 20281 3393 20327 3427
rect 20361 3393 20407 3427
rect 20441 3393 20482 3427
rect 20165 3359 20482 3393
rect 20165 3325 20167 3359
rect 20201 3325 20247 3359
rect 20281 3325 20327 3359
rect 20361 3325 20407 3359
rect 20441 3325 20482 3359
rect 20165 3291 20482 3325
rect 20165 3257 20167 3291
rect 20201 3257 20247 3291
rect 20281 3257 20327 3291
rect 20361 3257 20407 3291
rect 20441 3257 20482 3291
rect 20165 3223 20482 3257
rect 20165 3189 20167 3223
rect 20201 3189 20247 3223
rect 20281 3189 20327 3223
rect 20361 3189 20407 3223
rect 20441 3189 20482 3223
rect 20165 3155 20482 3189
rect 20165 3121 20167 3155
rect 20201 3121 20247 3155
rect 20281 3121 20327 3155
rect 20361 3121 20407 3155
rect 20441 3121 20482 3155
rect 20165 3087 20482 3121
rect 20165 3053 20167 3087
rect 20201 3053 20247 3087
rect 20281 3053 20327 3087
rect 20361 3053 20407 3087
rect 20441 3053 20482 3087
rect 20165 3019 20482 3053
rect 20165 2985 20167 3019
rect 20201 2985 20247 3019
rect 20281 2985 20327 3019
rect 20361 2985 20407 3019
rect 20441 2985 20482 3019
rect 20165 2951 20482 2985
rect 20165 2917 20167 2951
rect 20201 2917 20247 2951
rect 20281 2917 20327 2951
rect 20361 2917 20407 2951
rect 20441 2917 20482 2951
rect 20165 2883 20482 2917
rect 20165 2849 20167 2883
rect 20201 2849 20247 2883
rect 20281 2849 20327 2883
rect 20361 2849 20407 2883
rect 20441 2849 20482 2883
rect 20165 2815 20482 2849
rect 20165 2781 20167 2815
rect 20201 2781 20247 2815
rect 20281 2781 20327 2815
rect 20361 2781 20407 2815
rect 20441 2781 20482 2815
rect 20165 2747 20482 2781
rect 20165 2713 20167 2747
rect 20201 2713 20247 2747
rect 20281 2713 20327 2747
rect 20361 2713 20407 2747
rect 20441 2713 20482 2747
rect 20165 2678 20482 2713
rect 20165 2644 20167 2678
rect 20201 2644 20247 2678
rect 20281 2644 20327 2678
rect 20361 2644 20407 2678
rect 20441 2644 20482 2678
rect 20165 2637 20482 2644
rect 22522 3049 22789 3073
rect 22522 3015 22559 3049
rect 22593 3015 22657 3049
rect 22691 3015 22755 3049
rect 22522 2977 22789 3015
rect 22522 2943 22559 2977
rect 22593 2943 22657 2977
rect 22691 2943 22755 2977
rect 22522 2904 22789 2943
rect 22522 2870 22559 2904
rect 22593 2870 22657 2904
rect 22691 2870 22755 2904
rect 22522 2831 22789 2870
rect 22522 2797 22559 2831
rect 22593 2797 22657 2831
rect 22691 2797 22755 2831
rect 22522 2758 22789 2797
rect 22522 2724 22559 2758
rect 22593 2724 22657 2758
rect 22691 2724 22755 2758
rect 22522 2685 22789 2724
rect 22522 2651 22559 2685
rect 22593 2651 22657 2685
rect 22691 2651 22755 2685
rect 22522 2637 22789 2651
rect 20165 2612 22789 2637
rect 20165 2585 22559 2612
rect 17164 2551 18172 2585
rect 18206 2551 18241 2585
rect 18275 2551 18310 2585
rect 18344 2551 18379 2585
rect 18413 2551 18448 2585
rect 18482 2551 18517 2585
rect 18551 2551 18586 2585
rect 18620 2551 18655 2585
rect 18689 2551 18724 2585
rect 18758 2551 18793 2585
rect 18827 2551 18861 2585
rect 18895 2551 18929 2585
rect 18963 2551 18997 2585
rect 19031 2551 19065 2585
rect 19099 2551 19133 2585
rect 19167 2551 19201 2585
rect 19235 2551 19269 2585
rect 19303 2551 19337 2585
rect 19371 2551 19405 2585
rect 19439 2551 19473 2585
rect 19507 2551 19541 2585
rect 19575 2551 19609 2585
rect 19643 2551 19677 2585
rect 19711 2551 19745 2585
rect 19779 2551 19813 2585
rect 19847 2551 19881 2585
rect 19915 2551 19949 2585
rect 19983 2551 20017 2585
rect 20051 2551 20085 2585
rect 20119 2551 20153 2585
rect 20187 2551 20221 2585
rect 20255 2551 20289 2585
rect 20323 2551 20357 2585
rect 20391 2551 20425 2585
rect 20459 2551 20493 2585
rect 20527 2551 20561 2585
rect 20595 2551 20629 2585
rect 20663 2551 20697 2585
rect 20731 2551 20765 2585
rect 20799 2551 20833 2585
rect 20867 2551 20901 2585
rect 20935 2551 20969 2585
rect 21003 2551 21037 2585
rect 21071 2551 21105 2585
rect 21139 2551 21173 2585
rect 21207 2551 21241 2585
rect 21275 2551 21309 2585
rect 21343 2551 21377 2585
rect 21411 2551 21445 2585
rect 21479 2551 21513 2585
rect 21547 2551 21581 2585
rect 21615 2551 21649 2585
rect 21683 2551 21717 2585
rect 21751 2551 21785 2585
rect 21819 2551 21853 2585
rect 21887 2551 21921 2585
rect 21955 2551 21989 2585
rect 22023 2551 22057 2585
rect 22091 2551 22125 2585
rect 22159 2551 22193 2585
rect 22227 2551 22261 2585
rect 22295 2551 22329 2585
rect 22363 2551 22397 2585
rect 22431 2551 22465 2585
rect 22499 2578 22559 2585
rect 22593 2578 22657 2612
rect 22691 2578 22755 2612
rect 22499 2551 22789 2578
rect 17164 2539 22789 2551
rect 17164 2515 22559 2539
rect 16523 2481 16579 2515
rect 16613 2481 16650 2515
rect 16684 2481 16721 2515
rect 16755 2481 16792 2515
rect 16826 2481 16863 2515
rect 16897 2481 16933 2515
rect 16967 2481 17003 2515
rect 17037 2481 17073 2515
rect 17107 2481 17143 2515
rect 17177 2481 17213 2515
rect 17247 2481 17283 2515
rect 17317 2481 17353 2515
rect 17387 2481 17423 2515
rect 17457 2481 17493 2515
rect 17527 2481 17563 2515
rect 17597 2481 17633 2515
rect 17667 2481 17703 2515
rect 17737 2481 17773 2515
rect 17807 2481 17843 2515
rect 17877 2481 17913 2515
rect 17947 2481 17983 2515
rect 18017 2481 18053 2515
rect 18087 2481 18172 2515
rect 18206 2481 18241 2515
rect 18275 2481 18310 2515
rect 18344 2481 18379 2515
rect 18413 2481 18448 2515
rect 18482 2481 18517 2515
rect 18551 2481 18586 2515
rect 18620 2481 18655 2515
rect 18689 2481 18724 2515
rect 18758 2481 18793 2515
rect 18827 2481 18861 2515
rect 18895 2481 18929 2515
rect 18963 2481 18997 2515
rect 19031 2481 19065 2515
rect 19099 2481 19133 2515
rect 19167 2481 19201 2515
rect 19235 2481 19269 2515
rect 19303 2481 19337 2515
rect 19371 2481 19405 2515
rect 19439 2481 19473 2515
rect 19507 2481 19541 2515
rect 19575 2481 19609 2515
rect 19643 2481 19677 2515
rect 19711 2481 19745 2515
rect 19779 2481 19813 2515
rect 19847 2481 19881 2515
rect 19915 2481 19949 2515
rect 19983 2481 20017 2515
rect 20051 2481 20085 2515
rect 20119 2481 20153 2515
rect 20187 2481 20221 2515
rect 20255 2481 20289 2515
rect 20323 2481 20357 2515
rect 20391 2481 20425 2515
rect 20459 2481 20493 2515
rect 20527 2481 20561 2515
rect 20595 2481 20629 2515
rect 20663 2481 20697 2515
rect 20731 2481 20765 2515
rect 20799 2481 20833 2515
rect 20867 2481 20901 2515
rect 20935 2481 20969 2515
rect 21003 2481 21037 2515
rect 21071 2481 21105 2515
rect 21139 2481 21173 2515
rect 21207 2481 21241 2515
rect 21275 2481 21309 2515
rect 21343 2481 21377 2515
rect 21411 2481 21445 2515
rect 21479 2481 21513 2515
rect 21547 2481 21581 2515
rect 21615 2481 21649 2515
rect 21683 2481 21717 2515
rect 21751 2481 21785 2515
rect 21819 2481 21853 2515
rect 21887 2481 21921 2515
rect 21955 2481 21989 2515
rect 22023 2481 22057 2515
rect 22091 2481 22125 2515
rect 22159 2481 22193 2515
rect 22227 2481 22261 2515
rect 22295 2481 22329 2515
rect 22363 2481 22397 2515
rect 22431 2481 22465 2515
rect 22499 2505 22559 2515
rect 22593 2505 22657 2539
rect 22691 2505 22755 2539
rect 22499 2481 22789 2505
rect 16523 2462 22789 2481
rect 16523 2446 22405 2462
rect 22275 2428 22405 2446
rect 22439 2428 22507 2462
rect 22541 2428 22609 2462
rect 22643 2428 22789 2462
rect 22275 2403 22789 2428
rect 22275 2369 22347 2403
rect 22381 2387 22415 2403
rect 22381 2369 22405 2387
rect 22449 2369 22483 2403
rect 22517 2387 22551 2403
rect 22541 2369 22551 2387
rect 22585 2387 22619 2403
rect 22585 2369 22609 2387
rect 22653 2369 22687 2403
rect 22721 2369 22755 2403
rect 22275 2353 22405 2369
rect 22439 2353 22507 2369
rect 22541 2353 22609 2369
rect 22643 2353 22789 2369
rect 22275 2328 22789 2353
rect 22275 2294 22347 2328
rect 22381 2312 22415 2328
rect 22381 2294 22405 2312
rect 22449 2294 22483 2328
rect 22517 2312 22551 2328
rect 22541 2294 22551 2312
rect 22585 2312 22619 2328
rect 22585 2294 22609 2312
rect 22653 2294 22687 2328
rect 22721 2294 22755 2328
rect 22275 2278 22405 2294
rect 22439 2278 22507 2294
rect 22541 2278 22609 2294
rect 22643 2278 22789 2294
rect 22275 2252 22789 2278
rect 22275 2218 22347 2252
rect 22381 2237 22415 2252
rect 22381 2218 22405 2237
rect 22449 2218 22483 2252
rect 22517 2237 22551 2252
rect 22541 2218 22551 2237
rect 22585 2237 22619 2252
rect 22585 2218 22609 2237
rect 22653 2218 22687 2252
rect 22721 2218 22755 2252
rect 22275 2203 22405 2218
rect 22439 2203 22507 2218
rect 22541 2203 22609 2218
rect 22643 2203 22789 2218
rect 22275 2176 22789 2203
rect 22275 2142 22347 2176
rect 22381 2162 22415 2176
rect 22381 2142 22405 2162
rect 22449 2142 22483 2176
rect 22517 2162 22551 2176
rect 22541 2142 22551 2162
rect 22585 2162 22619 2176
rect 22585 2142 22609 2162
rect 22653 2142 22687 2176
rect 22721 2142 22755 2176
rect 22275 2128 22405 2142
rect 22439 2128 22507 2142
rect 22541 2128 22609 2142
rect 22643 2128 22789 2142
rect 22275 2100 22789 2128
rect 22275 2066 22347 2100
rect 22381 2087 22415 2100
rect 22381 2066 22405 2087
rect 22449 2066 22483 2100
rect 22517 2087 22551 2100
rect 22541 2066 22551 2087
rect 22585 2087 22619 2100
rect 22585 2066 22609 2087
rect 22653 2066 22687 2100
rect 22721 2066 22755 2100
rect 22275 2053 22405 2066
rect 22439 2053 22507 2066
rect 22541 2053 22609 2066
rect 22643 2053 22789 2066
rect 22275 2024 22789 2053
rect 22275 1990 22347 2024
rect 22381 2012 22415 2024
rect 22381 1990 22405 2012
rect 22449 1990 22483 2024
rect 22517 2012 22551 2024
rect 22541 1990 22551 2012
rect 22585 2012 22619 2024
rect 22585 1990 22609 2012
rect 22653 1990 22687 2024
rect 22721 1990 22755 2024
rect 22275 1978 22405 1990
rect 22439 1978 22507 1990
rect 22541 1978 22609 1990
rect 22643 1978 22789 1990
rect 22275 1948 22789 1978
rect 22275 1914 22347 1948
rect 22381 1936 22415 1948
rect 22381 1914 22405 1936
rect 22449 1914 22483 1948
rect 22517 1936 22551 1948
rect 22541 1914 22551 1936
rect 22585 1936 22619 1948
rect 22585 1914 22609 1936
rect 22653 1914 22687 1948
rect 22721 1914 22755 1948
rect 22275 1902 22405 1914
rect 22439 1902 22507 1914
rect 22541 1902 22609 1914
rect 22643 1902 22789 1914
rect 22275 1872 22789 1902
rect 22275 1838 22347 1872
rect 22381 1860 22415 1872
rect 22381 1838 22405 1860
rect 22449 1838 22483 1872
rect 22517 1860 22551 1872
rect 22541 1838 22551 1860
rect 22585 1860 22619 1872
rect 22585 1838 22609 1860
rect 22653 1838 22687 1872
rect 22721 1838 22755 1872
rect 22275 1826 22405 1838
rect 22439 1826 22507 1838
rect 22541 1826 22609 1838
rect 22643 1826 22789 1838
rect 22275 1796 22789 1826
rect 22275 1762 22347 1796
rect 22381 1784 22415 1796
rect 22381 1762 22405 1784
rect 22449 1762 22483 1796
rect 22517 1784 22551 1796
rect 22541 1762 22551 1784
rect 22585 1784 22619 1796
rect 22585 1762 22609 1784
rect 22653 1762 22687 1796
rect 22721 1762 22755 1796
rect 22275 1750 22405 1762
rect 22439 1750 22507 1762
rect 22541 1750 22609 1762
rect 22643 1750 22789 1762
rect 22275 1738 22789 1750
rect 26722 2273 28392 2348
rect 26722 2239 26787 2273
rect 26821 2239 26858 2273
rect 26892 2239 26929 2273
rect 26963 2239 27000 2273
rect 27034 2239 27071 2273
rect 27105 2239 27142 2273
rect 27176 2239 27213 2273
rect 27247 2239 27284 2273
rect 27318 2239 27354 2273
rect 27388 2239 27424 2273
rect 27458 2239 27494 2273
rect 27528 2239 27564 2273
rect 27598 2239 27634 2273
rect 27668 2239 27704 2273
rect 27738 2239 27774 2273
rect 27808 2239 27844 2273
rect 27878 2239 27914 2273
rect 27948 2239 27984 2273
rect 28018 2239 28054 2273
rect 28088 2239 28124 2273
rect 28158 2239 28194 2273
rect 28228 2239 28264 2273
rect 28298 2239 28334 2273
rect 28368 2239 28392 2273
rect 26722 2205 28392 2239
rect 26722 2171 26787 2205
rect 26821 2171 26858 2205
rect 26892 2171 26929 2205
rect 26963 2171 27000 2205
rect 27034 2171 27071 2205
rect 27105 2171 27142 2205
rect 27176 2171 27213 2205
rect 27247 2171 27284 2205
rect 27318 2171 27354 2205
rect 27388 2171 27424 2205
rect 27458 2171 27494 2205
rect 27528 2171 27564 2205
rect 27598 2171 27634 2205
rect 27668 2171 27704 2205
rect 27738 2171 27774 2205
rect 27808 2171 27844 2205
rect 27878 2171 27914 2205
rect 27948 2171 27984 2205
rect 28018 2171 28054 2205
rect 28088 2171 28124 2205
rect 28158 2171 28194 2205
rect 28228 2171 28264 2205
rect 28298 2171 28334 2205
rect 28368 2171 28392 2205
rect 26722 2137 28392 2171
rect 26722 2103 26787 2137
rect 26821 2103 26858 2137
rect 26892 2103 26929 2137
rect 26963 2103 27000 2137
rect 27034 2103 27071 2137
rect 27105 2103 27142 2137
rect 27176 2103 27213 2137
rect 27247 2103 27284 2137
rect 27318 2103 27354 2137
rect 27388 2103 27424 2137
rect 27458 2103 27494 2137
rect 27528 2103 27564 2137
rect 27598 2103 27634 2137
rect 27668 2103 27704 2137
rect 27738 2103 27774 2137
rect 27808 2103 27844 2137
rect 27878 2103 27914 2137
rect 27948 2103 27984 2137
rect 28018 2103 28054 2137
rect 28088 2103 28124 2137
rect 28158 2103 28194 2137
rect 28228 2103 28264 2137
rect 28298 2103 28334 2137
rect 28368 2103 28392 2137
rect 26722 2069 28392 2103
rect 26722 2035 26787 2069
rect 26821 2035 26858 2069
rect 26892 2035 26929 2069
rect 26963 2035 27000 2069
rect 27034 2035 27071 2069
rect 27105 2035 27142 2069
rect 27176 2035 27213 2069
rect 27247 2035 27284 2069
rect 27318 2035 27354 2069
rect 27388 2035 27424 2069
rect 27458 2035 27494 2069
rect 27528 2035 27564 2069
rect 27598 2035 27634 2069
rect 27668 2035 27704 2069
rect 27738 2035 27774 2069
rect 27808 2035 27844 2069
rect 27878 2035 27914 2069
rect 27948 2035 27984 2069
rect 28018 2035 28054 2069
rect 28088 2035 28124 2069
rect 28158 2035 28194 2069
rect 28228 2035 28264 2069
rect 28298 2035 28334 2069
rect 28368 2035 28392 2069
rect 26722 2001 28392 2035
rect 26722 1967 26787 2001
rect 26821 1967 26858 2001
rect 26892 1967 26929 2001
rect 26963 1967 27000 2001
rect 27034 1967 27071 2001
rect 27105 1967 27142 2001
rect 27176 1967 27213 2001
rect 27247 1967 27284 2001
rect 27318 1967 27354 2001
rect 27388 1967 27424 2001
rect 27458 1967 27494 2001
rect 27528 1967 27564 2001
rect 27598 1967 27634 2001
rect 27668 1967 27704 2001
rect 27738 1967 27774 2001
rect 27808 1967 27844 2001
rect 27878 1967 27914 2001
rect 27948 1967 27984 2001
rect 28018 1967 28054 2001
rect 28088 1967 28124 2001
rect 28158 1967 28194 2001
rect 28228 1967 28264 2001
rect 28298 1967 28334 2001
rect 28368 1967 28392 2001
rect 26722 1933 28392 1967
rect 26722 1899 26787 1933
rect 26821 1899 26858 1933
rect 26892 1899 26929 1933
rect 26963 1899 27000 1933
rect 27034 1899 27071 1933
rect 27105 1899 27142 1933
rect 27176 1899 27213 1933
rect 27247 1899 27284 1933
rect 27318 1899 27354 1933
rect 27388 1899 27424 1933
rect 27458 1899 27494 1933
rect 27528 1899 27564 1933
rect 27598 1899 27634 1933
rect 27668 1899 27704 1933
rect 27738 1899 27774 1933
rect 27808 1899 27844 1933
rect 27878 1899 27914 1933
rect 27948 1899 27984 1933
rect 28018 1899 28054 1933
rect 28088 1899 28124 1933
rect 28158 1899 28194 1933
rect 28228 1899 28264 1933
rect 28298 1899 28334 1933
rect 28368 1899 28392 1933
rect 26722 1865 28392 1899
rect 26722 1831 26787 1865
rect 26821 1831 26858 1865
rect 26892 1831 26929 1865
rect 26963 1831 27000 1865
rect 27034 1831 27071 1865
rect 27105 1831 27142 1865
rect 27176 1831 27213 1865
rect 27247 1831 27284 1865
rect 27318 1831 27354 1865
rect 27388 1831 27424 1865
rect 27458 1831 27494 1865
rect 27528 1831 27564 1865
rect 27598 1831 27634 1865
rect 27668 1831 27704 1865
rect 27738 1831 27774 1865
rect 27808 1831 27844 1865
rect 27878 1831 27914 1865
rect 27948 1831 27984 1865
rect 28018 1831 28054 1865
rect 28088 1831 28124 1865
rect 28158 1831 28194 1865
rect 28228 1831 28264 1865
rect 28298 1831 28334 1865
rect 28368 1831 28392 1865
rect 26722 1797 28392 1831
rect 26722 1763 26787 1797
rect 26821 1763 26858 1797
rect 26892 1763 26929 1797
rect 26963 1763 27000 1797
rect 27034 1763 27071 1797
rect 27105 1763 27142 1797
rect 27176 1763 27213 1797
rect 27247 1763 27284 1797
rect 27318 1763 27354 1797
rect 27388 1763 27424 1797
rect 27458 1763 27494 1797
rect 27528 1763 27564 1797
rect 27598 1763 27634 1797
rect 27668 1763 27704 1797
rect 27738 1763 27774 1797
rect 27808 1763 27844 1797
rect 27878 1763 27914 1797
rect 27948 1763 27984 1797
rect 28018 1763 28054 1797
rect 28088 1763 28124 1797
rect 28158 1763 28194 1797
rect 28228 1763 28264 1797
rect 28298 1763 28334 1797
rect 28368 1763 28392 1797
rect 26722 1729 28392 1763
rect 26722 1695 26787 1729
rect 26821 1695 26858 1729
rect 26892 1695 26929 1729
rect 26963 1695 27000 1729
rect 27034 1695 27071 1729
rect 27105 1695 27142 1729
rect 27176 1695 27213 1729
rect 27247 1695 27284 1729
rect 27318 1695 27354 1729
rect 27388 1695 27424 1729
rect 27458 1695 27494 1729
rect 27528 1695 27564 1729
rect 27598 1695 27634 1729
rect 27668 1695 27704 1729
rect 27738 1695 27774 1729
rect 27808 1695 27844 1729
rect 27878 1695 27914 1729
rect 27948 1695 27984 1729
rect 28018 1695 28054 1729
rect 28088 1695 28124 1729
rect 28158 1695 28194 1729
rect 28228 1695 28264 1729
rect 28298 1695 28334 1729
rect 28368 1695 28392 1729
rect 26722 1643 26979 1695
rect 26722 1609 26753 1643
rect 26787 1609 26849 1643
rect 26883 1609 26945 1643
rect 26722 1571 26979 1609
rect 26722 1537 26753 1571
rect 26787 1537 26849 1571
rect 26883 1537 26945 1571
rect 26722 1499 26979 1537
rect 26722 1465 26753 1499
rect 26787 1465 26849 1499
rect 26883 1465 26945 1499
rect 26722 1426 26979 1465
rect 26722 1392 26753 1426
rect 26787 1392 26849 1426
rect 26883 1392 26945 1426
rect 26722 1353 26979 1392
rect 26722 1319 26753 1353
rect 26787 1319 26849 1353
rect 26883 1319 26945 1353
rect 26722 1280 26979 1319
rect 26722 1246 26753 1280
rect 26787 1246 26849 1280
rect 26883 1246 26945 1280
rect 26722 1207 26979 1246
rect 26722 1173 26753 1207
rect 26787 1173 26849 1207
rect 26883 1173 26945 1207
rect 26722 1134 26979 1173
rect 26722 1100 26753 1134
rect 26787 1100 26849 1134
rect 26883 1100 26945 1134
rect 26722 1061 26979 1100
rect 26722 1027 26753 1061
rect 26787 1027 26849 1061
rect 26883 1027 26945 1061
rect 26722 988 26979 1027
rect 26722 954 26753 988
rect 26787 954 26849 988
rect 26883 954 26945 988
rect 26722 915 26979 954
rect 26722 881 26753 915
rect 26787 881 26849 915
rect 26883 881 26945 915
rect 26722 831 26979 881
<< viali >>
rect 448 33062 626 41880
rect 448 32989 482 33023
rect 520 32989 554 33023
rect 592 32989 626 33023
rect 448 32916 482 32950
rect 520 32916 554 32950
rect 592 32916 626 32950
rect 448 32843 482 32877
rect 520 32843 554 32877
rect 592 32843 626 32877
rect 448 32770 482 32804
rect 520 32770 554 32804
rect 592 32770 626 32804
rect 448 32697 482 32731
rect 520 32697 554 32731
rect 592 32697 626 32731
rect 448 32624 482 32658
rect 520 32624 554 32658
rect 592 32624 626 32658
rect 448 32551 482 32585
rect 520 32551 554 32585
rect 592 32551 626 32585
rect 448 32478 482 32512
rect 520 32478 554 32512
rect 592 32478 626 32512
rect 448 32405 482 32439
rect 520 32405 554 32439
rect 592 32405 626 32439
rect 448 32332 482 32366
rect 520 32332 554 32366
rect 592 32332 626 32366
rect 448 32259 482 32293
rect 520 32259 554 32293
rect 592 32259 626 32293
rect 448 32186 482 32220
rect 520 32186 554 32220
rect 592 32186 626 32220
rect 448 32113 482 32147
rect 520 32113 554 32147
rect 592 32113 626 32147
rect 448 32040 482 32074
rect 520 32040 554 32074
rect 592 32040 626 32074
rect 448 31967 482 32001
rect 520 31967 554 32001
rect 592 31967 626 32001
rect 448 31894 482 31928
rect 520 31894 554 31928
rect 592 31894 626 31928
rect 448 31821 482 31855
rect 520 31821 554 31855
rect 592 31821 626 31855
rect 448 31748 482 31782
rect 520 31748 554 31782
rect 592 31748 626 31782
rect 448 31675 482 31709
rect 520 31675 554 31709
rect 592 31675 626 31709
rect 448 31602 482 31636
rect 520 31602 554 31636
rect 592 31602 626 31636
rect 448 31529 482 31563
rect 520 31529 554 31563
rect 592 31529 626 31563
rect 448 31456 482 31490
rect 520 31456 554 31490
rect 592 31456 626 31490
rect 448 31383 482 31417
rect 520 31383 554 31417
rect 592 31383 626 31417
rect 448 31310 482 31344
rect 520 31310 554 31344
rect 592 31310 626 31344
rect 448 31237 482 31271
rect 520 31237 554 31271
rect 592 31237 626 31271
rect 448 31164 482 31198
rect 520 31164 554 31198
rect 592 31164 626 31198
rect 448 31091 482 31125
rect 520 31091 554 31125
rect 592 31091 626 31125
rect 448 31018 482 31052
rect 520 31018 554 31052
rect 592 31018 626 31052
rect 448 30945 482 30979
rect 520 30945 554 30979
rect 592 30945 626 30979
rect 448 30872 482 30906
rect 520 30872 554 30906
rect 592 30872 626 30906
rect 448 30799 482 30833
rect 520 30799 554 30833
rect 592 30799 626 30833
rect 448 30726 482 30760
rect 520 30726 554 30760
rect 592 30726 626 30760
rect 448 30653 482 30687
rect 520 30653 554 30687
rect 592 30653 626 30687
rect 448 30580 482 30614
rect 520 30580 554 30614
rect 592 30580 626 30614
rect 448 30507 482 30541
rect 520 30507 554 30541
rect 592 30507 626 30541
rect 448 30434 482 30468
rect 520 30434 554 30468
rect 592 30434 626 30468
rect 448 30361 482 30395
rect 520 30361 554 30395
rect 592 30361 626 30395
rect 26916 31540 26950 31574
rect 26996 31540 27030 31574
rect 27076 31540 27110 31574
rect 27156 31540 27190 31574
rect 27236 31540 27270 31574
rect 26916 31467 26950 31501
rect 26996 31467 27030 31501
rect 27076 31467 27110 31501
rect 27156 31467 27190 31501
rect 27236 31467 27270 31501
rect 26916 31394 26950 31428
rect 26996 31394 27030 31428
rect 27076 31394 27110 31428
rect 27156 31394 27190 31428
rect 27236 31394 27270 31428
rect 26916 31321 26950 31355
rect 26996 31321 27030 31355
rect 27076 31321 27110 31355
rect 27156 31321 27190 31355
rect 27236 31321 27270 31355
rect 26916 31248 26950 31282
rect 26996 31248 27030 31282
rect 27076 31248 27110 31282
rect 27156 31248 27190 31282
rect 27236 31248 27270 31282
rect 26916 31175 26950 31209
rect 26996 31175 27030 31209
rect 27076 31175 27110 31209
rect 27156 31175 27190 31209
rect 27236 31175 27270 31209
rect 26916 31102 26950 31136
rect 26996 31102 27030 31136
rect 27076 31102 27110 31136
rect 27156 31102 27190 31136
rect 27236 31102 27270 31136
rect 26916 31029 26950 31063
rect 26996 31029 27030 31063
rect 27076 31029 27110 31063
rect 27156 31029 27190 31063
rect 27236 31029 27270 31063
rect 26916 30956 26950 30990
rect 26996 30956 27030 30990
rect 27076 30956 27110 30990
rect 27156 30956 27190 30990
rect 27236 30956 27270 30990
rect 26916 30883 26950 30917
rect 26996 30883 27030 30917
rect 27076 30883 27110 30917
rect 27156 30883 27190 30917
rect 27236 30883 27270 30917
rect 26916 30810 26950 30844
rect 26996 30810 27030 30844
rect 27076 30810 27110 30844
rect 27156 30810 27190 30844
rect 27236 30810 27270 30844
rect 26916 30737 26950 30771
rect 26996 30737 27030 30771
rect 27076 30737 27110 30771
rect 27156 30737 27190 30771
rect 27236 30737 27270 30771
rect 26916 30664 26950 30698
rect 26996 30664 27030 30698
rect 27076 30664 27110 30698
rect 27156 30664 27190 30698
rect 27236 30664 27270 30698
rect 26916 30591 26950 30625
rect 26996 30591 27030 30625
rect 27076 30591 27110 30625
rect 27156 30591 27190 30625
rect 27236 30591 27270 30625
rect 26916 30517 26950 30551
rect 26996 30517 27030 30551
rect 27076 30517 27110 30551
rect 27156 30517 27190 30551
rect 27236 30517 27270 30551
rect 26916 30443 26950 30477
rect 26996 30443 27030 30477
rect 27076 30443 27110 30477
rect 27156 30443 27190 30477
rect 27236 30443 27270 30477
rect 26916 30369 26950 30403
rect 26996 30369 27030 30403
rect 27076 30369 27110 30403
rect 27156 30369 27190 30403
rect 27236 30369 27270 30403
rect 26916 30295 26950 30329
rect 26996 30295 27030 30329
rect 27076 30295 27110 30329
rect 27156 30295 27190 30329
rect 27236 30295 27270 30329
rect 439 30241 473 30275
rect 579 30241 613 30275
rect 439 30169 473 30203
rect 579 30169 613 30203
rect 439 30097 473 30131
rect 579 30097 613 30131
rect 439 30025 473 30059
rect 579 30025 613 30059
rect 439 29953 473 29987
rect 579 29953 613 29987
rect 439 29881 473 29915
rect 579 29881 613 29915
rect 439 29809 473 29843
rect 579 29809 613 29843
rect 439 29737 473 29771
rect 579 29737 613 29771
rect 439 29665 473 29699
rect 579 29665 613 29699
rect 439 29593 473 29627
rect 579 29593 613 29627
rect 439 29521 473 29555
rect 579 29521 613 29555
rect 439 29449 473 29483
rect 579 29449 613 29483
rect 439 29377 473 29411
rect 579 29377 613 29411
rect 439 29305 473 29339
rect 579 29305 613 29339
rect 439 29233 473 29267
rect 579 29233 613 29267
rect 439 29161 473 29195
rect 579 29161 613 29195
rect 439 29089 473 29123
rect 579 29089 613 29123
rect 439 29017 473 29051
rect 579 29017 613 29051
rect 439 28945 473 28979
rect 579 28945 613 28979
rect 439 28873 473 28907
rect 579 28873 613 28907
rect 439 28801 473 28835
rect 579 28801 613 28835
rect 439 28729 473 28763
rect 579 28729 613 28763
rect 439 28657 473 28691
rect 579 28657 613 28691
rect 439 28585 473 28619
rect 579 28585 613 28619
rect 439 28513 473 28547
rect 579 28513 613 28547
rect 26916 30221 26950 30255
rect 26996 30221 27030 30255
rect 27076 30221 27110 30255
rect 27156 30221 27190 30255
rect 27236 30221 27270 30255
rect 26916 30147 26950 30181
rect 26996 30147 27030 30181
rect 27076 30147 27110 30181
rect 27156 30147 27190 30181
rect 27236 30147 27270 30181
rect 26916 30073 26950 30107
rect 26996 30073 27030 30107
rect 27076 30073 27110 30107
rect 27156 30073 27190 30107
rect 27236 30073 27270 30107
rect 26916 29999 26950 30033
rect 26996 29999 27030 30033
rect 27076 29999 27110 30033
rect 27156 29999 27190 30033
rect 27236 29999 27270 30033
rect 26916 29925 26950 29959
rect 26996 29925 27030 29959
rect 27076 29925 27110 29959
rect 27156 29925 27190 29959
rect 27236 29925 27270 29959
rect 26916 29851 26950 29885
rect 26996 29851 27030 29885
rect 27076 29851 27110 29885
rect 27156 29851 27190 29885
rect 27236 29851 27270 29885
rect 26916 29777 26950 29811
rect 26996 29777 27030 29811
rect 27076 29777 27110 29811
rect 27156 29777 27190 29811
rect 27236 29777 27270 29811
rect 26916 29703 26950 29737
rect 26996 29703 27030 29737
rect 27076 29703 27110 29737
rect 27156 29703 27190 29737
rect 27236 29703 27270 29737
rect 26916 29629 26950 29663
rect 26996 29629 27030 29663
rect 27076 29629 27110 29663
rect 27156 29629 27190 29663
rect 27236 29629 27270 29663
rect 26916 29555 26950 29589
rect 26996 29555 27030 29589
rect 27076 29555 27110 29589
rect 27156 29555 27190 29589
rect 27236 29555 27270 29589
rect 26916 29481 26950 29515
rect 26996 29481 27030 29515
rect 27076 29481 27110 29515
rect 27156 29481 27190 29515
rect 27236 29481 27270 29515
rect 26916 29407 26950 29441
rect 26996 29407 27030 29441
rect 27076 29407 27110 29441
rect 27156 29407 27190 29441
rect 27236 29407 27270 29441
rect 26916 29333 26950 29367
rect 26996 29333 27030 29367
rect 27076 29333 27110 29367
rect 27156 29333 27190 29367
rect 27236 29333 27270 29367
rect 26916 29259 26950 29293
rect 26996 29259 27030 29293
rect 27076 29259 27110 29293
rect 27156 29259 27190 29293
rect 27236 29259 27270 29293
rect 26916 29185 26950 29219
rect 26996 29185 27030 29219
rect 27076 29185 27110 29219
rect 27156 29185 27190 29219
rect 27236 29185 27270 29219
rect 26916 29111 26950 29145
rect 26996 29111 27030 29145
rect 27076 29111 27110 29145
rect 27156 29111 27190 29145
rect 27236 29111 27270 29145
rect 26916 29037 26950 29071
rect 26996 29037 27030 29071
rect 27076 29037 27110 29071
rect 27156 29037 27190 29071
rect 27236 29037 27270 29071
rect 26916 28963 26950 28997
rect 26996 28963 27030 28997
rect 27076 28963 27110 28997
rect 27156 28963 27190 28997
rect 27236 28963 27270 28997
rect 26916 28889 26950 28923
rect 26996 28889 27030 28923
rect 27076 28889 27110 28923
rect 27156 28889 27190 28923
rect 27236 28889 27270 28923
rect 26916 28815 26950 28849
rect 26996 28815 27030 28849
rect 27076 28815 27110 28849
rect 27156 28815 27190 28849
rect 27236 28815 27270 28849
rect 26916 28741 26950 28775
rect 26996 28741 27030 28775
rect 27076 28741 27110 28775
rect 27156 28741 27190 28775
rect 27236 28741 27270 28775
rect 26916 28667 26950 28701
rect 26996 28667 27030 28701
rect 27076 28667 27110 28701
rect 27156 28667 27190 28701
rect 27236 28667 27270 28701
rect 26916 28593 26950 28627
rect 26996 28593 27030 28627
rect 27076 28593 27110 28627
rect 27156 28593 27190 28627
rect 27236 28593 27270 28627
rect 26916 28519 26950 28553
rect 26996 28519 27030 28553
rect 27076 28519 27110 28553
rect 27156 28519 27190 28553
rect 27236 28519 27270 28553
rect 439 28441 473 28475
rect 579 28441 613 28475
rect 439 28369 473 28403
rect 579 28369 613 28403
rect 439 28297 473 28331
rect 579 28297 613 28331
rect 439 28225 473 28259
rect 579 28225 613 28259
rect 439 28153 473 28187
rect 579 28153 613 28187
rect 439 28081 473 28115
rect 579 28081 613 28115
rect 439 28009 473 28043
rect 579 28009 613 28043
rect 439 27937 473 27971
rect 579 27937 613 27971
rect 439 27865 473 27899
rect 579 27865 613 27899
rect 439 27793 473 27827
rect 579 27793 613 27827
rect 439 27721 473 27755
rect 579 27721 613 27755
rect 439 27649 473 27683
rect 579 27649 613 27683
rect 439 27577 473 27611
rect 579 27577 613 27611
rect 439 27505 473 27539
rect 579 27505 613 27539
rect 439 27433 473 27467
rect 579 27433 613 27467
rect 439 27361 473 27395
rect 579 27361 613 27395
rect 439 27289 473 27323
rect 579 27289 613 27323
rect 439 27217 473 27251
rect 579 27217 613 27251
rect 439 27145 473 27179
rect 579 27145 613 27179
rect 439 27073 473 27107
rect 579 27073 613 27107
rect 439 27001 473 27035
rect 579 27001 613 27035
rect 439 26929 473 26963
rect 579 26929 613 26963
rect 439 26857 473 26891
rect 579 26857 613 26891
rect 439 26785 473 26819
rect 579 26785 613 26819
rect 439 26713 473 26747
rect 579 26713 613 26747
rect 439 26641 473 26675
rect 579 26641 613 26675
rect 439 26569 473 26603
rect 579 26569 613 26603
rect 439 26496 473 26530
rect 579 26496 613 26530
rect 439 26423 473 26457
rect 579 26423 613 26457
rect 439 26350 473 26384
rect 579 26350 613 26384
rect 439 26277 473 26311
rect 579 26277 613 26311
rect 439 26204 473 26238
rect 579 26204 613 26238
rect 439 26131 473 26165
rect 579 26131 613 26165
rect -2255 26037 -2221 26071
rect -2182 26037 -2148 26071
rect -2109 26037 -2075 26071
rect -2036 26037 -2002 26071
rect -1963 26037 -1929 26071
rect -1890 26037 -1856 26071
rect -1817 26037 -1783 26071
rect -1744 26037 -1710 26071
rect -1671 26037 -1637 26071
rect -1598 26037 -1564 26071
rect -1525 26037 -1491 26071
rect -1453 26037 -1419 26071
rect -2255 25963 -2221 25997
rect -2182 25963 -2148 25997
rect -2109 25963 -2075 25997
rect -2036 25963 -2002 25997
rect -1963 25963 -1929 25997
rect -1890 25963 -1856 25997
rect -1817 25963 -1783 25997
rect -1744 25963 -1710 25997
rect -1671 25963 -1637 25997
rect -1598 25963 -1564 25997
rect -1525 25963 -1491 25997
rect -1453 25963 -1419 25997
rect -2255 25889 -2221 25923
rect -2182 25889 -2148 25923
rect -2109 25889 -2075 25923
rect -2036 25889 -2002 25923
rect -1963 25889 -1929 25923
rect -1890 25889 -1856 25923
rect -1817 25889 -1783 25923
rect -1744 25889 -1710 25923
rect -1671 25889 -1637 25923
rect -1598 25889 -1564 25923
rect -1525 25889 -1491 25923
rect -1453 25889 -1419 25923
rect -2255 25815 -2221 25849
rect -2182 25815 -2148 25849
rect -2109 25815 -2075 25849
rect -2036 25815 -2002 25849
rect -1963 25815 -1929 25849
rect -1890 25815 -1856 25849
rect -1817 25815 -1783 25849
rect -1744 25815 -1710 25849
rect -1671 25815 -1637 25849
rect -1598 25815 -1564 25849
rect -1525 25815 -1491 25849
rect -1453 25815 -1419 25849
rect -2255 25741 -2221 25775
rect -2182 25741 -2148 25775
rect -2109 25741 -2075 25775
rect -2036 25741 -2002 25775
rect -1963 25741 -1929 25775
rect -1890 25741 -1856 25775
rect -1817 25741 -1783 25775
rect -1744 25741 -1710 25775
rect -1671 25741 -1637 25775
rect -1598 25741 -1564 25775
rect -1525 25741 -1491 25775
rect -1453 25741 -1419 25775
rect -2255 25667 -2221 25701
rect -2182 25667 -2148 25701
rect -2109 25667 -2075 25701
rect -2036 25667 -2002 25701
rect -1963 25667 -1929 25701
rect -1890 25667 -1856 25701
rect -1817 25667 -1783 25701
rect -1744 25667 -1710 25701
rect -1671 25667 -1637 25701
rect -1598 25667 -1564 25701
rect -1525 25667 -1491 25701
rect -1453 25667 -1419 25701
rect -2255 25593 -2221 25627
rect -2182 25593 -2148 25627
rect -2109 25593 -2075 25627
rect -2036 25593 -2002 25627
rect -1963 25593 -1929 25627
rect -1890 25593 -1856 25627
rect -1817 25593 -1783 25627
rect -1744 25593 -1710 25627
rect -1671 25593 -1637 25627
rect -1598 25593 -1564 25627
rect -1525 25593 -1491 25627
rect -1453 25593 -1419 25627
rect -1181 25881 -1147 25915
rect -1108 25881 -1074 25915
rect -1035 25881 -1001 25915
rect -962 25881 -928 25915
rect -889 25881 -855 25915
rect -816 25881 -782 25915
rect -743 25881 -709 25915
rect -670 25881 -636 25915
rect -597 25881 -563 25915
rect -524 25881 -490 25915
rect -1181 25809 -1147 25843
rect -1108 25809 -1074 25843
rect -1035 25809 -1001 25843
rect -962 25809 -928 25843
rect -889 25809 -855 25843
rect -816 25809 -782 25843
rect -743 25809 -709 25843
rect -670 25809 -636 25843
rect -597 25809 -563 25843
rect -524 25809 -490 25843
rect -1181 25737 -1147 25771
rect -1108 25737 -1074 25771
rect -1035 25737 -1001 25771
rect -962 25737 -928 25771
rect -889 25737 -855 25771
rect -816 25737 -782 25771
rect -743 25737 -709 25771
rect -670 25737 -636 25771
rect -597 25737 -563 25771
rect -524 25737 -490 25771
rect -1181 25665 -1147 25699
rect -1108 25665 -1074 25699
rect -1035 25665 -1001 25699
rect -962 25665 -928 25699
rect -889 25665 -855 25699
rect -816 25665 -782 25699
rect -743 25665 -709 25699
rect -670 25665 -636 25699
rect -597 25665 -563 25699
rect -524 25665 -490 25699
rect -1181 25593 -1147 25627
rect -1108 25593 -1074 25627
rect -1035 25593 -1001 25627
rect -962 25593 -928 25627
rect -889 25593 -855 25627
rect -816 25593 -782 25627
rect -743 25593 -709 25627
rect -670 25593 -636 25627
rect -597 25593 -563 25627
rect -524 25593 -490 25627
rect -451 25593 2679 25915
rect 31932 23611 31966 23645
rect 32020 23611 32054 23645
rect 31932 23536 31966 23570
rect 32020 23536 32054 23570
rect 31932 23461 31966 23495
rect 32020 23461 32054 23495
rect 17778 23395 17811 23429
rect 17811 23395 17812 23429
rect 17878 23395 17912 23429
rect 17978 23395 18012 23429
rect 17778 23322 17811 23356
rect 17811 23322 17812 23356
rect 17878 23322 17912 23356
rect 17978 23322 18012 23356
rect 17778 23249 17811 23283
rect 17811 23249 17812 23283
rect 17878 23249 17912 23283
rect 17978 23249 18012 23283
rect 31932 23386 31966 23420
rect 32020 23386 32054 23420
rect 31932 23311 31966 23345
rect 32020 23311 32054 23345
rect 31932 23236 31966 23270
rect 32020 23236 32054 23270
rect 17778 23176 17811 23210
rect 17811 23176 17812 23210
rect 17878 23176 17912 23210
rect 17978 23176 18012 23210
rect 17778 23103 17811 23137
rect 17811 23103 17812 23137
rect 17878 23103 17912 23137
rect 17978 23103 18012 23137
rect 17778 23030 17811 23064
rect 17811 23030 17812 23064
rect 17878 23030 17912 23064
rect 17978 23030 18012 23064
rect 17778 22957 17811 22991
rect 17811 22957 17812 22991
rect 17878 22957 17912 22991
rect 17978 22957 18012 22991
rect 17778 22884 17811 22918
rect 17811 22884 17812 22918
rect 17878 22884 17912 22918
rect 17978 22884 18012 22918
rect 17778 22811 17811 22845
rect 17811 22811 17812 22845
rect 17878 22811 17912 22845
rect 17978 22811 18012 22845
rect 17778 22738 17811 22772
rect 17811 22738 17812 22772
rect 17878 22738 17912 22772
rect 17978 22738 18012 22772
rect 17778 22665 17811 22699
rect 17811 22665 17812 22699
rect 17878 22665 17912 22699
rect 17978 22665 18012 22699
rect 17778 22592 17811 22626
rect 17811 22592 17812 22626
rect 17878 22592 17912 22626
rect 17978 22592 18012 22626
rect 17778 22519 17811 22553
rect 17811 22519 17812 22553
rect 17878 22519 17912 22553
rect 17978 22519 18012 22553
rect 17778 22479 17812 22480
rect 17878 22479 17912 22480
rect 17778 22446 17811 22479
rect 17811 22446 17812 22479
rect 17878 22446 17879 22479
rect 17879 22446 17912 22479
rect 17978 22446 18012 22480
rect 17778 22376 17811 22407
rect 17811 22376 17812 22407
rect 17878 22376 17879 22407
rect 17879 22376 17912 22407
rect 17778 22373 17812 22376
rect 17878 22373 17912 22376
rect 17978 22373 18012 22407
rect 17778 22307 17811 22334
rect 17811 22307 17812 22334
rect 17878 22307 17879 22334
rect 17879 22307 17912 22334
rect 17778 22300 17812 22307
rect 17878 22300 17912 22307
rect 17978 22300 18012 22334
rect 17778 22238 17811 22261
rect 17811 22238 17812 22261
rect 17878 22238 17879 22261
rect 17879 22238 17912 22261
rect 17778 22227 17812 22238
rect 17878 22227 17912 22238
rect 17978 22227 18012 22261
rect 17778 22169 17811 22188
rect 17811 22169 17812 22188
rect 17878 22169 17879 22188
rect 17879 22169 17912 22188
rect 17778 22154 17812 22169
rect 17878 22154 17912 22169
rect 17978 22154 18012 22188
rect 17778 22100 17811 22115
rect 17811 22100 17812 22115
rect 17878 22100 17879 22115
rect 17879 22100 17912 22115
rect 17778 22081 17812 22100
rect 17878 22081 17912 22100
rect 17978 22081 18012 22115
rect 17778 22031 17811 22042
rect 17811 22031 17812 22042
rect 17878 22031 17879 22042
rect 17879 22031 17912 22042
rect 17778 22008 17812 22031
rect 17878 22008 17912 22031
rect 17978 22008 18012 22042
rect 17778 21962 17811 21968
rect 17811 21962 17812 21968
rect 17878 21962 17879 21968
rect 17879 21962 17912 21968
rect 17778 21934 17812 21962
rect 17878 21934 17912 21962
rect 17978 21934 18012 21968
rect 17778 21893 17811 21894
rect 17811 21893 17812 21894
rect 17878 21893 17879 21894
rect 17879 21893 17912 21894
rect 17778 21860 17812 21893
rect 17878 21860 17912 21893
rect 17978 21860 18012 21894
rect 17778 21789 17812 21820
rect 17878 21789 17912 21820
rect 17778 21786 17811 21789
rect 17811 21786 17812 21789
rect 17878 21786 17879 21789
rect 17879 21786 17912 21789
rect 17978 21786 18012 21820
rect 17778 21720 17812 21746
rect 17878 21720 17912 21746
rect 17778 21712 17811 21720
rect 17811 21712 17812 21720
rect 17878 21712 17879 21720
rect 17879 21712 17912 21720
rect 17978 21712 18012 21746
rect 17778 21651 17812 21672
rect 17878 21651 17912 21672
rect 17778 21638 17811 21651
rect 17811 21638 17812 21651
rect 17878 21638 17879 21651
rect 17879 21638 17912 21651
rect 17978 21638 18012 21672
rect 17778 21582 17812 21598
rect 17878 21582 17912 21598
rect 17778 21564 17811 21582
rect 17811 21564 17812 21582
rect 17878 21564 17879 21582
rect 17879 21564 17912 21582
rect 17978 21564 18012 21598
rect 17778 21513 17812 21524
rect 17878 21513 17912 21524
rect 17778 21490 17811 21513
rect 17811 21490 17812 21513
rect 17878 21490 17879 21513
rect 17879 21490 17912 21513
rect 17978 21490 18012 21524
rect 17778 21444 17812 21450
rect 17878 21444 17912 21450
rect 17778 21416 17811 21444
rect 17811 21416 17812 21444
rect 17878 21416 17879 21444
rect 17879 21416 17912 21444
rect 17978 21416 18012 21450
rect 17778 21375 17812 21376
rect 17878 21375 17912 21376
rect 17778 21342 17811 21375
rect 17811 21342 17812 21375
rect 17878 21342 17879 21375
rect 17879 21342 17912 21375
rect 17978 21342 18012 21376
rect 17778 21272 17811 21302
rect 17811 21272 17812 21302
rect 17878 21272 17879 21302
rect 17879 21272 17912 21302
rect 17778 21268 17812 21272
rect 17878 21268 17912 21272
rect 17978 21268 18012 21302
rect 17778 21203 17811 21228
rect 17811 21203 17812 21228
rect 17878 21203 17879 21228
rect 17879 21203 17912 21228
rect 17778 21194 17812 21203
rect 17878 21194 17912 21203
rect 17978 21194 18012 21228
rect 17778 21134 17811 21154
rect 17811 21134 17812 21154
rect 17878 21134 17879 21154
rect 17879 21134 17912 21154
rect 17778 21120 17812 21134
rect 17878 21120 17912 21134
rect 17978 21120 18012 21154
rect 17778 21065 17811 21080
rect 17811 21065 17812 21080
rect 17878 21065 17879 21080
rect 17879 21065 17912 21080
rect 17778 21046 17812 21065
rect 17878 21046 17912 21065
rect 17978 21046 18012 21080
rect 17778 20996 17811 21006
rect 17811 20996 17812 21006
rect 17878 20996 17879 21006
rect 17879 20996 17912 21006
rect 17778 20972 17812 20996
rect 17878 20972 17912 20996
rect 17978 20972 18012 21006
rect 31724 23121 31758 23155
rect 31802 23121 31836 23155
rect 31880 23121 31914 23155
rect 31958 23121 31992 23155
rect 32036 23121 32070 23155
rect 31724 23047 31758 23081
rect 31802 23047 31836 23081
rect 31880 23047 31914 23081
rect 31958 23047 31992 23081
rect 32036 23047 32070 23081
rect 31724 22973 31758 23007
rect 31802 22973 31836 23007
rect 31880 22973 31914 23007
rect 31958 22973 31992 23007
rect 32036 22973 32070 23007
rect 31724 22899 31758 22933
rect 31802 22899 31836 22933
rect 31880 22899 31914 22933
rect 31958 22899 31992 22933
rect 32036 22899 32070 22933
rect 31724 22825 31758 22859
rect 31802 22825 31836 22859
rect 31880 22825 31914 22859
rect 31958 22825 31992 22859
rect 32036 22825 32070 22859
rect 31724 22751 31758 22785
rect 31802 22751 31836 22785
rect 31880 22751 31914 22785
rect 31958 22751 31992 22785
rect 32036 22751 32070 22785
rect 31724 22677 31758 22711
rect 31802 22677 31836 22711
rect 31880 22677 31914 22711
rect 31958 22677 31992 22711
rect 32036 22677 32070 22711
rect 31724 22603 31758 22637
rect 31802 22603 31836 22637
rect 31880 22603 31914 22637
rect 31958 22603 31992 22637
rect 32036 22603 32070 22637
rect 31724 22529 31758 22563
rect 31802 22529 31836 22563
rect 31880 22529 31914 22563
rect 31958 22529 31992 22563
rect 32036 22529 32070 22563
rect 31724 22455 31758 22489
rect 31802 22455 31836 22489
rect 31880 22455 31914 22489
rect 31958 22455 31992 22489
rect 32036 22455 32070 22489
rect 31724 22381 31758 22415
rect 31802 22381 31836 22415
rect 31880 22381 31914 22415
rect 31958 22381 31992 22415
rect 32036 22381 32070 22415
rect 31724 22307 31758 22341
rect 31802 22307 31836 22341
rect 31880 22307 31914 22341
rect 31958 22307 31992 22341
rect 32036 22307 32070 22341
rect 31724 22233 31758 22267
rect 31802 22233 31836 22267
rect 31880 22233 31914 22267
rect 31958 22233 31992 22267
rect 32036 22233 32070 22267
rect 31724 22159 31758 22193
rect 31802 22159 31836 22193
rect 31880 22159 31914 22193
rect 31958 22159 31992 22193
rect 32036 22159 32070 22193
rect 31724 22085 31758 22119
rect 31802 22085 31836 22119
rect 31880 22085 31914 22119
rect 31958 22085 31992 22119
rect 32036 22085 32070 22119
rect 31724 22011 31758 22045
rect 31802 22011 31836 22045
rect 31880 22011 31914 22045
rect 31958 22011 31992 22045
rect 32036 22011 32070 22045
rect 31724 21937 31758 21971
rect 31802 21937 31836 21971
rect 31880 21937 31914 21971
rect 31958 21937 31992 21971
rect 32036 21937 32070 21971
rect 31724 21863 31758 21897
rect 31802 21863 31836 21897
rect 31880 21863 31914 21897
rect 31958 21863 31992 21897
rect 32036 21863 32070 21897
rect 31724 21789 31758 21823
rect 31802 21789 31836 21823
rect 31880 21789 31914 21823
rect 31958 21789 31992 21823
rect 32036 21789 32070 21823
rect 31724 21715 31758 21749
rect 31802 21715 31836 21749
rect 31880 21715 31914 21749
rect 31958 21715 31992 21749
rect 32036 21715 32070 21749
rect 31724 21641 31758 21675
rect 31802 21641 31836 21675
rect 31880 21641 31914 21675
rect 31958 21641 31992 21675
rect 32036 21641 32070 21675
rect 31724 21567 31758 21601
rect 31802 21567 31836 21601
rect 31880 21567 31914 21601
rect 31958 21567 31992 21601
rect 32036 21567 32070 21601
rect 31724 21493 31758 21527
rect 31802 21493 31836 21527
rect 31880 21493 31914 21527
rect 31958 21493 31992 21527
rect 32036 21493 32070 21527
rect 31724 21418 31758 21452
rect 31802 21418 31836 21452
rect 31880 21418 31914 21452
rect 31958 21418 31992 21452
rect 32036 21418 32070 21452
rect 31724 21343 31758 21377
rect 31802 21343 31836 21377
rect 31880 21343 31914 21377
rect 31958 21343 31992 21377
rect 32036 21343 32070 21377
rect 31724 21268 31758 21302
rect 31802 21268 31836 21302
rect 31880 21268 31914 21302
rect 31958 21268 31992 21302
rect 32036 21268 32070 21302
rect 31724 21193 31758 21227
rect 31802 21193 31836 21227
rect 31880 21193 31914 21227
rect 31958 21193 31992 21227
rect 32036 21193 32070 21227
rect 31724 21118 31758 21152
rect 31802 21118 31836 21152
rect 31880 21118 31914 21152
rect 31958 21118 31992 21152
rect 32036 21118 32070 21152
rect 31724 21043 31758 21077
rect 31802 21043 31836 21077
rect 31880 21043 31914 21077
rect 31958 21043 31992 21077
rect 32036 21043 32070 21077
rect 31724 20968 31758 21002
rect 31802 20968 31836 21002
rect 31880 20968 31914 21002
rect 31958 20968 31992 21002
rect 32036 20968 32070 21002
rect 17778 20927 17811 20932
rect 17811 20927 17812 20932
rect 17878 20927 17879 20932
rect 17879 20927 17912 20932
rect 17778 20898 17812 20927
rect 17878 20898 17912 20927
rect 17978 20898 18012 20932
rect 17778 20824 17812 20858
rect 17878 20824 17912 20858
rect 17978 20824 18012 20858
rect 17778 20754 17812 20784
rect 17878 20754 17912 20784
rect 17778 20750 17811 20754
rect 17811 20750 17812 20754
rect 17878 20750 17879 20754
rect 17879 20750 17912 20754
rect 17978 20750 18012 20784
rect 17778 20685 17812 20710
rect 17878 20685 17912 20710
rect 17778 20676 17811 20685
rect 17811 20676 17812 20685
rect 17878 20676 17879 20685
rect 17879 20676 17912 20685
rect 17978 20676 18012 20710
rect 17778 20616 17812 20636
rect 17878 20616 17912 20636
rect 17778 20602 17811 20616
rect 17811 20602 17812 20616
rect 17878 20602 17879 20616
rect 17879 20602 17912 20616
rect 17978 20602 18012 20636
rect 17778 20547 17812 20562
rect 17878 20547 17912 20562
rect 17778 20528 17811 20547
rect 17811 20528 17812 20547
rect 17878 20528 17879 20547
rect 17879 20528 17912 20547
rect 17978 20528 18012 20562
rect 17778 20478 17812 20488
rect 17878 20478 17912 20488
rect 17778 20454 17811 20478
rect 17811 20454 17812 20478
rect 17878 20454 17879 20478
rect 17879 20454 17912 20478
rect 17978 20454 18012 20488
rect 17778 20409 17812 20414
rect 17878 20409 17912 20414
rect 17778 20380 17811 20409
rect 17811 20380 17812 20409
rect 17878 20380 17879 20409
rect 17879 20380 17912 20409
rect 17978 20380 18012 20414
rect 17778 20306 17811 20340
rect 17811 20306 17812 20340
rect 17878 20306 17879 20340
rect 17879 20306 17912 20340
rect 17978 20306 18012 20340
rect -2289 13313 -2255 13347
rect -2215 13313 -2181 13347
rect -2141 13313 -2107 13347
rect -2067 13313 -2033 13347
rect -1993 13313 -1959 13347
rect -1919 13313 -1885 13347
rect -1845 13313 -1811 13347
rect -1771 13313 -1737 13347
rect -1698 13313 -1664 13347
rect -1625 13313 -1591 13347
rect -1552 13313 -1518 13347
rect -2289 13229 -2255 13263
rect -2215 13229 -2181 13263
rect -2141 13229 -2107 13263
rect -2067 13229 -2033 13263
rect -1993 13229 -1959 13263
rect -1919 13229 -1885 13263
rect -1845 13229 -1811 13263
rect -1771 13229 -1737 13263
rect -1698 13229 -1664 13263
rect -1625 13229 -1591 13263
rect -1552 13229 -1518 13263
rect 28826 7430 28837 7439
rect 28837 7430 28860 7439
rect 28899 7430 28906 7439
rect 28906 7430 28933 7439
rect 28972 7430 28975 7439
rect 28975 7430 29006 7439
rect 28826 7405 28860 7430
rect 28899 7405 28933 7430
rect 28972 7405 29006 7430
rect 29045 7405 29079 7439
rect 29117 7430 29148 7439
rect 29148 7430 29151 7439
rect 29189 7430 29217 7439
rect 29217 7430 29223 7439
rect 29261 7430 29286 7439
rect 29286 7430 29295 7439
rect 29333 7430 29355 7439
rect 29355 7430 29367 7439
rect 29405 7430 29424 7439
rect 29424 7430 29439 7439
rect 29477 7430 29493 7439
rect 29493 7430 29511 7439
rect 29549 7430 29562 7439
rect 29562 7430 29583 7439
rect 29621 7430 29631 7439
rect 29631 7430 29655 7439
rect 29693 7430 29700 7439
rect 29700 7430 29727 7439
rect 29765 7430 29769 7439
rect 29769 7430 29799 7439
rect 29837 7430 29838 7439
rect 29838 7430 29871 7439
rect 29909 7430 29941 7439
rect 29941 7430 29943 7439
rect 29981 7430 30010 7439
rect 30010 7430 30015 7439
rect 30053 7430 30079 7439
rect 30079 7430 30087 7439
rect 30125 7430 30148 7439
rect 30148 7430 30159 7439
rect 30197 7430 30217 7439
rect 30217 7430 30231 7439
rect 30269 7430 30286 7439
rect 30286 7430 30303 7439
rect 30341 7430 30355 7439
rect 30355 7430 30375 7439
rect 30413 7430 30424 7439
rect 30424 7430 30447 7439
rect 30485 7430 30493 7439
rect 30493 7430 30519 7439
rect 30557 7430 30562 7439
rect 30562 7430 30591 7439
rect 29117 7405 29151 7430
rect 29189 7405 29223 7430
rect 29261 7405 29295 7430
rect 29333 7405 29367 7430
rect 29405 7405 29439 7430
rect 29477 7405 29511 7430
rect 29549 7405 29583 7430
rect 29621 7405 29655 7430
rect 29693 7405 29727 7430
rect 29765 7405 29799 7430
rect 29837 7405 29871 7430
rect 29909 7405 29943 7430
rect 29981 7405 30015 7430
rect 30053 7405 30087 7430
rect 30125 7405 30159 7430
rect 30197 7405 30231 7430
rect 30269 7405 30303 7430
rect 30341 7405 30375 7430
rect 30413 7405 30447 7430
rect 30485 7405 30519 7430
rect 30557 7405 30591 7430
rect 30629 7405 30663 7439
rect 30701 7405 30735 7439
rect 30773 7405 30807 7439
rect 30845 7405 30879 7439
rect 30917 7405 30951 7439
rect 28754 7362 28768 7364
rect 28768 7362 28788 7364
rect 28754 7330 28788 7362
rect 28866 7294 28872 7327
rect 28872 7294 28900 7327
rect 28940 7294 28941 7327
rect 28941 7294 28974 7327
rect 29014 7294 29044 7327
rect 29044 7294 29048 7327
rect 29088 7294 29113 7327
rect 29113 7294 29122 7327
rect 29162 7294 29182 7327
rect 29182 7294 29196 7327
rect 29236 7294 29251 7327
rect 29251 7294 29270 7327
rect 29310 7294 29320 7327
rect 29320 7294 29344 7327
rect 29384 7294 29389 7327
rect 29389 7294 29418 7327
rect 29457 7294 29458 7327
rect 29458 7294 29491 7327
rect 29530 7294 29562 7327
rect 29562 7294 29564 7327
rect 29603 7294 29631 7327
rect 29631 7294 29637 7327
rect 29676 7294 29700 7327
rect 29700 7294 29710 7327
rect 29749 7294 29769 7327
rect 29769 7294 29783 7327
rect 29822 7294 29838 7327
rect 29838 7294 29856 7327
rect 29895 7294 29907 7327
rect 29907 7294 29929 7327
rect 29968 7294 29976 7327
rect 29976 7294 30002 7327
rect 30041 7294 30045 7327
rect 30045 7294 30075 7327
rect 30114 7294 30148 7327
rect 30187 7294 30217 7327
rect 30217 7294 30221 7327
rect 30260 7294 30286 7327
rect 30286 7294 30294 7327
rect 30333 7294 30355 7327
rect 30355 7294 30367 7327
rect 30406 7294 30424 7327
rect 30424 7294 30440 7327
rect 30479 7294 30493 7327
rect 30493 7294 30513 7327
rect 30552 7294 30562 7327
rect 30562 7294 30586 7327
rect 30625 7294 30659 7327
rect 30698 7294 30732 7327
rect 30771 7294 30805 7327
rect 30844 7294 30878 7327
rect 30917 7294 30951 7327
rect 28866 7293 28900 7294
rect 28940 7293 28974 7294
rect 29014 7293 29048 7294
rect 29088 7293 29122 7294
rect 29162 7293 29196 7294
rect 29236 7293 29270 7294
rect 29310 7293 29344 7294
rect 29384 7293 29418 7294
rect 29457 7293 29491 7294
rect 29530 7293 29564 7294
rect 29603 7293 29637 7294
rect 29676 7293 29710 7294
rect 29749 7293 29783 7294
rect 29822 7293 29856 7294
rect 29895 7293 29929 7294
rect 29968 7293 30002 7294
rect 30041 7293 30075 7294
rect 30114 7293 30148 7294
rect 30187 7293 30221 7294
rect 30260 7293 30294 7294
rect 30333 7293 30367 7294
rect 30406 7293 30440 7294
rect 30479 7293 30513 7294
rect 30552 7293 30586 7294
rect 30625 7293 30659 7294
rect 30698 7293 30732 7294
rect 30771 7293 30805 7294
rect 30844 7293 30878 7294
rect 30917 7293 30951 7294
rect 28754 7255 28788 7289
rect 28754 7180 28788 7214
rect 28866 7212 28900 7246
rect 28754 7105 28788 7139
rect 28866 7131 28900 7165
rect 28754 7030 28788 7064
rect 28866 7049 28900 7083
rect 28754 6955 28788 6989
rect 28866 6967 28900 7001
rect 28754 6880 28788 6913
rect 28866 6885 28900 6919
rect 28754 6879 28777 6880
rect 28777 6879 28788 6880
rect 28754 6811 28788 6837
rect 28754 6803 28777 6811
rect 28777 6803 28788 6811
rect 28866 6803 28900 6837
rect 30216 5823 30248 5835
rect 30248 5823 30250 5835
rect 30291 5823 30317 5835
rect 30317 5823 30325 5835
rect 30366 5823 30386 5835
rect 30386 5823 30400 5835
rect 30441 5823 30455 5835
rect 30455 5823 30475 5835
rect 30516 5823 30524 5835
rect 30524 5823 30550 5835
rect 30591 5823 30593 5835
rect 30593 5823 30625 5835
rect 30666 5823 30697 5835
rect 30697 5823 30700 5835
rect 30741 5823 30766 5835
rect 30766 5823 30775 5835
rect 30816 5823 30835 5835
rect 30835 5823 30850 5835
rect 30891 5823 30904 5835
rect 30904 5823 30925 5835
rect 30966 5823 30973 5835
rect 30973 5823 31000 5835
rect 31041 5823 31042 5835
rect 31042 5823 31075 5835
rect 31116 5823 31145 5835
rect 31145 5823 31150 5835
rect 31191 5823 31214 5835
rect 31214 5823 31225 5835
rect 31266 5823 31283 5835
rect 31283 5823 31300 5835
rect 31341 5823 31352 5835
rect 31352 5823 31375 5835
rect 31416 5823 31421 5835
rect 31421 5823 31450 5835
rect 31491 5823 31523 5835
rect 31523 5823 31525 5835
rect 31566 5823 31591 5835
rect 31591 5823 31600 5835
rect 31640 5823 31659 5835
rect 31659 5823 31674 5835
rect 31714 5823 31727 5835
rect 31727 5823 31748 5835
rect 31788 5823 31795 5835
rect 31795 5823 31822 5835
rect 31862 5823 31863 5835
rect 31863 5823 31896 5835
rect 31936 5823 31965 5835
rect 31965 5823 31970 5835
rect 32010 5823 32033 5835
rect 32033 5823 32044 5835
rect 30216 5801 30250 5823
rect 30291 5801 30325 5823
rect 30366 5801 30400 5823
rect 30441 5801 30475 5823
rect 30516 5801 30550 5823
rect 30591 5801 30625 5823
rect 30666 5801 30700 5823
rect 30741 5801 30775 5823
rect 30816 5801 30850 5823
rect 30891 5801 30925 5823
rect 30966 5801 31000 5823
rect 31041 5801 31075 5823
rect 31116 5801 31150 5823
rect 31191 5801 31225 5823
rect 31266 5801 31300 5823
rect 31341 5801 31375 5823
rect 31416 5801 31450 5823
rect 31491 5801 31525 5823
rect 31566 5801 31600 5823
rect 31640 5801 31674 5823
rect 31714 5801 31748 5823
rect 31788 5801 31822 5823
rect 31862 5801 31896 5823
rect 31936 5801 31970 5823
rect 32010 5801 32044 5823
rect 16808 5511 16842 5545
rect 16881 5511 16915 5545
rect 16954 5511 16988 5545
rect 17027 5511 17061 5545
rect 17100 5511 17134 5545
rect 17173 5511 17207 5545
rect 17246 5511 17280 5545
rect 17319 5511 17353 5545
rect 17392 5511 17426 5545
rect 17465 5511 17499 5545
rect 17538 5511 17572 5545
rect 17611 5511 17645 5545
rect 17684 5511 17718 5545
rect 17757 5511 17791 5545
rect 17830 5511 17864 5545
rect 17903 5511 17937 5545
rect 17976 5511 18010 5545
rect 18049 5511 18083 5545
rect 18122 5511 18156 5545
rect 18195 5511 18229 5545
rect 18268 5511 18302 5545
rect 18341 5511 18375 5545
rect 18414 5511 18448 5545
rect 18487 5511 18521 5545
rect 18560 5511 18594 5545
rect 18633 5511 18667 5545
rect 18705 5511 18739 5545
rect 18777 5511 18811 5545
rect 18849 5511 18883 5545
rect 18921 5511 18955 5545
rect 16808 5433 16842 5467
rect 16881 5433 16915 5467
rect 16954 5433 16988 5467
rect 17027 5433 17061 5467
rect 17100 5433 17134 5467
rect 17173 5433 17207 5467
rect 17246 5433 17280 5467
rect 17319 5433 17353 5467
rect 17392 5433 17426 5467
rect 17465 5433 17499 5467
rect 17538 5433 17572 5467
rect 17611 5433 17645 5467
rect 17684 5433 17718 5467
rect 17757 5433 17791 5467
rect 17830 5433 17864 5467
rect 17903 5433 17937 5467
rect 17976 5433 18010 5467
rect 18049 5433 18083 5467
rect 18122 5433 18156 5467
rect 18195 5433 18229 5467
rect 18268 5433 18302 5467
rect 18341 5433 18375 5467
rect 18414 5433 18448 5467
rect 18487 5433 18521 5467
rect 18560 5433 18594 5467
rect 18633 5433 18667 5467
rect 18705 5433 18739 5467
rect 18777 5433 18811 5467
rect 18849 5433 18883 5467
rect 18921 5433 18955 5467
rect 16808 5355 16842 5389
rect 16881 5355 16915 5389
rect 16954 5355 16988 5389
rect 17027 5355 17061 5389
rect 17100 5355 17134 5389
rect 17173 5355 17207 5389
rect 17246 5355 17280 5389
rect 17319 5355 17353 5389
rect 17392 5355 17426 5389
rect 17465 5355 17499 5389
rect 17538 5355 17572 5389
rect 17611 5355 17645 5389
rect 17684 5355 17718 5389
rect 17757 5355 17791 5389
rect 17830 5355 17864 5389
rect 17903 5355 17937 5389
rect 17976 5355 18010 5389
rect 18049 5355 18083 5389
rect 18122 5355 18156 5389
rect 18195 5355 18229 5389
rect 18268 5355 18302 5389
rect 18341 5355 18375 5389
rect 18414 5355 18448 5389
rect 18487 5355 18521 5389
rect 18560 5355 18594 5389
rect 18633 5355 18667 5389
rect 18705 5355 18739 5389
rect 18777 5355 18811 5389
rect 18849 5355 18883 5389
rect 18921 5355 18955 5389
rect 16808 5277 16842 5311
rect 16881 5277 16915 5311
rect 16954 5277 16988 5311
rect 17027 5277 17061 5311
rect 17100 5277 17134 5311
rect 17173 5277 17207 5311
rect 17246 5277 17280 5311
rect 17319 5277 17353 5311
rect 17392 5277 17426 5311
rect 17465 5277 17499 5311
rect 17538 5277 17572 5311
rect 17611 5277 17645 5311
rect 17684 5277 17718 5311
rect 17757 5277 17791 5311
rect 17830 5277 17864 5311
rect 17903 5277 17937 5311
rect 17976 5277 18010 5311
rect 18049 5277 18083 5311
rect 18122 5277 18156 5311
rect 18195 5277 18229 5311
rect 18268 5277 18302 5311
rect 18341 5277 18375 5311
rect 18414 5277 18448 5311
rect 18487 5277 18521 5311
rect 18560 5277 18594 5311
rect 18633 5277 18667 5311
rect 18705 5277 18739 5311
rect 18777 5277 18811 5311
rect 18849 5277 18883 5311
rect 18921 5277 18955 5311
rect 27910 5101 27944 5135
rect 27988 5101 28022 5135
rect 28066 5101 28100 5135
rect 28144 5101 28178 5135
rect 28222 5101 28256 5135
rect 28300 5101 28334 5135
rect 28378 5101 28412 5135
rect 28456 5101 28490 5135
rect 28534 5101 28568 5135
rect 28612 5101 28646 5135
rect 27910 5024 27944 5058
rect 27988 5024 28022 5058
rect 28066 5024 28100 5058
rect 28144 5024 28178 5058
rect 28222 5024 28256 5058
rect 28300 5024 28334 5058
rect 28378 5024 28412 5058
rect 28456 5024 28490 5058
rect 28534 5024 28568 5058
rect 28612 5024 28646 5058
rect 27910 4946 27944 4980
rect 27988 4946 28022 4980
rect 28066 4946 28100 4980
rect 28144 4946 28178 4980
rect 28222 4946 28256 4980
rect 28300 4946 28334 4980
rect 28378 4946 28412 4980
rect 28456 4946 28490 4980
rect 28534 4946 28568 4980
rect 28612 4946 28646 4980
rect 27910 4868 27944 4902
rect 27988 4868 28022 4902
rect 28066 4868 28100 4902
rect 28144 4868 28178 4902
rect 28222 4868 28256 4902
rect 28300 4868 28334 4902
rect 28378 4868 28412 4902
rect 28456 4868 28490 4902
rect 28534 4868 28568 4902
rect 28612 4868 28646 4902
rect 27910 4790 27944 4824
rect 27988 4790 28022 4824
rect 28066 4790 28100 4824
rect 28144 4790 28178 4824
rect 28222 4790 28256 4824
rect 28300 4790 28334 4824
rect 28378 4790 28412 4824
rect 28456 4790 28490 4824
rect 28534 4790 28568 4824
rect 28612 4790 28646 4824
rect 27910 4712 27944 4746
rect 27988 4712 28022 4746
rect 28066 4712 28100 4746
rect 28144 4712 28178 4746
rect 28222 4712 28256 4746
rect 28300 4712 28334 4746
rect 28378 4712 28412 4746
rect 28456 4712 28490 4746
rect 28534 4712 28568 4746
rect 28612 4712 28646 4746
rect 27910 4634 27944 4668
rect 27988 4634 28022 4668
rect 28066 4634 28100 4668
rect 28144 4634 28178 4668
rect 28222 4634 28256 4668
rect 28300 4634 28334 4668
rect 28378 4634 28412 4668
rect 28456 4634 28490 4668
rect 28534 4634 28568 4668
rect 28612 4634 28646 4668
rect 26713 4581 26740 4615
rect 26740 4581 26747 4615
rect 26788 4581 26809 4615
rect 26809 4581 26822 4615
rect 26863 4581 26878 4615
rect 26878 4581 26897 4615
rect 26938 4581 26947 4615
rect 26947 4581 26972 4615
rect 27013 4581 27016 4615
rect 27016 4581 27047 4615
rect 27088 4581 27119 4615
rect 27119 4581 27122 4615
rect 27163 4581 27188 4615
rect 27188 4581 27197 4615
rect 27238 4581 27257 4615
rect 27257 4581 27272 4615
rect 27312 4581 27326 4615
rect 27326 4581 27346 4615
rect 27386 4581 27395 4615
rect 27395 4581 27420 4615
rect 27460 4581 27464 4615
rect 27464 4581 27494 4615
rect 27534 4581 27568 4615
rect 27608 4581 27642 4615
rect 27682 4581 27716 4615
rect 27756 4581 27790 4615
rect 27910 4556 27944 4590
rect 27988 4556 28022 4590
rect 28066 4556 28100 4590
rect 28144 4556 28178 4590
rect 28222 4556 28256 4590
rect 28300 4556 28334 4590
rect 28378 4556 28412 4590
rect 28456 4556 28490 4590
rect 28534 4556 28568 4590
rect 28612 4556 28646 4590
rect 26713 4513 26740 4535
rect 26740 4513 26747 4535
rect 26788 4513 26809 4535
rect 26809 4513 26822 4535
rect 26863 4513 26878 4535
rect 26878 4513 26897 4535
rect 26938 4513 26947 4535
rect 26947 4513 26972 4535
rect 27013 4513 27016 4535
rect 27016 4513 27047 4535
rect 27088 4513 27119 4535
rect 27119 4513 27122 4535
rect 27163 4513 27188 4535
rect 27188 4513 27197 4535
rect 27238 4513 27257 4535
rect 27257 4513 27272 4535
rect 27312 4513 27326 4535
rect 27326 4513 27346 4535
rect 27386 4513 27395 4535
rect 27395 4513 27420 4535
rect 27460 4513 27464 4535
rect 27464 4513 27494 4535
rect 26713 4501 26747 4513
rect 26788 4501 26822 4513
rect 26863 4501 26897 4513
rect 26938 4501 26972 4513
rect 27013 4501 27047 4513
rect 27088 4501 27122 4513
rect 27163 4501 27197 4513
rect 27238 4501 27272 4513
rect 27312 4501 27346 4513
rect 27386 4501 27420 4513
rect 27460 4501 27494 4513
rect 27534 4501 27568 4535
rect 27608 4501 27642 4535
rect 27682 4501 27716 4535
rect 27756 4501 27790 4535
rect 26713 4445 26740 4455
rect 26740 4445 26747 4455
rect 26788 4445 26809 4455
rect 26809 4445 26822 4455
rect 26863 4445 26878 4455
rect 26878 4445 26897 4455
rect 26938 4445 26947 4455
rect 26947 4445 26972 4455
rect 27013 4445 27016 4455
rect 27016 4445 27047 4455
rect 27088 4445 27119 4455
rect 27119 4445 27122 4455
rect 27163 4445 27188 4455
rect 27188 4445 27197 4455
rect 27238 4445 27257 4455
rect 27257 4445 27272 4455
rect 27312 4445 27326 4455
rect 27326 4445 27346 4455
rect 27386 4445 27395 4455
rect 27395 4445 27420 4455
rect 27460 4445 27464 4455
rect 27464 4445 27494 4455
rect 27910 4478 27944 4512
rect 27988 4478 28022 4512
rect 28066 4478 28100 4512
rect 28144 4478 28178 4512
rect 28222 4478 28256 4512
rect 28300 4478 28334 4512
rect 28378 4478 28412 4512
rect 28456 4478 28490 4512
rect 28534 4478 28568 4512
rect 28612 4478 28646 4512
rect 26713 4421 26747 4445
rect 26788 4421 26822 4445
rect 26863 4421 26897 4445
rect 26938 4421 26972 4445
rect 27013 4421 27047 4445
rect 27088 4421 27122 4445
rect 27163 4421 27197 4445
rect 27238 4421 27272 4445
rect 27312 4421 27346 4445
rect 27386 4421 27420 4445
rect 27460 4421 27494 4445
rect 27534 4421 27568 4455
rect 27608 4421 27642 4455
rect 27682 4421 27716 4455
rect 27756 4421 27790 4455
rect 27910 4400 27944 4434
rect 27988 4400 28022 4434
rect 28066 4400 28100 4434
rect 28144 4400 28178 4434
rect 28222 4400 28256 4434
rect 28300 4400 28334 4434
rect 28378 4400 28412 4434
rect 28456 4400 28490 4434
rect 28534 4400 28568 4434
rect 28612 4400 28646 4434
rect 26713 4343 26747 4375
rect 26788 4343 26822 4375
rect 26863 4343 26897 4375
rect 26938 4343 26972 4375
rect 27013 4343 27047 4375
rect 27088 4343 27122 4375
rect 27163 4343 27197 4375
rect 27238 4343 27272 4375
rect 27312 4343 27346 4375
rect 27386 4343 27420 4375
rect 27460 4343 27494 4375
rect 26713 4341 26740 4343
rect 26740 4341 26747 4343
rect 26788 4341 26809 4343
rect 26809 4341 26822 4343
rect 26863 4341 26878 4343
rect 26878 4341 26897 4343
rect 26938 4341 26947 4343
rect 26947 4341 26972 4343
rect 27013 4341 27016 4343
rect 27016 4341 27047 4343
rect 27088 4341 27119 4343
rect 27119 4341 27122 4343
rect 27163 4341 27188 4343
rect 27188 4341 27197 4343
rect 27238 4341 27257 4343
rect 27257 4341 27272 4343
rect 27312 4341 27326 4343
rect 27326 4341 27346 4343
rect 27386 4341 27395 4343
rect 27395 4341 27420 4343
rect 27460 4341 27464 4343
rect 27464 4341 27494 4343
rect 27534 4341 27568 4375
rect 27608 4341 27642 4375
rect 27682 4341 27716 4375
rect 27756 4341 27790 4375
rect 27910 4322 27944 4356
rect 27988 4322 28022 4356
rect 28066 4322 28100 4356
rect 28144 4322 28178 4356
rect 28222 4322 28256 4356
rect 28300 4322 28334 4356
rect 28378 4322 28412 4356
rect 28456 4322 28490 4356
rect 28534 4322 28568 4356
rect 28612 4322 28646 4356
rect 26713 4275 26747 4295
rect 26788 4275 26822 4295
rect 26863 4275 26897 4295
rect 26938 4275 26972 4295
rect 27013 4275 27047 4295
rect 27088 4275 27122 4295
rect 27163 4275 27197 4295
rect 27238 4275 27272 4295
rect 27312 4275 27346 4295
rect 27386 4275 27420 4295
rect 27460 4275 27494 4295
rect 26713 4261 26740 4275
rect 26740 4261 26747 4275
rect 26788 4261 26809 4275
rect 26809 4261 26822 4275
rect 26863 4261 26878 4275
rect 26878 4261 26897 4275
rect 26938 4261 26947 4275
rect 26947 4261 26972 4275
rect 27013 4261 27016 4275
rect 27016 4261 27047 4275
rect 27088 4261 27119 4275
rect 27119 4261 27122 4275
rect 27163 4261 27188 4275
rect 27188 4261 27197 4275
rect 27238 4261 27257 4275
rect 27257 4261 27272 4275
rect 27312 4261 27326 4275
rect 27326 4261 27346 4275
rect 27386 4261 27395 4275
rect 27395 4261 27420 4275
rect 27460 4261 27464 4275
rect 27464 4261 27494 4275
rect 27534 4261 27568 4295
rect 27608 4261 27642 4295
rect 27682 4261 27716 4295
rect 27756 4261 27790 4295
rect 27910 4244 27944 4278
rect 27988 4244 28022 4278
rect 28066 4244 28100 4278
rect 28144 4244 28178 4278
rect 28222 4244 28256 4278
rect 28300 4244 28334 4278
rect 28378 4244 28412 4278
rect 28456 4244 28490 4278
rect 28534 4244 28568 4278
rect 28612 4244 28646 4278
rect 26713 4181 26747 4215
rect 26788 4181 26822 4215
rect 26863 4181 26897 4215
rect 26938 4181 26972 4215
rect 27013 4181 27047 4215
rect 27088 4181 27122 4215
rect 27163 4181 27197 4215
rect 27238 4181 27272 4215
rect 27312 4181 27346 4215
rect 27386 4181 27420 4215
rect 27460 4181 27494 4215
rect 27534 4181 27568 4215
rect 27608 4181 27642 4215
rect 27682 4181 27716 4215
rect 27756 4181 27790 4215
rect 27910 4166 27944 4200
rect 27988 4166 28022 4200
rect 28066 4166 28100 4200
rect 28144 4166 28178 4200
rect 28222 4166 28256 4200
rect 28300 4166 28334 4200
rect 28378 4166 28412 4200
rect 28456 4166 28490 4200
rect 28534 4166 28568 4200
rect 28612 4166 28646 4200
rect 9109 3273 9143 3307
rect 9109 3201 9143 3235
rect 9281 3273 9315 3307
rect 9281 3201 9315 3235
rect 10769 3273 10803 3307
rect 10769 3201 10803 3235
rect 10941 3273 10975 3307
rect 10941 3201 10975 3235
rect 22405 2428 22439 2462
rect 22507 2428 22541 2462
rect 22609 2428 22643 2462
rect 22405 2369 22415 2387
rect 22415 2369 22439 2387
rect 22507 2369 22517 2387
rect 22517 2369 22541 2387
rect 22609 2369 22619 2387
rect 22619 2369 22643 2387
rect 22405 2353 22439 2369
rect 22507 2353 22541 2369
rect 22609 2353 22643 2369
rect 22405 2294 22415 2312
rect 22415 2294 22439 2312
rect 22507 2294 22517 2312
rect 22517 2294 22541 2312
rect 22609 2294 22619 2312
rect 22619 2294 22643 2312
rect 22405 2278 22439 2294
rect 22507 2278 22541 2294
rect 22609 2278 22643 2294
rect 22405 2218 22415 2237
rect 22415 2218 22439 2237
rect 22507 2218 22517 2237
rect 22517 2218 22541 2237
rect 22609 2218 22619 2237
rect 22619 2218 22643 2237
rect 22405 2203 22439 2218
rect 22507 2203 22541 2218
rect 22609 2203 22643 2218
rect 22405 2142 22415 2162
rect 22415 2142 22439 2162
rect 22507 2142 22517 2162
rect 22517 2142 22541 2162
rect 22609 2142 22619 2162
rect 22619 2142 22643 2162
rect 22405 2128 22439 2142
rect 22507 2128 22541 2142
rect 22609 2128 22643 2142
rect 22405 2066 22415 2087
rect 22415 2066 22439 2087
rect 22507 2066 22517 2087
rect 22517 2066 22541 2087
rect 22609 2066 22619 2087
rect 22619 2066 22643 2087
rect 22405 2053 22439 2066
rect 22507 2053 22541 2066
rect 22609 2053 22643 2066
rect 22405 1990 22415 2012
rect 22415 1990 22439 2012
rect 22507 1990 22517 2012
rect 22517 1990 22541 2012
rect 22609 1990 22619 2012
rect 22619 1990 22643 2012
rect 22405 1978 22439 1990
rect 22507 1978 22541 1990
rect 22609 1978 22643 1990
rect 22405 1914 22415 1936
rect 22415 1914 22439 1936
rect 22507 1914 22517 1936
rect 22517 1914 22541 1936
rect 22609 1914 22619 1936
rect 22619 1914 22643 1936
rect 22405 1902 22439 1914
rect 22507 1902 22541 1914
rect 22609 1902 22643 1914
rect 22405 1838 22415 1860
rect 22415 1838 22439 1860
rect 22507 1838 22517 1860
rect 22517 1838 22541 1860
rect 22609 1838 22619 1860
rect 22619 1838 22643 1860
rect 22405 1826 22439 1838
rect 22507 1826 22541 1838
rect 22609 1826 22643 1838
rect 22405 1762 22415 1784
rect 22415 1762 22439 1784
rect 22507 1762 22517 1784
rect 22517 1762 22541 1784
rect 22609 1762 22619 1784
rect 22619 1762 22643 1784
rect 22405 1750 22439 1762
rect 22507 1750 22541 1762
rect 22609 1750 22643 1762
<< metal1 >>
tri 433 41919 621 42107 se
rect 621 41919 677 42107
rect 433 41880 677 41919
rect 433 33062 448 41880
rect 626 33062 677 41880
rect 433 33023 677 33062
rect 433 32989 448 33023
rect 482 32989 520 33023
rect 554 32989 592 33023
rect 626 32989 677 33023
rect 433 32950 677 32989
rect 433 32916 448 32950
rect 482 32916 520 32950
rect 554 32916 592 32950
rect 626 32916 677 32950
rect 433 32877 677 32916
rect 433 32843 448 32877
rect 482 32843 520 32877
rect 554 32843 592 32877
rect 626 32843 677 32877
rect 433 32804 677 32843
rect 433 32770 448 32804
rect 482 32770 520 32804
rect 554 32770 592 32804
rect 626 32770 677 32804
rect 433 32731 677 32770
rect 433 32697 448 32731
rect 482 32697 520 32731
rect 554 32697 592 32731
rect 626 32697 677 32731
rect 433 32658 677 32697
rect 433 32624 448 32658
rect 482 32624 520 32658
rect 554 32624 592 32658
rect 626 32624 677 32658
rect 433 32585 677 32624
rect 433 32551 448 32585
rect 482 32551 520 32585
rect 554 32551 592 32585
rect 626 32551 677 32585
rect 433 32512 677 32551
rect 433 32478 448 32512
rect 482 32478 520 32512
rect 554 32478 592 32512
rect 626 32478 677 32512
rect 433 32439 677 32478
rect 433 32405 448 32439
rect 482 32405 520 32439
rect 554 32405 592 32439
rect 626 32405 677 32439
rect 433 32366 677 32405
rect 433 32332 448 32366
rect 482 32332 520 32366
rect 554 32332 592 32366
rect 626 32332 677 32366
rect 433 32293 677 32332
rect 433 32259 448 32293
rect 482 32259 520 32293
rect 554 32259 592 32293
rect 626 32259 677 32293
rect 433 32220 677 32259
rect 433 32186 448 32220
rect 482 32186 520 32220
rect 554 32186 592 32220
rect 626 32186 677 32220
rect 433 32147 677 32186
rect 433 32113 448 32147
rect 482 32113 520 32147
rect 554 32113 592 32147
rect 626 32113 677 32147
rect 433 32074 677 32113
rect 433 32040 448 32074
rect 482 32040 520 32074
rect 554 32040 592 32074
rect 626 32040 677 32074
rect 433 32001 677 32040
rect 433 31967 448 32001
rect 482 31967 520 32001
rect 554 31967 592 32001
rect 626 31967 677 32001
rect 433 31928 677 31967
rect 433 31894 448 31928
rect 482 31894 520 31928
rect 554 31894 592 31928
rect 626 31894 677 31928
rect 433 31855 677 31894
rect 433 31821 448 31855
rect 482 31821 520 31855
rect 554 31821 592 31855
rect 626 31821 677 31855
rect 433 31782 677 31821
rect 433 31748 448 31782
rect 482 31748 520 31782
rect 554 31748 592 31782
rect 626 31748 677 31782
rect 433 31709 677 31748
rect 433 31675 448 31709
rect 482 31675 520 31709
rect 554 31675 592 31709
rect 626 31675 677 31709
rect 433 31636 677 31675
rect 433 31602 448 31636
rect 482 31602 520 31636
rect 554 31602 592 31636
rect 626 31602 677 31636
rect 433 31563 677 31602
rect 433 31529 448 31563
rect 482 31529 520 31563
rect 554 31529 592 31563
rect 626 31529 677 31563
rect 433 31490 677 31529
rect 433 31456 448 31490
rect 482 31456 520 31490
rect 554 31456 592 31490
rect 626 31456 677 31490
rect 433 31417 677 31456
rect 433 31383 448 31417
rect 482 31383 520 31417
rect 554 31383 592 31417
rect 626 31383 677 31417
rect 433 31344 677 31383
rect 433 31310 448 31344
rect 482 31310 520 31344
rect 554 31310 592 31344
rect 626 31310 677 31344
rect 433 31271 677 31310
rect 433 31237 448 31271
rect 482 31237 520 31271
rect 554 31237 592 31271
rect 626 31237 677 31271
rect 433 31198 677 31237
rect 433 31164 448 31198
rect 482 31164 520 31198
rect 554 31164 592 31198
rect 626 31164 677 31198
rect 433 31125 677 31164
rect 433 31091 448 31125
rect 482 31091 520 31125
rect 554 31091 592 31125
rect 626 31091 677 31125
rect 433 31052 677 31091
rect 433 31018 448 31052
rect 482 31018 520 31052
rect 554 31018 592 31052
rect 626 31018 677 31052
rect 433 30979 677 31018
rect 433 30945 448 30979
rect 482 30945 520 30979
rect 554 30945 592 30979
rect 626 30945 677 30979
rect 433 30906 677 30945
rect 433 30872 448 30906
rect 482 30872 520 30906
rect 554 30872 592 30906
rect 626 30872 677 30906
rect 433 30833 677 30872
rect 433 30799 448 30833
rect 482 30799 520 30833
rect 554 30799 592 30833
rect 626 30799 677 30833
rect 433 30760 677 30799
rect 433 30726 448 30760
rect 482 30726 520 30760
rect 554 30726 592 30760
rect 626 30726 677 30760
rect 433 30687 677 30726
rect 433 30653 448 30687
rect 482 30653 520 30687
rect 554 30653 592 30687
rect 626 30653 677 30687
rect 433 30614 677 30653
rect 433 30580 448 30614
rect 482 30580 520 30614
rect 554 30580 592 30614
rect 626 30580 677 30614
rect 433 30541 677 30580
rect 433 30507 448 30541
rect 482 30507 520 30541
rect 554 30507 592 30541
rect 626 30507 677 30541
rect 433 30468 677 30507
rect 433 30434 448 30468
rect 482 30434 520 30468
rect 554 30434 592 30468
rect 626 30434 677 30468
rect 433 30395 677 30434
rect 433 30361 448 30395
rect 482 30361 520 30395
rect 554 30361 592 30395
rect 626 30361 677 30395
rect 433 30345 677 30361
rect 433 30329 661 30345
tri 661 30329 677 30345 nw
rect 26871 31574 27306 31622
rect 26871 31540 26916 31574
rect 26950 31540 26996 31574
rect 27030 31540 27076 31574
rect 27110 31540 27156 31574
rect 27190 31540 27236 31574
rect 27270 31540 27306 31574
rect 26871 31501 27306 31540
rect 26871 31467 26916 31501
rect 26950 31467 26996 31501
rect 27030 31467 27076 31501
rect 27110 31467 27156 31501
rect 27190 31467 27236 31501
rect 27270 31467 27306 31501
rect 26871 31428 27306 31467
rect 26871 31394 26916 31428
rect 26950 31394 26996 31428
rect 27030 31394 27076 31428
rect 27110 31394 27156 31428
rect 27190 31394 27236 31428
rect 27270 31394 27306 31428
rect 26871 31355 27306 31394
rect 26871 31321 26916 31355
rect 26950 31321 26996 31355
rect 27030 31321 27076 31355
rect 27110 31321 27156 31355
rect 27190 31321 27236 31355
rect 27270 31321 27306 31355
rect 26871 31282 27306 31321
rect 26871 31248 26916 31282
rect 26950 31248 26996 31282
rect 27030 31248 27076 31282
rect 27110 31248 27156 31282
rect 27190 31248 27236 31282
rect 27270 31248 27306 31282
rect 26871 31209 27306 31248
rect 26871 31175 26916 31209
rect 26950 31175 26996 31209
rect 27030 31175 27076 31209
rect 27110 31175 27156 31209
rect 27190 31175 27236 31209
rect 27270 31175 27306 31209
rect 26871 31136 27306 31175
rect 26871 31102 26916 31136
rect 26950 31102 26996 31136
rect 27030 31102 27076 31136
rect 27110 31102 27156 31136
rect 27190 31102 27236 31136
rect 27270 31102 27306 31136
rect 26871 31063 27306 31102
rect 26871 31029 26916 31063
rect 26950 31029 26996 31063
rect 27030 31029 27076 31063
rect 27110 31029 27156 31063
rect 27190 31029 27236 31063
rect 27270 31029 27306 31063
rect 26871 30990 27306 31029
rect 26871 30956 26916 30990
rect 26950 30956 26996 30990
rect 27030 30956 27076 30990
rect 27110 30956 27156 30990
rect 27190 30956 27236 30990
rect 27270 30956 27306 30990
rect 26871 30917 27306 30956
rect 26871 30883 26916 30917
rect 26950 30883 26996 30917
rect 27030 30883 27076 30917
rect 27110 30883 27156 30917
rect 27190 30883 27236 30917
rect 27270 30883 27306 30917
rect 26871 30844 27306 30883
rect 26871 30810 26916 30844
rect 26950 30810 26996 30844
rect 27030 30810 27076 30844
rect 27110 30810 27156 30844
rect 27190 30810 27236 30844
rect 27270 30810 27306 30844
rect 26871 30771 27306 30810
rect 26871 30737 26916 30771
rect 26950 30737 26996 30771
rect 27030 30737 27076 30771
rect 27110 30737 27156 30771
rect 27190 30737 27236 30771
rect 27270 30737 27306 30771
rect 26871 30698 27306 30737
rect 26871 30664 26916 30698
rect 26950 30664 26996 30698
rect 27030 30664 27076 30698
rect 27110 30664 27156 30698
rect 27190 30664 27236 30698
rect 27270 30664 27306 30698
rect 26871 30625 27306 30664
rect 26871 30591 26916 30625
rect 26950 30591 26996 30625
rect 27030 30591 27076 30625
rect 27110 30591 27156 30625
rect 27190 30591 27236 30625
rect 27270 30591 27306 30625
rect 26871 30551 27306 30591
rect 26871 30517 26916 30551
rect 26950 30517 26996 30551
rect 27030 30517 27076 30551
rect 27110 30517 27156 30551
rect 27190 30517 27236 30551
rect 27270 30517 27306 30551
rect 26871 30477 27306 30517
rect 26871 30443 26916 30477
rect 26950 30443 26996 30477
rect 27030 30443 27076 30477
rect 27110 30443 27156 30477
rect 27190 30443 27236 30477
rect 27270 30443 27306 30477
rect 26871 30403 27306 30443
rect 26871 30369 26916 30403
rect 26950 30369 26996 30403
rect 27030 30369 27076 30403
rect 27110 30369 27156 30403
rect 27190 30369 27236 30403
rect 27270 30369 27306 30403
rect 26871 30329 27306 30369
rect 433 30295 627 30329
tri 627 30295 661 30329 nw
rect 26871 30295 26916 30329
rect 26950 30295 26996 30329
rect 27030 30295 27076 30329
rect 27110 30295 27156 30329
rect 27190 30295 27236 30329
rect 27270 30295 27306 30329
rect 433 30275 619 30295
tri 619 30287 627 30295 nw
rect 433 30241 439 30275
rect 473 30241 579 30275
rect 613 30241 619 30275
rect 433 30203 619 30241
rect 433 30169 439 30203
rect 473 30169 579 30203
rect 613 30169 619 30203
rect 433 30131 619 30169
rect 433 30097 439 30131
rect 473 30097 579 30131
rect 613 30097 619 30131
rect 433 30059 619 30097
rect 433 30025 439 30059
rect 473 30025 579 30059
rect 613 30025 619 30059
rect 433 29987 619 30025
rect 433 29953 439 29987
rect 473 29953 579 29987
rect 613 29953 619 29987
rect 433 29915 619 29953
rect 433 29881 439 29915
rect 473 29881 579 29915
rect 613 29881 619 29915
rect 433 29843 619 29881
rect 433 29809 439 29843
rect 473 29809 579 29843
rect 613 29809 619 29843
rect 433 29771 619 29809
rect 433 29737 439 29771
rect 473 29737 579 29771
rect 613 29737 619 29771
rect 433 29699 619 29737
rect 433 29665 439 29699
rect 473 29665 579 29699
rect 613 29665 619 29699
rect 433 29627 619 29665
rect 433 29593 439 29627
rect 473 29593 579 29627
rect 613 29593 619 29627
rect 433 29555 619 29593
rect 433 29521 439 29555
rect 473 29521 579 29555
rect 613 29521 619 29555
rect 433 29483 619 29521
rect 433 29449 439 29483
rect 473 29449 579 29483
rect 613 29449 619 29483
rect 433 29411 619 29449
rect 433 29377 439 29411
rect 473 29377 579 29411
rect 613 29377 619 29411
rect 433 29339 619 29377
rect 433 29305 439 29339
rect 473 29305 579 29339
rect 613 29305 619 29339
rect 433 29267 619 29305
rect 433 29233 439 29267
rect 473 29233 579 29267
rect 613 29233 619 29267
rect 433 29195 619 29233
rect 433 29161 439 29195
rect 473 29161 579 29195
rect 613 29161 619 29195
rect 433 29123 619 29161
rect 433 29089 439 29123
rect 473 29089 579 29123
rect 613 29089 619 29123
rect 433 29051 619 29089
rect 433 29017 439 29051
rect 473 29017 579 29051
rect 613 29017 619 29051
rect 433 28979 619 29017
rect 433 28945 439 28979
rect 473 28945 579 28979
rect 613 28945 619 28979
rect 433 28907 619 28945
rect 433 28873 439 28907
rect 473 28873 579 28907
rect 613 28873 619 28907
rect 433 28835 619 28873
rect 433 28801 439 28835
rect 473 28801 579 28835
rect 613 28801 619 28835
rect 433 28763 619 28801
rect 433 28729 439 28763
rect 473 28729 579 28763
rect 613 28729 619 28763
rect 433 28691 619 28729
rect 433 28657 439 28691
rect 473 28657 579 28691
rect 613 28657 619 28691
rect 433 28619 619 28657
rect 433 28585 439 28619
rect 473 28585 579 28619
rect 613 28585 619 28619
rect 433 28547 619 28585
rect 433 28513 439 28547
rect 473 28513 579 28547
rect 613 28513 619 28547
rect 433 28475 619 28513
rect 433 28441 439 28475
rect 473 28441 579 28475
rect 613 28441 619 28475
rect 433 28403 619 28441
rect 433 28369 439 28403
rect 473 28369 579 28403
rect 613 28369 619 28403
rect 433 28331 619 28369
rect 433 28297 439 28331
rect 473 28297 579 28331
rect 613 28297 619 28331
rect 433 28259 619 28297
rect 26871 30255 27306 30295
rect 26871 30221 26916 30255
rect 26950 30221 26996 30255
rect 27030 30221 27076 30255
rect 27110 30221 27156 30255
rect 27190 30221 27236 30255
rect 27270 30221 27306 30255
rect 26871 30181 27306 30221
rect 26871 30147 26916 30181
rect 26950 30147 26996 30181
rect 27030 30147 27076 30181
rect 27110 30147 27156 30181
rect 27190 30147 27236 30181
rect 27270 30147 27306 30181
rect 26871 30107 27306 30147
rect 26871 30073 26916 30107
rect 26950 30073 26996 30107
rect 27030 30073 27076 30107
rect 27110 30073 27156 30107
rect 27190 30073 27236 30107
rect 27270 30073 27306 30107
rect 26871 30033 27306 30073
rect 26871 29999 26916 30033
rect 26950 29999 26996 30033
rect 27030 29999 27076 30033
rect 27110 29999 27156 30033
rect 27190 29999 27236 30033
rect 27270 29999 27306 30033
rect 26871 29959 27306 29999
rect 26871 29925 26916 29959
rect 26950 29925 26996 29959
rect 27030 29925 27076 29959
rect 27110 29925 27156 29959
rect 27190 29925 27236 29959
rect 27270 29925 27306 29959
rect 26871 29885 27306 29925
rect 26871 29851 26916 29885
rect 26950 29851 26996 29885
rect 27030 29851 27076 29885
rect 27110 29851 27156 29885
rect 27190 29851 27236 29885
rect 27270 29851 27306 29885
rect 26871 29811 27306 29851
rect 26871 29777 26916 29811
rect 26950 29777 26996 29811
rect 27030 29777 27076 29811
rect 27110 29777 27156 29811
rect 27190 29777 27236 29811
rect 27270 29777 27306 29811
rect 26871 29737 27306 29777
rect 26871 29703 26916 29737
rect 26950 29703 26996 29737
rect 27030 29703 27076 29737
rect 27110 29703 27156 29737
rect 27190 29703 27236 29737
rect 27270 29703 27306 29737
rect 26871 29663 27306 29703
rect 26871 29629 26916 29663
rect 26950 29629 26996 29663
rect 27030 29629 27076 29663
rect 27110 29629 27156 29663
rect 27190 29629 27236 29663
rect 27270 29629 27306 29663
rect 26871 29589 27306 29629
rect 26871 29555 26916 29589
rect 26950 29555 26996 29589
rect 27030 29555 27076 29589
rect 27110 29555 27156 29589
rect 27190 29555 27236 29589
rect 27270 29555 27306 29589
rect 26871 29515 27306 29555
rect 26871 29481 26916 29515
rect 26950 29481 26996 29515
rect 27030 29481 27076 29515
rect 27110 29481 27156 29515
rect 27190 29481 27236 29515
rect 27270 29481 27306 29515
rect 26871 29441 27306 29481
rect 26871 29407 26916 29441
rect 26950 29407 26996 29441
rect 27030 29407 27076 29441
rect 27110 29407 27156 29441
rect 27190 29407 27236 29441
rect 27270 29407 27306 29441
rect 26871 29367 27306 29407
rect 26871 29333 26916 29367
rect 26950 29333 26996 29367
rect 27030 29333 27076 29367
rect 27110 29333 27156 29367
rect 27190 29333 27236 29367
rect 27270 29333 27306 29367
rect 26871 29293 27306 29333
rect 26871 29259 26916 29293
rect 26950 29259 26996 29293
rect 27030 29259 27076 29293
rect 27110 29259 27156 29293
rect 27190 29259 27236 29293
rect 27270 29259 27306 29293
rect 26871 29219 27306 29259
rect 26871 29185 26916 29219
rect 26950 29185 26996 29219
rect 27030 29185 27076 29219
rect 27110 29185 27156 29219
rect 27190 29185 27236 29219
rect 27270 29185 27306 29219
rect 26871 29145 27306 29185
rect 26871 29111 26916 29145
rect 26950 29111 26996 29145
rect 27030 29111 27076 29145
rect 27110 29111 27156 29145
rect 27190 29111 27236 29145
rect 27270 29111 27306 29145
rect 26871 29071 27306 29111
rect 26871 29037 26916 29071
rect 26950 29037 26996 29071
rect 27030 29037 27076 29071
rect 27110 29037 27156 29071
rect 27190 29037 27236 29071
rect 27270 29037 27306 29071
rect 26871 28997 27306 29037
rect 26871 28963 26916 28997
rect 26950 28963 26996 28997
rect 27030 28963 27076 28997
rect 27110 28963 27156 28997
rect 27190 28963 27236 28997
rect 27270 28963 27306 28997
rect 26871 28923 27306 28963
rect 26871 28889 26916 28923
rect 26950 28889 26996 28923
rect 27030 28889 27076 28923
rect 27110 28889 27156 28923
rect 27190 28889 27236 28923
rect 27270 28889 27306 28923
rect 26871 28849 27306 28889
rect 26871 28815 26916 28849
rect 26950 28815 26996 28849
rect 27030 28815 27076 28849
rect 27110 28815 27156 28849
rect 27190 28815 27236 28849
rect 27270 28815 27306 28849
rect 26871 28775 27306 28815
rect 26871 28741 26916 28775
rect 26950 28741 26996 28775
rect 27030 28741 27076 28775
rect 27110 28741 27156 28775
rect 27190 28741 27236 28775
rect 27270 28741 27306 28775
rect 26871 28701 27306 28741
rect 26871 28667 26916 28701
rect 26950 28667 26996 28701
rect 27030 28667 27076 28701
rect 27110 28667 27156 28701
rect 27190 28667 27236 28701
rect 27270 28667 27306 28701
rect 26871 28627 27306 28667
rect 26871 28593 26916 28627
rect 26950 28593 26996 28627
rect 27030 28593 27076 28627
rect 27110 28593 27156 28627
rect 27190 28593 27236 28627
rect 27270 28593 27306 28627
rect 26871 28553 27306 28593
rect 26871 28519 26916 28553
rect 26950 28519 26996 28553
rect 27030 28519 27076 28553
rect 27110 28519 27156 28553
rect 27190 28519 27236 28553
rect 27270 28519 27306 28553
rect 26871 28507 27306 28519
rect 26871 28283 26890 28507
tri 26890 28283 27114 28507 nw
rect 433 28225 439 28259
rect 473 28225 579 28259
rect 613 28225 619 28259
rect 433 28187 619 28225
rect 433 28153 439 28187
rect 473 28153 579 28187
rect 613 28153 619 28187
rect 433 28115 619 28153
rect 433 28081 439 28115
rect 473 28081 579 28115
rect 613 28081 619 28115
rect 433 28043 619 28081
rect 433 28009 439 28043
rect 473 28009 579 28043
rect 613 28009 619 28043
rect 433 27971 619 28009
rect 433 27937 439 27971
rect 473 27937 579 27971
rect 613 27937 619 27971
rect 433 27899 619 27937
rect 433 27865 439 27899
rect 473 27865 579 27899
rect 613 27865 619 27899
rect 433 27827 619 27865
rect 433 27793 439 27827
rect 473 27793 579 27827
rect 613 27793 619 27827
rect 433 27755 619 27793
rect 433 27721 439 27755
rect 473 27721 579 27755
rect 613 27721 619 27755
rect 433 27683 619 27721
rect 433 27649 439 27683
rect 473 27649 579 27683
rect 613 27649 619 27683
rect 433 27611 619 27649
rect 433 27577 439 27611
rect 473 27577 579 27611
rect 613 27577 619 27611
rect 433 27539 619 27577
rect 433 27505 439 27539
rect 473 27505 579 27539
rect 613 27505 619 27539
rect 433 27467 619 27505
rect 433 27433 439 27467
rect 473 27433 579 27467
rect 613 27433 619 27467
rect 433 27395 619 27433
rect 433 27361 439 27395
rect 473 27361 579 27395
rect 613 27361 619 27395
rect 433 27323 619 27361
rect 433 27289 439 27323
rect 473 27289 579 27323
rect 613 27289 619 27323
rect 433 27251 619 27289
rect 433 27217 439 27251
rect 473 27217 579 27251
rect 613 27217 619 27251
rect 433 27179 619 27217
rect 433 27145 439 27179
rect 473 27145 579 27179
rect 613 27145 619 27179
rect 433 27107 619 27145
rect 433 27073 439 27107
rect 473 27073 579 27107
rect 613 27073 619 27107
rect 433 27035 619 27073
rect 433 27001 439 27035
rect 473 27001 579 27035
rect 613 27001 619 27035
rect 433 26963 619 27001
rect 433 26929 439 26963
rect 473 26929 579 26963
rect 613 26929 619 26963
rect 433 26891 619 26929
rect 433 26857 439 26891
rect 473 26857 579 26891
rect 613 26857 619 26891
rect 433 26819 619 26857
rect 433 26785 439 26819
rect 473 26785 579 26819
rect 613 26785 619 26819
rect 433 26747 619 26785
rect 433 26713 439 26747
rect 473 26713 579 26747
rect 613 26713 619 26747
rect 433 26675 619 26713
rect 433 26641 439 26675
rect 473 26641 579 26675
rect 613 26641 619 26675
rect 433 26603 619 26641
rect 433 26569 439 26603
rect 473 26569 579 26603
rect 613 26569 619 26603
rect 433 26530 619 26569
rect 433 26496 439 26530
rect 473 26496 579 26530
rect 613 26496 619 26530
rect 433 26457 619 26496
rect 433 26423 439 26457
rect 473 26423 579 26457
rect 613 26423 619 26457
rect 433 26384 619 26423
rect 433 26350 439 26384
rect 473 26350 579 26384
rect 613 26350 619 26384
rect 433 26311 619 26350
rect 433 26277 439 26311
rect 473 26277 579 26311
rect 613 26277 619 26311
rect 433 26238 619 26277
rect 433 26204 439 26238
rect 473 26204 579 26238
rect 613 26204 619 26238
rect 433 26165 619 26204
rect 433 26131 439 26165
rect 473 26131 579 26165
rect 613 26131 619 26165
tri 397 26083 433 26119 se
rect 433 26083 619 26131
tri 619 26083 655 26119 sw
rect -2267 26071 -1407 26079
rect -2267 26037 -2255 26071
rect -2221 26037 -2182 26071
rect -2148 26037 -2109 26071
rect -2075 26037 -2036 26071
rect -2002 26037 -1963 26071
rect -1929 26037 -1890 26071
rect -1856 26037 -1817 26071
rect -1783 26037 -1744 26071
rect -1710 26037 -1671 26071
rect -1637 26037 -1598 26071
rect -1564 26037 -1525 26071
rect -1491 26037 -1453 26071
rect -1419 26037 -1407 26071
rect -2267 25997 -1407 26037
rect -2267 25963 -2255 25997
rect -2221 25963 -2182 25997
rect -2148 25963 -2109 25997
rect -2075 25963 -2036 25997
rect -2002 25963 -1963 25997
rect -1929 25963 -1890 25997
rect -1856 25963 -1817 25997
rect -1783 25963 -1744 25997
rect -1710 25963 -1671 25997
rect -1637 25963 -1598 25997
rect -1564 25963 -1525 25997
rect -1491 25963 -1453 25997
rect -1419 25963 -1407 25997
rect -2267 25923 -1407 25963
rect -2267 25889 -2255 25923
rect -2221 25889 -2182 25923
rect -2148 25889 -2109 25923
rect -2075 25889 -2036 25923
rect -2002 25889 -1963 25923
rect -1929 25889 -1890 25923
rect -1856 25889 -1817 25923
rect -1783 25889 -1744 25923
rect -1710 25889 -1671 25923
rect -1637 25889 -1598 25923
rect -1564 25889 -1525 25923
rect -1491 25889 -1453 25923
rect -1419 25889 -1407 25923
rect -2267 25849 -1407 25889
rect -2267 25815 -2255 25849
rect -2221 25815 -2182 25849
rect -2148 25815 -2109 25849
rect -2075 25815 -2036 25849
rect -2002 25815 -1963 25849
rect -1929 25815 -1890 25849
rect -1856 25815 -1817 25849
rect -1783 25815 -1744 25849
rect -1710 25815 -1671 25849
rect -1637 25815 -1598 25849
rect -1564 25815 -1525 25849
rect -1491 25815 -1453 25849
rect -1419 25815 -1407 25849
rect -2267 25775 -1407 25815
rect -2267 25741 -2255 25775
rect -2221 25741 -2182 25775
rect -2148 25741 -2109 25775
rect -2075 25741 -2036 25775
rect -2002 25741 -1963 25775
rect -1929 25741 -1890 25775
rect -1856 25741 -1817 25775
rect -1783 25741 -1744 25775
rect -1710 25741 -1671 25775
rect -1637 25741 -1598 25775
rect -1564 25741 -1525 25775
rect -1491 25741 -1453 25775
rect -1419 25741 -1407 25775
rect -2267 25701 -1407 25741
rect -2267 25667 -2255 25701
rect -2221 25667 -2182 25701
rect -2148 25667 -2109 25701
rect -2075 25667 -2036 25701
rect -2002 25667 -1963 25701
rect -1929 25667 -1890 25701
rect -1856 25667 -1817 25701
rect -1783 25667 -1744 25701
rect -1710 25667 -1671 25701
rect -1637 25667 -1598 25701
rect -1564 25667 -1525 25701
rect -1491 25667 -1453 25701
rect -1419 25667 -1407 25701
rect -2267 25627 -1407 25667
rect -2267 25593 -2255 25627
rect -2221 25593 -2182 25627
rect -2148 25593 -2109 25627
rect -2075 25593 -2036 25627
rect -2002 25593 -1963 25627
rect -1929 25593 -1890 25627
rect -1856 25593 -1817 25627
rect -1783 25593 -1744 25627
rect -1710 25593 -1671 25627
rect -1637 25593 -1598 25627
rect -1564 25593 -1525 25627
rect -1491 25593 -1453 25627
rect -1419 25593 -1407 25627
rect -2267 25585 -1407 25593
rect -1193 25915 2691 25923
rect -1193 25881 -1181 25915
rect -1147 25881 -1108 25915
rect -1074 25881 -1035 25915
rect -1001 25881 -962 25915
rect -928 25881 -889 25915
rect -855 25881 -816 25915
rect -782 25881 -743 25915
rect -709 25881 -670 25915
rect -636 25881 -597 25915
rect -563 25881 -524 25915
rect -490 25881 -451 25915
rect -1193 25843 -451 25881
rect -1193 25809 -1181 25843
rect -1147 25809 -1108 25843
rect -1074 25809 -1035 25843
rect -1001 25809 -962 25843
rect -928 25809 -889 25843
rect -855 25809 -816 25843
rect -782 25809 -743 25843
rect -709 25809 -670 25843
rect -636 25809 -597 25843
rect -563 25809 -524 25843
rect -490 25809 -451 25843
rect -1193 25771 -451 25809
rect -1193 25737 -1181 25771
rect -1147 25737 -1108 25771
rect -1074 25737 -1035 25771
rect -1001 25737 -962 25771
rect -928 25737 -889 25771
rect -855 25737 -816 25771
rect -782 25737 -743 25771
rect -709 25737 -670 25771
rect -636 25737 -597 25771
rect -563 25737 -524 25771
rect -490 25737 -451 25771
rect -1193 25699 -451 25737
rect -1193 25665 -1181 25699
rect -1147 25665 -1108 25699
rect -1074 25665 -1035 25699
rect -1001 25665 -962 25699
rect -928 25665 -889 25699
rect -855 25665 -816 25699
rect -782 25665 -743 25699
rect -709 25665 -670 25699
rect -636 25665 -597 25699
rect -563 25665 -524 25699
rect -490 25665 -451 25699
rect -1193 25627 -451 25665
rect -1193 25593 -1181 25627
rect -1147 25593 -1108 25627
rect -1074 25593 -1035 25627
rect -1001 25593 -962 25627
rect -928 25593 -889 25627
rect -855 25593 -816 25627
rect -782 25593 -743 25627
rect -709 25593 -670 25627
rect -636 25593 -597 25627
rect -563 25593 -524 25627
rect -490 25593 -451 25627
rect 2679 25593 2691 25915
rect -1193 25585 2691 25593
tri 31968 23695 32040 23767 sw
tri 31756 23645 31806 23695 ne
rect 31806 23689 31891 23695
rect 31968 23689 32040 23695
tri 32040 23689 32046 23695 sw
rect 31806 23659 32046 23689
tri 32046 23659 32076 23689 sw
rect 31806 23645 32076 23659
tri 31806 23611 31840 23645 ne
rect 31840 23611 31932 23645
rect 31966 23611 32020 23645
rect 32054 23611 32076 23645
tri 31840 23574 31877 23611 ne
rect 31877 23570 32076 23611
rect 31877 23536 31932 23570
rect 31966 23536 32020 23570
rect 32054 23536 32076 23570
rect 31877 23495 32076 23536
rect 31877 23461 31932 23495
rect 31966 23461 32020 23495
rect 32054 23461 32076 23495
rect 17771 23429 18019 23441
rect 17771 23395 17778 23429
rect 17812 23395 17878 23429
rect 17912 23395 17978 23429
rect 18012 23395 18019 23429
rect 17771 23356 18019 23395
rect 17771 23322 17778 23356
rect 17812 23322 17878 23356
rect 17912 23322 17978 23356
rect 18012 23322 18019 23356
rect 31877 23420 32076 23461
rect 31877 23386 31932 23420
rect 31966 23386 32020 23420
rect 32054 23386 32076 23420
rect 31877 23345 32076 23386
rect 17771 23283 18019 23322
tri 31862 23311 31877 23326 se
rect 31877 23311 31932 23345
rect 31966 23311 32020 23345
rect 32054 23311 32076 23345
rect 17771 23249 17778 23283
rect 17812 23249 17878 23283
rect 17912 23249 17978 23283
rect 18012 23249 18019 23283
tri 31821 23270 31862 23311 se
rect 31862 23270 32076 23311
rect 17771 23210 18019 23249
tri 31787 23236 31821 23270 se
rect 31821 23236 31932 23270
rect 31966 23236 32020 23270
rect 32054 23236 32076 23270
rect 17771 23176 17778 23210
rect 17812 23176 17878 23210
rect 17912 23176 17978 23210
rect 18012 23176 18019 23210
rect 17771 23137 18019 23176
rect 17771 23103 17778 23137
rect 17812 23103 17878 23137
rect 17912 23103 17978 23137
rect 18012 23103 18019 23137
rect 17771 23064 18019 23103
rect 17771 23030 17778 23064
rect 17812 23030 17878 23064
rect 17912 23030 17978 23064
rect 18012 23030 18019 23064
rect 17771 22991 18019 23030
rect 17771 22957 17778 22991
rect 17812 22957 17878 22991
rect 17912 22957 17978 22991
rect 18012 22957 18019 22991
rect 17771 22918 18019 22957
rect 17771 22884 17778 22918
rect 17812 22884 17878 22918
rect 17912 22884 17978 22918
rect 18012 22884 18019 22918
rect 17771 22845 18019 22884
rect 17771 22811 17778 22845
rect 17812 22811 17878 22845
rect 17912 22811 17978 22845
rect 18012 22811 18019 22845
rect 17771 22772 18019 22811
rect 17771 22738 17778 22772
rect 17812 22738 17878 22772
rect 17912 22738 17978 22772
rect 18012 22738 18019 22772
rect 17771 22699 18019 22738
rect 17771 22665 17778 22699
rect 17812 22665 17878 22699
rect 17912 22665 17978 22699
rect 18012 22665 18019 22699
rect 17771 22626 18019 22665
rect 17771 22592 17778 22626
rect 17812 22592 17878 22626
rect 17912 22592 17978 22626
rect 18012 22592 18019 22626
rect 17771 22553 18019 22592
rect 17771 22519 17778 22553
rect 17812 22519 17878 22553
rect 17912 22519 17978 22553
rect 18012 22519 18019 22553
rect 17771 22480 18019 22519
rect 17771 22446 17778 22480
rect 17812 22446 17878 22480
rect 17912 22446 17978 22480
rect 18012 22446 18019 22480
rect 17771 22407 18019 22446
rect 17771 22373 17778 22407
rect 17812 22373 17878 22407
rect 17912 22373 17978 22407
rect 18012 22373 18019 22407
rect 17771 22334 18019 22373
rect 17771 22300 17778 22334
rect 17812 22300 17878 22334
rect 17912 22300 17978 22334
rect 18012 22300 18019 22334
rect 17771 22261 18019 22300
rect 17771 22227 17778 22261
rect 17812 22227 17878 22261
rect 17912 22227 17978 22261
rect 18012 22227 18019 22261
rect 17771 22188 18019 22227
rect 17771 22154 17778 22188
rect 17812 22154 17878 22188
rect 17912 22154 17978 22188
rect 18012 22154 18019 22188
rect 17771 22115 18019 22154
rect 17771 22081 17778 22115
rect 17812 22081 17878 22115
rect 17912 22081 17978 22115
rect 18012 22081 18019 22115
rect 17771 22042 18019 22081
rect 17771 22008 17778 22042
rect 17812 22008 17878 22042
rect 17912 22008 17978 22042
rect 18012 22008 18019 22042
rect 17771 21968 18019 22008
rect 17771 21934 17778 21968
rect 17812 21934 17878 21968
rect 17912 21934 17978 21968
rect 18012 21934 18019 21968
rect 17771 21894 18019 21934
rect 17771 21860 17778 21894
rect 17812 21860 17878 21894
rect 17912 21860 17978 21894
rect 18012 21860 18019 21894
rect 17771 21820 18019 21860
rect 17771 21786 17778 21820
rect 17812 21786 17878 21820
rect 17912 21786 17978 21820
rect 18012 21786 18019 21820
rect 17771 21746 18019 21786
rect 17771 21712 17778 21746
rect 17812 21712 17878 21746
rect 17912 21712 17978 21746
rect 18012 21712 18019 21746
rect 17771 21672 18019 21712
rect 17771 21638 17778 21672
rect 17812 21638 17878 21672
rect 17912 21638 17978 21672
rect 18012 21638 18019 21672
rect 17771 21598 18019 21638
rect 17771 21564 17778 21598
rect 17812 21564 17878 21598
rect 17912 21564 17978 21598
rect 18012 21564 18019 21598
rect 17771 21524 18019 21564
rect 17771 21490 17778 21524
rect 17812 21490 17878 21524
rect 17912 21490 17978 21524
rect 18012 21490 18019 21524
rect 17771 21450 18019 21490
rect 17771 21416 17778 21450
rect 17812 21416 17878 21450
rect 17912 21416 17978 21450
rect 18012 21416 18019 21450
rect 17771 21376 18019 21416
rect 17771 21342 17778 21376
rect 17812 21342 17878 21376
rect 17912 21342 17978 21376
rect 18012 21342 18019 21376
rect 17771 21302 18019 21342
rect 17771 21268 17778 21302
rect 17812 21268 17878 21302
rect 17912 21268 17978 21302
rect 18012 21268 18019 21302
rect 17771 21228 18019 21268
rect 17771 21194 17778 21228
rect 17812 21194 17878 21228
rect 17912 21194 17978 21228
rect 18012 21194 18019 21228
rect 17771 21154 18019 21194
rect 17771 21120 17778 21154
rect 17812 21120 17878 21154
rect 17912 21120 17978 21154
rect 18012 21120 18019 21154
rect 17771 21080 18019 21120
rect 17771 21046 17778 21080
rect 17812 21046 17878 21080
rect 17912 21046 17978 21080
rect 18012 21046 18019 21080
rect 17771 21006 18019 21046
rect 17771 20972 17778 21006
rect 17812 20972 17878 21006
rect 17912 20972 17978 21006
rect 18012 20972 18019 21006
rect 17771 20932 18019 20972
tri 31718 23167 31787 23236 se
rect 31787 23167 32076 23236
rect 31718 23155 32076 23167
rect 31718 23121 31724 23155
rect 31758 23121 31802 23155
rect 31836 23121 31880 23155
rect 31914 23121 31958 23155
rect 31992 23121 32036 23155
rect 32070 23121 32076 23155
rect 31718 23081 32076 23121
rect 31718 23047 31724 23081
rect 31758 23047 31802 23081
rect 31836 23047 31880 23081
rect 31914 23047 31958 23081
rect 31992 23047 32036 23081
rect 32070 23047 32076 23081
rect 31718 23007 32076 23047
rect 31718 22973 31724 23007
rect 31758 22973 31802 23007
rect 31836 22973 31880 23007
rect 31914 22973 31958 23007
rect 31992 22973 32036 23007
rect 32070 22973 32076 23007
rect 31718 22933 32076 22973
rect 31718 22899 31724 22933
rect 31758 22899 31802 22933
rect 31836 22899 31880 22933
rect 31914 22899 31958 22933
rect 31992 22899 32036 22933
rect 32070 22899 32076 22933
rect 31718 22859 32076 22899
rect 31718 22825 31724 22859
rect 31758 22825 31802 22859
rect 31836 22825 31880 22859
rect 31914 22825 31958 22859
rect 31992 22825 32036 22859
rect 32070 22825 32076 22859
rect 31718 22785 32076 22825
rect 31718 22751 31724 22785
rect 31758 22751 31802 22785
rect 31836 22751 31880 22785
rect 31914 22751 31958 22785
rect 31992 22751 32036 22785
rect 32070 22751 32076 22785
rect 31718 22711 32076 22751
rect 31718 22677 31724 22711
rect 31758 22677 31802 22711
rect 31836 22677 31880 22711
rect 31914 22677 31958 22711
rect 31992 22677 32036 22711
rect 32070 22677 32076 22711
rect 31718 22637 32076 22677
rect 31718 22603 31724 22637
rect 31758 22603 31802 22637
rect 31836 22603 31880 22637
rect 31914 22603 31958 22637
rect 31992 22603 32036 22637
rect 32070 22603 32076 22637
rect 31718 22563 32076 22603
rect 31718 22529 31724 22563
rect 31758 22529 31802 22563
rect 31836 22529 31880 22563
rect 31914 22529 31958 22563
rect 31992 22529 32036 22563
rect 32070 22529 32076 22563
rect 31718 22489 32076 22529
rect 31718 22455 31724 22489
rect 31758 22455 31802 22489
rect 31836 22455 31880 22489
rect 31914 22455 31958 22489
rect 31992 22455 32036 22489
rect 32070 22455 32076 22489
rect 31718 22415 32076 22455
rect 31718 22381 31724 22415
rect 31758 22381 31802 22415
rect 31836 22381 31880 22415
rect 31914 22381 31958 22415
rect 31992 22381 32036 22415
rect 32070 22381 32076 22415
rect 31718 22341 32076 22381
rect 31718 22307 31724 22341
rect 31758 22307 31802 22341
rect 31836 22307 31880 22341
rect 31914 22307 31958 22341
rect 31992 22307 32036 22341
rect 32070 22307 32076 22341
rect 31718 22267 32076 22307
rect 31718 22233 31724 22267
rect 31758 22233 31802 22267
rect 31836 22233 31880 22267
rect 31914 22233 31958 22267
rect 31992 22233 32036 22267
rect 32070 22233 32076 22267
rect 31718 22193 32076 22233
rect 31718 22159 31724 22193
rect 31758 22159 31802 22193
rect 31836 22159 31880 22193
rect 31914 22159 31958 22193
rect 31992 22159 32036 22193
rect 32070 22159 32076 22193
rect 31718 22119 32076 22159
rect 31718 22085 31724 22119
rect 31758 22085 31802 22119
rect 31836 22085 31880 22119
rect 31914 22085 31958 22119
rect 31992 22085 32036 22119
rect 32070 22085 32076 22119
rect 31718 22045 32076 22085
rect 31718 22011 31724 22045
rect 31758 22011 31802 22045
rect 31836 22011 31880 22045
rect 31914 22011 31958 22045
rect 31992 22011 32036 22045
rect 32070 22011 32076 22045
rect 31718 21971 32076 22011
rect 31718 21937 31724 21971
rect 31758 21937 31802 21971
rect 31836 21937 31880 21971
rect 31914 21937 31958 21971
rect 31992 21937 32036 21971
rect 32070 21937 32076 21971
rect 31718 21897 32076 21937
rect 31718 21863 31724 21897
rect 31758 21863 31802 21897
rect 31836 21863 31880 21897
rect 31914 21863 31958 21897
rect 31992 21863 32036 21897
rect 32070 21863 32076 21897
rect 31718 21823 32076 21863
rect 31718 21789 31724 21823
rect 31758 21789 31802 21823
rect 31836 21789 31880 21823
rect 31914 21789 31958 21823
rect 31992 21789 32036 21823
rect 32070 21789 32076 21823
rect 31718 21749 32076 21789
rect 31718 21715 31724 21749
rect 31758 21715 31802 21749
rect 31836 21715 31880 21749
rect 31914 21715 31958 21749
rect 31992 21715 32036 21749
rect 32070 21715 32076 21749
rect 31718 21675 32076 21715
rect 31718 21641 31724 21675
rect 31758 21641 31802 21675
rect 31836 21641 31880 21675
rect 31914 21641 31958 21675
rect 31992 21641 32036 21675
rect 32070 21641 32076 21675
rect 31718 21601 32076 21641
rect 31718 21567 31724 21601
rect 31758 21567 31802 21601
rect 31836 21567 31880 21601
rect 31914 21567 31958 21601
rect 31992 21567 32036 21601
rect 32070 21567 32076 21601
rect 31718 21527 32076 21567
rect 31718 21493 31724 21527
rect 31758 21493 31802 21527
rect 31836 21493 31880 21527
rect 31914 21493 31958 21527
rect 31992 21493 32036 21527
rect 32070 21493 32076 21527
rect 31718 21452 32076 21493
rect 31718 21418 31724 21452
rect 31758 21418 31802 21452
rect 31836 21418 31880 21452
rect 31914 21418 31958 21452
rect 31992 21418 32036 21452
rect 32070 21418 32076 21452
rect 31718 21377 32076 21418
rect 31718 21343 31724 21377
rect 31758 21343 31802 21377
rect 31836 21343 31880 21377
rect 31914 21343 31958 21377
rect 31992 21343 32036 21377
rect 32070 21343 32076 21377
rect 31718 21302 32076 21343
rect 31718 21268 31724 21302
rect 31758 21268 31802 21302
rect 31836 21268 31880 21302
rect 31914 21268 31958 21302
rect 31992 21268 32036 21302
rect 32070 21268 32076 21302
rect 31718 21227 32076 21268
rect 31718 21193 31724 21227
rect 31758 21193 31802 21227
rect 31836 21193 31880 21227
rect 31914 21193 31958 21227
rect 31992 21193 32036 21227
rect 32070 21193 32076 21227
rect 31718 21152 32076 21193
rect 31718 21118 31724 21152
rect 31758 21118 31802 21152
rect 31836 21118 31880 21152
rect 31914 21118 31958 21152
rect 31992 21118 32036 21152
rect 32070 21118 32076 21152
rect 31718 21077 32076 21118
rect 31718 21043 31724 21077
rect 31758 21043 31802 21077
rect 31836 21043 31880 21077
rect 31914 21043 31958 21077
rect 31992 21043 32036 21077
rect 32070 21043 32076 21077
rect 31718 21002 32076 21043
rect 31718 20968 31724 21002
rect 31758 20968 31802 21002
rect 31836 20968 31880 21002
rect 31914 20968 31958 21002
rect 31992 20968 32036 21002
rect 32070 20968 32076 21002
rect 31718 20956 32076 20968
rect 17771 20898 17778 20932
rect 17812 20898 17878 20932
rect 17912 20898 17978 20932
rect 18012 20898 18019 20932
rect 17771 20858 18019 20898
rect 17771 20824 17778 20858
rect 17812 20824 17878 20858
rect 17912 20824 17978 20858
rect 18012 20824 18019 20858
rect 17771 20784 18019 20824
rect 17771 20750 17778 20784
rect 17812 20750 17878 20784
rect 17912 20750 17978 20784
rect 18012 20750 18019 20784
rect 17771 20710 18019 20750
rect 17771 20676 17778 20710
rect 17812 20676 17878 20710
rect 17912 20676 17978 20710
rect 18012 20676 18019 20710
rect 17771 20636 18019 20676
rect 17771 20602 17778 20636
rect 17812 20602 17878 20636
rect 17912 20602 17978 20636
rect 18012 20602 18019 20636
rect 17771 20562 18019 20602
rect 17771 20528 17778 20562
rect 17812 20528 17878 20562
rect 17912 20528 17978 20562
rect 18012 20528 18019 20562
rect 17771 20488 18019 20528
rect 17771 20454 17778 20488
rect 17812 20454 17878 20488
rect 17912 20454 17978 20488
rect 18012 20454 18019 20488
rect 17771 20414 18019 20454
rect 17771 20380 17778 20414
rect 17812 20380 17878 20414
rect 17912 20380 17978 20414
rect 18012 20380 18019 20414
rect 17771 20340 18019 20380
rect 17771 20306 17778 20340
rect 17812 20306 17878 20340
rect 17912 20306 17978 20340
rect 18012 20306 18019 20340
rect 17771 20294 18019 20306
rect -2301 13347 -1506 13353
rect -2301 13313 -2289 13347
rect -2255 13313 -2215 13347
rect -2181 13313 -2141 13347
rect -2107 13313 -2067 13347
rect -2033 13313 -1993 13347
rect -1959 13313 -1919 13347
rect -1885 13313 -1845 13347
rect -1811 13313 -1771 13347
rect -1737 13313 -1698 13347
rect -1664 13313 -1625 13347
rect -1591 13313 -1552 13347
rect -1518 13313 -1506 13347
rect -2301 13263 -1506 13313
rect -2301 13229 -2289 13263
rect -2255 13229 -2215 13263
rect -2181 13229 -2141 13263
rect -2107 13229 -2067 13263
rect -2033 13229 -1993 13263
rect -1959 13229 -1919 13263
rect -1885 13229 -1845 13263
rect -1811 13229 -1771 13263
rect -1737 13229 -1698 13263
rect -1664 13229 -1625 13263
rect -1591 13229 -1552 13263
rect -1518 13229 -1506 13263
rect -2301 13223 -1506 13229
rect 15779 7802 15813 8070
rect 28748 7439 31001 7445
rect 28748 7405 28826 7439
rect 28860 7405 28899 7439
rect 28933 7405 28972 7439
rect 29006 7405 29045 7439
rect 29079 7405 29117 7439
rect 29151 7405 29189 7439
rect 29223 7405 29261 7439
rect 29295 7405 29333 7439
rect 29367 7405 29405 7439
rect 29439 7405 29477 7439
rect 29511 7405 29549 7439
rect 29583 7405 29621 7439
rect 29655 7405 29693 7439
rect 29727 7405 29765 7439
rect 29799 7405 29837 7439
rect 29871 7405 29909 7439
rect 29943 7405 29981 7439
rect 30015 7405 30053 7439
rect 30087 7405 30125 7439
rect 30159 7405 30197 7439
rect 30231 7405 30269 7439
rect 30303 7405 30341 7439
rect 30375 7405 30413 7439
rect 30447 7405 30485 7439
rect 30519 7405 30557 7439
rect 30591 7405 30629 7439
rect 30663 7405 30701 7439
rect 30735 7405 30773 7439
rect 30807 7405 30845 7439
rect 30879 7405 30917 7439
rect 30951 7405 31001 7439
rect 28748 7364 31001 7405
rect 28748 7330 28754 7364
rect 28788 7330 31001 7364
rect 28748 7327 31001 7330
rect 28748 7293 28866 7327
rect 28900 7293 28940 7327
rect 28974 7293 29014 7327
rect 29048 7293 29088 7327
rect 29122 7293 29162 7327
rect 29196 7293 29236 7327
rect 29270 7293 29310 7327
rect 29344 7293 29384 7327
rect 29418 7293 29457 7327
rect 29491 7293 29530 7327
rect 29564 7293 29603 7327
rect 29637 7293 29676 7327
rect 29710 7293 29749 7327
rect 29783 7293 29822 7327
rect 29856 7293 29895 7327
rect 29929 7293 29968 7327
rect 30002 7293 30041 7327
rect 30075 7293 30114 7327
rect 30148 7293 30187 7327
rect 30221 7293 30260 7327
rect 30294 7293 30333 7327
rect 30367 7293 30406 7327
rect 30440 7293 30479 7327
rect 30513 7293 30552 7327
rect 30586 7293 30625 7327
rect 30659 7293 30698 7327
rect 30732 7293 30771 7327
rect 30805 7293 30844 7327
rect 30878 7293 30917 7327
rect 30951 7293 31001 7327
rect 28748 7289 31001 7293
rect 28748 7255 28754 7289
rect 28788 7255 31001 7289
rect 28748 7246 31001 7255
rect 28748 7214 28866 7246
rect 28748 7180 28754 7214
rect 28788 7212 28866 7214
rect 28900 7212 31001 7246
rect 28788 7208 31001 7212
rect 28788 7180 28985 7208
rect 28748 7165 28985 7180
rect 28748 7139 28866 7165
rect 16426 7105 16891 7116
tri 16891 7105 16902 7116 sw
rect 28748 7105 28754 7139
rect 28788 7131 28866 7139
rect 28900 7131 28985 7165
rect 28788 7105 28985 7131
rect 16426 7083 16902 7105
tri 16902 7083 16924 7105 sw
rect 28748 7083 28985 7105
rect 478 6940 520 7070
rect 16426 7064 16924 7083
tri 16924 7064 16943 7083 sw
rect 28748 7064 28866 7083
rect 16426 7030 16943 7064
tri 16943 7030 16977 7064 sw
rect 28748 7030 28754 7064
rect 28788 7049 28866 7064
rect 28900 7049 28985 7083
rect 28788 7030 28985 7049
rect 16426 7001 16977 7030
tri 16977 7001 17006 7030 sw
rect 28748 7001 28985 7030
rect 16426 6989 17006 7001
tri 17006 6989 17018 7001 sw
rect 28748 6989 28866 7001
rect 16426 6955 17018 6989
tri 17018 6955 17052 6989 sw
rect 28748 6955 28754 6989
rect 28788 6967 28866 6989
rect 28900 6967 28985 7001
rect 28788 6955 28985 6967
rect 16426 6952 17052 6955
tri 17052 6952 17055 6955 sw
rect 16426 6948 17246 6952
tri 16490 6940 16498 6948 ne
rect 16498 6947 17246 6948
rect 16498 6940 17029 6947
tri 16498 6919 16519 6940 ne
rect 16519 6919 17029 6940
tri 16519 6913 16525 6919 ne
rect 16525 6913 17029 6919
tri 16525 6879 16559 6913 ne
rect 16559 6895 17029 6913
rect 17081 6895 17107 6947
rect 17159 6895 17185 6947
rect 17237 6895 17246 6947
rect 16559 6879 17246 6895
tri 16559 6837 16601 6879 ne
rect 16601 6837 17246 6879
tri 16601 6803 16635 6837 ne
rect 16635 6825 17246 6837
rect 16635 6803 17029 6825
tri 16635 6770 16668 6803 ne
rect 16668 6773 17029 6803
rect 17081 6773 17107 6825
rect 17159 6773 17185 6825
rect 17237 6773 17246 6825
rect 28748 6919 28985 6955
rect 28748 6913 28866 6919
rect 28748 6879 28754 6913
rect 28788 6885 28866 6913
rect 28900 6885 28985 6919
rect 28788 6879 28985 6885
rect 28748 6837 28985 6879
rect 28748 6803 28754 6837
rect 28788 6803 28866 6837
rect 28900 6803 28985 6837
rect 28748 6786 28985 6803
rect 16668 6770 17246 6773
tri 30167 5863 30178 5874 se
rect 30178 5863 32056 5874
rect 30094 5835 32056 5863
rect 30094 5811 30216 5835
tri 30149 5801 30159 5811 ne
rect 30159 5801 30216 5811
rect 30250 5801 30291 5835
rect 30325 5801 30366 5835
rect 30400 5801 30441 5835
rect 30475 5801 30516 5835
rect 30550 5801 30591 5835
rect 30625 5801 30666 5835
rect 30700 5801 30741 5835
rect 30775 5801 30816 5835
rect 30850 5801 30891 5835
rect 30925 5801 30966 5835
rect 31000 5801 31041 5835
rect 31075 5801 31116 5835
rect 31150 5801 31191 5835
rect 31225 5801 31266 5835
rect 31300 5801 31341 5835
rect 31375 5801 31416 5835
rect 31450 5801 31491 5835
rect 31525 5801 31566 5835
rect 31600 5801 31640 5835
rect 31674 5801 31714 5835
rect 31748 5801 31788 5835
rect 31822 5801 31862 5835
rect 31896 5801 31936 5835
rect 31970 5801 32010 5835
rect 32044 5801 32056 5835
tri 30159 5762 30198 5801 ne
rect 30198 5762 32056 5801
rect 16796 5545 18967 5552
rect 16796 5511 16808 5545
rect 16842 5511 16881 5545
rect 16915 5511 16954 5545
rect 16988 5511 17027 5545
rect 17061 5539 17100 5545
rect 17134 5539 17173 5545
rect 17207 5539 17246 5545
rect 17079 5511 17100 5539
rect 17159 5511 17173 5539
rect 17239 5511 17246 5539
rect 17280 5511 17319 5545
rect 17353 5511 17392 5545
rect 17426 5511 17465 5545
rect 17499 5511 17538 5545
rect 17572 5511 17611 5545
rect 17645 5511 17684 5545
rect 17718 5511 17757 5545
rect 17791 5511 17830 5545
rect 17864 5511 17903 5545
rect 17937 5511 17976 5545
rect 18010 5511 18049 5545
rect 18083 5511 18122 5545
rect 18156 5511 18195 5545
rect 18229 5511 18268 5545
rect 18302 5511 18341 5545
rect 18375 5511 18414 5545
rect 18448 5511 18487 5545
rect 18521 5511 18560 5545
rect 18594 5511 18633 5545
rect 18667 5511 18705 5545
rect 18739 5511 18777 5545
rect 18811 5511 18849 5545
rect 18883 5511 18921 5545
rect 18955 5511 18967 5545
rect 16796 5487 17027 5511
rect 17079 5487 17107 5511
rect 17159 5487 17187 5511
rect 17239 5487 18967 5511
rect 16796 5473 18967 5487
rect 16796 5467 17027 5473
rect 17079 5467 17107 5473
rect 17159 5467 17187 5473
rect 17239 5467 18967 5473
rect 16796 5433 16808 5467
rect 16842 5433 16881 5467
rect 16915 5433 16954 5467
rect 16988 5433 17027 5467
rect 17079 5433 17100 5467
rect 17159 5433 17173 5467
rect 17239 5433 17246 5467
rect 17280 5433 17319 5467
rect 17353 5433 17392 5467
rect 17426 5433 17465 5467
rect 17499 5433 17538 5467
rect 17572 5433 17611 5467
rect 17645 5433 17684 5467
rect 17718 5433 17757 5467
rect 17791 5433 17830 5467
rect 17864 5433 17903 5467
rect 17937 5433 17976 5467
rect 18010 5433 18049 5467
rect 18083 5433 18122 5467
rect 18156 5433 18195 5467
rect 18229 5433 18268 5467
rect 18302 5433 18341 5467
rect 18375 5433 18414 5467
rect 18448 5433 18487 5467
rect 18521 5433 18560 5467
rect 18594 5433 18633 5467
rect 18667 5433 18705 5467
rect 18739 5433 18777 5467
rect 18811 5433 18849 5467
rect 18883 5433 18921 5467
rect 18955 5433 18967 5467
rect 16796 5421 17027 5433
rect 17079 5421 17107 5433
rect 17159 5421 17187 5433
rect 17239 5421 18967 5433
rect 16796 5407 18967 5421
rect 16796 5389 17027 5407
rect 17079 5389 17107 5407
rect 17159 5389 17187 5407
rect 17239 5389 18967 5407
rect 16796 5355 16808 5389
rect 16842 5355 16881 5389
rect 16915 5355 16954 5389
rect 16988 5355 17027 5389
rect 17079 5355 17100 5389
rect 17159 5355 17173 5389
rect 17239 5355 17246 5389
rect 17280 5355 17319 5389
rect 17353 5355 17392 5389
rect 17426 5355 17465 5389
rect 17499 5355 17538 5389
rect 17572 5355 17611 5389
rect 17645 5355 17684 5389
rect 17718 5355 17757 5389
rect 17791 5355 17830 5389
rect 17864 5355 17903 5389
rect 17937 5355 17976 5389
rect 18010 5355 18049 5389
rect 18083 5355 18122 5389
rect 18156 5355 18195 5389
rect 18229 5355 18268 5389
rect 18302 5355 18341 5389
rect 18375 5355 18414 5389
rect 18448 5355 18487 5389
rect 18521 5355 18560 5389
rect 18594 5355 18633 5389
rect 18667 5355 18705 5389
rect 18739 5355 18777 5389
rect 18811 5355 18849 5389
rect 18883 5355 18921 5389
rect 18955 5355 18967 5389
rect 16796 5340 18967 5355
rect 16796 5311 17027 5340
rect 17079 5311 17107 5340
rect 17159 5311 17187 5340
rect 17239 5311 18967 5340
rect 16796 5277 16808 5311
rect 16842 5277 16881 5311
rect 16915 5277 16954 5311
rect 16988 5277 17027 5311
rect 17079 5288 17100 5311
rect 17159 5288 17173 5311
rect 17239 5288 17246 5311
rect 17061 5277 17100 5288
rect 17134 5277 17173 5288
rect 17207 5277 17246 5288
rect 17280 5277 17319 5311
rect 17353 5277 17392 5311
rect 17426 5277 17465 5311
rect 17499 5277 17538 5311
rect 17572 5277 17611 5311
rect 17645 5277 17684 5311
rect 17718 5277 17757 5311
rect 17791 5277 17830 5311
rect 17864 5277 17903 5311
rect 17937 5277 17976 5311
rect 18010 5277 18049 5311
rect 18083 5277 18122 5311
rect 18156 5277 18195 5311
rect 18229 5277 18268 5311
rect 18302 5277 18341 5311
rect 18375 5277 18414 5311
rect 18448 5277 18487 5311
rect 18521 5277 18560 5311
rect 18594 5277 18633 5311
rect 18667 5277 18705 5311
rect 18739 5277 18777 5311
rect 18811 5277 18849 5311
rect 18883 5277 18921 5311
rect 18955 5277 18967 5311
rect 16796 5270 18967 5277
rect 27866 5141 28690 5147
rect 27866 5135 28174 5141
rect 28226 5135 28262 5141
rect 28314 5135 28350 5141
rect 28402 5135 28690 5141
rect 27866 5101 27910 5135
rect 27944 5101 27988 5135
rect 28022 5101 28066 5135
rect 28100 5101 28144 5135
rect 28256 5101 28262 5135
rect 28334 5101 28350 5135
rect 28412 5101 28456 5135
rect 28490 5101 28534 5135
rect 28568 5101 28612 5135
rect 28646 5101 28690 5135
rect 27866 5089 28174 5101
rect 28226 5089 28262 5101
rect 28314 5089 28350 5101
rect 28402 5089 28690 5101
rect 27866 5063 28690 5089
rect 27866 5058 28174 5063
rect 28226 5058 28262 5063
rect 28314 5058 28350 5063
rect 28402 5058 28690 5063
rect 27866 5024 27910 5058
rect 27944 5024 27988 5058
rect 28022 5024 28066 5058
rect 28100 5024 28144 5058
rect 28256 5024 28262 5058
rect 28334 5024 28350 5058
rect 28412 5024 28456 5058
rect 28490 5024 28534 5058
rect 28568 5024 28612 5058
rect 28646 5024 28690 5058
rect 27866 5011 28174 5024
rect 28226 5011 28262 5024
rect 28314 5011 28350 5024
rect 28402 5011 28690 5024
rect 27866 4984 28690 5011
rect 27866 4980 28174 4984
rect 28226 4980 28262 4984
rect 28314 4980 28350 4984
rect 28402 4980 28690 4984
rect 27866 4946 27910 4980
rect 27944 4946 27988 4980
rect 28022 4946 28066 4980
rect 28100 4946 28144 4980
rect 28256 4946 28262 4980
rect 28334 4946 28350 4980
rect 28412 4946 28456 4980
rect 28490 4946 28534 4980
rect 28568 4946 28612 4980
rect 28646 4946 28690 4980
rect 27866 4932 28174 4946
rect 28226 4932 28262 4946
rect 28314 4932 28350 4946
rect 28402 4932 28690 4946
rect 27866 4905 28690 4932
rect 27866 4902 28174 4905
rect 28226 4902 28262 4905
rect 28314 4902 28350 4905
rect 28402 4902 28690 4905
rect 27866 4868 27910 4902
rect 27944 4868 27988 4902
rect 28022 4868 28066 4902
rect 28100 4868 28144 4902
rect 28256 4868 28262 4902
rect 28334 4868 28350 4902
rect 28412 4868 28456 4902
rect 28490 4868 28534 4902
rect 28568 4868 28612 4902
rect 28646 4868 28690 4902
rect 27866 4853 28174 4868
rect 28226 4853 28262 4868
rect 28314 4853 28350 4868
rect 28402 4853 28690 4868
rect 27866 4824 28690 4853
rect 27866 4790 27910 4824
rect 27944 4790 27988 4824
rect 28022 4790 28066 4824
rect 28100 4790 28144 4824
rect 28178 4790 28222 4824
rect 28256 4790 28300 4824
rect 28334 4790 28378 4824
rect 28412 4790 28456 4824
rect 28490 4790 28534 4824
rect 28568 4790 28612 4824
rect 28646 4790 28690 4824
tri 27838 4746 27866 4774 se
rect 27866 4766 28690 4790
rect 27866 4746 27980 4766
rect 28032 4746 28068 4766
rect 28120 4746 28156 4766
rect 28208 4746 28690 4766
tri 27804 4712 27838 4746 se
rect 27838 4712 27910 4746
rect 27944 4714 27980 4746
rect 28032 4714 28066 4746
rect 28120 4714 28144 4746
rect 28208 4714 28222 4746
rect 27944 4712 27988 4714
rect 28022 4712 28066 4714
rect 28100 4712 28144 4714
rect 28178 4712 28222 4714
rect 28256 4712 28300 4746
rect 28334 4712 28378 4746
rect 28412 4712 28456 4746
rect 28490 4712 28534 4746
rect 28568 4712 28612 4746
rect 28646 4712 28690 4746
tri 27760 4668 27804 4712 se
rect 27804 4700 28690 4712
rect 27804 4668 27980 4700
rect 28032 4668 28068 4700
rect 28120 4668 28156 4700
rect 28208 4668 28690 4700
tri 27726 4634 27760 4668 se
rect 27760 4634 27910 4668
rect 27944 4648 27980 4668
rect 28032 4648 28066 4668
rect 28120 4648 28144 4668
rect 28208 4648 28222 4668
rect 27944 4634 27988 4648
rect 28022 4634 28066 4648
rect 28100 4634 28144 4648
rect 28178 4634 28222 4648
rect 28256 4634 28300 4668
rect 28334 4634 28378 4668
rect 28412 4634 28456 4668
rect 28490 4634 28534 4668
rect 28568 4634 28612 4668
rect 28646 4634 28690 4668
tri 27716 4624 27726 4634 se
rect 27726 4624 27980 4634
rect 26701 4615 27980 4624
rect 26701 4581 26713 4615
rect 26747 4581 26788 4615
rect 26822 4581 26863 4615
rect 26897 4608 26938 4615
rect 26972 4608 27013 4615
rect 27047 4608 27088 4615
rect 27122 4608 27163 4615
rect 27197 4608 27238 4615
rect 27272 4608 27312 4615
rect 26922 4581 26938 4608
rect 27005 4581 27013 4608
rect 27087 4581 27088 4608
rect 27197 4581 27199 4608
rect 27272 4581 27281 4608
rect 27346 4581 27386 4615
rect 27420 4581 27460 4615
rect 27494 4581 27534 4615
rect 27568 4581 27608 4615
rect 27642 4581 27682 4615
rect 27716 4581 27756 4615
rect 27790 4590 27980 4615
rect 28032 4590 28068 4634
rect 28120 4590 28156 4634
rect 28208 4590 28690 4634
rect 27790 4581 27910 4590
rect 26701 4556 26870 4581
rect 26922 4556 26953 4581
rect 27005 4556 27035 4581
rect 27087 4556 27117 4581
rect 27169 4556 27199 4581
rect 27251 4556 27281 4581
rect 27333 4556 27910 4581
rect 27944 4582 27980 4590
rect 28032 4582 28066 4590
rect 28120 4582 28144 4590
rect 28208 4582 28222 4590
rect 27944 4568 27988 4582
rect 28022 4568 28066 4582
rect 28100 4568 28144 4582
rect 28178 4568 28222 4582
rect 27944 4556 27980 4568
rect 28032 4556 28066 4568
rect 28120 4556 28144 4568
rect 28208 4556 28222 4568
rect 28256 4556 28300 4590
rect 28334 4556 28378 4590
rect 28412 4556 28456 4590
rect 28490 4556 28534 4590
rect 28568 4556 28612 4590
rect 28646 4556 28690 4590
rect 26701 4535 27980 4556
rect 26701 4501 26713 4535
rect 26747 4501 26788 4535
rect 26822 4501 26863 4535
rect 26897 4512 26938 4535
rect 26972 4512 27013 4535
rect 27047 4512 27088 4535
rect 27122 4512 27163 4535
rect 27197 4512 27238 4535
rect 27272 4512 27312 4535
rect 26922 4501 26938 4512
rect 27005 4501 27013 4512
rect 27087 4501 27088 4512
rect 27197 4501 27199 4512
rect 27272 4501 27281 4512
rect 27346 4501 27386 4535
rect 27420 4501 27460 4535
rect 27494 4501 27534 4535
rect 27568 4501 27608 4535
rect 27642 4501 27682 4535
rect 27716 4501 27756 4535
rect 27790 4516 27980 4535
rect 28032 4516 28068 4556
rect 28120 4516 28156 4556
rect 28208 4516 28690 4556
rect 27790 4512 28690 4516
rect 27790 4501 27910 4512
rect 26701 4460 26870 4501
rect 26922 4460 26953 4501
rect 27005 4460 27035 4501
rect 27087 4460 27117 4501
rect 27169 4460 27199 4501
rect 27251 4460 27281 4501
rect 27333 4478 27910 4501
rect 27944 4502 27988 4512
rect 28022 4502 28066 4512
rect 28100 4502 28144 4512
rect 28178 4502 28222 4512
rect 27944 4478 27980 4502
rect 28032 4478 28066 4502
rect 28120 4478 28144 4502
rect 28208 4478 28222 4502
rect 28256 4478 28300 4512
rect 28334 4478 28378 4512
rect 28412 4478 28456 4512
rect 28490 4478 28534 4512
rect 28568 4478 28612 4512
rect 28646 4478 28690 4512
rect 27333 4460 27980 4478
rect 26701 4455 27980 4460
rect 26701 4421 26713 4455
rect 26747 4421 26788 4455
rect 26822 4421 26863 4455
rect 26897 4421 26938 4455
rect 26972 4421 27013 4455
rect 27047 4421 27088 4455
rect 27122 4421 27163 4455
rect 27197 4421 27238 4455
rect 27272 4421 27312 4455
rect 27346 4421 27386 4455
rect 27420 4421 27460 4455
rect 27494 4421 27534 4455
rect 27568 4421 27608 4455
rect 27642 4421 27682 4455
rect 27716 4421 27756 4455
rect 27790 4450 27980 4455
rect 28032 4450 28068 4478
rect 28120 4450 28156 4478
rect 28208 4450 28690 4478
rect 27790 4436 28690 4450
rect 27790 4434 27980 4436
rect 28032 4434 28068 4436
rect 28120 4434 28156 4436
rect 28208 4434 28690 4436
rect 27790 4421 27910 4434
rect 26701 4416 27910 4421
rect 26701 4375 26870 4416
rect 26922 4375 26953 4416
rect 27005 4375 27035 4416
rect 27087 4375 27117 4416
rect 27169 4375 27199 4416
rect 27251 4375 27281 4416
rect 27333 4400 27910 4416
rect 27944 4400 27980 4434
rect 28032 4400 28066 4434
rect 28120 4400 28144 4434
rect 28208 4400 28222 4434
rect 28256 4400 28300 4434
rect 28334 4400 28378 4434
rect 28412 4400 28456 4434
rect 28490 4400 28534 4434
rect 28568 4400 28612 4434
rect 28646 4400 28690 4434
rect 27333 4384 27980 4400
rect 28032 4384 28068 4400
rect 28120 4384 28156 4400
rect 28208 4384 28690 4400
rect 27333 4375 28690 4384
rect 26701 4341 26713 4375
rect 26747 4341 26788 4375
rect 26822 4341 26863 4375
rect 26922 4364 26938 4375
rect 27005 4364 27013 4375
rect 27087 4364 27088 4375
rect 27197 4364 27199 4375
rect 27272 4364 27281 4375
rect 26897 4341 26938 4364
rect 26972 4341 27013 4364
rect 27047 4341 27088 4364
rect 27122 4341 27163 4364
rect 27197 4341 27238 4364
rect 27272 4341 27312 4364
rect 27346 4341 27386 4375
rect 27420 4341 27460 4375
rect 27494 4341 27534 4375
rect 27568 4341 27608 4375
rect 27642 4341 27682 4375
rect 27716 4341 27756 4375
rect 27790 4369 28690 4375
rect 27790 4356 27980 4369
rect 28032 4356 28068 4369
rect 28120 4356 28156 4369
rect 28208 4356 28690 4369
rect 27790 4341 27910 4356
rect 26701 4322 27910 4341
rect 27944 4322 27980 4356
rect 28032 4322 28066 4356
rect 28120 4322 28144 4356
rect 28208 4322 28222 4356
rect 28256 4322 28300 4356
rect 28334 4322 28378 4356
rect 28412 4322 28456 4356
rect 28490 4322 28534 4356
rect 28568 4322 28612 4356
rect 28646 4322 28690 4356
rect 26701 4320 27980 4322
rect 26701 4295 26870 4320
rect 26922 4295 26953 4320
rect 27005 4295 27035 4320
rect 27087 4295 27117 4320
rect 27169 4295 27199 4320
rect 27251 4295 27281 4320
rect 27333 4317 27980 4320
rect 28032 4317 28068 4322
rect 28120 4317 28156 4322
rect 28208 4317 28690 4322
rect 27333 4302 28690 4317
rect 27333 4295 27980 4302
rect 26701 4261 26713 4295
rect 26747 4261 26788 4295
rect 26822 4261 26863 4295
rect 26922 4268 26938 4295
rect 27005 4268 27013 4295
rect 27087 4268 27088 4295
rect 27197 4268 27199 4295
rect 27272 4268 27281 4295
rect 26897 4261 26938 4268
rect 26972 4261 27013 4268
rect 27047 4261 27088 4268
rect 27122 4261 27163 4268
rect 27197 4261 27238 4268
rect 27272 4261 27312 4268
rect 27346 4261 27386 4295
rect 27420 4261 27460 4295
rect 27494 4261 27534 4295
rect 27568 4261 27608 4295
rect 27642 4261 27682 4295
rect 27716 4261 27756 4295
rect 27790 4278 27980 4295
rect 28032 4278 28068 4302
rect 28120 4278 28156 4302
rect 28208 4278 28690 4302
rect 27790 4261 27910 4278
rect 26701 4244 27910 4261
rect 27944 4250 27980 4278
rect 28032 4250 28066 4278
rect 28120 4250 28144 4278
rect 28208 4250 28222 4278
rect 27944 4244 27988 4250
rect 28022 4244 28066 4250
rect 28100 4244 28144 4250
rect 28178 4244 28222 4250
rect 28256 4244 28300 4278
rect 28334 4244 28378 4278
rect 28412 4244 28456 4278
rect 28490 4244 28534 4278
rect 28568 4244 28612 4278
rect 28646 4244 28690 4278
rect 26701 4235 28690 4244
rect 26701 4224 27980 4235
rect 26701 4215 26870 4224
rect 26922 4215 26953 4224
rect 27005 4215 27035 4224
rect 27087 4215 27117 4224
rect 27169 4215 27199 4224
rect 27251 4215 27281 4224
rect 27333 4215 27980 4224
rect 26701 4181 26713 4215
rect 26747 4181 26788 4215
rect 26822 4181 26863 4215
rect 26922 4181 26938 4215
rect 27005 4181 27013 4215
rect 27087 4181 27088 4215
rect 27197 4181 27199 4215
rect 27272 4181 27281 4215
rect 27346 4181 27386 4215
rect 27420 4181 27460 4215
rect 27494 4181 27534 4215
rect 27568 4181 27608 4215
rect 27642 4181 27682 4215
rect 27716 4181 27756 4215
rect 27790 4200 27980 4215
rect 28032 4200 28068 4235
rect 28120 4200 28156 4235
rect 28208 4200 28690 4235
rect 27790 4181 27910 4200
rect 26701 4172 26870 4181
rect 26922 4172 26953 4181
rect 27005 4172 27035 4181
rect 27087 4172 27117 4181
rect 27169 4172 27199 4181
rect 27251 4172 27281 4181
rect 27333 4172 27910 4181
rect 26701 4166 27910 4172
rect 27944 4183 27980 4200
rect 28032 4183 28066 4200
rect 28120 4183 28144 4200
rect 28208 4183 28222 4200
rect 27944 4166 27988 4183
rect 28022 4166 28066 4183
rect 28100 4166 28144 4183
rect 28178 4166 28222 4183
rect 28256 4166 28300 4200
rect 28334 4166 28378 4200
rect 28412 4166 28456 4200
rect 28490 4166 28534 4200
rect 28568 4166 28612 4200
rect 28646 4166 28690 4200
rect 26701 4154 28690 4166
rect 6715 3347 6755 3549
rect 16507 3347 16518 3549
rect 6715 3189 6755 3319
rect 9103 3307 9149 3319
rect 9103 3273 9109 3307
rect 9143 3273 9149 3307
rect 9103 3235 9149 3273
rect 9103 3201 9109 3235
rect 9143 3201 9149 3235
rect 9103 3189 9149 3201
rect 9275 3307 9321 3319
rect 9275 3273 9281 3307
rect 9315 3273 9321 3307
rect 9275 3235 9321 3273
rect 9275 3201 9281 3235
rect 9315 3201 9321 3235
rect 9275 3189 9321 3201
rect 10763 3307 10809 3319
rect 10763 3273 10769 3307
rect 10803 3273 10809 3307
rect 10763 3235 10809 3273
rect 10763 3201 10769 3235
rect 10803 3201 10809 3235
rect 10763 3189 10809 3201
rect 10935 3307 10981 3319
rect 10935 3273 10941 3307
rect 10975 3273 10981 3307
rect 10935 3235 10981 3273
rect 10935 3201 10941 3235
rect 10975 3201 10981 3235
rect 10935 3189 10981 3201
rect 16501 3189 16518 3319
rect 16508 2959 16518 3161
rect 4549 2556 4583 2590
rect 22399 2462 22649 2474
rect 22399 2428 22405 2462
rect 22439 2428 22507 2462
rect 22541 2428 22609 2462
rect 22643 2428 22649 2462
rect 6715 2198 6755 2400
rect 16505 2198 16519 2400
rect 22399 2387 22649 2428
rect 22399 2353 22405 2387
rect 22439 2353 22507 2387
rect 22541 2353 22609 2387
rect 22643 2353 22649 2387
rect 22399 2312 22649 2353
rect 22399 2278 22405 2312
rect 22439 2278 22507 2312
rect 22541 2278 22609 2312
rect 22643 2278 22649 2312
rect 22399 2237 22649 2278
rect 22399 2203 22405 2237
rect 22439 2203 22507 2237
rect 22541 2203 22609 2237
rect 22643 2203 22649 2237
rect 22399 2170 22649 2203
rect 2121 2130 2170 2163
rect 22306 2162 22649 2170
rect 22306 2128 22405 2162
rect 22439 2128 22507 2162
rect 22541 2128 22609 2162
rect 22643 2128 22649 2162
rect 22306 2087 22649 2128
rect 22306 2053 22405 2087
rect 22439 2053 22507 2087
rect 22541 2053 22609 2087
rect 22643 2053 22649 2087
rect 22306 2052 22649 2053
tri 22323 2012 22363 2052 ne
rect 22363 2012 22649 2052
tri 22363 2007 22368 2012 ne
rect 22368 1978 22405 2012
rect 22439 1978 22507 2012
rect 22541 1978 22609 2012
rect 22643 1978 22649 2012
rect 22368 1936 22649 1978
rect 22368 1902 22405 1936
rect 22439 1902 22507 1936
rect 22541 1902 22609 1936
rect 22643 1902 22649 1936
rect 22368 1860 22649 1902
rect 22368 1826 22405 1860
rect 22439 1826 22507 1860
rect 22541 1826 22609 1860
rect 22643 1826 22649 1860
rect 22368 1784 22649 1826
rect 22368 1750 22405 1784
rect 22439 1750 22507 1784
rect 22541 1750 22609 1784
rect 22643 1750 22649 1784
rect 15566 1743 15886 1749
rect 15566 1691 15572 1743
rect 15624 1691 15636 1743
rect 15688 1691 15700 1743
rect 15752 1691 15764 1743
rect 15816 1691 15828 1743
rect 15880 1691 15886 1743
rect 22368 1738 22649 1750
rect 15566 1675 15886 1691
rect 15566 1623 15572 1675
rect 15624 1623 15636 1675
rect 15688 1623 15700 1675
rect 15752 1623 15764 1675
rect 15816 1623 15828 1675
rect 15880 1623 15886 1675
rect 15566 1606 15886 1623
rect 15566 1554 15572 1606
rect 15624 1554 15636 1606
rect 15688 1554 15700 1606
rect 15752 1554 15764 1606
rect 15816 1554 15828 1606
rect 15880 1554 15886 1606
rect 15566 1537 15886 1554
rect 15566 1485 15572 1537
rect 15624 1485 15636 1537
rect 15688 1485 15700 1537
rect 15752 1485 15764 1537
rect 15816 1485 15828 1537
rect 15880 1485 15886 1537
rect 15566 1468 15886 1485
rect 15566 1416 15572 1468
rect 15624 1416 15636 1468
rect 15688 1416 15700 1468
rect 15752 1416 15764 1468
rect 15816 1416 15828 1468
rect 15880 1416 15886 1468
rect 15566 1410 15886 1416
rect 2714 1372 2766 1378
rect 9434 1339 9467 1372
rect 10606 1339 10640 1373
rect 2714 1308 2766 1320
rect 2766 1256 7896 1291
rect 2714 1251 7896 1256
rect 2714 1250 2766 1251
rect 5450 1175 5487 1209
rect 16623 731 16663 933
tri 23475 411 23481 417 se
rect 23481 411 23487 417
tri 19785 345 19851 411 se
rect 19851 365 23487 411
rect 23539 365 23551 417
rect 23603 365 23609 417
tri 19851 345 19871 365 nw
tri 19719 279 19785 345 se
tri 19785 279 19851 345 nw
tri 19653 213 19719 279 se
tri 19719 213 19785 279 nw
tri 19634 194 19653 213 se
rect 19653 194 19654 213
tri 15900 128 15966 194 se
rect 15966 148 19654 194
tri 19654 148 19719 213 nw
tri 15966 128 15986 148 nw
tri 15834 62 15900 128 se
tri 15900 62 15966 128 nw
tri 15768 -4 15834 62 se
tri 15834 -4 15900 62 nw
tri 15702 -70 15768 -4 se
tri 15768 -70 15834 -4 nw
tri 15636 -136 15702 -70 se
tri 15702 -136 15768 -70 nw
tri 15579 -193 15636 -136 se
rect 15636 -193 15645 -136
tri 15645 -193 15702 -136 nw
tri 15513 -454 15579 -388 se
rect 15579 -408 15625 -193
tri 15625 -213 15645 -193 nw
tri 15579 -454 15625 -408 nw
tri 15501 -466 15513 -454 se
rect 13175 -512 13386 -466
tri 13342 -556 13386 -512 ne
tri 13386 -540 13460 -466 sw
tri 15447 -520 15501 -466 se
rect 15501 -520 15513 -466
tri 15513 -520 15579 -454 nw
tri 15427 -540 15447 -520 se
rect 13386 -546 15447 -540
rect 13386 -556 13682 -546
tri 13386 -604 13434 -556 ne
rect 13434 -598 13682 -556
rect 13734 -598 13746 -546
rect 13798 -586 15447 -546
tri 15447 -586 15513 -520 nw
rect 13434 -604 13798 -598
tri 13798 -604 13816 -586 nw
rect 13682 -1165 13798 -1159
tri 10954 -1237 11004 -1187 se
rect 11004 -1217 13682 -1187
rect 13734 -1217 13746 -1165
rect 11004 -1223 13798 -1217
tri 11004 -1237 11018 -1223 nw
tri 10904 -1287 10954 -1237 se
tri 10954 -1287 11004 -1237 nw
tri 10854 -1337 10904 -1287 se
tri 10904 -1337 10954 -1287 nw
tri 10805 -1386 10854 -1337 se
rect 10854 -1386 10855 -1337
tri 10855 -1386 10904 -1337 nw
rect 10638 -1422 10819 -1386
tri 10819 -1422 10855 -1386 nw
<< via1 >>
rect 17029 6895 17081 6947
rect 17107 6895 17159 6947
rect 17185 6895 17237 6947
rect 17029 6773 17081 6825
rect 17107 6773 17159 6825
rect 17185 6773 17237 6825
rect 17027 5511 17061 5539
rect 17061 5511 17079 5539
rect 17107 5511 17134 5539
rect 17134 5511 17159 5539
rect 17187 5511 17207 5539
rect 17207 5511 17239 5539
rect 17027 5487 17079 5511
rect 17107 5487 17159 5511
rect 17187 5487 17239 5511
rect 17027 5467 17079 5473
rect 17107 5467 17159 5473
rect 17187 5467 17239 5473
rect 17027 5433 17061 5467
rect 17061 5433 17079 5467
rect 17107 5433 17134 5467
rect 17134 5433 17159 5467
rect 17187 5433 17207 5467
rect 17207 5433 17239 5467
rect 17027 5421 17079 5433
rect 17107 5421 17159 5433
rect 17187 5421 17239 5433
rect 17027 5389 17079 5407
rect 17107 5389 17159 5407
rect 17187 5389 17239 5407
rect 17027 5355 17061 5389
rect 17061 5355 17079 5389
rect 17107 5355 17134 5389
rect 17134 5355 17159 5389
rect 17187 5355 17207 5389
rect 17207 5355 17239 5389
rect 17027 5311 17079 5340
rect 17107 5311 17159 5340
rect 17187 5311 17239 5340
rect 17027 5288 17061 5311
rect 17061 5288 17079 5311
rect 17107 5288 17134 5311
rect 17134 5288 17159 5311
rect 17187 5288 17207 5311
rect 17207 5288 17239 5311
rect 28174 5135 28226 5141
rect 28262 5135 28314 5141
rect 28350 5135 28402 5141
rect 28174 5101 28178 5135
rect 28178 5101 28222 5135
rect 28222 5101 28226 5135
rect 28262 5101 28300 5135
rect 28300 5101 28314 5135
rect 28350 5101 28378 5135
rect 28378 5101 28402 5135
rect 28174 5089 28226 5101
rect 28262 5089 28314 5101
rect 28350 5089 28402 5101
rect 28174 5058 28226 5063
rect 28262 5058 28314 5063
rect 28350 5058 28402 5063
rect 28174 5024 28178 5058
rect 28178 5024 28222 5058
rect 28222 5024 28226 5058
rect 28262 5024 28300 5058
rect 28300 5024 28314 5058
rect 28350 5024 28378 5058
rect 28378 5024 28402 5058
rect 28174 5011 28226 5024
rect 28262 5011 28314 5024
rect 28350 5011 28402 5024
rect 28174 4980 28226 4984
rect 28262 4980 28314 4984
rect 28350 4980 28402 4984
rect 28174 4946 28178 4980
rect 28178 4946 28222 4980
rect 28222 4946 28226 4980
rect 28262 4946 28300 4980
rect 28300 4946 28314 4980
rect 28350 4946 28378 4980
rect 28378 4946 28402 4980
rect 28174 4932 28226 4946
rect 28262 4932 28314 4946
rect 28350 4932 28402 4946
rect 28174 4902 28226 4905
rect 28262 4902 28314 4905
rect 28350 4902 28402 4905
rect 28174 4868 28178 4902
rect 28178 4868 28222 4902
rect 28222 4868 28226 4902
rect 28262 4868 28300 4902
rect 28300 4868 28314 4902
rect 28350 4868 28378 4902
rect 28378 4868 28402 4902
rect 28174 4853 28226 4868
rect 28262 4853 28314 4868
rect 28350 4853 28402 4868
rect 27980 4746 28032 4766
rect 28068 4746 28120 4766
rect 28156 4746 28208 4766
rect 27980 4714 27988 4746
rect 27988 4714 28022 4746
rect 28022 4714 28032 4746
rect 28068 4714 28100 4746
rect 28100 4714 28120 4746
rect 28156 4714 28178 4746
rect 28178 4714 28208 4746
rect 27980 4668 28032 4700
rect 28068 4668 28120 4700
rect 28156 4668 28208 4700
rect 27980 4648 27988 4668
rect 27988 4648 28022 4668
rect 28022 4648 28032 4668
rect 28068 4648 28100 4668
rect 28100 4648 28120 4668
rect 28156 4648 28178 4668
rect 28178 4648 28208 4668
rect 26870 4581 26897 4608
rect 26897 4581 26922 4608
rect 26953 4581 26972 4608
rect 26972 4581 27005 4608
rect 27035 4581 27047 4608
rect 27047 4581 27087 4608
rect 27117 4581 27122 4608
rect 27122 4581 27163 4608
rect 27163 4581 27169 4608
rect 27199 4581 27238 4608
rect 27238 4581 27251 4608
rect 27281 4581 27312 4608
rect 27312 4581 27333 4608
rect 27980 4590 28032 4634
rect 28068 4590 28120 4634
rect 28156 4590 28208 4634
rect 26870 4556 26922 4581
rect 26953 4556 27005 4581
rect 27035 4556 27087 4581
rect 27117 4556 27169 4581
rect 27199 4556 27251 4581
rect 27281 4556 27333 4581
rect 27980 4582 27988 4590
rect 27988 4582 28022 4590
rect 28022 4582 28032 4590
rect 28068 4582 28100 4590
rect 28100 4582 28120 4590
rect 28156 4582 28178 4590
rect 28178 4582 28208 4590
rect 27980 4556 27988 4568
rect 27988 4556 28022 4568
rect 28022 4556 28032 4568
rect 28068 4556 28100 4568
rect 28100 4556 28120 4568
rect 28156 4556 28178 4568
rect 28178 4556 28208 4568
rect 26870 4501 26897 4512
rect 26897 4501 26922 4512
rect 26953 4501 26972 4512
rect 26972 4501 27005 4512
rect 27035 4501 27047 4512
rect 27047 4501 27087 4512
rect 27117 4501 27122 4512
rect 27122 4501 27163 4512
rect 27163 4501 27169 4512
rect 27199 4501 27238 4512
rect 27238 4501 27251 4512
rect 27281 4501 27312 4512
rect 27312 4501 27333 4512
rect 27980 4516 28032 4556
rect 28068 4516 28120 4556
rect 28156 4516 28208 4556
rect 26870 4460 26922 4501
rect 26953 4460 27005 4501
rect 27035 4460 27087 4501
rect 27117 4460 27169 4501
rect 27199 4460 27251 4501
rect 27281 4460 27333 4501
rect 27980 4478 27988 4502
rect 27988 4478 28022 4502
rect 28022 4478 28032 4502
rect 28068 4478 28100 4502
rect 28100 4478 28120 4502
rect 28156 4478 28178 4502
rect 28178 4478 28208 4502
rect 27980 4450 28032 4478
rect 28068 4450 28120 4478
rect 28156 4450 28208 4478
rect 27980 4434 28032 4436
rect 28068 4434 28120 4436
rect 28156 4434 28208 4436
rect 26870 4375 26922 4416
rect 26953 4375 27005 4416
rect 27035 4375 27087 4416
rect 27117 4375 27169 4416
rect 27199 4375 27251 4416
rect 27281 4375 27333 4416
rect 27980 4400 27988 4434
rect 27988 4400 28022 4434
rect 28022 4400 28032 4434
rect 28068 4400 28100 4434
rect 28100 4400 28120 4434
rect 28156 4400 28178 4434
rect 28178 4400 28208 4434
rect 27980 4384 28032 4400
rect 28068 4384 28120 4400
rect 28156 4384 28208 4400
rect 26870 4364 26897 4375
rect 26897 4364 26922 4375
rect 26953 4364 26972 4375
rect 26972 4364 27005 4375
rect 27035 4364 27047 4375
rect 27047 4364 27087 4375
rect 27117 4364 27122 4375
rect 27122 4364 27163 4375
rect 27163 4364 27169 4375
rect 27199 4364 27238 4375
rect 27238 4364 27251 4375
rect 27281 4364 27312 4375
rect 27312 4364 27333 4375
rect 27980 4356 28032 4369
rect 28068 4356 28120 4369
rect 28156 4356 28208 4369
rect 27980 4322 27988 4356
rect 27988 4322 28022 4356
rect 28022 4322 28032 4356
rect 28068 4322 28100 4356
rect 28100 4322 28120 4356
rect 28156 4322 28178 4356
rect 28178 4322 28208 4356
rect 26870 4295 26922 4320
rect 26953 4295 27005 4320
rect 27035 4295 27087 4320
rect 27117 4295 27169 4320
rect 27199 4295 27251 4320
rect 27281 4295 27333 4320
rect 27980 4317 28032 4322
rect 28068 4317 28120 4322
rect 28156 4317 28208 4322
rect 26870 4268 26897 4295
rect 26897 4268 26922 4295
rect 26953 4268 26972 4295
rect 26972 4268 27005 4295
rect 27035 4268 27047 4295
rect 27047 4268 27087 4295
rect 27117 4268 27122 4295
rect 27122 4268 27163 4295
rect 27163 4268 27169 4295
rect 27199 4268 27238 4295
rect 27238 4268 27251 4295
rect 27281 4268 27312 4295
rect 27312 4268 27333 4295
rect 27980 4278 28032 4302
rect 28068 4278 28120 4302
rect 28156 4278 28208 4302
rect 27980 4250 27988 4278
rect 27988 4250 28022 4278
rect 28022 4250 28032 4278
rect 28068 4250 28100 4278
rect 28100 4250 28120 4278
rect 28156 4250 28178 4278
rect 28178 4250 28208 4278
rect 26870 4215 26922 4224
rect 26953 4215 27005 4224
rect 27035 4215 27087 4224
rect 27117 4215 27169 4224
rect 27199 4215 27251 4224
rect 27281 4215 27333 4224
rect 26870 4181 26897 4215
rect 26897 4181 26922 4215
rect 26953 4181 26972 4215
rect 26972 4181 27005 4215
rect 27035 4181 27047 4215
rect 27047 4181 27087 4215
rect 27117 4181 27122 4215
rect 27122 4181 27163 4215
rect 27163 4181 27169 4215
rect 27199 4181 27238 4215
rect 27238 4181 27251 4215
rect 27281 4181 27312 4215
rect 27312 4181 27333 4215
rect 27980 4200 28032 4235
rect 28068 4200 28120 4235
rect 28156 4200 28208 4235
rect 26870 4172 26922 4181
rect 26953 4172 27005 4181
rect 27035 4172 27087 4181
rect 27117 4172 27169 4181
rect 27199 4172 27251 4181
rect 27281 4172 27333 4181
rect 27980 4183 27988 4200
rect 27988 4183 28022 4200
rect 28022 4183 28032 4200
rect 28068 4183 28100 4200
rect 28100 4183 28120 4200
rect 28156 4183 28178 4200
rect 28178 4183 28208 4200
rect 15572 1691 15624 1743
rect 15636 1691 15688 1743
rect 15700 1691 15752 1743
rect 15764 1691 15816 1743
rect 15828 1691 15880 1743
rect 15572 1623 15624 1675
rect 15636 1623 15688 1675
rect 15700 1623 15752 1675
rect 15764 1623 15816 1675
rect 15828 1623 15880 1675
rect 15572 1554 15624 1606
rect 15636 1554 15688 1606
rect 15700 1554 15752 1606
rect 15764 1554 15816 1606
rect 15828 1554 15880 1606
rect 15572 1485 15624 1537
rect 15636 1485 15688 1537
rect 15700 1485 15752 1537
rect 15764 1485 15816 1537
rect 15828 1485 15880 1537
rect 15572 1416 15624 1468
rect 15636 1416 15688 1468
rect 15700 1416 15752 1468
rect 15764 1416 15816 1468
rect 15828 1416 15880 1468
rect 2714 1320 2766 1372
rect 2714 1256 2766 1308
rect 23487 365 23539 417
rect 23551 365 23603 417
rect 13682 -598 13734 -546
rect 13746 -598 13798 -546
rect 13682 -1217 13734 -1165
rect 13746 -1217 13798 -1165
<< metal2 >>
rect 20600 23528 20822 23602
rect 31606 23371 31750 23506
rect 31830 23366 31958 23506
rect 32016 23366 32144 23506
rect 2967 13103 3235 13137
rect 17102 13103 17160 13161
rect 17328 13103 17648 13168
rect 17016 6947 17246 6952
rect 17016 6895 17029 6947
rect 17081 6895 17107 6947
rect 17159 6895 17185 6947
rect 17237 6895 17246 6947
rect 17016 6825 17246 6895
rect 17016 6773 17029 6825
rect 17081 6773 17107 6825
rect 17159 6773 17185 6825
rect 17237 6773 17246 6825
rect 17016 5539 17246 6773
rect 17016 5487 17027 5539
rect 17079 5487 17107 5539
rect 17159 5487 17187 5539
rect 17239 5487 17246 5539
rect 17016 5473 17246 5487
rect 17016 5421 17027 5473
rect 17079 5421 17107 5473
rect 17159 5421 17187 5473
rect 17239 5421 17246 5473
rect 17016 5407 17246 5421
rect 17016 5355 17027 5407
rect 17079 5355 17107 5407
rect 17159 5355 17187 5407
rect 17239 5355 17246 5407
rect 17016 5340 17246 5355
rect 17016 5288 17027 5340
rect 17079 5288 17107 5340
rect 17159 5288 17187 5340
rect 17239 5288 17246 5340
rect 17016 5277 17246 5288
rect 28173 5141 28403 5147
rect 28173 5089 28174 5141
rect 28226 5089 28262 5141
rect 28314 5089 28350 5141
rect 28402 5089 28403 5141
rect 28173 5063 28403 5089
rect 28173 5011 28174 5063
rect 28226 5011 28262 5063
rect 28314 5011 28350 5063
rect 28402 5011 28403 5063
rect 28173 4984 28403 5011
rect 28173 4932 28174 4984
rect 28226 4932 28262 4984
rect 28314 4932 28350 4984
rect 28402 4932 28403 4984
rect 28173 4905 28403 4932
rect 28173 4853 28174 4905
rect 28226 4853 28262 4905
rect 28314 4853 28350 4905
rect 28402 4853 28403 4905
rect 28173 4847 28403 4853
rect 27979 4766 28209 4772
rect 27979 4714 27980 4766
rect 28032 4714 28068 4766
rect 28120 4714 28156 4766
rect 28208 4714 28209 4766
rect 27979 4700 28209 4714
rect 27979 4648 27980 4700
rect 28032 4648 28068 4700
rect 28120 4648 28156 4700
rect 28208 4648 28209 4700
rect 27979 4634 28209 4648
rect 26864 4608 27339 4609
rect 26864 4556 26870 4608
rect 26922 4556 26953 4608
rect 27005 4556 27035 4608
rect 27087 4556 27117 4608
rect 27169 4556 27199 4608
rect 27251 4556 27281 4608
rect 27333 4556 27339 4608
rect 26864 4512 27339 4556
rect 26864 4460 26870 4512
rect 26922 4460 26953 4512
rect 27005 4460 27035 4512
rect 27087 4460 27117 4512
rect 27169 4460 27199 4512
rect 27251 4460 27281 4512
rect 27333 4460 27339 4512
rect 26864 4416 27339 4460
rect 26864 4364 26870 4416
rect 26922 4364 26953 4416
rect 27005 4364 27035 4416
rect 27087 4364 27117 4416
rect 27169 4364 27199 4416
rect 27251 4364 27281 4416
rect 27333 4364 27339 4416
rect 26864 4320 27339 4364
rect 26864 4268 26870 4320
rect 26922 4268 26953 4320
rect 27005 4268 27035 4320
rect 27087 4268 27117 4320
rect 27169 4268 27199 4320
rect 27251 4268 27281 4320
rect 27333 4268 27339 4320
rect 26864 4224 27339 4268
rect 26864 4172 26870 4224
rect 26922 4172 26953 4224
rect 27005 4172 27035 4224
rect 27087 4172 27117 4224
rect 27169 4172 27199 4224
rect 27251 4172 27281 4224
rect 27333 4172 27339 4224
rect 27979 4582 27980 4634
rect 28032 4582 28068 4634
rect 28120 4582 28156 4634
rect 28208 4582 28209 4634
rect 27979 4568 28209 4582
rect 27979 4516 27980 4568
rect 28032 4516 28068 4568
rect 28120 4516 28156 4568
rect 28208 4516 28209 4568
rect 27979 4502 28209 4516
rect 27979 4450 27980 4502
rect 28032 4450 28068 4502
rect 28120 4450 28156 4502
rect 28208 4450 28209 4502
rect 27979 4436 28209 4450
rect 27979 4384 27980 4436
rect 28032 4384 28068 4436
rect 28120 4384 28156 4436
rect 28208 4384 28209 4436
rect 27979 4369 28209 4384
rect 27979 4317 27980 4369
rect 28032 4317 28068 4369
rect 28120 4317 28156 4369
rect 28208 4317 28209 4369
rect 27979 4302 28209 4317
rect 27979 4250 27980 4302
rect 28032 4250 28068 4302
rect 28120 4250 28156 4302
rect 28208 4250 28209 4302
rect 27979 4235 28209 4250
rect 27979 4183 27980 4235
rect 28032 4183 28068 4235
rect 28120 4183 28156 4235
rect 28208 4183 28209 4235
rect 27979 4177 28209 4183
rect 26864 4171 27339 4172
rect 17328 2561 17648 2571
rect 18030 2561 18840 2577
rect 20241 2561 21066 2577
rect 22520 2561 22931 2571
rect 23069 2561 23261 2571
rect 15566 1743 15886 1749
rect 15566 1691 15572 1743
rect 15624 1691 15636 1743
rect 15688 1691 15700 1743
rect 15752 1691 15764 1743
rect 15816 1691 15828 1743
rect 15880 1691 15886 1743
rect 15566 1675 15886 1691
rect 15566 1623 15572 1675
rect 15624 1623 15636 1675
rect 15688 1623 15700 1675
rect 15752 1623 15764 1675
rect 15816 1623 15828 1675
rect 15880 1623 15886 1675
rect 15566 1606 15886 1623
rect 15566 1554 15572 1606
rect 15624 1554 15636 1606
rect 15688 1554 15700 1606
rect 15752 1554 15764 1606
rect 15816 1554 15828 1606
rect 15880 1554 15886 1606
rect 15566 1537 15886 1554
rect 15566 1485 15572 1537
rect 15624 1485 15636 1537
rect 15688 1485 15700 1537
rect 15752 1485 15764 1537
rect 15816 1485 15828 1537
rect 15880 1485 15886 1537
rect 15566 1468 15886 1485
rect 15566 1416 15572 1468
rect 15624 1416 15636 1468
rect 15688 1416 15700 1468
rect 15752 1416 15764 1468
rect 15816 1416 15828 1468
rect 15880 1416 15886 1468
rect 15566 1410 15886 1416
rect 2714 1372 2766 1378
rect 2714 1308 2766 1320
rect 1404 1210 1456 1259
rect 1484 1210 1814 1259
rect 1842 1210 1894 1259
rect 1922 1210 1974 1259
rect 9028 1259 9075 1299
rect 2714 1210 2766 1256
rect 2794 1210 2846 1253
rect 3030 1210 3082 1253
rect 6126 1210 6178 1253
rect 6362 1210 6414 1253
rect 12886 1192 13341 1224
tri 23532 417 23557 442 se
rect 23557 417 23609 2631
rect 23709 2561 24160 2571
rect 24250 2561 24442 2571
rect 24832 2561 25014 2571
rect 25070 2561 25777 2571
rect 25835 2561 25974 2571
rect 26263 2561 26676 2571
rect 28707 2543 29181 2571
rect 29294 2543 29614 2571
rect 31793 2543 32144 2571
rect 23481 365 23487 417
rect 23539 365 23551 417
rect 23603 365 23609 417
rect 13682 -546 13798 -540
rect 13734 -598 13746 -546
rect 13682 -604 13798 -598
tri 13695 -629 13720 -604 ne
tri 13695 -1159 13720 -1134 se
rect 13720 -1159 13760 -604
tri 13760 -629 13785 -604 nw
tri 13760 -1159 13785 -1134 sw
rect 13682 -1165 13798 -1159
rect 13734 -1217 13746 -1165
rect 13682 -1223 13798 -1217
<< metal3 >>
rect 1451 28291 1670 28505
<< metal4 >>
rect 9108 31750 9327 31964
rect 13991 23755 14416 24626
rect 8628 17004 9031 17032
rect 8298 16732 9031 17004
rect 8628 16675 9031 16732
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 1 0 23481 0 1 365
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform 0 -1 13798 1 0 -1223
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1704896540
transform 0 -1 13798 1 0 -604
box 0 0 1 1
use sky130_fd_io__sio_odrvr  sky130_fd_io__sio_odrvr_0
timestamp 1704896540
transform 1 0 141 0 1 152
box -3034 -367 33934 42251
use sky130_fd_io__sio_opath_sub  sky130_fd_io__sio_opath_sub_0
timestamp 1704896540
transform 1 0 478 0 1 -1111
box -2923 1361 23223 13618
<< labels >>
flabel metal1 s 17512 6272 17512 6272 3 FreeSans 200 0 0 0 vreg_en_h
flabel metal1 s 17512 6272 17512 6272 3 FreeSans 200 0 0 0 vreg_en_h
flabel metal1 s 2121 2130 2170 2163 3 FreeSans 300 0 0 0 hld_i_vpwr
port 3 nsew
flabel metal1 s 17455 6055 17455 6055 0 FreeSans 200 0 0 0 drvhi_h
flabel metal1 s 17511 6364 17511 6364 3 FreeSans 200 0 0 0 slow_h_n
flabel metal1 s 17511 6364 17511 6364 3 FreeSans 200 0 0 0 slow_h_n
flabel metal1 s 17526 6132 17526 6132 3 FreeSans 200 0 0 0 puen_reg_h
flabel metal1 s 17526 6132 17526 6132 3 FreeSans 200 0 0 0 puen_reg_h
flabel metal1 s 17521 7481 17521 7481 3 FreeSans 200 0 0 0 pu_h_n<5>
flabel metal1 s 17521 7481 17521 7481 3 FreeSans 200 0 0 0 pu_h_n<5>
flabel metal1 s 17521 7595 17521 7595 3 FreeSans 200 0 0 0 pu_h_n<4>
flabel metal1 s 17521 7595 17521 7595 3 FreeSans 200 0 0 0 pu_h_n<4>
flabel metal1 s 17521 7356 17521 7356 3 FreeSans 200 0 0 0 sio_reg_hifreq_h
flabel metal1 s 17521 7356 17521 7356 3 FreeSans 200 0 0 0 sio_reg_hifreq_h
flabel metal1 s 17526 6052 17526 6052 3 FreeSans 200 0 0 0 drvhi_h
flabel metal1 s 17526 6052 17526 6052 3 FreeSans 200 0 0 0 drvhi_h
flabel metal1 s 17249 4880 17249 4880 0 FreeSans 200 0 0 0 oe_hs_h
flabel metal1 s 17249 4880 17249 4880 0 FreeSans 200 0 0 0 oe_hs_h
flabel metal1 s 17455 6269 17455 6269 0 FreeSans 200 0 0 0 vreg_en_h
flabel metal1 s 16508 2959 16518 3161 7 FreeSans 200 0 0 0 vpwr_ka
port 4 nsew
flabel metal1 s 6715 3189 6755 3319 3 FreeSans 300 180 0 0 vgnd
port 5 nsew
flabel metal1 s 16501 3189 16518 3319 7 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal1 s 16623 731 16663 933 3 FreeSans 300 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 6715 3347 6755 3549 3 FreeSans 300 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 16507 3347 16518 3549 7 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 478 6940 520 7070 3 FreeSans 200 0 0 0 vgnd_io
port 6 nsew
flabel metal1 s 6715 2198 6755 2400 3 FreeSans 300 180 0 0 vgnd
port 5 nsew
flabel metal1 s 16505 2198 16519 2400 7 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal1 s 8812 12746 8812 12746 0 FreeSans 200 0 0 0 pd_h<0>
flabel metal1 s 6758 12746 6758 12746 0 FreeSans 200 0 0 0 pd_h<1>
flabel metal1 s 13726 6802 13726 6802 0 FreeSans 200 180 0 0 pd_h<2>
flabel metal1 s 13698 7910 13698 7910 0 FreeSans 200 0 0 0 pd_h<3>
flabel metal1 s 1880 12921 1880 12921 0 FreeSans 200 0 0 0 pu_h_n<0>
flabel metal1 s 106 11448 106 11448 0 FreeSans 200 0 0 0 pu_h_n<1>
flabel metal1 s 139 12292 139 12292 0 FreeSans 200 0 0 0 pu_h_n<2>
flabel metal1 s 137 12404 137 12404 0 FreeSans 200 0 0 0 pu_h_n<3>
flabel metal1 s 4549 2556 4583 2590 0 FreeSans 200 0 0 0 vreg_en
port 7 nsew
flabel metal1 s 9434 1339 9467 1372 0 FreeSans 200 0 0 0 oe_n
port 8 nsew
flabel metal1 s 5450 1175 5487 1209 0 FreeSans 200 0 0 0 hld_i_h_n
port 9 nsew
flabel metal1 s 10606 1339 10640 1373 0 FreeSans 400 0 0 0 din
port 10 nsew
flabel metal1 s 17455 7359 17455 7359 0 FreeSans 200 0 0 0 sio_reg_hifreq_h
flabel metal1 s 17455 7599 17455 7599 0 FreeSans 200 0 0 0 pu_h_n<4>
flabel metal1 s 15779 7802 15813 8070 3 FreeSans 200 90 0 0 vcc_io
port 2 nsew
flabel metal1 s 17455 7485 17455 7485 0 FreeSans 200 0 0 0 pu_h_n<5>
flabel metal1 s 17455 6134 17455 6134 0 FreeSans 200 0 0 0 puen_reg_h
flabel metal1 s 17455 6366 17455 6366 0 FreeSans 200 0 0 0 slow_h_n
flabel metal1 s 15796 7936 15796 7936 3 FreeSans 200 90 0 0 vcc_io
flabel metal1 s 15796 7936 15796 7936 0 FreeSans 400 0 0 0 vcc_io
flabel metal4 s 13991 23755 14416 24626 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal4 s 8628 16675 9031 17032 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal4 s 9108 31750 9327 31964 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal4 s 14023 23777 14404 24574 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal4 s 9117 31765 9312 31948 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal4 s 9217 31857 9217 31857 0 FreeSans 400 0 0 0 pad
flabel metal4 s 14204 24191 14204 24191 0 FreeSans 400 0 0 0 pad
flabel metal4 s 9217 31857 9217 31857 0 FreeSans 400 0 0 0 pad
flabel metal4 s 14204 24191 14204 24191 0 FreeSans 400 0 0 0 pad
flabel metal4 s 8298 16732 8634 17004 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal4 s 14213 24176 14213 24176 0 FreeSans 200 0 0 0 pad
flabel metal4 s 9215 31857 9215 31857 0 FreeSans 200 0 0 0 pad
flabel metal3 s 1451 28291 1670 28505 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal3 s 1472 28330 1647 28473 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal3 s 1561 28398 1561 28398 0 FreeSans 400 0 0 0 pad
flabel metal3 s 1561 28398 1561 28398 0 FreeSans 400 0 0 0 pad
flabel metal3 s 1559 28401 1559 28401 0 FreeSans 200 0 0 0 pad
flabel metal2 s 23557 2561 23609 2631 3 FreeSans 200 90 0 0 od_h
port 12 nsew
flabel metal2 s 23583 2596 23583 2596 3 FreeSans 200 90 0 0 od_h
flabel metal2 s 20600 23528 20822 23602 0 FreeSans 400 0 0 0 vgnd_io
port 6 nsew
flabel metal2 s 20711 23565 20711 23565 0 FreeSans 400 0 0 0 vgnd_io
flabel metal2 s 29294 2543 29614 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 26263 2561 26676 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 25070 2561 25777 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 23709 2561 24160 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 22520 2561 22931 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 9028 1259 9075 1299 3 FreeSans 300 0 0 0 hld_i_ovr_h
port 13 nsew
flabel metal2 s 29454 2557 29454 2557 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 26505 2566 26505 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 25430 2566 25430 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 23934 2566 23934 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 31793 2543 32144 2571 0 FreeSans 200 0 0 0 vpwr_ka
port 4 nsew
flabel metal2 s 31606 23371 31750 23506 0 FreeSans 200 0 0 0 vpwr_ka
port 4 nsew
flabel metal2 s 31968 2557 31968 2557 0 FreeSans 200 0 0 0 vpwr_ka
flabel metal2 s 31678 23438 31678 23438 0 FreeSans 200 0 0 0 vpwr_ka
flabel metal2 s 29454 2557 29454 2557 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 26505 2566 26505 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 25430 2566 25430 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 23934 2566 23934 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 22725 2566 22725 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 29454 2557 29454 2557 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 26505 2566 26505 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 25430 2566 25430 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 23934 2567 23934 2567 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 22725 2566 22725 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 20711 23565 20711 23565 0 FreeSans 400 0 0 0 vgnd_io
flabel metal2 s 22725 2566 22725 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 25835 2561 25974 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 24832 2561 25014 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 24250 2561 24442 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 23069 2561 23261 2571 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 20711 23565 20711 23565 0 FreeSans 400 0 0 0 vgnd_io
flabel metal2 s 20241 2561 21066 2577 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 25968 2566 25968 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 24928 2566 24928 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 24346 2566 24346 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 25968 2566 25968 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 24928 2566 24928 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 23165 2566 23165 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 20653 2569 20653 2569 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 31968 2557 31968 2557 0 FreeSans 200 0 0 0 vpwr_ka
flabel metal2 s 31678 23438 31678 23438 0 FreeSans 200 0 0 0 vpwr_ka
flabel metal2 s 31968 2557 31968 2557 0 FreeSans 200 0 0 0 vpwr_ka
flabel metal2 s 31678 23438 31678 23438 0 FreeSans 200 0 0 0 vpwr_ka
flabel metal2 s 31830 23366 31958 23506 7 FreeSans 200 90 0 0 voutref
port 14 nsew
flabel metal2 s 31894 23436 31894 23436 7 FreeSans 200 90 0 0 voutref
flabel metal2 s 28707 2543 29181 2571 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 18030 2561 18840 2577 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 2967 13103 3235 13137 3 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 28944 2557 28944 2557 0 FreeSans 200 0 0 0 vcc_io
flabel metal2 s 18435 2569 18435 2569 0 FreeSans 200 0 0 0 vcc_io
flabel metal2 s 17102 13103 17160 13161 3 FreeSans 200 90 0 0 tie_lo_esd
port 15 nsew
flabel metal2 s 17131 13132 17131 13132 3 FreeSans 200 90 0 0 tie_lo_esd
flabel metal2 s 16882 13131 16882 13131 3 FreeSans 200 90 0 0 pd_h<3>
flabel metal2 s 16882 13131 16882 13131 3 FreeSans 200 90 0 0 pd_h<3>
flabel metal2 s 16198 13131 16198 13131 3 FreeSans 200 90 0 0 pd_h<2>
flabel metal2 s 23583 2596 23583 2596 3 FreeSans 200 90 0 0 od_h
flabel metal2 s 23583 2596 23583 2596 3 FreeSans 200 90 0 0 od_h
flabel metal2 s 32016 23366 32144 23506 7 FreeSans 200 90 0 0 refleak_bias
port 16 nsew
flabel metal2 s 32080 23436 32080 23436 7 FreeSans 200 90 0 0 refleak_bias
flabel metal2 s 17328 2561 17648 2571 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal2 s 17328 13103 17648 13168 0 FreeSans 200 0 0 0 pad
port 11 nsew
flabel metal2 s 17488 2566 17488 2566 0 FreeSans 200 0 0 0 pad
flabel metal2 s 17488 13135 17488 13135 0 FreeSans 200 0 0 0 pad
flabel metal2 s 12886 1192 13341 1224 0 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal2 s 1842 1210 1894 1259 3 FreeSans 200 90 0 0 slow
port 17 nsew
flabel metal2 s 2714 1210 2766 1253 3 FreeSans 200 90 0 0 od_h
port 12 nsew
flabel metal2 s 6362 1210 6414 1253 3 FreeSans 200 90 0 0 dm_h_n<2>
port 18 nsew
flabel metal2 s 2794 1210 2846 1253 3 FreeSans 200 90 0 0 dm_h_n<1>
port 19 nsew
flabel metal2 s 1404 1210 1456 1259 3 FreeSans 200 90 0 0 dm_h_n<0>
port 20 nsew
flabel metal2 s 6126 1210 6178 1253 3 FreeSans 200 90 0 0 dm_h<2>
port 21 nsew
flabel metal2 s 3030 1210 3082 1253 3 FreeSans 200 90 0 0 dm_h<1>
port 22 nsew
flabel metal2 s 1922 1210 1974 1259 3 FreeSans 200 90 0 0 dm_h<0>
port 23 nsew
flabel metal2 s 18435 2569 18435 2569 0 FreeSans 200 0 0 0 vcc_io
flabel metal2 s 28944 2557 28944 2557 0 FreeSans 200 0 0 0 vcc_io
flabel metal2 s 18435 2569 18435 2569 0 FreeSans 200 0 0 0 vcc_io
flabel metal2 s 28944 2557 28944 2557 0 FreeSans 200 0 0 0 vcc_io
flabel metal2 s 20653 2569 20653 2569 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 23165 2566 23165 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 24346 2566 24346 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 24928 2566 24928 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 25968 2566 25968 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 20653 2569 20653 2569 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 23165 2566 23165 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 24346 2566 24346 2566 0 FreeSans 200 0 0 0 vgnd
flabel metal2 s 18435 2569 18435 2569 0 FreeSans 400 0 0 0 vcc_io
flabel metal2 s 24346 2566 24346 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 23165 2566 23165 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 20654 2569 20654 2569 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 17488 13136 17488 13136 0 FreeSans 400 0 0 0 pad
flabel metal2 s 17488 2566 17488 2566 0 FreeSans 400 0 0 0 pad
flabel metal2 s 32080 23436 32080 23436 0 FreeSans 400 0 0 0 refleak_bias
flabel metal2 s 23583 2596 23583 2596 0 FreeSans 400 0 0 0 od_h
flabel metal2 s 17131 13132 17131 13132 0 FreeSans 400 0 0 0 tie_lo_esd
flabel metal2 s 18435 2569 18435 2569 0 FreeSans 400 0 0 0 vcc_io
flabel metal2 s 28944 2557 28944 2557 0 FreeSans 400 0 0 0 vcc_io
flabel metal2 s 18435 2569 18435 2569 0 FreeSans 400 0 0 0 vcc_io
flabel metal2 s 28944 2557 28944 2557 0 FreeSans 400 0 0 0 vcc_io
flabel metal2 s 31894 23436 31894 23436 0 FreeSans 400 0 0 0 voutref
flabel metal2 s 31678 23439 31678 23439 0 FreeSans 400 0 0 0 vpwr_ka
flabel metal2 s 31969 2557 31969 2557 0 FreeSans 400 0 0 0 vpwr_ka
flabel metal2 s 20654 2569 20654 2569 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 22726 2566 22726 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 23935 2566 23935 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 25423 2566 25423 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 26470 2566 26470 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 29454 2557 29454 2557 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 20711 23565 20711 23565 0 FreeSans 400 0 0 0 vgnd_io
flabel metal2 s 20711 23565 20711 23565 0 FreeSans 400 0 0 0 vgnd_io
flabel metal2 s 23583 2596 23583 2596 0 FreeSans 400 0 0 0 od_h
flabel metal2 s 23583 2596 23583 2596 0 FreeSans 400 0 0 0 od_h
flabel metal2 s 24923 2566 24923 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 25905 2566 25905 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 23165 2566 23165 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 24346 2566 24346 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 24923 2566 24923 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 25905 2566 25905 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 20654 2569 20654 2569 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 23165 2566 23165 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 24346 2566 24346 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 24923 2566 24923 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 25905 2566 25905 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 20711 23565 20711 23565 0 FreeSans 400 0 0 0 vgnd_io
flabel metal2 s 22726 2566 22726 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 23935 2566 23935 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 25423 2566 25423 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 26470 2566 26470 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 29454 2557 29454 2557 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 31678 23439 31678 23439 0 FreeSans 400 0 0 0 vpwr_ka
flabel metal2 s 31969 2557 31969 2557 0 FreeSans 400 0 0 0 vpwr_ka
flabel metal2 s 31678 23439 31678 23439 0 FreeSans 400 0 0 0 vpwr_ka
flabel metal2 s 31969 2557 31969 2557 0 FreeSans 400 0 0 0 vpwr_ka
flabel metal2 s 22726 2566 22726 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 23935 2566 23935 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 25423 2566 25423 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 26470 2566 26470 2566 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 29454 2557 29454 2557 0 FreeSans 400 0 0 0 vgnd
flabel metal2 s 1484 1210 1814 1259 0 FreeSans 200 0 0 0 vpwr
port 24 nsew
flabel metal2 s 31830 23444 31958 23506 0 FreeSans 200 0 0 0 voutref
port 14 nsew
flabel metal2 s 32016 23442 32144 23506 0 FreeSans 200 0 0 0 refleak_bias
port 16 nsew
flabel metal2 s 28944 2557 28944 2557 0 FreeSans 400 0 0 0 vcc_io
<< properties >>
string GDS_END 100633310
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 100320590
string path 68.500 31.250 68.500 34.450 
<< end >>
