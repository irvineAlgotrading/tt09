magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< poly >>
rect 12348 -69 12485 -52
rect 14625 -69 14762 -52
rect 12348 -85 12551 -69
rect 12348 -119 12365 -85
rect 12399 -119 12433 -85
rect 12467 -119 12501 -85
rect 12535 -119 12551 -85
rect 12348 -135 12551 -119
rect 14559 -85 14762 -69
rect 14559 -119 14575 -85
rect 14609 -119 14643 -85
rect 14677 -119 14711 -85
rect 14745 -119 14762 -85
rect 14559 -135 14762 -119
rect 12348 -152 12485 -135
rect 14625 -152 14762 -135
<< polycont >>
rect 12365 -119 12399 -85
rect 12433 -119 12467 -85
rect 12501 -119 12535 -85
rect 14575 -119 14609 -85
rect 14643 -119 14677 -85
rect 14711 -119 14745 -85
<< locali >>
rect 14559 -38 14761 -32
rect 12349 -85 12551 -69
rect 12349 -95 12365 -85
rect 12349 -129 12362 -95
rect 12399 -119 12433 -85
rect 12467 -95 12501 -85
rect 12535 -89 12551 -85
rect 14559 -72 14571 -38
rect 14605 -72 14643 -38
rect 14677 -72 14715 -38
rect 14749 -72 14761 -38
rect 14559 -85 14761 -72
rect 12535 -95 12552 -89
rect 12468 -119 12501 -95
rect 12396 -129 12434 -119
rect 12468 -129 12506 -119
rect 12540 -129 12552 -95
rect 12349 -135 12552 -129
rect 14559 -119 14575 -85
rect 14609 -119 14643 -85
rect 14677 -119 14711 -85
rect 14745 -119 14761 -85
rect 14559 -120 14761 -119
rect 14559 -154 14571 -120
rect 14605 -154 14643 -120
rect 14677 -154 14715 -120
rect 14749 -154 14761 -120
rect 14559 -160 14761 -154
<< viali >>
rect 12362 -119 12365 -95
rect 12365 -119 12396 -95
rect 14571 -72 14605 -38
rect 14643 -72 14677 -38
rect 14715 -72 14749 -38
rect 12434 -119 12467 -95
rect 12467 -119 12468 -95
rect 12506 -119 12535 -95
rect 12535 -119 12540 -95
rect 12362 -129 12396 -119
rect 12434 -129 12468 -119
rect 12506 -129 12540 -119
rect 14571 -154 14605 -120
rect 14643 -154 14677 -120
rect 14715 -154 14749 -120
<< metal1 >>
rect 1427 1478 2325 1608
rect 2455 1478 2755 1608
rect 2885 1602 3747 1608
rect 2885 1550 3593 1602
rect 3645 1550 3671 1602
rect 3723 1550 3747 1602
rect 2885 1536 3747 1550
rect 2885 1484 3593 1536
rect 3645 1484 3671 1536
rect 3723 1484 3747 1536
rect 2885 1478 3747 1484
rect 4439 1478 5301 1608
rect 5431 1478 7285 1608
rect 7367 1556 8282 1608
rect 8334 1556 8349 1608
rect 8401 1556 8407 1608
rect 7367 1530 8407 1556
rect 7367 1478 8282 1530
rect 8334 1478 8349 1530
rect 8401 1478 8407 1530
rect 8837 1556 9132 1608
rect 9184 1556 9199 1608
rect 9251 1556 9267 1608
rect 9319 1556 9335 1608
rect 9387 1556 9403 1608
rect 9455 1556 9471 1608
rect 9523 1556 9539 1608
rect 9591 1556 9607 1608
rect 9659 1556 9675 1608
rect 9727 1556 9733 1608
rect 8837 1530 9733 1556
rect 8837 1478 9132 1530
rect 9184 1478 9199 1530
rect 9251 1478 9267 1530
rect 9319 1478 9335 1530
rect 9387 1478 9403 1530
rect 9455 1478 9471 1530
rect 9523 1478 9539 1530
rect 9591 1478 9607 1530
rect 9659 1478 9675 1530
rect 9727 1478 9733 1530
rect 10391 1556 10950 1608
rect 11002 1556 11025 1608
rect 11077 1556 11100 1608
rect 11152 1556 11175 1608
rect 11227 1556 11250 1608
rect 11302 1556 11325 1608
rect 11377 1556 11383 1608
rect 10391 1530 11383 1556
rect 10391 1478 10950 1530
rect 11002 1478 11025 1530
rect 11077 1478 11100 1530
rect 11152 1478 11175 1530
rect 11227 1478 11250 1530
rect 11302 1478 11325 1530
rect 11377 1478 11383 1530
rect 11745 1556 12371 1608
rect 12423 1556 12437 1608
rect 12489 1556 12503 1608
rect 12555 1556 12570 1608
rect 12622 1556 12637 1608
rect 12689 1556 12704 1608
rect 12756 1556 12771 1608
rect 12823 1556 12829 1608
rect 11745 1530 12829 1556
rect 11745 1478 12371 1530
rect 12423 1478 12437 1530
rect 12489 1478 12503 1530
rect 12555 1478 12570 1530
rect 12622 1478 12637 1530
rect 12689 1478 12704 1530
rect 12756 1478 12771 1530
rect 12823 1478 12829 1530
rect 13237 1601 13367 1608
rect 13237 1549 13243 1601
rect 13295 1549 13309 1601
rect 13361 1549 13367 1601
rect 13237 1537 13367 1549
rect 13237 1485 13243 1537
rect 13295 1485 13309 1537
rect 13361 1485 13367 1537
rect 13237 1478 13367 1485
rect 13667 1601 13797 1608
rect 13667 1549 13673 1601
rect 13725 1549 13739 1601
rect 13791 1549 13797 1601
rect 13667 1537 13797 1549
rect 13667 1485 13673 1537
rect 13725 1485 13739 1537
rect 13791 1485 13797 1537
rect 13667 1478 13797 1485
rect 14229 1601 14587 1608
rect 14229 1549 14235 1601
rect 14287 1549 14301 1601
rect 14353 1549 14587 1601
rect 14229 1537 14587 1549
rect 14229 1485 14235 1537
rect 14287 1485 14301 1537
rect 14353 1485 14587 1537
rect 14229 1478 14587 1485
rect 12712 661 12811 745
rect 11936 151 11942 203
rect 11994 151 12015 203
rect 12067 151 12087 203
rect 12139 151 14108 203
rect 11936 150 14108 151
tri 14108 150 14161 203 sw
rect 11936 123 14161 150
rect 11936 71 11942 123
rect 11994 71 12015 123
rect 12067 71 12087 123
rect 12139 71 14161 123
tri 14058 -32 14161 71 ne
tri 14161 -32 14343 150 sw
tri 14161 -38 14167 -32 ne
rect 14167 -38 14761 -32
tri 14167 -72 14201 -38 ne
rect 14201 -72 14571 -38
rect 14605 -72 14643 -38
rect 14677 -72 14715 -38
rect 14749 -72 14761 -38
tri 14201 -89 14218 -72 ne
rect 14218 -89 14761 -72
rect 12003 -141 12009 -89
rect 12061 -141 12073 -89
rect 12125 -95 12552 -89
rect 12125 -129 12362 -95
rect 12396 -129 12434 -95
rect 12468 -129 12506 -95
rect 12540 -129 12552 -95
tri 14218 -120 14249 -89 ne
rect 14249 -120 14761 -89
rect 12125 -141 12552 -129
tri 14249 -141 14270 -120 ne
rect 14270 -141 14571 -120
tri 14270 -154 14283 -141 ne
rect 14283 -154 14571 -141
rect 14605 -154 14643 -120
rect 14677 -154 14715 -120
rect 14749 -154 14761 -120
tri 14283 -160 14289 -154 ne
rect 14289 -160 14761 -154
tri 14471 -317 14498 -290 se
rect 14498 -317 14725 -290
tri 7986 -391 8060 -317 se
rect 8060 -369 10681 -317
rect 10733 -369 10745 -317
rect 10797 -369 11429 -317
rect 11481 -369 11493 -317
rect 11545 -369 12856 -317
rect 12908 -369 12920 -317
rect 12972 -369 13141 -317
rect 13193 -369 13207 -317
rect 13259 -369 14082 -317
rect 14134 -369 14146 -317
rect 14198 -342 14725 -317
rect 14777 -342 14789 -290
rect 14841 -342 14853 -290
rect 14905 -342 14917 -290
rect 14969 -342 14975 -290
rect 14198 -369 14550 -342
tri 14550 -369 14577 -342 nw
tri 8060 -391 8082 -369 nw
tri 14613 -391 14629 -375 se
rect 14629 -391 14905 -375
tri 7975 -402 7986 -391 se
rect 7986 -402 7997 -391
rect 7615 -454 7621 -402
rect 7673 -454 7685 -402
rect 7737 -454 7997 -402
tri 7997 -454 8060 -391 nw
tri 14602 -402 14613 -391 se
rect 14613 -402 14905 -391
rect 8246 -454 8252 -402
rect 8304 -454 8360 -402
rect 8412 -454 10446 -402
rect 10498 -454 10510 -402
rect 10562 -454 11194 -402
rect 11246 -454 11258 -402
rect 11310 -454 12615 -402
rect 12667 -454 12679 -402
rect 12731 -454 13845 -402
rect 13897 -454 13909 -402
rect 13961 -454 14539 -402
rect 14591 -454 14603 -402
rect 14655 -427 14905 -402
rect 14957 -427 14970 -375
rect 15022 -427 15028 -375
rect 14655 -454 14665 -427
tri 14665 -454 14692 -427 nw
tri 14689 -482 14716 -455 se
rect 14716 -461 14954 -455
rect 14716 -482 14902 -461
rect 7649 -534 10204 -482
rect 10256 -534 10268 -482
rect 10320 -534 10952 -482
rect 11004 -534 11016 -482
rect 11068 -534 12006 -482
rect 12058 -534 12070 -482
rect 12122 -534 12373 -482
rect 12425 -534 12437 -482
rect 12489 -534 13600 -482
rect 13652 -534 13664 -482
rect 13716 -534 14294 -482
rect 14346 -534 14358 -482
rect 14410 -507 14902 -482
rect 14410 -534 14753 -507
tri 14753 -534 14780 -507 nw
tri 14858 -534 14885 -507 ne
rect 14885 -513 14902 -507
rect 14885 -525 14954 -513
rect 14885 -534 14902 -525
tri 14885 -551 14902 -534 ne
rect 14902 -583 14954 -577
<< via1 >>
rect 3593 1550 3645 1602
rect 3671 1550 3723 1602
rect 3593 1484 3645 1536
rect 3671 1484 3723 1536
rect 8282 1556 8334 1608
rect 8349 1556 8401 1608
rect 8282 1478 8334 1530
rect 8349 1478 8401 1530
rect 9132 1556 9184 1608
rect 9199 1556 9251 1608
rect 9267 1556 9319 1608
rect 9335 1556 9387 1608
rect 9403 1556 9455 1608
rect 9471 1556 9523 1608
rect 9539 1556 9591 1608
rect 9607 1556 9659 1608
rect 9675 1556 9727 1608
rect 9132 1478 9184 1530
rect 9199 1478 9251 1530
rect 9267 1478 9319 1530
rect 9335 1478 9387 1530
rect 9403 1478 9455 1530
rect 9471 1478 9523 1530
rect 9539 1478 9591 1530
rect 9607 1478 9659 1530
rect 9675 1478 9727 1530
rect 10950 1556 11002 1608
rect 11025 1556 11077 1608
rect 11100 1556 11152 1608
rect 11175 1556 11227 1608
rect 11250 1556 11302 1608
rect 11325 1556 11377 1608
rect 10950 1478 11002 1530
rect 11025 1478 11077 1530
rect 11100 1478 11152 1530
rect 11175 1478 11227 1530
rect 11250 1478 11302 1530
rect 11325 1478 11377 1530
rect 12371 1556 12423 1608
rect 12437 1556 12489 1608
rect 12503 1556 12555 1608
rect 12570 1556 12622 1608
rect 12637 1556 12689 1608
rect 12704 1556 12756 1608
rect 12771 1556 12823 1608
rect 12371 1478 12423 1530
rect 12437 1478 12489 1530
rect 12503 1478 12555 1530
rect 12570 1478 12622 1530
rect 12637 1478 12689 1530
rect 12704 1478 12756 1530
rect 12771 1478 12823 1530
rect 13243 1549 13295 1601
rect 13309 1549 13361 1601
rect 13243 1485 13295 1537
rect 13309 1485 13361 1537
rect 13673 1549 13725 1601
rect 13739 1549 13791 1601
rect 13673 1485 13725 1537
rect 13739 1485 13791 1537
rect 14235 1549 14287 1601
rect 14301 1549 14353 1601
rect 14235 1485 14287 1537
rect 14301 1485 14353 1537
rect 11942 151 11994 203
rect 12015 151 12067 203
rect 12087 151 12139 203
rect 11942 71 11994 123
rect 12015 71 12067 123
rect 12087 71 12139 123
rect 12009 -141 12061 -89
rect 12073 -141 12125 -89
rect 10681 -369 10733 -317
rect 10745 -369 10797 -317
rect 11429 -369 11481 -317
rect 11493 -369 11545 -317
rect 12856 -369 12908 -317
rect 12920 -369 12972 -317
rect 13141 -369 13193 -317
rect 13207 -369 13259 -317
rect 14082 -369 14134 -317
rect 14146 -369 14198 -317
rect 14725 -342 14777 -290
rect 14789 -342 14841 -290
rect 14853 -342 14905 -290
rect 14917 -342 14969 -290
rect 7621 -454 7673 -402
rect 7685 -454 7737 -402
rect 8252 -454 8304 -402
rect 8360 -454 8412 -402
rect 10446 -454 10498 -402
rect 10510 -454 10562 -402
rect 11194 -454 11246 -402
rect 11258 -454 11310 -402
rect 12615 -454 12667 -402
rect 12679 -454 12731 -402
rect 13845 -454 13897 -402
rect 13909 -454 13961 -402
rect 14539 -454 14591 -402
rect 14603 -454 14655 -402
rect 14905 -427 14957 -375
rect 14970 -427 15022 -375
rect 10204 -534 10256 -482
rect 10268 -534 10320 -482
rect 10952 -534 11004 -482
rect 11016 -534 11068 -482
rect 12006 -534 12058 -482
rect 12070 -534 12122 -482
rect 12373 -534 12425 -482
rect 12437 -534 12489 -482
rect 13600 -534 13652 -482
rect 13664 -534 13716 -482
rect 14294 -534 14346 -482
rect 14358 -534 14410 -482
rect 14902 -513 14954 -461
rect 14902 -577 14954 -525
<< metal2 >>
rect 3593 1602 3723 1608
rect 3645 1550 3671 1602
rect 3593 1536 3723 1550
rect 3645 1484 3671 1536
rect 3593 -664 3723 1484
rect 8246 1556 8282 1608
rect 8334 1556 8349 1608
rect 8401 1556 8418 1608
rect 8246 1530 8418 1556
rect 8246 1478 8282 1530
rect 8334 1478 8349 1530
rect 8401 1478 8418 1530
rect 9126 1556 9132 1608
rect 9184 1556 9199 1608
rect 9251 1556 9267 1608
rect 9319 1556 9335 1608
rect 9387 1556 9403 1608
rect 9455 1556 9471 1608
rect 9523 1556 9539 1608
rect 9591 1556 9607 1608
rect 9659 1556 9675 1608
rect 9727 1556 10531 1608
rect 9126 1530 10531 1556
rect 9126 1478 9132 1530
rect 9184 1478 9199 1530
rect 9251 1478 9267 1530
rect 9319 1478 9335 1530
rect 9387 1478 9403 1530
rect 9455 1478 9471 1530
rect 9523 1478 9539 1530
rect 9591 1478 9607 1530
rect 9659 1478 9675 1530
rect 9727 1478 10531 1530
rect 8246 -402 8418 1478
tri 9939 1221 10196 1478 ne
rect 10196 260 10531 1478
rect 10944 1556 10950 1608
rect 11002 1556 11025 1608
rect 11077 1556 11100 1608
rect 11152 1556 11175 1608
rect 11227 1556 11250 1608
rect 11302 1556 11325 1608
rect 11377 1556 11383 1608
rect 10944 1530 11383 1556
rect 10944 1478 10950 1530
rect 11002 1478 11025 1530
rect 11077 1478 11100 1530
rect 11152 1478 11175 1530
rect 11227 1478 11250 1530
rect 11302 1478 11325 1530
rect 11377 1478 11383 1530
tri 10531 260 10803 532 sw
rect 10196 146 10803 260
rect 10196 123 10335 146
tri 10335 123 10358 146 nw
tri 10405 123 10428 146 ne
rect 10428 123 10577 146
tri 10577 123 10600 146 nw
tri 10639 123 10662 146 ne
rect 10662 123 10803 146
rect 10196 94 10326 123
tri 10326 114 10335 123 nw
tri 10428 114 10437 123 ne
rect 10437 114 10568 123
tri 10568 114 10577 123 nw
tri 10662 114 10671 123 ne
rect 10671 114 10803 123
tri 10437 113 10438 114 ne
rect 10197 92 10325 93
rect 10438 94 10568 114
tri 10671 112 10673 114 ne
rect 10439 92 10567 93
rect 10673 94 10803 114
rect 10674 92 10802 93
rect 10944 260 11383 1478
rect 12365 1556 12371 1608
rect 12423 1556 12437 1608
rect 12489 1556 12503 1608
rect 12555 1556 12570 1608
rect 12622 1556 12637 1608
rect 12689 1556 12704 1608
rect 12756 1556 12771 1608
rect 12823 1556 12829 1608
tri 13198 1601 13205 1608 se
rect 13205 1601 13367 1608
rect 12365 1530 12829 1556
tri 13146 1549 13198 1601 se
rect 13198 1549 13243 1601
rect 13295 1549 13309 1601
rect 13361 1549 13367 1601
rect 12365 1478 12371 1530
rect 12423 1478 12437 1530
rect 12489 1478 12503 1530
rect 12555 1478 12570 1530
rect 12622 1478 12637 1530
rect 12689 1478 12704 1530
rect 12756 1478 12771 1530
rect 12823 1478 12829 1530
tri 11383 260 11551 428 sw
rect 10944 146 11551 260
rect 12365 284 12829 1478
tri 13135 1538 13146 1549 se
rect 13146 1538 13367 1549
rect 13135 1537 13367 1538
rect 13135 1485 13243 1537
rect 13295 1485 13309 1537
rect 13361 1485 13367 1537
rect 13135 1478 13367 1485
rect 13667 1601 13797 1608
rect 13667 1549 13673 1601
rect 13725 1549 13739 1601
rect 13791 1549 13797 1601
rect 13667 1537 13797 1549
rect 13667 1485 13673 1537
rect 13725 1485 13739 1537
rect 13791 1485 13797 1537
tri 12829 284 12978 433 sw
rect 10944 123 11083 146
tri 11083 123 11106 146 nw
tri 11153 123 11176 146 ne
rect 11176 123 11325 146
tri 11325 123 11348 146 nw
tri 11387 123 11410 146 ne
rect 11410 123 11551 146
rect 10944 94 11074 123
tri 11074 114 11083 123 nw
tri 11176 114 11185 123 ne
rect 11185 114 11316 123
tri 11316 114 11325 123 nw
tri 11410 114 11419 123 ne
rect 11419 114 11551 123
tri 11185 113 11186 114 ne
rect 10945 92 11073 93
rect 11186 94 11316 114
tri 11419 112 11421 114 ne
rect 11187 92 11315 93
rect 11421 94 11551 114
rect 11422 92 11550 93
rect 11931 151 11940 207
rect 11996 203 12064 207
rect 12120 203 12145 207
rect 11996 151 12015 203
rect 12139 151 12145 203
rect 11931 123 12145 151
rect 11931 121 11942 123
rect 11994 121 12015 123
rect 12067 121 12087 123
rect 10673 -208 10803 92
rect 11186 -208 11316 92
rect 11931 65 11940 121
rect 11996 71 12015 121
rect 12139 71 12145 123
rect 11996 65 12064 71
rect 12120 65 12145 71
rect 12365 170 12978 284
rect 12365 118 12495 170
tri 12495 136 12529 170 nw
tri 12573 136 12607 170 ne
rect 12366 116 12494 117
rect 12607 118 12737 170
tri 12737 136 12771 170 nw
tri 12814 136 12848 170 ne
rect 12608 116 12736 117
rect 12848 118 12978 170
rect 12849 116 12977 117
rect 12003 -141 12009 -89
rect 12061 -141 12073 -89
rect 12125 -141 12131 -89
tri 12003 -179 12041 -141 ne
tri 7424 -454 7476 -402 se
rect 7476 -454 7621 -402
rect 7673 -454 7685 -402
rect 7737 -454 7743 -402
rect 8246 -454 8252 -402
rect 8304 -454 8360 -402
rect 8412 -454 8418 -402
rect 10197 -209 10325 -208
tri 7417 -461 7424 -454 se
rect 7424 -461 7491 -454
tri 7491 -461 7498 -454 nw
tri 7402 -476 7417 -461 se
rect 7417 -476 7476 -461
tri 7476 -476 7491 -461 nw
tri 7396 -482 7402 -476 se
rect 7402 -482 7470 -476
tri 7470 -482 7476 -476 nw
rect 10196 -482 10326 -210
rect 10439 -209 10567 -208
rect 10438 -402 10568 -210
rect 10674 -209 10802 -208
rect 10673 -317 10803 -210
rect 10673 -369 10681 -317
rect 10733 -369 10745 -317
rect 10797 -369 10803 -317
rect 10945 -209 11073 -208
rect 10438 -454 10446 -402
rect 10498 -454 10510 -402
rect 10562 -454 10568 -402
tri 7382 -496 7396 -482 se
rect 7396 -496 7418 -482
tri 4421 -534 4459 -496 se
rect 4459 -534 7418 -496
tri 7418 -534 7470 -482 nw
rect 10196 -534 10204 -482
rect 10256 -534 10268 -482
rect 10320 -534 10326 -482
rect 10944 -482 11074 -210
rect 11187 -209 11315 -208
rect 11186 -402 11316 -210
rect 11422 -209 11550 -208
rect 11421 -317 11551 -210
rect 11421 -369 11429 -317
rect 11481 -369 11493 -317
rect 11545 -369 11551 -317
rect 11186 -454 11194 -402
rect 11246 -454 11258 -402
rect 11310 -454 11316 -402
tri 12028 -454 12041 -441 se
rect 12041 -454 12093 -141
tri 12093 -179 12131 -141 nw
rect 12365 -184 12495 116
rect 12366 -185 12494 -184
tri 12093 -454 12100 -447 sw
tri 12021 -461 12028 -454 se
rect 12028 -461 12100 -454
tri 12100 -461 12107 -454 sw
rect 10944 -534 10952 -482
rect 11004 -534 11016 -482
rect 11068 -534 11074 -482
tri 12000 -482 12021 -461 se
rect 12021 -482 12107 -461
tri 12107 -482 12128 -461 sw
rect 12000 -534 12006 -482
rect 12058 -534 12070 -482
rect 12122 -534 12128 -482
rect 12365 -482 12495 -186
rect 12608 -185 12736 -184
rect 12607 -402 12737 -186
rect 12849 -185 12977 -184
rect 12848 -317 12978 -186
rect 12848 -369 12856 -317
rect 12908 -369 12920 -317
rect 12972 -369 12978 -317
rect 13135 -317 13265 1478
tri 13265 1408 13335 1478 nw
tri 13592 1147 13667 1222 se
rect 13667 1147 13797 1485
rect 14229 1601 14359 1608
rect 14229 1549 14235 1601
rect 14287 1549 14301 1601
rect 14353 1549 14359 1601
rect 14229 1537 14359 1549
rect 14229 1485 14235 1537
rect 14287 1485 14301 1537
rect 14353 1485 14359 1537
rect 14229 1357 14359 1485
tri 14229 1300 14286 1357 ne
rect 14286 1328 14359 1357
tri 14359 1328 14442 1411 sw
rect 13592 1126 13797 1147
tri 13797 1126 13893 1222 sw
rect 14286 1126 14442 1328
tri 14442 1126 14563 1247 sw
rect 13592 1012 14204 1126
rect 13592 960 13722 1012
tri 13722 978 13756 1012 nw
tri 13803 978 13837 1012 ne
rect 13593 958 13721 959
rect 13837 960 13967 1012
tri 13967 978 14001 1012 nw
tri 14040 978 14074 1012 ne
rect 13838 958 13966 959
rect 14074 960 14204 1012
rect 14075 958 14203 959
rect 14286 1012 14898 1126
rect 14286 960 14416 1012
tri 14416 978 14450 1012 nw
tri 14497 978 14531 1012 ne
rect 14287 958 14415 959
rect 14531 960 14661 1012
tri 14661 978 14695 1012 nw
tri 14734 978 14768 1012 ne
rect 14532 958 14660 959
rect 14768 960 14898 1012
rect 14769 958 14897 959
rect 13837 658 13967 958
rect 14286 658 14416 958
rect 13135 -369 13141 -317
rect 13193 -369 13207 -317
rect 13259 -369 13265 -317
rect 13593 657 13721 658
rect 12607 -454 12615 -402
rect 12667 -454 12679 -402
rect 12731 -454 12737 -402
rect 12365 -534 12373 -482
rect 12425 -534 12437 -482
rect 12489 -534 12495 -482
rect 13592 -482 13722 656
rect 13838 657 13966 658
rect 13837 -402 13967 656
rect 14075 657 14203 658
rect 14074 -317 14204 656
rect 14074 -369 14082 -317
rect 14134 -369 14146 -317
rect 14198 -369 14204 -317
rect 14287 657 14415 658
rect 13837 -454 13845 -402
rect 13897 -454 13909 -402
rect 13961 -454 13967 -402
rect 13592 -534 13600 -482
rect 13652 -534 13664 -482
rect 13716 -534 13722 -482
rect 14286 -482 14416 656
rect 14532 657 14660 658
rect 14531 -402 14661 656
rect 14769 657 14897 658
tri 14712 -290 14768 -234 se
rect 14768 -290 14898 656
tri 14898 -290 14972 -216 sw
rect 14712 -342 14725 -290
rect 14777 -342 14789 -290
rect 14841 -342 14853 -290
rect 14905 -342 14917 -290
rect 14969 -342 14975 -290
rect 14531 -454 14539 -402
rect 14591 -454 14603 -402
rect 14655 -454 14661 -402
rect 14899 -427 14905 -375
rect 14957 -427 14970 -375
rect 15022 -427 15028 -375
rect 14286 -534 14294 -482
rect 14346 -534 14358 -482
rect 14410 -534 14416 -482
rect 14902 -461 14954 -455
rect 14902 -525 14954 -513
tri 4385 -570 4421 -534 se
rect 4421 -548 7404 -534
tri 7404 -548 7418 -534 nw
rect 4421 -570 4459 -548
tri 4459 -570 4481 -548 nw
tri 4378 -577 4385 -570 se
rect 4385 -577 4452 -570
tri 4452 -577 4459 -570 nw
tri 4311 -644 4378 -577 se
rect 4378 -644 4385 -577
tri 4385 -644 4452 -577 nw
rect 14902 -583 14954 -577
tri 3593 -790 3719 -664 ne
rect 3719 -738 3723 -664
tri 4264 -691 4311 -644 se
tri 3723 -738 3770 -691 sw
tri 4237 -718 4264 -691 se
rect 4264 -718 4311 -691
tri 4311 -718 4385 -644 nw
tri 4217 -738 4237 -718 se
rect 4237 -738 4239 -718
rect 3719 -790 4239 -738
tri 4239 -790 4311 -718 nw
<< rmetal2 >>
rect 10196 93 10326 94
rect 10196 92 10197 93
rect 10325 92 10326 93
rect 10438 93 10568 94
rect 10438 92 10439 93
rect 10567 92 10568 93
rect 10673 93 10803 94
rect 10673 92 10674 93
rect 10802 92 10803 93
rect 10944 93 11074 94
rect 10944 92 10945 93
rect 11073 92 11074 93
rect 11186 93 11316 94
rect 11186 92 11187 93
rect 11315 92 11316 93
rect 11421 93 11551 94
rect 11421 92 11422 93
rect 11550 92 11551 93
rect 12365 117 12495 118
rect 12365 116 12366 117
rect 12494 116 12495 117
rect 12607 117 12737 118
rect 12607 116 12608 117
rect 12736 116 12737 117
rect 12848 117 12978 118
rect 12848 116 12849 117
rect 12977 116 12978 117
rect 10196 -209 10197 -208
rect 10325 -209 10326 -208
rect 10196 -210 10326 -209
rect 10438 -209 10439 -208
rect 10567 -209 10568 -208
rect 10438 -210 10568 -209
rect 10673 -209 10674 -208
rect 10802 -209 10803 -208
rect 10673 -210 10803 -209
rect 10944 -209 10945 -208
rect 11073 -209 11074 -208
rect 10944 -210 11074 -209
rect 11186 -209 11187 -208
rect 11315 -209 11316 -208
rect 11186 -210 11316 -209
rect 11421 -209 11422 -208
rect 11550 -209 11551 -208
rect 11421 -210 11551 -209
rect 12365 -185 12366 -184
rect 12494 -185 12495 -184
rect 12365 -186 12495 -185
rect 12607 -185 12608 -184
rect 12736 -185 12737 -184
rect 12607 -186 12737 -185
rect 12848 -185 12849 -184
rect 12977 -185 12978 -184
rect 12848 -186 12978 -185
rect 13592 959 13722 960
rect 13592 958 13593 959
rect 13721 958 13722 959
rect 13837 959 13967 960
rect 13837 958 13838 959
rect 13966 958 13967 959
rect 14074 959 14204 960
rect 14074 958 14075 959
rect 14203 958 14204 959
rect 14286 959 14416 960
rect 14286 958 14287 959
rect 14415 958 14416 959
rect 14531 959 14661 960
rect 14531 958 14532 959
rect 14660 958 14661 959
rect 14768 959 14898 960
rect 14768 958 14769 959
rect 14897 958 14898 959
rect 13592 657 13593 658
rect 13721 657 13722 658
rect 13592 656 13722 657
rect 13837 657 13838 658
rect 13966 657 13967 658
rect 13837 656 13967 657
rect 14074 657 14075 658
rect 14203 657 14204 658
rect 14074 656 14204 657
rect 14286 657 14287 658
rect 14415 657 14416 658
rect 14286 656 14416 657
rect 14531 657 14532 658
rect 14660 657 14661 658
rect 14531 656 14661 657
rect 14768 657 14769 658
rect 14897 657 14898 658
rect 14768 656 14898 657
<< via2 >>
rect 11940 203 11996 207
rect 12064 203 12120 207
rect 11940 151 11942 203
rect 11942 151 11994 203
rect 11994 151 11996 203
rect 12064 151 12067 203
rect 12067 151 12087 203
rect 12087 151 12120 203
rect 11940 71 11942 121
rect 11942 71 11994 121
rect 11994 71 11996 121
rect 12064 71 12067 121
rect 12067 71 12087 121
rect 12087 71 12120 121
rect 11940 65 11996 71
rect 12064 65 12120 71
<< metal3 >>
rect 11935 207 12125 212
rect 11935 151 11940 207
rect 11996 151 12064 207
rect 12120 151 12125 207
rect 11935 121 12125 151
rect 11935 65 11940 121
rect 11996 65 12064 121
rect 12120 65 12125 121
rect 11935 60 12125 65
use PYL1_C_CDNS_524688791850  PYL1_C_CDNS_524688791850_0
timestamp 1704896540
transform -1 0 14660 0 -1 -102
box 0 0 1 1
use PYL1_C_CDNS_524688791850  PYL1_C_CDNS_524688791850_1
timestamp 1704896540
transform 1 0 12450 0 -1 -102
box 0 0 1 1
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_0
timestamp 1704896540
transform 1 0 12535 0 1 -152
box -50 0 2090 100
use sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad  sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0
timestamp 1704896540
transform 1 0 457 0 1 346
box 36 -976 15097 5118
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_0
timestamp 1704896540
transform 0 1 12607 1 0 -238
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_1
timestamp 1704896540
transform 0 1 14768 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_2
timestamp 1704896540
transform 0 1 12848 1 0 -238
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_3
timestamp 1704896540
transform 0 1 10944 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_4
timestamp 1704896540
transform 0 1 11421 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_5
timestamp 1704896540
transform 0 1 10438 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_6
timestamp 1704896540
transform 0 1 10196 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_7
timestamp 1704896540
transform 0 1 13592 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_8
timestamp 1704896540
transform 0 1 14531 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_524688791854  sky130_fd_io__tk_em2o_CDNS_524688791854_9
timestamp 1704896540
transform 0 1 14074 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_0
timestamp 1704896540
transform 0 1 12365 1 0 -238
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_1
timestamp 1704896540
transform 0 1 11186 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_2
timestamp 1704896540
transform 0 1 10673 1 0 -262
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_3
timestamp 1704896540
transform 0 1 13837 1 0 604
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_524688791855  sky130_fd_io__tk_em2s_CDNS_524688791855_4
timestamp 1704896540
transform 0 1 14286 1 0 604
box 0 0 1 1
<< labels >>
flabel comment s 13504 -93 13504 -93 0 FreeSans 440 0 0 0 leaker
flabel metal1 s 12712 661 12811 745 3 FreeSans 520 0 0 0 vnb
port 1 nsew
flabel metal1 s 9905 -508 9905 -508 0 FreeSans 400 180 0 0 tie_hi_esd
flabel metal1 s 10299 -369 10384 -317 0 FreeSans 400 180 0 0 pu_h_n<2>
port 3 nsew
flabel metal1 s 10483 -454 10635 -402 0 FreeSans 400 180 0 0 pu_h_n<3>
port 4 nsew
<< properties >>
string GDS_END 13669710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 13650570
string path 298.375 3.400 303.125 3.400 
<< end >>
