magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -122 -66 714 1466
<< mvpmos >>
rect 0 0 160 1400
rect 216 0 376 1400
rect 432 0 592 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 592 0 642 1400
<< poly >>
rect 0 1400 160 1432
rect 0 -32 160 0
rect 216 1400 376 1432
rect 216 -32 376 0
rect 432 1400 592 1432
rect 432 -32 592 0
<< locali >>
rect -45 -4 -11 1354
rect 171 -4 205 1354
rect 387 -4 421 1354
rect 603 -4 637 1354
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_0
timestamp 1704896540
transform 1 0 376 0 1 0
box -36 -36 92 1436
use DFL1sd2_CDNS_5246887918574  DFL1sd2_CDNS_5246887918574_1
timestamp 1704896540
transform 1 0 160 0 1 0
box -36 -36 92 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 92 1436
use hvDFL1sd2_CDNS_5246887918575  hvDFL1sd2_CDNS_5246887918575_1
timestamp 1704896540
transform 1 0 592 0 1 0
box -36 -36 92 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 188 675 188 675 0 FreeSans 300 0 0 0 D
flabel comment s 404 675 404 675 0 FreeSans 300 0 0 0 S
flabel comment s 620 675 620 675 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85591968
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85589958
<< end >>
