magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< metal2 >>
rect 0 385 216 394
rect 0 0 216 9
<< via2 >>
rect 0 9 216 385
<< metal3 >>
rect -5 385 221 390
rect -5 9 0 385
rect 216 9 221 385
rect -5 4 221 9
<< properties >>
string GDS_END 91722180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91721088
<< end >>
