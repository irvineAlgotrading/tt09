magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 3444 626
<< mvnmos >>
rect 0 0 800 600
rect 856 0 1656 600
rect 1712 0 2512 600
rect 2568 0 3368 600
<< mvndiff >>
rect -50 0 0 600
rect 3368 0 3418 600
<< poly >>
rect 0 600 800 626
rect 0 -26 800 0
rect 856 600 1656 626
rect 856 -26 1656 0
rect 1712 600 2512 626
rect 1712 -26 2512 0
rect 2568 600 3368 626
rect 2568 -26 3368 0
<< locali >>
rect -45 -4 -11 538
<< metal1 >>
rect 805 -16 851 546
rect 1661 -16 1707 546
rect 2517 -16 2563 546
rect 3373 -16 3419 546
use hvDFL1sd_CDNS_52468879185311  hvDFL1sd_CDNS_52468879185311_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 626
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_0
timestamp 1704896540
transform 1 0 2512 0 1 0
box -26 -26 82 626
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_1
timestamp 1704896540
transform 1 0 1656 0 1 0
box -26 -26 82 626
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_2
timestamp 1704896540
transform 1 0 800 0 1 0
box -26 -26 82 626
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_0
timestamp 1704896540
transform 1 0 3368 0 1 0
box -26 -26 79 626
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 828 265 828 265 0 FreeSans 300 0 0 0 D
flabel comment s 1684 265 1684 265 0 FreeSans 300 0 0 0 S
flabel comment s 2540 265 2540 265 0 FreeSans 300 0 0 0 D
flabel comment s 3396 265 3396 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86900470
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86898080
<< end >>
