magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 876 2026
<< mvnnmos >>
rect 0 0 800 2000
<< mvndiff >>
rect -50 0 0 2000
rect 800 0 850 2000
<< poly >>
rect 0 2000 800 2026
rect 0 -26 800 0
<< locali >>
rect -113 -4 -11 1978
rect 811 -4 913 1978
use hvDFTPL1s_CDNS_52468879185835  hvDFTPL1s_CDNS_52468879185835_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 226 2026
use hvDFTPL1s_CDNS_52468879185835  hvDFTPL1s_CDNS_52468879185835_1
timestamp 1704896540
transform 1 0 800 0 1 0
box -26 -26 226 2026
<< labels >>
flabel comment s -62 987 -62 987 0 FreeSans 300 0 0 0 S
flabel comment s 862 987 862 987 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 96480924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96479966
<< end >>
