magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 4119 150
<< mvpmos >>
rect 0 0 4000 84
<< mvpdiff >>
rect -53 46 0 84
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 4000 46 4053 84
rect 4000 12 4011 46
rect 4045 12 4053 46
rect 4000 0 4053 12
<< mvpdiffc >>
rect -45 12 -11 46
rect 4011 12 4045 46
<< poly >>
rect 0 84 4000 116
rect 0 -32 4000 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 4011 46 4045 62
rect 4011 -4 4045 12
use DFL1sd_CDNS_52468879185322  DFL1sd_CDNS_52468879185322_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185322  DFL1sd_CDNS_52468879185322_1
timestamp 1704896540
transform 1 0 4000 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 4028 29 4028 29 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6071064
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6070050
<< end >>
