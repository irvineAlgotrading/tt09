magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 3 3 93
rect 93 3 96 93
<< via1 >>
rect 3 3 93 93
<< metal2 >>
rect 3 93 93 96
rect 3 0 93 3
<< properties >>
string FIXED_BBOX 0 0 96 96
string GDS_END 12233040
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 12232204
<< end >>
