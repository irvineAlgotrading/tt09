magic
tech sky130B
timestamp 1704896540
<< viali >>
rect 0 0 53 305
<< metal1 >>
rect -6 305 59 308
rect -6 0 0 305
rect 53 0 59 305
rect -6 -3 59 0
<< properties >>
string GDS_END 87999354
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87998070
<< end >>
