magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 131 0 160
rect -50 97 -34 131
rect -50 63 0 97
rect -50 29 -34 63
rect -50 0 0 29
rect -50 -637 0 -608
rect -50 -671 -34 -637
rect -50 -705 0 -671
rect -50 -739 -34 -705
rect -50 -768 0 -739
<< polycont >>
rect -34 97 0 131
rect -34 29 0 63
rect -34 -671 0 -637
rect -34 -739 0 -705
<< npolyres >>
rect 0 0 2523 160
rect 2363 -96 2523 0
rect -50 -256 2523 -96
rect -50 -352 110 -256
rect -50 -512 2523 -352
rect 2363 -608 2523 -512
rect 0 -768 2523 -608
<< locali >>
rect -34 131 0 147
rect -34 63 0 97
rect -34 13 0 29
rect -34 -637 0 -621
rect -34 -705 0 -671
rect -34 -755 0 -739
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 1 0 -50 0 1 -755
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 1 0 -50 0 1 13
box 0 0 1 1
<< properties >>
string GDS_END 90831050
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90829798
<< end >>
