magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 219 366
<< mvpmos >>
rect 0 0 100 300
<< mvpdiff >>
rect -50 0 0 300
rect 100 0 150 300
<< poly >>
rect 0 300 100 326
rect 0 -26 100 0
<< metal1 >>
rect -51 -16 -5 258
rect 105 -16 151 258
use DFM1sd_CDNS_524688791851302  DFM1sd_CDNS_524688791851302_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 336
use DFM1sd_CDNS_524688791851302  DFM1sd_CDNS_524688791851302_1
timestamp 1704896540
transform 1 0 100 0 1 0
box -36 -36 89 336
<< labels >>
flabel comment s -28 121 -28 121 0 FreeSans 300 0 0 0 S
flabel comment s 128 121 128 121 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86358660
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86357642
<< end >>
