magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< metal2 >>
rect 0 785 216 794
rect 0 0 216 9
<< via2 >>
rect 0 9 216 785
<< metal3 >>
rect -5 785 221 790
rect -5 9 0 785
rect 216 9 221 785
rect -5 4 221 9
<< properties >>
string GDS_END 98012434
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98010382
<< end >>
