magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 314
rect 253 0 256 314
<< via1 >>
rect 3 0 253 314
<< metal2 >>
rect 0 0 3 314
rect 253 0 256 314
<< properties >>
string GDS_END 88444466
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88439214
<< end >>
